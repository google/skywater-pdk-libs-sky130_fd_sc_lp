* File: sky130_fd_sc_lp__o211a_4.spice
* Created: Fri Aug 28 11:02:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o211a_4.pex.spice"
.subckt sky130_fd_sc_lp__o211a_4  VNB VPB B1 C1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1011 N_X_M1011_d N_A_80_21#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1014 N_X_M1011_d N_A_80_21#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1015 N_X_M1015_d N_A_80_21#_M1015_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1023 N_X_M1015_d N_A_80_21#_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_475_49#_M1004_d N_B1_M1004_g N_A_574_49#_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2898 AS=0.1176 PD=2.37 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6
+ SA=75000.3 SB=75003.5 A=0.126 P=1.98 MULT=1
MM1016 N_A_80_21#_M1016_d N_C1_M1016_g N_A_574_49#_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.21365 AS=0.1176 PD=1.44 PS=1.12 NRD=14.28 NRS=0 M=1 R=5.6
+ SA=75000.7 SB=75003.1 A=0.126 P=1.98 MULT=1
MM1020 N_A_80_21#_M1016_d N_C1_M1020_g N_A_574_49#_M1020_s VNB NSHORT L=0.15
+ W=0.84 AD=0.21365 AS=0.1176 PD=1.44 PS=1.12 NRD=14.28 NRS=0 M=1 R=5.6
+ SA=75001.3 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1008 N_A_475_49#_M1008_d N_B1_M1008_g N_A_574_49#_M1020_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6
+ SA=75001.7 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A1_M1001_g N_A_475_49#_M1008_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1344 PD=1.23 PS=1.16 NRD=5.712 NRS=0 M=1 R=5.6 SA=75002.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1006 N_A_475_49#_M1006_d N_A2_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1638 PD=1.12 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.8
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1018 N_A_475_49#_M1006_d N_A2_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1018_s N_A1_M1003_g N_A_475_49#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_80_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.5 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_80_21#_M1009_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6 SB=75005
+ A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1009_d N_A_80_21#_M1012_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.6 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1021_d N_A_80_21#_M1021_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75004.2 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1021_d N_B1_M1005_g N_A_80_21#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4284 PD=1.54 PS=1.94 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_C1_M1010_g N_A_80_21#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4284 PD=1.54 PS=1.94 NRD=0 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1010_d N_C1_M1022_g N_A_80_21#_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2457 PD=1.54 PS=1.65 NRD=0 NRS=10.9335 M=1 R=8.4 SA=75003.2
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_B1_M1017_g N_A_80_21#_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.2457 PD=1.58 PS=1.65 NRD=0 NRS=6.2449 M=1 R=8.4 SA=75003.7
+ SB=75002 A=0.189 P=2.82 MULT=1
MM1000 N_A_986_367#_M1000_d N_A1_M1000_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=6.2449 M=1 R=8.4
+ SA=75004.2 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1007 N_A_986_367#_M1000_d N_A2_M1007_g N_A_80_21#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1013 N_A_986_367#_M1013_d N_A2_M1013_g N_A_80_21#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1019 N_A_986_367#_M1013_d N_A1_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75005.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.2415 P=17.93
*
.include "sky130_fd_sc_lp__o211a_4.pxi.spice"
*
.ends
*
*
