# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.385000 1.775000 2.130000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.195000 0.365000 10.465000 3.075000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.495000 2.735000 1.795000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.145000 1.285000 1.475000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.255000 1.175000 3.695000 2.215000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.245000 10.560000 3.415000 ;
      RECT 0.095000  0.635000  0.620000 0.965000 ;
      RECT 0.095000  0.965000  0.265000 1.655000 ;
      RECT 0.095000  1.655000  1.235000 1.985000 ;
      RECT 0.450000  1.985000  1.235000 2.300000 ;
      RECT 0.450000  2.300000  2.235000 2.470000 ;
      RECT 0.450000  2.470000  0.780000 3.045000 ;
      RECT 0.840000  0.085000  1.050000 0.925000 ;
      RECT 0.950000  2.640000  1.245000 3.245000 ;
      RECT 1.750000  2.640000  2.585000 2.970000 ;
      RECT 1.945000  0.685000  2.195000 1.155000 ;
      RECT 1.945000  1.155000  3.075000 1.325000 ;
      RECT 1.995000  1.965000  2.235000 2.300000 ;
      RECT 2.415000  2.035000  3.075000 2.205000 ;
      RECT 2.415000  2.205000  2.725000 2.490000 ;
      RECT 2.415000  2.490000  2.585000 2.640000 ;
      RECT 2.655000  0.085000  2.945000 0.935000 ;
      RECT 2.755000  2.660000  2.945000 3.245000 ;
      RECT 2.905000  1.325000  3.075000 2.035000 ;
      RECT 3.115000  0.715000  4.235000 0.985000 ;
      RECT 3.115000  2.385000  4.235000 2.555000 ;
      RECT 3.115000  2.555000  3.445000 3.045000 ;
      RECT 3.635000  2.725000  3.895000 3.245000 ;
      RECT 3.660000  0.085000  3.920000 0.545000 ;
      RECT 3.865000  0.985000  4.235000 2.385000 ;
      RECT 4.065000  2.555000  4.235000 2.895000 ;
      RECT 4.065000  2.895000  5.930000 3.065000 ;
      RECT 4.090000  0.265000  5.850000 0.485000 ;
      RECT 4.405000  0.485000  4.595000 2.725000 ;
      RECT 4.765000  0.665000  5.095000 0.995000 ;
      RECT 4.765000  0.995000  4.935000 2.225000 ;
      RECT 4.765000  2.225000  5.170000 2.555000 ;
      RECT 5.115000  1.175000  6.820000 1.345000 ;
      RECT 5.115000  1.345000  5.285000 1.875000 ;
      RECT 5.115000  1.875000  5.590000 2.045000 ;
      RECT 5.265000  0.655000  5.510000 1.175000 ;
      RECT 5.340000  2.045000  5.590000 2.615000 ;
      RECT 5.465000  1.515000  5.930000 1.705000 ;
      RECT 5.680000  0.485000  5.850000 0.815000 ;
      RECT 5.680000  0.815000  6.905000 0.985000 ;
      RECT 5.760000  1.705000  5.930000 2.635000 ;
      RECT 5.760000  2.635000  7.520000 2.805000 ;
      RECT 5.760000  2.805000  5.930000 2.895000 ;
      RECT 6.100000  1.685000  7.170000 2.465000 ;
      RECT 6.225000  0.085000  6.555000 0.635000 ;
      RECT 6.330000  2.975000  6.660000 3.245000 ;
      RECT 6.650000  1.345000  6.820000 1.505000 ;
      RECT 6.735000  0.385000  7.765000 0.555000 ;
      RECT 6.735000  0.555000  6.905000 0.815000 ;
      RECT 7.000000  1.165000  7.265000 1.335000 ;
      RECT 7.000000  1.335000  7.170000 1.685000 ;
      RECT 7.075000  0.735000  7.265000 1.165000 ;
      RECT 7.350000  1.755000  7.605000 2.085000 ;
      RECT 7.350000  2.085000  7.520000 2.635000 ;
      RECT 7.435000  0.555000  7.765000 1.125000 ;
      RECT 7.435000  1.295000  8.250000 1.465000 ;
      RECT 7.435000  1.465000  7.605000 1.755000 ;
      RECT 7.690000  2.515000  7.955000 2.845000 ;
      RECT 7.785000  1.645000  9.220000 1.815000 ;
      RECT 7.785000  1.815000  7.955000 2.515000 ;
      RECT 7.945000  0.345000  8.590000 0.675000 ;
      RECT 7.990000  0.855000  8.250000 1.295000 ;
      RECT 8.285000  1.985000  9.570000 2.175000 ;
      RECT 8.420000  0.675000  8.590000 1.305000 ;
      RECT 8.420000  1.305000  9.220000 1.645000 ;
      RECT 8.755000  2.345000  9.085000 3.245000 ;
      RECT 8.810000  0.085000  9.020000 0.975000 ;
      RECT 9.240000  0.315000  9.570000 0.985000 ;
      RECT 9.265000  2.175000  9.570000 2.910000 ;
      RECT 9.400000  0.985000  9.570000 1.415000 ;
      RECT 9.400000  1.415000  9.780000 1.645000 ;
      RECT 9.400000  1.645000  9.570000 1.985000 ;
      RECT 9.740000  0.085000 10.025000 1.245000 ;
      RECT 9.740000  1.815000  9.975000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  2.320000  2.725000 2.490000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  2.320000  5.125000 2.490000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
    LAYER met1 ;
      RECT 2.495000 2.290000 2.785000 2.335000 ;
      RECT 2.495000 2.335000 5.185000 2.475000 ;
      RECT 2.495000 2.475000 2.785000 2.520000 ;
      RECT 4.895000 2.290000 5.185000 2.335000 ;
      RECT 4.895000 2.475000 5.185000 2.520000 ;
  END
END sky130_fd_sc_lp__sdfxtp_1
END LIBRARY
