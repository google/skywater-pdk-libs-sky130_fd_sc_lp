* File: sky130_fd_sc_lp__or4b_4.pex.spice
* Created: Fri Aug 28 11:25:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4B_4%A_83_21# 1 2 3 12 16 20 24 28 32 36 40 42 51
+ 52 53 56 58 62 66 68 72 73 75 82
c128 75 0 3.41083e-19 $X=3.972 $Y=1.815
c129 51 0 5.1554e-20 $X=1.82 $Y=1.355
r130 79 80 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.92 $Y=1.44
+ $X2=1.35 $Y2=1.44
r131 73 74 19.6322 $w=1.74e-07 $l=2.8e-07 $layer=LI1_cond $X=3.665 $Y=1.085
+ $X2=3.945 $Y2=1.085
r132 68 70 45.6073 $w=2.33e-07 $l=9.3e-07 $layer=LI1_cond $X=3.972 $Y=1.98
+ $X2=3.972 $Y2=2.91
r133 66 75 6.39787 $w=2.33e-07 $l=1.17e-07 $layer=LI1_cond $X=3.972 $Y=1.932
+ $X2=3.972 $Y2=1.815
r134 66 68 2.35393 $w=2.33e-07 $l=4.8e-08 $layer=LI1_cond $X=3.972 $Y=1.932
+ $X2=3.972 $Y2=1.98
r135 64 74 0.508694 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=3.945 $Y=1.175
+ $X2=3.945 $Y2=1.085
r136 64 75 39.4343 $w=1.78e-07 $l=6.4e-07 $layer=LI1_cond $X=3.945 $Y=1.175
+ $X2=3.945 $Y2=1.815
r137 60 73 0.172717 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=3.665 $Y=0.995
+ $X2=3.665 $Y2=1.085
r138 60 62 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=3.665 $Y=0.995
+ $X2=3.665 $Y2=0.42
r139 59 72 5.86152 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=2.56 $Y=1.085
+ $X2=2.455 $Y2=1.085
r140 58 73 6.43889 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.57 $Y=1.085
+ $X2=3.665 $Y2=1.085
r141 58 59 62.2323 $w=1.78e-07 $l=1.01e-06 $layer=LI1_cond $X=3.57 $Y=1.085
+ $X2=2.56 $Y2=1.085
r142 54 72 0.793806 $w=2.1e-07 $l=9e-08 $layer=LI1_cond $X=2.455 $Y=0.995
+ $X2=2.455 $Y2=1.085
r143 54 56 30.368 $w=2.08e-07 $l=5.75e-07 $layer=LI1_cond $X=2.455 $Y=0.995
+ $X2=2.455 $Y2=0.42
r144 52 72 5.86152 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=2.35 $Y=1.085
+ $X2=2.455 $Y2=1.085
r145 52 53 27.4192 $w=1.78e-07 $l=4.45e-07 $layer=LI1_cond $X=2.35 $Y=1.085
+ $X2=1.905 $Y2=1.085
r146 50 53 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.82 $Y=1.175
+ $X2=1.905 $Y2=1.085
r147 50 51 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.82 $Y=1.175
+ $X2=1.82 $Y2=1.355
r148 49 82 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.69 $Y=1.44 $X2=1.78
+ $Y2=1.44
r149 49 80 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.69 $Y=1.44
+ $X2=1.35 $Y2=1.44
r150 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.44 $X2=1.69 $Y2=1.44
r151 45 79 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.67 $Y=1.44
+ $X2=0.92 $Y2=1.44
r152 45 76 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.67 $Y=1.44
+ $X2=0.49 $Y2=1.44
r153 44 48 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.67 $Y=1.44
+ $X2=1.69 $Y2=1.44
r154 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.67
+ $Y=1.44 $X2=0.67 $Y2=1.44
r155 42 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.735 $Y=1.44
+ $X2=1.82 $Y2=1.355
r156 42 48 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.735 $Y=1.44
+ $X2=1.69 $Y2=1.44
r157 38 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.605
+ $X2=1.78 $Y2=1.44
r158 38 40 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.78 $Y=1.605
+ $X2=1.78 $Y2=2.465
r159 34 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.275
+ $X2=1.78 $Y2=1.44
r160 34 36 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.78 $Y=1.275
+ $X2=1.78 $Y2=0.655
r161 30 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.605
+ $X2=1.35 $Y2=1.44
r162 30 32 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.35 $Y=1.605
+ $X2=1.35 $Y2=2.465
r163 26 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.275
+ $X2=1.35 $Y2=1.44
r164 26 28 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.35 $Y=1.275
+ $X2=1.35 $Y2=0.655
r165 22 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.605
+ $X2=0.92 $Y2=1.44
r166 22 24 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.92 $Y=1.605
+ $X2=0.92 $Y2=2.465
r167 18 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.275
+ $X2=0.92 $Y2=1.44
r168 18 20 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.92 $Y=1.275
+ $X2=0.92 $Y2=0.655
r169 14 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.605
+ $X2=0.49 $Y2=1.44
r170 14 16 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.49 $Y=1.605
+ $X2=0.49 $Y2=2.465
r171 10 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.275
+ $X2=0.49 $Y2=1.44
r172 10 12 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.49 $Y=1.275
+ $X2=0.49 $Y2=0.655
r173 3 70 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.835
+ $Y=1.835 $X2=3.975 $Y2=2.91
r174 3 68 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.835
+ $Y=1.835 $X2=3.975 $Y2=1.98
r175 2 62 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.525
+ $Y=0.235 $X2=3.665 $Y2=0.42
r176 1 56 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.235 $X2=2.465 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_4%A 3 7 9 12 13
c38 12 0 5.1554e-20 $X=2.23 $Y=1.51
r39 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.51
+ $X2=2.23 $Y2=1.675
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.51
+ $X2=2.23 $Y2=1.345
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.51 $X2=2.23 $Y2=1.51
r42 9 13 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=1.51
r43 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.32 $Y=2.465
+ $X2=2.32 $Y2=1.675
r44 3 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.25 $Y=0.655
+ $X2=2.25 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_4%B 3 7 9 10 11 12 18 19
r41 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.51
+ $X2=2.77 $Y2=1.675
r42 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.51
+ $X2=2.77 $Y2=1.345
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.51 $X2=2.77 $Y2=1.51
r44 11 12 9.41594 $w=4.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.405
+ $X2=2.62 $Y2=2.775
r45 11 27 6.36212 $w=4.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.62 $Y=2.405
+ $X2=2.62 $Y2=2.155
r46 10 27 3.05382 $w=4.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.62 $Y=2.035
+ $X2=2.62 $Y2=2.155
r47 10 34 3.5012 $w=4.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.62 $Y=2.035
+ $X2=2.62 $Y2=1.92
r48 9 34 7.94251 $w=3.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.67 $Y=1.665
+ $X2=2.67 $Y2=1.92
r49 9 19 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.67 $Y=1.665
+ $X2=2.67 $Y2=1.51
r50 7 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.68 $Y=2.465
+ $X2=2.68 $Y2=1.675
r51 3 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.68 $Y=0.655
+ $X2=2.68 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_4%C 1 3 5 7 8 9 10 11 26
c36 3 0 7.92674e-20 $X=3.22 $Y=2.465
r37 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.31
+ $Y=1.43 $X2=3.31 $Y2=1.43
r38 10 11 6.70529 $w=6.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.355 $Y=2.405
+ $X2=3.355 $Y2=2.775
r39 9 10 6.70529 $w=6.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.355 $Y=2.035
+ $X2=3.355 $Y2=2.405
r40 8 9 6.70529 $w=6.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.355 $Y=1.665
+ $X2=3.355 $Y2=2.035
r41 8 26 4.25876 $w=6.58e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=1.665
+ $X2=3.355 $Y2=1.43
r42 5 25 49.8417 $w=3.48e-07 $l=2.96985e-07 $layer=POLY_cond $X=3.45 $Y=1.185
+ $X2=3.335 $Y2=1.43
r43 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.45 $Y=1.185 $X2=3.45
+ $Y2=0.655
r44 1 25 38.7612 $w=3.48e-07 $l=2.14942e-07 $layer=POLY_cond $X=3.22 $Y=1.595
+ $X2=3.335 $Y2=1.43
r45 1 3 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=3.22 $Y=1.595 $X2=3.22
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_4%A_737_315# 1 2 7 9 10 12 14 15 17 18 21 25 27
+ 34
c61 34 0 1.81959e-19 $X=3.88 $Y=1.455
r62 31 34 42.175 $w=4.8e-07 $l=4.2e-07 $layer=POLY_cond $X=4.3 $Y=1.455 $X2=3.88
+ $Y2=1.455
r63 30 32 5.73858 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=4.387 $Y=1.35
+ $X2=4.387 $Y2=1.515
r64 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.3
+ $Y=1.35 $X2=4.3 $Y2=1.35
r65 27 30 2.67233 $w=3.43e-07 $l=8e-08 $layer=LI1_cond $X=4.387 $Y=1.27
+ $X2=4.387 $Y2=1.35
r66 23 25 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=5.055 $Y=2.545
+ $X2=5.055 $Y2=2.835
r67 19 21 14.1839 $w=2.58e-07 $l=3.2e-07 $layer=LI1_cond $X=5 $Y=1.185 $X2=5
+ $Y2=0.865
r68 17 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.925 $Y=2.46
+ $X2=5.055 $Y2=2.545
r69 17 18 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.925 $Y=2.46
+ $X2=4.56 $Y2=2.46
r70 16 27 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.56 $Y=1.27
+ $X2=4.387 $Y2=1.27
r71 15 19 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.87 $Y=1.27
+ $X2=5 $Y2=1.185
r72 15 16 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.87 $Y=1.27
+ $X2=4.56 $Y2=1.27
r73 14 18 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=4.41 $Y=2.375
+ $X2=4.56 $Y2=2.46
r74 14 32 33.0367 $w=2.98e-07 $l=8.6e-07 $layer=LI1_cond $X=4.41 $Y=2.375
+ $X2=4.41 $Y2=1.515
r75 10 34 30.3798 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.88 $Y=1.185
+ $X2=3.88 $Y2=1.455
r76 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.88 $Y=1.185
+ $X2=3.88 $Y2=0.655
r77 7 34 12.05 $w=4.8e-07 $l=3.245e-07 $layer=POLY_cond $X=3.76 $Y=1.725
+ $X2=3.88 $Y2=1.455
r78 7 9 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.76 $Y=1.725 $X2=3.76
+ $Y2=2.465
r79 2 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=2.625 $X2=5.02 $Y2=2.835
r80 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.655 $X2=4.965 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_4%D_N 3 7 11 13 14 15 19
c33 14 0 1.81959e-19 $X=5.04 $Y=1.665
c34 3 0 1.30707e-19 $X=4.75 $Y=0.865
r35 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.895
+ $Y=1.7 $X2=4.895 $Y2=1.7
r36 15 20 8.61691 $w=4.63e-07 $l=3.35e-07 $layer=LI1_cond $X=4.962 $Y=2.035
+ $X2=4.962 $Y2=1.7
r37 14 20 0.900274 $w=4.63e-07 $l=3.5e-08 $layer=LI1_cond $X=4.962 $Y=1.665
+ $X2=4.962 $Y2=1.7
r38 12 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.895 $Y=2.04
+ $X2=4.895 $Y2=1.7
r39 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.895 $Y=2.04
+ $X2=4.895 $Y2=2.205
r40 11 19 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.895 $Y=1.685
+ $X2=4.895 $Y2=1.7
r41 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.867 $Y=1.535
+ $X2=4.867 $Y2=1.685
r42 7 13 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=4.805 $Y=2.835
+ $X2=4.805 $Y2=2.205
r43 3 10 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=4.75 $Y=0.865
+ $X2=4.75 $Y2=1.535
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_4%VPWR 1 2 3 4 13 15 21 27 33 35 37 42 47 54 55
+ 61 64 67
r74 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r77 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r78 55 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r79 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r80 52 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=3.33
+ $X2=4.59 $Y2=3.33
r81 52 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.755 $Y=3.33
+ $X2=5.04 $Y2=3.33
r82 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r83 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r84 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.05 $Y2=3.33
r85 48 50 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 47 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.59 $Y2=3.33
r87 47 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 46 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r89 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r90 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 43 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.135 $Y2=3.33
r92 43 45 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=1.68
+ $Y2=3.33
r93 42 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=2.05 $Y2=3.33
r94 42 45 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.68 $Y2=3.33
r95 41 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r96 41 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r97 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 38 58 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r99 38 40 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 37 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.135 $Y2=3.33
r101 37 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 35 51 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r103 35 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 31 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=3.245
+ $X2=4.59 $Y2=3.33
r105 31 33 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=4.59 $Y=3.245
+ $X2=4.59 $Y2=2.84
r106 27 30 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=2.05 $Y=2.005
+ $X2=2.05 $Y2=2.95
r107 25 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=3.245
+ $X2=2.05 $Y2=3.33
r108 25 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.05 $Y=3.245
+ $X2=2.05 $Y2=2.95
r109 21 24 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.135 $Y=2.12
+ $X2=1.135 $Y2=2.95
r110 19 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=3.33
r111 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=2.95
r112 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.275 $Y=2.12
+ $X2=0.275 $Y2=2.95
r113 13 58 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r114 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.95
r115 4 33 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=4.465
+ $Y=2.625 $X2=4.59 $Y2=2.84
r116 3 30 400 $w=1.7e-07 $l=1.20857e-06 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=2.05 $Y2=2.95
r117 3 27 400 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=2.05 $Y2=2.005
r118 2 24 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.95
r119 2 21 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.12
r120 1 18 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.95
r121 1 15 400 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_4%X 1 2 3 4 13 14 15 19 27 31 33 37 43 45 49 50
+ 54 59
r59 54 59 1.41115 $w=2.43e-07 $l=3e-08 $layer=LI1_cond $X=0.212 $Y=1.695
+ $X2=0.212 $Y2=1.665
r60 50 54 2.90557 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.212 $Y=1.78
+ $X2=0.212 $Y2=1.695
r61 50 59 1.31708 $w=2.43e-07 $l=2.8e-08 $layer=LI1_cond $X=0.212 $Y=1.637
+ $X2=0.212 $Y2=1.665
r62 49 50 16.0872 $w=2.43e-07 $l=3.42e-07 $layer=LI1_cond $X=0.212 $Y=1.295
+ $X2=0.212 $Y2=1.637
r63 45 47 4.75325 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=1.575 $Y=0.65
+ $X2=1.575 $Y2=0.74
r64 41 49 5.64462 $w=2.43e-07 $l=1.2e-07 $layer=LI1_cond $X=0.212 $Y=1.175
+ $X2=0.212 $Y2=1.295
r65 37 39 43.7458 $w=2.43e-07 $l=9.3e-07 $layer=LI1_cond $X=1.592 $Y=1.98
+ $X2=1.592 $Y2=2.91
r66 35 37 5.40943 $w=2.43e-07 $l=1.15e-07 $layer=LI1_cond $X=1.592 $Y=1.865
+ $X2=1.592 $Y2=1.98
r67 34 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.8 $Y=1.78 $X2=0.705
+ $Y2=1.78
r68 33 35 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=1.47 $Y=1.78
+ $X2=1.592 $Y2=1.865
r69 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.47 $Y=1.78 $X2=0.8
+ $Y2=1.78
r70 32 42 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.8 $Y=0.74 $X2=0.705
+ $Y2=0.74
r71 31 47 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.47 $Y=0.74
+ $X2=1.575 $Y2=0.74
r72 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.47 $Y=0.74 $X2=0.8
+ $Y2=0.74
r73 27 29 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.705 $Y=1.98
+ $X2=0.705 $Y2=2.91
r74 25 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.865
+ $X2=0.705 $Y2=1.78
r75 25 27 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=0.705 $Y=1.865
+ $X2=0.705 $Y2=1.98
r76 22 24 4.62121 $w=1.78e-07 $l=7.5e-08 $layer=LI1_cond $X=0.7 $Y=1.005 $X2=0.7
+ $Y2=0.93
r77 21 42 4.81226 $w=1.85e-07 $l=8.74643e-08 $layer=LI1_cond $X=0.7 $Y=0.825
+ $X2=0.705 $Y2=0.74
r78 21 24 6.4697 $w=1.78e-07 $l=1.05e-07 $layer=LI1_cond $X=0.7 $Y=0.825 $X2=0.7
+ $Y2=0.93
r79 17 42 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.655
+ $X2=0.705 $Y2=0.74
r80 17 19 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=0.705 $Y=0.655
+ $X2=0.705 $Y2=0.42
r81 16 50 4.20453 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.335 $Y=1.78
+ $X2=0.212 $Y2=1.78
r82 15 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.61 $Y=1.78
+ $X2=0.705 $Y2=1.78
r83 15 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.61 $Y=1.78
+ $X2=0.335 $Y2=1.78
r84 14 41 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.335 $Y=1.09
+ $X2=0.212 $Y2=1.175
r85 13 22 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.61 $Y=1.09
+ $X2=0.7 $Y2=1.005
r86 13 14 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.61 $Y=1.09
+ $X2=0.335 $Y2=1.09
r87 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=2.91
r88 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=1.98
r89 3 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.91
r90 3 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=1.98
r91 2 45 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=1.425
+ $Y=0.235 $X2=1.565 $Y2=0.65
r92 1 24 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.705 $Y2=0.93
r93 1 19 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.705 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_4%VGND 1 2 3 4 5 16 18 22 26 30 33 34 35 37 46
+ 50 57 58 64 67 75
r83 75 77 8.83448 $w=7.25e-07 $l=5.25e-07 $layer=LI1_cond $X=4.315 $Y=0.38
+ $X2=4.315 $Y2=0.905
r84 71 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r85 70 75 6.39448 $w=7.25e-07 $l=3.8e-07 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.315
+ $Y2=0.38
r86 70 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r87 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r88 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r89 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r90 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r91 58 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r92 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r93 55 70 9.55322 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=4.7 $Y=0 $X2=4.315
+ $Y2=0
r94 55 57 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.7 $Y=0 $X2=5.04
+ $Y2=0
r95 54 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r96 54 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r97 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r98 51 67 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.065
+ $Y2=0
r99 51 53 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.6 $Y2=0
r100 50 70 9.55322 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=3.93 $Y=0 $X2=4.315
+ $Y2=0
r101 50 53 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.93 $Y=0 $X2=3.6
+ $Y2=0
r102 46 67 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.73 $Y=0 $X2=3.065
+ $Y2=0
r103 46 48 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.73 $Y=0 $X2=2.64
+ $Y2=0
r104 45 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r105 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r106 42 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.135
+ $Y2=0
r107 42 44 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.68
+ $Y2=0
r108 41 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r109 41 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r110 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r111 38 61 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r112 38 40 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.72
+ $Y2=0
r113 37 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.135
+ $Y2=0
r114 37 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.72
+ $Y2=0
r115 35 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r116 35 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r117 35 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r118 33 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.68
+ $Y2=0
r119 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.015
+ $Y2=0
r120 32 48 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.64
+ $Y2=0
r121 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.015
+ $Y2=0
r122 28 67 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.065 $Y2=0
r123 28 30 4.90928 $w=6.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.065 $Y2=0.36
r124 24 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0
r125 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0.36
r126 20 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0
r127 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0.36
r128 16 61 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r129 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.38
r130 5 77 182 $w=1.7e-07 $l=9.1515e-07 $layer=licon1_NDIFF $count=1 $X=3.955
+ $Y=0.235 $X2=4.535 $Y2=0.905
r131 5 75 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.955
+ $Y=0.235 $X2=4.095 $Y2=0.38
r132 4 30 45.5 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=4 $X=2.755
+ $Y=0.235 $X2=3.235 $Y2=0.36
r133 3 26 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=1.855
+ $Y=0.235 $X2=2.015 $Y2=0.36
r134 2 22 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.235 $X2=1.135 $Y2=0.36
r135 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.38
.ends

