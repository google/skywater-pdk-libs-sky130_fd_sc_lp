* File: sky130_fd_sc_lp__a221oi_4.pxi.spice
* Created: Fri Aug 28 09:53:32 2020
* 
x_PM_SKY130_FD_SC_LP__A221OI_4%C1 N_C1_M1016_g N_C1_c_144_n N_C1_M1007_g
+ N_C1_M1022_g N_C1_c_146_n N_C1_M1025_g N_C1_M1031_g N_C1_c_148_n N_C1_M1028_g
+ N_C1_M1037_g N_C1_c_150_n N_C1_M1036_g C1 C1 C1 C1 C1 N_C1_c_152_n
+ N_C1_c_153_n PM_SKY130_FD_SC_LP__A221OI_4%C1
x_PM_SKY130_FD_SC_LP__A221OI_4%B2 N_B2_M1001_g N_B2_M1004_g N_B2_M1002_g
+ N_B2_M1008_g N_B2_M1021_g N_B2_M1023_g N_B2_M1032_g N_B2_M1034_g N_B2_c_287_p
+ N_B2_c_262_p N_B2_c_242_n N_B2_c_254_p N_B2_c_294_p B2 N_B2_c_235_n
+ N_B2_c_236_n N_B2_c_237_n B2 PM_SKY130_FD_SC_LP__A221OI_4%B2
x_PM_SKY130_FD_SC_LP__A221OI_4%B1 N_B1_M1006_g N_B1_M1003_g N_B1_M1012_g
+ N_B1_M1011_g N_B1_M1026_g N_B1_M1030_g N_B1_M1027_g N_B1_M1035_g B1 B1 B1 B1
+ N_B1_c_371_n PM_SKY130_FD_SC_LP__A221OI_4%B1
x_PM_SKY130_FD_SC_LP__A221OI_4%A2 N_A2_M1005_g N_A2_M1013_g N_A2_c_441_n
+ N_A2_M1015_g N_A2_M1014_g N_A2_c_443_n N_A2_M1018_g N_A2_M1019_g N_A2_c_445_n
+ N_A2_M1029_g N_A2_M1033_g N_A2_c_447_n N_A2_c_448_n N_A2_c_449_n N_A2_c_450_n
+ N_A2_c_451_n A2 A2 A2 A2 N_A2_c_453_n PM_SKY130_FD_SC_LP__A221OI_4%A2
x_PM_SKY130_FD_SC_LP__A221OI_4%A1 N_A1_c_565_n N_A1_M1000_g N_A1_M1009_g
+ N_A1_c_567_n N_A1_M1017_g N_A1_M1010_g N_A1_c_569_n N_A1_M1020_g N_A1_c_577_n
+ N_A1_M1024_g N_A1_c_570_n N_A1_c_571_n N_A1_c_572_n N_A1_M1039_g N_A1_c_579_n
+ N_A1_M1038_g A1 A1 A1 N_A1_c_574_n PM_SKY130_FD_SC_LP__A221OI_4%A1
x_PM_SKY130_FD_SC_LP__A221OI_4%A_85_367# N_A_85_367#_M1016_s N_A_85_367#_M1022_s
+ N_A_85_367#_M1037_s N_A_85_367#_M1004_s N_A_85_367#_M1023_s
+ N_A_85_367#_M1011_s N_A_85_367#_M1035_s N_A_85_367#_c_650_n
+ N_A_85_367#_c_651_n N_A_85_367#_c_659_n N_A_85_367#_c_691_p
+ N_A_85_367#_c_661_n N_A_85_367#_c_652_n N_A_85_367#_c_653_n
+ N_A_85_367#_c_654_n N_A_85_367#_c_706_p N_A_85_367#_c_671_n
+ N_A_85_367#_c_714_p N_A_85_367#_c_655_n PM_SKY130_FD_SC_LP__A221OI_4%A_85_367#
x_PM_SKY130_FD_SC_LP__A221OI_4%Y N_Y_M1007_s N_Y_M1028_s N_Y_M1006_s N_Y_M1026_s
+ N_Y_M1000_s N_Y_M1020_s N_Y_M1016_d N_Y_M1031_d N_Y_c_739_n N_Y_c_843_p
+ N_Y_c_727_n N_Y_c_728_n N_Y_c_750_n N_Y_c_754_n N_Y_c_756_n N_Y_c_844_p
+ N_Y_c_729_n N_Y_c_762_n N_Y_c_730_n N_Y_c_731_n N_Y_c_732_n N_Y_c_808_n
+ N_Y_c_809_n N_Y_c_733_n N_Y_c_771_n N_Y_c_734_n N_Y_c_793_n Y Y Y Y
+ N_Y_c_735_n N_Y_c_736_n PM_SKY130_FD_SC_LP__A221OI_4%Y
x_PM_SKY130_FD_SC_LP__A221OI_4%A_533_367# N_A_533_367#_M1004_d
+ N_A_533_367#_M1008_d N_A_533_367#_M1003_d N_A_533_367#_M1030_d
+ N_A_533_367#_M1032_d N_A_533_367#_M1009_d N_A_533_367#_M1024_d
+ N_A_533_367#_M1014_d N_A_533_367#_M1033_d N_A_533_367#_c_877_n
+ N_A_533_367#_c_888_n N_A_533_367#_c_878_n N_A_533_367#_c_894_n
+ N_A_533_367#_c_961_p N_A_533_367#_c_896_n N_A_533_367#_c_903_n
+ N_A_533_367#_c_897_n N_A_533_367#_c_962_p N_A_533_367#_c_909_n
+ N_A_533_367#_c_956_p N_A_533_367#_c_910_n N_A_533_367#_c_879_n
+ N_A_533_367#_c_963_p N_A_533_367#_c_875_n N_A_533_367#_c_876_n
+ N_A_533_367#_c_881_n N_A_533_367#_c_927_n N_A_533_367#_c_928_n
+ N_A_533_367#_c_929_n PM_SKY130_FD_SC_LP__A221OI_4%A_533_367#
x_PM_SKY130_FD_SC_LP__A221OI_4%VPWR N_VPWR_M1005_s N_VPWR_M1010_s N_VPWR_M1038_s
+ N_VPWR_M1019_s N_VPWR_c_982_n N_VPWR_c_983_n N_VPWR_c_984_n N_VPWR_c_985_n
+ N_VPWR_c_986_n N_VPWR_c_987_n N_VPWR_c_988_n N_VPWR_c_989_n N_VPWR_c_990_n
+ VPWR N_VPWR_c_991_n N_VPWR_c_992_n N_VPWR_c_981_n N_VPWR_c_994_n
+ N_VPWR_c_995_n PM_SKY130_FD_SC_LP__A221OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A221OI_4%VGND N_VGND_M1007_d N_VGND_M1025_d N_VGND_M1036_d
+ N_VGND_M1002_s N_VGND_M1034_s N_VGND_M1015_d N_VGND_M1029_d N_VGND_c_1100_n
+ N_VGND_c_1101_n N_VGND_c_1102_n N_VGND_c_1103_n N_VGND_c_1104_n
+ N_VGND_c_1105_n N_VGND_c_1106_n N_VGND_c_1107_n N_VGND_c_1108_n
+ N_VGND_c_1109_n N_VGND_c_1110_n N_VGND_c_1111_n N_VGND_c_1112_n
+ N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n VGND N_VGND_c_1116_n
+ N_VGND_c_1117_n N_VGND_c_1118_n N_VGND_c_1119_n N_VGND_c_1120_n
+ N_VGND_c_1121_n PM_SKY130_FD_SC_LP__A221OI_4%VGND
x_PM_SKY130_FD_SC_LP__A221OI_4%A_546_47# N_A_546_47#_M1001_d N_A_546_47#_M1021_d
+ N_A_546_47#_M1012_d N_A_546_47#_M1027_d N_A_546_47#_c_1237_n
+ N_A_546_47#_c_1239_n N_A_546_47#_c_1255_n N_A_546_47#_c_1243_n
+ PM_SKY130_FD_SC_LP__A221OI_4%A_546_47#
x_PM_SKY130_FD_SC_LP__A221OI_4%A_1334_47# N_A_1334_47#_M1013_s
+ N_A_1334_47#_M1017_d N_A_1334_47#_M1039_d N_A_1334_47#_M1018_s
+ N_A_1334_47#_c_1273_n N_A_1334_47#_c_1297_n N_A_1334_47#_c_1274_n
+ N_A_1334_47#_c_1277_n N_A_1334_47#_c_1301_n
+ PM_SKY130_FD_SC_LP__A221OI_4%A_1334_47#
cc_1 VNB N_C1_M1016_g 0.0109769f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=2.465
cc_2 VNB N_C1_c_144_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.185
cc_3 VNB N_C1_M1022_g 0.00665511f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=2.465
cc_4 VNB N_C1_c_146_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.185
cc_5 VNB N_C1_M1031_g 0.00665511f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=2.465
cc_6 VNB N_C1_c_148_n 0.0160037f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.185
cc_7 VNB N_C1_M1037_g 0.00754919f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=2.465
cc_8 VNB N_C1_c_150_n 0.0161688f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.185
cc_9 VNB C1 0.0190386f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_10 VNB N_C1_c_152_n 0.0659072f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.35
cc_11 VNB N_C1_c_153_n 0.0868839f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.35
cc_12 VNB N_B2_M1001_g 0.0222432f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=2.465
cc_13 VNB N_B2_M1002_g 0.0225787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B2_M1021_g 0.0261986f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.185
cc_15 VNB N_B2_M1034_g 0.028209f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_16 VNB N_B2_c_235_n 0.0683684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B2_c_236_n 0.0248393f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.322
cc_18 VNB N_B2_c_237_n 0.00435502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_M1006_g 0.0271034f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=2.465
cc_20 VNB N_B1_M1012_g 0.0233885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_M1026_g 0.0233885f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.185
cc_22 VNB N_B1_M1027_g 0.0256501f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.655
cc_23 VNB B1 0.00652666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_c_371_n 0.0649774f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=1.35
cc_25 VNB N_A2_M1013_g 0.0264901f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.655
cc_26 VNB N_A2_c_441_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=2.465
cc_27 VNB N_A2_M1014_g 0.00727234f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.655
cc_28 VNB N_A2_c_443_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=2.465
cc_29 VNB N_A2_M1019_g 0.00665779f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.655
cc_30 VNB N_A2_c_445_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=2.465
cc_31 VNB N_A2_M1033_g 0.0100771f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.655
cc_32 VNB N_A2_c_447_n 0.00739997f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_33 VNB N_A2_c_448_n 0.00285936f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_34 VNB N_A2_c_449_n 0.00549961f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_35 VNB N_A2_c_450_n 0.0012932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A2_c_451_n 0.0258995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB A2 0.0132101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A2_c_453_n 0.0921595f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.322
cc_39 VNB N_A1_c_565_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.515
cc_40 VNB N_A1_M1009_g 0.00650355f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.655
cc_41 VNB N_A1_c_567_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.515
cc_42 VNB N_A1_M1010_g 0.00674291f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.655
cc_43 VNB N_A1_c_569_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.515
cc_44 VNB N_A1_c_570_n 0.0163505f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.655
cc_45 VNB N_A1_c_571_n 0.0107967f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=2.465
cc_46 VNB N_A1_c_572_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB A1 0.00582647f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_48 VNB N_A1_c_574_n 0.0556033f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.35
cc_49 VNB N_Y_c_727_n 0.00223696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_Y_c_728_n 0.00228659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_Y_c_729_n 0.00302899f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.35
cc_52 VNB N_Y_c_730_n 0.00280369f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.35
cc_53 VNB N_Y_c_731_n 0.00710553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_Y_c_732_n 0.0020833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_Y_c_733_n 0.00228659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Y_c_734_n 0.00177903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Y_c_735_n 0.00638811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Y_c_736_n 0.0068064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_533_367#_c_875_n 0.00678475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_533_367#_c_876_n 0.00186209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VPWR_c_981_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1100_n 0.0338983f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=2.465
cc_63 VNB N_VGND_c_1101_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.655
cc_64 VNB N_VGND_c_1102_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_65 VNB N_VGND_c_1103_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1104_n 0.002833f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.35
cc_67 VNB N_VGND_c_1105_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.35
cc_68 VNB N_VGND_c_1106_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.35
cc_69 VNB N_VGND_c_1107_n 0.034011f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.35
cc_70 VNB N_VGND_c_1108_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=1.35
cc_71 VNB N_VGND_c_1109_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=1.35
cc_72 VNB N_VGND_c_1110_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.35
cc_73 VNB N_VGND_c_1111_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1112_n 0.0129195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1113_n 0.0043639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1114_n 0.0597532f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.322
cc_77 VNB N_VGND_c_1115_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1116_n 0.0198045f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.322
cc_79 VNB N_VGND_c_1117_n 0.0538181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1118_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1119_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1120_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1121_n 0.486338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VPB N_C1_M1016_g 0.0264961f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=2.465
cc_85 VPB N_C1_M1022_g 0.0185149f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=2.465
cc_86 VPB N_C1_M1031_g 0.0185149f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=2.465
cc_87 VPB N_C1_M1037_g 0.0246251f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=2.465
cc_88 VPB N_B2_M1004_g 0.0236566f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.655
cc_89 VPB N_B2_M1008_g 0.0186926f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=1.515
cc_90 VPB N_B2_M1023_g 0.0183617f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=2.465
cc_91 VPB N_B2_M1032_g 0.019617f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=0.655
cc_92 VPB N_B2_c_242_n 0.00142004f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.35
cc_93 VPB B2 0.00127504f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=1.35
cc_94 VPB N_B2_c_235_n 0.0187599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_B2_c_236_n 0.00634987f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.322
cc_96 VPB N_B2_c_237_n 0.00284809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_B1_M1003_g 0.0182364f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.655
cc_98 VPB N_B1_M1011_g 0.0180542f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=1.515
cc_99 VPB N_B1_M1030_g 0.018053f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=2.465
cc_100 VPB N_B1_M1035_g 0.0182238f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_101 VPB B1 0.0114892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_B1_c_371_n 0.014175f $X=-0.19 $Y=1.655 $X2=2.09 $Y2=1.35
cc_103 VPB N_A2_M1005_g 0.0194847f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=2.465
cc_104 VPB N_A2_M1014_g 0.0191179f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=0.655
cc_105 VPB N_A2_M1019_g 0.0185652f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=0.655
cc_106 VPB N_A2_M1033_g 0.0232847f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=0.655
cc_107 VPB N_A2_c_447_n 0.0124445f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_108 VPB N_A2_c_450_n 0.00203732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A2_c_451_n 0.00632332f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A1_M1009_g 0.0189179f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.655
cc_111 VPB N_A1_M1010_g 0.0185384f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=0.655
cc_112 VPB N_A1_c_577_n 0.0155213f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A1_c_571_n 0.00697523f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=2.465
cc_114 VPB N_A1_c_579_n 0.0156118f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=0.655
cc_115 VPB N_A1_c_574_n 0.00204448f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=1.35
cc_116 VPB N_A_85_367#_c_650_n 0.00746637f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=1.515
cc_117 VPB N_A_85_367#_c_651_n 0.0435127f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=2.465
cc_118 VPB N_A_85_367#_c_652_n 6.27129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_85_367#_c_653_n 0.00985145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_85_367#_c_654_n 0.0102866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_85_367#_c_655_n 0.00230215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_Y_c_727_n 0.00488423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_Y_c_729_n 0.0074522f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=1.35
cc_124 VPB N_A_533_367#_c_877_n 0.00462239f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_125 VPB N_A_533_367#_c_878_n 0.0030329f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_126 VPB N_A_533_367#_c_879_n 4.98048e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_533_367#_c_875_n 0.0110324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_533_367#_c_881_n 0.0498589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_982_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=1.625 $Y2=1.515
cc_130 VPB N_VPWR_c_983_n 3.12649e-19 $X=-0.19 $Y=1.655 $X2=1.795 $Y2=1.185
cc_131 VPB N_VPWR_c_984_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=0.655
cc_132 VPB N_VPWR_c_985_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_986_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_134 VPB N_VPWR_c_987_n 0.155096f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_988_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_989_n 0.0134822f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_990_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_991_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=1.35
cc_139 VPB N_VPWR_c_992_n 0.0153631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_981_n 0.0665856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_994_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_995_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.322
cc_143 N_C1_c_150_n N_B2_M1001_g 0.0225415f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_144 C1 N_B2_M1001_g 2.10368e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_145 N_C1_M1037_g N_B2_c_235_n 0.00354542f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_146 N_C1_c_153_n N_B2_c_235_n 0.0225415f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_147 N_C1_M1016_g N_A_85_367#_c_651_n 0.00335189f $X=0.765 $Y=2.465 $X2=0
+ $Y2=0
cc_148 C1 N_A_85_367#_c_651_n 0.0116679f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_149 N_C1_c_152_n N_A_85_367#_c_651_n 0.00581571f $X=0.69 $Y=1.35 $X2=0 $Y2=0
cc_150 N_C1_M1016_g N_A_85_367#_c_659_n 0.0115031f $X=0.765 $Y=2.465 $X2=0 $Y2=0
cc_151 N_C1_M1022_g N_A_85_367#_c_659_n 0.0115031f $X=1.195 $Y=2.465 $X2=0 $Y2=0
cc_152 N_C1_M1031_g N_A_85_367#_c_661_n 0.0115031f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_153 N_C1_M1037_g N_A_85_367#_c_661_n 0.0115031f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_154 N_C1_M1016_g N_Y_c_739_n 0.0125173f $X=0.765 $Y=2.465 $X2=0 $Y2=0
cc_155 N_C1_M1022_g N_Y_c_739_n 0.0119581f $X=1.195 $Y=2.465 $X2=0 $Y2=0
cc_156 N_C1_M1031_g N_Y_c_739_n 6.58347e-19 $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_157 N_C1_M1022_g N_Y_c_727_n 0.01115f $X=1.195 $Y=2.465 $X2=0 $Y2=0
cc_158 N_C1_M1031_g N_Y_c_727_n 0.01115f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_159 C1 N_Y_c_727_n 0.0376973f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_160 N_C1_c_153_n N_Y_c_727_n 0.00289453f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_161 N_C1_M1016_g N_Y_c_728_n 0.0104117f $X=0.765 $Y=2.465 $X2=0 $Y2=0
cc_162 N_C1_M1022_g N_Y_c_728_n 0.00279308f $X=1.195 $Y=2.465 $X2=0 $Y2=0
cc_163 C1 N_Y_c_728_n 0.0268977f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_164 N_C1_c_153_n N_Y_c_728_n 0.00299787f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_165 N_C1_c_146_n N_Y_c_750_n 0.0122595f $X=1.365 $Y=1.185 $X2=0 $Y2=0
cc_166 N_C1_c_148_n N_Y_c_750_n 0.0122129f $X=1.795 $Y=1.185 $X2=0 $Y2=0
cc_167 C1 N_Y_c_750_n 0.039834f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_168 N_C1_c_153_n N_Y_c_750_n 0.00271364f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_169 C1 N_Y_c_754_n 0.0142048f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_170 N_C1_c_153_n N_Y_c_754_n 0.00280606f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_171 N_C1_M1022_g N_Y_c_756_n 6.58347e-19 $X=1.195 $Y=2.465 $X2=0 $Y2=0
cc_172 N_C1_M1031_g N_Y_c_756_n 0.0119581f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_173 N_C1_M1037_g N_Y_c_756_n 0.0167624f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_174 N_C1_M1037_g N_Y_c_729_n 0.0125165f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_175 C1 N_Y_c_729_n 0.0184815f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_176 N_C1_c_153_n N_Y_c_729_n 0.00508426f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_177 N_C1_c_150_n N_Y_c_762_n 0.0125637f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_178 C1 N_Y_c_762_n 0.00952471f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_179 N_C1_M1037_g N_Y_c_730_n 0.00173663f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_180 C1 N_Y_c_730_n 0.0144348f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_181 N_C1_c_153_n N_Y_c_730_n 0.00327775f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_182 N_C1_M1031_g N_Y_c_733_n 0.00279308f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_183 N_C1_M1037_g N_Y_c_733_n 0.00279308f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_184 C1 N_Y_c_733_n 0.0268977f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_185 N_C1_c_153_n N_Y_c_733_n 0.00299787f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_186 C1 N_Y_c_771_n 0.0142048f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_187 N_C1_c_153_n N_Y_c_771_n 0.00280606f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_188 N_C1_c_150_n N_Y_c_734_n 0.00531522f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_189 C1 N_Y_c_734_n 0.00392261f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_190 N_C1_M1016_g N_VPWR_c_987_n 0.00357877f $X=0.765 $Y=2.465 $X2=0 $Y2=0
cc_191 N_C1_M1022_g N_VPWR_c_987_n 0.00357877f $X=1.195 $Y=2.465 $X2=0 $Y2=0
cc_192 N_C1_M1031_g N_VPWR_c_987_n 0.00357877f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_193 N_C1_M1037_g N_VPWR_c_987_n 0.00357877f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_194 N_C1_M1016_g N_VPWR_c_981_n 0.00646653f $X=0.765 $Y=2.465 $X2=0 $Y2=0
cc_195 N_C1_M1022_g N_VPWR_c_981_n 0.00541285f $X=1.195 $Y=2.465 $X2=0 $Y2=0
cc_196 N_C1_M1031_g N_VPWR_c_981_n 0.00541285f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_197 N_C1_M1037_g N_VPWR_c_981_n 0.00665089f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_198 N_C1_c_144_n N_VGND_c_1100_n 0.0165374f $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_199 N_C1_c_146_n N_VGND_c_1100_n 6.24191e-19 $X=1.365 $Y=1.185 $X2=0 $Y2=0
cc_200 C1 N_VGND_c_1100_n 0.0237475f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_201 N_C1_c_152_n N_VGND_c_1100_n 0.00778396f $X=0.69 $Y=1.35 $X2=0 $Y2=0
cc_202 N_C1_c_144_n N_VGND_c_1101_n 5.75816e-19 $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_203 N_C1_c_146_n N_VGND_c_1101_n 0.0105703f $X=1.365 $Y=1.185 $X2=0 $Y2=0
cc_204 N_C1_c_148_n N_VGND_c_1101_n 0.0105703f $X=1.795 $Y=1.185 $X2=0 $Y2=0
cc_205 N_C1_c_150_n N_VGND_c_1101_n 5.75816e-19 $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_206 N_C1_c_148_n N_VGND_c_1102_n 5.75816e-19 $X=1.795 $Y=1.185 $X2=0 $Y2=0
cc_207 N_C1_c_150_n N_VGND_c_1102_n 0.0104941f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_208 N_C1_c_144_n N_VGND_c_1108_n 0.00486043f $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_209 N_C1_c_146_n N_VGND_c_1108_n 0.00486043f $X=1.365 $Y=1.185 $X2=0 $Y2=0
cc_210 N_C1_c_148_n N_VGND_c_1110_n 0.00486043f $X=1.795 $Y=1.185 $X2=0 $Y2=0
cc_211 N_C1_c_150_n N_VGND_c_1110_n 0.00486043f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_212 N_C1_c_144_n N_VGND_c_1121_n 0.00824727f $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_213 N_C1_c_146_n N_VGND_c_1121_n 0.00824727f $X=1.365 $Y=1.185 $X2=0 $Y2=0
cc_214 N_C1_c_148_n N_VGND_c_1121_n 0.00824727f $X=1.795 $Y=1.185 $X2=0 $Y2=0
cc_215 N_C1_c_150_n N_VGND_c_1121_n 0.00824727f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_216 N_B2_M1021_g N_B1_M1006_g 0.0177659f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_217 N_B2_M1023_g N_B1_M1003_g 0.054301f $X=3.865 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B2_c_242_n N_B1_M1003_g 9.0036e-19 $X=3.73 $Y=1.93 $X2=0 $Y2=0
cc_219 N_B2_c_254_p N_B1_M1003_g 0.010446f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_220 N_B2_c_254_p N_B1_M1011_g 0.0104926f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_221 N_B2_c_254_p N_B1_M1030_g 0.0104926f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_222 N_B2_M1034_g N_B1_M1027_g 0.0296173f $X=6.085 $Y=0.655 $X2=0 $Y2=0
cc_223 N_B2_M1032_g N_B1_M1035_g 0.0527509f $X=6.015 $Y=2.465 $X2=0 $Y2=0
cc_224 N_B2_c_254_p N_B1_M1035_g 0.010446f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_225 B2 N_B1_M1035_g 0.00402468f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_226 N_B2_M1032_g B1 2.72953e-19 $X=6.015 $Y=2.465 $X2=0 $Y2=0
cc_227 N_B2_c_262_p B1 0.0178283f $X=3.73 $Y=1.625 $X2=0 $Y2=0
cc_228 N_B2_c_242_n B1 0.0107418f $X=3.73 $Y=1.93 $X2=0 $Y2=0
cc_229 N_B2_c_254_p B1 0.114702f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_230 N_B2_c_235_n B1 0.00510205f $X=3.865 $Y=1.51 $X2=0 $Y2=0
cc_231 N_B2_c_236_n B1 0.00118708f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_232 N_B2_c_237_n B1 0.035542f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_233 N_B2_c_254_p N_B1_c_371_n 0.00196281f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_234 N_B2_c_235_n N_B1_c_371_n 0.0218533f $X=3.865 $Y=1.51 $X2=0 $Y2=0
cc_235 N_B2_c_236_n N_B1_c_371_n 0.0179851f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_236 N_B2_c_237_n N_B1_c_371_n 0.00109469f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_237 N_B2_M1032_g N_A2_M1005_g 0.03315f $X=6.015 $Y=2.465 $X2=0 $Y2=0
cc_238 B2 N_A2_M1005_g 9.50204e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_239 N_B2_M1034_g N_A2_M1013_g 0.0349269f $X=6.085 $Y=0.655 $X2=0 $Y2=0
cc_240 N_B2_M1032_g N_A2_c_450_n 7.33524e-19 $X=6.015 $Y=2.465 $X2=0 $Y2=0
cc_241 B2 N_A2_c_450_n 0.00511231f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_242 N_B2_c_236_n N_A2_c_450_n 0.00115083f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_243 N_B2_c_237_n N_A2_c_450_n 0.0205723f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_244 N_B2_c_236_n N_A2_c_451_n 0.0201104f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_245 N_B2_c_237_n N_A2_c_451_n 0.00114905f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_246 N_B2_c_254_p N_A_85_367#_M1023_s 0.0035116f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_247 N_B2_c_254_p N_A_85_367#_M1011_s 0.00333608f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_248 N_B2_c_254_p N_A_85_367#_M1035_s 0.00679813f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_249 B2 N_A_85_367#_M1035_s 0.00114953f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_250 N_B2_M1004_g N_A_85_367#_c_653_n 0.00447454f $X=3.005 $Y=2.465 $X2=0
+ $Y2=0
cc_251 N_B2_M1004_g N_A_85_367#_c_654_n 0.0125958f $X=3.005 $Y=2.465 $X2=0 $Y2=0
cc_252 N_B2_c_287_p N_A_85_367#_c_654_n 0.00933996f $X=3.645 $Y=1.525 $X2=0
+ $Y2=0
cc_253 N_B2_c_235_n N_A_85_367#_c_654_n 0.00921295f $X=3.865 $Y=1.51 $X2=0 $Y2=0
cc_254 N_B2_M1008_g N_A_85_367#_c_671_n 0.0149596f $X=3.435 $Y=2.465 $X2=0 $Y2=0
cc_255 N_B2_M1023_g N_A_85_367#_c_671_n 0.0125991f $X=3.865 $Y=2.465 $X2=0 $Y2=0
cc_256 N_B2_M1032_g N_A_85_367#_c_671_n 0.00406236f $X=6.015 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_B2_c_287_p N_A_85_367#_c_671_n 0.00664216f $X=3.645 $Y=1.525 $X2=0
+ $Y2=0
cc_258 N_B2_c_254_p N_A_85_367#_c_671_n 0.117148f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_259 N_B2_c_294_p N_A_85_367#_c_671_n 0.00939762f $X=3.815 $Y=2.015 $X2=0
+ $Y2=0
cc_260 N_B2_c_235_n N_A_85_367#_c_671_n 9.44648e-19 $X=3.865 $Y=1.51 $X2=0 $Y2=0
cc_261 N_B2_M1004_g N_A_85_367#_c_655_n 0.00868052f $X=3.005 $Y=2.465 $X2=0
+ $Y2=0
cc_262 N_B2_M1008_g N_A_85_367#_c_655_n 7.69038e-19 $X=3.435 $Y=2.465 $X2=0
+ $Y2=0
cc_263 N_B2_c_287_p N_A_85_367#_c_655_n 0.0214139f $X=3.645 $Y=1.525 $X2=0 $Y2=0
cc_264 N_B2_c_242_n N_A_85_367#_c_655_n 0.00412561f $X=3.73 $Y=1.93 $X2=0 $Y2=0
cc_265 N_B2_c_235_n N_A_85_367#_c_655_n 0.00280798f $X=3.865 $Y=1.51 $X2=0 $Y2=0
cc_266 N_B2_M1004_g N_Y_c_729_n 0.00358178f $X=3.005 $Y=2.465 $X2=0 $Y2=0
cc_267 N_B2_c_287_p N_Y_c_729_n 0.00160837f $X=3.645 $Y=1.525 $X2=0 $Y2=0
cc_268 N_B2_c_235_n N_Y_c_729_n 0.00536343f $X=3.865 $Y=1.51 $X2=0 $Y2=0
cc_269 N_B2_M1001_g N_Y_c_730_n 0.00237569f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_270 N_B2_M1002_g N_Y_c_730_n 4.59734e-19 $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_271 N_B2_c_287_p N_Y_c_730_n 0.0137548f $X=3.645 $Y=1.525 $X2=0 $Y2=0
cc_272 N_B2_c_235_n N_Y_c_730_n 0.00959614f $X=3.865 $Y=1.51 $X2=0 $Y2=0
cc_273 N_B2_M1001_g N_Y_c_731_n 0.0132965f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_274 N_B2_M1002_g N_Y_c_731_n 0.0131372f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_275 N_B2_M1021_g N_Y_c_731_n 0.0144966f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_276 N_B2_c_287_p N_Y_c_731_n 0.0612922f $X=3.645 $Y=1.525 $X2=0 $Y2=0
cc_277 N_B2_c_262_p N_Y_c_731_n 0.00405481f $X=3.73 $Y=1.625 $X2=0 $Y2=0
cc_278 N_B2_c_235_n N_Y_c_731_n 0.00796581f $X=3.865 $Y=1.51 $X2=0 $Y2=0
cc_279 N_B2_M1034_g N_Y_c_732_n 0.00253831f $X=6.085 $Y=0.655 $X2=0 $Y2=0
cc_280 N_B2_c_236_n N_Y_c_732_n 5.80146e-19 $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_281 N_B2_c_237_n N_Y_c_732_n 0.00556632f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_282 N_B2_M1001_g N_Y_c_734_n 0.00958029f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_283 N_B2_M1002_g N_Y_c_734_n 7.0069e-19 $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_284 N_B2_M1034_g N_Y_c_793_n 0.0135731f $X=6.085 $Y=0.655 $X2=0 $Y2=0
cc_285 N_B2_c_237_n N_Y_c_793_n 0.0088351f $X=6.035 $Y=1.51 $X2=0 $Y2=0
cc_286 N_B2_M1021_g N_Y_c_736_n 0.00393366f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_287 N_B2_c_262_p N_Y_c_736_n 0.00987737f $X=3.73 $Y=1.625 $X2=0 $Y2=0
cc_288 N_B2_c_235_n N_Y_c_736_n 0.00873501f $X=3.865 $Y=1.51 $X2=0 $Y2=0
cc_289 N_B2_c_242_n N_A_533_367#_M1008_d 0.00100696f $X=3.73 $Y=1.93 $X2=0 $Y2=0
cc_290 N_B2_c_294_p N_A_533_367#_M1008_d 0.00286639f $X=3.815 $Y=2.015 $X2=0
+ $Y2=0
cc_291 N_B2_c_254_p N_A_533_367#_M1003_d 0.00333608f $X=5.85 $Y=2.015 $X2=0
+ $Y2=0
cc_292 N_B2_c_254_p N_A_533_367#_M1030_d 0.00333608f $X=5.85 $Y=2.015 $X2=0
+ $Y2=0
cc_293 N_B2_M1004_g N_A_533_367#_c_877_n 0.00922548f $X=3.005 $Y=2.465 $X2=0
+ $Y2=0
cc_294 N_B2_M1008_g N_A_533_367#_c_877_n 7.61713e-19 $X=3.435 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_B2_M1004_g N_A_533_367#_c_888_n 0.0118334f $X=3.005 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_B2_M1008_g N_A_533_367#_c_888_n 0.0112455f $X=3.435 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_B2_M1023_g N_A_533_367#_c_888_n 0.0111475f $X=3.865 $Y=2.465 $X2=0
+ $Y2=0
cc_298 N_B2_M1032_g N_A_533_367#_c_888_n 0.0174506f $X=6.015 $Y=2.465 $X2=0
+ $Y2=0
cc_299 N_B2_c_254_p N_A_533_367#_c_888_n 0.0030166f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_300 N_B2_M1004_g N_A_533_367#_c_878_n 8.94866e-19 $X=3.005 $Y=2.465 $X2=0
+ $Y2=0
cc_301 N_B2_c_236_n N_A_533_367#_c_894_n 3.49628e-19 $X=6.035 $Y=1.51 $X2=0
+ $Y2=0
cc_302 N_B2_c_237_n N_A_533_367#_c_894_n 0.00175636f $X=6.035 $Y=1.51 $X2=0
+ $Y2=0
cc_303 N_B2_M1032_g N_A_533_367#_c_896_n 0.00325588f $X=6.015 $Y=2.465 $X2=0
+ $Y2=0
cc_304 N_B2_M1032_g N_A_533_367#_c_897_n 0.00183621f $X=6.015 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_B2_c_254_p N_A_533_367#_c_897_n 0.0126736f $X=5.85 $Y=2.015 $X2=0 $Y2=0
cc_306 N_B2_M1032_g N_VPWR_c_982_n 0.00124613f $X=6.015 $Y=2.465 $X2=0 $Y2=0
cc_307 N_B2_M1004_g N_VPWR_c_987_n 0.00357842f $X=3.005 $Y=2.465 $X2=0 $Y2=0
cc_308 N_B2_M1008_g N_VPWR_c_987_n 0.00357877f $X=3.435 $Y=2.465 $X2=0 $Y2=0
cc_309 N_B2_M1023_g N_VPWR_c_987_n 0.00357877f $X=3.865 $Y=2.465 $X2=0 $Y2=0
cc_310 N_B2_M1032_g N_VPWR_c_987_n 0.00357877f $X=6.015 $Y=2.465 $X2=0 $Y2=0
cc_311 N_B2_M1004_g N_VPWR_c_981_n 0.00665087f $X=3.005 $Y=2.465 $X2=0 $Y2=0
cc_312 N_B2_M1008_g N_VPWR_c_981_n 0.0053512f $X=3.435 $Y=2.465 $X2=0 $Y2=0
cc_313 N_B2_M1023_g N_VPWR_c_981_n 0.00537849f $X=3.865 $Y=2.465 $X2=0 $Y2=0
cc_314 N_B2_M1032_g N_VPWR_c_981_n 0.00575852f $X=6.015 $Y=2.465 $X2=0 $Y2=0
cc_315 N_B2_M1001_g N_VGND_c_1102_n 0.0123289f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_316 N_B2_M1002_g N_VGND_c_1102_n 0.00120563f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_317 N_B2_M1001_g N_VGND_c_1103_n 0.00115725f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_318 N_B2_M1002_g N_VGND_c_1103_n 0.00867619f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_319 N_B2_M1021_g N_VGND_c_1103_n 0.00815384f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_320 N_B2_M1034_g N_VGND_c_1104_n 0.0128677f $X=6.085 $Y=0.655 $X2=0 $Y2=0
cc_321 N_B2_M1001_g N_VGND_c_1112_n 0.00486043f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_322 N_B2_M1002_g N_VGND_c_1112_n 0.00358332f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_323 N_B2_M1021_g N_VGND_c_1114_n 0.00358332f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_324 N_B2_M1034_g N_VGND_c_1114_n 0.00486043f $X=6.085 $Y=0.655 $X2=0 $Y2=0
cc_325 N_B2_M1001_g N_VGND_c_1121_n 0.00835506f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_326 N_B2_M1002_g N_VGND_c_1121_n 0.00427377f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_327 N_B2_M1021_g N_VGND_c_1121_n 0.00475663f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_328 N_B2_M1034_g N_VGND_c_1121_n 0.00484087f $X=6.085 $Y=0.655 $X2=0 $Y2=0
cc_329 N_B2_M1002_g N_A_546_47#_c_1237_n 0.00965692f $X=3.085 $Y=0.655 $X2=0
+ $Y2=0
cc_330 N_B2_M1021_g N_A_546_47#_c_1237_n 0.0112968f $X=3.515 $Y=0.655 $X2=0
+ $Y2=0
cc_331 N_B1_M1003_g N_A_85_367#_c_671_n 0.0127052f $X=4.295 $Y=2.465 $X2=0 $Y2=0
cc_332 N_B1_M1011_g N_A_85_367#_c_671_n 0.0127052f $X=4.725 $Y=2.465 $X2=0 $Y2=0
cc_333 N_B1_M1030_g N_A_85_367#_c_671_n 0.0127052f $X=5.155 $Y=2.465 $X2=0 $Y2=0
cc_334 N_B1_M1035_g N_A_85_367#_c_671_n 0.0127052f $X=5.585 $Y=2.465 $X2=0 $Y2=0
cc_335 N_B1_M1027_g N_Y_c_732_n 0.0167399f $X=5.515 $Y=0.655 $X2=0 $Y2=0
cc_336 B1 N_Y_c_732_n 0.0200139f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_337 N_B1_c_371_n N_Y_c_732_n 2.31066e-19 $X=5.515 $Y=1.51 $X2=0 $Y2=0
cc_338 N_B1_M1006_g N_Y_c_735_n 0.00805022f $X=4.225 $Y=0.655 $X2=0 $Y2=0
cc_339 N_B1_M1012_g N_Y_c_735_n 0.0166676f $X=4.655 $Y=0.655 $X2=0 $Y2=0
cc_340 N_B1_M1026_g N_Y_c_735_n 0.0166377f $X=5.085 $Y=0.655 $X2=0 $Y2=0
cc_341 B1 N_Y_c_735_n 0.0958482f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_342 N_B1_c_371_n N_Y_c_735_n 0.00780147f $X=5.515 $Y=1.51 $X2=0 $Y2=0
cc_343 N_B1_M1006_g N_Y_c_736_n 0.0116544f $X=4.225 $Y=0.655 $X2=0 $Y2=0
cc_344 B1 N_Y_c_736_n 0.0182099f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_345 N_B1_M1003_g N_A_533_367#_c_888_n 0.0111616f $X=4.295 $Y=2.465 $X2=0
+ $Y2=0
cc_346 N_B1_M1011_g N_A_533_367#_c_888_n 0.0112455f $X=4.725 $Y=2.465 $X2=0
+ $Y2=0
cc_347 N_B1_M1030_g N_A_533_367#_c_888_n 0.0112455f $X=5.155 $Y=2.465 $X2=0
+ $Y2=0
cc_348 N_B1_M1035_g N_A_533_367#_c_888_n 0.0111616f $X=5.585 $Y=2.465 $X2=0
+ $Y2=0
cc_349 N_B1_M1003_g N_VPWR_c_987_n 0.00357877f $X=4.295 $Y=2.465 $X2=0 $Y2=0
cc_350 N_B1_M1011_g N_VPWR_c_987_n 0.00357877f $X=4.725 $Y=2.465 $X2=0 $Y2=0
cc_351 N_B1_M1030_g N_VPWR_c_987_n 0.00357877f $X=5.155 $Y=2.465 $X2=0 $Y2=0
cc_352 N_B1_M1035_g N_VPWR_c_987_n 0.00357877f $X=5.585 $Y=2.465 $X2=0 $Y2=0
cc_353 N_B1_M1003_g N_VPWR_c_981_n 0.00537849f $X=4.295 $Y=2.465 $X2=0 $Y2=0
cc_354 N_B1_M1011_g N_VPWR_c_981_n 0.0053512f $X=4.725 $Y=2.465 $X2=0 $Y2=0
cc_355 N_B1_M1030_g N_VPWR_c_981_n 0.0053512f $X=5.155 $Y=2.465 $X2=0 $Y2=0
cc_356 N_B1_M1035_g N_VPWR_c_981_n 0.00537849f $X=5.585 $Y=2.465 $X2=0 $Y2=0
cc_357 N_B1_M1006_g N_VGND_c_1103_n 7.74631e-19 $X=4.225 $Y=0.655 $X2=0 $Y2=0
cc_358 N_B1_M1027_g N_VGND_c_1104_n 0.00164616f $X=5.515 $Y=0.655 $X2=0 $Y2=0
cc_359 N_B1_M1006_g N_VGND_c_1114_n 0.00357877f $X=4.225 $Y=0.655 $X2=0 $Y2=0
cc_360 N_B1_M1012_g N_VGND_c_1114_n 0.00357877f $X=4.655 $Y=0.655 $X2=0 $Y2=0
cc_361 N_B1_M1026_g N_VGND_c_1114_n 0.00357877f $X=5.085 $Y=0.655 $X2=0 $Y2=0
cc_362 N_B1_M1027_g N_VGND_c_1114_n 0.00357877f $X=5.515 $Y=0.655 $X2=0 $Y2=0
cc_363 N_B1_M1006_g N_VGND_c_1121_n 0.00602315f $X=4.225 $Y=0.655 $X2=0 $Y2=0
cc_364 N_B1_M1012_g N_VGND_c_1121_n 0.0053512f $X=4.655 $Y=0.655 $X2=0 $Y2=0
cc_365 N_B1_M1026_g N_VGND_c_1121_n 0.0053512f $X=5.085 $Y=0.655 $X2=0 $Y2=0
cc_366 N_B1_M1027_g N_VGND_c_1121_n 0.00577254f $X=5.515 $Y=0.655 $X2=0 $Y2=0
cc_367 N_B1_M1006_g N_A_546_47#_c_1239_n 0.0171609f $X=4.225 $Y=0.655 $X2=0
+ $Y2=0
cc_368 N_B1_M1012_g N_A_546_47#_c_1239_n 0.0119021f $X=4.655 $Y=0.655 $X2=0
+ $Y2=0
cc_369 N_B1_M1026_g N_A_546_47#_c_1239_n 0.0119021f $X=5.085 $Y=0.655 $X2=0
+ $Y2=0
cc_370 N_B1_M1027_g N_A_546_47#_c_1239_n 0.0166096f $X=5.515 $Y=0.655 $X2=0
+ $Y2=0
cc_371 N_B1_M1006_g N_A_546_47#_c_1243_n 0.00385562f $X=4.225 $Y=0.655 $X2=0
+ $Y2=0
cc_372 N_A2_M1013_g N_A1_c_565_n 0.0419856f $X=6.595 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_373 N_A2_M1005_g N_A1_M1009_g 0.0333392f $X=6.565 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A2_c_447_n N_A1_M1009_g 0.0102122f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_375 N_A2_c_447_n N_A1_M1010_g 0.0105539f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_376 N_A2_c_447_n N_A1_c_577_n 0.00424188f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_377 N_A2_c_447_n N_A1_c_570_n 8.13109e-19 $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_378 N_A2_c_448_n N_A1_c_570_n 0.0131912f $X=8.365 $Y=1.435 $X2=0 $Y2=0
cc_379 N_A2_c_453_n N_A1_c_570_n 0.0102387f $X=9.785 $Y=1.35 $X2=0 $Y2=0
cc_380 N_A2_M1014_g N_A1_c_571_n 0.0403844f $X=8.745 $Y=2.465 $X2=0 $Y2=0
cc_381 N_A2_c_447_n N_A1_c_571_n 0.00945338f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_382 N_A2_c_449_n N_A1_c_571_n 0.00392986f $X=8.365 $Y=1.615 $X2=0 $Y2=0
cc_383 N_A2_c_441_n N_A1_c_572_n 0.0146005f $X=8.745 $Y=1.185 $X2=0 $Y2=0
cc_384 N_A2_c_447_n N_A1_c_579_n 0.0039366f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_385 N_A2_M1013_g A1 0.00400963f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_386 N_A2_c_447_n A1 0.0861325f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_387 N_A2_c_448_n A1 0.0198573f $X=8.365 $Y=1.435 $X2=0 $Y2=0
cc_388 N_A2_c_450_n A1 0.00736506f $X=6.575 $Y=1.51 $X2=0 $Y2=0
cc_389 N_A2_c_451_n A1 6.4198e-19 $X=6.575 $Y=1.51 $X2=0 $Y2=0
cc_390 N_A2_c_453_n A1 4.49811e-19 $X=9.785 $Y=1.35 $X2=0 $Y2=0
cc_391 N_A2_c_447_n N_A1_c_574_n 0.00985409f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_392 N_A2_c_449_n N_A1_c_574_n 0.00120228f $X=8.365 $Y=1.615 $X2=0 $Y2=0
cc_393 N_A2_c_450_n N_A1_c_574_n 0.00115456f $X=6.575 $Y=1.51 $X2=0 $Y2=0
cc_394 N_A2_c_451_n N_A1_c_574_n 0.0217495f $X=6.575 $Y=1.51 $X2=0 $Y2=0
cc_395 N_A2_c_453_n N_A1_c_574_n 7.8558e-19 $X=9.785 $Y=1.35 $X2=0 $Y2=0
cc_396 N_A2_M1013_g N_Y_c_808_n 7.68343e-19 $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_397 N_A2_c_448_n N_Y_c_809_n 7.52138e-19 $X=8.365 $Y=1.435 $X2=0 $Y2=0
cc_398 N_A2_M1013_g N_Y_c_793_n 0.0131906f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_399 N_A2_c_447_n N_Y_c_793_n 0.00784112f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_400 N_A2_c_450_n N_Y_c_793_n 0.0100412f $X=6.575 $Y=1.51 $X2=0 $Y2=0
cc_401 N_A2_c_451_n N_Y_c_793_n 0.00178367f $X=6.575 $Y=1.51 $X2=0 $Y2=0
cc_402 N_A2_M1005_g N_A_533_367#_c_903_n 0.0126836f $X=6.565 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A2_c_447_n N_A_533_367#_c_903_n 0.0294876f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_404 N_A2_c_450_n N_A_533_367#_c_903_n 0.0133469f $X=6.575 $Y=1.51 $X2=0 $Y2=0
cc_405 N_A2_c_451_n N_A_533_367#_c_903_n 3.60177e-19 $X=6.575 $Y=1.51 $X2=0
+ $Y2=0
cc_406 N_A2_c_450_n N_A_533_367#_c_897_n 0.00292251f $X=6.575 $Y=1.51 $X2=0
+ $Y2=0
cc_407 N_A2_c_451_n N_A_533_367#_c_897_n 2.10792e-19 $X=6.575 $Y=1.51 $X2=0
+ $Y2=0
cc_408 N_A2_c_447_n N_A_533_367#_c_909_n 0.0402256f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_409 N_A2_M1014_g N_A_533_367#_c_910_n 0.0118088f $X=8.745 $Y=2.465 $X2=0
+ $Y2=0
cc_410 N_A2_c_447_n N_A_533_367#_c_910_n 0.0185646f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_411 A2 N_A_533_367#_c_910_n 0.00854407f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_412 N_A2_c_453_n N_A_533_367#_c_910_n 0.00111203f $X=9.785 $Y=1.35 $X2=0
+ $Y2=0
cc_413 N_A2_M1014_g N_A_533_367#_c_879_n 0.00367383f $X=8.745 $Y=2.465 $X2=0
+ $Y2=0
cc_414 N_A2_M1019_g N_A_533_367#_c_879_n 8.32811e-19 $X=9.175 $Y=2.465 $X2=0
+ $Y2=0
cc_415 N_A2_c_447_n N_A_533_367#_c_879_n 5.0837e-19 $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_416 N_A2_M1019_g N_A_533_367#_c_875_n 0.0143398f $X=9.175 $Y=2.465 $X2=0
+ $Y2=0
cc_417 N_A2_M1033_g N_A_533_367#_c_875_n 0.0157274f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_418 A2 N_A_533_367#_c_875_n 0.0692282f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_419 N_A2_c_453_n N_A_533_367#_c_875_n 0.00934834f $X=9.785 $Y=1.35 $X2=0
+ $Y2=0
cc_420 N_A2_M1014_g N_A_533_367#_c_876_n 0.00466344f $X=8.745 $Y=2.465 $X2=0
+ $Y2=0
cc_421 N_A2_c_447_n N_A_533_367#_c_876_n 0.00908491f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_422 N_A2_c_449_n N_A_533_367#_c_876_n 4.95511e-19 $X=8.365 $Y=1.615 $X2=0
+ $Y2=0
cc_423 A2 N_A_533_367#_c_876_n 0.0211316f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_424 N_A2_c_453_n N_A_533_367#_c_876_n 0.00256759f $X=9.785 $Y=1.35 $X2=0
+ $Y2=0
cc_425 N_A2_M1033_g N_A_533_367#_c_881_n 0.0046421f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_426 N_A2_c_447_n N_A_533_367#_c_927_n 0.0150119f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_427 N_A2_c_447_n N_A_533_367#_c_928_n 0.0146338f $X=8.245 $Y=1.7 $X2=0 $Y2=0
cc_428 N_A2_M1014_g N_A_533_367#_c_929_n 0.00154209f $X=8.745 $Y=2.465 $X2=0
+ $Y2=0
cc_429 N_A2_M1005_g N_VPWR_c_982_n 0.01469f $X=6.565 $Y=2.465 $X2=0 $Y2=0
cc_430 N_A2_M1014_g N_VPWR_c_985_n 0.014044f $X=8.745 $Y=2.465 $X2=0 $Y2=0
cc_431 N_A2_M1019_g N_VPWR_c_985_n 6.7059e-19 $X=9.175 $Y=2.465 $X2=0 $Y2=0
cc_432 N_A2_M1014_g N_VPWR_c_986_n 7.18684e-19 $X=8.745 $Y=2.465 $X2=0 $Y2=0
cc_433 N_A2_M1019_g N_VPWR_c_986_n 0.0174002f $X=9.175 $Y=2.465 $X2=0 $Y2=0
cc_434 N_A2_M1033_g N_VPWR_c_986_n 0.0194824f $X=9.605 $Y=2.465 $X2=0 $Y2=0
cc_435 N_A2_M1005_g N_VPWR_c_987_n 0.00525069f $X=6.565 $Y=2.465 $X2=0 $Y2=0
cc_436 N_A2_M1014_g N_VPWR_c_991_n 0.00486043f $X=8.745 $Y=2.465 $X2=0 $Y2=0
cc_437 N_A2_M1019_g N_VPWR_c_991_n 0.00486043f $X=9.175 $Y=2.465 $X2=0 $Y2=0
cc_438 N_A2_M1033_g N_VPWR_c_992_n 0.00486043f $X=9.605 $Y=2.465 $X2=0 $Y2=0
cc_439 N_A2_M1005_g N_VPWR_c_981_n 0.00928218f $X=6.565 $Y=2.465 $X2=0 $Y2=0
cc_440 N_A2_M1014_g N_VPWR_c_981_n 0.00824727f $X=8.745 $Y=2.465 $X2=0 $Y2=0
cc_441 N_A2_M1019_g N_VPWR_c_981_n 0.00824727f $X=9.175 $Y=2.465 $X2=0 $Y2=0
cc_442 N_A2_M1033_g N_VPWR_c_981_n 0.00917987f $X=9.605 $Y=2.465 $X2=0 $Y2=0
cc_443 N_A2_M1013_g N_VGND_c_1104_n 0.00539808f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_444 N_A2_c_441_n N_VGND_c_1105_n 0.0117408f $X=8.745 $Y=1.185 $X2=0 $Y2=0
cc_445 N_A2_c_443_n N_VGND_c_1105_n 0.0105703f $X=9.175 $Y=1.185 $X2=0 $Y2=0
cc_446 N_A2_c_445_n N_VGND_c_1105_n 5.75816e-19 $X=9.605 $Y=1.185 $X2=0 $Y2=0
cc_447 N_A2_c_443_n N_VGND_c_1107_n 6.24191e-19 $X=9.175 $Y=1.185 $X2=0 $Y2=0
cc_448 N_A2_c_445_n N_VGND_c_1107_n 0.0165374f $X=9.605 $Y=1.185 $X2=0 $Y2=0
cc_449 A2 N_VGND_c_1107_n 0.0239165f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_450 N_A2_c_453_n N_VGND_c_1107_n 0.00629958f $X=9.785 $Y=1.35 $X2=0 $Y2=0
cc_451 N_A2_M1013_g N_VGND_c_1117_n 0.00547467f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_452 N_A2_c_441_n N_VGND_c_1117_n 0.00486043f $X=8.745 $Y=1.185 $X2=0 $Y2=0
cc_453 N_A2_c_443_n N_VGND_c_1118_n 0.00486043f $X=9.175 $Y=1.185 $X2=0 $Y2=0
cc_454 N_A2_c_445_n N_VGND_c_1118_n 0.00486043f $X=9.605 $Y=1.185 $X2=0 $Y2=0
cc_455 N_A2_M1013_g N_VGND_c_1121_n 0.00644606f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_456 N_A2_c_441_n N_VGND_c_1121_n 0.0082726f $X=8.745 $Y=1.185 $X2=0 $Y2=0
cc_457 N_A2_c_443_n N_VGND_c_1121_n 0.00824727f $X=9.175 $Y=1.185 $X2=0 $Y2=0
cc_458 N_A2_c_445_n N_VGND_c_1121_n 0.00824727f $X=9.605 $Y=1.185 $X2=0 $Y2=0
cc_459 N_A2_M1013_g N_A_1334_47#_c_1273_n 0.00355848f $X=6.595 $Y=0.655 $X2=0
+ $Y2=0
cc_460 N_A2_c_448_n N_A_1334_47#_c_1274_n 0.004454f $X=8.365 $Y=1.435 $X2=0
+ $Y2=0
cc_461 A2 N_A_1334_47#_c_1274_n 0.0111312f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_462 N_A2_c_453_n N_A_1334_47#_c_1274_n 5.61757e-19 $X=9.785 $Y=1.35 $X2=0
+ $Y2=0
cc_463 N_A2_c_441_n N_A_1334_47#_c_1277_n 0.0121992f $X=8.745 $Y=1.185 $X2=0
+ $Y2=0
cc_464 N_A2_c_443_n N_A_1334_47#_c_1277_n 0.0122129f $X=9.175 $Y=1.185 $X2=0
+ $Y2=0
cc_465 A2 N_A_1334_47#_c_1277_n 0.0540388f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_466 N_A2_c_453_n N_A_1334_47#_c_1277_n 0.00470965f $X=9.785 $Y=1.35 $X2=0
+ $Y2=0
cc_467 N_A1_c_565_n N_Y_c_808_n 0.00419931f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_468 N_A1_c_574_n N_Y_c_808_n 0.00231647f $X=7.885 $Y=1.455 $X2=0 $Y2=0
cc_469 N_A1_c_567_n N_Y_c_809_n 0.0127021f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_470 N_A1_c_569_n N_Y_c_809_n 0.0127021f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_471 N_A1_c_570_n N_Y_c_809_n 0.00235915f $X=8.24 $Y=1.26 $X2=0 $Y2=0
cc_472 N_A1_c_571_n N_Y_c_809_n 4.8938e-19 $X=8.24 $Y=1.65 $X2=0 $Y2=0
cc_473 N_A1_c_572_n N_Y_c_809_n 0.00341274f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_474 N_A1_c_574_n N_Y_c_809_n 0.00231911f $X=7.885 $Y=1.455 $X2=0 $Y2=0
cc_475 N_A1_c_565_n N_Y_c_793_n 0.00712505f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_476 A1 N_Y_c_793_n 0.079349f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_477 N_A1_M1009_g N_A_533_367#_c_903_n 0.012941f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_478 N_A1_M1010_g N_A_533_367#_c_909_n 0.0122595f $X=7.455 $Y=2.465 $X2=0
+ $Y2=0
cc_479 N_A1_c_577_n N_A_533_367#_c_909_n 0.0122595f $X=7.885 $Y=1.725 $X2=0
+ $Y2=0
cc_480 N_A1_c_579_n N_A_533_367#_c_910_n 0.0119024f $X=8.315 $Y=1.725 $X2=0
+ $Y2=0
cc_481 N_A1_c_579_n N_A_533_367#_c_879_n 8.37992e-19 $X=8.315 $Y=1.725 $X2=0
+ $Y2=0
cc_482 N_A1_c_571_n N_A_533_367#_c_928_n 6.85025e-19 $X=8.24 $Y=1.65 $X2=0 $Y2=0
cc_483 N_A1_M1009_g N_VPWR_c_982_n 0.0125055f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_484 N_A1_M1010_g N_VPWR_c_982_n 6.56668e-19 $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_485 N_A1_M1009_g N_VPWR_c_983_n 6.78754e-19 $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_486 N_A1_M1010_g N_VPWR_c_983_n 0.0141705f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_487 N_A1_c_577_n N_VPWR_c_983_n 0.0141241f $X=7.885 $Y=1.725 $X2=0 $Y2=0
cc_488 N_A1_c_579_n N_VPWR_c_983_n 6.7059e-19 $X=8.315 $Y=1.725 $X2=0 $Y2=0
cc_489 N_A1_c_577_n N_VPWR_c_984_n 0.00486043f $X=7.885 $Y=1.725 $X2=0 $Y2=0
cc_490 N_A1_c_579_n N_VPWR_c_984_n 0.00486043f $X=8.315 $Y=1.725 $X2=0 $Y2=0
cc_491 N_A1_c_577_n N_VPWR_c_985_n 6.7059e-19 $X=7.885 $Y=1.725 $X2=0 $Y2=0
cc_492 N_A1_c_579_n N_VPWR_c_985_n 0.014044f $X=8.315 $Y=1.725 $X2=0 $Y2=0
cc_493 N_A1_M1009_g N_VPWR_c_989_n 0.00564095f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_494 N_A1_M1010_g N_VPWR_c_989_n 0.00486043f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_495 N_A1_M1009_g N_VPWR_c_981_n 0.00948291f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_496 N_A1_M1010_g N_VPWR_c_981_n 0.00824727f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_497 N_A1_c_577_n N_VPWR_c_981_n 0.00824727f $X=7.885 $Y=1.725 $X2=0 $Y2=0
cc_498 N_A1_c_579_n N_VPWR_c_981_n 0.00824727f $X=8.315 $Y=1.725 $X2=0 $Y2=0
cc_499 N_A1_c_572_n N_VGND_c_1105_n 0.00109252f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_500 N_A1_c_565_n N_VGND_c_1117_n 0.00357877f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_501 N_A1_c_567_n N_VGND_c_1117_n 0.00357877f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_502 N_A1_c_569_n N_VGND_c_1117_n 0.00357877f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_503 N_A1_c_572_n N_VGND_c_1117_n 0.00357877f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_504 N_A1_c_565_n N_VGND_c_1121_n 0.00537654f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_505 N_A1_c_567_n N_VGND_c_1121_n 0.0053512f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_506 N_A1_c_569_n N_VGND_c_1121_n 0.0053512f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_507 N_A1_c_572_n N_VGND_c_1121_n 0.00537654f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_508 N_A1_c_565_n N_A_1334_47#_c_1273_n 0.0116856f $X=7.025 $Y=1.185 $X2=0
+ $Y2=0
cc_509 N_A1_c_567_n N_A_1334_47#_c_1273_n 0.0104569f $X=7.455 $Y=1.185 $X2=0
+ $Y2=0
cc_510 N_A1_c_569_n N_A_1334_47#_c_1273_n 0.0103812f $X=7.885 $Y=1.185 $X2=0
+ $Y2=0
cc_511 N_A1_c_572_n N_A_1334_47#_c_1273_n 0.0148497f $X=8.315 $Y=1.185 $X2=0
+ $Y2=0
cc_512 N_A_85_367#_c_659_n N_Y_M1016_d 0.00332344f $X=1.315 $Y=2.99 $X2=0 $Y2=0
cc_513 N_A_85_367#_c_661_n N_Y_M1031_d 0.00332344f $X=2.175 $Y=2.99 $X2=0 $Y2=0
cc_514 N_A_85_367#_c_651_n N_Y_c_739_n 0.0352831f $X=0.55 $Y=1.98 $X2=0 $Y2=0
cc_515 N_A_85_367#_c_659_n N_Y_c_739_n 0.0159805f $X=1.315 $Y=2.99 $X2=0 $Y2=0
cc_516 N_A_85_367#_c_691_p N_Y_c_727_n 0.0145583f $X=1.41 $Y=2.11 $X2=0 $Y2=0
cc_517 N_A_85_367#_c_661_n N_Y_c_756_n 0.0159805f $X=2.175 $Y=2.99 $X2=0 $Y2=0
cc_518 N_A_85_367#_c_652_n N_Y_c_729_n 0.0209937f $X=2.305 $Y=2.115 $X2=0 $Y2=0
cc_519 N_A_85_367#_c_654_n N_Y_c_729_n 0.0168539f $X=3.055 $Y=2.03 $X2=0 $Y2=0
cc_520 N_A_85_367#_c_654_n N_A_533_367#_M1004_d 0.0055232f $X=3.055 $Y=2.03
+ $X2=-0.19 $Y2=1.655
cc_521 N_A_85_367#_c_671_n N_A_533_367#_M1008_d 0.00416883f $X=5.8 $Y=2.435
+ $X2=0 $Y2=0
cc_522 N_A_85_367#_c_671_n N_A_533_367#_M1003_d 0.00347245f $X=5.8 $Y=2.435
+ $X2=0 $Y2=0
cc_523 N_A_85_367#_c_671_n N_A_533_367#_M1030_d 0.00347245f $X=5.8 $Y=2.435
+ $X2=0 $Y2=0
cc_524 N_A_85_367#_c_653_n N_A_533_367#_c_877_n 0.0366457f $X=2.305 $Y=2.905
+ $X2=0 $Y2=0
cc_525 N_A_85_367#_c_654_n N_A_533_367#_c_877_n 0.0220026f $X=3.055 $Y=2.03
+ $X2=0 $Y2=0
cc_526 N_A_85_367#_M1004_s N_A_533_367#_c_888_n 0.00338379f $X=3.08 $Y=1.835
+ $X2=0 $Y2=0
cc_527 N_A_85_367#_M1023_s N_A_533_367#_c_888_n 0.00338818f $X=3.94 $Y=1.835
+ $X2=0 $Y2=0
cc_528 N_A_85_367#_M1011_s N_A_533_367#_c_888_n 0.00338818f $X=4.8 $Y=1.835
+ $X2=0 $Y2=0
cc_529 N_A_85_367#_M1035_s N_A_533_367#_c_888_n 0.00337733f $X=5.66 $Y=1.835
+ $X2=0 $Y2=0
cc_530 N_A_85_367#_c_654_n N_A_533_367#_c_888_n 0.00229198f $X=3.055 $Y=2.03
+ $X2=0 $Y2=0
cc_531 N_A_85_367#_c_706_p N_A_533_367#_c_888_n 0.0135088f $X=3.225 $Y=2.27
+ $X2=0 $Y2=0
cc_532 N_A_85_367#_c_671_n N_A_533_367#_c_888_n 0.14238f $X=5.8 $Y=2.435 $X2=0
+ $Y2=0
cc_533 N_A_85_367#_c_655_n N_A_533_367#_c_888_n 5.68856e-19 $X=3.22 $Y=1.96
+ $X2=0 $Y2=0
cc_534 N_A_85_367#_c_653_n N_A_533_367#_c_878_n 0.0255317f $X=2.305 $Y=2.905
+ $X2=0 $Y2=0
cc_535 N_A_85_367#_c_650_n N_VPWR_c_987_n 0.0179183f $X=0.515 $Y=2.905 $X2=0
+ $Y2=0
cc_536 N_A_85_367#_c_659_n N_VPWR_c_987_n 0.0361172f $X=1.315 $Y=2.99 $X2=0
+ $Y2=0
cc_537 N_A_85_367#_c_661_n N_VPWR_c_987_n 0.0361172f $X=2.175 $Y=2.99 $X2=0
+ $Y2=0
cc_538 N_A_85_367#_c_653_n N_VPWR_c_987_n 0.0179183f $X=2.305 $Y=2.905 $X2=0
+ $Y2=0
cc_539 N_A_85_367#_c_714_p N_VPWR_c_987_n 0.0125234f $X=1.41 $Y=2.99 $X2=0 $Y2=0
cc_540 N_A_85_367#_M1016_s N_VPWR_c_981_n 0.00215161f $X=0.425 $Y=1.835 $X2=0
+ $Y2=0
cc_541 N_A_85_367#_M1022_s N_VPWR_c_981_n 0.00223565f $X=1.27 $Y=1.835 $X2=0
+ $Y2=0
cc_542 N_A_85_367#_M1037_s N_VPWR_c_981_n 0.00215161f $X=2.13 $Y=1.835 $X2=0
+ $Y2=0
cc_543 N_A_85_367#_M1004_s N_VPWR_c_981_n 0.00225186f $X=3.08 $Y=1.835 $X2=0
+ $Y2=0
cc_544 N_A_85_367#_M1023_s N_VPWR_c_981_n 0.00225186f $X=3.94 $Y=1.835 $X2=0
+ $Y2=0
cc_545 N_A_85_367#_M1011_s N_VPWR_c_981_n 0.00225186f $X=4.8 $Y=1.835 $X2=0
+ $Y2=0
cc_546 N_A_85_367#_M1035_s N_VPWR_c_981_n 0.00225186f $X=5.66 $Y=1.835 $X2=0
+ $Y2=0
cc_547 N_A_85_367#_c_650_n N_VPWR_c_981_n 0.0101029f $X=0.515 $Y=2.905 $X2=0
+ $Y2=0
cc_548 N_A_85_367#_c_659_n N_VPWR_c_981_n 0.023676f $X=1.315 $Y=2.99 $X2=0 $Y2=0
cc_549 N_A_85_367#_c_661_n N_VPWR_c_981_n 0.023676f $X=2.175 $Y=2.99 $X2=0 $Y2=0
cc_550 N_A_85_367#_c_653_n N_VPWR_c_981_n 0.0101082f $X=2.305 $Y=2.905 $X2=0
+ $Y2=0
cc_551 N_A_85_367#_c_714_p N_VPWR_c_981_n 0.00738676f $X=1.41 $Y=2.99 $X2=0
+ $Y2=0
cc_552 N_Y_M1016_d N_VPWR_c_981_n 0.00225186f $X=0.84 $Y=1.835 $X2=0 $Y2=0
cc_553 N_Y_M1031_d N_VPWR_c_981_n 0.00225186f $X=1.7 $Y=1.835 $X2=0 $Y2=0
cc_554 N_Y_c_750_n N_VGND_M1025_d 0.00329816f $X=1.915 $Y=0.955 $X2=0 $Y2=0
cc_555 N_Y_c_762_n N_VGND_M1036_d 0.00220534f $X=2.435 $Y=0.955 $X2=0 $Y2=0
cc_556 N_Y_c_734_n N_VGND_M1036_d 0.00144333f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_557 N_Y_c_731_n N_VGND_M1002_s 0.00178782f $X=3.695 $Y=1.135 $X2=0 $Y2=0
cc_558 N_Y_c_793_n N_VGND_M1034_s 0.0105792f $X=7.075 $Y=0.865 $X2=0 $Y2=0
cc_559 N_Y_c_750_n N_VGND_c_1101_n 0.0170777f $X=1.915 $Y=0.955 $X2=0 $Y2=0
cc_560 N_Y_c_762_n N_VGND_c_1102_n 0.00809557f $X=2.435 $Y=0.955 $X2=0 $Y2=0
cc_561 N_Y_c_734_n N_VGND_c_1102_n 0.00992353f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_562 N_Y_c_793_n N_VGND_c_1104_n 0.0213572f $X=7.075 $Y=0.865 $X2=0 $Y2=0
cc_563 N_Y_c_843_p N_VGND_c_1108_n 0.0124525f $X=1.15 $Y=0.42 $X2=0 $Y2=0
cc_564 N_Y_c_844_p N_VGND_c_1110_n 0.0124525f $X=2.01 $Y=0.42 $X2=0 $Y2=0
cc_565 N_Y_M1007_s N_VGND_c_1121_n 0.00536646f $X=1.01 $Y=0.235 $X2=0 $Y2=0
cc_566 N_Y_M1028_s N_VGND_c_1121_n 0.00536646f $X=1.87 $Y=0.235 $X2=0 $Y2=0
cc_567 N_Y_M1006_s N_VGND_c_1121_n 0.00225186f $X=4.3 $Y=0.235 $X2=0 $Y2=0
cc_568 N_Y_M1026_s N_VGND_c_1121_n 0.00225186f $X=5.16 $Y=0.235 $X2=0 $Y2=0
cc_569 N_Y_M1000_s N_VGND_c_1121_n 0.00225186f $X=7.1 $Y=0.235 $X2=0 $Y2=0
cc_570 N_Y_M1020_s N_VGND_c_1121_n 0.00225186f $X=7.96 $Y=0.235 $X2=0 $Y2=0
cc_571 N_Y_c_843_p N_VGND_c_1121_n 0.00730901f $X=1.15 $Y=0.42 $X2=0 $Y2=0
cc_572 N_Y_c_844_p N_VGND_c_1121_n 0.00730901f $X=2.01 $Y=0.42 $X2=0 $Y2=0
cc_573 N_Y_c_732_n N_VGND_c_1121_n 0.00124096f $X=5.965 $Y=0.945 $X2=0 $Y2=0
cc_574 N_Y_c_793_n N_VGND_c_1121_n 0.0103847f $X=7.075 $Y=0.865 $X2=0 $Y2=0
cc_575 N_Y_c_731_n N_A_546_47#_M1001_d 0.00178346f $X=3.695 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_576 N_Y_c_731_n N_A_546_47#_M1021_d 5.04957e-19 $X=3.695 $Y=1.135 $X2=0 $Y2=0
cc_577 N_Y_c_736_n N_A_546_47#_M1021_d 0.00958745f $X=4.2 $Y=0.97 $X2=0 $Y2=0
cc_578 N_Y_c_735_n N_A_546_47#_M1012_d 0.00178117f $X=5.39 $Y=0.97 $X2=0 $Y2=0
cc_579 N_Y_c_732_n N_A_546_47#_M1027_d 0.0127565f $X=5.965 $Y=0.945 $X2=0 $Y2=0
cc_580 N_Y_c_731_n N_A_546_47#_c_1237_n 0.0332304f $X=3.695 $Y=1.135 $X2=0 $Y2=0
cc_581 N_Y_M1006_s N_A_546_47#_c_1239_n 0.00339639f $X=4.3 $Y=0.235 $X2=0 $Y2=0
cc_582 N_Y_M1026_s N_A_546_47#_c_1239_n 0.00339639f $X=5.16 $Y=0.235 $X2=0 $Y2=0
cc_583 N_Y_c_732_n N_A_546_47#_c_1239_n 0.0346386f $X=5.965 $Y=0.945 $X2=0 $Y2=0
cc_584 N_Y_c_735_n N_A_546_47#_c_1239_n 0.0686814f $X=5.39 $Y=0.97 $X2=0 $Y2=0
cc_585 N_Y_c_736_n N_A_546_47#_c_1239_n 0.0188632f $X=4.2 $Y=0.97 $X2=0 $Y2=0
cc_586 N_Y_c_731_n N_A_546_47#_c_1255_n 0.0130987f $X=3.695 $Y=1.135 $X2=0 $Y2=0
cc_587 N_Y_c_731_n N_A_546_47#_c_1243_n 0.00391474f $X=3.695 $Y=1.135 $X2=0
+ $Y2=0
cc_588 N_Y_c_736_n N_A_546_47#_c_1243_n 0.0172002f $X=4.2 $Y=0.97 $X2=0 $Y2=0
cc_589 N_Y_c_793_n N_A_1334_47#_M1013_s 0.00499536f $X=7.075 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_590 N_Y_c_809_n N_A_1334_47#_M1017_d 0.00332201f $X=8.1 $Y=0.865 $X2=0 $Y2=0
cc_591 N_Y_M1000_s N_A_1334_47#_c_1273_n 0.00329779f $X=7.1 $Y=0.235 $X2=0 $Y2=0
cc_592 N_Y_M1020_s N_A_1334_47#_c_1273_n 0.00329779f $X=7.96 $Y=0.235 $X2=0
+ $Y2=0
cc_593 N_Y_c_808_n N_A_1334_47#_c_1273_n 0.0616052f $X=7.24 $Y=0.865 $X2=0 $Y2=0
cc_594 N_Y_c_793_n N_A_1334_47#_c_1273_n 0.0106197f $X=7.075 $Y=0.865 $X2=0
+ $Y2=0
cc_595 N_A_533_367#_c_903_n N_VPWR_M1005_s 0.0040891f $X=7.135 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_596 N_A_533_367#_c_909_n N_VPWR_M1010_s 0.00339614f $X=8.005 $Y=2.04 $X2=0
+ $Y2=0
cc_597 N_A_533_367#_c_910_n N_VPWR_M1038_s 0.00448631f $X=8.795 $Y=2.04 $X2=0
+ $Y2=0
cc_598 N_A_533_367#_c_903_n N_VPWR_c_982_n 0.0172332f $X=7.135 $Y=2.04 $X2=0
+ $Y2=0
cc_599 N_A_533_367#_c_909_n N_VPWR_c_983_n 0.0170777f $X=8.005 $Y=2.04 $X2=0
+ $Y2=0
cc_600 N_A_533_367#_c_956_p N_VPWR_c_984_n 0.0124525f $X=8.1 $Y=2.475 $X2=0
+ $Y2=0
cc_601 N_A_533_367#_c_910_n N_VPWR_c_985_n 0.0170777f $X=8.795 $Y=2.04 $X2=0
+ $Y2=0
cc_602 N_A_533_367#_c_875_n N_VPWR_c_986_n 0.0216087f $X=9.725 $Y=1.69 $X2=0
+ $Y2=0
cc_603 N_A_533_367#_c_888_n N_VPWR_c_987_n 0.181339f $X=6.135 $Y=2.922 $X2=0
+ $Y2=0
cc_604 N_A_533_367#_c_878_n N_VPWR_c_987_n 0.0211865f $X=2.955 $Y=2.922 $X2=0
+ $Y2=0
cc_605 N_A_533_367#_c_961_p N_VPWR_c_987_n 0.0213157f $X=6.295 $Y=2.77 $X2=0
+ $Y2=0
cc_606 N_A_533_367#_c_962_p N_VPWR_c_989_n 0.0128073f $X=7.24 $Y=2.475 $X2=0
+ $Y2=0
cc_607 N_A_533_367#_c_963_p N_VPWR_c_991_n 0.0124525f $X=8.96 $Y=2.44 $X2=0
+ $Y2=0
cc_608 N_A_533_367#_c_881_n N_VPWR_c_992_n 0.0178111f $X=9.82 $Y=1.98 $X2=0
+ $Y2=0
cc_609 N_A_533_367#_M1004_d N_VPWR_c_981_n 0.00215158f $X=2.665 $Y=1.835 $X2=0
+ $Y2=0
cc_610 N_A_533_367#_M1008_d N_VPWR_c_981_n 0.00223577f $X=3.51 $Y=1.835 $X2=0
+ $Y2=0
cc_611 N_A_533_367#_M1003_d N_VPWR_c_981_n 0.00223577f $X=4.37 $Y=1.835 $X2=0
+ $Y2=0
cc_612 N_A_533_367#_M1030_d N_VPWR_c_981_n 0.00223577f $X=5.23 $Y=1.835 $X2=0
+ $Y2=0
cc_613 N_A_533_367#_M1032_d N_VPWR_c_981_n 0.00444771f $X=6.09 $Y=1.835 $X2=0
+ $Y2=0
cc_614 N_A_533_367#_M1009_d N_VPWR_c_981_n 0.00501859f $X=7.1 $Y=1.835 $X2=0
+ $Y2=0
cc_615 N_A_533_367#_M1024_d N_VPWR_c_981_n 0.00536646f $X=7.96 $Y=1.835 $X2=0
+ $Y2=0
cc_616 N_A_533_367#_M1014_d N_VPWR_c_981_n 0.00536646f $X=8.82 $Y=1.835 $X2=0
+ $Y2=0
cc_617 N_A_533_367#_M1033_d N_VPWR_c_981_n 0.00371702f $X=9.68 $Y=1.835 $X2=0
+ $Y2=0
cc_618 N_A_533_367#_c_888_n N_VPWR_c_981_n 0.115318f $X=6.135 $Y=2.922 $X2=0
+ $Y2=0
cc_619 N_A_533_367#_c_878_n N_VPWR_c_981_n 0.0126421f $X=2.955 $Y=2.922 $X2=0
+ $Y2=0
cc_620 N_A_533_367#_c_961_p N_VPWR_c_981_n 0.0124409f $X=6.295 $Y=2.77 $X2=0
+ $Y2=0
cc_621 N_A_533_367#_c_962_p N_VPWR_c_981_n 0.00769778f $X=7.24 $Y=2.475 $X2=0
+ $Y2=0
cc_622 N_A_533_367#_c_956_p N_VPWR_c_981_n 0.00730901f $X=8.1 $Y=2.475 $X2=0
+ $Y2=0
cc_623 N_A_533_367#_c_963_p N_VPWR_c_981_n 0.00730901f $X=8.96 $Y=2.44 $X2=0
+ $Y2=0
cc_624 N_A_533_367#_c_881_n N_VPWR_c_981_n 0.0100304f $X=9.82 $Y=1.98 $X2=0
+ $Y2=0
cc_625 N_VGND_c_1121_n N_A_546_47#_M1001_d 0.00437356f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_626 N_VGND_c_1121_n N_A_546_47#_M1021_d 0.00473013f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_627 N_VGND_c_1121_n N_A_546_47#_M1012_d 0.00223577f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_628 N_VGND_c_1121_n N_A_546_47#_M1027_d 0.00497397f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_629 N_VGND_M1002_s N_A_546_47#_c_1237_n 0.00335844f $X=3.16 $Y=0.235 $X2=0
+ $Y2=0
cc_630 N_VGND_c_1103_n N_A_546_47#_c_1237_n 0.0161939f $X=3.3 $Y=0.38 $X2=0
+ $Y2=0
cc_631 N_VGND_c_1112_n N_A_546_47#_c_1237_n 0.00224524f $X=3.135 $Y=0 $X2=0
+ $Y2=0
cc_632 N_VGND_c_1114_n N_A_546_47#_c_1237_n 0.00225133f $X=6.135 $Y=0 $X2=0
+ $Y2=0
cc_633 N_VGND_c_1121_n N_A_546_47#_c_1237_n 0.00952646f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_634 N_VGND_c_1114_n N_A_546_47#_c_1239_n 0.126445f $X=6.135 $Y=0 $X2=0 $Y2=0
cc_635 N_VGND_c_1121_n N_A_546_47#_c_1239_n 0.0787666f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_636 N_VGND_c_1112_n N_A_546_47#_c_1255_n 0.00446942f $X=3.135 $Y=0 $X2=0
+ $Y2=0
cc_637 N_VGND_c_1121_n N_A_546_47#_c_1255_n 0.00609473f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_638 N_VGND_c_1114_n N_A_546_47#_c_1243_n 0.0120113f $X=6.135 $Y=0 $X2=0 $Y2=0
cc_639 N_VGND_c_1121_n N_A_546_47#_c_1243_n 0.00689462f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_640 N_VGND_c_1121_n N_A_1334_47#_M1013_s 0.00223577f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_641 N_VGND_c_1121_n N_A_1334_47#_M1017_d 0.00223577f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_642 N_VGND_c_1121_n N_A_1334_47#_M1039_d 0.00376626f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_643 N_VGND_c_1121_n N_A_1334_47#_M1018_s 0.00536646f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_644 N_VGND_c_1117_n N_A_1334_47#_c_1273_n 0.100358f $X=8.795 $Y=0 $X2=0 $Y2=0
cc_645 N_VGND_c_1121_n N_A_1334_47#_c_1273_n 0.0644219f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_646 N_VGND_c_1117_n N_A_1334_47#_c_1297_n 0.0128782f $X=8.795 $Y=0 $X2=0
+ $Y2=0
cc_647 N_VGND_c_1121_n N_A_1334_47#_c_1297_n 0.00777554f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_648 N_VGND_M1015_d N_A_1334_47#_c_1277_n 0.00329816f $X=8.82 $Y=0.235 $X2=0
+ $Y2=0
cc_649 N_VGND_c_1105_n N_A_1334_47#_c_1277_n 0.0170777f $X=8.96 $Y=0.575 $X2=0
+ $Y2=0
cc_650 N_VGND_c_1118_n N_A_1334_47#_c_1301_n 0.0124525f $X=9.655 $Y=0 $X2=0
+ $Y2=0
cc_651 N_VGND_c_1121_n N_A_1334_47#_c_1301_n 0.00730901f $X=9.84 $Y=0 $X2=0
+ $Y2=0
