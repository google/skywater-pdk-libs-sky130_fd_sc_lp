* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_313_365# A3 a_615_365# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VGND A2 a_155_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_155_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_313_365# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_155_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_615_365# A3 a_313_365# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Y A4 a_313_365# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND A4 a_155_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_155_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VPWR A1 a_808_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_808_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_615_365# A2 a_808_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 Y B1 a_155_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_808_367# A2 a_615_365# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_155_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VGND A3 a_155_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 VGND A1 a_155_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_155_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
