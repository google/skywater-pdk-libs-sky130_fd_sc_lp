* File: sky130_fd_sc_lp__a2111o_m.pex.spice
* Created: Fri Aug 28 09:46:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111O_M%A_85_21# 1 2 3 12 16 20 21 24 25 27 28 33
+ 36 37 38 41
c89 16 0 1.34772e-19 $X=0.5 $Y=2.745
r90 39 41 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.225 $Y=0.725
+ $X2=2.225 $Y2=0.51
r91 38 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.81
+ $X2=1.56 $Y2=0.81
r92 37 39 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.12 $Y=0.81
+ $X2=2.225 $Y2=0.725
r93 37 38 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.12 $Y=0.81
+ $X2=1.645 $Y2=0.81
r94 35 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=0.895
+ $X2=1.56 $Y2=0.81
r95 35 36 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=1.56 $Y=0.895
+ $X2=1.56 $Y2=1.93
r96 31 45 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.365 $Y=0.81
+ $X2=1.56 $Y2=0.81
r97 31 33 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.365 $Y=0.725
+ $X2=1.365 $Y2=0.51
r98 28 30 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=1.045 $Y2=2.035
r99 27 36 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.475 $Y=2.035
+ $X2=1.56 $Y2=1.93
r100 27 30 22.71 $w=2.08e-07 $l=4.3e-07 $layer=LI1_cond $X=1.475 $Y=2.035
+ $X2=1.045 $Y2=2.035
r101 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.635 $X2=0.59 $Y2=1.635
r102 22 28 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.59 $Y=1.93
+ $X2=0.675 $Y2=2.035
r103 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.59 $Y=1.93
+ $X2=0.59 $Y2=1.635
r104 20 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.59 $Y=1.975
+ $X2=0.59 $Y2=1.635
r105 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.975
+ $X2=0.59 $Y2=2.14
r106 19 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.47
+ $X2=0.59 $Y2=1.635
r107 16 21 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=0.5 $Y=2.745
+ $X2=0.5 $Y2=2.14
r108 12 19 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=0.5 $Y=0.445
+ $X2=0.5 $Y2=1.47
r109 3 30 600 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_PDIFF $count=1 $X=0.92
+ $Y=1.845 $X2=1.045 $Y2=2.035
r110 2 41 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.235 $X2=2.225 $Y2=0.51
r111 1 33 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.235 $X2=1.365 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_M%D1 3 7 12 13 14 15 19 20
r45 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.13
+ $Y=1.18 $X2=1.13 $Y2=1.18
r46 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.13 $Y=1.295
+ $X2=1.13 $Y2=1.665
r47 14 20 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.13 $Y=1.295
+ $X2=1.13 $Y2=1.18
r48 12 19 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.13 $Y=1.535
+ $X2=1.13 $Y2=1.18
r49 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.15 $Y=1.535
+ $X2=1.15 $Y2=1.685
r50 10 19 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.015
+ $X2=1.13 $Y2=1.18
r51 7 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.26 $Y=2.055
+ $X2=1.26 $Y2=1.685
r52 3 10 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.15 $Y=0.445
+ $X2=1.15 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_M%C1 3 8 10 11 12 13
c47 12 0 1.13753e-19 $X=1.2 $Y=2.405
r48 13 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=2.8 $X2=1.165 $Y2=2.8
r49 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.165 $Y=2.405
+ $X2=1.165 $Y2=2.775
r50 11 17 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=1.545 $Y=2.8
+ $X2=1.165 $Y2=2.8
r51 9 10 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.6 $Y=1.145 $X2=1.6
+ $Y2=1.295
r52 8 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.62 $Y=2.055
+ $X2=1.62 $Y2=1.295
r53 6 11 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.62 $Y=2.635
+ $X2=1.545 $Y2=2.8
r54 6 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.62 $Y=2.635 $X2=1.62
+ $Y2=2.055
r55 3 9 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=1.58 $Y=0.445 $X2=1.58
+ $Y2=1.145
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_M%B1 4 7 10 11 12 18 19 22
c51 19 0 7.15014e-20 $X=2.07 $Y=2.9
c52 18 0 1.13753e-19 $X=2.07 $Y=2.9
r53 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=2.9
+ $X2=2.07 $Y2=2.735
r54 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=2.9 $X2=2.07 $Y2=2.9
r55 12 22 3.83311 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=1.632 $Y=2.9
+ $X2=1.632 $Y2=2.735
r56 12 19 8.94118 $w=4.53e-07 $l=3.05e-07 $layer=LI1_cond $X=1.765 $Y=2.9
+ $X2=2.07 $Y2=2.9
r57 12 22 1.00023 $w=2.63e-07 $l=2.3e-08 $layer=LI1_cond $X=1.632 $Y=2.712
+ $X2=1.632 $Y2=2.735
r58 11 12 13.3509 $w=2.63e-07 $l=3.07e-07 $layer=LI1_cond $X=1.632 $Y=2.405
+ $X2=1.632 $Y2=2.712
r59 9 10 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.995 $Y=1.585
+ $X2=1.995 $Y2=1.735
r60 7 9 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=2.01 $Y=0.445
+ $X2=2.01 $Y2=1.585
r61 4 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.98 $Y=2.055
+ $X2=1.98 $Y2=2.735
r62 4 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.98 $Y=2.055
+ $X2=1.98 $Y2=1.735
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_M%A1 4 7 10 12 15 17 18
c49 18 0 3.5305e-20 $X=3.12 $Y=2.775
c50 15 0 1.5666e-19 $X=2.52 $Y=2.45
c51 12 0 1.42179e-19 $X=2.425 $Y=1.635
c52 10 0 8.15188e-20 $X=2.52 $Y=2.665
r53 25 31 1.01705 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=3.047 $Y=2.665
+ $X2=3.047 $Y2=2.83
r54 24 31 9.1497 $w=3.28e-07 $l=2.62e-07 $layer=LI1_cond $X=2.785 $Y=2.83
+ $X2=3.047 $Y2=2.83
r55 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.785
+ $Y=2.83 $X2=2.785 $Y2=2.83
r56 18 31 2.54934 $w=3.28e-07 $l=7.3e-08 $layer=LI1_cond $X=3.12 $Y=2.83
+ $X2=3.047 $Y2=2.83
r57 17 25 9.51223 $w=3.13e-07 $l=2.6e-07 $layer=LI1_cond $X=3.047 $Y=2.405
+ $X2=3.047 $Y2=2.665
r58 13 15 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=2.41 $Y=2.45
+ $X2=2.52 $Y2=2.45
r59 11 12 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.425 $Y=1.485
+ $X2=2.425 $Y2=1.635
r60 10 23 47.839 $w=2.67e-07 $l=3.37565e-07 $layer=POLY_cond $X=2.52 $Y=2.665
+ $X2=2.785 $Y2=2.83
r61 9 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.52 $Y=2.525
+ $X2=2.52 $Y2=2.45
r62 9 10 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.52 $Y=2.525
+ $X2=2.52 $Y2=2.665
r63 7 11 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.44 $Y=0.445
+ $X2=2.44 $Y2=1.485
r64 4 12 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.41 $Y=2.055
+ $X2=2.41 $Y2=1.635
r65 2 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.41 $Y=2.375
+ $X2=2.41 $Y2=2.45
r66 2 4 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.41 $Y=2.375 $X2=2.41
+ $Y2=2.055
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_M%A2 3 6 9 10 11 12 14 21
r30 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.89
+ $Y=0.93 $X2=2.89 $Y2=0.93
r31 14 22 5.09441 $w=5.38e-07 $l=2.3e-07 $layer=LI1_cond $X=3.12 $Y=1.11
+ $X2=2.89 $Y2=1.11
r32 12 22 5.5374 $w=5.38e-07 $l=2.5e-07 $layer=LI1_cond $X=2.64 $Y=1.11 $X2=2.89
+ $Y2=1.11
r33 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.89 $Y=1.27
+ $X2=2.89 $Y2=0.93
r34 10 11 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=1.27
+ $X2=2.89 $Y2=1.435
r35 9 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=0.765
+ $X2=2.89 $Y2=0.93
r36 6 11 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.88 $Y=2.055
+ $X2=2.88 $Y2=1.435
r37 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.8 $Y=0.445 $X2=2.8
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_M%X 1 2 7 8 9 10 11 12 13
c16 13 0 1.34772e-19 $X=0.24 $Y=2.775
r17 13 40 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=2.695
+ $X2=0.272 $Y2=2.53
r18 12 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=2.405
+ $X2=0.24 $Y2=2.53
r19 11 12 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.405
r20 10 11 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r21 9 10 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295 $X2=0.24
+ $Y2=1.665
r22 8 9 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925 $X2=0.24
+ $Y2=1.295
r23 8 37 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=0.675
r24 7 37 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=0.51
+ $X2=0.272 $Y2=0.675
r25 2 13 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.535 $X2=0.285 $Y2=2.695
r26 1 7 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_M%VPWR 1 2 9 12 15 19 22 23 24 26 39 40 43
c57 40 0 1.5666e-19 $X=3.12 $Y=3.33
c58 19 0 1.2895e-19 $X=2.615 $Y=2.4
r59 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 34 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r65 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 31 43 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.715 $Y2=3.33
r67 31 33 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33 $X2=1.2
+ $Y2=3.33
r68 29 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r70 26 43 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.61 $Y=3.33
+ $X2=0.715 $Y2=3.33
r71 26 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.61 $Y=3.33 $X2=0.24
+ $Y2=3.33
r72 24 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r73 24 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r74 22 36 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 22 23 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=2.435 $Y2=3.33
r76 21 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.53 $Y=3.33 $X2=3.12
+ $Y2=3.33
r77 21 23 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.53 $Y=3.33
+ $X2=2.435 $Y2=3.33
r78 17 19 10.5072 $w=1.88e-07 $l=1.8e-07 $layer=LI1_cond $X=2.435 $Y=2.4
+ $X2=2.615 $Y2=2.4
r79 13 19 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.615 $Y=2.305
+ $X2=2.615 $Y2=2.4
r80 13 15 10.799 $w=1.88e-07 $l=1.85e-07 $layer=LI1_cond $X=2.615 $Y=2.305
+ $X2=2.615 $Y2=2.12
r81 12 23 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=3.245
+ $X2=2.435 $Y2=3.33
r82 11 17 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.435 $Y=2.495
+ $X2=2.435 $Y2=2.4
r83 11 12 43.7799 $w=1.88e-07 $l=7.5e-07 $layer=LI1_cond $X=2.435 $Y=2.495
+ $X2=2.435 $Y2=3.245
r84 7 43 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=3.33
r85 7 9 22.974 $w=2.08e-07 $l=4.35e-07 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=2.81
r86 2 15 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.845 $X2=2.625 $Y2=2.12
r87 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.535 $X2=0.715 $Y2=2.81
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_M%A_411_369# 1 2 9 11 12 13
c30 13 0 5.85507e-20 $X=3.095 $Y=1.69
r31 13 16 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.095 $Y=1.69
+ $X2=3.095 $Y2=1.99
r32 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=1.69
+ $X2=3.095 $Y2=1.69
r33 11 12 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.93 $Y=1.69 $X2=2.3
+ $Y2=1.69
r34 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.195 $Y=1.775
+ $X2=2.3 $Y2=1.69
r35 7 9 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=2.195 $Y=1.775
+ $X2=2.195 $Y2=1.97
r36 2 16 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.845 $X2=3.095 $Y2=1.99
r37 1 9 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.845 $X2=2.195 $Y2=1.97
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_M%VGND 1 2 3 12 16 18 20 23 24 25 27 36 41 45
r46 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r49 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r50 36 44 4.60552 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=3.105
+ $Y2=0
r51 36 38 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=2.64
+ $Y2=0
r52 32 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=0.735
+ $Y2=0
r53 32 34 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=1.68
+ $Y2=0
r54 30 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r55 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r56 27 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.735
+ $Y2=0
r57 27 29 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.24
+ $Y2=0
r58 25 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r59 25 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r60 25 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r61 23 34 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.69 $Y=0 $X2=1.68
+ $Y2=0
r62 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.69 $Y=0 $X2=1.795
+ $Y2=0
r63 22 38 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=2.64
+ $Y2=0
r64 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=1.795
+ $Y2=0
r65 18 44 3.16065 $w=3.3e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.105 $Y2=0
r66 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0.38
r67 14 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=0.085
+ $X2=1.795 $Y2=0
r68 14 16 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.795 $Y=0.085
+ $X2=1.795 $Y2=0.38
r69 10 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0
r70 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0.38
r71 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.235 $X2=3.015 $Y2=0.38
r72 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.235 $X2=1.795 $Y2=0.38
r73 1 12 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.735 $Y2=0.38
.ends

