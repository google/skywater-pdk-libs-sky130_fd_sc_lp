* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 VGND A3 a_132_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 Y A3 a_49_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VGND A3 a_132_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR A1 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND A2 a_132_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND A1 a_132_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_132_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR A1 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_132_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_132_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_49_367# A2 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 Y B1 a_132_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND A2 a_132_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_132_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_132_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_49_367# A2 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_49_367# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 Y A3 a_49_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_132_367# A2 a_49_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_132_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_132_367# A2 a_49_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_49_367# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_132_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_132_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VGND A1 a_132_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 Y B1 a_132_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 a_132_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 a_132_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
