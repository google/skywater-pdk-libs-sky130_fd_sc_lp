* File: sky130_fd_sc_lp__nor2b_lp.pex.spice
* Created: Wed Sep  2 10:08:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2B_LP%A 3 7 11 15 17 18 20 22 31
c35 22 0 1.69014e-19 $X=1.2 $Y=1.665
r36 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.99
+ $Y=1.275 $X2=0.99 $Y2=1.275
r37 22 32 3.7489 $w=6.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.2 $Y=1.445 $X2=0.99
+ $Y2=1.445
r38 20 32 4.82002 $w=6.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.72 $Y=1.445
+ $X2=0.99 $Y2=1.445
r39 18 20 8.56892 $w=6.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.445
+ $X2=0.72 $Y2=1.445
r40 16 31 34.6051 $w=4.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.05 $Y=1.555
+ $X2=1.05 $Y2=1.275
r41 16 17 38.7081 $w=4.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.05 $Y=1.555
+ $X2=1.05 $Y2=1.78
r42 15 31 1.85385 $w=4.5e-07 $l=1.5e-08 $layer=POLY_cond $X=1.05 $Y=1.26
+ $X2=1.05 $Y2=1.275
r43 7 17 188.825 $w=2.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.15 $Y=2.54 $X2=1.15
+ $Y2=1.78
r44 1 15 24.7324 $w=4.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.08 $Y=1.11 $X2=1.08
+ $Y2=1.26
r45 1 11 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.26 $Y=1.11
+ $X2=1.26 $Y2=0.495
r46 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.9 $Y=1.11 $X2=0.9
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_LP%A_303_300# 1 2 7 9 13 17 21 23 24 26 29 30
+ 32 33 36 40 44 46 47
c89 13 0 1.69014e-19 $X=1.69 $Y=0.495
r90 46 47 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=3.057 $Y=2.19
+ $X2=3.057 $Y2=2.025
r91 42 44 3.67481 $w=2.52e-07 $l=1.19499e-07 $layer=LI1_cond $X=3.14 $Y=0.995
+ $X2=3.057 $Y2=0.91
r92 42 47 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.14 $Y=0.995
+ $X2=3.14 $Y2=2.025
r93 38 46 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=3.057 $Y=2.192
+ $X2=3.057 $Y2=2.19
r94 38 40 24.3561 $w=3.33e-07 $l=7.08e-07 $layer=LI1_cond $X=3.057 $Y=2.192
+ $X2=3.057 $Y2=2.9
r95 34 44 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=3.057 $Y=0.825
+ $X2=3.057 $Y2=0.91
r96 34 36 11.3524 $w=3.33e-07 $l=3.3e-07 $layer=LI1_cond $X=3.057 $Y=0.825
+ $X2=3.057 $Y2=0.495
r97 32 44 2.79892 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.89 $Y=0.91
+ $X2=3.057 $Y2=0.91
r98 32 33 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.89 $Y=0.91
+ $X2=2.305 $Y2=0.91
r99 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.14
+ $Y=1.335 $X2=2.14 $Y2=1.335
r100 27 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.14 $Y=0.995
+ $X2=2.305 $Y2=0.91
r101 27 29 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.14 $Y=0.995
+ $X2=2.14 $Y2=1.335
r102 25 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.14 $Y=1.32
+ $X2=2.14 $Y2=1.335
r103 25 26 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=2.14 $Y=1.32
+ $X2=2.14 $Y2=1.245
r104 19 26 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.05 $Y=1.17
+ $X2=2.14 $Y2=1.245
r105 19 21 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.05 $Y=1.17
+ $X2=2.05 $Y2=0.495
r106 18 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.245
+ $X2=1.69 $Y2=1.245
r107 17 26 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=1.245
+ $X2=2.14 $Y2=1.245
r108 17 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.975 $Y=1.245
+ $X2=1.765 $Y2=1.245
r109 15 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.32
+ $X2=1.69 $Y2=1.245
r110 15 23 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.69 $Y=1.32
+ $X2=1.69 $Y2=1.5
r111 11 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.17
+ $X2=1.69 $Y2=1.245
r112 11 13 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.69 $Y=1.17
+ $X2=1.69 $Y2=0.495
r113 7 23 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.64 $Y=1.625
+ $X2=1.64 $Y2=1.5
r114 7 9 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=1.64 $Y=1.625
+ $X2=1.64 $Y2=2.54
r115 2 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.915
+ $Y=2.045 $X2=3.055 $Y2=2.19
r116 2 40 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.915
+ $Y=2.045 $X2=3.055 $Y2=2.9
r117 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.285 $X2=3.055 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_LP%B_N 1 3 5 6 7 10 12 14 17 18 19 20 24 26
c49 5 0 1.57071e-19 $X=2.73 $Y=1.66
r50 24 26 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.34
+ $X2=2.73 $Y2=1.175
r51 19 20 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.7 $Y=1.295 $X2=2.7
+ $Y2=1.665
r52 19 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.71
+ $Y=1.34 $X2=2.71 $Y2=1.34
r53 15 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.84 $Y=0.93
+ $X2=2.84 $Y2=0.855
r54 15 26 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=2.84 $Y=0.93
+ $X2=2.84 $Y2=1.175
r55 12 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.84 $Y=0.78
+ $X2=2.84 $Y2=0.855
r56 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.84 $Y=0.78 $X2=2.84
+ $Y2=0.495
r57 10 17 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.79 $Y=2.545 $X2=2.79
+ $Y2=1.845
r58 6 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.765 $Y=0.855
+ $X2=2.84 $Y2=0.855
r59 6 7 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.765 $Y=0.855
+ $X2=2.555 $Y2=0.855
r60 5 17 34.9505 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.73 $Y=1.66
+ $X2=2.73 $Y2=1.845
r61 4 24 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=2.73 $Y=1.36 $X2=2.73
+ $Y2=1.34
r62 4 5 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=2.73 $Y=1.36 $X2=2.73
+ $Y2=1.66
r63 1 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.48 $Y=0.78
+ $X2=2.555 $Y2=0.855
r64 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.48 $Y=0.78 $X2=2.48
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_LP%VPWR 1 2 11 17 22 23 24 34 35 38
r29 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r31 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 29 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 28 31 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r35 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 26 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.05 $Y=3.33
+ $X2=0.885 $Y2=3.33
r37 26 28 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.05 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 24 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 22 31 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=3.33 $X2=2.16
+ $Y2=3.33
r41 22 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.525 $Y2=3.33
r42 21 34 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 21 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=2.525 $Y2=3.33
r44 17 20 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.525 $Y=2.19
+ $X2=2.525 $Y2=2.9
r45 15 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=3.33
r46 15 20 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=2.9
r47 11 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.885 $Y=2.185
+ $X2=0.885 $Y2=2.895
r48 9 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=3.245
+ $X2=0.885 $Y2=3.33
r49 9 14 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.885 $Y=3.245
+ $X2=0.885 $Y2=2.895
r50 2 20 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=2.045 $X2=2.525 $Y2=2.9
r51 2 17 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=2.045 $X2=2.525 $Y2=2.19
r52 1 14 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.74
+ $Y=2.04 $X2=0.885 $Y2=2.895
r53 1 11 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.74
+ $Y=2.04 $X2=0.885 $Y2=2.185
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_LP%Y 1 2 7 8 9 10 11 12 13 40 46
r38 46 47 3.94059 $w=5.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.817 $Y=2.035
+ $X2=1.817 $Y2=2.02
r39 31 50 2.06057 $w=5.03e-07 $l=8.7e-08 $layer=LI1_cond $X=1.817 $Y=2.272
+ $X2=1.817 $Y2=2.185
r40 13 37 2.84217 $w=5.03e-07 $l=1.2e-07 $layer=LI1_cond $X=1.817 $Y=2.775
+ $X2=1.817 $Y2=2.895
r41 12 13 8.76335 $w=5.03e-07 $l=3.7e-07 $layer=LI1_cond $X=1.817 $Y=2.405
+ $X2=1.817 $Y2=2.775
r42 12 31 3.15007 $w=5.03e-07 $l=1.33e-07 $layer=LI1_cond $X=1.817 $Y=2.405
+ $X2=1.817 $Y2=2.272
r43 11 50 2.72374 $w=5.03e-07 $l=1.15e-07 $layer=LI1_cond $X=1.817 $Y=2.07
+ $X2=1.817 $Y2=2.185
r44 11 46 0.828965 $w=5.03e-07 $l=3.5e-08 $layer=LI1_cond $X=1.817 $Y=2.07
+ $X2=1.817 $Y2=2.035
r45 11 47 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=1.985
+ $X2=1.68 $Y2=2.02
r46 10 11 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.985
r47 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=1.295
+ $X2=1.68 $Y2=1.665
r48 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=0.925 $X2=1.68
+ $Y2=1.295
r49 8 44 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=1.68 $Y=0.925 $X2=1.68
+ $Y2=0.725
r50 7 44 7.5165 $w=4.83e-07 $l=1.7e-07 $layer=LI1_cond $X=1.552 $Y=0.555
+ $X2=1.552 $Y2=0.725
r51 7 40 1.47968 $w=4.83e-07 $l=6e-08 $layer=LI1_cond $X=1.552 $Y=0.555
+ $X2=1.552 $Y2=0.495
r52 2 50 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=2.04 $X2=1.905 $Y2=2.185
r53 2 37 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=2.04 $X2=1.905 $Y2=2.895
r54 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.335
+ $Y=0.285 $X2=1.475 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r41 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.265
+ $Y2=0
r46 27 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=3.12
+ $Y2=0
r47 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=0 $X2=0.685
+ $Y2=0
r50 23 25 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.85 $Y=0 $X2=1.2
+ $Y2=0
r51 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=2.265
+ $Y2=0
r52 22 25 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=1.2 $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.52 $Y=0 $X2=0.685
+ $Y2=0
r56 17 19 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.52 $Y=0 $X2=0.24
+ $Y2=0
r57 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r58 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.265 $Y=0.085
+ $X2=2.265 $Y2=0
r60 11 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.265 $Y=0.085
+ $X2=2.265 $Y2=0.455
r61 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.085
+ $X2=0.685 $Y2=0
r62 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.685 $Y=0.085
+ $X2=0.685 $Y2=0.495
r63 2 13 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=2.125
+ $Y=0.285 $X2=2.265 $Y2=0.455
r64 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.54
+ $Y=0.285 $X2=0.685 $Y2=0.495
.ends

