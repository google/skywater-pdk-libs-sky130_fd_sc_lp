* NGSPICE file created from sky130_fd_sc_lp__dlybuf4s18kapwr_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlybuf4s18kapwr_1 A KAPWR VGND VNB VPB VPWR X
M1000 a_282_52# a_27_52# KAPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.65e+11p pd=2.53e+06u as=1.49e+12p ps=7.76e+06u
M1001 X a_394_52# KAPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1002 KAPWR a_282_52# a_394_52# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1003 a_282_52# a_27_52# VGND VNB nshort w=1e+06u l=180000u
+  ad=2.65e+11p pd=2.53e+06u as=1.2324e+12p ps=6.72e+06u
M1004 VGND A a_27_52# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 X a_394_52# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 VGND a_282_52# a_394_52# VNB nshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1007 KAPWR A a_27_52# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

