* File: sky130_fd_sc_lp__dlxtp_lp2.pxi.spice
* Created: Fri Aug 28 10:29:04 2020
* 
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%D N_D_c_138_n N_D_M1009_g N_D_M1004_g
+ N_D_M1002_g N_D_c_140_n N_D_c_141_n D D N_D_c_142_n N_D_c_143_n
+ PM_SKY130_FD_SC_LP__DLXTP_LP2%D
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%GATE N_GATE_c_181_n N_GATE_M1014_g
+ N_GATE_M1011_g N_GATE_c_176_n N_GATE_M1012_g N_GATE_c_182_n N_GATE_c_178_n
+ GATE GATE N_GATE_c_180_n PM_SKY130_FD_SC_LP__DLXTP_LP2%GATE
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%A_240_409# N_A_240_409#_M1012_d
+ N_A_240_409#_M1014_d N_A_240_409#_c_230_n N_A_240_409#_c_231_n
+ N_A_240_409#_c_232_n N_A_240_409#_M1013_g N_A_240_409#_M1017_g
+ N_A_240_409#_M1010_g N_A_240_409#_M1015_g N_A_240_409#_M1000_g
+ N_A_240_409#_c_246_n N_A_240_409#_c_236_n N_A_240_409#_c_247_n
+ N_A_240_409#_c_237_n N_A_240_409#_c_238_n N_A_240_409#_c_239_n
+ N_A_240_409#_c_240_n PM_SKY130_FD_SC_LP__DLXTP_LP2%A_240_409#
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%A_27_57# N_A_27_57#_M1009_s N_A_27_57#_M1004_s
+ N_A_27_57#_M1018_g N_A_27_57#_M1003_g N_A_27_57#_c_351_n N_A_27_57#_c_352_n
+ N_A_27_57#_c_353_n N_A_27_57#_c_362_n N_A_27_57#_c_354_n N_A_27_57#_c_355_n
+ N_A_27_57#_c_347_n N_A_27_57#_c_348_n N_A_27_57#_c_357_n N_A_27_57#_c_368_n
+ N_A_27_57#_c_349_n PM_SKY130_FD_SC_LP__DLXTP_LP2%A_27_57#
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%A_452_419# N_A_452_419#_M1017_s
+ N_A_452_419#_M1013_s N_A_452_419#_M1021_g N_A_452_419#_M1019_g
+ N_A_452_419#_c_449_n N_A_452_419#_c_438_n N_A_452_419#_c_439_n
+ N_A_452_419#_c_440_n N_A_452_419#_c_441_n N_A_452_419#_c_442_n
+ N_A_452_419#_c_443_n N_A_452_419#_c_444_n N_A_452_419#_c_445_n
+ N_A_452_419#_c_446_n N_A_452_419#_c_447_n
+ PM_SKY130_FD_SC_LP__DLXTP_LP2%A_452_419#
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%A_928_21# N_A_928_21#_M1001_d
+ N_A_928_21#_M1020_d N_A_928_21#_c_530_n N_A_928_21#_M1005_g
+ N_A_928_21#_c_531_n N_A_928_21#_c_532_n N_A_928_21#_M1016_g
+ N_A_928_21#_c_533_n N_A_928_21#_c_534_n N_A_928_21#_M1006_g
+ N_A_928_21#_M1007_g N_A_928_21#_M1008_g N_A_928_21#_c_538_n
+ N_A_928_21#_c_539_n N_A_928_21#_c_540_n N_A_928_21#_c_549_n
+ N_A_928_21#_c_550_n N_A_928_21#_c_541_n N_A_928_21#_c_542_n
+ N_A_928_21#_c_552_n N_A_928_21#_c_553_n N_A_928_21#_c_543_n
+ N_A_928_21#_c_544_n N_A_928_21#_c_545_n
+ PM_SKY130_FD_SC_LP__DLXTP_LP2%A_928_21#
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%A_778_47# N_A_778_47#_M1021_d
+ N_A_778_47#_M1015_d N_A_778_47#_M1022_g N_A_778_47#_M1020_g
+ N_A_778_47#_M1001_g N_A_778_47#_c_656_n N_A_778_47#_c_657_n
+ N_A_778_47#_c_668_n N_A_778_47#_c_665_n N_A_778_47#_c_658_n
+ N_A_778_47#_c_659_n N_A_778_47#_c_660_n N_A_778_47#_c_667_n
+ N_A_778_47#_c_661_n N_A_778_47#_c_662_n N_A_778_47#_c_663_n
+ PM_SKY130_FD_SC_LP__DLXTP_LP2%A_778_47#
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%VPWR N_VPWR_M1004_d N_VPWR_M1013_d
+ N_VPWR_M1016_d N_VPWR_M1007_s N_VPWR_c_760_n N_VPWR_c_761_n N_VPWR_c_762_n
+ VPWR N_VPWR_c_763_n N_VPWR_c_764_n N_VPWR_c_765_n N_VPWR_c_766_n
+ N_VPWR_c_759_n N_VPWR_c_768_n N_VPWR_c_769_n N_VPWR_c_770_n N_VPWR_c_771_n
+ PM_SKY130_FD_SC_LP__DLXTP_LP2%VPWR
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%Q N_Q_M1008_d N_Q_M1007_d Q Q Q Q Q Q Q
+ N_Q_c_839_n PM_SKY130_FD_SC_LP__DLXTP_LP2%Q
x_PM_SKY130_FD_SC_LP__DLXTP_LP2%VGND N_VGND_M1002_d N_VGND_M1010_d
+ N_VGND_M1005_d N_VGND_M1006_s N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n
+ N_VGND_c_861_n N_VGND_c_862_n VGND N_VGND_c_863_n N_VGND_c_864_n
+ N_VGND_c_865_n N_VGND_c_866_n N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n
+ N_VGND_c_870_n N_VGND_c_871_n PM_SKY130_FD_SC_LP__DLXTP_LP2%VGND
cc_1 VNB N_D_c_138_n 0.0326953f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.785
cc_2 VNB N_D_M1004_g 0.00525719f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_3 VNB N_D_c_140_n 0.022494f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.935
cc_4 VNB N_D_c_141_n 0.0177981f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.575
cc_5 VNB N_D_c_142_n 0.0356897f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.07
cc_6 VNB N_D_c_143_n 0.00623391f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.07
cc_7 VNB N_GATE_M1011_g 0.0343644f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_8 VNB N_GATE_c_176_n 0.0284486f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.785
cc_9 VNB N_GATE_M1012_g 0.0408324f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.785
cc_10 VNB N_GATE_c_178_n 0.0126107f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB GATE 0.00224742f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_12 VNB N_GATE_c_180_n 0.0264205f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.07
cc_13 VNB N_A_240_409#_c_230_n 0.0222696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_240_409#_c_231_n 0.0118098f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.785
cc_15 VNB N_A_240_409#_c_232_n 0.0392982f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_16 VNB N_A_240_409#_M1017_g 0.0480031f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.575
cc_17 VNB N_A_240_409#_M1010_g 0.0382859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_240_409#_M1000_g 0.0516381f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.665
cc_19 VNB N_A_240_409#_c_236_n 0.01887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_240_409#_c_237_n 0.0275078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_240_409#_c_238_n 3.73352e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_240_409#_c_239_n 0.00186136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_240_409#_c_240_n 0.0296477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_57#_M1018_g 0.0645408f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_25 VNB N_A_27_57#_c_347_n 0.0251105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_57#_c_348_n 0.0434461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_57#_c_349_n 0.0138264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_452_419#_c_438_n 0.00720411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_452_419#_c_439_n 0.00645886f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.07
cc_30 VNB N_A_452_419#_c_440_n 0.0145351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_452_419#_c_441_n 0.00174403f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.665
cc_32 VNB N_A_452_419#_c_442_n 0.0320358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_452_419#_c_443_n 0.00237049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_452_419#_c_444_n 0.0357886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_452_419#_c_445_n 0.00223764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_452_419#_c_446_n 0.0242336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_452_419#_c_447_n 0.0169948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_928_21#_c_530_n 0.0173894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_928_21#_c_531_n 0.0389097f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_40 VNB N_A_928_21#_c_532_n 0.00672488f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=0.935
cc_41 VNB N_A_928_21#_c_533_n 0.0138477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_928_21#_c_534_n 0.0173885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_928_21#_M1006_g 0.0233771f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.07
cc_44 VNB N_A_928_21#_M1007_g 0.0337887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_928_21#_M1008_g 0.0244697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_928_21#_c_538_n 0.02068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_928_21#_c_539_n 0.00251773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_928_21#_c_540_n 0.0465721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_928_21#_c_541_n 0.008013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_928_21#_c_542_n 0.0201442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_928_21#_c_543_n 0.0038902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_928_21#_c_544_n 0.0311384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_928_21#_c_545_n 0.0224001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_778_47#_M1022_g 0.0245479f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_55 VNB N_A_778_47#_M1020_g 0.00897645f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.935
cc_56 VNB N_A_778_47#_M1001_g 0.0232686f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_57 VNB N_A_778_47#_c_656_n 0.0257202f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.07
cc_58 VNB N_A_778_47#_c_657_n 0.0147077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_778_47#_c_658_n 0.00174008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_778_47#_c_659_n 0.00412328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_778_47#_c_660_n 0.0176878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_778_47#_c_661_n 0.00115699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_778_47#_c_662_n 0.001548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_778_47#_c_663_n 0.0290391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VPWR_c_759_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB Q 0.0454498f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.785
cc_67 VNB N_Q_c_839_n 0.0166981f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.07
cc_68 VNB N_VGND_c_858_n 0.00833355f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.575
cc_69 VNB N_VGND_c_859_n 0.0495794f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_70 VNB N_VGND_c_860_n 0.00345358f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.07
cc_71 VNB N_VGND_c_861_n 0.00884771f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.295
cc_72 VNB N_VGND_c_862_n 0.01602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_863_n 0.0271986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_864_n 0.0524784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_865_n 0.0347785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_866_n 0.0267209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_867_n 0.439831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_868_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_869_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_870_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_871_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VPB N_D_M1004_g 0.0463329f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_83 VPB N_D_c_143_n 0.0036938f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.07
cc_84 VPB N_GATE_c_181_n 0.0236547f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.785
cc_85 VPB N_GATE_c_182_n 0.0327043f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.388
cc_86 VPB GATE 0.00171359f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_87 VPB N_GATE_c_180_n 0.00188746f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.07
cc_88 VPB N_A_240_409#_c_230_n 0.0175592f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_240_409#_c_231_n 0.00562653f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.785
cc_90 VPB N_A_240_409#_c_232_n 0.0328072f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.495
cc_91 VPB N_A_240_409#_M1013_g 0.0330542f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=0.935
cc_92 VPB N_A_240_409#_M1015_g 0.0427369f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.07
cc_93 VPB N_A_240_409#_c_246_n 0.0211551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_240_409#_c_247_n 0.0512543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_240_409#_c_238_n 0.0048479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_240_409#_c_239_n 0.00105578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_240_409#_c_240_n 0.00295026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_27_57#_M1003_g 0.0295061f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.935
cc_99 VPB N_A_27_57#_c_351_n 0.00998646f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_27_57#_c_352_n 0.0118411f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.07
cc_101 VPB N_A_27_57#_c_353_n 0.0189994f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.07
cc_102 VPB N_A_27_57#_c_354_n 0.0266693f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.665
cc_103 VPB N_A_27_57#_c_355_n 0.00227719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_27_57#_c_348_n 0.0175744f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_27_57#_c_357_n 0.00704942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_27_57#_c_349_n 0.0327118f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_452_419#_M1019_g 0.0288285f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.785
cc_108 VPB N_A_452_419#_c_449_n 0.0141455f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.575
cc_109 VPB N_A_452_419#_c_439_n 0.00945331f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.07
cc_110 VPB N_A_452_419#_c_444_n 0.00535196f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_928_21#_M1016_g 0.0309863f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_112 VPB N_A_928_21#_M1007_g 0.040962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_928_21#_c_540_n 0.0239791f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_928_21#_c_549_n 0.022477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_928_21#_c_550_n 0.00242083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_928_21#_c_542_n 0.0197449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_928_21#_c_552_n 0.0169982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_928_21#_c_553_n 0.00524078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_928_21#_c_544_n 0.0127871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_778_47#_M1020_g 0.0508229f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.935
cc_121 VPB N_A_778_47#_c_665_n 0.00479404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_778_47#_c_659_n 0.00319282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_778_47#_c_667_n 0.00935447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_760_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_125 VPB N_VPWR_c_761_n 0.00537225f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.07
cc_126 VPB N_VPWR_c_762_n 0.0333348f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.665
cc_127 VPB N_VPWR_c_763_n 0.0497246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_764_n 0.0645029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_765_n 0.0339021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_766_n 0.0266596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_759_n 0.0848832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_768_n 0.0231183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_769_n 0.0112407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_770_n 0.00513801f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_771_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB Q 0.0702779f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.785
cc_137 N_D_c_138_n N_GATE_M1011_g 0.0193566f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_138 N_D_c_142_n N_GATE_M1011_g 0.00589521f $X=0.63 $Y=1.07 $X2=0 $Y2=0
cc_139 N_D_c_143_n N_GATE_M1011_g 0.00493178f $X=0.63 $Y=1.07 $X2=0 $Y2=0
cc_140 N_D_M1004_g N_GATE_c_182_n 0.0469034f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_141 N_D_c_142_n N_GATE_c_178_n 0.0100071f $X=0.63 $Y=1.07 $X2=0 $Y2=0
cc_142 N_D_c_143_n N_GATE_c_178_n 0.00421358f $X=0.63 $Y=1.07 $X2=0 $Y2=0
cc_143 N_D_M1004_g GATE 6.08032e-19 $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_144 N_D_c_142_n GATE 4.75068e-19 $X=0.63 $Y=1.07 $X2=0 $Y2=0
cc_145 N_D_c_143_n GATE 0.0404826f $X=0.63 $Y=1.07 $X2=0 $Y2=0
cc_146 N_D_M1004_g N_GATE_c_180_n 0.00810991f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_147 N_D_c_141_n N_GATE_c_180_n 0.0100071f $X=0.607 $Y=1.575 $X2=0 $Y2=0
cc_148 N_D_M1004_g N_A_240_409#_c_246_n 0.0010579f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_149 N_D_M1004_g N_A_27_57#_c_351_n 0.00533154f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_150 N_D_M1004_g N_A_27_57#_c_352_n 0.00497631f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_151 N_D_M1004_g N_A_27_57#_c_353_n 0.00855612f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_152 N_D_M1004_g N_A_27_57#_c_362_n 0.0175147f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_153 N_D_c_143_n N_A_27_57#_c_362_n 0.00917312f $X=0.63 $Y=1.07 $X2=0 $Y2=0
cc_154 N_D_c_138_n N_A_27_57#_c_347_n 0.0113742f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_155 N_D_c_138_n N_A_27_57#_c_348_n 0.0333303f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_156 N_D_c_143_n N_A_27_57#_c_348_n 0.0634302f $X=0.63 $Y=1.07 $X2=0 $Y2=0
cc_157 N_D_M1004_g N_A_27_57#_c_357_n 3.84191e-19 $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_158 N_D_M1004_g N_A_27_57#_c_368_n 5.33974e-19 $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_159 N_D_M1004_g N_VPWR_c_760_n 0.00983558f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_160 N_D_M1004_g N_VPWR_c_759_n 0.00762765f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_161 N_D_M1004_g N_VPWR_c_768_n 0.00580736f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_162 N_D_c_138_n N_VGND_c_858_n 0.0153894f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_163 N_D_c_138_n N_VGND_c_863_n 0.00947719f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_164 N_D_c_138_n N_VGND_c_867_n 0.0180243f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_165 N_D_c_140_n N_VGND_c_867_n 7.9244e-19 $X=0.675 $Y=0.935 $X2=0 $Y2=0
cc_166 N_GATE_c_176_n N_A_240_409#_c_231_n 0.00116165f $X=1.57 $Y=1.25 $X2=0
+ $Y2=0
cc_167 GATE N_A_240_409#_c_231_n 0.00106029f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_168 N_GATE_c_180_n N_A_240_409#_c_231_n 0.00460354f $X=1.215 $Y=1.34 $X2=0
+ $Y2=0
cc_169 N_GATE_c_181_n N_A_240_409#_c_246_n 0.0064589f $X=1.075 $Y=1.97 $X2=0
+ $Y2=0
cc_170 N_GATE_c_182_n N_A_240_409#_c_246_n 0.00126755f $X=1.215 $Y=1.68 $X2=0
+ $Y2=0
cc_171 GATE N_A_240_409#_c_246_n 0.0159377f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_172 N_GATE_M1011_g N_A_240_409#_c_236_n 0.00350406f $X=1.285 $Y=0.495 $X2=0
+ $Y2=0
cc_173 N_GATE_c_176_n N_A_240_409#_c_236_n 0.0066104f $X=1.57 $Y=1.25 $X2=0
+ $Y2=0
cc_174 N_GATE_M1012_g N_A_240_409#_c_236_n 0.0258005f $X=1.645 $Y=0.495 $X2=0
+ $Y2=0
cc_175 N_GATE_c_182_n N_A_240_409#_c_236_n 0.00102978f $X=1.215 $Y=1.68 $X2=0
+ $Y2=0
cc_176 GATE N_A_240_409#_c_236_n 0.0318088f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_177 N_GATE_c_180_n N_A_240_409#_c_236_n 0.00674633f $X=1.215 $Y=1.34 $X2=0
+ $Y2=0
cc_178 N_GATE_c_182_n N_A_240_409#_c_247_n 0.0121824f $X=1.215 $Y=1.68 $X2=0
+ $Y2=0
cc_179 N_GATE_c_181_n N_A_27_57#_c_352_n 0.00184553f $X=1.075 $Y=1.97 $X2=0
+ $Y2=0
cc_180 N_GATE_c_181_n N_A_27_57#_c_353_n 6.30887e-19 $X=1.075 $Y=1.97 $X2=0
+ $Y2=0
cc_181 N_GATE_c_181_n N_A_27_57#_c_362_n 0.0175989f $X=1.075 $Y=1.97 $X2=0 $Y2=0
cc_182 GATE N_A_27_57#_c_362_n 0.00273719f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_183 N_GATE_c_181_n N_A_27_57#_c_354_n 9.86509e-19 $X=1.075 $Y=1.97 $X2=0
+ $Y2=0
cc_184 N_GATE_c_181_n N_A_27_57#_c_368_n 0.0107217f $X=1.075 $Y=1.97 $X2=0 $Y2=0
cc_185 GATE N_A_27_57#_c_368_n 5.215e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_186 N_GATE_M1012_g N_A_452_419#_c_438_n 0.0016802f $X=1.645 $Y=0.495 $X2=0
+ $Y2=0
cc_187 N_GATE_M1012_g N_A_452_419#_c_439_n 9.23893e-19 $X=1.645 $Y=0.495 $X2=0
+ $Y2=0
cc_188 N_GATE_M1012_g N_A_452_419#_c_445_n 7.2158e-19 $X=1.645 $Y=0.495 $X2=0
+ $Y2=0
cc_189 N_GATE_c_181_n N_VPWR_c_760_n 0.0168697f $X=1.075 $Y=1.97 $X2=0 $Y2=0
cc_190 N_GATE_c_181_n N_VPWR_c_763_n 0.00586345f $X=1.075 $Y=1.97 $X2=0 $Y2=0
cc_191 N_GATE_c_181_n N_VPWR_c_759_n 0.00791681f $X=1.075 $Y=1.97 $X2=0 $Y2=0
cc_192 N_GATE_M1011_g N_VGND_c_858_n 0.0127712f $X=1.285 $Y=0.495 $X2=0 $Y2=0
cc_193 N_GATE_M1012_g N_VGND_c_858_n 0.002112f $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_194 N_GATE_c_178_n N_VGND_c_858_n 0.00108472f $X=1.215 $Y=1.25 $X2=0 $Y2=0
cc_195 GATE N_VGND_c_858_n 0.0077292f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_196 N_GATE_M1011_g N_VGND_c_859_n 0.00445056f $X=1.285 $Y=0.495 $X2=0 $Y2=0
cc_197 N_GATE_M1012_g N_VGND_c_859_n 0.00502664f $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_198 N_GATE_M1011_g N_VGND_c_867_n 0.00796275f $X=1.285 $Y=0.495 $X2=0 $Y2=0
cc_199 N_GATE_M1012_g N_VGND_c_867_n 0.010303f $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_200 N_A_240_409#_c_232_n N_A_27_57#_M1018_g 0.0168139f $X=2.67 $Y=1.935 $X2=0
+ $Y2=0
cc_201 N_A_240_409#_M1010_g N_A_27_57#_M1018_g 0.0366025f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_202 N_A_240_409#_c_237_n N_A_27_57#_M1018_g 0.0119529f $X=4.07 $Y=1.35 $X2=0
+ $Y2=0
cc_203 N_A_240_409#_c_238_n N_A_27_57#_M1018_g 0.00106764f $X=2.915 $Y=1.43
+ $X2=0 $Y2=0
cc_204 N_A_240_409#_c_239_n N_A_27_57#_M1018_g 0.00106741f $X=4.235 $Y=1.35
+ $X2=0 $Y2=0
cc_205 N_A_240_409#_c_240_n N_A_27_57#_M1018_g 0.0054193f $X=4.235 $Y=1.5 $X2=0
+ $Y2=0
cc_206 N_A_240_409#_M1015_g N_A_27_57#_M1003_g 0.0464877f $X=4.195 $Y=2.595
+ $X2=0 $Y2=0
cc_207 N_A_240_409#_M1014_d N_A_27_57#_c_354_n 0.00621637f $X=1.2 $Y=2.045 $X2=0
+ $Y2=0
cc_208 N_A_240_409#_c_232_n N_A_27_57#_c_354_n 0.00120194f $X=2.67 $Y=1.935
+ $X2=0 $Y2=0
cc_209 N_A_240_409#_M1013_g N_A_27_57#_c_354_n 0.0270548f $X=2.67 $Y=2.595 $X2=0
+ $Y2=0
cc_210 N_A_240_409#_M1015_g N_A_27_57#_c_354_n 4.99054e-19 $X=4.195 $Y=2.595
+ $X2=0 $Y2=0
cc_211 N_A_240_409#_c_246_n N_A_27_57#_c_354_n 0.0351957f $X=1.695 $Y=2.15 $X2=0
+ $Y2=0
cc_212 N_A_240_409#_c_247_n N_A_27_57#_c_354_n 0.00202888f $X=1.86 $Y=1.77 $X2=0
+ $Y2=0
cc_213 N_A_240_409#_c_238_n N_A_27_57#_c_354_n 0.00799373f $X=2.915 $Y=1.43
+ $X2=0 $Y2=0
cc_214 N_A_240_409#_c_232_n N_A_27_57#_c_355_n 0.00132466f $X=2.67 $Y=1.935
+ $X2=0 $Y2=0
cc_215 N_A_240_409#_M1013_g N_A_27_57#_c_355_n 0.0175426f $X=2.67 $Y=2.595 $X2=0
+ $Y2=0
cc_216 N_A_240_409#_c_237_n N_A_27_57#_c_355_n 0.0245309f $X=4.07 $Y=1.35 $X2=0
+ $Y2=0
cc_217 N_A_240_409#_c_238_n N_A_27_57#_c_355_n 0.0182306f $X=2.915 $Y=1.43 $X2=0
+ $Y2=0
cc_218 N_A_240_409#_c_239_n N_A_27_57#_c_355_n 0.00180728f $X=4.235 $Y=1.35
+ $X2=0 $Y2=0
cc_219 N_A_240_409#_c_240_n N_A_27_57#_c_355_n 0.00356088f $X=4.235 $Y=1.5 $X2=0
+ $Y2=0
cc_220 N_A_240_409#_M1014_d N_A_27_57#_c_368_n 0.00727888f $X=1.2 $Y=2.045 $X2=0
+ $Y2=0
cc_221 N_A_240_409#_c_246_n N_A_27_57#_c_368_n 0.00674878f $X=1.695 $Y=2.15
+ $X2=0 $Y2=0
cc_222 N_A_240_409#_c_232_n N_A_27_57#_c_349_n 0.0185824f $X=2.67 $Y=1.935 $X2=0
+ $Y2=0
cc_223 N_A_240_409#_c_237_n N_A_27_57#_c_349_n 0.00989014f $X=4.07 $Y=1.35 $X2=0
+ $Y2=0
cc_224 N_A_240_409#_c_238_n N_A_27_57#_c_349_n 0.00135255f $X=2.915 $Y=1.43
+ $X2=0 $Y2=0
cc_225 N_A_240_409#_c_239_n N_A_27_57#_c_349_n 2.9337e-19 $X=4.235 $Y=1.35 $X2=0
+ $Y2=0
cc_226 N_A_240_409#_c_240_n N_A_27_57#_c_349_n 0.0464877f $X=4.235 $Y=1.5 $X2=0
+ $Y2=0
cc_227 N_A_240_409#_M1017_g N_A_452_419#_c_438_n 0.0163907f $X=2.635 $Y=0.445
+ $X2=0 $Y2=0
cc_228 N_A_240_409#_M1010_g N_A_452_419#_c_438_n 0.00231534f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_229 N_A_240_409#_c_236_n N_A_452_419#_c_438_n 0.0460377f $X=1.86 $Y=0.495
+ $X2=0 $Y2=0
cc_230 N_A_240_409#_c_230_n N_A_452_419#_c_439_n 0.0191052f $X=2.545 $Y=1.68
+ $X2=0 $Y2=0
cc_231 N_A_240_409#_c_232_n N_A_452_419#_c_439_n 0.0207447f $X=2.67 $Y=1.935
+ $X2=0 $Y2=0
cc_232 N_A_240_409#_M1013_g N_A_452_419#_c_439_n 0.0236068f $X=2.67 $Y=2.595
+ $X2=0 $Y2=0
cc_233 N_A_240_409#_M1017_g N_A_452_419#_c_439_n 0.00652566f $X=2.635 $Y=0.445
+ $X2=0 $Y2=0
cc_234 N_A_240_409#_M1010_g N_A_452_419#_c_439_n 8.67864e-19 $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_235 N_A_240_409#_c_246_n N_A_452_419#_c_439_n 0.0175733f $X=1.695 $Y=2.15
+ $X2=0 $Y2=0
cc_236 N_A_240_409#_c_236_n N_A_452_419#_c_439_n 0.0638949f $X=1.86 $Y=0.495
+ $X2=0 $Y2=0
cc_237 N_A_240_409#_c_247_n N_A_452_419#_c_439_n 0.00352861f $X=1.86 $Y=1.77
+ $X2=0 $Y2=0
cc_238 N_A_240_409#_c_238_n N_A_452_419#_c_439_n 0.0487642f $X=2.915 $Y=1.43
+ $X2=0 $Y2=0
cc_239 N_A_240_409#_M1000_g N_A_452_419#_c_440_n 0.0173733f $X=4.325 $Y=0.445
+ $X2=0 $Y2=0
cc_240 N_A_240_409#_c_239_n N_A_452_419#_c_440_n 0.0254231f $X=4.235 $Y=1.35
+ $X2=0 $Y2=0
cc_241 N_A_240_409#_c_240_n N_A_452_419#_c_440_n 0.00108118f $X=4.235 $Y=1.5
+ $X2=0 $Y2=0
cc_242 N_A_240_409#_M1000_g N_A_452_419#_c_442_n 0.0213634f $X=4.325 $Y=0.445
+ $X2=0 $Y2=0
cc_243 N_A_240_409#_c_237_n N_A_452_419#_c_442_n 0.00616629f $X=4.07 $Y=1.35
+ $X2=0 $Y2=0
cc_244 N_A_240_409#_M1015_g N_A_452_419#_c_443_n 0.00150575f $X=4.195 $Y=2.595
+ $X2=0 $Y2=0
cc_245 N_A_240_409#_M1000_g N_A_452_419#_c_443_n 0.00646079f $X=4.325 $Y=0.445
+ $X2=0 $Y2=0
cc_246 N_A_240_409#_c_239_n N_A_452_419#_c_443_n 0.024934f $X=4.235 $Y=1.35
+ $X2=0 $Y2=0
cc_247 N_A_240_409#_M1015_g N_A_452_419#_c_444_n 0.0393409f $X=4.195 $Y=2.595
+ $X2=0 $Y2=0
cc_248 N_A_240_409#_M1000_g N_A_452_419#_c_444_n 0.0266774f $X=4.325 $Y=0.445
+ $X2=0 $Y2=0
cc_249 N_A_240_409#_c_239_n N_A_452_419#_c_444_n 0.00139253f $X=4.235 $Y=1.35
+ $X2=0 $Y2=0
cc_250 N_A_240_409#_M1017_g N_A_452_419#_c_445_n 0.0046518f $X=2.635 $Y=0.445
+ $X2=0 $Y2=0
cc_251 N_A_240_409#_c_236_n N_A_452_419#_c_445_n 0.0127463f $X=1.86 $Y=0.495
+ $X2=0 $Y2=0
cc_252 N_A_240_409#_c_232_n N_A_452_419#_c_446_n 2.75182e-19 $X=2.67 $Y=1.935
+ $X2=0 $Y2=0
cc_253 N_A_240_409#_M1017_g N_A_452_419#_c_446_n 0.0144626f $X=2.635 $Y=0.445
+ $X2=0 $Y2=0
cc_254 N_A_240_409#_M1010_g N_A_452_419#_c_446_n 0.0139129f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_255 N_A_240_409#_c_237_n N_A_452_419#_c_446_n 0.0703f $X=4.07 $Y=1.35 $X2=0
+ $Y2=0
cc_256 N_A_240_409#_c_238_n N_A_452_419#_c_446_n 0.0246567f $X=2.915 $Y=1.43
+ $X2=0 $Y2=0
cc_257 N_A_240_409#_M1000_g N_A_452_419#_c_447_n 0.0167095f $X=4.325 $Y=0.445
+ $X2=0 $Y2=0
cc_258 N_A_240_409#_M1000_g N_A_928_21#_c_530_n 0.0437277f $X=4.325 $Y=0.445
+ $X2=0 $Y2=0
cc_259 N_A_240_409#_M1000_g N_A_778_47#_c_668_n 0.0106725f $X=4.325 $Y=0.445
+ $X2=0 $Y2=0
cc_260 N_A_240_409#_M1000_g N_A_778_47#_c_659_n 3.07502e-19 $X=4.325 $Y=0.445
+ $X2=0 $Y2=0
cc_261 N_A_240_409#_M1015_g N_A_778_47#_c_667_n 0.024011f $X=4.195 $Y=2.595
+ $X2=0 $Y2=0
cc_262 N_A_240_409#_c_239_n N_A_778_47#_c_667_n 0.00410784f $X=4.235 $Y=1.35
+ $X2=0 $Y2=0
cc_263 N_A_240_409#_c_240_n N_A_778_47#_c_667_n 5.49786e-19 $X=4.235 $Y=1.5
+ $X2=0 $Y2=0
cc_264 N_A_240_409#_M1000_g N_A_778_47#_c_661_n 4.6246e-19 $X=4.325 $Y=0.445
+ $X2=0 $Y2=0
cc_265 N_A_240_409#_M1013_g N_VPWR_c_763_n 0.00693303f $X=2.67 $Y=2.595 $X2=0
+ $Y2=0
cc_266 N_A_240_409#_M1015_g N_VPWR_c_764_n 0.00954582f $X=4.195 $Y=2.595 $X2=0
+ $Y2=0
cc_267 N_A_240_409#_M1013_g N_VPWR_c_759_n 0.0113938f $X=2.67 $Y=2.595 $X2=0
+ $Y2=0
cc_268 N_A_240_409#_M1015_g N_VPWR_c_759_n 0.0165468f $X=4.195 $Y=2.595 $X2=0
+ $Y2=0
cc_269 N_A_240_409#_M1013_g N_VPWR_c_769_n 0.00812485f $X=2.67 $Y=2.595 $X2=0
+ $Y2=0
cc_270 N_A_240_409#_c_236_n N_VGND_c_858_n 0.0153904f $X=1.86 $Y=0.495 $X2=0
+ $Y2=0
cc_271 N_A_240_409#_M1017_g N_VGND_c_859_n 0.00549284f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_272 N_A_240_409#_M1010_g N_VGND_c_859_n 0.00486043f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_273 N_A_240_409#_c_236_n N_VGND_c_859_n 0.0220321f $X=1.86 $Y=0.495 $X2=0
+ $Y2=0
cc_274 N_A_240_409#_M1017_g N_VGND_c_860_n 0.00239794f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_275 N_A_240_409#_M1010_g N_VGND_c_860_n 0.0128479f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_276 N_A_240_409#_M1000_g N_VGND_c_864_n 0.00366111f $X=4.325 $Y=0.445 $X2=0
+ $Y2=0
cc_277 N_A_240_409#_M1017_g N_VGND_c_867_n 0.0112805f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_278 N_A_240_409#_M1010_g N_VGND_c_867_n 0.00814425f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_279 N_A_240_409#_M1000_g N_VGND_c_867_n 0.00548904f $X=4.325 $Y=0.445 $X2=0
+ $Y2=0
cc_280 N_A_240_409#_c_236_n N_VGND_c_867_n 0.0125808f $X=1.86 $Y=0.495 $X2=0
+ $Y2=0
cc_281 N_A_27_57#_c_354_n N_A_452_419#_M1013_s 0.0071475f $X=3.32 $Y=2.67 $X2=0
+ $Y2=0
cc_282 N_A_27_57#_c_354_n N_A_452_419#_c_439_n 0.02102f $X=3.32 $Y=2.67 $X2=0
+ $Y2=0
cc_283 N_A_27_57#_M1018_g N_A_452_419#_c_441_n 9.83442e-19 $X=3.425 $Y=0.445
+ $X2=0 $Y2=0
cc_284 N_A_27_57#_M1018_g N_A_452_419#_c_442_n 0.0206263f $X=3.425 $Y=0.445
+ $X2=0 $Y2=0
cc_285 N_A_27_57#_c_349_n N_A_452_419#_c_442_n 0.00218158f $X=3.705 $Y=1.77
+ $X2=0 $Y2=0
cc_286 N_A_27_57#_M1018_g N_A_452_419#_c_446_n 0.013919f $X=3.425 $Y=0.445 $X2=0
+ $Y2=0
cc_287 N_A_27_57#_M1018_g N_A_452_419#_c_447_n 0.0353429f $X=3.425 $Y=0.445
+ $X2=0 $Y2=0
cc_288 N_A_27_57#_M1003_g N_A_778_47#_c_667_n 0.00311375f $X=3.705 $Y=2.595
+ $X2=0 $Y2=0
cc_289 N_A_27_57#_c_354_n N_A_778_47#_c_667_n 0.00438731f $X=3.32 $Y=2.67 $X2=0
+ $Y2=0
cc_290 N_A_27_57#_c_355_n N_A_778_47#_c_667_n 0.0126395f $X=3.485 $Y=1.77 $X2=0
+ $Y2=0
cc_291 N_A_27_57#_c_362_n N_VPWR_M1004_d 0.00627257f $X=1.155 $Y=2.54 $X2=-0.19
+ $Y2=-0.245
cc_292 N_A_27_57#_c_354_n N_VPWR_M1013_d 0.0262573f $X=3.32 $Y=2.67 $X2=0 $Y2=0
cc_293 N_A_27_57#_c_355_n N_VPWR_M1013_d 0.0103916f $X=3.485 $Y=1.77 $X2=0 $Y2=0
cc_294 N_A_27_57#_c_353_n N_VPWR_c_760_n 0.0171316f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_295 N_A_27_57#_c_362_n N_VPWR_c_760_n 0.0155262f $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_296 N_A_27_57#_c_362_n N_VPWR_c_763_n 0.00250321f $X=1.155 $Y=2.54 $X2=0
+ $Y2=0
cc_297 N_A_27_57#_c_354_n N_VPWR_c_763_n 0.0299159f $X=3.32 $Y=2.67 $X2=0 $Y2=0
cc_298 N_A_27_57#_c_368_n N_VPWR_c_763_n 0.00291601f $X=1.24 $Y=2.54 $X2=0 $Y2=0
cc_299 N_A_27_57#_M1003_g N_VPWR_c_764_n 0.00896513f $X=3.705 $Y=2.595 $X2=0
+ $Y2=0
cc_300 N_A_27_57#_c_354_n N_VPWR_c_764_n 0.00935983f $X=3.32 $Y=2.67 $X2=0 $Y2=0
cc_301 N_A_27_57#_M1003_g N_VPWR_c_759_n 0.0161276f $X=3.705 $Y=2.595 $X2=0
+ $Y2=0
cc_302 N_A_27_57#_c_353_n N_VPWR_c_759_n 0.0125808f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_303 N_A_27_57#_c_362_n N_VPWR_c_759_n 0.00975551f $X=1.155 $Y=2.54 $X2=0
+ $Y2=0
cc_304 N_A_27_57#_c_354_n N_VPWR_c_759_n 0.0603989f $X=3.32 $Y=2.67 $X2=0 $Y2=0
cc_305 N_A_27_57#_c_368_n N_VPWR_c_759_n 0.00492279f $X=1.24 $Y=2.54 $X2=0 $Y2=0
cc_306 N_A_27_57#_c_353_n N_VPWR_c_768_n 0.0220321f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_307 N_A_27_57#_c_362_n N_VPWR_c_768_n 0.00277646f $X=1.155 $Y=2.54 $X2=0
+ $Y2=0
cc_308 N_A_27_57#_M1003_g N_VPWR_c_769_n 0.00732785f $X=3.705 $Y=2.595 $X2=0
+ $Y2=0
cc_309 N_A_27_57#_c_354_n N_VPWR_c_769_n 0.0231925f $X=3.32 $Y=2.67 $X2=0 $Y2=0
cc_310 N_A_27_57#_c_347_n N_VGND_c_858_n 0.0153904f $X=0.28 $Y=0.495 $X2=0 $Y2=0
cc_311 N_A_27_57#_M1018_g N_VGND_c_860_n 0.0136303f $X=3.425 $Y=0.445 $X2=0
+ $Y2=0
cc_312 N_A_27_57#_c_347_n N_VGND_c_863_n 0.0217285f $X=0.28 $Y=0.495 $X2=0 $Y2=0
cc_313 N_A_27_57#_M1018_g N_VGND_c_864_n 0.00486043f $X=3.425 $Y=0.445 $X2=0
+ $Y2=0
cc_314 N_A_27_57#_M1018_g N_VGND_c_867_n 0.00827383f $X=3.425 $Y=0.445 $X2=0
+ $Y2=0
cc_315 N_A_27_57#_c_347_n N_VGND_c_867_n 0.0125175f $X=0.28 $Y=0.495 $X2=0 $Y2=0
cc_316 N_A_452_419#_c_440_n N_A_928_21#_c_531_n 0.00443311f $X=4.61 $Y=0.925
+ $X2=0 $Y2=0
cc_317 N_A_452_419#_c_440_n N_A_928_21#_c_532_n 0.00716998f $X=4.61 $Y=0.925
+ $X2=0 $Y2=0
cc_318 N_A_452_419#_c_444_n N_A_928_21#_c_532_n 0.0108565f $X=4.775 $Y=1.39
+ $X2=0 $Y2=0
cc_319 N_A_452_419#_M1019_g N_A_928_21#_M1016_g 0.0520244f $X=4.735 $Y=2.595
+ $X2=0 $Y2=0
cc_320 N_A_452_419#_c_449_n N_A_928_21#_M1016_g 0.0175277f $X=4.775 $Y=1.895
+ $X2=0 $Y2=0
cc_321 N_A_452_419#_c_443_n N_A_928_21#_c_540_n 6.18803e-19 $X=4.775 $Y=1.39
+ $X2=0 $Y2=0
cc_322 N_A_452_419#_c_444_n N_A_928_21#_c_540_n 0.0175277f $X=4.775 $Y=1.39
+ $X2=0 $Y2=0
cc_323 N_A_452_419#_c_440_n N_A_928_21#_c_545_n 0.00122954f $X=4.61 $Y=0.925
+ $X2=0 $Y2=0
cc_324 N_A_452_419#_c_443_n N_A_928_21#_c_545_n 7.57295e-19 $X=4.775 $Y=1.39
+ $X2=0 $Y2=0
cc_325 N_A_452_419#_c_440_n N_A_778_47#_c_668_n 0.0594098f $X=4.61 $Y=0.925
+ $X2=0 $Y2=0
cc_326 N_A_452_419#_c_442_n N_A_778_47#_c_668_n 0.00213932f $X=3.875 $Y=0.93
+ $X2=0 $Y2=0
cc_327 N_A_452_419#_M1019_g N_A_778_47#_c_665_n 0.0188025f $X=4.735 $Y=2.595
+ $X2=0 $Y2=0
cc_328 N_A_452_419#_c_449_n N_A_778_47#_c_665_n 0.00261165f $X=4.775 $Y=1.895
+ $X2=0 $Y2=0
cc_329 N_A_452_419#_c_443_n N_A_778_47#_c_665_n 0.0177883f $X=4.775 $Y=1.39
+ $X2=0 $Y2=0
cc_330 N_A_452_419#_c_440_n N_A_778_47#_c_658_n 0.00651431f $X=4.61 $Y=0.925
+ $X2=0 $Y2=0
cc_331 N_A_452_419#_M1019_g N_A_778_47#_c_659_n 0.00371872f $X=4.735 $Y=2.595
+ $X2=0 $Y2=0
cc_332 N_A_452_419#_c_440_n N_A_778_47#_c_659_n 0.00482953f $X=4.61 $Y=0.925
+ $X2=0 $Y2=0
cc_333 N_A_452_419#_c_443_n N_A_778_47#_c_659_n 0.0579205f $X=4.775 $Y=1.39
+ $X2=0 $Y2=0
cc_334 N_A_452_419#_c_444_n N_A_778_47#_c_659_n 0.00428512f $X=4.775 $Y=1.39
+ $X2=0 $Y2=0
cc_335 N_A_452_419#_M1019_g N_A_778_47#_c_667_n 0.0215896f $X=4.735 $Y=2.595
+ $X2=0 $Y2=0
cc_336 N_A_452_419#_c_443_n N_A_778_47#_c_667_n 0.00193953f $X=4.775 $Y=1.39
+ $X2=0 $Y2=0
cc_337 N_A_452_419#_c_440_n N_A_778_47#_c_661_n 0.0150623f $X=4.61 $Y=0.925
+ $X2=0 $Y2=0
cc_338 N_A_452_419#_M1019_g N_VPWR_c_761_n 0.00450239f $X=4.735 $Y=2.595 $X2=0
+ $Y2=0
cc_339 N_A_452_419#_M1019_g N_VPWR_c_764_n 0.00939541f $X=4.735 $Y=2.595 $X2=0
+ $Y2=0
cc_340 N_A_452_419#_M1013_s N_VPWR_c_759_n 0.00310908f $X=2.26 $Y=2.095 $X2=0
+ $Y2=0
cc_341 N_A_452_419#_M1019_g N_VPWR_c_759_n 0.0163871f $X=4.735 $Y=2.595 $X2=0
+ $Y2=0
cc_342 N_A_452_419#_c_438_n N_VGND_c_859_n 0.0207998f $X=2.42 $Y=0.47 $X2=0
+ $Y2=0
cc_343 N_A_452_419#_c_438_n N_VGND_c_860_n 0.0137643f $X=2.42 $Y=0.47 $X2=0
+ $Y2=0
cc_344 N_A_452_419#_c_446_n N_VGND_c_860_n 0.021341f $X=3.71 $Y=0.925 $X2=0
+ $Y2=0
cc_345 N_A_452_419#_c_447_n N_VGND_c_860_n 0.00268757f $X=3.875 $Y=0.765 $X2=0
+ $Y2=0
cc_346 N_A_452_419#_c_442_n N_VGND_c_864_n 0.00154485f $X=3.875 $Y=0.93 $X2=0
+ $Y2=0
cc_347 N_A_452_419#_c_447_n N_VGND_c_864_n 0.00585385f $X=3.875 $Y=0.765 $X2=0
+ $Y2=0
cc_348 N_A_452_419#_M1017_s N_VGND_c_867_n 0.00232985f $X=2.275 $Y=0.235 $X2=0
+ $Y2=0
cc_349 N_A_452_419#_c_438_n N_VGND_c_867_n 0.0131612f $X=2.42 $Y=0.47 $X2=0
+ $Y2=0
cc_350 N_A_452_419#_c_441_n N_VGND_c_867_n 0.00890193f $X=3.87 $Y=0.925 $X2=0
+ $Y2=0
cc_351 N_A_452_419#_c_442_n N_VGND_c_867_n 0.00201388f $X=3.875 $Y=0.93 $X2=0
+ $Y2=0
cc_352 N_A_452_419#_c_447_n N_VGND_c_867_n 0.00648686f $X=3.875 $Y=0.765 $X2=0
+ $Y2=0
cc_353 N_A_928_21#_c_531_n N_A_778_47#_M1022_g 0.00462318f $X=5.18 $Y=0.805
+ $X2=0 $Y2=0
cc_354 N_A_928_21#_c_543_n N_A_778_47#_M1022_g 0.00121823f $X=6.535 $Y=0.47
+ $X2=0 $Y2=0
cc_355 N_A_928_21#_M1016_g N_A_778_47#_M1020_g 0.0177151f $X=5.305 $Y=2.595
+ $X2=0 $Y2=0
cc_356 N_A_928_21#_c_539_n N_A_778_47#_M1020_g 0.00121992f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_357 N_A_928_21#_c_540_n N_A_778_47#_M1020_g 0.0200998f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_358 N_A_928_21#_c_549_n N_A_778_47#_M1020_g 0.023114f $X=6.395 $Y=1.79 $X2=0
+ $Y2=0
cc_359 N_A_928_21#_c_542_n N_A_778_47#_M1020_g 0.00481152f $X=6.48 $Y=1.875
+ $X2=0 $Y2=0
cc_360 N_A_928_21#_c_552_n N_A_778_47#_M1020_g 0.0252795f $X=6.305 $Y=2.24 $X2=0
+ $Y2=0
cc_361 N_A_928_21#_c_553_n N_A_778_47#_M1020_g 0.00677868f $X=6.352 $Y=2.075
+ $X2=0 $Y2=0
cc_362 N_A_928_21#_c_544_n N_A_778_47#_M1020_g 0.00360249f $X=6.8 $Y=1.2 $X2=0
+ $Y2=0
cc_363 N_A_928_21#_c_541_n N_A_778_47#_M1001_g 0.0125202f $X=6.547 $Y=1.035
+ $X2=0 $Y2=0
cc_364 N_A_928_21#_c_543_n N_A_778_47#_M1001_g 0.00948209f $X=6.535 $Y=0.47
+ $X2=0 $Y2=0
cc_365 N_A_928_21#_c_545_n N_A_778_47#_c_656_n 0.00462318f $X=5.427 $Y=1.205
+ $X2=0 $Y2=0
cc_366 N_A_928_21#_c_549_n N_A_778_47#_c_657_n 5.35956e-19 $X=6.395 $Y=1.79
+ $X2=0 $Y2=0
cc_367 N_A_928_21#_c_544_n N_A_778_47#_c_657_n 0.00591381f $X=6.8 $Y=1.2 $X2=0
+ $Y2=0
cc_368 N_A_928_21#_c_530_n N_A_778_47#_c_668_n 0.0169753f $X=4.715 $Y=0.73 $X2=0
+ $Y2=0
cc_369 N_A_928_21#_c_531_n N_A_778_47#_c_668_n 0.00836647f $X=5.18 $Y=0.805
+ $X2=0 $Y2=0
cc_370 N_A_928_21#_M1016_g N_A_778_47#_c_665_n 0.00805041f $X=5.305 $Y=2.595
+ $X2=0 $Y2=0
cc_371 N_A_928_21#_c_530_n N_A_778_47#_c_658_n 0.00442924f $X=4.715 $Y=0.73
+ $X2=0 $Y2=0
cc_372 N_A_928_21#_c_531_n N_A_778_47#_c_658_n 0.00976527f $X=5.18 $Y=0.805
+ $X2=0 $Y2=0
cc_373 N_A_928_21#_M1016_g N_A_778_47#_c_659_n 0.00617324f $X=5.305 $Y=2.595
+ $X2=0 $Y2=0
cc_374 N_A_928_21#_c_539_n N_A_778_47#_c_659_n 0.0334796f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_375 N_A_928_21#_c_540_n N_A_778_47#_c_659_n 0.0162683f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_376 N_A_928_21#_c_550_n N_A_778_47#_c_659_n 0.0123662f $X=5.675 $Y=1.79 $X2=0
+ $Y2=0
cc_377 N_A_928_21#_c_545_n N_A_778_47#_c_659_n 0.00697815f $X=5.427 $Y=1.205
+ $X2=0 $Y2=0
cc_378 N_A_928_21#_c_531_n N_A_778_47#_c_660_n 0.0027586f $X=5.18 $Y=0.805 $X2=0
+ $Y2=0
cc_379 N_A_928_21#_c_539_n N_A_778_47#_c_660_n 0.0200997f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_380 N_A_928_21#_c_540_n N_A_778_47#_c_660_n 0.00513507f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_381 N_A_928_21#_c_545_n N_A_778_47#_c_660_n 0.00836963f $X=5.427 $Y=1.205
+ $X2=0 $Y2=0
cc_382 N_A_928_21#_M1016_g N_A_778_47#_c_667_n 0.00349872f $X=5.305 $Y=2.595
+ $X2=0 $Y2=0
cc_383 N_A_928_21#_c_531_n N_A_778_47#_c_661_n 0.00362689f $X=5.18 $Y=0.805
+ $X2=0 $Y2=0
cc_384 N_A_928_21#_c_545_n N_A_778_47#_c_661_n 0.00308318f $X=5.427 $Y=1.205
+ $X2=0 $Y2=0
cc_385 N_A_928_21#_c_534_n N_A_778_47#_c_662_n 4.38387e-19 $X=6.965 $Y=1.11
+ $X2=0 $Y2=0
cc_386 N_A_928_21#_c_539_n N_A_778_47#_c_662_n 0.0199127f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_387 N_A_928_21#_c_540_n N_A_778_47#_c_662_n 0.00120219f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_388 N_A_928_21#_c_549_n N_A_778_47#_c_662_n 0.0241241f $X=6.395 $Y=1.79 $X2=0
+ $Y2=0
cc_389 N_A_928_21#_c_541_n N_A_778_47#_c_662_n 0.0142152f $X=6.547 $Y=1.035
+ $X2=0 $Y2=0
cc_390 N_A_928_21#_c_542_n N_A_778_47#_c_662_n 0.0389719f $X=6.48 $Y=1.875 $X2=0
+ $Y2=0
cc_391 N_A_928_21#_c_545_n N_A_778_47#_c_662_n 6.66499e-19 $X=5.427 $Y=1.205
+ $X2=0 $Y2=0
cc_392 N_A_928_21#_c_534_n N_A_778_47#_c_663_n 0.00591381f $X=6.965 $Y=1.11
+ $X2=0 $Y2=0
cc_393 N_A_928_21#_c_539_n N_A_778_47#_c_663_n 0.00111281f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_394 N_A_928_21#_c_540_n N_A_778_47#_c_663_n 0.020087f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_395 N_A_928_21#_c_541_n N_A_778_47#_c_663_n 3.64472e-19 $X=6.547 $Y=1.035
+ $X2=0 $Y2=0
cc_396 N_A_928_21#_c_542_n N_A_778_47#_c_663_n 0.00419843f $X=6.48 $Y=1.875
+ $X2=0 $Y2=0
cc_397 N_A_928_21#_M1016_g N_VPWR_c_761_n 0.0258135f $X=5.305 $Y=2.595 $X2=0
+ $Y2=0
cc_398 N_A_928_21#_c_540_n N_VPWR_c_761_n 0.00188061f $X=5.51 $Y=1.37 $X2=0
+ $Y2=0
cc_399 N_A_928_21#_c_549_n N_VPWR_c_761_n 0.00478574f $X=6.395 $Y=1.79 $X2=0
+ $Y2=0
cc_400 N_A_928_21#_c_550_n N_VPWR_c_761_n 0.0207009f $X=5.675 $Y=1.79 $X2=0
+ $Y2=0
cc_401 N_A_928_21#_c_552_n N_VPWR_c_761_n 0.0405136f $X=6.305 $Y=2.24 $X2=0
+ $Y2=0
cc_402 N_A_928_21#_c_533_n N_VPWR_c_762_n 0.00214633f $X=7.235 $Y=1.11 $X2=0
+ $Y2=0
cc_403 N_A_928_21#_M1007_g N_VPWR_c_762_n 0.0278632f $X=7.36 $Y=2.405 $X2=0
+ $Y2=0
cc_404 N_A_928_21#_c_542_n N_VPWR_c_762_n 0.00289924f $X=6.48 $Y=1.875 $X2=0
+ $Y2=0
cc_405 N_A_928_21#_c_553_n N_VPWR_c_762_n 0.0583964f $X=6.352 $Y=2.075 $X2=0
+ $Y2=0
cc_406 N_A_928_21#_c_544_n N_VPWR_c_762_n 2.64278e-19 $X=6.8 $Y=1.2 $X2=0 $Y2=0
cc_407 N_A_928_21#_M1016_g N_VPWR_c_764_n 0.00895812f $X=5.305 $Y=2.595 $X2=0
+ $Y2=0
cc_408 N_A_928_21#_c_552_n N_VPWR_c_765_n 0.0261633f $X=6.305 $Y=2.24 $X2=0
+ $Y2=0
cc_409 N_A_928_21#_M1007_g N_VPWR_c_766_n 0.00781729f $X=7.36 $Y=2.405 $X2=0
+ $Y2=0
cc_410 N_A_928_21#_M1020_d N_VPWR_c_759_n 0.0023218f $X=6.165 $Y=2.095 $X2=0
+ $Y2=0
cc_411 N_A_928_21#_M1016_g N_VPWR_c_759_n 0.014976f $X=5.305 $Y=2.595 $X2=0
+ $Y2=0
cc_412 N_A_928_21#_M1007_g N_VPWR_c_759_n 0.00796052f $X=7.36 $Y=2.405 $X2=0
+ $Y2=0
cc_413 N_A_928_21#_c_552_n N_VPWR_c_759_n 0.0161839f $X=6.305 $Y=2.24 $X2=0
+ $Y2=0
cc_414 N_A_928_21#_M1006_g Q 0.0060281f $X=7.31 $Y=0.625 $X2=0 $Y2=0
cc_415 N_A_928_21#_M1007_g Q 0.0544493f $X=7.36 $Y=2.405 $X2=0 $Y2=0
cc_416 N_A_928_21#_M1008_g Q 0.0100885f $X=7.67 $Y=0.625 $X2=0 $Y2=0
cc_417 N_A_928_21#_c_538_n Q 0.0181573f $X=7.67 $Y=1.11 $X2=0 $Y2=0
cc_418 N_A_928_21#_c_542_n Q 0.0229454f $X=6.48 $Y=1.875 $X2=0 $Y2=0
cc_419 N_A_928_21#_c_544_n Q 4.7897e-19 $X=6.8 $Y=1.2 $X2=0 $Y2=0
cc_420 N_A_928_21#_M1006_g N_Q_c_839_n 0.00225544f $X=7.31 $Y=0.625 $X2=0 $Y2=0
cc_421 N_A_928_21#_M1008_g N_Q_c_839_n 0.00903368f $X=7.67 $Y=0.625 $X2=0 $Y2=0
cc_422 N_A_928_21#_c_530_n N_VGND_c_861_n 0.00397845f $X=4.715 $Y=0.73 $X2=0
+ $Y2=0
cc_423 N_A_928_21#_c_543_n N_VGND_c_861_n 0.011309f $X=6.535 $Y=0.47 $X2=0 $Y2=0
cc_424 N_A_928_21#_c_533_n N_VGND_c_862_n 0.012228f $X=7.235 $Y=1.11 $X2=0 $Y2=0
cc_425 N_A_928_21#_c_534_n N_VGND_c_862_n 2.64278e-19 $X=6.965 $Y=1.11 $X2=0
+ $Y2=0
cc_426 N_A_928_21#_M1006_g N_VGND_c_862_n 0.0124337f $X=7.31 $Y=0.625 $X2=0
+ $Y2=0
cc_427 N_A_928_21#_M1008_g N_VGND_c_862_n 0.00101745f $X=7.67 $Y=0.625 $X2=0
+ $Y2=0
cc_428 N_A_928_21#_c_542_n N_VGND_c_862_n 0.00289924f $X=6.48 $Y=1.875 $X2=0
+ $Y2=0
cc_429 N_A_928_21#_c_543_n N_VGND_c_862_n 0.0396717f $X=6.535 $Y=0.47 $X2=0
+ $Y2=0
cc_430 N_A_928_21#_c_530_n N_VGND_c_864_n 0.00366111f $X=4.715 $Y=0.73 $X2=0
+ $Y2=0
cc_431 N_A_928_21#_c_531_n N_VGND_c_864_n 0.00267712f $X=5.18 $Y=0.805 $X2=0
+ $Y2=0
cc_432 N_A_928_21#_c_543_n N_VGND_c_865_n 0.0197343f $X=6.535 $Y=0.47 $X2=0
+ $Y2=0
cc_433 N_A_928_21#_M1006_g N_VGND_c_866_n 0.00452954f $X=7.31 $Y=0.625 $X2=0
+ $Y2=0
cc_434 N_A_928_21#_M1008_g N_VGND_c_866_n 0.00396337f $X=7.67 $Y=0.625 $X2=0
+ $Y2=0
cc_435 N_A_928_21#_M1001_d N_VGND_c_867_n 0.00232985f $X=6.395 $Y=0.235 $X2=0
+ $Y2=0
cc_436 N_A_928_21#_c_530_n N_VGND_c_867_n 0.00675335f $X=4.715 $Y=0.73 $X2=0
+ $Y2=0
cc_437 N_A_928_21#_c_531_n N_VGND_c_867_n 0.00275062f $X=5.18 $Y=0.805 $X2=0
+ $Y2=0
cc_438 N_A_928_21#_M1006_g N_VGND_c_867_n 0.0044646f $X=7.31 $Y=0.625 $X2=0
+ $Y2=0
cc_439 N_A_928_21#_M1008_g N_VGND_c_867_n 0.005315f $X=7.67 $Y=0.625 $X2=0 $Y2=0
cc_440 N_A_928_21#_c_543_n N_VGND_c_867_n 0.0125687f $X=6.535 $Y=0.47 $X2=0
+ $Y2=0
cc_441 N_A_778_47#_M1020_g N_VPWR_c_761_n 0.0144784f $X=6.04 $Y=2.595 $X2=0
+ $Y2=0
cc_442 N_A_778_47#_c_665_n N_VPWR_c_761_n 0.0129587f $X=5.06 $Y=2.16 $X2=0 $Y2=0
cc_443 N_A_778_47#_c_667_n N_VPWR_c_764_n 0.0178162f $X=4.47 $Y=2.24 $X2=0 $Y2=0
cc_444 N_A_778_47#_M1020_g N_VPWR_c_765_n 0.00939541f $X=6.04 $Y=2.595 $X2=0
+ $Y2=0
cc_445 N_A_778_47#_M1015_d N_VPWR_c_759_n 0.0023187f $X=4.32 $Y=2.095 $X2=0
+ $Y2=0
cc_446 N_A_778_47#_M1020_g N_VPWR_c_759_n 0.0180059f $X=6.04 $Y=2.595 $X2=0
+ $Y2=0
cc_447 N_A_778_47#_c_667_n N_VPWR_c_759_n 0.0123708f $X=4.47 $Y=2.24 $X2=0 $Y2=0
cc_448 N_A_778_47#_c_665_n A_972_419# 0.00826005f $X=5.06 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_449 N_A_778_47#_c_668_n N_VGND_M1005_d 0.0131703f $X=5.06 $Y=0.44 $X2=0 $Y2=0
cc_450 N_A_778_47#_c_658_n N_VGND_M1005_d 0.00156129f $X=5.145 $Y=0.855 $X2=0
+ $Y2=0
cc_451 N_A_778_47#_M1022_g N_VGND_c_861_n 0.0154129f $X=5.96 $Y=0.445 $X2=0
+ $Y2=0
cc_452 N_A_778_47#_c_668_n N_VGND_c_861_n 0.0236638f $X=5.06 $Y=0.44 $X2=0 $Y2=0
cc_453 N_A_778_47#_c_658_n N_VGND_c_861_n 0.00661526f $X=5.145 $Y=0.855 $X2=0
+ $Y2=0
cc_454 N_A_778_47#_c_660_n N_VGND_c_861_n 0.0259511f $X=5.885 $Y=0.94 $X2=0
+ $Y2=0
cc_455 N_A_778_47#_M1001_g N_VGND_c_862_n 0.00336443f $X=6.32 $Y=0.445 $X2=0
+ $Y2=0
cc_456 N_A_778_47#_c_668_n N_VGND_c_864_n 0.0618319f $X=5.06 $Y=0.44 $X2=0 $Y2=0
cc_457 N_A_778_47#_M1022_g N_VGND_c_865_n 0.00585385f $X=5.96 $Y=0.445 $X2=0
+ $Y2=0
cc_458 N_A_778_47#_M1001_g N_VGND_c_865_n 0.00549284f $X=6.32 $Y=0.445 $X2=0
+ $Y2=0
cc_459 N_A_778_47#_M1021_d N_VGND_c_867_n 0.00321357f $X=3.89 $Y=0.235 $X2=0
+ $Y2=0
cc_460 N_A_778_47#_M1022_g N_VGND_c_867_n 0.00775723f $X=5.96 $Y=0.445 $X2=0
+ $Y2=0
cc_461 N_A_778_47#_M1001_g N_VGND_c_867_n 0.0112805f $X=6.32 $Y=0.445 $X2=0
+ $Y2=0
cc_462 N_A_778_47#_c_668_n N_VGND_c_867_n 0.0464445f $X=5.06 $Y=0.44 $X2=0 $Y2=0
cc_463 N_A_778_47#_c_660_n N_VGND_c_867_n 0.0118433f $X=5.885 $Y=0.94 $X2=0
+ $Y2=0
cc_464 N_A_778_47#_c_662_n N_VGND_c_867_n 0.0109709f $X=6.05 $Y=1.02 $X2=0 $Y2=0
cc_465 N_A_778_47#_c_668_n A_880_47# 0.00270787f $X=5.06 $Y=0.44 $X2=-0.19
+ $Y2=-0.245
cc_466 N_VPWR_c_759_n A_766_419# 0.010279f $X=7.92 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_467 N_VPWR_c_759_n A_972_419# 0.0137053f $X=7.92 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_468 N_VPWR_c_762_n Q 0.071709f $X=7.095 $Y=2.05 $X2=0 $Y2=0
cc_469 N_VPWR_c_766_n Q 0.0214072f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_470 N_VPWR_c_759_n Q 0.0209596f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_471 Q N_VGND_c_862_n 0.00860144f $X=7.835 $Y=0.84 $X2=0 $Y2=0
cc_472 N_Q_c_839_n N_VGND_c_862_n 0.0227507f $X=7.755 $Y=0.735 $X2=0 $Y2=0
cc_473 N_Q_c_839_n N_VGND_c_866_n 0.0195834f $X=7.755 $Y=0.735 $X2=0 $Y2=0
cc_474 N_Q_c_839_n N_VGND_c_867_n 0.0207724f $X=7.755 $Y=0.735 $X2=0 $Y2=0
cc_475 Q A_1477_83# 8.93626e-19 $X=7.835 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_476 N_Q_c_839_n A_1477_83# 0.00374071f $X=7.755 $Y=0.735 $X2=-0.19 $Y2=-0.245
cc_477 N_VGND_c_867_n A_542_47# 0.00899413f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
cc_478 N_VGND_c_867_n A_700_47# 0.00940065f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
cc_479 N_VGND_c_867_n A_880_47# 0.00194865f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
cc_480 N_VGND_c_867_n A_1207_47# 0.00396395f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
