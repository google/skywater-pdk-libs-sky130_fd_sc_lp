* File: sky130_fd_sc_lp__a21boi_0.pxi.spice
* Created: Fri Aug 28 09:49:45 2020
* 
x_PM_SKY130_FD_SC_LP__A21BOI_0%B1_N N_B1_N_M1002_g N_B1_N_c_62_n N_B1_N_M1004_g
+ N_B1_N_c_64_n B1_N B1_N B1_N N_B1_N_c_66_n PM_SKY130_FD_SC_LP__A21BOI_0%B1_N
x_PM_SKY130_FD_SC_LP__A21BOI_0%A_27_47# N_A_27_47#_M1002_s N_A_27_47#_M1004_s
+ N_A_27_47#_c_96_n N_A_27_47#_c_97_n N_A_27_47#_c_98_n N_A_27_47#_M1006_g
+ N_A_27_47#_c_104_n N_A_27_47#_c_105_n N_A_27_47#_M1001_g N_A_27_47#_c_99_n
+ N_A_27_47#_c_100_n N_A_27_47#_c_101_n N_A_27_47#_c_102_n
+ PM_SKY130_FD_SC_LP__A21BOI_0%A_27_47#
x_PM_SKY130_FD_SC_LP__A21BOI_0%A1 N_A1_M1000_g N_A1_c_162_n N_A1_M1005_g A1 A1
+ A1 PM_SKY130_FD_SC_LP__A21BOI_0%A1
x_PM_SKY130_FD_SC_LP__A21BOI_0%A2 N_A2_M1007_g N_A2_c_205_n N_A2_c_206_n
+ N_A2_M1003_g N_A2_c_208_n A2 A2 A2 N_A2_c_210_n
+ PM_SKY130_FD_SC_LP__A21BOI_0%A2
x_PM_SKY130_FD_SC_LP__A21BOI_0%VPWR N_VPWR_M1004_d N_VPWR_M1005_d N_VPWR_c_239_n
+ N_VPWR_c_240_n VPWR N_VPWR_c_241_n N_VPWR_c_242_n N_VPWR_c_243_n
+ N_VPWR_c_238_n N_VPWR_c_245_n N_VPWR_c_246_n PM_SKY130_FD_SC_LP__A21BOI_0%VPWR
x_PM_SKY130_FD_SC_LP__A21BOI_0%Y N_Y_M1006_d N_Y_M1001_s N_Y_c_284_n Y Y Y Y
+ N_Y_c_276_n PM_SKY130_FD_SC_LP__A21BOI_0%Y
x_PM_SKY130_FD_SC_LP__A21BOI_0%A_324_483# N_A_324_483#_M1001_d
+ N_A_324_483#_M1003_d N_A_324_483#_c_311_n N_A_324_483#_c_312_n
+ N_A_324_483#_c_313_n N_A_324_483#_c_314_n
+ PM_SKY130_FD_SC_LP__A21BOI_0%A_324_483#
x_PM_SKY130_FD_SC_LP__A21BOI_0%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_c_335_n
+ VGND N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n N_VGND_c_339_n
+ N_VGND_c_340_n PM_SKY130_FD_SC_LP__A21BOI_0%VGND
cc_1 VNB N_B1_N_M1002_g 0.0721776f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_2 VNB B1_N 0.00336351f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_A_27_47#_c_96_n 0.0819332f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.345
cc_4 VNB N_A_27_47#_c_97_n 0.0125511f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_5 VNB N_A_27_47#_c_98_n 0.0184689f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_6 VNB N_A_27_47#_c_99_n 0.0208551f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.84
cc_7 VNB N_A_27_47#_c_100_n 0.0130772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_101_n 0.00432805f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=2.405
cc_9 VNB N_A_27_47#_c_102_n 0.0289089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_M1000_g 0.0389487f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_11 VNB N_A1_c_162_n 0.0506582f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.872
cc_12 VNB A1 0.0100447f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_13 VNB N_A2_M1007_g 0.0238873f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_14 VNB N_A2_c_205_n 0.0365301f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.872
cc_15 VNB N_A2_c_206_n 0.00666448f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=2.148
cc_16 VNB N_A2_M1003_g 0.00912821f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_17 VNB N_A2_c_208_n 0.0200975f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_18 VNB A2 0.0404124f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_19 VNB N_A2_c_210_n 0.0334055f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.675
cc_20 VNB N_VPWR_c_238_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB Y 0.00285875f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_22 VNB N_Y_c_276_n 0.0121362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_335_n 0.0175746f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_24 VNB N_VGND_c_336_n 0.0356726f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_25 VNB N_VGND_c_337_n 0.0260593f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.84
cc_26 VNB N_VGND_c_338_n 0.0169405f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=1.84
cc_27 VNB N_VGND_c_339_n 0.172691f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=2.035
cc_28 VNB N_VGND_c_340_n 0.00510915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_B1_N_M1002_g 0.00110475f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_30 VPB N_B1_N_c_62_n 0.0216433f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=2.148
cc_31 VPB N_B1_N_M1004_g 0.0300489f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_32 VPB N_B1_N_c_64_n 0.0233482f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=2.345
cc_33 VPB B1_N 0.00911832f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_34 VPB N_B1_N_c_66_n 0.0219801f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.84
cc_35 VPB N_A_27_47#_c_97_n 0.022251f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_36 VPB N_A_27_47#_c_104_n 0.0264151f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_37 VPB N_A_27_47#_c_105_n 0.00872638f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_38 VPB N_A_27_47#_M1001_g 0.022372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_100_n 0.0655735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A1_c_162_n 0.0304223f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.872
cc_41 VPB N_A1_M1005_g 0.0407902f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.345
cc_42 VPB A1 0.00519045f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_43 VPB N_A2_M1003_g 0.0632568f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_44 VPB A2 0.0117702f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_45 VPB N_VPWR_c_239_n 0.00935902f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_46 VPB N_VPWR_c_240_n 0.00912313f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_47 VPB N_VPWR_c_241_n 0.0164641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_242_n 0.0321579f $X=-0.19 $Y=1.655 $X2=0.712 $Y2=1.665
cc_49 VPB N_VPWR_c_243_n 0.0172605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_238_n 0.0654286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_245_n 0.00598038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_246_n 0.00507132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB Y 0.00183012f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_54 VPB Y 0.0203612f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_55 VPB N_A_324_483#_c_311_n 0.00492707f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_56 VPB N_A_324_483#_c_312_n 0.0187627f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=2.345
cc_57 VPB N_A_324_483#_c_313_n 0.00320584f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_58 VPB N_A_324_483#_c_314_n 0.0365357f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 N_B1_N_M1002_g N_A_27_47#_c_96_n 0.0435681f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_60 B1_N N_A_27_47#_c_96_n 0.00319916f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_61 N_B1_N_c_66_n N_A_27_47#_c_96_n 0.00193775f $X=0.63 $Y=1.84 $X2=0 $Y2=0
cc_62 N_B1_N_M1002_g N_A_27_47#_c_97_n 0.00550057f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_63 B1_N N_A_27_47#_c_97_n 0.00252242f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_64 N_B1_N_c_66_n N_A_27_47#_c_97_n 0.0127506f $X=0.63 $Y=1.84 $X2=0 $Y2=0
cc_65 N_B1_N_M1002_g N_A_27_47#_c_98_n 0.0056502f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_66 N_B1_N_c_62_n N_A_27_47#_c_105_n 0.0127506f $X=0.597 $Y=2.148 $X2=0 $Y2=0
cc_67 N_B1_N_c_64_n N_A_27_47#_M1001_g 8.37917e-19 $X=0.597 $Y=2.345 $X2=0 $Y2=0
cc_68 B1_N N_A_27_47#_M1001_g 4.94949e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_69 N_B1_N_M1002_g N_A_27_47#_c_99_n 0.00561773f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_70 N_B1_N_M1002_g N_A_27_47#_c_100_n 0.0348284f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_71 B1_N N_A_27_47#_c_100_n 0.0731454f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_72 N_B1_N_M1002_g N_A_27_47#_c_101_n 0.037174f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_73 B1_N N_A_27_47#_c_101_n 0.0336917f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_74 N_B1_N_c_66_n N_A_27_47#_c_101_n 0.00126457f $X=0.63 $Y=1.84 $X2=0 $Y2=0
cc_75 N_B1_N_M1004_g N_VPWR_c_239_n 0.0111694f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_76 N_B1_N_c_64_n N_VPWR_c_239_n 0.00119629f $X=0.597 $Y=2.345 $X2=0 $Y2=0
cc_77 B1_N N_VPWR_c_239_n 0.0266711f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_78 N_B1_N_M1004_g N_VPWR_c_241_n 0.00396895f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_79 N_B1_N_M1004_g N_VPWR_c_238_n 0.00789173f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_80 B1_N N_VPWR_c_238_n 0.00299306f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_81 N_B1_N_M1002_g Y 2.21541e-19 $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_82 B1_N Y 0.0799292f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_83 N_B1_N_c_66_n Y 9.8656e-19 $X=0.63 $Y=1.84 $X2=0 $Y2=0
cc_84 N_B1_N_c_62_n Y 9.8656e-19 $X=0.597 $Y=2.148 $X2=0 $Y2=0
cc_85 N_B1_N_M1004_g Y 0.00513287f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_86 N_B1_N_M1002_g N_VGND_c_336_n 0.00991559f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_87 N_B1_N_M1002_g N_VGND_c_339_n 0.00780787f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_96_n N_A1_M1000_g 0.00547701f $X=1.16 $Y=1.435 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_98_n N_A1_M1000_g 0.0214029f $X=1.245 $Y=0.765 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_96_n N_A1_c_162_n 0.0283947f $X=1.16 $Y=1.435 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_104_n N_A1_c_162_n 0.00774427f $X=1.47 $Y=2.19 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_97_n N_A1_M1005_g 0.00262645f $X=1.16 $Y=2.115 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_104_n N_A1_M1005_g 0.0178451f $X=1.47 $Y=2.19 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_97_n A1 2.1137e-19 $X=1.16 $Y=2.115 $X2=0 $Y2=0
cc_95 N_A_27_47#_M1001_g N_VPWR_c_239_n 0.00234177f $X=1.545 $Y=2.735 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_c_100_n N_VPWR_c_239_n 0.0131449f $X=0.26 $Y=2.795 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_100_n N_VPWR_c_241_n 0.0125145f $X=0.26 $Y=2.795 $X2=0 $Y2=0
cc_98 N_A_27_47#_M1001_g N_VPWR_c_242_n 0.00525778f $X=1.545 $Y=2.735 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_M1001_g N_VPWR_c_238_n 0.0110397f $X=1.545 $Y=2.735 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_100_n N_VPWR_c_238_n 0.00964185f $X=0.26 $Y=2.795 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_98_n N_Y_c_284_n 0.00305845f $X=1.245 $Y=0.765 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_96_n Y 0.00293354f $X=1.16 $Y=1.435 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_97_n Y 0.0137245f $X=1.16 $Y=2.115 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_101_n Y 0.00165124f $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_97_n Y 0.0107549f $X=1.16 $Y=2.115 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_104_n Y 0.016193f $X=1.47 $Y=2.19 $X2=0 $Y2=0
cc_107 N_A_27_47#_c_105_n Y 0.00642263f $X=1.235 $Y=2.19 $X2=0 $Y2=0
cc_108 N_A_27_47#_M1001_g Y 0.0107494f $X=1.545 $Y=2.735 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_96_n N_Y_c_276_n 0.0135461f $X=1.16 $Y=1.435 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_98_n N_Y_c_276_n 0.00688411f $X=1.245 $Y=0.765 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_101_n N_Y_c_276_n 0.0388231f $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_104_n N_A_324_483#_c_311_n 0.00154463f $X=1.47 $Y=2.19 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_104_n N_A_324_483#_c_313_n 0.00108951f $X=1.47 $Y=2.19 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_96_n N_VGND_c_336_n 0.0109008f $X=1.16 $Y=1.435 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_98_n N_VGND_c_336_n 0.00386375f $X=1.245 $Y=0.765 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_99_n N_VGND_c_336_n 0.0161226f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_101_n N_VGND_c_336_n 0.0436037f $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_96_n N_VGND_c_337_n 4.96289e-19 $X=1.16 $Y=1.435 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_98_n N_VGND_c_337_n 0.0057945f $X=1.245 $Y=0.765 $X2=0 $Y2=0
cc_120 N_A_27_47#_M1002_s N_VGND_c_339_n 0.00227481f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_c_96_n N_VGND_c_339_n 6.69668e-19 $X=1.16 $Y=1.435 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_98_n N_VGND_c_339_n 0.0113118f $X=1.245 $Y=0.765 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_99_n N_VGND_c_339_n 0.0108688f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_101_n N_VGND_c_339_n 0.00783385f $X=0.925 $Y=0.93 $X2=0
+ $Y2=0
cc_125 N_A1_M1000_g N_A2_M1007_g 0.0531201f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_126 A1 N_A2_M1007_g 0.00496689f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_127 A1 N_A2_c_205_n 0.00971705f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_128 N_A1_c_162_n N_A2_c_206_n 0.00499022f $X=1.975 $Y=1.875 $X2=0 $Y2=0
cc_129 A1 N_A2_c_206_n 0.00594249f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_130 N_A1_M1005_g N_A2_c_208_n 0.0291624f $X=1.975 $Y=2.735 $X2=0 $Y2=0
cc_131 N_A1_c_162_n A2 5.08847e-19 $X=1.975 $Y=1.875 $X2=0 $Y2=0
cc_132 A1 A2 0.0885427f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_133 N_A1_M1000_g N_A2_c_210_n 0.00326168f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A1_c_162_n N_A2_c_210_n 0.0291624f $X=1.975 $Y=1.875 $X2=0 $Y2=0
cc_135 A1 N_A2_c_210_n 0.00868077f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_136 N_A1_M1005_g N_VPWR_c_240_n 0.00305256f $X=1.975 $Y=2.735 $X2=0 $Y2=0
cc_137 N_A1_M1005_g N_VPWR_c_242_n 0.00545548f $X=1.975 $Y=2.735 $X2=0 $Y2=0
cc_138 N_A1_M1005_g N_VPWR_c_238_n 0.0103212f $X=1.975 $Y=2.735 $X2=0 $Y2=0
cc_139 N_A1_M1000_g N_Y_c_284_n 0.00657543f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A1_c_162_n N_Y_c_284_n 0.00167601f $X=1.975 $Y=1.875 $X2=0 $Y2=0
cc_141 N_A1_M1005_g Y 0.00423225f $X=1.975 $Y=2.735 $X2=0 $Y2=0
cc_142 N_A1_M1000_g N_Y_c_276_n 0.00677724f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A1_c_162_n N_Y_c_276_n 0.00691217f $X=1.975 $Y=1.875 $X2=0 $Y2=0
cc_144 A1 N_Y_c_276_n 0.0682438f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_145 N_A1_M1005_g N_A_324_483#_c_311_n 0.00267012f $X=1.975 $Y=2.735 $X2=0
+ $Y2=0
cc_146 N_A1_M1005_g N_A_324_483#_c_312_n 0.0150291f $X=1.975 $Y=2.735 $X2=0
+ $Y2=0
cc_147 A1 N_A_324_483#_c_312_n 0.0285683f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_148 N_A1_c_162_n N_A_324_483#_c_313_n 0.00443365f $X=1.975 $Y=1.875 $X2=0
+ $Y2=0
cc_149 A1 N_A_324_483#_c_313_n 0.0139995f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_150 N_A1_M1000_g N_VGND_c_335_n 0.00225543f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_151 A1 N_VGND_c_335_n 0.0122038f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_152 N_A1_M1000_g N_VGND_c_337_n 0.0054978f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_153 N_A1_M1000_g N_VGND_c_339_n 0.00906239f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_154 A1 N_VGND_c_339_n 0.0146292f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_155 N_A2_M1003_g N_VPWR_c_240_n 0.00302473f $X=2.405 $Y=2.735 $X2=0 $Y2=0
cc_156 N_A2_M1003_g N_VPWR_c_243_n 0.00545548f $X=2.405 $Y=2.735 $X2=0 $Y2=0
cc_157 N_A2_M1003_g N_VPWR_c_238_n 0.0110328f $X=2.405 $Y=2.735 $X2=0 $Y2=0
cc_158 N_A2_M1007_g N_Y_c_284_n 8.98642e-19 $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A2_M1003_g N_A_324_483#_c_312_n 0.01941f $X=2.405 $Y=2.735 $X2=0 $Y2=0
cc_160 N_A2_c_208_n N_A_324_483#_c_312_n 7.45206e-19 $X=2.502 $Y=1.51 $X2=0
+ $Y2=0
cc_161 A2 N_A_324_483#_c_312_n 0.0289557f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_162 N_A2_M1003_g N_A_324_483#_c_314_n 0.00590286f $X=2.405 $Y=2.735 $X2=0
+ $Y2=0
cc_163 N_A2_M1007_g N_VGND_c_335_n 0.0125719f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A2_c_205_n N_VGND_c_335_n 0.007757f $X=2.33 $Y=0.89 $X2=0 $Y2=0
cc_165 N_A2_M1007_g N_VGND_c_337_n 0.00486043f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A2_M1007_g N_VGND_c_339_n 0.00432334f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A2_c_205_n N_VGND_c_339_n 3.11509e-19 $X=2.33 $Y=0.89 $X2=0 $Y2=0
cc_168 A2 N_VGND_c_339_n 0.0153012f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_169 N_VPWR_c_239_n Y 0.0283963f $X=0.69 $Y=2.795 $X2=0 $Y2=0
cc_170 N_VPWR_c_242_n Y 0.0277978f $X=2.055 $Y=3.33 $X2=0 $Y2=0
cc_171 N_VPWR_c_238_n Y 0.0159158f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_240_n N_A_324_483#_c_311_n 0.00143344f $X=2.19 $Y=2.57 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_242_n N_A_324_483#_c_311_n 0.0153728f $X=2.055 $Y=3.33 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_238_n N_A_324_483#_c_311_n 0.00882204f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_240_n N_A_324_483#_c_312_n 0.0213307f $X=2.19 $Y=2.57 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_240_n N_A_324_483#_c_314_n 0.00146069f $X=2.19 $Y=2.57 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_243_n N_A_324_483#_c_314_n 0.0197554f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_238_n N_A_324_483#_c_314_n 0.0113371f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_179 Y N_A_324_483#_c_311_n 0.0403648f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_180 Y N_A_324_483#_c_313_n 0.0148191f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_181 N_Y_c_284_n N_VGND_c_335_n 0.0109883f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_182 N_Y_c_284_n N_VGND_c_337_n 0.0149222f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_183 N_Y_M1006_d N_VGND_c_339_n 0.00226149f $X=1.32 $Y=0.235 $X2=0 $Y2=0
cc_184 N_Y_c_284_n N_VGND_c_339_n 0.0115755f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_185 N_VGND_c_339_n A_350_47# 0.00288969f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
