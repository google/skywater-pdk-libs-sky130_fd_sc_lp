* File: sky130_fd_sc_lp__srdlxtp_1.pxi.spice
* Created: Fri Aug 28 11:33:22 2020
* 
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%A_84_153# N_A_84_153#_M1023_s
+ N_A_84_153#_M1026_d N_A_84_153#_M1013_g N_A_84_153#_M1004_g
+ N_A_84_153#_c_185_n N_A_84_153#_M1015_g N_A_84_153#_M1024_g
+ N_A_84_153#_c_186_n N_A_84_153#_M1006_g N_A_84_153#_c_188_n
+ N_A_84_153#_c_189_n N_A_84_153#_c_205_n N_A_84_153#_c_190_n
+ N_A_84_153#_c_207_n N_A_84_153#_c_225_p N_A_84_153#_c_345_p
+ N_A_84_153#_c_208_n N_A_84_153#_c_255_p N_A_84_153#_c_191_n
+ N_A_84_153#_c_257_p N_A_84_153#_c_210_n N_A_84_153#_c_192_n
+ N_A_84_153#_c_211_n N_A_84_153#_c_193_n N_A_84_153#_c_194_n
+ N_A_84_153#_c_195_n N_A_84_153#_c_355_p N_A_84_153#_c_196_n
+ N_A_84_153#_c_258_p N_A_84_153#_c_197_n N_A_84_153#_c_198_n
+ PM_SKY130_FD_SC_LP__SRDLXTP_1%A_84_153#
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%D N_D_M1022_g N_D_M1014_g N_D_c_420_n
+ N_D_c_421_n D PM_SKY130_FD_SC_LP__SRDLXTP_1%D
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%A_226_491# N_A_226_491#_M1014_s
+ N_A_226_491#_M1022_s N_A_226_491#_c_471_n N_A_226_491#_c_465_n
+ N_A_226_491#_M1025_g N_A_226_491#_c_472_n N_A_226_491#_M1012_g
+ N_A_226_491#_c_473_n N_A_226_491#_c_474_n N_A_226_491#_c_475_n
+ N_A_226_491#_c_466_n N_A_226_491#_c_476_n N_A_226_491#_c_477_n
+ N_A_226_491#_c_467_n N_A_226_491#_c_468_n N_A_226_491#_c_469_n
+ N_A_226_491#_c_470_n PM_SKY130_FD_SC_LP__SRDLXTP_1%A_226_491#
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%A_114_179# N_A_114_179#_M1013_d
+ N_A_114_179#_M1004_d N_A_114_179#_M1002_g N_A_114_179#_c_570_n
+ N_A_114_179#_M1003_g N_A_114_179#_c_572_n N_A_114_179#_c_573_n
+ N_A_114_179#_c_574_n N_A_114_179#_c_585_n N_A_114_179#_M1020_g
+ N_A_114_179#_c_575_n N_A_114_179#_c_576_n N_A_114_179#_c_577_n
+ N_A_114_179#_c_578_n N_A_114_179#_c_579_n N_A_114_179#_c_588_n
+ N_A_114_179#_c_580_n N_A_114_179#_c_581_n N_A_114_179#_c_582_n
+ PM_SKY130_FD_SC_LP__SRDLXTP_1%A_114_179#
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%A_831_21# N_A_831_21#_M1005_d
+ N_A_831_21#_M1021_s N_A_831_21#_M1007_g N_A_831_21#_c_701_n
+ N_A_831_21#_c_702_n N_A_831_21#_M1001_g N_A_831_21#_M1009_g
+ N_A_831_21#_c_704_n N_A_831_21#_c_705_n N_A_831_21#_c_706_n
+ N_A_831_21#_c_707_n N_A_831_21#_c_708_n N_A_831_21#_c_709_n
+ PM_SKY130_FD_SC_LP__SRDLXTP_1%A_831_21#
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%GATE N_GATE_c_777_n N_GATE_M1026_g
+ N_GATE_M1023_g N_GATE_c_779_n GATE GATE N_GATE_c_780_n N_GATE_c_781_n
+ PM_SKY130_FD_SC_LP__SRDLXTP_1%GATE
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%SLEEP_B N_SLEEP_B_M1017_g N_SLEEP_B_M1018_g
+ N_SLEEP_B_c_821_n N_SLEEP_B_M1019_g SLEEP_B SLEEP_B N_SLEEP_B_c_823_n
+ PM_SKY130_FD_SC_LP__SRDLXTP_1%SLEEP_B
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%A_662_47# N_A_662_47#_M1003_d
+ N_A_662_47#_M1024_d N_A_662_47#_M1016_g N_A_662_47#_M1005_g
+ N_A_662_47#_M1021_g N_A_662_47#_c_881_n N_A_662_47#_c_882_n
+ N_A_662_47#_c_868_n N_A_662_47#_c_884_n N_A_662_47#_c_869_n
+ N_A_662_47#_c_870_n N_A_662_47#_c_871_n N_A_662_47#_M1000_g
+ N_A_662_47#_M1011_g N_A_662_47#_c_873_n N_A_662_47#_c_886_n
+ N_A_662_47#_c_874_n N_A_662_47#_c_887_n N_A_662_47#_c_888_n
+ N_A_662_47#_c_875_n N_A_662_47#_c_876_n N_A_662_47#_c_877_n
+ N_A_662_47#_c_878_n N_A_662_47#_c_879_n
+ PM_SKY130_FD_SC_LP__SRDLXTP_1%A_662_47#
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%A_1530_367# N_A_1530_367#_M1011_s
+ N_A_1530_367#_M1000_s N_A_1530_367#_M1010_g N_A_1530_367#_M1008_g
+ N_A_1530_367#_c_1033_n N_A_1530_367#_c_1026_n N_A_1530_367#_c_1027_n
+ N_A_1530_367#_c_1028_n N_A_1530_367#_c_1029_n N_A_1530_367#_c_1030_n
+ N_A_1530_367#_c_1031_n PM_SKY130_FD_SC_LP__SRDLXTP_1%A_1530_367#
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%VPWR N_VPWR_M1004_s N_VPWR_M1022_d
+ N_VPWR_M1000_d N_VPWR_c_1084_n N_VPWR_c_1085_n N_VPWR_c_1086_n N_VPWR_c_1087_n
+ VPWR N_VPWR_c_1088_n N_VPWR_c_1089_n N_VPWR_c_1090_n N_VPWR_c_1083_n
+ N_VPWR_c_1092_n N_VPWR_c_1093_n PM_SKY130_FD_SC_LP__SRDLXTP_1%VPWR
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%A_476_47# N_A_476_47#_M1025_d
+ N_A_476_47#_M1012_d N_A_476_47#_c_1172_n N_A_476_47#_c_1173_n
+ N_A_476_47#_c_1174_n N_A_476_47#_c_1176_n N_A_476_47#_c_1177_n
+ N_A_476_47#_c_1175_n PM_SKY130_FD_SC_LP__SRDLXTP_1%A_476_47#
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%KAPWR N_KAPWR_M1001_d N_KAPWR_M1021_d
+ N_KAPWR_M1018_d N_KAPWR_c_1242_n N_KAPWR_c_1243_n N_KAPWR_c_1244_n
+ N_KAPWR_c_1245_n KAPWR N_KAPWR_c_1246_n N_KAPWR_c_1247_n
+ PM_SKY130_FD_SC_LP__SRDLXTP_1%KAPWR
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%Q N_Q_M1010_d N_Q_M1008_d N_Q_c_1339_n
+ N_Q_c_1340_n N_Q_c_1336_n Q Q N_Q_c_1338_n Q PM_SKY130_FD_SC_LP__SRDLXTP_1%Q
x_PM_SKY130_FD_SC_LP__SRDLXTP_1%VGND N_VGND_M1013_s N_VGND_M1014_d
+ N_VGND_M1009_d N_VGND_M1019_d N_VGND_M1011_d N_VGND_c_1356_n N_VGND_c_1357_n
+ N_VGND_c_1358_n N_VGND_c_1359_n N_VGND_c_1360_n N_VGND_c_1361_n
+ N_VGND_c_1362_n N_VGND_c_1363_n N_VGND_c_1364_n N_VGND_c_1365_n
+ N_VGND_c_1366_n N_VGND_c_1367_n VGND N_VGND_c_1368_n N_VGND_c_1369_n
+ N_VGND_c_1370_n N_VGND_c_1371_n PM_SKY130_FD_SC_LP__SRDLXTP_1%VGND
cc_1 VNB N_A_84_153#_M1013_g 0.0415426f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.105
cc_2 VNB N_A_84_153#_c_185_n 0.00854066f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.7
cc_3 VNB N_A_84_153#_c_186_n 0.0486161f $X=-0.19 $Y=-0.245 $X2=3.84 $Y2=1.185
cc_4 VNB N_A_84_153#_M1006_g 0.0411708f $X=-0.19 $Y=-0.245 $X2=3.84 $Y2=0.445
cc_5 VNB N_A_84_153#_c_188_n 0.00213573f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.7
cc_6 VNB N_A_84_153#_c_189_n 0.0202524f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.79
cc_7 VNB N_A_84_153#_c_190_n 0.00661097f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.71
cc_8 VNB N_A_84_153#_c_191_n 0.00251061f $X=-0.19 $Y=-0.245 $X2=4.29 $Y2=2.075
cc_9 VNB N_A_84_153#_c_192_n 0.00480307f $X=-0.19 $Y=-0.245 $X2=6.58 $Y2=0.59
cc_10 VNB N_A_84_153#_c_193_n 0.00794943f $X=-0.19 $Y=-0.245 $X2=6.665 $Y2=1.82
cc_11 VNB N_A_84_153#_c_194_n 0.00260266f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.71
cc_12 VNB N_A_84_153#_c_195_n 0.00302073f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.71
cc_13 VNB N_A_84_153#_c_196_n 0.00410343f $X=-0.19 $Y=-0.245 $X2=4.21 $Y2=1.35
cc_14 VNB N_A_84_153#_c_197_n 0.00601898f $X=-0.19 $Y=-0.245 $X2=6.155 $Y2=0.465
cc_15 VNB N_A_84_153#_c_198_n 0.00893232f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.7
cc_16 VNB N_D_M1022_g 0.036406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_D_M1014_g 0.0254026f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.625
cc_18 VNB N_D_c_420_n 0.0447453f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.105
cc_19 VNB N_D_c_421_n 0.0155921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB D 0.00271789f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.775
cc_21 VNB N_A_226_491#_c_465_n 0.0198916f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.775
cc_22 VNB N_A_226_491#_c_466_n 0.00319274f $X=-0.19 $Y=-0.245 $X2=3.525
+ $Y2=2.775
cc_23 VNB N_A_226_491#_c_467_n 0.0151331f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.79
cc_24 VNB N_A_226_491#_c_468_n 0.00294575f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.13
cc_25 VNB N_A_226_491#_c_469_n 0.0511094f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.71
cc_26 VNB N_A_226_491#_c_470_n 0.0369897f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=2.99
cc_27 VNB N_A_114_179#_M1002_g 0.0330522f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.105
cc_28 VNB N_A_114_179#_c_570_n 0.00827357f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.775
cc_29 VNB N_A_114_179#_M1003_g 0.0402896f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.7
cc_30 VNB N_A_114_179#_c_572_n 0.0117911f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.775
cc_31 VNB N_A_114_179#_c_573_n 0.00712254f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.775
cc_32 VNB N_A_114_179#_c_574_n 0.00299402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_114_179#_c_575_n 0.0217876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_114_179#_c_576_n 0.00664455f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=1.79
cc_35 VNB N_A_114_179#_c_577_n 0.00921217f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.71
cc_36 VNB N_A_114_179#_c_578_n 0.0342506f $X=-0.19 $Y=-0.245 $X2=3.312 $Y2=2.905
cc_37 VNB N_A_114_179#_c_579_n 0.00120897f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.13
cc_38 VNB N_A_114_179#_c_580_n 0.00580575f $X=-0.19 $Y=-0.245 $X2=4.205 $Y2=2.99
cc_39 VNB N_A_114_179#_c_581_n 0.00571351f $X=-0.19 $Y=-0.245 $X2=4.29 $Y2=1.515
cc_40 VNB N_A_114_179#_c_582_n 0.0320113f $X=-0.19 $Y=-0.245 $X2=4.29 $Y2=2.075
cc_41 VNB N_A_831_21#_M1007_g 0.0167461f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.105
cc_42 VNB N_A_831_21#_c_701_n 0.00914164f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.775
cc_43 VNB N_A_831_21#_c_702_n 0.00618076f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.735
cc_44 VNB N_A_831_21#_M1009_g 0.0168164f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.775
cc_45 VNB N_A_831_21#_c_704_n 0.045665f $X=-0.19 $Y=-0.245 $X2=3.525 $Y2=2.775
cc_46 VNB N_A_831_21#_c_705_n 0.00914104f $X=-0.19 $Y=-0.245 $X2=3.525 $Y2=2.775
cc_47 VNB N_A_831_21#_c_706_n 0.0030293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_831_21#_c_707_n 0.0149981f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=1.79
cc_49 VNB N_A_831_21#_c_708_n 0.00571827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_831_21#_c_709_n 0.012649f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=1.955
cc_51 VNB N_GATE_c_777_n 0.0216089f $X=-0.19 $Y=-0.245 $X2=6.385 $Y2=1.675
cc_52 VNB N_GATE_M1023_g 0.0247835f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.105
cc_53 VNB N_GATE_c_779_n 0.011743f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.775
cc_54 VNB N_GATE_c_780_n 0.0202831f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.295
cc_55 VNB N_GATE_c_781_n 0.00990985f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.775
cc_56 VNB N_SLEEP_B_M1017_g 0.0206776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_SLEEP_B_M1018_g 0.0230491f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.625
cc_58 VNB N_SLEEP_B_c_821_n 0.0192814f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.105
cc_59 VNB SLEEP_B 0.0187774f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.735
cc_60 VNB N_SLEEP_B_c_823_n 0.0504894f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.775
cc_61 VNB N_A_662_47#_M1016_g 0.019145f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.105
cc_62 VNB N_A_662_47#_M1005_g 0.0239909f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.735
cc_63 VNB N_A_662_47#_M1021_g 0.0232001f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.775
cc_64 VNB N_A_662_47#_c_868_n 0.00507677f $X=-0.19 $Y=-0.245 $X2=3.525 $Y2=2.775
cc_65 VNB N_A_662_47#_c_869_n 0.0173719f $X=-0.19 $Y=-0.245 $X2=3.84 $Y2=0.445
cc_66 VNB N_A_662_47#_c_870_n 0.0298934f $X=-0.19 $Y=-0.245 $X2=3.84 $Y2=0.445
cc_67 VNB N_A_662_47#_c_871_n 0.0123106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_662_47#_M1011_g 0.0283957f $X=-0.19 $Y=-0.245 $X2=3.45 $Y2=2.13
cc_69 VNB N_A_662_47#_c_873_n 0.0238564f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.905
cc_70 VNB N_A_662_47#_c_874_n 0.00193638f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.13
cc_71 VNB N_A_662_47#_c_875_n 0.0190067f $X=-0.19 $Y=-0.245 $X2=4.29 $Y2=2.905
cc_72 VNB N_A_662_47#_c_876_n 0.00530144f $X=-0.19 $Y=-0.245 $X2=4.375 $Y2=2.16
cc_73 VNB N_A_662_47#_c_877_n 0.00760689f $X=-0.19 $Y=-0.245 $X2=6.58 $Y2=0.59
cc_74 VNB N_A_662_47#_c_878_n 0.00488356f $X=-0.19 $Y=-0.245 $X2=6.32 $Y2=0.59
cc_75 VNB N_A_662_47#_c_879_n 0.0681492f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.79
cc_76 VNB N_A_1530_367#_M1010_g 0.0284723f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.105
cc_77 VNB N_A_1530_367#_M1008_g 6.10221e-19 $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=2.735
cc_78 VNB N_A_1530_367#_c_1026_n 0.00739702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1530_367#_c_1027_n 0.0120223f $X=-0.19 $Y=-0.245 $X2=3.84
+ $Y2=1.185
cc_80 VNB N_A_1530_367#_c_1028_n 0.0420777f $X=-0.19 $Y=-0.245 $X2=3.84
+ $Y2=0.445
cc_81 VNB N_A_1530_367#_c_1029_n 2.14189e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1530_367#_c_1030_n 0.00560529f $X=-0.19 $Y=-0.245 $X2=3.03
+ $Y2=1.79
cc_83 VNB N_A_1530_367#_c_1031_n 0.00591987f $X=-0.19 $Y=-0.245 $X2=3.03
+ $Y2=2.13
cc_84 VNB N_VPWR_c_1083_n 0.382608f $X=-0.19 $Y=-0.245 $X2=3.312 $Y2=2.905
cc_85 VNB N_A_476_47#_c_1172_n 0.00620369f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.625
cc_86 VNB N_A_476_47#_c_1173_n 0.0134178f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.735
cc_87 VNB N_A_476_47#_c_1174_n 0.00461988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_476_47#_c_1175_n 7.291e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_Q_c_1336_n 0.0242086f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.7
cc_90 VNB Q 0.008411f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.295
cc_91 VNB N_Q_c_1338_n 0.0294022f $X=-0.19 $Y=-0.245 $X2=3.525 $Y2=2.775
cc_92 VNB N_VGND_c_1356_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.7
cc_93 VNB N_VGND_c_1357_n 0.0812624f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=2.775
cc_94 VNB N_VGND_c_1358_n 0.00457095f $X=-0.19 $Y=-0.245 $X2=3.525 $Y2=2.775
cc_95 VNB N_VGND_c_1359_n 0.00288245f $X=-0.19 $Y=-0.245 $X2=3.84 $Y2=0.445
cc_96 VNB N_VGND_c_1360_n 0.00639987f $X=-0.19 $Y=-0.245 $X2=3.03 $Y2=1.79
cc_97 VNB N_VGND_c_1361_n 0.0115604f $X=-0.19 $Y=-0.245 $X2=3.105 $Y2=2.13
cc_98 VNB N_VGND_c_1362_n 0.040836f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.905
cc_99 VNB N_VGND_c_1363_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=2.99
cc_100 VNB N_VGND_c_1364_n 0.0679255f $X=-0.19 $Y=-0.245 $X2=3.312 $Y2=2.905
cc_101 VNB N_VGND_c_1365_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.312 $Y2=2.13
cc_102 VNB N_VGND_c_1366_n 0.0575224f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.13
cc_103 VNB N_VGND_c_1367_n 0.00510891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1368_n 0.0213849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1369_n 0.0188185f $X=-0.19 $Y=-0.245 $X2=4.21 $Y2=1.35
cc_106 VNB N_VGND_c_1370_n 0.479075f $X=-0.19 $Y=-0.245 $X2=4.21 $Y2=1.35
cc_107 VNB N_VGND_c_1371_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=6.155 $Y2=0.465
cc_108 VPB N_A_84_153#_M1004_g 0.0709968f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.735
cc_109 VPB N_A_84_153#_c_185_n 0.0128301f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.7
cc_110 VPB N_A_84_153#_M1015_g 0.0187799f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=2.775
cc_111 VPB N_A_84_153#_M1024_g 0.0201955f $X=-0.19 $Y=1.655 $X2=3.525 $Y2=2.775
cc_112 VPB N_A_84_153#_c_188_n 0.00854292f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.7
cc_113 VPB N_A_84_153#_c_189_n 0.0634419f $X=-0.19 $Y=1.655 $X2=2.955 $Y2=1.79
cc_114 VPB N_A_84_153#_c_205_n 0.0381795f $X=-0.19 $Y=1.655 $X2=3.45 $Y2=2.13
cc_115 VPB N_A_84_153#_c_190_n 0.0106135f $X=-0.19 $Y=1.655 $X2=2.31 $Y2=1.71
cc_116 VPB N_A_84_153#_c_207_n 0.00557266f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=2.905
cc_117 VPB N_A_84_153#_c_208_n 0.0044091f $X=-0.19 $Y=1.655 $X2=3.31 $Y2=2.13
cc_118 VPB N_A_84_153#_c_191_n 0.00376031f $X=-0.19 $Y=1.655 $X2=4.29 $Y2=2.075
cc_119 VPB N_A_84_153#_c_210_n 0.0131759f $X=-0.19 $Y=1.655 $X2=6.58 $Y2=2.16
cc_120 VPB N_A_84_153#_c_211_n 0.0016888f $X=-0.19 $Y=1.655 $X2=6.705 $Y2=2.075
cc_121 VPB N_A_84_153#_c_193_n 0.00133796f $X=-0.19 $Y=1.655 $X2=6.665 $Y2=1.82
cc_122 VPB N_A_84_153#_c_194_n 0.010079f $X=-0.19 $Y=1.655 $X2=1.04 $Y2=1.71
cc_123 VPB N_A_84_153#_c_195_n 0.00389565f $X=-0.19 $Y=1.655 $X2=2.475 $Y2=1.71
cc_124 VPB N_A_84_153#_c_198_n 0.0272647f $X=-0.19 $Y=1.655 $X2=1.04 $Y2=1.7
cc_125 VPB N_D_M1022_g 0.0691894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_226_491#_c_471_n 0.0357621f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.105
cc_127 VPB N_A_226_491#_c_472_n 0.0193983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_226_491#_c_473_n 0.00333304f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=2.775
cc_129 VPB N_A_226_491#_c_474_n 0.00357867f $X=-0.19 $Y=1.655 $X2=3.525
+ $Y2=2.295
cc_130 VPB N_A_226_491#_c_475_n 0.0061641f $X=-0.19 $Y=1.655 $X2=3.525 $Y2=2.775
cc_131 VPB N_A_226_491#_c_476_n 0.0032807f $X=-0.19 $Y=1.655 $X2=3.84 $Y2=0.445
cc_132 VPB N_A_226_491#_c_477_n 0.0398556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_226_491#_c_470_n 0.0156361f $X=-0.19 $Y=1.655 $X2=3.15 $Y2=2.99
cc_134 VPB N_A_114_179#_c_573_n 0.00785461f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=2.775
cc_135 VPB N_A_114_179#_c_574_n 0.00519628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_114_179#_c_585_n 0.0198692f $X=-0.19 $Y=1.655 $X2=3.525 $Y2=2.295
cc_137 VPB N_A_114_179#_M1020_g 0.0295372f $X=-0.19 $Y=1.655 $X2=3.84 $Y2=1.185
cc_138 VPB N_A_114_179#_c_576_n 0.0143636f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=1.79
cc_139 VPB N_A_114_179#_c_588_n 0.0105369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_114_179#_c_580_n 0.0161626f $X=-0.19 $Y=1.655 $X2=4.205 $Y2=2.99
cc_141 VPB N_A_831_21#_M1001_g 0.0350597f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.7
cc_142 VPB N_A_831_21#_c_706_n 0.0109445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_831_21#_c_707_n 0.00271393f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=1.79
cc_144 VPB N_A_831_21#_c_709_n 0.0312065f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=1.955
cc_145 VPB N_GATE_M1026_g 0.0196051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_GATE_c_779_n 0.00780196f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.775
cc_147 VPB N_GATE_c_781_n 0.00241972f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=2.775
cc_148 VPB N_SLEEP_B_M1018_g 0.0222069f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.625
cc_149 VPB N_A_662_47#_M1021_g 0.0226739f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=2.775
cc_150 VPB N_A_662_47#_c_881_n 0.119756f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=2.775
cc_151 VPB N_A_662_47#_c_882_n 0.0169834f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_662_47#_c_868_n 0.0737822f $X=-0.19 $Y=1.655 $X2=3.525 $Y2=2.775
cc_153 VPB N_A_662_47#_c_884_n 0.0344096f $X=-0.19 $Y=1.655 $X2=3.525 $Y2=2.775
cc_154 VPB N_A_662_47#_M1000_g 0.0292253f $X=-0.19 $Y=1.655 $X2=2.955 $Y2=1.79
cc_155 VPB N_A_662_47#_c_886_n 0.00749069f $X=-0.19 $Y=1.655 $X2=2.48 $Y2=2.99
cc_156 VPB N_A_662_47#_c_887_n 0.00282757f $X=-0.19 $Y=1.655 $X2=3.475 $Y2=2.99
cc_157 VPB N_A_662_47#_c_888_n 0.00150946f $X=-0.19 $Y=1.655 $X2=4.29 $Y2=2.075
cc_158 VPB N_A_662_47#_c_877_n 0.00440203f $X=-0.19 $Y=1.655 $X2=6.58 $Y2=0.59
cc_159 VPB N_A_1530_367#_M1008_g 0.0289051f $X=-0.19 $Y=1.655 $X2=0.495
+ $Y2=2.735
cc_160 VPB N_A_1530_367#_c_1033_n 0.0113743f $X=-0.19 $Y=1.655 $X2=3.03
+ $Y2=2.295
cc_161 VPB N_A_1530_367#_c_1029_n 0.00208648f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1084_n 0.0106488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1085_n 0.0354032f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.735
cc_164 VPB N_VPWR_c_1086_n 0.00558649f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.7
cc_165 VPB N_VPWR_c_1087_n 0.0196639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1088_n 0.0323966f $X=-0.19 $Y=1.655 $X2=3.84 $Y2=0.445
cc_167 VPB N_VPWR_c_1089_n 0.161633f $X=-0.19 $Y=1.655 $X2=2.955 $Y2=1.79
cc_168 VPB N_VPWR_c_1090_n 0.0185039f $X=-0.19 $Y=1.655 $X2=2.48 $Y2=2.99
cc_169 VPB N_VPWR_c_1083_n 0.0650118f $X=-0.19 $Y=1.655 $X2=3.312 $Y2=2.905
cc_170 VPB N_VPWR_c_1092_n 0.0063162f $X=-0.19 $Y=1.655 $X2=3.475 $Y2=2.99
cc_171 VPB N_VPWR_c_1093_n 0.00631825f $X=-0.19 $Y=1.655 $X2=4.29 $Y2=2.245
cc_172 VPB N_A_476_47#_c_1176_n 0.0018326f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=2.775
cc_173 VPB N_A_476_47#_c_1177_n 0.00470395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_476_47#_c_1175_n 0.00250392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_KAPWR_c_1242_n 0.00761913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_KAPWR_c_1243_n 0.0280423f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.735
cc_177 VPB N_KAPWR_c_1244_n 0.0167901f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.7
cc_178 VPB N_KAPWR_c_1245_n 0.00521908f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=2.775
cc_179 VPB N_KAPWR_c_1246_n 0.0606338f $X=-0.19 $Y=1.655 $X2=3.03 $Y2=1.79
cc_180 VPB N_KAPWR_c_1247_n 0.0143533f $X=-0.19 $Y=1.655 $X2=2.955 $Y2=1.79
cc_181 VPB N_Q_c_1339_n 0.008411f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.105
cc_182 VPB N_Q_c_1340_n 0.0350919f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.775
cc_183 VPB N_Q_c_1336_n 0.00753674f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.7
cc_184 N_A_84_153#_c_190_n N_D_M1022_g 0.0122101f $X=2.31 $Y=1.71 $X2=0 $Y2=0
cc_185 N_A_84_153#_c_194_n N_D_M1022_g 0.00118187f $X=1.04 $Y=1.71 $X2=0 $Y2=0
cc_186 N_A_84_153#_c_198_n N_D_M1022_g 0.0213066f $X=1.04 $Y=1.7 $X2=0 $Y2=0
cc_187 N_A_84_153#_M1013_g N_D_c_420_n 0.00591664f $X=0.495 $Y=1.105 $X2=0 $Y2=0
cc_188 N_A_84_153#_c_198_n N_D_c_420_n 0.00386649f $X=1.04 $Y=1.7 $X2=0 $Y2=0
cc_189 N_A_84_153#_M1013_g D 4.41487e-19 $X=0.495 $Y=1.105 $X2=0 $Y2=0
cc_190 N_A_84_153#_c_189_n N_A_226_491#_c_471_n 0.035905f $X=2.955 $Y=1.79 $X2=0
+ $Y2=0
cc_191 N_A_84_153#_c_190_n N_A_226_491#_c_471_n 0.00548845f $X=2.31 $Y=1.71
+ $X2=0 $Y2=0
cc_192 N_A_84_153#_c_207_n N_A_226_491#_c_471_n 0.0122433f $X=2.395 $Y=2.905
+ $X2=0 $Y2=0
cc_193 N_A_84_153#_c_225_p N_A_226_491#_c_471_n 6.46131e-19 $X=3.15 $Y=2.99
+ $X2=0 $Y2=0
cc_194 N_A_84_153#_c_195_n N_A_226_491#_c_471_n 0.0011548f $X=2.475 $Y=1.71
+ $X2=0 $Y2=0
cc_195 N_A_84_153#_M1015_g N_A_226_491#_c_472_n 0.0157471f $X=3.03 $Y=2.775
+ $X2=0 $Y2=0
cc_196 N_A_84_153#_c_207_n N_A_226_491#_c_472_n 0.0114889f $X=2.395 $Y=2.905
+ $X2=0 $Y2=0
cc_197 N_A_84_153#_c_225_p N_A_226_491#_c_472_n 0.0119716f $X=3.15 $Y=2.99 $X2=0
+ $Y2=0
cc_198 N_A_84_153#_M1004_g N_A_226_491#_c_473_n 6.59467e-19 $X=0.495 $Y=2.735
+ $X2=0 $Y2=0
cc_199 N_A_84_153#_c_190_n N_A_226_491#_c_474_n 0.00906195f $X=2.31 $Y=1.71
+ $X2=0 $Y2=0
cc_200 N_A_84_153#_c_207_n N_A_226_491#_c_474_n 0.0120957f $X=2.395 $Y=2.905
+ $X2=0 $Y2=0
cc_201 N_A_84_153#_c_190_n N_A_226_491#_c_475_n 0.0076104f $X=2.31 $Y=1.71 $X2=0
+ $Y2=0
cc_202 N_A_84_153#_c_194_n N_A_226_491#_c_475_n 0.00363901f $X=1.04 $Y=1.71
+ $X2=0 $Y2=0
cc_203 N_A_84_153#_c_198_n N_A_226_491#_c_475_n 6.24746e-19 $X=1.04 $Y=1.7 $X2=0
+ $Y2=0
cc_204 N_A_84_153#_c_190_n N_A_226_491#_c_476_n 0.0255244f $X=2.31 $Y=1.71 $X2=0
+ $Y2=0
cc_205 N_A_84_153#_c_207_n N_A_226_491#_c_476_n 0.0304621f $X=2.395 $Y=2.905
+ $X2=0 $Y2=0
cc_206 N_A_84_153#_c_190_n N_A_226_491#_c_477_n 0.00125175f $X=2.31 $Y=1.71
+ $X2=0 $Y2=0
cc_207 N_A_84_153#_c_207_n N_A_226_491#_c_477_n 0.00503937f $X=2.395 $Y=2.905
+ $X2=0 $Y2=0
cc_208 N_A_84_153#_c_189_n N_A_226_491#_c_469_n 7.03598e-19 $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_209 N_A_84_153#_c_189_n N_A_226_491#_c_470_n 0.0129246f $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_210 N_A_84_153#_c_190_n N_A_226_491#_c_470_n 0.0103509f $X=2.31 $Y=1.71 $X2=0
+ $Y2=0
cc_211 N_A_84_153#_c_195_n N_A_226_491#_c_470_n 0.00366586f $X=2.475 $Y=1.71
+ $X2=0 $Y2=0
cc_212 N_A_84_153#_c_189_n N_A_114_179#_c_570_n 0.013731f $X=2.955 $Y=1.79 $X2=0
+ $Y2=0
cc_213 N_A_84_153#_c_205_n N_A_114_179#_c_570_n 0.00360282f $X=3.45 $Y=2.13
+ $X2=0 $Y2=0
cc_214 N_A_84_153#_M1006_g N_A_114_179#_M1003_g 0.0197973f $X=3.84 $Y=0.445
+ $X2=0 $Y2=0
cc_215 N_A_84_153#_c_189_n N_A_114_179#_c_574_n 0.00538577f $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_216 N_A_84_153#_c_205_n N_A_114_179#_c_574_n 0.0121975f $X=3.45 $Y=2.13 $X2=0
+ $Y2=0
cc_217 N_A_84_153#_c_208_n N_A_114_179#_c_574_n 9.25755e-19 $X=3.31 $Y=2.13
+ $X2=0 $Y2=0
cc_218 N_A_84_153#_c_186_n N_A_114_179#_c_585_n 0.0214984f $X=3.84 $Y=1.185
+ $X2=0 $Y2=0
cc_219 N_A_84_153#_c_191_n N_A_114_179#_c_585_n 0.0048861f $X=4.29 $Y=2.075
+ $X2=0 $Y2=0
cc_220 N_A_84_153#_c_196_n N_A_114_179#_c_585_n 0.00122569f $X=4.21 $Y=1.35
+ $X2=0 $Y2=0
cc_221 N_A_84_153#_c_205_n N_A_114_179#_M1020_g 0.0286778f $X=3.45 $Y=2.13 $X2=0
+ $Y2=0
cc_222 N_A_84_153#_c_208_n N_A_114_179#_M1020_g 0.00145852f $X=3.31 $Y=2.13
+ $X2=0 $Y2=0
cc_223 N_A_84_153#_c_255_p N_A_114_179#_M1020_g 0.0142836f $X=4.205 $Y=2.99
+ $X2=0 $Y2=0
cc_224 N_A_84_153#_c_191_n N_A_114_179#_M1020_g 0.00485587f $X=4.29 $Y=2.075
+ $X2=0 $Y2=0
cc_225 N_A_84_153#_c_257_p N_A_114_179#_M1020_g 0.0162083f $X=4.29 $Y=2.905
+ $X2=0 $Y2=0
cc_226 N_A_84_153#_c_258_p N_A_114_179#_M1020_g 0.00490948f $X=4.29 $Y=2.16
+ $X2=0 $Y2=0
cc_227 N_A_84_153#_c_186_n N_A_114_179#_c_575_n 0.00739409f $X=3.84 $Y=1.185
+ $X2=0 $Y2=0
cc_228 N_A_84_153#_c_208_n N_A_114_179#_c_575_n 3.07471e-19 $X=3.31 $Y=2.13
+ $X2=0 $Y2=0
cc_229 N_A_84_153#_c_186_n N_A_114_179#_c_576_n 0.00386389f $X=3.84 $Y=1.185
+ $X2=0 $Y2=0
cc_230 N_A_84_153#_c_189_n N_A_114_179#_c_576_n 0.00319482f $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_231 N_A_84_153#_c_191_n N_A_114_179#_c_576_n 8.61869e-19 $X=4.29 $Y=2.075
+ $X2=0 $Y2=0
cc_232 N_A_84_153#_M1013_g N_A_114_179#_c_577_n 0.00656956f $X=0.495 $Y=1.105
+ $X2=0 $Y2=0
cc_233 N_A_84_153#_c_185_n N_A_114_179#_c_578_n 0.00274226f $X=0.875 $Y=1.7
+ $X2=0 $Y2=0
cc_234 N_A_84_153#_c_189_n N_A_114_179#_c_578_n 0.00196908f $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_235 N_A_84_153#_c_190_n N_A_114_179#_c_578_n 0.0809511f $X=2.31 $Y=1.71 $X2=0
+ $Y2=0
cc_236 N_A_84_153#_c_194_n N_A_114_179#_c_578_n 0.0247729f $X=1.04 $Y=1.71 $X2=0
+ $Y2=0
cc_237 N_A_84_153#_c_195_n N_A_114_179#_c_578_n 0.0240978f $X=2.475 $Y=1.71
+ $X2=0 $Y2=0
cc_238 N_A_84_153#_c_198_n N_A_114_179#_c_578_n 0.00159846f $X=1.04 $Y=1.7 $X2=0
+ $Y2=0
cc_239 N_A_84_153#_M1013_g N_A_114_179#_c_579_n 0.0100628f $X=0.495 $Y=1.105
+ $X2=0 $Y2=0
cc_240 N_A_84_153#_c_185_n N_A_114_179#_c_579_n 0.0035961f $X=0.875 $Y=1.7 $X2=0
+ $Y2=0
cc_241 N_A_84_153#_M1004_g N_A_114_179#_c_588_n 0.00769019f $X=0.495 $Y=2.735
+ $X2=0 $Y2=0
cc_242 N_A_84_153#_c_185_n N_A_114_179#_c_588_n 0.00432518f $X=0.875 $Y=1.7
+ $X2=0 $Y2=0
cc_243 N_A_84_153#_M1013_g N_A_114_179#_c_580_n 0.00977678f $X=0.495 $Y=1.105
+ $X2=0 $Y2=0
cc_244 N_A_84_153#_M1004_g N_A_114_179#_c_580_n 0.0342773f $X=0.495 $Y=2.735
+ $X2=0 $Y2=0
cc_245 N_A_84_153#_c_185_n N_A_114_179#_c_580_n 0.0103261f $X=0.875 $Y=1.7 $X2=0
+ $Y2=0
cc_246 N_A_84_153#_c_188_n N_A_114_179#_c_580_n 0.00617699f $X=0.495 $Y=1.7
+ $X2=0 $Y2=0
cc_247 N_A_84_153#_c_194_n N_A_114_179#_c_580_n 0.0242401f $X=1.04 $Y=1.71 $X2=0
+ $Y2=0
cc_248 N_A_84_153#_c_198_n N_A_114_179#_c_580_n 0.00117139f $X=1.04 $Y=1.7 $X2=0
+ $Y2=0
cc_249 N_A_84_153#_c_189_n N_A_114_179#_c_581_n 0.00513175f $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_250 N_A_84_153#_c_195_n N_A_114_179#_c_581_n 0.00146077f $X=2.475 $Y=1.71
+ $X2=0 $Y2=0
cc_251 N_A_84_153#_c_189_n N_A_114_179#_c_582_n 0.013731f $X=2.955 $Y=1.79 $X2=0
+ $Y2=0
cc_252 N_A_84_153#_c_210_n N_A_831_21#_M1021_s 0.00715571f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_253 N_A_84_153#_M1006_g N_A_831_21#_M1007_g 0.0462131f $X=3.84 $Y=0.445 $X2=0
+ $Y2=0
cc_254 N_A_84_153#_c_186_n N_A_831_21#_c_702_n 0.0121273f $X=3.84 $Y=1.185 $X2=0
+ $Y2=0
cc_255 N_A_84_153#_c_196_n N_A_831_21#_c_702_n 2.3783e-19 $X=4.21 $Y=1.35 $X2=0
+ $Y2=0
cc_256 N_A_84_153#_c_255_p N_A_831_21#_M1001_g 0.00161295f $X=4.205 $Y=2.99
+ $X2=0 $Y2=0
cc_257 N_A_84_153#_c_257_p N_A_831_21#_M1001_g 0.00741802f $X=4.29 $Y=2.905
+ $X2=0 $Y2=0
cc_258 N_A_84_153#_c_210_n N_A_831_21#_M1001_g 0.0208408f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_259 N_A_84_153#_c_186_n N_A_831_21#_c_704_n 0.0217281f $X=3.84 $Y=1.185 $X2=0
+ $Y2=0
cc_260 N_A_84_153#_M1006_g N_A_831_21#_c_704_n 0.00459277f $X=3.84 $Y=0.445
+ $X2=0 $Y2=0
cc_261 N_A_84_153#_c_191_n N_A_831_21#_c_704_n 0.00197078f $X=4.29 $Y=2.075
+ $X2=0 $Y2=0
cc_262 N_A_84_153#_c_196_n N_A_831_21#_c_704_n 0.00220005f $X=4.21 $Y=1.35 $X2=0
+ $Y2=0
cc_263 N_A_84_153#_c_191_n N_A_831_21#_c_706_n 0.0223345f $X=4.29 $Y=2.075 $X2=0
+ $Y2=0
cc_264 N_A_84_153#_c_210_n N_A_831_21#_c_706_n 0.0658204f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_265 N_A_84_153#_c_210_n N_A_831_21#_c_707_n 0.00897969f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_266 N_A_84_153#_c_197_n N_A_831_21#_c_708_n 0.0283157f $X=6.155 $Y=0.465
+ $X2=0 $Y2=0
cc_267 N_A_84_153#_c_191_n N_A_831_21#_c_709_n 0.00594588f $X=4.29 $Y=2.075
+ $X2=0 $Y2=0
cc_268 N_A_84_153#_c_210_n N_A_831_21#_c_709_n 0.0040357f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_269 N_A_84_153#_c_210_n N_GATE_M1026_g 0.0121708f $X=6.58 $Y=2.16 $X2=0 $Y2=0
cc_270 N_A_84_153#_c_211_n N_GATE_M1026_g 0.0020738f $X=6.705 $Y=2.075 $X2=0
+ $Y2=0
cc_271 N_A_84_153#_c_193_n N_GATE_M1026_g 0.00769832f $X=6.665 $Y=1.82 $X2=0
+ $Y2=0
cc_272 N_A_84_153#_c_192_n N_GATE_M1023_g 0.0091533f $X=6.58 $Y=0.59 $X2=0 $Y2=0
cc_273 N_A_84_153#_c_193_n N_GATE_M1023_g 0.00862558f $X=6.665 $Y=1.82 $X2=0
+ $Y2=0
cc_274 N_A_84_153#_c_197_n N_GATE_M1023_g 0.00642652f $X=6.155 $Y=0.465 $X2=0
+ $Y2=0
cc_275 N_A_84_153#_c_210_n N_GATE_c_779_n 0.00110294f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_276 N_A_84_153#_c_197_n N_GATE_c_780_n 0.00160731f $X=6.155 $Y=0.465 $X2=0
+ $Y2=0
cc_277 N_A_84_153#_c_210_n N_GATE_c_781_n 0.022554f $X=6.58 $Y=2.16 $X2=0 $Y2=0
cc_278 N_A_84_153#_c_192_n N_GATE_c_781_n 0.00659917f $X=6.58 $Y=0.59 $X2=0
+ $Y2=0
cc_279 N_A_84_153#_c_193_n N_GATE_c_781_n 0.0711678f $X=6.665 $Y=1.82 $X2=0
+ $Y2=0
cc_280 N_A_84_153#_c_197_n N_GATE_c_781_n 0.0277968f $X=6.155 $Y=0.465 $X2=0
+ $Y2=0
cc_281 N_A_84_153#_c_192_n N_SLEEP_B_M1017_g 0.00705548f $X=6.58 $Y=0.59 $X2=0
+ $Y2=0
cc_282 N_A_84_153#_c_193_n N_SLEEP_B_M1017_g 0.00546096f $X=6.665 $Y=1.82 $X2=0
+ $Y2=0
cc_283 N_A_84_153#_c_197_n N_SLEEP_B_M1017_g 0.00133263f $X=6.155 $Y=0.465 $X2=0
+ $Y2=0
cc_284 N_A_84_153#_c_211_n N_SLEEP_B_M1018_g 0.00312633f $X=6.705 $Y=2.075 $X2=0
+ $Y2=0
cc_285 N_A_84_153#_c_193_n N_SLEEP_B_M1018_g 0.0190621f $X=6.665 $Y=1.82 $X2=0
+ $Y2=0
cc_286 N_A_84_153#_c_192_n N_SLEEP_B_c_821_n 8.45271e-19 $X=6.58 $Y=0.59 $X2=0
+ $Y2=0
cc_287 N_A_84_153#_c_193_n N_SLEEP_B_c_821_n 0.00308424f $X=6.665 $Y=1.82 $X2=0
+ $Y2=0
cc_288 N_A_84_153#_c_193_n SLEEP_B 0.0473771f $X=6.665 $Y=1.82 $X2=0 $Y2=0
cc_289 N_A_84_153#_c_193_n N_SLEEP_B_c_823_n 0.008947f $X=6.665 $Y=1.82 $X2=0
+ $Y2=0
cc_290 N_A_84_153#_c_255_p N_A_662_47#_M1024_d 0.00470752f $X=4.205 $Y=2.99
+ $X2=0 $Y2=0
cc_291 N_A_84_153#_c_197_n N_A_662_47#_M1005_g 8.05639e-19 $X=6.155 $Y=0.465
+ $X2=0 $Y2=0
cc_292 N_A_84_153#_c_210_n N_A_662_47#_M1021_g 0.0264876f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_293 N_A_84_153#_c_210_n N_A_662_47#_c_881_n 7.78776e-19 $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_294 N_A_84_153#_c_193_n N_A_662_47#_c_873_n 0.00124368f $X=6.665 $Y=1.82
+ $X2=0 $Y2=0
cc_295 N_A_84_153#_M1006_g N_A_662_47#_c_874_n 0.0134732f $X=3.84 $Y=0.445 $X2=0
+ $Y2=0
cc_296 N_A_84_153#_c_205_n N_A_662_47#_c_887_n 0.00275551f $X=3.45 $Y=2.13 $X2=0
+ $Y2=0
cc_297 N_A_84_153#_c_258_p N_A_662_47#_c_887_n 0.0126407f $X=4.29 $Y=2.16 $X2=0
+ $Y2=0
cc_298 N_A_84_153#_M1024_g N_A_662_47#_c_888_n 0.00275551f $X=3.525 $Y=2.775
+ $X2=0 $Y2=0
cc_299 N_A_84_153#_c_255_p N_A_662_47#_c_888_n 0.0209818f $X=4.205 $Y=2.99 $X2=0
+ $Y2=0
cc_300 N_A_84_153#_c_257_p N_A_662_47#_c_888_n 0.0322178f $X=4.29 $Y=2.905 $X2=0
+ $Y2=0
cc_301 N_A_84_153#_c_186_n N_A_662_47#_c_875_n 0.00591794f $X=3.84 $Y=1.185
+ $X2=0 $Y2=0
cc_302 N_A_84_153#_M1006_g N_A_662_47#_c_875_n 0.00673985f $X=3.84 $Y=0.445
+ $X2=0 $Y2=0
cc_303 N_A_84_153#_c_196_n N_A_662_47#_c_875_n 0.0255146f $X=4.21 $Y=1.35 $X2=0
+ $Y2=0
cc_304 N_A_84_153#_M1006_g N_A_662_47#_c_876_n 0.00587054f $X=3.84 $Y=0.445
+ $X2=0 $Y2=0
cc_305 N_A_84_153#_c_186_n N_A_662_47#_c_877_n 0.00717966f $X=3.84 $Y=1.185
+ $X2=0 $Y2=0
cc_306 N_A_84_153#_M1006_g N_A_662_47#_c_877_n 0.0092114f $X=3.84 $Y=0.445 $X2=0
+ $Y2=0
cc_307 N_A_84_153#_c_189_n N_A_662_47#_c_877_n 0.00302335f $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_308 N_A_84_153#_c_205_n N_A_662_47#_c_877_n 0.00172187f $X=3.45 $Y=2.13 $X2=0
+ $Y2=0
cc_309 N_A_84_153#_c_208_n N_A_662_47#_c_877_n 0.049415f $X=3.31 $Y=2.13 $X2=0
+ $Y2=0
cc_310 N_A_84_153#_c_191_n N_A_662_47#_c_877_n 0.0238137f $X=4.29 $Y=2.075 $X2=0
+ $Y2=0
cc_311 N_A_84_153#_c_196_n N_A_662_47#_c_877_n 0.0227038f $X=4.21 $Y=1.35 $X2=0
+ $Y2=0
cc_312 N_A_84_153#_c_207_n N_VPWR_M1022_d 0.00938163f $X=2.395 $Y=2.905 $X2=0
+ $Y2=0
cc_313 N_A_84_153#_c_345_p N_VPWR_M1022_d 0.00432904f $X=2.48 $Y=2.99 $X2=0
+ $Y2=0
cc_314 N_A_84_153#_M1004_g N_VPWR_c_1085_n 0.00502318f $X=0.495 $Y=2.735 $X2=0
+ $Y2=0
cc_315 N_A_84_153#_c_207_n N_VPWR_c_1086_n 0.00387428f $X=2.395 $Y=2.905 $X2=0
+ $Y2=0
cc_316 N_A_84_153#_c_345_p N_VPWR_c_1086_n 0.00745042f $X=2.48 $Y=2.99 $X2=0
+ $Y2=0
cc_317 N_A_84_153#_M1004_g N_VPWR_c_1088_n 0.00497111f $X=0.495 $Y=2.735 $X2=0
+ $Y2=0
cc_318 N_A_84_153#_M1015_g N_VPWR_c_1089_n 0.00357877f $X=3.03 $Y=2.775 $X2=0
+ $Y2=0
cc_319 N_A_84_153#_M1024_g N_VPWR_c_1089_n 0.00357842f $X=3.525 $Y=2.775 $X2=0
+ $Y2=0
cc_320 N_A_84_153#_c_225_p N_VPWR_c_1089_n 0.0361696f $X=3.15 $Y=2.99 $X2=0
+ $Y2=0
cc_321 N_A_84_153#_c_345_p N_VPWR_c_1089_n 0.0115003f $X=2.48 $Y=2.99 $X2=0
+ $Y2=0
cc_322 N_A_84_153#_c_255_p N_VPWR_c_1089_n 0.0522343f $X=4.205 $Y=2.99 $X2=0
+ $Y2=0
cc_323 N_A_84_153#_c_355_p N_VPWR_c_1089_n 0.020362f $X=3.312 $Y=2.99 $X2=0
+ $Y2=0
cc_324 N_A_84_153#_M1004_g N_VPWR_c_1083_n 0.00643301f $X=0.495 $Y=2.735 $X2=0
+ $Y2=0
cc_325 N_A_84_153#_M1015_g N_VPWR_c_1083_n 0.00502013f $X=3.03 $Y=2.775 $X2=0
+ $Y2=0
cc_326 N_A_84_153#_M1024_g N_VPWR_c_1083_n 0.00529158f $X=3.525 $Y=2.775 $X2=0
+ $Y2=0
cc_327 N_A_84_153#_c_225_p N_VPWR_c_1083_n 0.00513225f $X=3.15 $Y=2.99 $X2=0
+ $Y2=0
cc_328 N_A_84_153#_c_345_p N_VPWR_c_1083_n 0.00158693f $X=2.48 $Y=2.99 $X2=0
+ $Y2=0
cc_329 N_A_84_153#_c_255_p N_VPWR_c_1083_n 0.00713478f $X=4.205 $Y=2.99 $X2=0
+ $Y2=0
cc_330 N_A_84_153#_c_355_p N_VPWR_c_1083_n 0.00301708f $X=3.312 $Y=2.99 $X2=0
+ $Y2=0
cc_331 N_A_84_153#_c_225_p N_A_476_47#_M1012_d 0.00234113f $X=3.15 $Y=2.99 $X2=0
+ $Y2=0
cc_332 N_A_84_153#_M1006_g N_A_476_47#_c_1173_n 6.14494e-19 $X=3.84 $Y=0.445
+ $X2=0 $Y2=0
cc_333 N_A_84_153#_M1015_g N_A_476_47#_c_1176_n 0.00303902f $X=3.03 $Y=2.775
+ $X2=0 $Y2=0
cc_334 N_A_84_153#_c_189_n N_A_476_47#_c_1176_n 0.00395295f $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_335 N_A_84_153#_c_207_n N_A_476_47#_c_1176_n 0.0119845f $X=2.395 $Y=2.905
+ $X2=0 $Y2=0
cc_336 N_A_84_153#_c_225_p N_A_476_47#_c_1176_n 0.0189111f $X=3.15 $Y=2.99 $X2=0
+ $Y2=0
cc_337 N_A_84_153#_M1015_g N_A_476_47#_c_1177_n 0.00260157f $X=3.03 $Y=2.775
+ $X2=0 $Y2=0
cc_338 N_A_84_153#_M1024_g N_A_476_47#_c_1177_n 3.27735e-19 $X=3.525 $Y=2.775
+ $X2=0 $Y2=0
cc_339 N_A_84_153#_c_189_n N_A_476_47#_c_1177_n 0.0258401f $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_340 N_A_84_153#_c_207_n N_A_476_47#_c_1177_n 0.0226608f $X=2.395 $Y=2.905
+ $X2=0 $Y2=0
cc_341 N_A_84_153#_c_208_n N_A_476_47#_c_1177_n 0.0468206f $X=3.31 $Y=2.13 $X2=0
+ $Y2=0
cc_342 N_A_84_153#_c_195_n N_A_476_47#_c_1177_n 0.011426f $X=2.475 $Y=1.71 $X2=0
+ $Y2=0
cc_343 N_A_84_153#_c_189_n N_A_476_47#_c_1175_n 0.0173013f $X=2.955 $Y=1.79
+ $X2=0 $Y2=0
cc_344 N_A_84_153#_c_205_n N_A_476_47#_c_1175_n 0.00174555f $X=3.45 $Y=2.13
+ $X2=0 $Y2=0
cc_345 N_A_84_153#_c_208_n N_A_476_47#_c_1175_n 0.0111083f $X=3.31 $Y=2.13 $X2=0
+ $Y2=0
cc_346 N_A_84_153#_c_195_n N_A_476_47#_c_1175_n 0.0130452f $X=2.475 $Y=1.71
+ $X2=0 $Y2=0
cc_347 N_A_84_153#_c_208_n A_621_491# 0.00150044f $X=3.31 $Y=2.13 $X2=-0.19
+ $Y2=-0.245
cc_348 N_A_84_153#_c_355_p A_621_491# 0.00225871f $X=3.312 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_349 N_A_84_153#_c_255_p A_849_419# 0.00251825f $X=4.205 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_350 N_A_84_153#_c_257_p A_849_419# 0.00668156f $X=4.29 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_351 N_A_84_153#_c_210_n A_849_419# 8.93923e-19 $X=6.58 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_352 N_A_84_153#_c_210_n N_KAPWR_M1001_d 0.00321751f $X=6.58 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_353 N_A_84_153#_c_210_n N_KAPWR_M1021_d 0.00672024f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_354 N_A_84_153#_c_210_n N_KAPWR_c_1242_n 0.0128679f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_355 N_A_84_153#_c_210_n N_KAPWR_c_1243_n 0.0174838f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_356 N_A_84_153#_c_211_n N_KAPWR_c_1243_n 0.0177264f $X=6.705 $Y=2.075 $X2=0
+ $Y2=0
cc_357 N_A_84_153#_c_211_n N_KAPWR_c_1244_n 0.0112106f $X=6.705 $Y=2.075 $X2=0
+ $Y2=0
cc_358 N_A_84_153#_c_193_n N_KAPWR_c_1244_n 0.0158575f $X=6.665 $Y=1.82 $X2=0
+ $Y2=0
cc_359 N_A_84_153#_c_210_n N_KAPWR_c_1245_n 0.0204088f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_360 N_A_84_153#_M1004_g N_KAPWR_c_1246_n 0.00570827f $X=0.495 $Y=2.735 $X2=0
+ $Y2=0
cc_361 N_A_84_153#_M1015_g N_KAPWR_c_1246_n 0.00780991f $X=3.03 $Y=2.775 $X2=0
+ $Y2=0
cc_362 N_A_84_153#_M1024_g N_KAPWR_c_1246_n 0.00691921f $X=3.525 $Y=2.775 $X2=0
+ $Y2=0
cc_363 N_A_84_153#_c_207_n N_KAPWR_c_1246_n 0.0194873f $X=2.395 $Y=2.905 $X2=0
+ $Y2=0
cc_364 N_A_84_153#_c_225_p N_KAPWR_c_1246_n 0.0185991f $X=3.15 $Y=2.99 $X2=0
+ $Y2=0
cc_365 N_A_84_153#_c_345_p N_KAPWR_c_1246_n 0.00284371f $X=2.48 $Y=2.99 $X2=0
+ $Y2=0
cc_366 N_A_84_153#_c_208_n N_KAPWR_c_1246_n 0.0322625f $X=3.31 $Y=2.13 $X2=0
+ $Y2=0
cc_367 N_A_84_153#_c_255_p N_KAPWR_c_1246_n 0.0232083f $X=4.205 $Y=2.99 $X2=0
+ $Y2=0
cc_368 N_A_84_153#_c_257_p N_KAPWR_c_1246_n 0.0226674f $X=4.29 $Y=2.905 $X2=0
+ $Y2=0
cc_369 N_A_84_153#_c_210_n N_KAPWR_c_1246_n 0.0315671f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_370 N_A_84_153#_c_211_n N_KAPWR_c_1246_n 0.00148909f $X=6.705 $Y=2.075 $X2=0
+ $Y2=0
cc_371 N_A_84_153#_c_355_p N_KAPWR_c_1246_n 0.00407551f $X=3.312 $Y=2.99 $X2=0
+ $Y2=0
cc_372 N_A_84_153#_c_255_p N_KAPWR_c_1247_n 0.00775792f $X=4.205 $Y=2.99 $X2=0
+ $Y2=0
cc_373 N_A_84_153#_c_257_p N_KAPWR_c_1247_n 0.0189043f $X=4.29 $Y=2.905 $X2=0
+ $Y2=0
cc_374 N_A_84_153#_c_210_n N_KAPWR_c_1247_n 0.0303449f $X=6.58 $Y=2.16 $X2=0
+ $Y2=0
cc_375 N_A_84_153#_M1013_g N_VGND_c_1357_n 0.00482327f $X=0.495 $Y=1.105 $X2=0
+ $Y2=0
cc_376 N_A_84_153#_M1013_g N_VGND_c_1362_n 0.00297774f $X=0.495 $Y=1.105 $X2=0
+ $Y2=0
cc_377 N_A_84_153#_M1006_g N_VGND_c_1364_n 0.0054895f $X=3.84 $Y=0.445 $X2=0
+ $Y2=0
cc_378 N_A_84_153#_c_192_n N_VGND_c_1366_n 0.0108219f $X=6.58 $Y=0.59 $X2=0
+ $Y2=0
cc_379 N_A_84_153#_c_197_n N_VGND_c_1366_n 0.0204006f $X=6.155 $Y=0.465 $X2=0
+ $Y2=0
cc_380 N_A_84_153#_M1023_s N_VGND_c_1370_n 0.00232718f $X=6.01 $Y=0.235 $X2=0
+ $Y2=0
cc_381 N_A_84_153#_M1013_g N_VGND_c_1370_n 0.00400849f $X=0.495 $Y=1.105 $X2=0
+ $Y2=0
cc_382 N_A_84_153#_M1006_g N_VGND_c_1370_n 0.00668652f $X=3.84 $Y=0.445 $X2=0
+ $Y2=0
cc_383 N_A_84_153#_c_192_n N_VGND_c_1370_n 0.0151606f $X=6.58 $Y=0.59 $X2=0
+ $Y2=0
cc_384 N_A_84_153#_c_197_n N_VGND_c_1370_n 0.0124872f $X=6.155 $Y=0.465 $X2=0
+ $Y2=0
cc_385 N_A_84_153#_c_192_n A_1289_47# 0.00140799f $X=6.58 $Y=0.59 $X2=-0.19
+ $Y2=-0.245
cc_386 N_D_M1014_g N_A_226_491#_c_465_n 0.00905596f $X=1.545 $Y=0.445 $X2=0
+ $Y2=0
cc_387 N_D_M1022_g N_A_226_491#_c_473_n 0.0104312f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_388 N_D_M1022_g N_A_226_491#_c_474_n 0.0120962f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_389 N_D_M1022_g N_A_226_491#_c_475_n 0.00364124f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_390 N_D_M1022_g N_A_226_491#_c_476_n 0.00571191f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_391 N_D_M1022_g N_A_226_491#_c_477_n 0.0250933f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_392 N_D_M1014_g N_A_226_491#_c_467_n 0.0215898f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_393 N_D_c_420_n N_A_226_491#_c_467_n 0.00759333f $X=1.415 $Y=0.95 $X2=0 $Y2=0
cc_394 N_D_c_421_n N_A_226_491#_c_467_n 0.00303099f $X=1.415 $Y=0.785 $X2=0
+ $Y2=0
cc_395 D N_A_226_491#_c_467_n 0.0114718f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_396 N_D_M1014_g N_A_226_491#_c_468_n 2.55261e-19 $X=1.545 $Y=0.445 $X2=0
+ $Y2=0
cc_397 N_D_c_421_n N_A_226_491#_c_468_n 0.0015036f $X=1.415 $Y=0.785 $X2=0 $Y2=0
cc_398 D N_A_226_491#_c_468_n 0.00892814f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_399 N_D_M1014_g N_A_226_491#_c_469_n 0.0100141f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_400 N_D_c_421_n N_A_226_491#_c_469_n 0.0232949f $X=1.415 $Y=0.785 $X2=0 $Y2=0
cc_401 D N_A_226_491#_c_469_n 8.79005e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_402 N_D_M1022_g N_A_226_491#_c_470_n 0.0232949f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_403 N_D_M1022_g N_A_114_179#_c_577_n 0.00381924f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_404 N_D_c_420_n N_A_114_179#_c_577_n 9.06786e-19 $X=1.415 $Y=0.95 $X2=0 $Y2=0
cc_405 D N_A_114_179#_c_577_n 0.0168252f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_406 N_D_M1022_g N_A_114_179#_c_578_n 0.0143563f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_407 N_D_c_420_n N_A_114_179#_c_578_n 0.0071327f $X=1.415 $Y=0.95 $X2=0 $Y2=0
cc_408 N_D_c_421_n N_A_114_179#_c_578_n 0.00132179f $X=1.415 $Y=0.785 $X2=0
+ $Y2=0
cc_409 D N_A_114_179#_c_578_n 0.0248017f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_410 N_D_M1022_g N_A_114_179#_c_588_n 0.00247337f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_411 N_D_M1022_g N_VPWR_c_1086_n 0.010618f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_412 N_D_M1022_g N_VPWR_c_1088_n 0.00426006f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_413 N_D_M1022_g N_VPWR_c_1083_n 0.00768781f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_414 N_D_M1022_g N_KAPWR_c_1246_n 0.00619908f $X=1.49 $Y=2.775 $X2=0 $Y2=0
cc_415 D N_VGND_c_1357_n 0.00256299f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_416 N_D_M1014_g N_VGND_c_1358_n 0.00362591f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_417 N_D_M1014_g N_VGND_c_1362_n 0.00357668f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_418 N_D_M1014_g N_VGND_c_1370_n 0.00740789f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_419 N_D_c_420_n N_VGND_c_1370_n 0.00421544f $X=1.415 $Y=0.95 $X2=0 $Y2=0
cc_420 D N_VGND_c_1370_n 0.00648315f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_421 N_A_226_491#_c_465_n N_A_114_179#_M1002_g 0.0176273f $X=2.305 $Y=0.765
+ $X2=0 $Y2=0
cc_422 N_A_226_491#_c_468_n N_A_114_179#_M1002_g 0.00130573f $X=2.025 $Y=0.7
+ $X2=0 $Y2=0
cc_423 N_A_226_491#_c_469_n N_A_114_179#_M1002_g 0.00299518f $X=2.025 $Y=0.93
+ $X2=0 $Y2=0
cc_424 N_A_226_491#_c_466_n N_A_114_179#_c_578_n 0.00730044f $X=1.86 $Y=0.7
+ $X2=0 $Y2=0
cc_425 N_A_226_491#_c_467_n N_A_114_179#_c_578_n 0.00949484f $X=1.33 $Y=0.435
+ $X2=0 $Y2=0
cc_426 N_A_226_491#_c_468_n N_A_114_179#_c_578_n 0.0228712f $X=2.025 $Y=0.7
+ $X2=0 $Y2=0
cc_427 N_A_226_491#_c_469_n N_A_114_179#_c_578_n 0.00639981f $X=2.025 $Y=0.93
+ $X2=0 $Y2=0
cc_428 N_A_226_491#_c_470_n N_A_114_179#_c_578_n 0.012165f $X=1.94 $Y=1.965
+ $X2=0 $Y2=0
cc_429 N_A_226_491#_c_473_n N_A_114_179#_c_588_n 0.027449f $X=1.275 $Y=2.755
+ $X2=0 $Y2=0
cc_430 N_A_226_491#_c_475_n N_A_114_179#_c_588_n 0.0119736f $X=1.44 $Y=2.52
+ $X2=0 $Y2=0
cc_431 N_A_226_491#_c_468_n N_A_114_179#_c_581_n 0.00141768f $X=2.025 $Y=0.7
+ $X2=0 $Y2=0
cc_432 N_A_226_491#_c_470_n N_A_114_179#_c_581_n 0.00113096f $X=1.94 $Y=1.965
+ $X2=0 $Y2=0
cc_433 N_A_226_491#_c_469_n N_A_114_179#_c_582_n 0.00101665f $X=2.025 $Y=0.93
+ $X2=0 $Y2=0
cc_434 N_A_226_491#_c_470_n N_A_114_179#_c_582_n 0.00548518f $X=1.94 $Y=1.965
+ $X2=0 $Y2=0
cc_435 N_A_226_491#_c_474_n N_VPWR_M1022_d 0.00897404f $X=1.775 $Y=2.52 $X2=0
+ $Y2=0
cc_436 N_A_226_491#_c_472_n N_VPWR_c_1086_n 0.00304924f $X=2.6 $Y=2.345 $X2=0
+ $Y2=0
cc_437 N_A_226_491#_c_473_n N_VPWR_c_1086_n 0.0134857f $X=1.275 $Y=2.755 $X2=0
+ $Y2=0
cc_438 N_A_226_491#_c_474_n N_VPWR_c_1086_n 0.021586f $X=1.775 $Y=2.52 $X2=0
+ $Y2=0
cc_439 N_A_226_491#_c_477_n N_VPWR_c_1086_n 5.85992e-19 $X=1.94 $Y=2.13 $X2=0
+ $Y2=0
cc_440 N_A_226_491#_c_473_n N_VPWR_c_1088_n 0.0209673f $X=1.275 $Y=2.755 $X2=0
+ $Y2=0
cc_441 N_A_226_491#_c_474_n N_VPWR_c_1088_n 0.00177689f $X=1.775 $Y=2.52 $X2=0
+ $Y2=0
cc_442 N_A_226_491#_c_472_n N_VPWR_c_1089_n 0.00357877f $X=2.6 $Y=2.345 $X2=0
+ $Y2=0
cc_443 N_A_226_491#_c_474_n N_VPWR_c_1089_n 0.00218011f $X=1.775 $Y=2.52 $X2=0
+ $Y2=0
cc_444 N_A_226_491#_M1022_s N_VPWR_c_1083_n 0.00119809f $X=1.13 $Y=2.455 $X2=0
+ $Y2=0
cc_445 N_A_226_491#_c_472_n N_VPWR_c_1083_n 0.00624787f $X=2.6 $Y=2.345 $X2=0
+ $Y2=0
cc_446 N_A_226_491#_c_473_n N_VPWR_c_1083_n 0.00303603f $X=1.275 $Y=2.755 $X2=0
+ $Y2=0
cc_447 N_A_226_491#_c_465_n N_A_476_47#_c_1174_n 0.011054f $X=2.305 $Y=0.765
+ $X2=0 $Y2=0
cc_448 N_A_226_491#_c_468_n N_A_476_47#_c_1174_n 0.00304184f $X=2.025 $Y=0.7
+ $X2=0 $Y2=0
cc_449 N_A_226_491#_c_472_n N_A_476_47#_c_1176_n 0.00356654f $X=2.6 $Y=2.345
+ $X2=0 $Y2=0
cc_450 N_A_226_491#_c_471_n N_A_476_47#_c_1177_n 0.00218424f $X=2.525 $Y=2.27
+ $X2=0 $Y2=0
cc_451 N_A_226_491#_c_472_n N_KAPWR_c_1246_n 0.00925987f $X=2.6 $Y=2.345 $X2=0
+ $Y2=0
cc_452 N_A_226_491#_c_473_n N_KAPWR_c_1246_n 0.0363334f $X=1.275 $Y=2.755 $X2=0
+ $Y2=0
cc_453 N_A_226_491#_c_474_n N_KAPWR_c_1246_n 0.0235788f $X=1.775 $Y=2.52 $X2=0
+ $Y2=0
cc_454 N_A_226_491#_c_477_n N_KAPWR_c_1246_n 0.0053823f $X=1.94 $Y=2.13 $X2=0
+ $Y2=0
cc_455 N_A_226_491#_c_466_n N_VGND_M1014_d 0.00296385f $X=1.86 $Y=0.7 $X2=0
+ $Y2=0
cc_456 N_A_226_491#_c_468_n N_VGND_M1014_d 0.00348441f $X=2.025 $Y=0.7 $X2=0
+ $Y2=0
cc_457 N_A_226_491#_c_465_n N_VGND_c_1358_n 0.00582901f $X=2.305 $Y=0.765 $X2=0
+ $Y2=0
cc_458 N_A_226_491#_c_466_n N_VGND_c_1358_n 0.00257529f $X=1.86 $Y=0.7 $X2=0
+ $Y2=0
cc_459 N_A_226_491#_c_468_n N_VGND_c_1358_n 0.0239155f $X=2.025 $Y=0.7 $X2=0
+ $Y2=0
cc_460 N_A_226_491#_c_469_n N_VGND_c_1358_n 0.00156301f $X=2.025 $Y=0.93 $X2=0
+ $Y2=0
cc_461 N_A_226_491#_c_466_n N_VGND_c_1362_n 0.00291965f $X=1.86 $Y=0.7 $X2=0
+ $Y2=0
cc_462 N_A_226_491#_c_467_n N_VGND_c_1362_n 0.0299351f $X=1.33 $Y=0.435 $X2=0
+ $Y2=0
cc_463 N_A_226_491#_c_465_n N_VGND_c_1364_n 0.0055654f $X=2.305 $Y=0.765 $X2=0
+ $Y2=0
cc_464 N_A_226_491#_c_468_n N_VGND_c_1364_n 5.08778e-19 $X=2.025 $Y=0.7 $X2=0
+ $Y2=0
cc_465 N_A_226_491#_c_469_n N_VGND_c_1364_n 7.42015e-19 $X=2.025 $Y=0.93 $X2=0
+ $Y2=0
cc_466 N_A_226_491#_M1014_s N_VGND_c_1370_n 0.00231914f $X=1.185 $Y=0.235 $X2=0
+ $Y2=0
cc_467 N_A_226_491#_c_465_n N_VGND_c_1370_n 0.011238f $X=2.305 $Y=0.765 $X2=0
+ $Y2=0
cc_468 N_A_226_491#_c_466_n N_VGND_c_1370_n 0.00512809f $X=1.86 $Y=0.7 $X2=0
+ $Y2=0
cc_469 N_A_226_491#_c_467_n N_VGND_c_1370_n 0.0180531f $X=1.33 $Y=0.435 $X2=0
+ $Y2=0
cc_470 N_A_226_491#_c_468_n N_VGND_c_1370_n 0.00257211f $X=2.025 $Y=0.7 $X2=0
+ $Y2=0
cc_471 N_A_226_491#_c_469_n N_VGND_c_1370_n 8.89392e-19 $X=2.025 $Y=0.93 $X2=0
+ $Y2=0
cc_472 N_A_114_179#_M1020_g N_A_831_21#_M1001_g 0.0396504f $X=4.12 $Y=2.595
+ $X2=0 $Y2=0
cc_473 N_A_114_179#_c_585_n N_A_831_21#_c_709_n 0.040709f $X=3.995 $Y=1.8 $X2=0
+ $Y2=0
cc_474 N_A_114_179#_M1003_g N_A_662_47#_c_874_n 0.00917469f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_475 N_A_114_179#_c_585_n N_A_662_47#_c_887_n 0.00529447f $X=3.995 $Y=1.8
+ $X2=0 $Y2=0
cc_476 N_A_114_179#_M1020_g N_A_662_47#_c_887_n 0.00565927f $X=4.12 $Y=2.595
+ $X2=0 $Y2=0
cc_477 N_A_114_179#_M1020_g N_A_662_47#_c_888_n 0.00947597f $X=4.12 $Y=2.595
+ $X2=0 $Y2=0
cc_478 N_A_114_179#_M1003_g N_A_662_47#_c_876_n 0.00143852f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_479 N_A_114_179#_c_573_n N_A_662_47#_c_876_n 0.00532527f $X=3.685 $Y=1.65
+ $X2=0 $Y2=0
cc_480 N_A_114_179#_c_575_n N_A_662_47#_c_876_n 0.00153734f $X=3.42 $Y=1.31
+ $X2=0 $Y2=0
cc_481 N_A_114_179#_M1003_g N_A_662_47#_c_877_n 0.00146206f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_482 N_A_114_179#_c_585_n N_A_662_47#_c_877_n 0.00413688f $X=3.995 $Y=1.8
+ $X2=0 $Y2=0
cc_483 N_A_114_179#_M1020_g N_A_662_47#_c_877_n 0.00338606f $X=4.12 $Y=2.595
+ $X2=0 $Y2=0
cc_484 N_A_114_179#_c_575_n N_A_662_47#_c_877_n 0.00407058f $X=3.42 $Y=1.31
+ $X2=0 $Y2=0
cc_485 N_A_114_179#_c_576_n N_A_662_47#_c_877_n 0.0170135f $X=3.76 $Y=1.65 $X2=0
+ $Y2=0
cc_486 N_A_114_179#_c_588_n N_VPWR_c_1085_n 0.0305639f $X=0.71 $Y=2.56 $X2=0
+ $Y2=0
cc_487 N_A_114_179#_c_588_n N_VPWR_c_1088_n 0.0241106f $X=0.71 $Y=2.56 $X2=0
+ $Y2=0
cc_488 N_A_114_179#_M1020_g N_VPWR_c_1089_n 0.00596406f $X=4.12 $Y=2.595 $X2=0
+ $Y2=0
cc_489 N_A_114_179#_M1020_g N_VPWR_c_1083_n 0.00712107f $X=4.12 $Y=2.595 $X2=0
+ $Y2=0
cc_490 N_A_114_179#_c_588_n N_VPWR_c_1083_n 0.0031395f $X=0.71 $Y=2.56 $X2=0
+ $Y2=0
cc_491 N_A_114_179#_M1002_g N_A_476_47#_c_1172_n 0.0114201f $X=2.875 $Y=0.445
+ $X2=0 $Y2=0
cc_492 N_A_114_179#_c_570_n N_A_476_47#_c_1172_n 6.84032e-19 $X=3.16 $Y=1.31
+ $X2=0 $Y2=0
cc_493 N_A_114_179#_M1003_g N_A_476_47#_c_1172_n 0.00686676f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_494 N_A_114_179#_c_581_n N_A_476_47#_c_1172_n 0.0102852f $X=2.785 $Y=1.22
+ $X2=0 $Y2=0
cc_495 N_A_114_179#_c_582_n N_A_476_47#_c_1172_n 6.49923e-19 $X=2.785 $Y=1.22
+ $X2=0 $Y2=0
cc_496 N_A_114_179#_M1002_g N_A_476_47#_c_1173_n 0.00849585f $X=2.875 $Y=0.445
+ $X2=0 $Y2=0
cc_497 N_A_114_179#_c_570_n N_A_476_47#_c_1173_n 0.00314365f $X=3.16 $Y=1.31
+ $X2=0 $Y2=0
cc_498 N_A_114_179#_M1003_g N_A_476_47#_c_1173_n 0.0121858f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_499 N_A_114_179#_c_572_n N_A_476_47#_c_1173_n 0.00626951f $X=3.42 $Y=1.575
+ $X2=0 $Y2=0
cc_500 N_A_114_179#_c_575_n N_A_476_47#_c_1173_n 0.00599604f $X=3.42 $Y=1.31
+ $X2=0 $Y2=0
cc_501 N_A_114_179#_c_581_n N_A_476_47#_c_1173_n 0.0297899f $X=2.785 $Y=1.22
+ $X2=0 $Y2=0
cc_502 N_A_114_179#_M1002_g N_A_476_47#_c_1174_n 0.007068f $X=2.875 $Y=0.445
+ $X2=0 $Y2=0
cc_503 N_A_114_179#_c_578_n N_A_476_47#_c_1174_n 0.00853898f $X=2.62 $Y=1.37
+ $X2=0 $Y2=0
cc_504 N_A_114_179#_c_581_n N_A_476_47#_c_1174_n 0.00307339f $X=2.785 $Y=1.22
+ $X2=0 $Y2=0
cc_505 N_A_114_179#_c_582_n N_A_476_47#_c_1174_n 4.50311e-19 $X=2.785 $Y=1.22
+ $X2=0 $Y2=0
cc_506 N_A_114_179#_c_570_n N_A_476_47#_c_1175_n 6.0824e-19 $X=3.16 $Y=1.31
+ $X2=0 $Y2=0
cc_507 N_A_114_179#_c_574_n N_A_476_47#_c_1175_n 0.00121779f $X=3.495 $Y=1.65
+ $X2=0 $Y2=0
cc_508 N_A_114_179#_c_576_n N_A_476_47#_c_1175_n 6.61092e-19 $X=3.76 $Y=1.65
+ $X2=0 $Y2=0
cc_509 N_A_114_179#_c_581_n N_A_476_47#_c_1175_n 0.010718f $X=2.785 $Y=1.22
+ $X2=0 $Y2=0
cc_510 N_A_114_179#_c_582_n N_A_476_47#_c_1175_n 0.00130405f $X=2.785 $Y=1.22
+ $X2=0 $Y2=0
cc_511 N_A_114_179#_M1020_g N_KAPWR_c_1246_n 0.00956062f $X=4.12 $Y=2.595 $X2=0
+ $Y2=0
cc_512 N_A_114_179#_c_588_n N_KAPWR_c_1246_n 0.0368757f $X=0.71 $Y=2.56 $X2=0
+ $Y2=0
cc_513 N_A_114_179#_M1020_g N_KAPWR_c_1247_n 6.92853e-19 $X=4.12 $Y=2.595 $X2=0
+ $Y2=0
cc_514 N_A_114_179#_c_577_n N_VGND_c_1357_n 0.0155541f $X=0.71 $Y=1.105 $X2=0
+ $Y2=0
cc_515 N_A_114_179#_c_579_n N_VGND_c_1357_n 0.00286735f $X=0.665 $Y=1.37 $X2=0
+ $Y2=0
cc_516 N_A_114_179#_M1002_g N_VGND_c_1364_n 0.00404693f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_517 N_A_114_179#_M1003_g N_VGND_c_1364_n 0.00428641f $X=3.235 $Y=0.445 $X2=0
+ $Y2=0
cc_518 N_A_114_179#_M1002_g N_VGND_c_1370_n 0.00586992f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_519 N_A_114_179#_M1003_g N_VGND_c_1370_n 0.00663699f $X=3.235 $Y=0.445 $X2=0
+ $Y2=0
cc_520 N_A_831_21#_c_707_n N_GATE_M1026_g 6.51883e-19 $X=5.53 $Y=1.575 $X2=0
+ $Y2=0
cc_521 N_A_831_21#_c_707_n N_GATE_M1023_g 0.00342284f $X=5.53 $Y=1.575 $X2=0
+ $Y2=0
cc_522 N_A_831_21#_c_708_n N_GATE_M1023_g 8.05639e-19 $X=5.595 $Y=0.465 $X2=0
+ $Y2=0
cc_523 N_A_831_21#_c_707_n N_GATE_c_780_n 8.33715e-19 $X=5.53 $Y=1.575 $X2=0
+ $Y2=0
cc_524 N_A_831_21#_c_707_n N_GATE_c_781_n 0.0505069f $X=5.53 $Y=1.575 $X2=0
+ $Y2=0
cc_525 N_A_831_21#_M1009_g N_A_662_47#_M1016_g 0.0141741f $X=4.59 $Y=0.445 $X2=0
+ $Y2=0
cc_526 N_A_831_21#_c_705_n N_A_662_47#_M1016_g 0.0128372f $X=4.625 $Y=0.87 $X2=0
+ $Y2=0
cc_527 N_A_831_21#_c_707_n N_A_662_47#_M1016_g 8.27828e-19 $X=5.53 $Y=1.575
+ $X2=0 $Y2=0
cc_528 N_A_831_21#_c_708_n N_A_662_47#_M1016_g 0.00114317f $X=5.595 $Y=0.465
+ $X2=0 $Y2=0
cc_529 N_A_831_21#_c_707_n N_A_662_47#_M1005_g 0.0054859f $X=5.53 $Y=1.575 $X2=0
+ $Y2=0
cc_530 N_A_831_21#_c_708_n N_A_662_47#_M1005_g 0.00822864f $X=5.595 $Y=0.465
+ $X2=0 $Y2=0
cc_531 N_A_831_21#_c_707_n N_A_662_47#_M1021_g 0.0211913f $X=5.53 $Y=1.575 $X2=0
+ $Y2=0
cc_532 N_A_831_21#_c_709_n N_A_662_47#_M1021_g 0.00228899f $X=4.66 $Y=1.74 $X2=0
+ $Y2=0
cc_533 N_A_831_21#_M1007_g N_A_662_47#_c_874_n 0.00295602f $X=4.23 $Y=0.445
+ $X2=0 $Y2=0
cc_534 N_A_831_21#_c_701_n N_A_662_47#_c_875_n 0.00928871f $X=4.515 $Y=0.87
+ $X2=0 $Y2=0
cc_535 N_A_831_21#_c_702_n N_A_662_47#_c_875_n 0.006683f $X=4.305 $Y=0.87 $X2=0
+ $Y2=0
cc_536 N_A_831_21#_c_704_n N_A_662_47#_c_875_n 0.00689747f $X=4.66 $Y=1.575
+ $X2=0 $Y2=0
cc_537 N_A_831_21#_c_705_n N_A_662_47#_c_875_n 0.00785649f $X=4.625 $Y=0.87
+ $X2=0 $Y2=0
cc_538 N_A_831_21#_c_706_n N_A_662_47#_c_875_n 0.0105558f $X=5.445 $Y=1.74 $X2=0
+ $Y2=0
cc_539 N_A_831_21#_c_709_n N_A_662_47#_c_875_n 0.00299399f $X=4.66 $Y=1.74 $X2=0
+ $Y2=0
cc_540 N_A_831_21#_c_704_n N_A_662_47#_c_878_n 0.00107336f $X=4.66 $Y=1.575
+ $X2=0 $Y2=0
cc_541 N_A_831_21#_c_706_n N_A_662_47#_c_878_n 0.0137633f $X=5.445 $Y=1.74 $X2=0
+ $Y2=0
cc_542 N_A_831_21#_c_707_n N_A_662_47#_c_878_n 0.0235661f $X=5.53 $Y=1.575 $X2=0
+ $Y2=0
cc_543 N_A_831_21#_c_704_n N_A_662_47#_c_879_n 0.0128372f $X=4.66 $Y=1.575 $X2=0
+ $Y2=0
cc_544 N_A_831_21#_c_706_n N_A_662_47#_c_879_n 0.00799362f $X=5.445 $Y=1.74
+ $X2=0 $Y2=0
cc_545 N_A_831_21#_c_707_n N_A_662_47#_c_879_n 0.0186512f $X=5.53 $Y=1.575 $X2=0
+ $Y2=0
cc_546 N_A_831_21#_c_708_n N_A_662_47#_c_879_n 0.00542049f $X=5.595 $Y=0.465
+ $X2=0 $Y2=0
cc_547 N_A_831_21#_M1001_g N_VPWR_c_1089_n 0.00937723f $X=4.61 $Y=2.595 $X2=0
+ $Y2=0
cc_548 N_A_831_21#_M1001_g N_VPWR_c_1083_n 0.00909986f $X=4.61 $Y=2.595 $X2=0
+ $Y2=0
cc_549 N_A_831_21#_M1021_s N_KAPWR_c_1246_n 0.00328907f $X=5.305 $Y=1.675 $X2=0
+ $Y2=0
cc_550 N_A_831_21#_M1001_g N_KAPWR_c_1246_n 0.00728819f $X=4.61 $Y=2.595 $X2=0
+ $Y2=0
cc_551 N_A_831_21#_M1001_g N_KAPWR_c_1247_n 0.0160558f $X=4.61 $Y=2.595 $X2=0
+ $Y2=0
cc_552 N_A_831_21#_M1007_g N_VGND_c_1359_n 0.0033384f $X=4.23 $Y=0.445 $X2=0
+ $Y2=0
cc_553 N_A_831_21#_M1009_g N_VGND_c_1359_n 0.0133392f $X=4.59 $Y=0.445 $X2=0
+ $Y2=0
cc_554 N_A_831_21#_c_705_n N_VGND_c_1359_n 0.00202389f $X=4.625 $Y=0.87 $X2=0
+ $Y2=0
cc_555 N_A_831_21#_c_708_n N_VGND_c_1359_n 0.0140521f $X=5.595 $Y=0.465 $X2=0
+ $Y2=0
cc_556 N_A_831_21#_M1007_g N_VGND_c_1364_n 0.00585385f $X=4.23 $Y=0.445 $X2=0
+ $Y2=0
cc_557 N_A_831_21#_M1009_g N_VGND_c_1364_n 0.00486043f $X=4.59 $Y=0.445 $X2=0
+ $Y2=0
cc_558 N_A_831_21#_c_708_n N_VGND_c_1366_n 0.0206712f $X=5.595 $Y=0.465 $X2=0
+ $Y2=0
cc_559 N_A_831_21#_M1005_d N_VGND_c_1370_n 0.00232718f $X=5.455 $Y=0.235 $X2=0
+ $Y2=0
cc_560 N_A_831_21#_M1007_g N_VGND_c_1370_n 0.00625395f $X=4.23 $Y=0.445 $X2=0
+ $Y2=0
cc_561 N_A_831_21#_c_701_n N_VGND_c_1370_n 6.27631e-19 $X=4.515 $Y=0.87 $X2=0
+ $Y2=0
cc_562 N_A_831_21#_M1009_g N_VGND_c_1370_n 0.00441898f $X=4.59 $Y=0.445 $X2=0
+ $Y2=0
cc_563 N_A_831_21#_c_708_n N_VGND_c_1370_n 0.0125675f $X=5.595 $Y=0.465 $X2=0
+ $Y2=0
cc_564 N_GATE_M1023_g N_SLEEP_B_M1017_g 0.0311653f $X=6.37 $Y=0.445 $X2=0 $Y2=0
cc_565 N_GATE_c_781_n N_SLEEP_B_M1017_g 2.61225e-19 $X=6.245 $Y=1.01 $X2=0 $Y2=0
cc_566 N_GATE_c_777_n N_SLEEP_B_M1018_g 0.0123717f $X=6.262 $Y=1.333 $X2=0 $Y2=0
cc_567 N_GATE_M1026_g N_SLEEP_B_M1018_g 0.0149839f $X=6.31 $Y=1.995 $X2=0 $Y2=0
cc_568 N_GATE_c_781_n N_SLEEP_B_M1018_g 7.59447e-19 $X=6.245 $Y=1.01 $X2=0 $Y2=0
cc_569 N_GATE_c_780_n N_SLEEP_B_c_823_n 0.0311653f $X=6.245 $Y=1.01 $X2=0 $Y2=0
cc_570 N_GATE_c_777_n N_A_662_47#_M1021_g 0.0127467f $X=6.262 $Y=1.333 $X2=0
+ $Y2=0
cc_571 N_GATE_M1026_g N_A_662_47#_M1021_g 0.0273824f $X=6.31 $Y=1.995 $X2=0
+ $Y2=0
cc_572 N_GATE_M1026_g N_A_662_47#_c_881_n 0.00555199f $X=6.31 $Y=1.995 $X2=0
+ $Y2=0
cc_573 N_GATE_c_780_n N_A_662_47#_c_879_n 0.0150099f $X=6.245 $Y=1.01 $X2=0
+ $Y2=0
cc_574 N_GATE_c_781_n N_A_662_47#_c_879_n 0.00819386f $X=6.245 $Y=1.01 $X2=0
+ $Y2=0
cc_575 N_GATE_c_781_n N_KAPWR_M1021_d 0.0047707f $X=6.245 $Y=1.01 $X2=0 $Y2=0
cc_576 N_GATE_M1026_g N_KAPWR_c_1243_n 0.00163523f $X=6.31 $Y=1.995 $X2=0 $Y2=0
cc_577 N_GATE_M1026_g N_KAPWR_c_1245_n 8.19255e-19 $X=6.31 $Y=1.995 $X2=0 $Y2=0
cc_578 N_GATE_M1023_g N_VGND_c_1366_n 0.00398374f $X=6.37 $Y=0.445 $X2=0 $Y2=0
cc_579 N_GATE_M1023_g N_VGND_c_1370_n 0.00690137f $X=6.37 $Y=0.445 $X2=0 $Y2=0
cc_580 N_GATE_c_781_n N_VGND_c_1370_n 0.0047984f $X=6.245 $Y=1.01 $X2=0 $Y2=0
cc_581 N_SLEEP_B_M1018_g N_A_662_47#_c_881_n 0.00555199f $X=6.88 $Y=1.995 $X2=0
+ $Y2=0
cc_582 N_SLEEP_B_M1018_g N_A_662_47#_c_869_n 0.00231926f $X=6.88 $Y=1.995 $X2=0
+ $Y2=0
cc_583 SLEEP_B N_A_662_47#_c_871_n 0.00510295f $X=7.355 $Y=0.84 $X2=0 $Y2=0
cc_584 N_SLEEP_B_c_823_n N_A_662_47#_c_871_n 0.00958177f $X=7.09 $Y=0.955 $X2=0
+ $Y2=0
cc_585 SLEEP_B N_A_662_47#_M1011_g 4.70621e-19 $X=7.355 $Y=0.84 $X2=0 $Y2=0
cc_586 N_SLEEP_B_c_823_n N_A_662_47#_M1011_g 0.00165661f $X=7.09 $Y=0.955 $X2=0
+ $Y2=0
cc_587 N_SLEEP_B_M1018_g N_A_662_47#_c_873_n 0.0204843f $X=6.88 $Y=1.995 $X2=0
+ $Y2=0
cc_588 SLEEP_B N_A_662_47#_c_873_n 0.0121688f $X=7.355 $Y=0.84 $X2=0 $Y2=0
cc_589 N_SLEEP_B_c_821_n N_A_1530_367#_c_1026_n 0.0037531f $X=7.09 $Y=0.775
+ $X2=0 $Y2=0
cc_590 SLEEP_B N_A_1530_367#_c_1026_n 0.0357363f $X=7.355 $Y=0.84 $X2=0 $Y2=0
cc_591 N_SLEEP_B_c_823_n N_A_1530_367#_c_1026_n 5.18064e-19 $X=7.09 $Y=0.955
+ $X2=0 $Y2=0
cc_592 SLEEP_B N_A_1530_367#_c_1031_n 0.00663793f $X=7.355 $Y=0.84 $X2=0 $Y2=0
cc_593 N_SLEEP_B_M1018_g N_KAPWR_c_1243_n 0.00347912f $X=6.88 $Y=1.995 $X2=0
+ $Y2=0
cc_594 N_SLEEP_B_M1018_g N_KAPWR_c_1244_n 0.00793003f $X=6.88 $Y=1.995 $X2=0
+ $Y2=0
cc_595 SLEEP_B N_KAPWR_c_1244_n 0.0225539f $X=7.355 $Y=0.84 $X2=0 $Y2=0
cc_596 N_SLEEP_B_c_823_n N_KAPWR_c_1244_n 0.00180625f $X=7.09 $Y=0.955 $X2=0
+ $Y2=0
cc_597 N_SLEEP_B_M1017_g N_VGND_c_1360_n 0.00258772f $X=6.73 $Y=0.445 $X2=0
+ $Y2=0
cc_598 N_SLEEP_B_c_821_n N_VGND_c_1360_n 0.0121757f $X=7.09 $Y=0.775 $X2=0 $Y2=0
cc_599 SLEEP_B N_VGND_c_1360_n 0.0255818f $X=7.355 $Y=0.84 $X2=0 $Y2=0
cc_600 N_SLEEP_B_c_823_n N_VGND_c_1360_n 0.00124832f $X=7.09 $Y=0.955 $X2=0
+ $Y2=0
cc_601 N_SLEEP_B_M1017_g N_VGND_c_1366_n 0.00404527f $X=6.73 $Y=0.445 $X2=0
+ $Y2=0
cc_602 N_SLEEP_B_c_821_n N_VGND_c_1366_n 0.00486043f $X=7.09 $Y=0.775 $X2=0
+ $Y2=0
cc_603 N_SLEEP_B_M1017_g N_VGND_c_1370_n 0.0053493f $X=6.73 $Y=0.445 $X2=0 $Y2=0
cc_604 N_SLEEP_B_c_821_n N_VGND_c_1370_n 0.00425456f $X=7.09 $Y=0.775 $X2=0
+ $Y2=0
cc_605 SLEEP_B N_VGND_c_1370_n 0.00897228f $X=7.355 $Y=0.84 $X2=0 $Y2=0
cc_606 N_A_662_47#_M1011_g N_A_1530_367#_M1010_g 0.0144833f $X=8.08 $Y=0.485
+ $X2=0 $Y2=0
cc_607 N_A_662_47#_M1000_g N_A_1530_367#_M1008_g 0.0242157f $X=8.01 $Y=2.155
+ $X2=0 $Y2=0
cc_608 N_A_662_47#_c_868_n N_A_1530_367#_c_1033_n 0.00720759f $X=7.5 $Y=2.785
+ $X2=0 $Y2=0
cc_609 N_A_662_47#_c_884_n N_A_1530_367#_c_1033_n 0.00575963f $X=7.935 $Y=2.86
+ $X2=0 $Y2=0
cc_610 N_A_662_47#_M1000_g N_A_1530_367#_c_1033_n 0.00866019f $X=8.01 $Y=2.155
+ $X2=0 $Y2=0
cc_611 N_A_662_47#_c_873_n N_A_1530_367#_c_1033_n 0.004149f $X=7.66 $Y=1.42
+ $X2=0 $Y2=0
cc_612 N_A_662_47#_c_869_n N_A_1530_367#_c_1026_n 0.00554149f $X=7.66 $Y=1.345
+ $X2=0 $Y2=0
cc_613 N_A_662_47#_c_870_n N_A_1530_367#_c_1026_n 0.0167322f $X=8.005 $Y=1 $X2=0
+ $Y2=0
cc_614 N_A_662_47#_M1011_g N_A_1530_367#_c_1026_n 0.00867117f $X=8.08 $Y=0.485
+ $X2=0 $Y2=0
cc_615 N_A_662_47#_c_870_n N_A_1530_367#_c_1027_n 0.00434987f $X=8.005 $Y=1
+ $X2=0 $Y2=0
cc_616 N_A_662_47#_M1000_g N_A_1530_367#_c_1027_n 0.00186809f $X=8.01 $Y=2.155
+ $X2=0 $Y2=0
cc_617 N_A_662_47#_c_869_n N_A_1530_367#_c_1028_n 0.00227652f $X=7.66 $Y=1.345
+ $X2=0 $Y2=0
cc_618 N_A_662_47#_c_868_n N_A_1530_367#_c_1029_n 0.00230726f $X=7.5 $Y=2.785
+ $X2=0 $Y2=0
cc_619 N_A_662_47#_M1000_g N_A_1530_367#_c_1029_n 0.00361693f $X=8.01 $Y=2.155
+ $X2=0 $Y2=0
cc_620 N_A_662_47#_c_871_n N_A_1530_367#_c_1030_n 0.00299933f $X=7.735 $Y=1
+ $X2=0 $Y2=0
cc_621 N_A_662_47#_M1011_g N_A_1530_367#_c_1030_n 0.00454219f $X=8.08 $Y=0.485
+ $X2=0 $Y2=0
cc_622 N_A_662_47#_c_868_n N_A_1530_367#_c_1031_n 0.00585849f $X=7.5 $Y=2.785
+ $X2=0 $Y2=0
cc_623 N_A_662_47#_c_869_n N_A_1530_367#_c_1031_n 0.00445375f $X=7.66 $Y=1.345
+ $X2=0 $Y2=0
cc_624 N_A_662_47#_M1000_g N_A_1530_367#_c_1031_n 0.00272336f $X=8.01 $Y=2.155
+ $X2=0 $Y2=0
cc_625 N_A_662_47#_M1000_g N_VPWR_c_1087_n 0.0176007f $X=8.01 $Y=2.155 $X2=0
+ $Y2=0
cc_626 N_A_662_47#_c_882_n N_VPWR_c_1089_n 0.0415852f $X=5.84 $Y=2.86 $X2=0
+ $Y2=0
cc_627 N_A_662_47#_M1024_d N_VPWR_c_1083_n 0.00162345f $X=3.6 $Y=2.455 $X2=0
+ $Y2=0
cc_628 N_A_662_47#_c_882_n N_VPWR_c_1083_n 0.0141595f $X=5.84 $Y=2.86 $X2=0
+ $Y2=0
cc_629 N_A_662_47#_c_874_n N_A_476_47#_c_1172_n 0.0139054f $X=3.625 $Y=0.465
+ $X2=0 $Y2=0
cc_630 N_A_662_47#_c_874_n N_A_476_47#_c_1173_n 0.0127603f $X=3.625 $Y=0.465
+ $X2=0 $Y2=0
cc_631 N_A_662_47#_c_876_n N_A_476_47#_c_1173_n 0.0137158f $X=3.66 $Y=0.93 $X2=0
+ $Y2=0
cc_632 N_A_662_47#_c_877_n N_A_476_47#_c_1173_n 0.0237243f $X=3.855 $Y=2.075
+ $X2=0 $Y2=0
cc_633 N_A_662_47#_c_877_n N_A_476_47#_c_1175_n 0.00695625f $X=3.855 $Y=2.075
+ $X2=0 $Y2=0
cc_634 N_A_662_47#_M1021_g N_KAPWR_c_1242_n 0.00674166f $X=5.715 $Y=2.175 $X2=0
+ $Y2=0
cc_635 N_A_662_47#_c_882_n N_KAPWR_c_1242_n 0.00604835f $X=5.84 $Y=2.86 $X2=0
+ $Y2=0
cc_636 N_A_662_47#_c_881_n N_KAPWR_c_1243_n 0.0222609f $X=7.425 $Y=2.86 $X2=0
+ $Y2=0
cc_637 N_A_662_47#_c_868_n N_KAPWR_c_1243_n 0.00737094f $X=7.5 $Y=2.785 $X2=0
+ $Y2=0
cc_638 N_A_662_47#_c_868_n N_KAPWR_c_1244_n 0.0113724f $X=7.5 $Y=2.785 $X2=0
+ $Y2=0
cc_639 N_A_662_47#_M1021_g N_KAPWR_c_1245_n 0.00968924f $X=5.715 $Y=2.175 $X2=0
+ $Y2=0
cc_640 N_A_662_47#_c_881_n N_KAPWR_c_1245_n 0.0116711f $X=7.425 $Y=2.86 $X2=0
+ $Y2=0
cc_641 N_A_662_47#_c_882_n N_KAPWR_c_1245_n 3.67318e-19 $X=5.84 $Y=2.86 $X2=0
+ $Y2=0
cc_642 N_A_662_47#_M1024_d N_KAPWR_c_1246_n 0.00368344f $X=3.6 $Y=2.455 $X2=0
+ $Y2=0
cc_643 N_A_662_47#_M1021_g N_KAPWR_c_1246_n 0.00367573f $X=5.715 $Y=2.175 $X2=0
+ $Y2=0
cc_644 N_A_662_47#_c_881_n N_KAPWR_c_1246_n 0.0294035f $X=7.425 $Y=2.86 $X2=0
+ $Y2=0
cc_645 N_A_662_47#_c_882_n N_KAPWR_c_1246_n 0.0027285f $X=5.84 $Y=2.86 $X2=0
+ $Y2=0
cc_646 N_A_662_47#_c_868_n N_KAPWR_c_1246_n 0.00984461f $X=7.5 $Y=2.785 $X2=0
+ $Y2=0
cc_647 N_A_662_47#_c_884_n N_KAPWR_c_1246_n 0.0105717f $X=7.935 $Y=2.86 $X2=0
+ $Y2=0
cc_648 N_A_662_47#_M1000_g N_KAPWR_c_1246_n 0.00825874f $X=8.01 $Y=2.155 $X2=0
+ $Y2=0
cc_649 N_A_662_47#_c_886_n N_KAPWR_c_1246_n 0.00219234f $X=7.5 $Y=2.86 $X2=0
+ $Y2=0
cc_650 N_A_662_47#_c_888_n N_KAPWR_c_1246_n 0.0251148f $X=3.855 $Y=2.405 $X2=0
+ $Y2=0
cc_651 N_A_662_47#_M1021_g N_KAPWR_c_1247_n 0.00571051f $X=5.715 $Y=2.175 $X2=0
+ $Y2=0
cc_652 N_A_662_47#_c_882_n N_KAPWR_c_1247_n 8.95819e-19 $X=5.84 $Y=2.86 $X2=0
+ $Y2=0
cc_653 N_A_662_47#_M1016_g N_VGND_c_1359_n 0.0127481f $X=5.02 $Y=0.445 $X2=0
+ $Y2=0
cc_654 N_A_662_47#_M1005_g N_VGND_c_1359_n 0.002375f $X=5.38 $Y=0.445 $X2=0
+ $Y2=0
cc_655 N_A_662_47#_c_875_n N_VGND_c_1359_n 0.0246782f $X=4.945 $Y=0.93 $X2=0
+ $Y2=0
cc_656 N_A_662_47#_c_878_n N_VGND_c_1359_n 0.00180432f $X=5.11 $Y=0.93 $X2=0
+ $Y2=0
cc_657 N_A_662_47#_M1011_g N_VGND_c_1360_n 0.00239065f $X=8.08 $Y=0.485 $X2=0
+ $Y2=0
cc_658 N_A_662_47#_M1011_g N_VGND_c_1361_n 0.00981658f $X=8.08 $Y=0.485 $X2=0
+ $Y2=0
cc_659 N_A_662_47#_c_874_n N_VGND_c_1364_n 0.0210258f $X=3.625 $Y=0.465 $X2=0
+ $Y2=0
cc_660 N_A_662_47#_M1016_g N_VGND_c_1366_n 0.00486043f $X=5.02 $Y=0.445 $X2=0
+ $Y2=0
cc_661 N_A_662_47#_M1005_g N_VGND_c_1366_n 0.0054895f $X=5.38 $Y=0.445 $X2=0
+ $Y2=0
cc_662 N_A_662_47#_M1011_g N_VGND_c_1368_n 0.00511358f $X=8.08 $Y=0.485 $X2=0
+ $Y2=0
cc_663 N_A_662_47#_M1003_d N_VGND_c_1370_n 0.00894382f $X=3.31 $Y=0.235 $X2=0
+ $Y2=0
cc_664 N_A_662_47#_M1016_g N_VGND_c_1370_n 0.00441689f $X=5.02 $Y=0.445 $X2=0
+ $Y2=0
cc_665 N_A_662_47#_M1005_g N_VGND_c_1370_n 0.0112803f $X=5.38 $Y=0.445 $X2=0
+ $Y2=0
cc_666 N_A_662_47#_M1011_g N_VGND_c_1370_n 0.0108382f $X=8.08 $Y=0.485 $X2=0
+ $Y2=0
cc_667 N_A_662_47#_c_874_n N_VGND_c_1370_n 0.0126421f $X=3.625 $Y=0.465 $X2=0
+ $Y2=0
cc_668 N_A_662_47#_c_875_n N_VGND_c_1370_n 0.0246964f $X=4.945 $Y=0.93 $X2=0
+ $Y2=0
cc_669 N_A_662_47#_c_876_n N_VGND_c_1370_n 0.00220932f $X=3.66 $Y=0.93 $X2=0
+ $Y2=0
cc_670 N_A_662_47#_c_878_n N_VGND_c_1370_n 0.00964872f $X=5.11 $Y=0.93 $X2=0
+ $Y2=0
cc_671 N_A_1530_367#_M1008_g N_VPWR_c_1087_n 0.0152899f $X=8.625 $Y=2.465 $X2=0
+ $Y2=0
cc_672 N_A_1530_367#_c_1033_n N_VPWR_c_1087_n 0.0440983f $X=7.795 $Y=1.98 $X2=0
+ $Y2=0
cc_673 N_A_1530_367#_c_1027_n N_VPWR_c_1087_n 0.0283177f $X=8.5 $Y=1.48 $X2=0
+ $Y2=0
cc_674 N_A_1530_367#_c_1028_n N_VPWR_c_1087_n 0.00393697f $X=8.5 $Y=1.48 $X2=0
+ $Y2=0
cc_675 N_A_1530_367#_M1008_g N_VPWR_c_1090_n 0.0054895f $X=8.625 $Y=2.465 $X2=0
+ $Y2=0
cc_676 N_A_1530_367#_M1008_g N_VPWR_c_1083_n 0.00743814f $X=8.625 $Y=2.465 $X2=0
+ $Y2=0
cc_677 N_A_1530_367#_c_1033_n N_KAPWR_c_1244_n 0.0380639f $X=7.795 $Y=1.98 $X2=0
+ $Y2=0
cc_678 N_A_1530_367#_c_1029_n N_KAPWR_c_1244_n 0.00631642f $X=7.795 $Y=1.815
+ $X2=0 $Y2=0
cc_679 N_A_1530_367#_M1008_g N_KAPWR_c_1246_n 0.00882038f $X=8.625 $Y=2.465
+ $X2=0 $Y2=0
cc_680 N_A_1530_367#_c_1033_n N_KAPWR_c_1246_n 0.0179056f $X=7.795 $Y=1.98 $X2=0
+ $Y2=0
cc_681 N_A_1530_367#_M1008_g N_Q_c_1339_n 0.00278259f $X=8.625 $Y=2.465 $X2=0
+ $Y2=0
cc_682 N_A_1530_367#_M1008_g N_Q_c_1340_n 0.013676f $X=8.625 $Y=2.465 $X2=0
+ $Y2=0
cc_683 N_A_1530_367#_M1010_g N_Q_c_1336_n 0.0167529f $X=8.625 $Y=0.695 $X2=0
+ $Y2=0
cc_684 N_A_1530_367#_c_1027_n N_Q_c_1336_n 0.0262113f $X=8.5 $Y=1.48 $X2=0 $Y2=0
cc_685 N_A_1530_367#_M1010_g Q 0.00283148f $X=8.625 $Y=0.695 $X2=0 $Y2=0
cc_686 N_A_1530_367#_M1010_g N_Q_c_1338_n 0.0113242f $X=8.625 $Y=0.695 $X2=0
+ $Y2=0
cc_687 N_A_1530_367#_c_1030_n N_VGND_c_1360_n 0.0235965f $X=7.865 $Y=0.43 $X2=0
+ $Y2=0
cc_688 N_A_1530_367#_M1010_g N_VGND_c_1361_n 0.00403375f $X=8.625 $Y=0.695 $X2=0
+ $Y2=0
cc_689 N_A_1530_367#_c_1027_n N_VGND_c_1361_n 0.0204044f $X=8.5 $Y=1.48 $X2=0
+ $Y2=0
cc_690 N_A_1530_367#_c_1028_n N_VGND_c_1361_n 0.00368575f $X=8.5 $Y=1.48 $X2=0
+ $Y2=0
cc_691 N_A_1530_367#_c_1030_n N_VGND_c_1361_n 0.0559102f $X=7.865 $Y=0.43 $X2=0
+ $Y2=0
cc_692 N_A_1530_367#_c_1030_n N_VGND_c_1368_n 0.0231227f $X=7.865 $Y=0.43 $X2=0
+ $Y2=0
cc_693 N_A_1530_367#_M1010_g N_VGND_c_1369_n 0.00511358f $X=8.625 $Y=0.695 $X2=0
+ $Y2=0
cc_694 N_A_1530_367#_M1010_g N_VGND_c_1370_n 0.0104744f $X=8.625 $Y=0.695 $X2=0
+ $Y2=0
cc_695 N_A_1530_367#_c_1030_n N_VGND_c_1370_n 0.0125851f $X=7.865 $Y=0.43 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_1083_n N_A_476_47#_M1012_d 0.00114246f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_697 N_VPWR_c_1083_n A_621_491# 0.0014076f $X=8.88 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_698 N_VPWR_c_1083_n A_849_419# 0.00142282f $X=8.88 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_699 N_VPWR_c_1083_n N_KAPWR_M1001_d 0.00119816f $X=8.88 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_700 N_VPWR_c_1089_n N_KAPWR_c_1242_n 0.0215072f $X=8.175 $Y=3.33 $X2=0 $Y2=0
cc_701 N_VPWR_c_1083_n N_KAPWR_c_1242_n 0.00295526f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_702 N_VPWR_c_1089_n N_KAPWR_c_1243_n 0.0233418f $X=8.175 $Y=3.33 $X2=0 $Y2=0
cc_703 N_VPWR_c_1083_n N_KAPWR_c_1243_n 0.00330232f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_704 N_VPWR_c_1089_n N_KAPWR_c_1245_n 0.0100325f $X=8.175 $Y=3.33 $X2=0 $Y2=0
cc_705 N_VPWR_c_1083_n N_KAPWR_c_1245_n 0.00201631f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_706 N_VPWR_M1004_s N_KAPWR_c_1246_n 0.00240507f $X=0.135 $Y=2.415 $X2=0 $Y2=0
cc_707 N_VPWR_M1022_d N_KAPWR_c_1246_n 0.0121562f $X=1.565 $Y=2.455 $X2=0 $Y2=0
cc_708 N_VPWR_M1000_d N_KAPWR_c_1246_n 0.00199666f $X=8.085 $Y=1.835 $X2=0 $Y2=0
cc_709 N_VPWR_c_1084_n N_KAPWR_c_1246_n 2.42196e-19 $X=0.24 $Y=3.245 $X2=0 $Y2=0
cc_710 N_VPWR_c_1085_n N_KAPWR_c_1246_n 0.0312731f $X=0.28 $Y=2.56 $X2=0 $Y2=0
cc_711 N_VPWR_c_1086_n N_KAPWR_c_1246_n 0.017079f $X=1.775 $Y=2.945 $X2=0 $Y2=0
cc_712 N_VPWR_c_1087_n N_KAPWR_c_1246_n 0.0448539f $X=8.34 $Y=1.98 $X2=0 $Y2=0
cc_713 N_VPWR_c_1088_n N_KAPWR_c_1246_n 0.00309978f $X=1.61 $Y=3.33 $X2=0 $Y2=0
cc_714 N_VPWR_c_1089_n N_KAPWR_c_1246_n 0.0160618f $X=8.175 $Y=3.33 $X2=0 $Y2=0
cc_715 N_VPWR_c_1090_n N_KAPWR_c_1246_n 0.00133521f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_716 N_VPWR_c_1083_n N_KAPWR_c_1246_n 0.950197f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_717 N_VPWR_c_1089_n N_KAPWR_c_1247_n 0.0291833f $X=8.175 $Y=3.33 $X2=0 $Y2=0
cc_718 N_VPWR_c_1083_n N_KAPWR_c_1247_n 0.00414336f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_719 N_VPWR_c_1083_n N_Q_M1008_d 0.00119401f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_720 N_VPWR_c_1087_n N_Q_c_1339_n 0.0515713f $X=8.34 $Y=1.98 $X2=0 $Y2=0
cc_721 N_VPWR_c_1090_n N_Q_c_1340_n 0.0210192f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_722 N_VPWR_c_1083_n N_Q_c_1340_n 0.00303861f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_723 N_A_476_47#_c_1176_n N_KAPWR_c_1246_n 0.0236122f $X=2.815 $Y=2.61 $X2=0
+ $Y2=0
cc_724 N_A_476_47#_c_1174_n N_VGND_c_1358_n 0.01277f $X=2.525 $Y=0.465 $X2=0
+ $Y2=0
cc_725 N_A_476_47#_c_1172_n N_VGND_c_1364_n 0.0125713f $X=3.12 $Y=0.59 $X2=0
+ $Y2=0
cc_726 N_A_476_47#_c_1174_n N_VGND_c_1364_n 0.0203872f $X=2.525 $Y=0.465 $X2=0
+ $Y2=0
cc_727 N_A_476_47#_M1025_d N_VGND_c_1370_n 0.00359114f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_728 N_A_476_47#_c_1172_n N_VGND_c_1370_n 0.0178392f $X=3.12 $Y=0.59 $X2=0
+ $Y2=0
cc_729 N_A_476_47#_c_1174_n N_VGND_c_1370_n 0.0125101f $X=2.525 $Y=0.465 $X2=0
+ $Y2=0
cc_730 N_A_476_47#_c_1172_n A_590_47# 0.00141055f $X=3.12 $Y=0.59 $X2=-0.19
+ $Y2=-0.245
cc_731 A_621_491# N_KAPWR_c_1246_n 0.001781f $X=3.105 $Y=2.455 $X2=3.03 $Y2=1.79
cc_732 A_849_419# N_KAPWR_c_1246_n 0.00180861f $X=4.245 $Y=2.095 $X2=3.03
+ $Y2=1.79
cc_733 N_KAPWR_c_1246_n N_Q_c_1340_n 0.0391576f $X=5.04 $Y=2.82 $X2=0 $Y2=0
cc_734 N_Q_c_1338_n N_VGND_c_1361_n 0.0329605f $X=8.84 $Y=0.42 $X2=0 $Y2=0
cc_735 N_Q_c_1338_n N_VGND_c_1369_n 0.0234289f $X=8.84 $Y=0.42 $X2=0 $Y2=0
cc_736 N_Q_c_1338_n N_VGND_c_1370_n 0.0126421f $X=8.84 $Y=0.42 $X2=0 $Y2=0
cc_737 N_VGND_c_1370_n A_590_47# 0.00207295f $X=8.88 $Y=0 $X2=-0.19 $Y2=-0.245
cc_738 N_VGND_c_1370_n A_783_47# 0.00353984f $X=8.88 $Y=0 $X2=-0.19 $Y2=-0.245
cc_739 N_VGND_c_1370_n A_861_47# 0.00309736f $X=8.88 $Y=0 $X2=-0.19 $Y2=-0.245
cc_740 N_VGND_c_1370_n A_1019_47# 0.00396516f $X=8.88 $Y=0 $X2=-0.19 $Y2=-0.245
cc_741 N_VGND_c_1370_n A_1289_47# 0.00207252f $X=8.88 $Y=0 $X2=-0.19 $Y2=-0.245
cc_742 N_VGND_c_1370_n A_1361_47# 0.00816993f $X=8.88 $Y=0 $X2=-0.19 $Y2=-0.245
