* File: sky130_fd_sc_lp__clkinv_2.spice
* Created: Wed Sep  2 09:40:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkinv_2.pex.spice"
.subckt sky130_fd_sc_lp__clkinv_2  VNB VPB A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1001_d N_A_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX5_noxref VNB VPB NWDIODE A=4.2895 P=8.33
*
.include "sky130_fd_sc_lp__clkinv_2.pxi.spice"
*
.ends
*
*
