* File: sky130_fd_sc_lp__o2111a_m.pxi.spice
* Created: Fri Aug 28 11:00:30 2020
* 
x_PM_SKY130_FD_SC_LP__O2111A_M%A_80_21# N_A_80_21#_M1000_s N_A_80_21#_M1011_d
+ N_A_80_21#_M1010_d N_A_80_21#_M1004_g N_A_80_21#_c_90_n N_A_80_21#_M1001_g
+ N_A_80_21#_c_92_n N_A_80_21#_c_93_n N_A_80_21#_c_94_n N_A_80_21#_c_95_n
+ N_A_80_21#_c_96_n N_A_80_21#_c_101_n N_A_80_21#_c_102_n N_A_80_21#_c_97_n
+ N_A_80_21#_c_103_n N_A_80_21#_c_104_n N_A_80_21#_c_105_n N_A_80_21#_c_106_n
+ N_A_80_21#_c_98_n PM_SKY130_FD_SC_LP__O2111A_M%A_80_21#
x_PM_SKY130_FD_SC_LP__O2111A_M%D1 N_D1_M1011_g N_D1_c_182_n N_D1_c_183_n
+ N_D1_c_184_n N_D1_M1000_g N_D1_c_185_n N_D1_c_186_n N_D1_c_191_n D1 D1 D1
+ N_D1_c_188_n PM_SKY130_FD_SC_LP__O2111A_M%D1
x_PM_SKY130_FD_SC_LP__O2111A_M%C1 N_C1_M1008_g N_C1_M1007_g N_C1_c_238_n
+ N_C1_c_242_n C1 C1 C1 C1 N_C1_c_240_n PM_SKY130_FD_SC_LP__O2111A_M%C1
x_PM_SKY130_FD_SC_LP__O2111A_M%B1 N_B1_c_288_n N_B1_M1010_g N_B1_M1009_g
+ N_B1_c_290_n B1 B1 B1 B1 N_B1_c_287_n PM_SKY130_FD_SC_LP__O2111A_M%B1
x_PM_SKY130_FD_SC_LP__O2111A_M%A2 N_A2_M1003_g N_A2_M1002_g N_A2_c_333_n
+ N_A2_c_338_n A2 A2 A2 N_A2_c_335_n PM_SKY130_FD_SC_LP__O2111A_M%A2
x_PM_SKY130_FD_SC_LP__O2111A_M%A1 N_A1_M1005_g N_A1_M1006_g N_A1_c_383_n
+ N_A1_c_378_n N_A1_c_379_n A1 A1 A1 A1 N_A1_c_381_n
+ PM_SKY130_FD_SC_LP__O2111A_M%A1
x_PM_SKY130_FD_SC_LP__O2111A_M%X N_X_M1004_s N_X_M1001_s N_X_c_411_n X X X X X X
+ X N_X_c_412_n N_X_c_410_n X PM_SKY130_FD_SC_LP__O2111A_M%X
x_PM_SKY130_FD_SC_LP__O2111A_M%VPWR N_VPWR_M1001_d N_VPWR_M1008_d N_VPWR_M1005_d
+ N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_434_n
+ N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n VPWR
+ N_VPWR_c_439_n N_VPWR_c_429_n PM_SKY130_FD_SC_LP__O2111A_M%VPWR
x_PM_SKY130_FD_SC_LP__O2111A_M%VGND N_VGND_M1004_d N_VGND_M1002_d N_VGND_c_486_n
+ N_VGND_c_487_n N_VGND_c_488_n N_VGND_c_489_n VGND N_VGND_c_490_n
+ N_VGND_c_491_n N_VGND_c_492_n N_VGND_c_493_n PM_SKY130_FD_SC_LP__O2111A_M%VGND
x_PM_SKY130_FD_SC_LP__O2111A_M%A_492_47# N_A_492_47#_M1009_d N_A_492_47#_M1006_d
+ N_A_492_47#_c_541_n N_A_492_47#_c_542_n N_A_492_47#_c_543_n
+ N_A_492_47#_c_544_n PM_SKY130_FD_SC_LP__O2111A_M%A_492_47#
cc_1 VNB N_A_80_21#_c_90_n 0.0242191f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.238
cc_2 VNB N_A_80_21#_M1001_g 0.0133235f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.885
cc_3 VNB N_A_80_21#_c_92_n 0.0269457f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.435
cc_4 VNB N_A_80_21#_c_93_n 0.00206039f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_5 VNB N_A_80_21#_c_94_n 0.0236159f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_6 VNB N_A_80_21#_c_95_n 0.0147104f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=0.81
cc_7 VNB N_A_80_21#_c_96_n 0.00165376f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.81
cc_8 VNB N_A_80_21#_c_97_n 0.00169333f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=0.51
cc_9 VNB N_A_80_21#_c_98_n 0.0231791f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=0.765
cc_10 VNB N_D1_c_182_n 0.0288562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_D1_c_183_n 0.00948712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_D1_c_184_n 0.0190876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D1_c_185_n 0.0190778f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=0.962
cc_14 VNB N_D1_c_186_n 0.0190547f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.238
cc_15 VNB D1 0.00118305f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.885
cc_16 VNB N_D1_c_188_n 0.0164179f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_17 VNB N_C1_M1007_g 0.0351152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C1_c_238_n 0.0359442f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_19 VNB C1 0.00584594f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.885
cc_20 VNB N_C1_c_240_n 0.0257084f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=0.81
cc_21 VNB N_B1_M1009_g 0.0527027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB B1 0.00682271f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_23 VNB N_B1_c_287_n 0.0134898f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.435
cc_24 VNB N_A2_M1002_g 0.0397982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A2_c_333_n 0.0181584f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_26 VNB A2 0.00540242f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=0.962
cc_27 VNB N_A2_c_335_n 0.0158878f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.895
cc_28 VNB N_A1_M1006_g 0.0227014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A1_c_378_n 0.0226623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_c_379_n 0.045551f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.435
cc_31 VNB A1 0.0233272f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_32 VNB N_A1_c_381_n 0.00973022f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=0.51
cc_33 VNB N_X_c_410_n 0.0492017f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.52
cc_34 VNB N_VPWR_c_429_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_486_n 0.00495479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_487_n 0.00494119f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=0.962
cc_37 VNB N_VGND_c_488_n 0.0625758f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.885
cc_38 VNB N_VGND_c_489_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.885
cc_39 VNB N_VGND_c_490_n 0.0186951f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.895
cc_40 VNB N_VGND_c_491_n 0.0221109f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=0.51
cc_41 VNB N_VGND_c_492_n 0.219847f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=0.51
cc_42 VNB N_VGND_c_493_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.82
cc_43 VNB N_A_492_47#_c_541_n 0.00131266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_492_47#_c_542_n 0.0193833f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_45 VNB N_A_492_47#_c_543_n 0.0050734f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_46 VNB N_A_492_47#_c_544_n 0.00300716f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.435
cc_47 VPB N_A_80_21#_M1001_g 0.0777058f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.885
cc_48 VPB N_A_80_21#_c_93_n 0.00729566f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.93
cc_49 VPB N_A_80_21#_c_101_n 0.0127956f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.52
cc_50 VPB N_A_80_21#_c_102_n 0.00250302f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.52
cc_51 VPB N_A_80_21#_c_103_n 0.00126234f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.82
cc_52 VPB N_A_80_21#_c_104_n 0.027312f $X=-0.19 $Y=1.655 $X2=2.425 $Y2=2.52
cc_53 VPB N_A_80_21#_c_105_n 0.0014249f $X=-0.19 $Y=1.655 $X2=2.53 $Y2=2.82
cc_54 VPB N_A_80_21#_c_106_n 0.00743452f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.52
cc_55 VPB N_D1_M1011_g 0.0504312f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.675
cc_56 VPB N_D1_c_186_n 0.0040295f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.238
cc_57 VPB N_D1_c_191_n 0.0171604f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.435
cc_58 VPB D1 0.00445054f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.885
cc_59 VPB N_C1_M1008_g 0.0590213f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.675
cc_60 VPB N_C1_c_242_n 0.0169534f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.435
cc_61 VPB C1 0.0034188f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.885
cc_62 VPB N_B1_c_288_n 0.021f $X=-0.19 $Y=1.655 $X2=1.265 $Y2=2.675
cc_63 VPB N_B1_M1010_g 0.0385612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_B1_c_290_n 0.0201032f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_65 VPB B1 0.00643674f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_66 VPB N_B1_c_287_n 0.00512564f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.435
cc_67 VPB N_A2_M1003_g 0.0494773f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.675
cc_68 VPB N_A2_c_333_n 0.00383996f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_69 VPB N_A2_c_338_n 0.0180086f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_70 VPB A2 0.0117077f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=0.962
cc_71 VPB N_A1_M1005_g 0.0387916f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.675
cc_72 VPB N_A1_c_383_n 0.0737942f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.238
cc_73 VPB A1 0.0391302f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.93
cc_74 VPB N_A1_c_381_n 0.00918478f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=0.51
cc_75 VPB N_X_c_411_n 7.1609e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_X_c_412_n 0.0115598f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.81
cc_77 VPB N_X_c_410_n 0.0565832f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.52
cc_78 VPB N_VPWR_c_430_n 0.00437582f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_79 VPB N_VPWR_c_431_n 0.00288248f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.885
cc_80 VPB N_VPWR_c_432_n 0.0126648f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.895
cc_81 VPB N_VPWR_c_433_n 0.0243744f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.93
cc_82 VPB N_VPWR_c_434_n 0.00401177f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.93
cc_83 VPB N_VPWR_c_435_n 0.0157189f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.81
cc_84 VPB N_VPWR_c_436_n 0.00522083f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.52
cc_85 VPB N_VPWR_c_437_n 0.0318538f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=0.725
cc_86 VPB N_VPWR_c_438_n 0.00510247f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=0.51
cc_87 VPB N_VPWR_c_439_n 0.0134401f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_429_n 0.0536083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 N_A_80_21#_M1001_g N_D1_M1011_g 0.0388769f $X=0.72 $Y=2.885 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_93_n N_D1_M1011_g 0.00191704f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_101_n N_D1_M1011_g 0.0131819f $X=1.3 $Y=2.52 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_103_n N_D1_M1011_g 0.0017418f $X=1.405 $Y=2.82 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_93_n N_D1_c_183_n 0.00159788f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_94_n N_D1_c_183_n 0.00742662f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_95_n N_D1_c_183_n 0.0130241f $X=1.11 $Y=0.81 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_95_n N_D1_c_184_n 0.00146205f $X=1.11 $Y=0.81 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_97_n N_D1_c_184_n 0.0119675f $X=1.215 $Y=0.51 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_90_n N_D1_c_185_n 0.00742662f $X=0.597 $Y=1.238 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_92_n N_D1_c_186_n 0.0135117f $X=0.597 $Y=1.435 $X2=0 $Y2=0
cc_100 N_A_80_21#_M1001_g N_D1_c_191_n 0.0135117f $X=0.72 $Y=2.885 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_101_n N_D1_c_191_n 0.00285165f $X=1.3 $Y=2.52 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_106_n N_D1_c_191_n 0.00110061f $X=1.405 $Y=2.52 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_90_n D1 0.00201882f $X=0.597 $Y=1.238 $X2=0 $Y2=0
cc_104 N_A_80_21#_M1001_g D1 0.00159489f $X=0.72 $Y=2.885 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_93_n D1 0.0342995f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_95_n D1 0.0103338f $X=1.11 $Y=0.81 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_101_n D1 0.00959922f $X=1.3 $Y=2.52 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_90_n N_D1_c_188_n 0.0135117f $X=0.597 $Y=1.238 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_93_n N_D1_c_188_n 0.00217681f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_95_n N_D1_c_188_n 0.00352419f $X=1.11 $Y=0.81 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_103_n N_C1_M1008_g 0.0017418f $X=1.405 $Y=2.82 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_104_n N_C1_M1008_g 0.0152449f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_95_n N_C1_M1007_g 2.34157e-19 $X=1.11 $Y=0.81 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_104_n N_C1_c_242_n 0.00246819f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_95_n C1 0.00287981f $X=1.11 $Y=0.81 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_104_n C1 0.0100372f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_104_n N_B1_M1010_g 0.0148008f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_105_n N_B1_M1010_g 0.0017418f $X=2.53 $Y=2.82 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_104_n N_B1_c_290_n 0.00394173f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_104_n B1 0.0166467f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_104_n N_A2_M1003_g 0.00551383f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_105_n N_A2_M1003_g 0.0017418f $X=2.53 $Y=2.82 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_104_n A2 0.00473482f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_124 N_A_80_21#_M1001_g N_X_c_411_n 0.00280495f $X=0.72 $Y=2.885 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_102_n N_X_c_411_n 0.00732621f $X=0.715 $Y=2.52 $X2=0 $Y2=0
cc_126 N_A_80_21#_M1001_g N_X_c_410_n 0.0107964f $X=0.72 $Y=2.885 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_93_n N_X_c_410_n 0.110997f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_96_n N_X_c_410_n 0.0131664f $X=0.715 $Y=0.81 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_102_n N_X_c_410_n 0.013988f $X=0.715 $Y=2.52 $X2=0 $Y2=0
cc_130 N_A_80_21#_c_98_n N_X_c_410_n 0.022766f $X=0.597 $Y=0.765 $X2=0 $Y2=0
cc_131 N_A_80_21#_M1001_g N_VPWR_c_430_n 0.00283606f $X=0.72 $Y=2.885 $X2=0
+ $Y2=0
cc_132 N_A_80_21#_c_101_n N_VPWR_c_430_n 0.0156577f $X=1.3 $Y=2.52 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_104_n N_VPWR_c_431_n 0.0173089f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_134 N_A_80_21#_M1001_g N_VPWR_c_433_n 0.00427177f $X=0.72 $Y=2.885 $X2=0
+ $Y2=0
cc_135 N_A_80_21#_c_101_n N_VPWR_c_433_n 0.00189187f $X=1.3 $Y=2.52 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_102_n N_VPWR_c_433_n 6.55542e-19 $X=0.715 $Y=2.52 $X2=0
+ $Y2=0
cc_137 N_A_80_21#_c_101_n N_VPWR_c_435_n 0.00335753f $X=1.3 $Y=2.52 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_103_n N_VPWR_c_435_n 0.008231f $X=1.405 $Y=2.82 $X2=0 $Y2=0
cc_139 N_A_80_21#_c_104_n N_VPWR_c_435_n 0.00245444f $X=2.425 $Y=2.52 $X2=0
+ $Y2=0
cc_140 N_A_80_21#_c_104_n N_VPWR_c_437_n 0.00586637f $X=2.425 $Y=2.52 $X2=0
+ $Y2=0
cc_141 N_A_80_21#_c_105_n N_VPWR_c_437_n 0.008231f $X=2.53 $Y=2.82 $X2=0 $Y2=0
cc_142 N_A_80_21#_M1011_d N_VPWR_c_429_n 0.0026421f $X=1.265 $Y=2.675 $X2=0
+ $Y2=0
cc_143 N_A_80_21#_M1010_d N_VPWR_c_429_n 0.00373063f $X=2.39 $Y=2.675 $X2=0
+ $Y2=0
cc_144 N_A_80_21#_M1001_g N_VPWR_c_429_n 0.00720937f $X=0.72 $Y=2.885 $X2=0
+ $Y2=0
cc_145 N_A_80_21#_c_101_n N_VPWR_c_429_n 0.009565f $X=1.3 $Y=2.52 $X2=0 $Y2=0
cc_146 N_A_80_21#_c_102_n N_VPWR_c_429_n 0.00131868f $X=0.715 $Y=2.52 $X2=0
+ $Y2=0
cc_147 N_A_80_21#_c_103_n N_VPWR_c_429_n 0.00765087f $X=1.405 $Y=2.82 $X2=0
+ $Y2=0
cc_148 N_A_80_21#_c_104_n N_VPWR_c_429_n 0.0156374f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_149 N_A_80_21#_c_105_n N_VPWR_c_429_n 0.00765087f $X=2.53 $Y=2.82 $X2=0 $Y2=0
cc_150 N_A_80_21#_c_94_n N_VGND_c_486_n 0.00139795f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_151 N_A_80_21#_c_95_n N_VGND_c_486_n 0.00594593f $X=1.11 $Y=0.81 $X2=0 $Y2=0
cc_152 N_A_80_21#_c_96_n N_VGND_c_486_n 0.0099165f $X=0.715 $Y=0.81 $X2=0 $Y2=0
cc_153 N_A_80_21#_c_97_n N_VGND_c_486_n 0.00952885f $X=1.215 $Y=0.51 $X2=0 $Y2=0
cc_154 N_A_80_21#_c_98_n N_VGND_c_486_n 0.00460896f $X=0.597 $Y=0.765 $X2=0
+ $Y2=0
cc_155 N_A_80_21#_c_95_n N_VGND_c_488_n 0.00477439f $X=1.11 $Y=0.81 $X2=0 $Y2=0
cc_156 N_A_80_21#_c_97_n N_VGND_c_488_n 0.00908451f $X=1.215 $Y=0.51 $X2=0 $Y2=0
cc_157 N_A_80_21#_c_96_n N_VGND_c_490_n 6.60115e-19 $X=0.715 $Y=0.81 $X2=0 $Y2=0
cc_158 N_A_80_21#_c_98_n N_VGND_c_490_n 0.00580462f $X=0.597 $Y=0.765 $X2=0
+ $Y2=0
cc_159 N_A_80_21#_M1000_s N_VGND_c_492_n 0.00746268f $X=1.09 $Y=0.235 $X2=0
+ $Y2=0
cc_160 N_A_80_21#_c_95_n N_VGND_c_492_n 0.00873461f $X=1.11 $Y=0.81 $X2=0 $Y2=0
cc_161 N_A_80_21#_c_96_n N_VGND_c_492_n 0.00165007f $X=0.715 $Y=0.81 $X2=0 $Y2=0
cc_162 N_A_80_21#_c_97_n N_VGND_c_492_n 0.00765087f $X=1.215 $Y=0.51 $X2=0 $Y2=0
cc_163 N_A_80_21#_c_98_n N_VGND_c_492_n 0.0126384f $X=0.597 $Y=0.765 $X2=0 $Y2=0
cc_164 N_D1_M1011_g N_C1_M1008_g 0.0459454f $X=1.19 $Y=2.885 $X2=0 $Y2=0
cc_165 N_D1_c_191_n N_C1_M1008_g 0.011291f $X=1.17 $Y=1.88 $X2=0 $Y2=0
cc_166 D1 N_C1_M1008_g 0.00146687f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_167 N_D1_c_184_n N_C1_M1007_g 0.0528208f $X=1.665 $Y=0.765 $X2=0 $Y2=0
cc_168 N_D1_c_185_n N_C1_M1007_g 0.00261233f $X=1.17 $Y=1.21 $X2=0 $Y2=0
cc_169 N_D1_c_182_n N_C1_c_238_n 0.0113788f $X=1.59 $Y=0.84 $X2=0 $Y2=0
cc_170 N_D1_c_185_n N_C1_c_238_n 0.011291f $X=1.17 $Y=1.21 $X2=0 $Y2=0
cc_171 D1 N_C1_c_238_n 0.00224428f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_172 N_D1_c_186_n N_C1_c_242_n 0.011291f $X=1.17 $Y=1.715 $X2=0 $Y2=0
cc_173 N_D1_M1011_g C1 2.81375e-19 $X=1.19 $Y=2.885 $X2=0 $Y2=0
cc_174 N_D1_c_182_n C1 0.00862051f $X=1.59 $Y=0.84 $X2=0 $Y2=0
cc_175 N_D1_c_185_n C1 0.00780227f $X=1.17 $Y=1.21 $X2=0 $Y2=0
cc_176 D1 C1 0.0399423f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_177 N_D1_c_188_n N_C1_c_240_n 0.011291f $X=1.17 $Y=1.375 $X2=0 $Y2=0
cc_178 N_D1_M1011_g N_VPWR_c_430_n 0.00151816f $X=1.19 $Y=2.885 $X2=0 $Y2=0
cc_179 N_D1_M1011_g N_VPWR_c_431_n 7.42935e-19 $X=1.19 $Y=2.885 $X2=0 $Y2=0
cc_180 N_D1_M1011_g N_VPWR_c_435_n 0.00437852f $X=1.19 $Y=2.885 $X2=0 $Y2=0
cc_181 N_D1_M1011_g N_VPWR_c_429_n 0.00619633f $X=1.19 $Y=2.885 $X2=0 $Y2=0
cc_182 N_D1_c_183_n N_VGND_c_488_n 0.00456946f $X=1.335 $Y=0.84 $X2=0 $Y2=0
cc_183 N_D1_c_184_n N_VGND_c_488_n 0.00585385f $X=1.665 $Y=0.765 $X2=0 $Y2=0
cc_184 N_D1_c_183_n N_VGND_c_492_n 0.00582457f $X=1.335 $Y=0.84 $X2=0 $Y2=0
cc_185 N_D1_c_184_n N_VGND_c_492_n 0.00794076f $X=1.665 $Y=0.765 $X2=0 $Y2=0
cc_186 N_C1_M1008_g N_B1_c_288_n 0.0110593f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_187 N_C1_c_242_n N_B1_c_288_n 0.00876784f $X=1.71 $Y=1.825 $X2=0 $Y2=0
cc_188 C1 N_B1_c_288_n 0.00108539f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_189 N_C1_M1008_g N_B1_M1010_g 0.0184997f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_190 N_C1_M1007_g N_B1_M1009_g 0.0769794f $X=2.025 $Y=0.445 $X2=0 $Y2=0
cc_191 C1 N_B1_M1009_g 2.95357e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_192 N_C1_c_240_n N_B1_M1009_g 0.00547019f $X=1.71 $Y=1.32 $X2=0 $Y2=0
cc_193 N_C1_M1008_g B1 0.00269366f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_194 N_C1_M1007_g B1 0.00768042f $X=2.025 $Y=0.445 $X2=0 $Y2=0
cc_195 N_C1_c_238_n B1 0.00483066f $X=2.025 $Y=1.23 $X2=0 $Y2=0
cc_196 C1 B1 0.066594f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_197 N_C1_c_240_n B1 0.0039996f $X=1.71 $Y=1.32 $X2=0 $Y2=0
cc_198 N_C1_c_238_n N_B1_c_287_n 8.31396e-19 $X=2.025 $Y=1.23 $X2=0 $Y2=0
cc_199 C1 N_B1_c_287_n 3.09496e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_200 N_C1_c_240_n N_B1_c_287_n 0.00876784f $X=1.71 $Y=1.32 $X2=0 $Y2=0
cc_201 N_C1_M1008_g N_VPWR_c_431_n 0.00685182f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_202 N_C1_M1008_g N_VPWR_c_435_n 0.00422464f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_203 N_C1_M1008_g N_VPWR_c_429_n 0.00500951f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_204 N_C1_M1007_g N_VGND_c_488_n 0.00585385f $X=2.025 $Y=0.445 $X2=0 $Y2=0
cc_205 N_C1_M1007_g N_VGND_c_492_n 0.00993297f $X=2.025 $Y=0.445 $X2=0 $Y2=0
cc_206 C1 N_VGND_c_492_n 0.00669775f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_207 N_B1_M1010_g N_A2_M1003_g 0.0307692f $X=2.315 $Y=2.885 $X2=0 $Y2=0
cc_208 N_B1_c_290_n N_A2_M1003_g 0.0154041f $X=2.272 $Y=2.215 $X2=0 $Y2=0
cc_209 B1 N_A2_M1003_g 4.78281e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_210 N_B1_M1009_g N_A2_M1002_g 0.0338672f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_211 B1 N_A2_M1002_g 0.00158213f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_212 N_B1_c_287_n N_A2_c_333_n 0.0154041f $X=2.25 $Y=1.71 $X2=0 $Y2=0
cc_213 N_B1_c_288_n N_A2_c_338_n 0.0154041f $X=2.272 $Y=2.028 $X2=0 $Y2=0
cc_214 N_B1_M1009_g A2 0.00661768f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_215 B1 A2 0.0587842f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_216 N_B1_M1009_g N_A2_c_335_n 0.0154041f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_217 B1 N_A2_c_335_n 7.78597e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_218 N_B1_M1010_g N_VPWR_c_431_n 0.00638576f $X=2.315 $Y=2.885 $X2=0 $Y2=0
cc_219 N_B1_M1010_g N_VPWR_c_437_n 0.00437852f $X=2.315 $Y=2.885 $X2=0 $Y2=0
cc_220 N_B1_M1010_g N_VPWR_c_429_n 0.00685069f $X=2.315 $Y=2.885 $X2=0 $Y2=0
cc_221 N_B1_M1009_g N_VGND_c_488_n 0.00585385f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_222 N_B1_M1009_g N_VGND_c_492_n 0.0101282f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_223 B1 N_VGND_c_492_n 0.00980315f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_224 N_B1_M1009_g N_A_492_47#_c_541_n 0.001666f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_225 N_B1_M1009_g N_A_492_47#_c_543_n 0.0040947f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_226 B1 N_A_492_47#_c_543_n 0.00437109f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_227 N_A2_M1002_g N_A1_M1006_g 0.0244165f $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_228 N_A2_M1003_g N_A1_c_383_n 0.0749869f $X=2.745 $Y=2.885 $X2=0 $Y2=0
cc_229 N_A2_c_338_n N_A1_c_383_n 0.00920498f $X=2.835 $Y=1.88 $X2=0 $Y2=0
cc_230 A2 N_A1_c_383_n 0.00207181f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_231 N_A2_M1002_g N_A1_c_379_n 0.00879051f $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_232 A2 N_A1_c_379_n 0.0022152f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_233 N_A2_c_335_n N_A1_c_379_n 0.00920498f $X=2.835 $Y=1.375 $X2=0 $Y2=0
cc_234 N_A2_M1003_g A1 7.42563e-19 $X=2.745 $Y=2.885 $X2=0 $Y2=0
cc_235 A2 A1 0.0320878f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_236 N_A2_c_335_n A1 0.00239899f $X=2.835 $Y=1.375 $X2=0 $Y2=0
cc_237 N_A2_c_333_n N_A1_c_381_n 0.00920498f $X=2.835 $Y=1.715 $X2=0 $Y2=0
cc_238 N_A2_M1003_g N_VPWR_c_432_n 0.00207709f $X=2.745 $Y=2.885 $X2=0 $Y2=0
cc_239 N_A2_M1003_g N_VPWR_c_437_n 0.00585385f $X=2.745 $Y=2.885 $X2=0 $Y2=0
cc_240 N_A2_M1003_g N_VPWR_c_429_n 0.0108402f $X=2.745 $Y=2.885 $X2=0 $Y2=0
cc_241 N_A2_M1002_g N_VGND_c_487_n 0.00288714f $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A2_M1002_g N_VGND_c_488_n 0.00437852f $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_243 N_A2_M1002_g N_VGND_c_492_n 0.00604796f $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_244 N_A2_M1002_g N_A_492_47#_c_541_n 9.325e-19 $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_245 N_A2_M1002_g N_A_492_47#_c_542_n 0.0125212f $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_246 A2 N_A_492_47#_c_542_n 0.0101515f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_247 N_A2_c_335_n N_A_492_47#_c_542_n 0.00324177f $X=2.835 $Y=1.375 $X2=0
+ $Y2=0
cc_248 A2 N_A_492_47#_c_543_n 0.00876354f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_249 N_A2_c_335_n N_A_492_47#_c_543_n 2.46176e-19 $X=2.835 $Y=1.375 $X2=0
+ $Y2=0
cc_250 N_A1_M1005_g N_VPWR_c_432_n 0.0113246f $X=3.105 $Y=2.885 $X2=0 $Y2=0
cc_251 N_A1_c_383_n N_VPWR_c_432_n 0.00505397f $X=3.455 $Y=2.12 $X2=0 $Y2=0
cc_252 A1 N_VPWR_c_432_n 0.00537346f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_253 N_A1_M1005_g N_VPWR_c_437_n 0.00486043f $X=3.105 $Y=2.885 $X2=0 $Y2=0
cc_254 N_A1_M1005_g N_VPWR_c_429_n 0.00818711f $X=3.105 $Y=2.885 $X2=0 $Y2=0
cc_255 A1 N_VPWR_c_429_n 0.00850174f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_256 N_A1_M1006_g N_VGND_c_487_n 0.00288714f $X=3.245 $Y=0.445 $X2=0 $Y2=0
cc_257 N_A1_M1006_g N_VGND_c_491_n 0.00437852f $X=3.245 $Y=0.445 $X2=0 $Y2=0
cc_258 N_A1_M1006_g N_VGND_c_492_n 0.00712774f $X=3.245 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A1_M1006_g N_A_492_47#_c_542_n 0.00798445f $X=3.245 $Y=0.445 $X2=0
+ $Y2=0
cc_260 N_A1_c_378_n N_A_492_47#_c_542_n 0.0159076f $X=3.365 $Y=0.895 $X2=0 $Y2=0
cc_261 A1 N_A_492_47#_c_542_n 0.0109849f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_262 N_A1_M1006_g N_A_492_47#_c_544_n 0.0020107f $X=3.245 $Y=0.445 $X2=0 $Y2=0
cc_263 N_X_c_411_n N_VPWR_c_433_n 0.0118624f $X=0.505 $Y=2.89 $X2=0 $Y2=0
cc_264 N_X_c_412_n N_VPWR_c_433_n 0.00992309f $X=0.26 $Y=2.785 $X2=0 $Y2=0
cc_265 N_X_M1001_s N_VPWR_c_429_n 0.00221771f $X=0.38 $Y=2.675 $X2=0 $Y2=0
cc_266 N_X_c_411_n N_VPWR_c_429_n 0.0107681f $X=0.505 $Y=2.89 $X2=0 $Y2=0
cc_267 N_X_c_412_n N_VPWR_c_429_n 0.00781253f $X=0.26 $Y=2.785 $X2=0 $Y2=0
cc_268 N_X_c_410_n N_VGND_c_490_n 0.0130576f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_269 N_X_M1004_s N_VGND_c_492_n 0.00410163f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_270 N_X_c_410_n N_VGND_c_492_n 0.00804818f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_271 N_VPWR_c_429_n A_564_535# 0.00899413f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_272 N_VGND_c_492_n A_348_47# 0.00747298f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_273 N_VGND_c_492_n A_420_47# 0.00307853f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_274 N_VGND_c_492_n N_A_492_47#_M1009_d 0.00442034f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_275 N_VGND_c_492_n N_A_492_47#_M1006_d 0.00311677f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_488_n N_A_492_47#_c_541_n 0.00776392f $X=2.925 $Y=0 $X2=0 $Y2=0
cc_277 N_VGND_c_492_n N_A_492_47#_c_541_n 0.00690901f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_487_n N_A_492_47#_c_542_n 0.0139569f $X=3.03 $Y=0.38 $X2=0 $Y2=0
cc_279 N_VGND_c_488_n N_A_492_47#_c_542_n 0.00305343f $X=2.925 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_491_n N_A_492_47#_c_542_n 0.00305343f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_492_n N_A_492_47#_c_542_n 0.0109462f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_491_n N_A_492_47#_c_544_n 0.00865775f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_492_n N_A_492_47#_c_544_n 0.00765087f $X=3.6 $Y=0 $X2=0 $Y2=0
