# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a41o_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a41o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.890000 1.210000 4.700000 1.585000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.870000 1.185000 5.170000 1.515000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.365000 1.210000 6.085000 1.520000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.395000 1.210000 7.580000 1.575000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.765000 1.195000 3.720000 1.535000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.055000 1.780000 1.225000 ;
        RECT 0.100000 1.225000 0.420000 1.755000 ;
        RECT 0.100000 1.755000 1.780000 1.925000 ;
        RECT 0.695000 0.255000 0.885000 1.055000 ;
        RECT 0.695000 1.925000 0.885000 3.075000 ;
        RECT 1.555000 0.255000 1.780000 1.055000 ;
        RECT 1.555000 1.925000 1.780000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.195000  0.085000 0.525000 0.885000 ;
      RECT 0.195000  2.095000 0.525000 3.245000 ;
      RECT 0.590000  1.405000 2.595000 1.575000 ;
      RECT 1.055000  0.085000 1.385000 0.885000 ;
      RECT 1.055000  2.095000 1.385000 3.245000 ;
      RECT 1.950000  0.085000 2.210000 1.105000 ;
      RECT 1.950000  1.815000 2.235000 3.245000 ;
      RECT 2.380000  0.255000 2.605000 0.685000 ;
      RECT 2.380000  0.685000 3.985000 1.015000 ;
      RECT 2.380000  1.015000 2.595000 1.405000 ;
      RECT 2.405000  1.575000 2.595000 1.705000 ;
      RECT 2.405000  1.705000 3.195000 1.875000 ;
      RECT 2.435000  2.045000 2.695000 2.905000 ;
      RECT 2.435000  2.905000 3.555000 3.075000 ;
      RECT 2.775000  0.085000 3.105000 0.515000 ;
      RECT 2.865000  1.875000 3.195000 2.735000 ;
      RECT 3.295000  0.255000 4.425000 0.505000 ;
      RECT 3.365000  1.755000 7.110000 1.925000 ;
      RECT 3.365000  1.925000 3.555000 2.905000 ;
      RECT 3.725000  2.095000 4.055000 3.245000 ;
      RECT 4.155000  0.505000 4.425000 0.765000 ;
      RECT 4.155000  0.765000 5.345000 1.015000 ;
      RECT 4.225000  1.925000 4.415000 3.075000 ;
      RECT 4.595000  0.265000 6.235000 0.595000 ;
      RECT 4.605000  2.095000 4.935000 3.245000 ;
      RECT 5.110000  1.925000 5.320000 3.075000 ;
      RECT 5.490000  2.095000 5.820000 3.245000 ;
      RECT 5.535000  0.765000 6.655000 0.870000 ;
      RECT 5.535000  0.870000 7.585000 1.040000 ;
      RECT 5.990000  1.925000 6.180000 3.075000 ;
      RECT 6.350000  2.095000 6.680000 3.245000 ;
      RECT 6.405000  0.255000 6.655000 0.765000 ;
      RECT 6.825000  0.085000 7.155000 0.700000 ;
      RECT 6.850000  1.925000 7.110000 3.075000 ;
      RECT 7.325000  0.255000 7.585000 0.870000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__a41o_4
END LIBRARY
