* File: sky130_fd_sc_lp__clkinvlp_8.spice
* Created: Wed Sep  2 09:41:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkinvlp_8.pex.spice"
.subckt sky130_fd_sc_lp__clkinvlp_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_A_M1014_g A_268_67# VNB NSHORT L=0.15 W=0.55 AD=0.14575
+ AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.2
+ SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1001 A_268_67# N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.5 SB=75002.6
+ A=0.0825 P=1.4 MULT=1
MM1004 A_426_67# N_A_M1004_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75001 SB=75002.1
+ A=0.0825 P=1.4 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g A_426_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001.3
+ SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1013 N_VGND_M1003_d N_A_M1013_g A_110_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001.8
+ SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1007 A_110_67# N_A_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75002.1 SB=75001
+ A=0.0825 P=1.4 MULT=1
MM1009 A_584_67# N_A_M1009_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75002.6 SB=75000.5
+ A=0.0825 P=1.4 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g A_584_67# VNB NSHORT L=0.15 W=0.55 AD=0.14575
+ AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75002.9
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125004 A=0.25 P=2.5
+ MULT=1
MM1002 N_Y_M1000_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125003 A=0.25 P=2.5
+ MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VPWR_M1002_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125003 A=0.25 P=2.5
+ MULT=1
MM1006 N_Y_M1005_d N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VPWR_M1006_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1011 N_Y_M1008_d N_A_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1012 N_Y_M1012_d N_A_M1012_g N_VPWR_M1011_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1015 N_Y_M1012_d N_A_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125000 A=0.25 P=2.5
+ MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__clkinvlp_8.pxi.spice"
*
.ends
*
*
