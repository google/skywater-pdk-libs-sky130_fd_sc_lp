* File: sky130_fd_sc_lp__o21ba_m.pxi.spice
* Created: Wed Sep  2 10:17:11 2020
* 
x_PM_SKY130_FD_SC_LP__O21BA_M%A_88_41# N_A_88_41#_M1007_s N_A_88_41#_M1009_d
+ N_A_88_41#_M1004_g N_A_88_41#_M1000_g N_A_88_41#_c_75_n N_A_88_41#_c_76_n
+ N_A_88_41#_c_77_n N_A_88_41#_c_78_n N_A_88_41#_c_89_p
+ PM_SKY130_FD_SC_LP__O21BA_M%A_88_41#
x_PM_SKY130_FD_SC_LP__O21BA_M%B1_N N_B1_N_M1008_g N_B1_N_M1005_g B1_N B1_N
+ N_B1_N_c_135_n N_B1_N_c_136_n PM_SKY130_FD_SC_LP__O21BA_M%B1_N
x_PM_SKY130_FD_SC_LP__O21BA_M%A_256_79# N_A_256_79#_M1008_d N_A_256_79#_M1005_d
+ N_A_256_79#_M1009_g N_A_256_79#_c_171_n N_A_256_79#_M1007_g
+ N_A_256_79#_c_172_n N_A_256_79#_c_173_n N_A_256_79#_c_180_n
+ N_A_256_79#_c_181_n N_A_256_79#_c_174_n N_A_256_79#_c_175_n
+ N_A_256_79#_c_176_n N_A_256_79#_c_177_n N_A_256_79#_c_178_n
+ PM_SKY130_FD_SC_LP__O21BA_M%A_256_79#
x_PM_SKY130_FD_SC_LP__O21BA_M%A2 N_A2_c_229_n N_A2_M1003_g N_A2_M1002_g
+ N_A2_c_235_n A2 A2 A2 A2 N_A2_c_232_n PM_SKY130_FD_SC_LP__O21BA_M%A2
x_PM_SKY130_FD_SC_LP__O21BA_M%A1 N_A1_M1001_g N_A1_M1006_g N_A1_c_274_n A1 A1 A1
+ A1 N_A1_c_272_n PM_SKY130_FD_SC_LP__O21BA_M%A1
x_PM_SKY130_FD_SC_LP__O21BA_M%X N_X_M1004_s N_X_M1000_s N_X_c_301_n N_X_c_302_n
+ X X X X X PM_SKY130_FD_SC_LP__O21BA_M%X
x_PM_SKY130_FD_SC_LP__O21BA_M%VPWR N_VPWR_M1000_d N_VPWR_M1009_s N_VPWR_M1001_d
+ N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n
+ N_VPWR_c_327_n N_VPWR_c_328_n VPWR N_VPWR_c_329_n N_VPWR_c_330_n
+ N_VPWR_c_321_n N_VPWR_c_332_n PM_SKY130_FD_SC_LP__O21BA_M%VPWR
x_PM_SKY130_FD_SC_LP__O21BA_M%VGND N_VGND_M1004_d N_VGND_M1002_d N_VGND_c_366_n
+ N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n N_VGND_c_382_n N_VGND_c_370_n
+ N_VGND_c_371_n N_VGND_c_372_n VGND N_VGND_c_373_n N_VGND_c_374_n
+ PM_SKY130_FD_SC_LP__O21BA_M%VGND
x_PM_SKY130_FD_SC_LP__O21BA_M%A_500_49# N_A_500_49#_M1007_d N_A_500_49#_M1006_d
+ N_A_500_49#_c_418_n N_A_500_49#_c_419_n N_A_500_49#_c_420_n
+ N_A_500_49#_c_421_n PM_SKY130_FD_SC_LP__O21BA_M%A_500_49#
cc_1 VNB N_A_88_41#_M1004_g 0.0404733f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.025
cc_2 VNB N_A_88_41#_c_75_n 0.0435128f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.37
cc_3 VNB N_A_88_41#_c_76_n 0.00771554f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=2.715
cc_4 VNB N_A_88_41#_c_77_n 0.0223813f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=0.39
cc_5 VNB N_A_88_41#_c_78_n 0.00249342f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=0.39
cc_6 VNB B1_N 0.00482179f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.025
cc_7 VNB N_B1_N_c_135_n 0.0303713f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=0.37
cc_8 VNB N_B1_N_c_136_n 0.0192902f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.37
cc_9 VNB N_A_256_79#_M1009_g 0.0117502f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.025
cc_10 VNB N_A_256_79#_c_171_n 0.0202399f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.045
cc_11 VNB N_A_256_79#_c_172_n 0.0459597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_256_79#_c_173_n 0.0310748f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=0.39
cc_13 VNB N_A_256_79#_c_174_n 0.0103112f $X=-0.19 $Y=-0.245 $X2=2.37 $Y2=2.82
cc_14 VNB N_A_256_79#_c_175_n 0.0156931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_256_79#_c_176_n 0.00186468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_256_79#_c_177_n 0.0278181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_256_79#_c_178_n 0.0045176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_229_n 0.0194379f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=2.675
cc_19 VNB N_A2_M1002_g 0.0406092f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.025
cc_20 VNB A2 0.00239073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_c_232_n 0.0264546f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=0.39
cc_22 VNB N_A1_M1006_g 0.0747211f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.535
cc_23 VNB A1 0.0206584f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.37
cc_24 VNB N_A1_c_272_n 0.0112101f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=2.82
cc_25 VNB N_X_c_301_n 0.0110556f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.535
cc_26 VNB N_X_c_302_n 7.32923e-19 $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.025
cc_27 VNB X 0.0228128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_321_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_366_n 0.00834176f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.535
cc_30 VNB N_VGND_c_367_n 0.0241493f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.025
cc_31 VNB N_VGND_c_368_n 0.00901417f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.025
cc_32 VNB N_VGND_c_369_n 0.0116434f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.045
cc_33 VNB N_VGND_c_370_n 0.00527464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_371_n 0.0658105f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=0.39
cc_35 VNB N_VGND_c_372_n 0.00401211f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=0.39
cc_36 VNB N_VGND_c_373_n 0.020886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_374_n 0.225281f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.37
cc_38 VNB N_A_500_49#_c_418_n 0.00108772f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.025
cc_39 VNB N_A_500_49#_c_419_n 0.0231031f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.045
cc_40 VNB N_A_500_49#_c_420_n 0.0028134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_500_49#_c_421_n 0.00317049f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.37
cc_42 VPB N_A_88_41#_M1004_g 0.0268504f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.025
cc_43 VPB N_A_88_41#_c_76_n 0.00676648f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=2.715
cc_44 VPB N_B1_N_M1005_g 0.0256955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB B1_N 0.0102593f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.025
cc_46 VPB N_B1_N_c_135_n 0.00662171f $X=-0.19 $Y=1.655 $X2=2.045 $Y2=0.37
cc_47 VPB N_A_256_79#_M1009_g 0.0706919f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.025
cc_48 VPB N_A_256_79#_c_180_n 0.00226677f $X=-0.19 $Y=1.655 $X2=2.21 $Y2=0.39
cc_49 VPB N_A_256_79#_c_181_n 0.0128109f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=0.39
cc_50 VPB N_A_256_79#_c_178_n 0.00584576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A2_c_229_n 0.00114646f $X=-0.19 $Y=1.655 $X2=2.23 $Y2=2.675
cc_52 VPB N_A2_M1003_g 0.0496936f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A2_c_235_n 0.0272533f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.045
cc_54 VPB A2 0.00650861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A1_M1001_g 0.03845f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A1_c_274_n 0.0838485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB A1 0.0192497f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.37
cc_58 VPB N_A1_c_272_n 0.0107424f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=2.82
cc_59 VPB X 0.017561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB X 0.0412882f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.37
cc_61 VPB X 0.011459f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.535
cc_62 VPB N_VPWR_c_322_n 0.00495479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_323_n 0.00484226f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=0.495
cc_64 VPB N_VPWR_c_324_n 0.0126648f $X=-0.19 $Y=1.655 $X2=2.045 $Y2=0.39
cc_65 VPB N_VPWR_c_325_n 0.0273869f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=2.82
cc_66 VPB N_VPWR_c_326_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_327_n 0.0212602f $X=-0.19 $Y=1.655 $X2=2.37 $Y2=2.82
cc_68 VPB N_VPWR_c_328_n 0.00362723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_329_n 0.0274415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_330_n 0.0185316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_321_n 0.0834225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_332_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 N_A_88_41#_M1004_g N_B1_N_M1005_g 0.0176165f $X=0.68 $Y=1.025 $X2=0 $Y2=0
cc_74 N_A_88_41#_M1004_g B1_N 0.0189224f $X=0.68 $Y=1.025 $X2=0 $Y2=0
cc_75 N_A_88_41#_M1004_g N_B1_N_c_135_n 0.0215825f $X=0.68 $Y=1.025 $X2=0 $Y2=0
cc_76 N_A_88_41#_M1004_g N_B1_N_c_136_n 0.0196272f $X=0.68 $Y=1.025 $X2=0 $Y2=0
cc_77 N_A_88_41#_c_75_n N_B1_N_c_136_n 0.00982868f $X=0.605 $Y=0.37 $X2=0 $Y2=0
cc_78 N_A_88_41#_c_77_n N_B1_N_c_136_n 0.0155763f $X=2.045 $Y=0.39 $X2=0 $Y2=0
cc_79 N_A_88_41#_c_77_n N_A_256_79#_M1008_d 0.00259556f $X=2.045 $Y=0.39
+ $X2=-0.19 $Y2=-0.245
cc_80 N_A_88_41#_c_76_n N_A_256_79#_M1009_g 0.0347265f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_81 N_A_88_41#_c_89_p N_A_256_79#_M1009_g 0.00333127f $X=2.37 $Y=2.82 $X2=0
+ $Y2=0
cc_82 N_A_88_41#_c_76_n N_A_256_79#_c_171_n 0.00628966f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_83 N_A_88_41#_c_78_n N_A_256_79#_c_171_n 0.00302238f $X=2.29 $Y=0.39 $X2=0
+ $Y2=0
cc_84 N_A_88_41#_c_76_n N_A_256_79#_c_172_n 0.012183f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_85 N_A_88_41#_c_77_n N_A_256_79#_c_172_n 0.00458438f $X=2.045 $Y=0.39 $X2=0
+ $Y2=0
cc_86 N_A_88_41#_c_78_n N_A_256_79#_c_172_n 0.00657218f $X=2.29 $Y=0.39 $X2=0
+ $Y2=0
cc_87 N_A_88_41#_c_76_n N_A_256_79#_c_173_n 0.00534309f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_88 N_A_88_41#_c_89_p N_A_256_79#_c_181_n 0.00221737f $X=2.37 $Y=2.82 $X2=0
+ $Y2=0
cc_89 N_A_88_41#_M1004_g N_A_256_79#_c_174_n 3.6599e-19 $X=0.68 $Y=1.025 $X2=0
+ $Y2=0
cc_90 N_A_88_41#_c_76_n N_A_256_79#_c_174_n 0.00454617f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_91 N_A_88_41#_c_77_n N_A_256_79#_c_174_n 0.0231547f $X=2.045 $Y=0.39 $X2=0
+ $Y2=0
cc_92 N_A_88_41#_c_76_n N_A_256_79#_c_175_n 0.012149f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_93 N_A_88_41#_c_76_n N_A_256_79#_c_176_n 0.03221f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_94 N_A_88_41#_c_77_n N_A_256_79#_c_176_n 0.00736287f $X=2.045 $Y=0.39 $X2=0
+ $Y2=0
cc_95 N_A_88_41#_c_76_n N_A_256_79#_c_177_n 0.00825357f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_96 N_A_88_41#_c_76_n N_A_256_79#_c_178_n 0.0381826f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_97 N_A_88_41#_c_89_p N_A2_M1003_g 0.00495015f $X=2.37 $Y=2.82 $X2=0 $Y2=0
cc_98 N_A_88_41#_c_76_n N_A2_M1002_g 0.00526649f $X=2.29 $Y=2.715 $X2=0 $Y2=0
cc_99 N_A_88_41#_c_76_n A2 0.0888087f $X=2.29 $Y=2.715 $X2=0 $Y2=0
cc_100 N_A_88_41#_c_76_n N_A2_c_232_n 0.0130919f $X=2.29 $Y=2.715 $X2=0 $Y2=0
cc_101 N_A_88_41#_c_89_p N_A1_M1001_g 8.63638e-19 $X=2.37 $Y=2.82 $X2=0 $Y2=0
cc_102 N_A_88_41#_M1004_g N_X_c_302_n 0.00423838f $X=0.68 $Y=1.025 $X2=0 $Y2=0
cc_103 N_A_88_41#_M1004_g X 0.0186761f $X=0.68 $Y=1.025 $X2=0 $Y2=0
cc_104 N_A_88_41#_M1004_g X 0.00513084f $X=0.68 $Y=1.025 $X2=0 $Y2=0
cc_105 N_A_88_41#_M1004_g X 0.00491774f $X=0.68 $Y=1.025 $X2=0 $Y2=0
cc_106 N_A_88_41#_M1004_g N_VPWR_c_322_n 0.00231568f $X=0.68 $Y=1.025 $X2=0
+ $Y2=0
cc_107 N_A_88_41#_c_89_p N_VPWR_c_324_n 0.0026493f $X=2.37 $Y=2.82 $X2=0 $Y2=0
cc_108 N_A_88_41#_c_89_p N_VPWR_c_329_n 0.00909174f $X=2.37 $Y=2.82 $X2=0 $Y2=0
cc_109 N_A_88_41#_M1009_d N_VPWR_c_321_n 0.00246398f $X=2.23 $Y=2.675 $X2=0
+ $Y2=0
cc_110 N_A_88_41#_c_89_p N_VPWR_c_321_n 0.0110299f $X=2.37 $Y=2.82 $X2=0 $Y2=0
cc_111 N_A_88_41#_c_77_n N_VGND_M1004_d 0.00354661f $X=2.045 $Y=0.39 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_88_41#_M1004_g N_VGND_c_367_n 0.00281355f $X=0.68 $Y=1.025 $X2=0
+ $Y2=0
cc_113 N_A_88_41#_c_75_n N_VGND_c_367_n 0.00682244f $X=0.605 $Y=0.37 $X2=0 $Y2=0
cc_114 N_A_88_41#_c_77_n N_VGND_c_367_n 0.0128545f $X=2.045 $Y=0.39 $X2=0 $Y2=0
cc_115 N_A_88_41#_M1004_g N_VGND_c_368_n 0.0141611f $X=0.68 $Y=1.025 $X2=0 $Y2=0
cc_116 N_A_88_41#_c_75_n N_VGND_c_368_n 0.00440824f $X=0.605 $Y=0.37 $X2=0 $Y2=0
cc_117 N_A_88_41#_c_77_n N_VGND_c_368_n 0.0385433f $X=2.045 $Y=0.39 $X2=0 $Y2=0
cc_118 N_A_88_41#_M1004_g N_VGND_c_382_n 2.19257e-19 $X=0.68 $Y=1.025 $X2=0
+ $Y2=0
cc_119 N_A_88_41#_c_75_n N_VGND_c_371_n 0.00634371f $X=0.605 $Y=0.37 $X2=0 $Y2=0
cc_120 N_A_88_41#_c_77_n N_VGND_c_371_n 0.102145f $X=2.045 $Y=0.39 $X2=0 $Y2=0
cc_121 N_A_88_41#_M1007_s N_VGND_c_374_n 0.002136f $X=2.085 $Y=0.245 $X2=0 $Y2=0
cc_122 N_A_88_41#_c_75_n N_VGND_c_374_n 0.00909824f $X=0.605 $Y=0.37 $X2=0 $Y2=0
cc_123 N_A_88_41#_c_77_n N_VGND_c_374_n 0.0696775f $X=2.045 $Y=0.39 $X2=0 $Y2=0
cc_124 N_A_88_41#_c_76_n N_A_500_49#_c_418_n 0.0102683f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_125 N_A_88_41#_c_76_n N_A_500_49#_c_420_n 0.0131052f $X=2.29 $Y=2.715 $X2=0
+ $Y2=0
cc_126 N_B1_N_c_136_n N_A_256_79#_c_172_n 0.00604367f $X=1.13 $Y=1.345 $X2=0
+ $Y2=0
cc_127 N_B1_N_c_135_n N_A_256_79#_c_173_n 0.001985f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_128 B1_N N_A_256_79#_c_174_n 0.00353952f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_129 N_B1_N_c_135_n N_A_256_79#_c_174_n 0.00241355f $X=1.13 $Y=1.51 $X2=0
+ $Y2=0
cc_130 N_B1_N_c_136_n N_A_256_79#_c_174_n 0.0112552f $X=1.13 $Y=1.345 $X2=0
+ $Y2=0
cc_131 N_B1_N_M1005_g N_A_256_79#_c_178_n 0.00601781f $X=1.205 $Y=2.465 $X2=0
+ $Y2=0
cc_132 B1_N N_A_256_79#_c_178_n 0.0235061f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_133 N_B1_N_c_135_n N_A_256_79#_c_178_n 0.00159907f $X=1.13 $Y=1.51 $X2=0
+ $Y2=0
cc_134 N_B1_N_c_136_n N_X_c_302_n 2.45758e-19 $X=1.13 $Y=1.345 $X2=0 $Y2=0
cc_135 B1_N X 0.0163879f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_136 N_B1_N_M1005_g X 4.82427e-19 $X=1.205 $Y=2.465 $X2=0 $Y2=0
cc_137 N_B1_N_M1005_g N_VPWR_c_322_n 0.00460896f $X=1.205 $Y=2.465 $X2=0 $Y2=0
cc_138 B1_N N_VPWR_c_322_n 0.0100766f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_139 N_B1_N_c_135_n N_VPWR_c_322_n 7.32048e-19 $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_140 N_B1_N_M1005_g N_VPWR_c_323_n 0.0051578f $X=1.205 $Y=2.465 $X2=0 $Y2=0
cc_141 N_B1_N_M1005_g N_VPWR_c_327_n 0.00585385f $X=1.205 $Y=2.465 $X2=0 $Y2=0
cc_142 N_B1_N_M1005_g N_VPWR_c_321_n 0.0133979f $X=1.205 $Y=2.465 $X2=0 $Y2=0
cc_143 B1_N N_VGND_c_368_n 0.0046802f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_144 N_B1_N_c_136_n N_VGND_c_368_n 0.00182165f $X=1.13 $Y=1.345 $X2=0 $Y2=0
cc_145 B1_N N_VGND_c_382_n 0.0114286f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_146 N_B1_N_c_135_n N_VGND_c_382_n 0.00126544f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_147 N_B1_N_c_136_n N_VGND_c_382_n 0.00266144f $X=1.13 $Y=1.345 $X2=0 $Y2=0
cc_148 N_B1_N_c_136_n N_VGND_c_371_n 0.00387882f $X=1.13 $Y=1.345 $X2=0 $Y2=0
cc_149 N_B1_N_c_136_n N_VGND_c_374_n 0.00537853f $X=1.13 $Y=1.345 $X2=0 $Y2=0
cc_150 N_A_256_79#_c_173_n N_A2_c_229_n 0.0237889f $X=2.002 $Y=1.445 $X2=0 $Y2=0
cc_151 N_A_256_79#_c_171_n N_A2_M1002_g 0.0209081f $X=2.425 $Y=0.775 $X2=0 $Y2=0
cc_152 N_A_256_79#_c_177_n N_A2_M1002_g 0.00447202f $X=1.94 $Y=0.94 $X2=0 $Y2=0
cc_153 N_A_256_79#_M1009_g N_A2_c_235_n 0.0237889f $X=2.155 $Y=2.885 $X2=0 $Y2=0
cc_154 N_A_256_79#_c_177_n A2 0.00120809f $X=1.94 $Y=0.94 $X2=0 $Y2=0
cc_155 N_A_256_79#_c_177_n N_A2_c_232_n 0.0237889f $X=1.94 $Y=0.94 $X2=0 $Y2=0
cc_156 N_A_256_79#_c_174_n N_X_c_302_n 0.001836f $X=1.56 $Y=1.445 $X2=0 $Y2=0
cc_157 N_A_256_79#_M1009_g N_VPWR_c_323_n 0.00442088f $X=2.155 $Y=2.885 $X2=0
+ $Y2=0
cc_158 N_A_256_79#_c_181_n N_VPWR_c_323_n 0.0111816f $X=1.42 $Y=2.095 $X2=0
+ $Y2=0
cc_159 N_A_256_79#_c_181_n N_VPWR_c_327_n 0.0115814f $X=1.42 $Y=2.095 $X2=0
+ $Y2=0
cc_160 N_A_256_79#_M1009_g N_VPWR_c_329_n 0.00552362f $X=2.155 $Y=2.885 $X2=0
+ $Y2=0
cc_161 N_A_256_79#_M1005_d N_VPWR_c_321_n 0.0042376f $X=1.28 $Y=1.835 $X2=0
+ $Y2=0
cc_162 N_A_256_79#_M1009_g N_VPWR_c_321_n 0.011165f $X=2.155 $Y=2.885 $X2=0
+ $Y2=0
cc_163 N_A_256_79#_c_181_n N_VPWR_c_321_n 0.0110901f $X=1.42 $Y=2.095 $X2=0
+ $Y2=0
cc_164 N_A_256_79#_c_174_n N_VGND_c_368_n 0.0104554f $X=1.56 $Y=1.445 $X2=0
+ $Y2=0
cc_165 N_A_256_79#_c_174_n N_VGND_c_382_n 0.0189935f $X=1.56 $Y=1.445 $X2=0
+ $Y2=0
cc_166 N_A_256_79#_c_171_n N_VGND_c_371_n 0.00538845f $X=2.425 $Y=0.775 $X2=0
+ $Y2=0
cc_167 N_A_256_79#_c_171_n N_VGND_c_374_n 0.0112526f $X=2.425 $Y=0.775 $X2=0
+ $Y2=0
cc_168 N_A_256_79#_c_171_n N_A_500_49#_c_418_n 4.98848e-19 $X=2.425 $Y=0.775
+ $X2=0 $Y2=0
cc_169 N_A_256_79#_c_171_n N_A_500_49#_c_420_n 0.00164017f $X=2.425 $Y=0.775
+ $X2=0 $Y2=0
cc_170 N_A2_M1002_g N_A1_M1006_g 0.0526964f $X=2.855 $Y=0.455 $X2=0 $Y2=0
cc_171 A2 N_A1_M1006_g 3.1139e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_172 N_A2_M1003_g N_A1_c_274_n 0.0731335f $X=2.585 $Y=2.885 $X2=0 $Y2=0
cc_173 N_A2_c_235_n N_A1_c_274_n 0.0118515f $X=2.72 $Y=1.88 $X2=0 $Y2=0
cc_174 A2 N_A1_c_274_n 0.00344018f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A2_M1003_g A1 9.98415e-19 $X=2.585 $Y=2.885 $X2=0 $Y2=0
cc_176 A2 A1 0.0711054f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A2_c_232_n A1 0.00616034f $X=2.675 $Y=1.375 $X2=0 $Y2=0
cc_178 N_A2_c_229_n N_A1_c_272_n 0.00740875f $X=2.72 $Y=1.67 $X2=0 $Y2=0
cc_179 A2 N_A1_c_272_n 2.29219e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A2_M1003_g N_VPWR_c_324_n 0.0022041f $X=2.585 $Y=2.885 $X2=0 $Y2=0
cc_181 N_A2_M1003_g N_VPWR_c_329_n 0.00552362f $X=2.585 $Y=2.885 $X2=0 $Y2=0
cc_182 N_A2_M1003_g N_VPWR_c_321_n 0.00684977f $X=2.585 $Y=2.885 $X2=0 $Y2=0
cc_183 A2 N_VPWR_c_321_n 0.00720306f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A2_M1002_g N_VGND_c_370_n 0.00279829f $X=2.855 $Y=0.455 $X2=0 $Y2=0
cc_185 N_A2_M1002_g N_VGND_c_371_n 0.00430555f $X=2.855 $Y=0.455 $X2=0 $Y2=0
cc_186 N_A2_M1002_g N_VGND_c_374_n 0.00602213f $X=2.855 $Y=0.455 $X2=0 $Y2=0
cc_187 N_A2_M1002_g N_A_500_49#_c_418_n 9.325e-19 $X=2.855 $Y=0.455 $X2=0 $Y2=0
cc_188 N_A2_M1002_g N_A_500_49#_c_419_n 0.0163196f $X=2.855 $Y=0.455 $X2=0 $Y2=0
cc_189 A2 N_A_500_49#_c_419_n 6.95622e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A2_c_232_n N_A_500_49#_c_419_n 8.30955e-19 $X=2.675 $Y=1.375 $X2=0
+ $Y2=0
cc_191 A2 N_A_500_49#_c_420_n 0.0106851f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A2_c_232_n N_A_500_49#_c_420_n 0.00133524f $X=2.675 $Y=1.375 $X2=0
+ $Y2=0
cc_193 N_A1_M1001_g N_VPWR_c_324_n 0.0112663f $X=2.945 $Y=2.885 $X2=0 $Y2=0
cc_194 N_A1_c_274_n N_VPWR_c_324_n 0.0012529f $X=3.335 $Y=2.12 $X2=0 $Y2=0
cc_195 A1 N_VPWR_c_324_n 0.0125401f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A1_M1001_g N_VPWR_c_329_n 0.00486043f $X=2.945 $Y=2.885 $X2=0 $Y2=0
cc_197 N_A1_M1001_g N_VPWR_c_321_n 0.00818711f $X=2.945 $Y=2.885 $X2=0 $Y2=0
cc_198 A1 N_VPWR_c_321_n 0.00531513f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_199 N_A1_M1006_g N_VGND_c_370_n 0.00279829f $X=3.285 $Y=0.455 $X2=0 $Y2=0
cc_200 N_A1_M1006_g N_VGND_c_373_n 0.00430555f $X=3.285 $Y=0.455 $X2=0 $Y2=0
cc_201 N_A1_M1006_g N_VGND_c_374_n 0.00699676f $X=3.285 $Y=0.455 $X2=0 $Y2=0
cc_202 N_A1_M1006_g N_A_500_49#_c_419_n 0.0142025f $X=3.285 $Y=0.455 $X2=0 $Y2=0
cc_203 A1 N_A_500_49#_c_419_n 0.0203402f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_204 N_A1_c_272_n N_A_500_49#_c_419_n 0.00251671f $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A1_M1006_g N_A_500_49#_c_421_n 0.0020107f $X=3.285 $Y=0.455 $X2=0 $Y2=0
cc_206 X N_VPWR_c_322_n 0.044752f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_207 X N_VPWR_c_325_n 0.0141816f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_208 X N_VPWR_c_321_n 0.0161584f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_209 N_X_c_301_n N_VGND_c_368_n 0.00523553f $X=0.325 $Y=1.09 $X2=0 $Y2=0
cc_210 N_X_c_302_n N_VGND_c_368_n 0.0197332f $X=0.465 $Y=1.09 $X2=0 $Y2=0
cc_211 N_X_c_301_n N_VGND_c_369_n 0.00944503f $X=0.325 $Y=1.09 $X2=0 $Y2=0
cc_212 N_VPWR_c_321_n A_532_535# 0.00620535f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_213 N_VGND_c_374_n N_A_500_49#_M1007_d 0.00443725f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_214 N_VGND_c_374_n N_A_500_49#_M1006_d 0.00310634f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_c_371_n N_A_500_49#_c_418_n 0.00745539f $X=2.965 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_374_n N_A_500_49#_c_418_n 0.00686654f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_370_n N_A_500_49#_c_419_n 0.0139953f $X=3.07 $Y=0.39 $X2=0 $Y2=0
cc_218 N_VGND_c_371_n N_A_500_49#_c_419_n 0.00299122f $X=2.965 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_373_n N_A_500_49#_c_419_n 0.00299122f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_374_n N_A_500_49#_c_419_n 0.0108442f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_c_373_n N_A_500_49#_c_421_n 0.00831344f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_374_n N_A_500_49#_c_421_n 0.00760397f $X=3.6 $Y=0 $X2=0 $Y2=0
