# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a32o_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a32o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.180000 1.435000 6.085000 1.750000 ;
        RECT 5.425000 1.355000 6.085000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.455000 1.415000 4.205000 1.750000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.540000 1.425000 3.245000 1.750000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.615000 1.425000 7.045000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.355000 1.425000 8.005000 1.750000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.045000 1.820000 1.215000 ;
        RECT 0.100000 1.215000 0.335000 1.755000 ;
        RECT 0.100000 1.755000 1.970000 1.925000 ;
        RECT 0.700000 0.255000 0.890000 1.045000 ;
        RECT 0.880000 1.925000 1.070000 3.075000 ;
        RECT 1.560000 0.255000 1.820000 1.045000 ;
        RECT 1.740000 1.925000 1.970000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.200000  0.085000 0.530000 0.875000 ;
      RECT 0.380000  2.095000 0.710000 3.245000 ;
      RECT 0.505000  1.385000 2.195000 1.585000 ;
      RECT 1.060000  0.085000 1.390000 0.875000 ;
      RECT 1.240000  2.095000 1.570000 3.245000 ;
      RECT 2.010000  0.085000 2.340000 0.905000 ;
      RECT 2.025000  1.075000 4.520000 1.095000 ;
      RECT 2.025000  1.095000 6.760000 1.175000 ;
      RECT 2.025000  1.175000 5.255000 1.245000 ;
      RECT 2.025000  1.245000 2.195000 1.385000 ;
      RECT 2.140000  1.815000 2.370000 3.245000 ;
      RECT 2.530000  0.255000 2.860000 0.735000 ;
      RECT 2.530000  0.735000 3.580000 0.905000 ;
      RECT 2.540000  1.920000 6.085000 2.090000 ;
      RECT 2.540000  2.090000 2.790000 3.075000 ;
      RECT 2.960000  2.260000 3.290000 3.245000 ;
      RECT 3.030000  0.085000 3.240000 0.565000 ;
      RECT 3.410000  0.255000 4.520000 0.515000 ;
      RECT 3.410000  0.515000 3.580000 0.735000 ;
      RECT 3.760000  0.685000 4.895000 0.895000 ;
      RECT 3.865000  2.090000 4.240000 3.075000 ;
      RECT 4.350000  1.245000 5.255000 1.265000 ;
      RECT 4.410000  2.260000 4.740000 3.245000 ;
      RECT 4.690000  0.255000 5.810000 0.445000 ;
      RECT 4.690000  0.445000 4.895000 0.685000 ;
      RECT 4.690000  0.895000 4.895000 0.925000 ;
      RECT 4.910000  2.090000 5.100000 3.075000 ;
      RECT 5.065000  0.615000 5.310000 1.005000 ;
      RECT 5.065000  1.005000 6.760000 1.095000 ;
      RECT 5.270000  2.260000 5.600000 3.245000 ;
      RECT 5.480000  0.445000 5.810000 0.835000 ;
      RECT 5.770000  2.090000 6.085000 2.905000 ;
      RECT 5.770000  2.905000 8.040000 3.075000 ;
      RECT 6.000000  0.255000 7.120000 0.425000 ;
      RECT 6.000000  0.425000 6.260000 0.835000 ;
      RECT 6.255000  1.175000 6.435000 1.920000 ;
      RECT 6.255000  1.920000 7.610000 2.100000 ;
      RECT 6.255000  2.100000 6.535000 2.735000 ;
      RECT 6.430000  0.595000 6.760000 1.005000 ;
      RECT 6.775000  2.270000 7.105000 2.905000 ;
      RECT 6.930000  0.425000 7.120000 1.075000 ;
      RECT 6.930000  1.075000 8.050000 1.245000 ;
      RECT 7.280000  2.100000 7.610000 2.735000 ;
      RECT 7.290000  0.085000 7.620000 0.905000 ;
      RECT 7.780000  1.920000 8.040000 2.905000 ;
      RECT 7.790000  0.255000 8.050000 1.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__a32o_4
