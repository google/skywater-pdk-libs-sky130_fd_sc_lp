* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_lp A0 A1 S VGND VNB VPB VPWR X
X0 a_704_55# S a_200_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_84_29# a_123_527# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VPWR a_200_367# a_281_527# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_84_29# A1 a_516_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_516_55# S VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND S a_704_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_307_55# A0 a_84_29# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_281_527# A1 a_84_29# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR S a_702_527# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_702_527# S a_200_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_84_29# A0 a_445_527# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_114_55# a_84_29# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_200_367# a_307_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_445_527# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 X a_84_29# a_114_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_123_527# a_84_29# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
