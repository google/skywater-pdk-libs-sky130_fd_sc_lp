# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__einvp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705000 1.425000 4.375000 1.750000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.819000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.210000 3.240000 1.430000 ;
        RECT 2.875000 1.065000 3.240000 1.210000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  1.520400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.455000 0.605000 3.785000 1.085000 ;
        RECT 3.455000 1.085000 4.795000 1.255000 ;
        RECT 3.965000 1.920000 5.225000 2.090000 ;
        RECT 3.965000 2.090000 4.265000 2.735000 ;
        RECT 4.465000 0.615000 4.795000 1.085000 ;
        RECT 4.545000 1.255000 4.795000 1.385000 ;
        RECT 4.545000 1.385000 5.665000 1.555000 ;
        RECT 4.545000 1.555000 5.225000 1.920000 ;
        RECT 4.935000 2.090000 5.225000 2.735000 ;
        RECT 5.365000 0.325000 5.665000 1.385000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.135000  0.255000 0.430000 1.420000 ;
      RECT 0.135000  1.420000 1.345000 1.645000 ;
      RECT 0.135000  1.645000 0.430000 3.075000 ;
      RECT 0.600000  0.085000 0.860000 1.115000 ;
      RECT 0.600000  1.815000 0.895000 3.245000 ;
      RECT 1.030000  0.255000 1.255000 0.870000 ;
      RECT 1.030000  0.870000 3.190000 0.895000 ;
      RECT 1.030000  0.895000 2.705000 1.040000 ;
      RECT 1.065000  1.645000 1.345000 2.245000 ;
      RECT 1.425000  0.085000 1.755000 0.700000 ;
      RECT 1.515000  1.755000 3.535000 1.920000 ;
      RECT 1.515000  1.920000 3.795000 1.925000 ;
      RECT 1.515000  1.925000 1.725000 3.075000 ;
      RECT 1.895000  2.095000 2.225000 3.245000 ;
      RECT 1.925000  0.255000 2.115000 0.725000 ;
      RECT 1.925000  0.725000 3.190000 0.870000 ;
      RECT 2.285000  0.085000 2.615000 0.555000 ;
      RECT 2.395000  1.925000 2.585000 3.075000 ;
      RECT 2.755000  2.105000 3.085000 3.245000 ;
      RECT 2.840000  0.265000 5.195000 0.435000 ;
      RECT 2.840000  0.435000 3.190000 0.725000 ;
      RECT 3.255000  1.925000 3.795000 2.905000 ;
      RECT 3.255000  2.905000 5.665000 3.075000 ;
      RECT 3.965000  0.435000 4.295000 0.895000 ;
      RECT 4.435000  2.260000 4.765000 2.905000 ;
      RECT 4.965000  0.435000 5.195000 1.215000 ;
      RECT 5.395000  1.815000 5.665000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__einvp_4
END LIBRARY
