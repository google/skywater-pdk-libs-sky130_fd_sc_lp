* File: sky130_fd_sc_lp__a31o_4.pex.spice
* Created: Wed Sep  2 09:26:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31O_4%B1 3 7 9 13 17 19 20 21 25
r45 28 29 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=0.362 $Y=1.465
+ $X2=0.362 $Y2=1.54
r46 25 28 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=0.362 $Y=1.375
+ $X2=0.362 $Y2=1.465
r47 25 27 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=1.375
+ $X2=0.362 $Y2=1.21
r48 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.375 $X2=0.34 $Y2=1.375
r49 21 26 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=1.375
r50 20 26 3.41465 $w=2.68e-07 $l=8e-08 $layer=LI1_cond $X=0.29 $Y=1.295 $X2=0.29
+ $Y2=1.375
r51 15 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.54
+ $X2=0.905 $Y2=1.465
r52 15 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.905 $Y=1.54
+ $X2=0.905 $Y2=2.465
r53 11 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.39
+ $X2=0.905 $Y2=1.465
r54 11 13 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=0.905 $Y=1.39
+ $X2=0.905 $Y2=0.655
r55 10 28 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=0.55 $Y=1.465
+ $X2=0.362 $Y2=1.465
r56 9 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.465
+ $X2=0.905 $Y2=1.465
r57 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.465
+ $X2=0.55 $Y2=1.465
r58 7 29 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.54
r59 3 27 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.475 $Y=0.655
+ $X2=0.475 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%A_110_47# 1 2 3 12 14 15 18 20 22 25 27 29 32
+ 34 36 37 38 39 41 44 48 52 54 63 64 68 70 71
c167 71 0 1.9094e-19 $X=3.165 $Y=1.16
c168 32 0 1.65438e-19 $X=3.045 $Y=0.655
r169 78 79 35.3298 $w=3.82e-07 $l=2.8e-07 $layer=POLY_cond $X=2.765 $Y=1.52
+ $X2=3.045 $Y2=1.52
r170 77 78 42.9005 $w=3.82e-07 $l=3.4e-07 $layer=POLY_cond $X=2.425 $Y=1.52
+ $X2=2.765 $Y2=1.52
r171 76 77 11.356 $w=3.82e-07 $l=9e-08 $layer=POLY_cond $X=2.335 $Y=1.52
+ $X2=2.425 $Y2=1.52
r172 66 68 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=6.03 $Y=1.075
+ $X2=6.03 $Y2=0.71
r173 65 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=1.16
+ $X2=3.165 $Y2=1.16
r174 64 66 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.865 $Y=1.16
+ $X2=6.03 $Y2=1.075
r175 64 65 170.604 $w=1.68e-07 $l=2.615e-06 $layer=LI1_cond $X=5.865 $Y=1.16
+ $X2=3.25 $Y2=1.16
r176 63 71 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=1.075
+ $X2=3.165 $Y2=1.16
r177 62 63 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.165 $Y=0.805
+ $X2=3.165 $Y2=1.075
r178 61 81 15.1414 $w=3.82e-07 $l=1.2e-07 $layer=POLY_cond $X=3.075 $Y=1.52
+ $X2=3.195 $Y2=1.52
r179 61 79 3.78534 $w=3.82e-07 $l=3e-08 $layer=POLY_cond $X=3.075 $Y=1.52
+ $X2=3.045 $Y2=1.52
r180 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.075
+ $Y=1.48 $X2=3.075 $Y2=1.48
r181 57 76 35.3298 $w=3.82e-07 $l=2.8e-07 $layer=POLY_cond $X=2.055 $Y=1.52
+ $X2=2.335 $Y2=1.52
r182 57 74 7.57068 $w=3.82e-07 $l=6e-08 $layer=POLY_cond $X=2.055 $Y=1.52
+ $X2=1.995 $Y2=1.52
r183 56 60 40.5342 $w=2.88e-07 $l=1.02e-06 $layer=LI1_cond $X=2.055 $Y=1.5
+ $X2=3.075 $Y2=1.5
r184 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.055
+ $Y=1.48 $X2=2.055 $Y2=1.48
r185 54 71 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.165 $Y=1.5
+ $X2=3.165 $Y2=1.16
r186 54 60 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=3.08 $Y=1.5
+ $X2=3.075 $Y2=1.5
r187 53 70 2.36881 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.855 $Y=0.72
+ $X2=0.725 $Y2=0.72
r188 52 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.08 $Y=0.72
+ $X2=3.165 $Y2=0.805
r189 52 53 145.16 $w=1.68e-07 $l=2.225e-06 $layer=LI1_cond $X=3.08 $Y=0.72
+ $X2=0.855 $Y2=0.72
r190 48 50 49.4221 $w=2.58e-07 $l=1.115e-06 $layer=LI1_cond $X=0.725 $Y=0.865
+ $X2=0.725 $Y2=1.98
r191 46 70 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=0.72
r192 46 48 2.65948 $w=2.58e-07 $l=6e-08 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=0.865
r193 42 70 4.06715 $w=2.25e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.69 $Y=0.635
+ $X2=0.725 $Y2=0.72
r194 42 44 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=0.69 $Y=0.635
+ $X2=0.69 $Y2=0.42
r195 39 41 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.625 $Y=1.725
+ $X2=3.625 $Y2=2.465
r196 38 81 27.8964 $w=3.82e-07 $l=1.63248e-07 $layer=POLY_cond $X=3.27 $Y=1.65
+ $X2=3.195 $Y2=1.52
r197 37 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.55 $Y=1.65
+ $X2=3.625 $Y2=1.725
r198 37 38 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.55 $Y=1.65
+ $X2=3.27 $Y2=1.65
r199 34 81 24.74 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=3.195 $Y=1.725
+ $X2=3.195 $Y2=1.52
r200 34 36 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.195 $Y=1.725
+ $X2=3.195 $Y2=2.465
r201 30 79 24.74 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=3.045 $Y=1.315
+ $X2=3.045 $Y2=1.52
r202 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.045 $Y=1.315
+ $X2=3.045 $Y2=0.655
r203 27 78 24.74 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.765 $Y=1.725
+ $X2=2.765 $Y2=1.52
r204 27 29 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.765 $Y=1.725
+ $X2=2.765 $Y2=2.465
r205 23 77 24.74 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.425 $Y=1.315
+ $X2=2.425 $Y2=1.52
r206 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.425 $Y=1.315
+ $X2=2.425 $Y2=0.655
r207 20 76 24.74 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.335 $Y=1.725
+ $X2=2.335 $Y2=1.52
r208 20 22 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.335 $Y=1.725
+ $X2=2.335 $Y2=2.465
r209 16 74 24.74 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=1.995 $Y=1.315
+ $X2=1.995 $Y2=1.52
r210 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.995 $Y=1.315
+ $X2=1.995 $Y2=0.655
r211 14 74 31.6817 $w=3.82e-07 $l=1.74786e-07 $layer=POLY_cond $X=1.89 $Y=1.39
+ $X2=1.995 $Y2=1.52
r212 14 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.89 $Y=1.39
+ $X2=1.41 $Y2=1.39
r213 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.315
+ $X2=1.41 $Y2=1.39
r214 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.315
+ $X2=1.335 $Y2=0.655
r215 3 50 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=1.98
r216 2 68 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=5.89
+ $Y=0.335 $X2=6.03 $Y2=0.71
r217 1 48 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.865
r218 1 44 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%A3 1 3 4 5 6 8 11 13 17 20 22 23 24 25 30
c75 22 0 2.9237e-20 $X=4.075 $Y=1.6
c76 17 0 5.21438e-20 $X=4.485 $Y=2.465
c77 1 0 1.61703e-19 $X=3.555 $Y=1.185
r78 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.075
+ $Y=1.51 $X2=4.075 $Y2=1.51
r79 24 25 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.582
+ $X2=4.56 $Y2=1.582
r80 24 31 0.172006 $w=3.33e-07 $l=5e-09 $layer=LI1_cond $X=4.08 $Y=1.582
+ $X2=4.075 $Y2=1.582
r81 23 31 16.3406 $w=3.33e-07 $l=4.75e-07 $layer=LI1_cond $X=3.6 $Y=1.582
+ $X2=4.075 $Y2=1.582
r82 21 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.075 $Y=1.525
+ $X2=4.075 $Y2=1.51
r83 21 22 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.075 $Y=1.525
+ $X2=4.075 $Y2=1.6
r84 19 30 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=4.075 $Y=1.335
+ $X2=4.075 $Y2=1.51
r85 19 20 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.075 $Y=1.335
+ $X2=4.075 $Y2=1.26
r86 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.485 $Y=1.675
+ $X2=4.485 $Y2=2.465
r87 14 22 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.24 $Y=1.6
+ $X2=4.075 $Y2=1.6
r88 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.41 $Y=1.6
+ $X2=4.485 $Y2=1.675
r89 13 14 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.41 $Y=1.6 $X2=4.24
+ $Y2=1.6
r90 9 22 13.5877 $w=2.4e-07 $l=8.44097e-08 $layer=POLY_cond $X=4.055 $Y=1.675
+ $X2=4.075 $Y2=1.6
r91 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.055 $Y=1.675
+ $X2=4.055 $Y2=2.465
r92 6 20 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.985 $Y=1.185
+ $X2=4.075 $Y2=1.26
r93 6 8 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.985 $Y=1.185
+ $X2=3.985 $Y2=0.655
r94 4 20 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.91 $Y=1.26
+ $X2=4.075 $Y2=1.26
r95 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.91 $Y=1.26 $X2=3.63
+ $Y2=1.26
r96 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.555 $Y=1.185
+ $X2=3.63 $Y2=1.26
r97 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.555 $Y=1.185
+ $X2=3.555 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%A2 3 7 11 15 17 18 26
c49 18 0 5.21438e-20 $X=5.52 $Y=1.665
r50 24 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.295 $Y=1.51
+ $X2=5.385 $Y2=1.51
r51 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.295
+ $Y=1.51 $X2=5.295 $Y2=1.51
r52 21 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.955 $Y=1.51
+ $X2=5.295 $Y2=1.51
r53 18 25 7.51593 $w=3.43e-07 $l=2.25e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.295 $Y2=1.587
r54 17 25 8.51806 $w=3.43e-07 $l=2.55e-07 $layer=LI1_cond $X=5.04 $Y=1.587
+ $X2=5.295 $Y2=1.587
r55 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=1.51
r56 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=2.465
r57 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.345
+ $X2=5.385 $Y2=1.51
r58 9 11 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.385 $Y=1.345
+ $X2=5.385 $Y2=0.755
r59 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=4.955 $Y2=1.51
r60 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=4.955 $Y2=2.465
r61 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.955 $Y=1.345
+ $X2=4.955 $Y2=1.51
r62 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.955 $Y=1.345
+ $X2=4.955 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%A1 3 7 11 15 17 18 26
r41 24 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.155 $Y=1.51
+ $X2=6.245 $Y2=1.51
r42 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.155
+ $Y=1.51 $X2=6.155 $Y2=1.51
r43 21 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.815 $Y=1.51
+ $X2=6.155 $Y2=1.51
r44 18 25 10.8563 $w=3.43e-07 $l=3.25e-07 $layer=LI1_cond $X=6.48 $Y=1.587
+ $X2=6.155 $Y2=1.587
r45 17 25 5.17764 $w=3.43e-07 $l=1.55e-07 $layer=LI1_cond $X=6 $Y=1.587
+ $X2=6.155 $Y2=1.587
r46 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.675
+ $X2=6.245 $Y2=1.51
r47 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.245 $Y=1.675
+ $X2=6.245 $Y2=2.465
r48 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.345
+ $X2=6.245 $Y2=1.51
r49 9 11 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.245 $Y=1.345
+ $X2=6.245 $Y2=0.755
r50 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.815 $Y2=1.51
r51 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.815 $Y2=2.465
r52 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.345
+ $X2=5.815 $Y2=1.51
r53 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.815 $Y=1.345
+ $X2=5.815 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%A_27_367# 1 2 3 4 5 16 18 20 24 27 28 30 31
+ 34 36 40 42 44 46 50 55 57
r81 44 59 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=2.1 $X2=6.03
+ $Y2=2.015
r82 44 46 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=6.03 $Y=2.1 $X2=6.03
+ $Y2=2.91
r83 43 57 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.265 $Y=2.015
+ $X2=5.16 $Y2=2.015
r84 42 59 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.935 $Y=2.015
+ $X2=6.03 $Y2=2.015
r85 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.935 $Y=2.015
+ $X2=5.265 $Y2=2.015
r86 38 57 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=2.1 $X2=5.16
+ $Y2=2.015
r87 38 40 42.7792 $w=2.08e-07 $l=8.1e-07 $layer=LI1_cond $X=5.16 $Y=2.1 $X2=5.16
+ $Y2=2.91
r88 37 54 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.385 $Y=2.015
+ $X2=4.245 $Y2=2.015
r89 36 57 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.055 $Y=2.015
+ $X2=5.16 $Y2=2.015
r90 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.055 $Y=2.015
+ $X2=4.385 $Y2=2.015
r91 32 55 3.77418 $w=2.45e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.28 $Y=2.61
+ $X2=4.245 $Y2=2.525
r92 32 34 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=4.28 $Y=2.61 $X2=4.28
+ $Y2=2.91
r93 31 55 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=2.44
+ $X2=4.245 $Y2=2.525
r94 30 54 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=2.1
+ $X2=4.245 $Y2=2.015
r95 30 31 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=4.245 $Y=2.1
+ $X2=4.245 $Y2=2.44
r96 29 50 2.53056 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.285 $Y=2.525
+ $X2=1.155 $Y2=2.525
r97 28 55 2.68609 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.105 $Y=2.525
+ $X2=4.245 $Y2=2.525
r98 28 29 183.979 $w=1.68e-07 $l=2.82e-06 $layer=LI1_cond $X=4.105 $Y=2.525
+ $X2=1.285 $Y2=2.525
r99 27 52 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=2.905
+ $X2=1.155 $Y2=2.99
r100 26 50 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=2.61
+ $X2=1.155 $Y2=2.525
r101 26 27 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.155 $Y=2.61
+ $X2=1.155 $Y2=2.905
r102 22 50 3.91525 $w=2.35e-07 $l=9.66954e-08 $layer=LI1_cond $X=1.13 $Y=2.44
+ $X2=1.155 $Y2=2.525
r103 22 24 18.2208 $w=2.08e-07 $l=3.45e-07 $layer=LI1_cond $X=1.13 $Y=2.44
+ $X2=1.13 $Y2=2.095
r104 21 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=2.99
+ $X2=0.26 $Y2=2.99
r105 20 52 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.025 $Y=2.99
+ $X2=1.155 $Y2=2.99
r106 20 21 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.025 $Y=2.99
+ $X2=0.425 $Y2=2.99
r107 16 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.905
+ $X2=0.26 $Y2=2.99
r108 16 18 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=0.26 $Y=2.905
+ $X2=0.26 $Y2=2.095
r109 5 59 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=1.835 $X2=6.03 $Y2=2.095
r110 5 46 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=1.835 $X2=6.03 $Y2=2.91
r111 4 57 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=5.03
+ $Y=1.835 $X2=5.17 $Y2=2.095
r112 4 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.03
+ $Y=1.835 $X2=5.17 $Y2=2.91
r113 3 54 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=4.13
+ $Y=1.835 $X2=4.27 $Y2=2.095
r114 3 34 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.13
+ $Y=1.835 $X2=4.27 $Y2=2.91
r115 2 52 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.91
r116 2 24 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.095
r117 1 49 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r118 1 18 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%VPWR 1 2 3 4 5 6 21 25 29 31 35 39 41 43 48
+ 49 50 51 52 54 69 74 80 83 86 90
r105 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r106 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r107 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r108 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 78 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r110 78 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r111 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r112 75 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.6 $Y2=3.33
r113 75 77 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=6 $Y2=3.33
r114 74 89 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=6.295 $Y=3.33
+ $X2=6.507 $Y2=3.33
r115 74 77 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.295 $Y=3.33 $X2=6
+ $Y2=3.33
r116 73 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r117 73 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 70 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.885 $Y=3.33
+ $X2=4.72 $Y2=3.33
r120 70 72 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.885 $Y=3.33
+ $X2=5.04 $Y2=3.33
r121 69 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.6 $Y2=3.33
r122 69 72 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 68 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r124 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r125 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r127 62 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.12 $Y2=3.33
r128 62 64 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 61 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r131 57 61 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r132 56 60 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r133 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r134 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=2.12 $Y2=3.33
r135 54 60 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.68 $Y2=3.33
r136 52 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r137 52 65 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 50 67 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=3.6 $Y2=3.33
r139 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=3.84 $Y2=3.33
r140 48 64 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.64 $Y2=3.33
r141 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.98 $Y2=3.33
r142 47 67 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=3.6 $Y2=3.33
r143 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=2.98 $Y2=3.33
r144 43 46 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=6.46 $Y=2.015
+ $X2=6.46 $Y2=2.95
r145 41 89 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.46 $Y=3.245
+ $X2=6.507 $Y2=3.33
r146 41 46 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.46 $Y=3.245
+ $X2=6.46 $Y2=2.95
r147 37 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.6 $Y=3.245 $X2=5.6
+ $Y2=3.33
r148 37 39 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.6 $Y=3.245
+ $X2=5.6 $Y2=2.385
r149 33 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.72 $Y=3.245
+ $X2=4.72 $Y2=3.33
r150 33 35 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.72 $Y=3.245
+ $X2=4.72 $Y2=2.385
r151 32 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=3.33
+ $X2=3.84 $Y2=3.33
r152 31 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.555 $Y=3.33
+ $X2=4.72 $Y2=3.33
r153 31 32 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.555 $Y=3.33
+ $X2=4.005 $Y2=3.33
r154 27 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=3.245
+ $X2=3.84 $Y2=3.33
r155 27 29 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.84 $Y=3.245
+ $X2=3.84 $Y2=2.915
r156 23 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=3.245
+ $X2=2.98 $Y2=3.33
r157 23 25 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.98 $Y=3.245
+ $X2=2.98 $Y2=2.915
r158 19 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=3.33
r159 19 21 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.915
r160 6 46 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.95
r161 6 43 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.015
r162 5 39 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.385
r163 4 35 300 $w=1.7e-07 $l=6.249e-07 $layer=licon1_PDIFF $count=2 $X=4.56
+ $Y=1.835 $X2=4.72 $Y2=2.385
r164 3 29 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=1.835 $X2=3.84 $Y2=2.915
r165 2 25 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=2.84
+ $Y=1.835 $X2=2.98 $Y2=2.915
r166 1 21 600 $w=1.7e-07 $l=1.14079e-06 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.835 $X2=2.12 $Y2=2.915
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%X 1 2 3 4 14 17 19 23 25 26 30
r58 26 36 5.69422 $w=6.63e-07 $l=9.5e-08 $layer=LI1_cond $X=1.357 $Y=1.665
+ $X2=1.357 $Y2=1.76
r59 25 26 6.65487 $w=6.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.357 $Y=1.295
+ $X2=1.357 $Y2=1.665
r60 25 30 4.22674 $w=6.63e-07 $l=2.35e-07 $layer=LI1_cond $X=1.357 $Y=1.295
+ $X2=1.357 $Y2=1.06
r61 21 23 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.55 $Y=2.095
+ $X2=3.41 $Y2=2.095
r62 19 21 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=1.69 $Y=2.095
+ $X2=2.55 $Y2=2.095
r63 15 30 7.62298 $w=2.1e-07 $l=3.42854e-07 $layer=LI1_cond $X=1.69 $Y=1.08
+ $X2=1.357 $Y2=1.06
r64 15 17 55.1905 $w=2.08e-07 $l=1.045e-06 $layer=LI1_cond $X=1.69 $Y=1.08
+ $X2=2.735 $Y2=1.08
r65 14 19 6.86407 $w=3.3e-07 $l=2.25433e-07 $layer=LI1_cond $X=1.547 $Y=1.93
+ $X2=1.69 $Y2=2.095
r66 14 36 6.87422 $w=2.83e-07 $l=1.7e-07 $layer=LI1_cond $X=1.547 $Y=1.93
+ $X2=1.547 $Y2=1.76
r67 4 23 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=1.835 $X2=3.41 $Y2=2.095
r68 3 21 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.835 $X2=2.55 $Y2=2.095
r69 2 17 182 $w=1.7e-07 $l=9.35147e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.235 $X2=2.735 $Y2=1.06
r70 1 30 182 $w=1.7e-07 $l=9.43928e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.665 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%VGND 1 2 3 4 5 16 18 22 26 28 32 36 39 40 41
+ 43 48 61 62 68 71 74
r91 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r92 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r93 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r94 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r95 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r96 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r97 59 62 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r98 58 61 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r99 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r100 56 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r101 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r102 53 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.26
+ $Y2=0
r103 53 55 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.425 $Y=0
+ $X2=4.08 $Y2=0
r104 52 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r105 52 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r106 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r107 49 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r108 49 51 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.68 $Y2=0
r109 48 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=2.21
+ $Y2=0
r110 48 51 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=1.68 $Y2=0
r111 47 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r112 47 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r113 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r114 44 65 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r115 44 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r116 43 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r117 43 46 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=0
+ $X2=0.72 $Y2=0
r118 41 56 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r119 41 75 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r120 39 55 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.08
+ $Y2=0
r121 39 40 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.205
+ $Y2=0
r122 38 58 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.305 $Y=0
+ $X2=4.56 $Y2=0
r123 38 40 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.205
+ $Y2=0
r124 34 40 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=0.085
+ $X2=4.205 $Y2=0
r125 34 36 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=4.205 $Y=0.085
+ $X2=4.205 $Y2=0.38
r126 30 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=0.085
+ $X2=3.26 $Y2=0
r127 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.26 $Y=0.085
+ $X2=3.26 $Y2=0.36
r128 29 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.21
+ $Y2=0
r129 28 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=3.26
+ $Y2=0
r130 28 29 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.095 $Y=0
+ $X2=2.375 $Y2=0
r131 24 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r132 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.36
r133 20 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r134 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.36
r135 16 65 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r136 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r137 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.235 $X2=4.2 $Y2=0.38
r138 4 32 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.12
+ $Y=0.235 $X2=3.26 $Y2=0.36
r139 3 26 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.235 $X2=2.21 $Y2=0.36
r140 2 22 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.36
r141 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%A_726_47# 1 2 9 11 13
c31 11 0 1.65438e-19 $X=3.935 $Y=0.815
r32 11 13 76.096 $w=1.78e-07 $l=1.235e-06 $layer=LI1_cond $X=3.935 $Y=0.815
+ $X2=5.17 $Y2=0.815
r33 7 11 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.77 $Y=0.725
+ $X2=3.935 $Y2=0.815
r34 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.77 $Y=0.725
+ $X2=3.77 $Y2=0.45
r35 2 13 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.335 $X2=5.17 $Y2=0.81
r36 1 9 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=3.63
+ $Y=0.235 $X2=3.77 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_4%A_919_67# 1 2 3 14 18 22 23
r27 21 23 6.35851 $w=3.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.6 $Y=0.46
+ $X2=5.695 $Y2=0.46
r28 21 22 3.3566 $w=3.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.6 $Y=0.46 $X2=5.515
+ $Y2=0.46
r29 16 18 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=6.495 $Y=0.445
+ $X2=6.495 $Y2=0.48
r30 14 16 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.365 $Y=0.36
+ $X2=6.495 $Y2=0.445
r31 14 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.365 $Y=0.36
+ $X2=5.695 $Y2=0.36
r32 12 22 31.898 $w=2.78e-07 $l=7.75e-07 $layer=LI1_cond $X=4.74 $Y=0.415
+ $X2=5.515 $Y2=0.415
r33 3 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.32
+ $Y=0.335 $X2=6.46 $Y2=0.48
r34 2 21 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.335 $X2=5.6 $Y2=0.46
r35 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.595
+ $Y=0.335 $X2=4.74 $Y2=0.46
.ends

