* File: sky130_fd_sc_lp__dfxbp_lp.spice
* Created: Wed Sep  2 09:45:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfxbp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dfxbp_lp  VNB VPB CLK D VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1018 A_125_85# N_CLK_M1018_g N_A_27_403#_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_CLK_M1006_g A_125_85# VNB NSHORT L=0.15 W=0.42 AD=0.0735
+ AS=0.0441 PD=0.77 PS=0.63 NRD=19.992 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75002.7
+ A=0.063 P=1.14 MULT=1
MM1000 A_297_85# N_D_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0735 PD=0.63 PS=0.77 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_239_403#_M1002_d N_D_M1002_g A_297_85# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1016 N_A_455_85#_M1016_d N_A_27_403#_M1016_g N_A_239_403#_M1002_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.11705 AS=0.0588 PD=1.03 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1029 A_573_119# N_A_511_218#_M1029_g N_A_455_85#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.11705 PD=0.63 PS=1.03 NRD=14.28 NRS=22.848 M=1 R=2.8
+ SA=75001.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_615_93#_M1019_g A_573_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1098 AS=0.0441 PD=0.98 PS=0.63 NRD=24.276 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1030 A_763_119# N_A_455_85#_M1030_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1098 PD=0.63 PS=0.98 NRD=14.28 NRS=24.276 M=1 R=2.8 SA=75002.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_A_615_93#_M1020_d N_A_455_85#_M1020_g A_763_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75002.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1034 A_1049_125# N_A_27_403#_M1034_g N_A_511_218#_M1034_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1736 PD=0.63 PS=1.71 NRD=14.28 NRS=24.276 M=1 R=2.8
+ SA=75000.3 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_27_403#_M1009_g A_1049_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_A_1339_153#_M1022_d N_A_27_403#_M1022_g N_A_1232_153#_M1022_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.098325 AS=0.1617 PD=0.96 PS=1.61 NRD=49.992
+ NRS=28.56 M=1 R=2.8 SA=75000.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1031 N_A_615_93#_M1031_d N_A_511_218#_M1031_g N_A_1339_153#_M1022_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1176 AS=0.098325 PD=1.4 PS=0.96 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1507_321#_M1010_g N_A_1232_153#_M1010_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1024 A_1742_57# N_A_1339_153#_M1024_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_A_1507_321#_M1015_d N_A_1339_153#_M1015_g A_1742_57# VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 A_2010_127# N_A_1507_321#_M1011_g N_Q_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_1507_321#_M1017_g A_2010_127# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_2168_127# N_A_1507_321#_M1003_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_2062_367#_M1012_d N_A_1507_321#_M1012_g A_2168_127# VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 A_2436_57# N_A_2062_367#_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_Q_N_M1025_d N_A_2062_367#_M1025_g A_2436_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_CLK_M1013_g N_A_27_403#_M1013_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1028 N_A_239_403#_M1028_d N_D_M1028_g N_VPWR_M1013_d VPB PHIGHVT L=0.25 W=1
+ AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000 A=0.25
+ P=2.5 MULT=1
MM1026 N_A_455_85#_M1026_d N_A_27_403#_M1026_g N_A_349_323#_M1026_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1008 N_A_239_403#_M1008_d N_A_511_218#_M1008_g N_A_455_85#_M1026_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_615_93#_M1004_g N_A_349_323#_M1004_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1027 N_A_615_93#_M1027_d N_A_455_85#_M1027_g N_VPWR_M1004_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1033 N_VPWR_M1033_d N_A_27_403#_M1033_g N_A_511_218#_M1033_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1023 N_A_1339_153#_M1023_d N_A_27_403#_M1023_g N_A_615_93#_M1023_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1005 A_1445_419# N_A_511_218#_M1005_g N_A_1339_153#_M1023_d VPB PHIGHVT L=0.25
+ W=1 AD=0.155 AS=0.14 PD=1.31 PS=1.28 NRD=19.6803 NRS=0 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1021 N_VPWR_M1021_d N_A_1507_321#_M1021_g A_1445_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.29 AS=0.155 PD=1.58 PS=1.31 NRD=6.8753 NRS=19.6803 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1035 N_A_1507_321#_M1035_d N_A_1339_153#_M1035_g N_VPWR_M1021_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.29 PD=2.57 PS=1.58 NRD=0 NRS=52.1853 M=1 R=4
+ SA=125002 SB=125000 A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A_1507_321#_M1007_g N_Q_M1007_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1014 N_A_2062_367#_M1014_d N_A_1507_321#_M1014_g N_VPWR_M1007_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1001 N_Q_N_M1001_d N_A_2062_367#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX36_noxref VNB VPB NWDIODE A=25.5606 P=30.91
*
.include "sky130_fd_sc_lp__dfxbp_lp.pxi.spice"
*
.ends
*
*
