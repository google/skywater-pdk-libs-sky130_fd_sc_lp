* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
X0 a_247_367# a_329_269# a_367_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_33_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_1708_411# a_359_367# a_1758_87# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 a_1340_412# CI VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_359_367# B a_33_367# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 a_1034_380# a_367_119# COUT_N VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 a_33_367# a_329_269# a_359_367# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 COUT_N a_359_367# a_1340_412# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_1571_367# a_359_367# a_1758_87# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 VPWR CI a_1571_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND a_33_367# a_247_367# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 COUT_N a_367_119# a_1340_412# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_329_269# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_33_367# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_1758_87# a_367_119# a_1571_367# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 VPWR a_1758_87# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_33_367# a_329_269# a_367_119# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_329_269# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_1708_411# a_1571_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND CI a_1571_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VGND a_1758_87# SUM VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_1708_411# a_1571_367# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 VPWR a_33_367# a_247_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_359_367# B a_247_367# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 VGND B a_1034_380# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_1034_380# a_359_367# COUT_N VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 a_247_367# a_329_269# a_359_367# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 a_1340_412# CI VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 a_367_119# B a_247_367# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X29 a_1758_87# a_367_119# a_1708_411# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 VPWR B a_1034_380# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_367_119# B a_33_367# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
