* File: sky130_fd_sc_lp__dfrbp_1.pxi.spice
* Created: Fri Aug 28 10:21:33 2020
* 
x_PM_SKY130_FD_SC_LP__DFRBP_1%CLK N_CLK_M1027_g N_CLK_M1012_g CLK CLK
+ N_CLK_c_248_n PM_SKY130_FD_SC_LP__DFRBP_1%CLK
x_PM_SKY130_FD_SC_LP__DFRBP_1%D N_D_M1022_g N_D_M1013_g N_D_c_280_n N_D_c_281_n
+ N_D_c_286_n D D N_D_c_283_n PM_SKY130_FD_SC_LP__DFRBP_1%D
x_PM_SKY130_FD_SC_LP__DFRBP_1%A_197_108# N_A_197_108#_M1014_d
+ N_A_197_108#_M1028_d N_A_197_108#_c_327_n N_A_197_108#_M1018_g
+ N_A_197_108#_c_328_n N_A_197_108#_M1019_g N_A_197_108#_c_329_n
+ N_A_197_108#_M1021_g N_A_197_108#_c_330_n N_A_197_108#_M1002_g
+ N_A_197_108#_c_348_n N_A_197_108#_c_349_n N_A_197_108#_c_331_n
+ N_A_197_108#_c_350_n N_A_197_108#_c_332_n N_A_197_108#_c_333_n
+ N_A_197_108#_c_334_n N_A_197_108#_c_335_n N_A_197_108#_c_336_n
+ N_A_197_108#_c_337_n N_A_197_108#_c_338_n N_A_197_108#_c_352_n
+ N_A_197_108#_c_339_n N_A_197_108#_c_353_n N_A_197_108#_c_340_n
+ N_A_197_108#_c_341_n N_A_197_108#_c_342_n N_A_197_108#_c_343_n
+ PM_SKY130_FD_SC_LP__DFRBP_1%A_197_108#
x_PM_SKY130_FD_SC_LP__DFRBP_1%A_804_328# N_A_804_328#_M1020_d
+ N_A_804_328#_M1032_d N_A_804_328#_M1010_g N_A_804_328#_M1009_g
+ N_A_804_328#_c_520_n N_A_804_328#_c_521_n N_A_804_328#_c_522_n
+ N_A_804_328#_c_523_n N_A_804_328#_c_524_n N_A_804_328#_c_531_n
+ N_A_804_328#_c_532_n N_A_804_328#_c_525_n N_A_804_328#_c_534_n
+ N_A_804_328#_c_526_n N_A_804_328#_c_548_n
+ PM_SKY130_FD_SC_LP__DFRBP_1%A_804_328#
x_PM_SKY130_FD_SC_LP__DFRBP_1%RESET_B N_RESET_B_M1025_g N_RESET_B_M1000_g
+ N_RESET_B_c_629_n N_RESET_B_c_630_n N_RESET_B_M1026_g N_RESET_B_M1015_g
+ N_RESET_B_M1017_g N_RESET_B_M1016_g N_RESET_B_c_633_n N_RESET_B_c_641_n
+ N_RESET_B_c_642_n N_RESET_B_c_643_n N_RESET_B_c_644_n N_RESET_B_c_645_n
+ RESET_B N_RESET_B_c_634_n N_RESET_B_c_635_n N_RESET_B_c_648_n
+ N_RESET_B_c_649_n N_RESET_B_c_650_n N_RESET_B_c_651_n
+ PM_SKY130_FD_SC_LP__DFRBP_1%RESET_B
x_PM_SKY130_FD_SC_LP__DFRBP_1%A_603_191# N_A_603_191#_M1003_d
+ N_A_603_191#_M1018_d N_A_603_191#_M1015_d N_A_603_191#_c_827_n
+ N_A_603_191#_M1020_g N_A_603_191#_M1032_g N_A_603_191#_c_828_n
+ N_A_603_191#_c_866_n N_A_603_191#_c_833_n N_A_603_191#_c_834_n
+ N_A_603_191#_c_846_n N_A_603_191#_c_829_n N_A_603_191#_c_849_n
+ N_A_603_191#_c_879_n N_A_603_191#_c_830_n
+ PM_SKY130_FD_SC_LP__DFRBP_1%A_603_191#
x_PM_SKY130_FD_SC_LP__DFRBP_1%A_28_108# N_A_28_108#_M1027_s N_A_28_108#_M1012_s
+ N_A_28_108#_M1014_g N_A_28_108#_M1028_g N_A_28_108#_c_928_n
+ N_A_28_108#_c_929_n N_A_28_108#_c_939_n N_A_28_108#_c_940_n
+ N_A_28_108#_c_930_n N_A_28_108#_M1003_g N_A_28_108#_c_943_n
+ N_A_28_108#_M1011_g N_A_28_108#_c_945_n N_A_28_108#_M1029_g
+ N_A_28_108#_M1005_g N_A_28_108#_c_947_n N_A_28_108#_c_948_n
+ N_A_28_108#_c_949_n N_A_28_108#_c_933_n N_A_28_108#_c_934_n
+ N_A_28_108#_c_935_n N_A_28_108#_c_936_n N_A_28_108#_c_937_n
+ PM_SKY130_FD_SC_LP__DFRBP_1%A_28_108#
x_PM_SKY130_FD_SC_LP__DFRBP_1%A_1440_304# N_A_1440_304#_M1024_d
+ N_A_1440_304#_M1016_d N_A_1440_304#_M1001_g N_A_1440_304#_M1033_g
+ N_A_1440_304#_c_1086_n N_A_1440_304#_c_1087_n N_A_1440_304#_c_1079_n
+ N_A_1440_304#_c_1080_n N_A_1440_304#_c_1081_n N_A_1440_304#_c_1082_n
+ N_A_1440_304#_c_1090_n N_A_1440_304#_c_1091_n N_A_1440_304#_c_1083_n
+ N_A_1440_304#_c_1084_n PM_SKY130_FD_SC_LP__DFRBP_1%A_1440_304#
x_PM_SKY130_FD_SC_LP__DFRBP_1%A_1245_128# N_A_1245_128#_M1021_d
+ N_A_1245_128#_M1029_d N_A_1245_128#_c_1173_n N_A_1245_128#_M1024_g
+ N_A_1245_128#_M1006_g N_A_1245_128#_M1031_g N_A_1245_128#_M1030_g
+ N_A_1245_128#_M1023_g N_A_1245_128#_M1008_g N_A_1245_128#_c_1177_n
+ N_A_1245_128#_c_1204_n N_A_1245_128#_c_1205_n N_A_1245_128#_c_1206_n
+ N_A_1245_128#_c_1178_n N_A_1245_128#_c_1179_n N_A_1245_128#_c_1180_n
+ N_A_1245_128#_c_1181_n N_A_1245_128#_c_1182_n N_A_1245_128#_c_1183_n
+ N_A_1245_128#_c_1184_n N_A_1245_128#_c_1185_n N_A_1245_128#_c_1186_n
+ N_A_1245_128#_c_1187_n N_A_1245_128#_c_1188_n N_A_1245_128#_c_1189_n
+ N_A_1245_128#_c_1190_n N_A_1245_128#_c_1191_n N_A_1245_128#_c_1192_n
+ N_A_1245_128#_c_1193_n N_A_1245_128#_c_1194_n N_A_1245_128#_c_1195_n
+ N_A_1245_128#_c_1196_n N_A_1245_128#_c_1197_n N_A_1245_128#_c_1198_n
+ N_A_1245_128#_c_1199_n PM_SKY130_FD_SC_LP__DFRBP_1%A_1245_128#
x_PM_SKY130_FD_SC_LP__DFRBP_1%A_1796_139# N_A_1796_139#_M1031_s
+ N_A_1796_139#_M1030_s N_A_1796_139#_M1007_g N_A_1796_139#_c_1375_n
+ N_A_1796_139#_M1004_g N_A_1796_139#_c_1376_n N_A_1796_139#_c_1377_n
+ N_A_1796_139#_c_1383_n N_A_1796_139#_c_1384_n N_A_1796_139#_c_1385_n
+ N_A_1796_139#_c_1386_n N_A_1796_139#_c_1378_n N_A_1796_139#_c_1379_n
+ PM_SKY130_FD_SC_LP__DFRBP_1%A_1796_139#
x_PM_SKY130_FD_SC_LP__DFRBP_1%VPWR N_VPWR_M1012_d N_VPWR_M1025_d N_VPWR_M1009_d
+ N_VPWR_M1032_s N_VPWR_M1001_d N_VPWR_M1006_d N_VPWR_M1030_d N_VPWR_M1004_d
+ N_VPWR_c_1458_n N_VPWR_c_1459_n N_VPWR_c_1460_n N_VPWR_c_1461_n
+ N_VPWR_c_1462_n N_VPWR_c_1463_n N_VPWR_c_1464_n N_VPWR_c_1465_n
+ N_VPWR_c_1466_n N_VPWR_c_1467_n N_VPWR_c_1468_n N_VPWR_c_1469_n
+ N_VPWR_c_1470_n N_VPWR_c_1471_n VPWR N_VPWR_c_1472_n N_VPWR_c_1473_n
+ N_VPWR_c_1474_n N_VPWR_c_1475_n N_VPWR_c_1476_n N_VPWR_c_1477_n
+ N_VPWR_c_1457_n N_VPWR_c_1479_n N_VPWR_c_1480_n N_VPWR_c_1481_n
+ N_VPWR_c_1482_n N_VPWR_c_1483_n PM_SKY130_FD_SC_LP__DFRBP_1%VPWR
x_PM_SKY130_FD_SC_LP__DFRBP_1%A_304_463# N_A_304_463#_M1022_d
+ N_A_304_463#_M1025_s N_A_304_463#_M1013_d N_A_304_463#_M1018_s
+ N_A_304_463#_c_1603_n N_A_304_463#_c_1599_n N_A_304_463#_c_1601_n
+ N_A_304_463#_c_1608_n N_A_304_463#_c_1602_n
+ PM_SKY130_FD_SC_LP__DFRBP_1%A_304_463#
x_PM_SKY130_FD_SC_LP__DFRBP_1%Q N_Q_M1007_d N_Q_M1004_s N_Q_c_1650_n Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DFRBP_1%Q
x_PM_SKY130_FD_SC_LP__DFRBP_1%Q_N N_Q_N_M1008_d N_Q_N_M1023_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1683_n Q_N Q_N PM_SKY130_FD_SC_LP__DFRBP_1%Q_N
x_PM_SKY130_FD_SC_LP__DFRBP_1%VGND N_VGND_M1027_d N_VGND_M1000_s N_VGND_M1026_d
+ N_VGND_M1033_d N_VGND_M1031_d N_VGND_M1008_s N_VGND_c_1703_n N_VGND_c_1704_n
+ N_VGND_c_1705_n N_VGND_c_1706_n N_VGND_c_1707_n N_VGND_c_1708_n
+ N_VGND_c_1709_n N_VGND_c_1710_n VGND N_VGND_c_1711_n N_VGND_c_1712_n
+ N_VGND_c_1713_n N_VGND_c_1714_n N_VGND_c_1715_n N_VGND_c_1716_n
+ N_VGND_c_1717_n N_VGND_c_1718_n N_VGND_c_1719_n N_VGND_c_1720_n
+ N_VGND_c_1721_n N_VGND_c_1722_n PM_SKY130_FD_SC_LP__DFRBP_1%VGND
cc_1 VNB N_CLK_M1027_g 0.0543851f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.75
cc_2 VNB CLK 0.00340066f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_CLK_c_248_n 0.00727691f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.805
cc_4 VNB N_D_c_280_n 0.0146013f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_5 VNB N_D_c_281_n 0.00439427f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_6 VNB D 0.00238816f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.805
cc_7 VNB N_D_c_283_n 0.01534f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.97
cc_8 VNB N_A_197_108#_c_327_n 0.0408163f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.68
cc_9 VNB N_A_197_108#_c_328_n 0.0152662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_197_108#_c_329_n 0.0187936f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.805
cc_11 VNB N_A_197_108#_c_330_n 0.0196671f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.97
cc_12 VNB N_A_197_108#_c_331_n 0.00224464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_197_108#_c_332_n 0.00702301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_197_108#_c_333_n 0.0105577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_197_108#_c_334_n 0.0210839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_197_108#_c_335_n 0.00772868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_197_108#_c_336_n 0.0351452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_197_108#_c_337_n 0.0072662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_197_108#_c_338_n 0.00164008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_197_108#_c_339_n 0.0128953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_197_108#_c_340_n 0.00377967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_197_108#_c_341_n 0.00236147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_197_108#_c_342_n 9.94774e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_197_108#_c_343_n 0.0314405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_804_328#_M1010_g 0.0222254f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_26 VNB N_A_804_328#_c_520_n 4.88773e-19 $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.97
cc_27 VNB N_A_804_328#_c_521_n 0.0105578f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.665
cc_28 VNB N_A_804_328#_c_522_n 0.0157463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_804_328#_c_523_n 0.00207767f $X=-0.19 $Y=-0.245 $X2=0.722
+ $Y2=1.805
cc_30 VNB N_A_804_328#_c_524_n 0.00236129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_804_328#_c_525_n 0.00246865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_804_328#_c_526_n 0.00181111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_RESET_B_M1000_g 0.0279719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_RESET_B_c_629_n 0.135146f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_35 VNB N_RESET_B_c_630_n 0.00872874f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_36 VNB N_RESET_B_M1026_g 0.0452928f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.805
cc_37 VNB N_RESET_B_M1017_g 0.0383638f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.805
cc_38 VNB N_RESET_B_c_633_n 0.0284986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_RESET_B_c_634_n 0.00610837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_RESET_B_c_635_n 0.00573509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_603_191#_c_827_n 0.0183742f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_42 VNB N_A_603_191#_c_828_n 0.00295285f $X=-0.19 $Y=-0.245 $X2=0.722
+ $Y2=1.665
cc_43 VNB N_A_603_191#_c_829_n 0.004564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_603_191#_c_830_n 0.0346718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_28_108#_M1014_g 0.0249026f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_46 VNB N_A_28_108#_c_928_n 0.435506f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.805
cc_47 VNB N_A_28_108#_c_929_n 0.0125018f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.64
cc_48 VNB N_A_28_108#_c_930_n 0.0156854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_28_108#_M1003_g 0.0274938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_28_108#_M1005_g 0.0434183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_28_108#_c_933_n 0.0195622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_28_108#_c_934_n 0.0128535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_28_108#_c_935_n 0.00457742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_28_108#_c_936_n 0.0370724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_28_108#_c_937_n 0.0167985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1440_304#_M1033_g 0.0377893f $X=-0.19 $Y=-0.245 $X2=0.592
+ $Y2=1.805
cc_57 VNB N_A_1440_304#_c_1079_n 0.0101336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1440_304#_c_1080_n 0.0126465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1440_304#_c_1081_n 4.57574e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1440_304#_c_1082_n 0.0137528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1440_304#_c_1083_n 0.00499034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1440_304#_c_1084_n 0.00266861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1245_128#_c_1173_n 0.0205761f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.68
cc_64 VNB N_A_1245_128#_M1006_g 0.0104047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1245_128#_M1031_g 0.0250038f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.64
cc_66 VNB N_A_1245_128#_M1023_g 0.00826167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1245_128#_c_1177_n 0.0121125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1245_128#_c_1178_n 0.00206495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1245_128#_c_1179_n 0.0264918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1245_128#_c_1180_n 0.0022574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1245_128#_c_1181_n 0.0225149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1245_128#_c_1182_n 0.00305626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1245_128#_c_1183_n 0.00119275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1245_128#_c_1184_n 0.00354838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1245_128#_c_1185_n 0.00144766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1245_128#_c_1186_n 0.00113942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1245_128#_c_1187_n 0.017694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1245_128#_c_1188_n 0.0143163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1245_128#_c_1189_n 0.00255324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1245_128#_c_1190_n 0.001778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1245_128#_c_1191_n 0.00102037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1245_128#_c_1192_n 0.0172897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1245_128#_c_1193_n 0.00209164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1245_128#_c_1194_n 0.00124146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1245_128#_c_1195_n 0.0015064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1245_128#_c_1196_n 0.041584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1245_128#_c_1197_n 0.0013953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1245_128#_c_1198_n 0.0439506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1245_128#_c_1199_n 0.0222104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1796_139#_M1007_g 0.0251298f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_91 VNB N_A_1796_139#_c_1375_n 0.0236871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1796_139#_c_1376_n 0.00542107f $X=-0.19 $Y=-0.245 $X2=0.592
+ $Y2=1.97
cc_93 VNB N_A_1796_139#_c_1377_n 0.00798375f $X=-0.19 $Y=-0.245 $X2=0.722
+ $Y2=1.665
cc_94 VNB N_A_1796_139#_c_1378_n 0.00209865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1796_139#_c_1379_n 0.0263323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VPWR_c_1457_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_304_463#_c_1599_n 0.00211387f $X=-0.19 $Y=-0.245 $X2=0.592
+ $Y2=1.64
cc_98 VNB N_Q_c_1650_n 0.00254822f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_99 VNB Q 0.00668751f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.805
cc_100 VNB Q_N 0.00617949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB Q_N 0.0289342f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_102 VNB N_Q_N_c_1683_n 0.0272323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1703_n 0.0172278f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.805
cc_104 VNB N_VGND_c_1704_n 0.0167178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1705_n 0.0199285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1706_n 0.0180421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1707_n 0.0127933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1708_n 0.00636224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1709_n 0.0563798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1710_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1711_n 0.0196239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1712_n 0.0203368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1713_n 0.0905011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1714_n 0.0488524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1715_n 0.0200035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1716_n 0.0152818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1717_n 0.575757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1718_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1719_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1720_n 0.00436638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1721_n 0.00631381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1722_n 0.00510065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VPB N_CLK_M1012_g 0.0352707f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.68
cc_124 VPB CLK 0.00556834f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_125 VPB N_CLK_c_248_n 0.0295174f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.805
cc_126 VPB N_D_M1013_g 0.0203377f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.68
cc_127 VPB N_D_c_281_n 0.0186592f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_128 VPB N_D_c_286_n 0.0156029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB D 0.0071827f $X=-0.19 $Y=1.655 $X2=0.592 $Y2=1.805
cc_130 VPB N_A_197_108#_c_327_n 0.0216591f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.68
cc_131 VPB N_A_197_108#_M1018_g 0.0315989f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_132 VPB N_A_197_108#_c_330_n 0.0128033f $X=-0.19 $Y=1.655 $X2=0.592 $Y2=1.97
cc_133 VPB N_A_197_108#_M1002_g 0.0444667f $X=-0.19 $Y=1.655 $X2=0.722 $Y2=1.805
cc_134 VPB N_A_197_108#_c_348_n 0.00231305f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_197_108#_c_349_n 0.00944566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_197_108#_c_350_n 0.00211549f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_197_108#_c_338_n 0.00116442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_197_108#_c_352_n 0.00351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_197_108#_c_353_n 0.00291651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_197_108#_c_342_n 0.00257657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_197_108#_c_343_n 0.015659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_804_328#_M1009_g 0.0290994f $X=-0.19 $Y=1.655 $X2=0.592 $Y2=1.805
cc_143 VPB N_A_804_328#_c_520_n 7.97285e-19 $X=-0.19 $Y=1.655 $X2=0.592 $Y2=1.97
cc_144 VPB N_A_804_328#_c_521_n 0.0249525f $X=-0.19 $Y=1.655 $X2=0.722 $Y2=1.665
cc_145 VPB N_A_804_328#_c_524_n 0.00465647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_804_328#_c_531_n 0.00458022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_804_328#_c_532_n 0.00369927f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_804_328#_c_525_n 0.00470065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_804_328#_c_534_n 0.00155678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_M1025_g 0.022151f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.75
cc_151 VPB N_RESET_B_M1026_g 0.00428474f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.805
cc_152 VPB N_RESET_B_M1015_g 0.0262624f $X=-0.19 $Y=1.655 $X2=0.592 $Y2=1.97
cc_153 VPB N_RESET_B_M1017_g 0.0111639f $X=-0.19 $Y=1.655 $X2=0.722 $Y2=1.805
cc_154 VPB N_RESET_B_M1016_g 0.0221339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_RESET_B_c_641_n 0.0172538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_RESET_B_c_642_n 0.0270215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_RESET_B_c_643_n 0.00443677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_RESET_B_c_644_n 0.029004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_RESET_B_c_645_n 0.00339961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_c_634_n 0.0210606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_RESET_B_c_635_n 0.00427478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_RESET_B_c_648_n 0.0416059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_RESET_B_c_649_n 0.00308769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_RESET_B_c_650_n 0.00140938f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_RESET_B_c_651_n 0.0359634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_603_191#_M1032_g 0.023071f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.805
cc_167 VPB N_A_603_191#_c_828_n 0.00956442f $X=-0.19 $Y=1.655 $X2=0.722
+ $Y2=1.665
cc_168 VPB N_A_603_191#_c_833_n 0.00792034f $X=-0.19 $Y=1.655 $X2=0.722
+ $Y2=1.805
cc_169 VPB N_A_603_191#_c_834_n 0.00189327f $X=-0.19 $Y=1.655 $X2=0.722
+ $Y2=2.035
cc_170 VPB N_A_603_191#_c_829_n 0.00151023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_603_191#_c_830_n 0.0148336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_28_108#_M1028_g 0.00924361f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.805
cc_173 VPB N_A_28_108#_c_939_n 0.136129f $X=-0.19 $Y=1.655 $X2=0.592 $Y2=1.97
cc_174 VPB N_A_28_108#_c_940_n 0.0107679f $X=-0.19 $Y=1.655 $X2=0.722 $Y2=1.665
cc_175 VPB N_A_28_108#_c_930_n 0.0250061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_28_108#_M1003_g 0.0738999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_28_108#_c_943_n 0.0528886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_28_108#_M1011_g 0.0361143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_28_108#_c_945_n 0.190742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_28_108#_M1029_g 0.025817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_28_108#_c_947_n 0.0218858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_28_108#_c_948_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_28_108#_c_949_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_28_108#_c_934_n 0.0639424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1440_304#_M1001_g 0.0218928f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_186 VPB N_A_1440_304#_c_1086_n 0.0213368f $X=-0.19 $Y=1.655 $X2=0.592
+ $Y2=1.97
cc_187 VPB N_A_1440_304#_c_1087_n 0.0154481f $X=-0.19 $Y=1.655 $X2=0.722
+ $Y2=1.665
cc_188 VPB N_A_1440_304#_c_1081_n 0.00276896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1440_304#_c_1082_n 0.00166117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_1440_304#_c_1090_n 0.00128987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_1440_304#_c_1091_n 0.00288055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_1440_304#_c_1083_n 0.00695162f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_1440_304#_c_1084_n 0.00939396f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_1245_128#_M1006_g 0.051983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_1245_128#_M1030_g 0.0448978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1245_128#_M1023_g 0.0243223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_1245_128#_c_1177_n 0.0157175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_1245_128#_c_1204_n 0.0201831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_1245_128#_c_1205_n 0.00353693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_1245_128#_c_1206_n 0.00697592f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1245_128#_c_1186_n 0.00455141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1245_128#_c_1189_n 0.00733717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1796_139#_c_1375_n 0.0092796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1796_139#_M1004_g 0.024046f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.805
cc_205 VPB N_A_1796_139#_c_1377_n 0.0111582f $X=-0.19 $Y=1.655 $X2=0.722
+ $Y2=1.665
cc_206 VPB N_A_1796_139#_c_1383_n 0.0104996f $X=-0.19 $Y=1.655 $X2=0.722
+ $Y2=1.805
cc_207 VPB N_A_1796_139#_c_1384_n 0.0216885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_1796_139#_c_1385_n 0.0090318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_1796_139#_c_1386_n 0.00794669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_1796_139#_c_1378_n 0.00201399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_1796_139#_c_1379_n 0.0125336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1458_n 0.00377124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1459_n 0.0111049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1460_n 0.0139596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1461_n 0.0191964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1462_n 0.0197944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1463_n 0.0132799f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1464_n 0.00945407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1465_n 0.0132218f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1466_n 0.017651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1467_n 0.00449427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1468_n 0.0176342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1469_n 0.00526006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1470_n 0.0217289f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1471_n 0.00506466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1472_n 0.0164079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1473_n 0.029476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1474_n 0.0560743f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1475_n 0.0182786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1476_n 0.0475998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1477_n 0.0191114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1457_n 0.102779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1479_n 0.0048079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1480_n 0.00463502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1481_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1482_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1483_n 0.0128614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_304_463#_c_1599_n 0.00203976f $X=-0.19 $Y=1.655 $X2=0.592
+ $Y2=1.64
cc_239 VPB N_A_304_463#_c_1601_n 0.00172661f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_304_463#_c_1602_n 0.0126702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB Q 0.00133701f $X=-0.19 $Y=1.655 $X2=0.592 $Y2=1.805
cc_242 VPB Q_N 0.00882992f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_243 VPB Q_N 0.0121582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB Q_N 0.0452598f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 CLK N_A_197_108#_c_331_n 0.0425329f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_246 N_CLK_c_248_n N_A_197_108#_c_331_n 2.69717e-19 $X=0.615 $Y=1.805 $X2=0
+ $Y2=0
cc_247 N_CLK_M1012_g N_A_197_108#_c_352_n 3.9525e-19 $X=0.48 $Y=2.68 $X2=0 $Y2=0
cc_248 N_CLK_M1027_g N_A_28_108#_M1014_g 0.0104606f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_249 N_CLK_M1027_g N_A_28_108#_c_930_n 0.00576321f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_250 N_CLK_M1012_g N_A_28_108#_c_930_n 0.0031545f $X=0.48 $Y=2.68 $X2=0 $Y2=0
cc_251 CLK N_A_28_108#_c_930_n 0.00422718f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_252 N_CLK_c_248_n N_A_28_108#_c_930_n 0.019325f $X=0.615 $Y=1.805 $X2=0 $Y2=0
cc_253 N_CLK_M1012_g N_A_28_108#_c_947_n 0.0157729f $X=0.48 $Y=2.68 $X2=0 $Y2=0
cc_254 CLK N_A_28_108#_c_947_n 0.00615732f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_255 N_CLK_M1027_g N_A_28_108#_c_933_n 0.00917402f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_256 N_CLK_M1027_g N_A_28_108#_c_934_n 0.0300419f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_257 CLK N_A_28_108#_c_934_n 0.0470522f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_258 N_CLK_M1027_g N_A_28_108#_c_935_n 0.0176028f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_259 CLK N_A_28_108#_c_935_n 0.0313842f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_260 N_CLK_c_248_n N_A_28_108#_c_935_n 0.00133533f $X=0.615 $Y=1.805 $X2=0
+ $Y2=0
cc_261 N_CLK_M1027_g N_A_28_108#_c_936_n 0.0213485f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_262 CLK N_A_28_108#_c_936_n 0.00349388f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_263 N_CLK_c_248_n N_A_28_108#_c_936_n 7.91557e-19 $X=0.615 $Y=1.805 $X2=0
+ $Y2=0
cc_264 N_CLK_M1027_g N_A_28_108#_c_937_n 0.00874187f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_265 N_CLK_M1012_g N_VPWR_c_1458_n 0.0133671f $X=0.48 $Y=2.68 $X2=0 $Y2=0
cc_266 CLK N_VPWR_c_1458_n 0.030015f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_267 N_CLK_c_248_n N_VPWR_c_1458_n 0.00110114f $X=0.615 $Y=1.805 $X2=0 $Y2=0
cc_268 N_CLK_M1012_g N_VPWR_c_1472_n 0.00411131f $X=0.48 $Y=2.68 $X2=0 $Y2=0
cc_269 N_CLK_M1012_g N_VPWR_c_1457_n 0.00816709f $X=0.48 $Y=2.68 $X2=0 $Y2=0
cc_270 N_CLK_M1027_g N_VGND_c_1703_n 0.0032504f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_271 N_CLK_M1027_g N_VGND_c_1711_n 0.00445346f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_272 N_CLK_M1027_g N_VGND_c_1717_n 0.00493565f $X=0.48 $Y=0.75 $X2=0 $Y2=0
cc_273 D N_A_197_108#_c_333_n 0.00114263f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_274 N_D_c_280_n N_A_197_108#_c_334_n 0.00201794f $X=2.49 $Y=1.485 $X2=0 $Y2=0
cc_275 D N_A_197_108#_c_334_n 0.00684317f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_276 D N_A_197_108#_c_339_n 0.00669563f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_277 N_D_c_280_n N_A_197_108#_c_340_n 0.00406294f $X=2.49 $Y=1.485 $X2=0 $Y2=0
cc_278 D N_A_197_108#_c_340_n 0.0127505f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_279 N_D_M1013_g N_RESET_B_M1025_g 0.0185316f $X=2.43 $Y=2.525 $X2=0 $Y2=0
cc_280 N_D_c_280_n N_RESET_B_M1000_g 0.0246294f $X=2.49 $Y=1.485 $X2=0 $Y2=0
cc_281 D N_RESET_B_M1000_g 0.00999707f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_282 N_D_c_280_n N_RESET_B_c_629_n 0.00881753f $X=2.49 $Y=1.485 $X2=0 $Y2=0
cc_283 D N_RESET_B_c_633_n 0.00665232f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_284 N_D_c_283_n N_RESET_B_c_633_n 0.0246294f $X=2.49 $Y=1.65 $X2=0 $Y2=0
cc_285 N_D_c_281_n N_RESET_B_c_641_n 0.00741205f $X=2.49 $Y=1.99 $X2=0 $Y2=0
cc_286 N_D_c_281_n N_RESET_B_c_642_n 0.00309776f $X=2.49 $Y=1.99 $X2=0 $Y2=0
cc_287 N_D_c_286_n N_RESET_B_c_642_n 0.0012229f $X=2.49 $Y=2.155 $X2=0 $Y2=0
cc_288 D N_RESET_B_c_642_n 0.0444737f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_289 D N_RESET_B_c_643_n 6.81234e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_290 D N_RESET_B_c_634_n 0.00463703f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_291 N_D_c_283_n N_RESET_B_c_634_n 0.00741205f $X=2.49 $Y=1.65 $X2=0 $Y2=0
cc_292 D N_RESET_B_c_635_n 0.0543685f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_293 N_D_c_283_n N_RESET_B_c_635_n 5.11581e-19 $X=2.49 $Y=1.65 $X2=0 $Y2=0
cc_294 N_D_M1013_g N_A_28_108#_c_939_n 0.0100449f $X=2.43 $Y=2.525 $X2=0 $Y2=0
cc_295 N_D_M1013_g N_A_28_108#_M1003_g 0.016434f $X=2.43 $Y=2.525 $X2=0 $Y2=0
cc_296 N_D_c_280_n N_A_28_108#_M1003_g 0.0122459f $X=2.49 $Y=1.485 $X2=0 $Y2=0
cc_297 D N_A_28_108#_M1003_g 9.91214e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_298 N_D_c_283_n N_A_28_108#_M1003_g 0.042099f $X=2.49 $Y=1.65 $X2=0 $Y2=0
cc_299 N_D_M1013_g N_VPWR_c_1459_n 0.00430022f $X=2.43 $Y=2.525 $X2=0 $Y2=0
cc_300 N_D_M1013_g N_VPWR_c_1457_n 9.39239e-19 $X=2.43 $Y=2.525 $X2=0 $Y2=0
cc_301 N_D_M1013_g N_A_304_463#_c_1603_n 0.00847642f $X=2.43 $Y=2.525 $X2=0
+ $Y2=0
cc_302 D N_A_304_463#_c_1603_n 0.0351743f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_303 N_D_c_280_n N_A_304_463#_c_1599_n 0.0015814f $X=2.49 $Y=1.485 $X2=0 $Y2=0
cc_304 D N_A_304_463#_c_1599_n 0.0567295f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_305 N_D_c_283_n N_A_304_463#_c_1599_n 0.00371532f $X=2.49 $Y=1.65 $X2=0 $Y2=0
cc_306 D N_A_304_463#_c_1608_n 0.00585036f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_307 N_D_c_283_n N_A_304_463#_c_1608_n 0.00348504f $X=2.49 $Y=1.65 $X2=0 $Y2=0
cc_308 N_D_M1013_g N_A_304_463#_c_1602_n 0.00394045f $X=2.43 $Y=2.525 $X2=0
+ $Y2=0
cc_309 N_D_c_286_n N_A_304_463#_c_1602_n 0.00407922f $X=2.49 $Y=2.155 $X2=0
+ $Y2=0
cc_310 D N_A_304_463#_c_1602_n 0.00515405f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_311 D A_423_191# 0.00105575f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_312 N_A_197_108#_c_337_n N_A_804_328#_M1020_d 0.00433831f $X=6.27 $Y=0.805
+ $X2=-0.19 $Y2=-0.245
cc_313 N_A_197_108#_c_327_n N_A_804_328#_M1010_g 4.07574e-19 $X=3.44 $Y=1.945
+ $X2=0 $Y2=0
cc_314 N_A_197_108#_c_328_n N_A_804_328#_M1010_g 0.0357342f $X=3.735 $Y=1.45
+ $X2=0 $Y2=0
cc_315 N_A_197_108#_c_336_n N_A_804_328#_M1010_g 0.00244906f $X=4.54 $Y=0.715
+ $X2=0 $Y2=0
cc_316 N_A_197_108#_M1018_g N_A_804_328#_M1009_g 0.00300256f $X=3.44 $Y=2.525
+ $X2=0 $Y2=0
cc_317 N_A_197_108#_c_327_n N_A_804_328#_c_521_n 0.00601212f $X=3.44 $Y=1.945
+ $X2=0 $Y2=0
cc_318 N_A_197_108#_M1018_g N_A_804_328#_c_521_n 4.31082e-19 $X=3.44 $Y=2.525
+ $X2=0 $Y2=0
cc_319 N_A_197_108#_c_328_n N_A_804_328#_c_523_n 6.13034e-19 $X=3.735 $Y=1.45
+ $X2=0 $Y2=0
cc_320 N_A_197_108#_c_329_n N_A_804_328#_c_525_n 0.00122536f $X=6.15 $Y=1.39
+ $X2=0 $Y2=0
cc_321 N_A_197_108#_c_343_n N_A_804_328#_c_525_n 0.00818838f $X=6.53 $Y=1.555
+ $X2=0 $Y2=0
cc_322 N_A_197_108#_c_329_n N_A_804_328#_c_526_n 0.00356187f $X=6.15 $Y=1.39
+ $X2=0 $Y2=0
cc_323 N_A_197_108#_c_337_n N_A_804_328#_c_526_n 0.0164806f $X=6.27 $Y=0.805
+ $X2=0 $Y2=0
cc_324 N_A_197_108#_c_338_n N_A_804_328#_c_526_n 0.0386635f $X=6.365 $Y=1.555
+ $X2=0 $Y2=0
cc_325 N_A_197_108#_c_343_n N_A_804_328#_c_548_n 0.00215396f $X=6.53 $Y=1.555
+ $X2=0 $Y2=0
cc_326 N_A_197_108#_c_348_n N_RESET_B_M1025_g 0.00266628f $X=1.19 $Y=2.51 $X2=0
+ $Y2=0
cc_327 N_A_197_108#_c_352_n N_RESET_B_M1025_g 0.00334426f $X=1.19 $Y=2.35 $X2=0
+ $Y2=0
cc_328 N_A_197_108#_c_332_n N_RESET_B_M1000_g 0.00272505f $X=1.3 $Y=1.04 $X2=0
+ $Y2=0
cc_329 N_A_197_108#_c_333_n N_RESET_B_M1000_g 0.010305f $X=2.045 $Y=0.955 $X2=0
+ $Y2=0
cc_330 N_A_197_108#_c_334_n N_RESET_B_M1000_g 9.38622e-19 $X=3.095 $Y=0.715
+ $X2=0 $Y2=0
cc_331 N_A_197_108#_c_339_n N_RESET_B_M1000_g 0.00744497f $X=1.252 $Y=1.58 $X2=0
+ $Y2=0
cc_332 N_A_197_108#_c_340_n N_RESET_B_M1000_g 0.0134597f $X=2.15 $Y=0.715 $X2=0
+ $Y2=0
cc_333 N_A_197_108#_c_328_n N_RESET_B_c_629_n 0.00881753f $X=3.735 $Y=1.45 $X2=0
+ $Y2=0
cc_334 N_A_197_108#_c_334_n N_RESET_B_c_629_n 0.0187279f $X=3.095 $Y=0.715 $X2=0
+ $Y2=0
cc_335 N_A_197_108#_c_336_n N_RESET_B_c_629_n 0.0290173f $X=4.54 $Y=0.715 $X2=0
+ $Y2=0
cc_336 N_A_197_108#_c_340_n N_RESET_B_c_629_n 0.00147306f $X=2.15 $Y=0.715 $X2=0
+ $Y2=0
cc_337 N_A_197_108#_c_341_n N_RESET_B_c_629_n 0.0053441f $X=3.18 $Y=0.715 $X2=0
+ $Y2=0
cc_338 N_A_197_108#_c_336_n N_RESET_B_M1026_g 0.0174015f $X=4.54 $Y=0.715 $X2=0
+ $Y2=0
cc_339 N_A_197_108#_c_337_n N_RESET_B_M1026_g 0.00167209f $X=6.27 $Y=0.805 $X2=0
+ $Y2=0
cc_340 N_A_197_108#_c_333_n N_RESET_B_c_633_n 0.00375722f $X=2.045 $Y=0.955
+ $X2=0 $Y2=0
cc_341 N_A_197_108#_c_339_n N_RESET_B_c_633_n 7.8527e-19 $X=1.252 $Y=1.58 $X2=0
+ $Y2=0
cc_342 N_A_197_108#_c_350_n N_RESET_B_c_641_n 7.8527e-19 $X=1.252 $Y=1.958 $X2=0
+ $Y2=0
cc_343 N_A_197_108#_c_352_n N_RESET_B_c_641_n 2.09777e-19 $X=1.19 $Y=2.35 $X2=0
+ $Y2=0
cc_344 N_A_197_108#_c_327_n N_RESET_B_c_642_n 0.00737392f $X=3.44 $Y=1.945 $X2=0
+ $Y2=0
cc_345 N_A_197_108#_M1018_g N_RESET_B_c_642_n 0.0112828f $X=3.44 $Y=2.525 $X2=0
+ $Y2=0
cc_346 N_A_197_108#_c_342_n N_RESET_B_c_642_n 0.0159879f $X=3.405 $Y=1.78 $X2=0
+ $Y2=0
cc_347 N_A_197_108#_c_350_n N_RESET_B_c_643_n 0.00612529f $X=1.252 $Y=1.958
+ $X2=0 $Y2=0
cc_348 N_A_197_108#_c_352_n N_RESET_B_c_643_n 0.00149644f $X=1.19 $Y=2.35 $X2=0
+ $Y2=0
cc_349 N_A_197_108#_M1002_g N_RESET_B_c_644_n 0.0102691f $X=6.915 $Y=2.57 $X2=0
+ $Y2=0
cc_350 N_A_197_108#_c_338_n N_RESET_B_c_644_n 0.00749067f $X=6.365 $Y=1.555
+ $X2=0 $Y2=0
cc_351 N_A_197_108#_c_343_n N_RESET_B_c_644_n 0.00704629f $X=6.53 $Y=1.555 $X2=0
+ $Y2=0
cc_352 N_A_197_108#_c_331_n N_RESET_B_c_634_n 7.8527e-19 $X=1.252 $Y=1.722 $X2=0
+ $Y2=0
cc_353 N_A_197_108#_c_333_n N_RESET_B_c_635_n 0.0117024f $X=2.045 $Y=0.955 $X2=0
+ $Y2=0
cc_354 N_A_197_108#_c_352_n N_RESET_B_c_635_n 0.0026035f $X=1.19 $Y=2.35 $X2=0
+ $Y2=0
cc_355 N_A_197_108#_c_339_n N_RESET_B_c_635_n 0.0439368f $X=1.252 $Y=1.58 $X2=0
+ $Y2=0
cc_356 N_A_197_108#_c_335_n N_A_603_191#_M1003_d 0.0104839f $X=3.18 $Y=1.615
+ $X2=-0.19 $Y2=-0.245
cc_357 N_A_197_108#_c_329_n N_A_603_191#_c_827_n 0.0259894f $X=6.15 $Y=1.39
+ $X2=0 $Y2=0
cc_358 N_A_197_108#_c_337_n N_A_603_191#_c_827_n 0.0170041f $X=6.27 $Y=0.805
+ $X2=0 $Y2=0
cc_359 N_A_197_108#_c_327_n N_A_603_191#_c_828_n 0.0125906f $X=3.44 $Y=1.945
+ $X2=0 $Y2=0
cc_360 N_A_197_108#_M1018_g N_A_603_191#_c_828_n 0.00536835f $X=3.44 $Y=2.525
+ $X2=0 $Y2=0
cc_361 N_A_197_108#_c_328_n N_A_603_191#_c_828_n 0.00494252f $X=3.735 $Y=1.45
+ $X2=0 $Y2=0
cc_362 N_A_197_108#_c_335_n N_A_603_191#_c_828_n 0.0108796f $X=3.18 $Y=1.615
+ $X2=0 $Y2=0
cc_363 N_A_197_108#_c_342_n N_A_603_191#_c_828_n 0.024198f $X=3.405 $Y=1.78
+ $X2=0 $Y2=0
cc_364 N_A_197_108#_M1018_g N_A_603_191#_c_834_n 5.74657e-19 $X=3.44 $Y=2.525
+ $X2=0 $Y2=0
cc_365 N_A_197_108#_c_336_n N_A_603_191#_c_846_n 0.0285421f $X=4.54 $Y=0.715
+ $X2=0 $Y2=0
cc_366 N_A_197_108#_c_337_n N_A_603_191#_c_846_n 0.0621646f $X=6.27 $Y=0.805
+ $X2=0 $Y2=0
cc_367 N_A_197_108#_c_343_n N_A_603_191#_c_829_n 2.6234e-19 $X=6.53 $Y=1.555
+ $X2=0 $Y2=0
cc_368 N_A_197_108#_c_327_n N_A_603_191#_c_849_n 0.007238f $X=3.44 $Y=1.945
+ $X2=0 $Y2=0
cc_369 N_A_197_108#_c_328_n N_A_603_191#_c_849_n 0.0106639f $X=3.735 $Y=1.45
+ $X2=0 $Y2=0
cc_370 N_A_197_108#_c_335_n N_A_603_191#_c_849_n 0.0265677f $X=3.18 $Y=1.615
+ $X2=0 $Y2=0
cc_371 N_A_197_108#_c_336_n N_A_603_191#_c_849_n 0.0528169f $X=4.54 $Y=0.715
+ $X2=0 $Y2=0
cc_372 N_A_197_108#_c_342_n N_A_603_191#_c_849_n 0.00314451f $X=3.405 $Y=1.78
+ $X2=0 $Y2=0
cc_373 N_A_197_108#_c_337_n N_A_603_191#_c_830_n 7.37384e-19 $X=6.27 $Y=0.805
+ $X2=0 $Y2=0
cc_374 N_A_197_108#_c_343_n N_A_603_191#_c_830_n 0.015211f $X=6.53 $Y=1.555
+ $X2=0 $Y2=0
cc_375 N_A_197_108#_c_332_n N_A_28_108#_M1014_g 0.00749509f $X=1.3 $Y=1.04 $X2=0
+ $Y2=0
cc_376 N_A_197_108#_c_339_n N_A_28_108#_M1014_g 9.53246e-19 $X=1.252 $Y=1.58
+ $X2=0 $Y2=0
cc_377 N_A_197_108#_c_348_n N_A_28_108#_M1028_g 6.7294e-19 $X=1.19 $Y=2.51 $X2=0
+ $Y2=0
cc_378 N_A_197_108#_c_352_n N_A_28_108#_M1028_g 0.0023971f $X=1.19 $Y=2.35 $X2=0
+ $Y2=0
cc_379 N_A_197_108#_c_329_n N_A_28_108#_c_928_n 0.00788265f $X=6.15 $Y=1.39
+ $X2=0 $Y2=0
cc_380 N_A_197_108#_c_332_n N_A_28_108#_c_928_n 0.00643416f $X=1.3 $Y=1.04 $X2=0
+ $Y2=0
cc_381 N_A_197_108#_c_333_n N_A_28_108#_c_928_n 0.00640947f $X=2.045 $Y=0.955
+ $X2=0 $Y2=0
cc_382 N_A_197_108#_c_336_n N_A_28_108#_c_928_n 0.0038404f $X=4.54 $Y=0.715
+ $X2=0 $Y2=0
cc_383 N_A_197_108#_c_337_n N_A_28_108#_c_928_n 0.0183871f $X=6.27 $Y=0.805
+ $X2=0 $Y2=0
cc_384 N_A_197_108#_c_340_n N_A_28_108#_c_928_n 8.87392e-19 $X=2.15 $Y=0.715
+ $X2=0 $Y2=0
cc_385 N_A_197_108#_c_349_n N_A_28_108#_c_939_n 0.0066165f $X=1.125 $Y=2.515
+ $X2=0 $Y2=0
cc_386 N_A_197_108#_c_331_n N_A_28_108#_c_930_n 0.00422718f $X=1.252 $Y=1.722
+ $X2=0 $Y2=0
cc_387 N_A_197_108#_c_350_n N_A_28_108#_c_930_n 0.0056781f $X=1.252 $Y=1.958
+ $X2=0 $Y2=0
cc_388 N_A_197_108#_c_352_n N_A_28_108#_c_930_n 4.282e-19 $X=1.19 $Y=2.35 $X2=0
+ $Y2=0
cc_389 N_A_197_108#_c_353_n N_A_28_108#_c_930_n 0.00349711f $X=1.252 $Y=2.1
+ $X2=0 $Y2=0
cc_390 N_A_197_108#_c_327_n N_A_28_108#_M1003_g 0.0265682f $X=3.44 $Y=1.945
+ $X2=0 $Y2=0
cc_391 N_A_197_108#_M1018_g N_A_28_108#_M1003_g 0.0252709f $X=3.44 $Y=2.525
+ $X2=0 $Y2=0
cc_392 N_A_197_108#_c_328_n N_A_28_108#_M1003_g 0.00438269f $X=3.735 $Y=1.45
+ $X2=0 $Y2=0
cc_393 N_A_197_108#_c_334_n N_A_28_108#_M1003_g 0.00275942f $X=3.095 $Y=0.715
+ $X2=0 $Y2=0
cc_394 N_A_197_108#_c_335_n N_A_28_108#_M1003_g 0.0101791f $X=3.18 $Y=1.615
+ $X2=0 $Y2=0
cc_395 N_A_197_108#_c_342_n N_A_28_108#_M1003_g 0.00213363f $X=3.405 $Y=1.78
+ $X2=0 $Y2=0
cc_396 N_A_197_108#_M1018_g N_A_28_108#_c_943_n 0.0104164f $X=3.44 $Y=2.525
+ $X2=0 $Y2=0
cc_397 N_A_197_108#_c_327_n N_A_28_108#_M1011_g 2.29185e-19 $X=3.44 $Y=1.945
+ $X2=0 $Y2=0
cc_398 N_A_197_108#_M1018_g N_A_28_108#_M1011_g 0.0131134f $X=3.44 $Y=2.525
+ $X2=0 $Y2=0
cc_399 N_A_197_108#_M1002_g N_A_28_108#_M1029_g 0.015997f $X=6.915 $Y=2.57 $X2=0
+ $Y2=0
cc_400 N_A_197_108#_c_338_n N_A_28_108#_M1029_g 0.00102182f $X=6.365 $Y=1.555
+ $X2=0 $Y2=0
cc_401 N_A_197_108#_c_343_n N_A_28_108#_M1029_g 0.01018f $X=6.53 $Y=1.555 $X2=0
+ $Y2=0
cc_402 N_A_197_108#_c_330_n N_A_28_108#_M1005_g 0.00114155f $X=6.84 $Y=1.645
+ $X2=0 $Y2=0
cc_403 N_A_197_108#_c_348_n N_A_28_108#_c_947_n 0.00425104f $X=1.19 $Y=2.51
+ $X2=0 $Y2=0
cc_404 N_A_197_108#_c_352_n N_A_28_108#_c_947_n 0.00626068f $X=1.19 $Y=2.35
+ $X2=0 $Y2=0
cc_405 N_A_197_108#_c_332_n N_A_28_108#_c_935_n 0.00222341f $X=1.3 $Y=1.04 $X2=0
+ $Y2=0
cc_406 N_A_197_108#_c_339_n N_A_28_108#_c_935_n 0.0264207f $X=1.252 $Y=1.58
+ $X2=0 $Y2=0
cc_407 N_A_197_108#_c_332_n N_A_28_108#_c_936_n 0.0053534f $X=1.3 $Y=1.04 $X2=0
+ $Y2=0
cc_408 N_A_197_108#_c_339_n N_A_28_108#_c_936_n 0.0144255f $X=1.252 $Y=1.58
+ $X2=0 $Y2=0
cc_409 N_A_197_108#_M1002_g N_A_1440_304#_c_1087_n 0.0408174f $X=6.915 $Y=2.57
+ $X2=0 $Y2=0
cc_410 N_A_197_108#_c_330_n N_A_1440_304#_c_1081_n 7.04468e-19 $X=6.84 $Y=1.645
+ $X2=0 $Y2=0
cc_411 N_A_197_108#_M1002_g N_A_1440_304#_c_1081_n 0.00154361f $X=6.915 $Y=2.57
+ $X2=0 $Y2=0
cc_412 N_A_197_108#_c_330_n N_A_1440_304#_c_1082_n 0.0408174f $X=6.84 $Y=1.645
+ $X2=0 $Y2=0
cc_413 N_A_197_108#_c_343_n N_A_1440_304#_c_1082_n 5.64085e-19 $X=6.53 $Y=1.555
+ $X2=0 $Y2=0
cc_414 N_A_197_108#_c_337_n N_A_1245_128#_M1021_d 0.00483246f $X=6.27 $Y=0.805
+ $X2=-0.19 $Y2=-0.245
cc_415 N_A_197_108#_c_338_n N_A_1245_128#_M1021_d 0.00552282f $X=6.365 $Y=1.555
+ $X2=-0.19 $Y2=-0.245
cc_416 N_A_197_108#_c_343_n N_A_1245_128#_c_1205_n 0.00327665f $X=6.53 $Y=1.555
+ $X2=0 $Y2=0
cc_417 N_A_197_108#_c_329_n N_A_1245_128#_c_1178_n 0.00376224f $X=6.15 $Y=1.39
+ $X2=0 $Y2=0
cc_418 N_A_197_108#_c_337_n N_A_1245_128#_c_1178_n 0.0139839f $X=6.27 $Y=0.805
+ $X2=0 $Y2=0
cc_419 N_A_197_108#_c_338_n N_A_1245_128#_c_1178_n 0.0265092f $X=6.365 $Y=1.555
+ $X2=0 $Y2=0
cc_420 N_A_197_108#_c_330_n N_A_1245_128#_c_1179_n 0.00640978f $X=6.84 $Y=1.645
+ $X2=0 $Y2=0
cc_421 N_A_197_108#_c_330_n N_A_1245_128#_c_1189_n 0.0164635f $X=6.84 $Y=1.645
+ $X2=0 $Y2=0
cc_422 N_A_197_108#_M1002_g N_A_1245_128#_c_1189_n 0.0177792f $X=6.915 $Y=2.57
+ $X2=0 $Y2=0
cc_423 N_A_197_108#_c_338_n N_A_1245_128#_c_1189_n 0.0204881f $X=6.365 $Y=1.555
+ $X2=0 $Y2=0
cc_424 N_A_197_108#_c_343_n N_A_1245_128#_c_1189_n 0.00302632f $X=6.53 $Y=1.555
+ $X2=0 $Y2=0
cc_425 N_A_197_108#_c_338_n N_A_1245_128#_c_1190_n 0.0150159f $X=6.365 $Y=1.555
+ $X2=0 $Y2=0
cc_426 N_A_197_108#_c_343_n N_A_1245_128#_c_1190_n 0.00109421f $X=6.53 $Y=1.555
+ $X2=0 $Y2=0
cc_427 N_A_197_108#_c_348_n N_VPWR_c_1458_n 0.0262995f $X=1.19 $Y=2.51 $X2=0
+ $Y2=0
cc_428 N_A_197_108#_c_349_n N_VPWR_c_1459_n 0.00959822f $X=1.125 $Y=2.515 $X2=0
+ $Y2=0
cc_429 N_A_197_108#_M1002_g N_VPWR_c_1462_n 0.00140117f $X=6.915 $Y=2.57 $X2=0
+ $Y2=0
cc_430 N_A_197_108#_c_349_n N_VPWR_c_1473_n 0.0168758f $X=1.125 $Y=2.515 $X2=0
+ $Y2=0
cc_431 N_A_197_108#_M1002_g N_VPWR_c_1476_n 0.00457115f $X=6.915 $Y=2.57 $X2=0
+ $Y2=0
cc_432 N_A_197_108#_M1018_g N_VPWR_c_1457_n 9.39239e-19 $X=3.44 $Y=2.525 $X2=0
+ $Y2=0
cc_433 N_A_197_108#_M1002_g N_VPWR_c_1457_n 0.00490658f $X=6.915 $Y=2.57 $X2=0
+ $Y2=0
cc_434 N_A_197_108#_c_349_n N_VPWR_c_1457_n 0.0107452f $X=1.125 $Y=2.515 $X2=0
+ $Y2=0
cc_435 N_A_197_108#_c_327_n N_A_304_463#_c_1599_n 4.13985e-19 $X=3.44 $Y=1.945
+ $X2=0 $Y2=0
cc_436 N_A_197_108#_M1018_g N_A_304_463#_c_1599_n 0.00115052f $X=3.44 $Y=2.525
+ $X2=0 $Y2=0
cc_437 N_A_197_108#_c_335_n N_A_304_463#_c_1599_n 0.0280455f $X=3.18 $Y=1.615
+ $X2=0 $Y2=0
cc_438 N_A_197_108#_c_342_n N_A_304_463#_c_1599_n 0.0253146f $X=3.405 $Y=1.78
+ $X2=0 $Y2=0
cc_439 N_A_197_108#_c_352_n N_A_304_463#_c_1601_n 0.0322342f $X=1.19 $Y=2.35
+ $X2=0 $Y2=0
cc_440 N_A_197_108#_c_334_n N_A_304_463#_c_1608_n 0.0280398f $X=3.095 $Y=0.715
+ $X2=0 $Y2=0
cc_441 N_A_197_108#_c_335_n N_A_304_463#_c_1608_n 0.0180638f $X=3.18 $Y=1.615
+ $X2=0 $Y2=0
cc_442 N_A_197_108#_c_327_n N_A_304_463#_c_1602_n 0.00230862f $X=3.44 $Y=1.945
+ $X2=0 $Y2=0
cc_443 N_A_197_108#_M1018_g N_A_304_463#_c_1602_n 0.00226731f $X=3.44 $Y=2.525
+ $X2=0 $Y2=0
cc_444 N_A_197_108#_c_342_n N_A_304_463#_c_1602_n 0.00890159f $X=3.405 $Y=1.78
+ $X2=0 $Y2=0
cc_445 N_A_197_108#_c_333_n N_VGND_M1000_s 0.0103358f $X=2.045 $Y=0.955 $X2=0
+ $Y2=0
cc_446 N_A_197_108#_c_337_n N_VGND_M1026_d 0.0141895f $X=6.27 $Y=0.805 $X2=0
+ $Y2=0
cc_447 N_A_197_108#_c_332_n N_VGND_c_1704_n 0.00975225f $X=1.3 $Y=1.04 $X2=0
+ $Y2=0
cc_448 N_A_197_108#_c_333_n N_VGND_c_1704_n 0.0268035f $X=2.045 $Y=0.955 $X2=0
+ $Y2=0
cc_449 N_A_197_108#_c_340_n N_VGND_c_1704_n 0.00536328f $X=2.15 $Y=0.715 $X2=0
+ $Y2=0
cc_450 N_A_197_108#_c_337_n N_VGND_c_1705_n 0.025714f $X=6.27 $Y=0.805 $X2=0
+ $Y2=0
cc_451 N_A_197_108#_c_337_n N_VGND_c_1709_n 0.0114527f $X=6.27 $Y=0.805 $X2=0
+ $Y2=0
cc_452 N_A_197_108#_c_332_n N_VGND_c_1712_n 0.00782093f $X=1.3 $Y=1.04 $X2=0
+ $Y2=0
cc_453 N_A_197_108#_c_334_n N_VGND_c_1713_n 0.0153767f $X=3.095 $Y=0.715 $X2=0
+ $Y2=0
cc_454 N_A_197_108#_c_336_n N_VGND_c_1713_n 0.0270999f $X=4.54 $Y=0.715 $X2=0
+ $Y2=0
cc_455 N_A_197_108#_c_337_n N_VGND_c_1713_n 0.00719708f $X=6.27 $Y=0.805 $X2=0
+ $Y2=0
cc_456 N_A_197_108#_c_340_n N_VGND_c_1713_n 0.00393693f $X=2.15 $Y=0.715 $X2=0
+ $Y2=0
cc_457 N_A_197_108#_c_341_n N_VGND_c_1713_n 0.00345508f $X=3.18 $Y=0.715 $X2=0
+ $Y2=0
cc_458 N_A_197_108#_c_329_n N_VGND_c_1717_n 9.54497e-19 $X=6.15 $Y=1.39 $X2=0
+ $Y2=0
cc_459 N_A_197_108#_c_332_n N_VGND_c_1717_n 0.0106024f $X=1.3 $Y=1.04 $X2=0
+ $Y2=0
cc_460 N_A_197_108#_c_334_n N_VGND_c_1717_n 0.0207833f $X=3.095 $Y=0.715 $X2=0
+ $Y2=0
cc_461 N_A_197_108#_c_336_n N_VGND_c_1717_n 0.0367639f $X=4.54 $Y=0.715 $X2=0
+ $Y2=0
cc_462 N_A_197_108#_c_337_n N_VGND_c_1717_n 0.032528f $X=6.27 $Y=0.805 $X2=0
+ $Y2=0
cc_463 N_A_197_108#_c_340_n N_VGND_c_1717_n 0.00529326f $X=2.15 $Y=0.715 $X2=0
+ $Y2=0
cc_464 N_A_197_108#_c_341_n N_VGND_c_1717_n 0.00450883f $X=3.18 $Y=0.715 $X2=0
+ $Y2=0
cc_465 N_A_197_108#_c_340_n A_423_191# 0.00173182f $X=2.15 $Y=0.715 $X2=-0.19
+ $Y2=-0.245
cc_466 N_A_804_328#_M1010_g N_RESET_B_c_629_n 0.00881753f $X=4.165 $Y=1.165
+ $X2=0 $Y2=0
cc_467 N_A_804_328#_M1010_g N_RESET_B_M1026_g 0.0324094f $X=4.165 $Y=1.165 $X2=0
+ $Y2=0
cc_468 N_A_804_328#_c_520_n N_RESET_B_M1026_g 0.00147578f $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_469 N_A_804_328#_c_521_n N_RESET_B_M1026_g 0.0209145f $X=4.185 $Y=1.805 $X2=0
+ $Y2=0
cc_470 N_A_804_328#_c_522_n N_RESET_B_M1026_g 0.0119116f $X=5.07 $Y=1.525 $X2=0
+ $Y2=0
cc_471 N_A_804_328#_c_524_n N_RESET_B_M1026_g 0.00400789f $X=5.155 $Y=1.9 $X2=0
+ $Y2=0
cc_472 N_A_804_328#_M1009_g N_RESET_B_M1015_g 0.0212826f $X=4.23 $Y=2.525 $X2=0
+ $Y2=0
cc_473 N_A_804_328#_M1009_g N_RESET_B_c_642_n 0.00300379f $X=4.23 $Y=2.525 $X2=0
+ $Y2=0
cc_474 N_A_804_328#_c_520_n N_RESET_B_c_642_n 0.0173224f $X=4.185 $Y=1.805 $X2=0
+ $Y2=0
cc_475 N_A_804_328#_c_521_n N_RESET_B_c_642_n 0.00207391f $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_476 N_A_804_328#_c_522_n N_RESET_B_c_642_n 0.00431406f $X=5.07 $Y=1.525 $X2=0
+ $Y2=0
cc_477 N_A_804_328#_M1032_d N_RESET_B_c_644_n 0.0116193f $X=5.805 $Y=1.895 $X2=0
+ $Y2=0
cc_478 N_A_804_328#_c_522_n N_RESET_B_c_644_n 0.00717483f $X=5.07 $Y=1.525 $X2=0
+ $Y2=0
cc_479 N_A_804_328#_c_531_n N_RESET_B_c_644_n 0.0361186f $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_480 N_A_804_328#_c_532_n N_RESET_B_c_644_n 0.0144162f $X=5.24 $Y=1.985 $X2=0
+ $Y2=0
cc_481 N_A_804_328#_c_534_n N_RESET_B_c_644_n 0.013839f $X=6.04 $Y=2.745 $X2=0
+ $Y2=0
cc_482 N_A_804_328#_c_548_n N_RESET_B_c_644_n 0.0140294f $X=6.04 $Y=2.065 $X2=0
+ $Y2=0
cc_483 N_A_804_328#_M1009_g N_RESET_B_c_645_n 7.38414e-19 $X=4.23 $Y=2.525 $X2=0
+ $Y2=0
cc_484 N_A_804_328#_c_520_n N_RESET_B_c_645_n 0.00135705f $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_485 N_A_804_328#_c_521_n N_RESET_B_c_645_n 7.38429e-19 $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_486 N_A_804_328#_c_522_n N_RESET_B_c_645_n 0.00370171f $X=5.07 $Y=1.525 $X2=0
+ $Y2=0
cc_487 N_A_804_328#_c_532_n N_RESET_B_c_645_n 2.44103e-19 $X=5.24 $Y=1.985 $X2=0
+ $Y2=0
cc_488 N_A_804_328#_M1009_g N_RESET_B_c_648_n 0.00789243f $X=4.23 $Y=2.525 $X2=0
+ $Y2=0
cc_489 N_A_804_328#_c_520_n N_RESET_B_c_648_n 2.71604e-19 $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_490 N_A_804_328#_c_522_n N_RESET_B_c_648_n 0.0073991f $X=5.07 $Y=1.525 $X2=0
+ $Y2=0
cc_491 N_A_804_328#_c_524_n N_RESET_B_c_648_n 0.00139817f $X=5.155 $Y=1.9 $X2=0
+ $Y2=0
cc_492 N_A_804_328#_c_532_n N_RESET_B_c_648_n 0.00193902f $X=5.24 $Y=1.985 $X2=0
+ $Y2=0
cc_493 N_A_804_328#_M1009_g N_RESET_B_c_649_n 0.00101763f $X=4.23 $Y=2.525 $X2=0
+ $Y2=0
cc_494 N_A_804_328#_c_520_n N_RESET_B_c_649_n 0.0168504f $X=4.185 $Y=1.805 $X2=0
+ $Y2=0
cc_495 N_A_804_328#_c_521_n N_RESET_B_c_649_n 0.00111747f $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_496 N_A_804_328#_c_522_n N_RESET_B_c_649_n 0.0283076f $X=5.07 $Y=1.525 $X2=0
+ $Y2=0
cc_497 N_A_804_328#_c_524_n N_RESET_B_c_649_n 0.00835538f $X=5.155 $Y=1.9 $X2=0
+ $Y2=0
cc_498 N_A_804_328#_c_532_n N_RESET_B_c_649_n 0.0127666f $X=5.24 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_A_804_328#_c_525_n N_A_603_191#_c_827_n 5.41282e-19 $X=6.015 $Y=1.9
+ $X2=0 $Y2=0
cc_500 N_A_804_328#_c_526_n N_A_603_191#_c_827_n 0.00417094f $X=5.935 $Y=1.155
+ $X2=0 $Y2=0
cc_501 N_A_804_328#_c_524_n N_A_603_191#_M1032_g 0.00380112f $X=5.155 $Y=1.9
+ $X2=0 $Y2=0
cc_502 N_A_804_328#_c_531_n N_A_603_191#_M1032_g 0.0176376f $X=5.93 $Y=1.985
+ $X2=0 $Y2=0
cc_503 N_A_804_328#_c_534_n N_A_603_191#_M1032_g 0.0101559f $X=6.04 $Y=2.745
+ $X2=0 $Y2=0
cc_504 N_A_804_328#_M1010_g N_A_603_191#_c_828_n 0.0020553f $X=4.165 $Y=1.165
+ $X2=0 $Y2=0
cc_505 N_A_804_328#_M1009_g N_A_603_191#_c_828_n 0.00288413f $X=4.23 $Y=2.525
+ $X2=0 $Y2=0
cc_506 N_A_804_328#_c_520_n N_A_603_191#_c_828_n 0.0294923f $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_507 N_A_804_328#_c_521_n N_A_603_191#_c_828_n 0.00282041f $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_508 N_A_804_328#_c_523_n N_A_603_191#_c_828_n 0.0138373f $X=4.295 $Y=1.525
+ $X2=0 $Y2=0
cc_509 N_A_804_328#_c_521_n N_A_603_191#_c_866_n 5.43954e-19 $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_510 N_A_804_328#_M1009_g N_A_603_191#_c_833_n 0.0114126f $X=4.23 $Y=2.525
+ $X2=0 $Y2=0
cc_511 N_A_804_328#_c_520_n N_A_603_191#_c_833_n 0.0096138f $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_512 N_A_804_328#_c_521_n N_A_603_191#_c_833_n 0.00234116f $X=4.185 $Y=1.805
+ $X2=0 $Y2=0
cc_513 N_A_804_328#_c_532_n N_A_603_191#_c_833_n 0.00127506f $X=5.24 $Y=1.985
+ $X2=0 $Y2=0
cc_514 N_A_804_328#_M1010_g N_A_603_191#_c_846_n 0.00365977f $X=4.165 $Y=1.165
+ $X2=0 $Y2=0
cc_515 N_A_804_328#_c_522_n N_A_603_191#_c_846_n 0.0641347f $X=5.07 $Y=1.525
+ $X2=0 $Y2=0
cc_516 N_A_804_328#_c_531_n N_A_603_191#_c_846_n 0.00479835f $X=5.93 $Y=1.985
+ $X2=0 $Y2=0
cc_517 N_A_804_328#_c_522_n N_A_603_191#_c_829_n 0.0138148f $X=5.07 $Y=1.525
+ $X2=0 $Y2=0
cc_518 N_A_804_328#_c_524_n N_A_603_191#_c_829_n 0.00789367f $X=5.155 $Y=1.9
+ $X2=0 $Y2=0
cc_519 N_A_804_328#_c_531_n N_A_603_191#_c_829_n 0.0127445f $X=5.93 $Y=1.985
+ $X2=0 $Y2=0
cc_520 N_A_804_328#_c_525_n N_A_603_191#_c_829_n 0.0178407f $X=6.015 $Y=1.9
+ $X2=0 $Y2=0
cc_521 N_A_804_328#_c_526_n N_A_603_191#_c_829_n 0.00374369f $X=5.935 $Y=1.155
+ $X2=0 $Y2=0
cc_522 N_A_804_328#_M1010_g N_A_603_191#_c_879_n 0.0110153f $X=4.165 $Y=1.165
+ $X2=0 $Y2=0
cc_523 N_A_804_328#_c_523_n N_A_603_191#_c_879_n 0.0157236f $X=4.295 $Y=1.525
+ $X2=0 $Y2=0
cc_524 N_A_804_328#_c_522_n N_A_603_191#_c_830_n 0.00225529f $X=5.07 $Y=1.525
+ $X2=0 $Y2=0
cc_525 N_A_804_328#_c_524_n N_A_603_191#_c_830_n 0.00134653f $X=5.155 $Y=1.9
+ $X2=0 $Y2=0
cc_526 N_A_804_328#_c_531_n N_A_603_191#_c_830_n 0.00321696f $X=5.93 $Y=1.985
+ $X2=0 $Y2=0
cc_527 N_A_804_328#_c_525_n N_A_603_191#_c_830_n 0.00938041f $X=6.015 $Y=1.9
+ $X2=0 $Y2=0
cc_528 N_A_804_328#_c_526_n N_A_603_191#_c_830_n 3.54818e-19 $X=5.935 $Y=1.155
+ $X2=0 $Y2=0
cc_529 N_A_804_328#_M1009_g N_A_28_108#_M1011_g 0.0416336f $X=4.23 $Y=2.525
+ $X2=0 $Y2=0
cc_530 N_A_804_328#_M1009_g N_A_28_108#_c_945_n 0.0100709f $X=4.23 $Y=2.525
+ $X2=0 $Y2=0
cc_531 N_A_804_328#_c_534_n N_A_28_108#_c_945_n 0.00483184f $X=6.04 $Y=2.745
+ $X2=0 $Y2=0
cc_532 N_A_804_328#_c_534_n N_A_28_108#_M1029_g 0.00888318f $X=6.04 $Y=2.745
+ $X2=0 $Y2=0
cc_533 N_A_804_328#_c_548_n N_A_28_108#_M1029_g 0.00143143f $X=6.04 $Y=2.065
+ $X2=0 $Y2=0
cc_534 N_A_804_328#_c_534_n N_A_1245_128#_c_1205_n 0.0186837f $X=6.04 $Y=2.745
+ $X2=0 $Y2=0
cc_535 N_A_804_328#_c_548_n N_A_1245_128#_c_1205_n 9.06256e-19 $X=6.04 $Y=2.065
+ $X2=0 $Y2=0
cc_536 N_A_804_328#_c_525_n N_A_1245_128#_c_1189_n 0.0063049f $X=6.015 $Y=1.9
+ $X2=0 $Y2=0
cc_537 N_A_804_328#_c_548_n N_A_1245_128#_c_1189_n 0.00429906f $X=6.04 $Y=2.065
+ $X2=0 $Y2=0
cc_538 N_A_804_328#_c_531_n N_VPWR_M1032_s 0.00366342f $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_539 N_A_804_328#_M1009_g N_VPWR_c_1460_n 0.00429952f $X=4.23 $Y=2.525 $X2=0
+ $Y2=0
cc_540 N_A_804_328#_c_531_n N_VPWR_c_1461_n 0.0200875f $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_541 N_A_804_328#_c_534_n N_VPWR_c_1461_n 0.0376436f $X=6.04 $Y=2.745 $X2=0
+ $Y2=0
cc_542 N_A_804_328#_c_534_n N_VPWR_c_1476_n 0.00739966f $X=6.04 $Y=2.745 $X2=0
+ $Y2=0
cc_543 N_A_804_328#_M1009_g N_VPWR_c_1457_n 9.39239e-19 $X=4.23 $Y=2.525 $X2=0
+ $Y2=0
cc_544 N_A_804_328#_c_534_n N_VPWR_c_1457_n 0.00667223f $X=6.04 $Y=2.745 $X2=0
+ $Y2=0
cc_545 N_RESET_B_c_644_n N_A_603_191#_M1032_g 0.0061151f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_546 N_RESET_B_c_648_n N_A_603_191#_M1032_g 0.00407373f $X=4.805 $Y=1.955
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_642_n N_A_603_191#_c_828_n 0.0239787f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_548 N_RESET_B_c_645_n N_A_603_191#_c_828_n 0.00137304f $X=4.705 $Y=2.035
+ $X2=0 $Y2=0
cc_549 N_RESET_B_c_649_n N_A_603_191#_c_828_n 0.0015005f $X=4.805 $Y=1.955 $X2=0
+ $Y2=0
cc_550 N_RESET_B_M1015_g N_A_603_191#_c_833_n 0.014344f $X=4.78 $Y=2.525 $X2=0
+ $Y2=0
cc_551 N_RESET_B_c_642_n N_A_603_191#_c_833_n 0.0145661f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_552 N_RESET_B_c_644_n N_A_603_191#_c_833_n 0.0100818f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_645_n N_A_603_191#_c_833_n 0.00942075f $X=4.705 $Y=2.035
+ $X2=0 $Y2=0
cc_554 N_RESET_B_c_648_n N_A_603_191#_c_833_n 0.0065767f $X=4.805 $Y=1.955 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_649_n N_A_603_191#_c_833_n 0.0262231f $X=4.805 $Y=1.955 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_642_n N_A_603_191#_c_834_n 0.0121646f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_557 N_RESET_B_M1026_g N_A_603_191#_c_846_n 0.0143331f $X=4.635 $Y=1.165 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_644_n N_A_603_191#_c_829_n 0.00128557f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_559 N_RESET_B_M1026_g N_A_603_191#_c_879_n 5.1029e-19 $X=4.635 $Y=1.165 $X2=0
+ $Y2=0
cc_560 N_RESET_B_M1026_g N_A_603_191#_c_830_n 0.00464925f $X=4.635 $Y=1.165
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_630_n N_A_28_108#_c_928_n 0.161575f $X=2.115 $Y=0.54 $X2=0
+ $Y2=0
cc_562 N_RESET_B_M1025_g N_A_28_108#_c_939_n 0.0100449f $X=1.86 $Y=2.525 $X2=0
+ $Y2=0
cc_563 N_RESET_B_c_633_n N_A_28_108#_c_930_n 0.00705208f $X=2.04 $Y=1.56 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_635_n N_A_28_108#_c_930_n 0.00119066f $X=1.775 $Y=1.65 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_629_n N_A_28_108#_M1003_g 0.00881753f $X=4.56 $Y=0.54 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_642_n N_A_28_108#_M1003_g 0.00552326f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_642_n N_A_28_108#_M1011_g 0.00252676f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_568 N_RESET_B_M1015_g N_A_28_108#_c_945_n 0.0100824f $X=4.78 $Y=2.525 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_644_n N_A_28_108#_M1029_g 0.0101661f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_570 N_RESET_B_M1025_g N_A_28_108#_c_947_n 0.00153424f $X=1.86 $Y=2.525 $X2=0
+ $Y2=0
cc_571 N_RESET_B_c_634_n N_A_28_108#_c_947_n 0.00705208f $X=1.775 $Y=1.65 $X2=0
+ $Y2=0
cc_572 N_RESET_B_M1016_g N_A_1440_304#_M1001_g 0.0059701f $X=8.055 $Y=2.57 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_651_n N_A_1440_304#_M1001_g 2.72506e-19 $X=8.055 $Y=2.035
+ $X2=0 $Y2=0
cc_574 N_RESET_B_M1017_g N_A_1440_304#_M1033_g 0.0295409f $X=7.815 $Y=0.85 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_644_n N_A_1440_304#_c_1086_n 5.85404e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_576 N_RESET_B_c_650_n N_A_1440_304#_c_1086_n 8.50765e-19 $X=7.905 $Y=2.035
+ $X2=0 $Y2=0
cc_577 N_RESET_B_c_651_n N_A_1440_304#_c_1086_n 0.0220627f $X=8.055 $Y=2.035
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_644_n N_A_1440_304#_c_1087_n 7.93769e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_579 N_RESET_B_M1017_g N_A_1440_304#_c_1079_n 2.56934e-19 $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_580 N_RESET_B_M1017_g N_A_1440_304#_c_1081_n 0.00117449f $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_644_n N_A_1440_304#_c_1081_n 0.0231381f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_582 RESET_B N_A_1440_304#_c_1081_n 0.00130672f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_583 N_RESET_B_c_650_n N_A_1440_304#_c_1081_n 0.0137133f $X=7.905 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_651_n N_A_1440_304#_c_1081_n 4.12896e-19 $X=8.055 $Y=2.035
+ $X2=0 $Y2=0
cc_585 N_RESET_B_M1017_g N_A_1440_304#_c_1082_n 0.0220627f $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_586 N_RESET_B_M1016_g N_A_1440_304#_c_1090_n 4.40496e-19 $X=8.055 $Y=2.57
+ $X2=0 $Y2=0
cc_587 RESET_B N_A_1440_304#_c_1091_n 0.0012972f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_588 N_RESET_B_c_650_n N_A_1440_304#_c_1091_n 0.0152563f $X=7.905 $Y=2.035
+ $X2=0 $Y2=0
cc_589 N_RESET_B_c_651_n N_A_1440_304#_c_1091_n 0.00482257f $X=8.055 $Y=2.035
+ $X2=0 $Y2=0
cc_590 N_RESET_B_M1017_g N_A_1440_304#_c_1083_n 0.0109185f $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_591 N_RESET_B_c_644_n N_A_1440_304#_c_1083_n 0.00662159f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_592 RESET_B N_A_1440_304#_c_1083_n 0.00698294f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_593 N_RESET_B_c_650_n N_A_1440_304#_c_1083_n 0.0204735f $X=7.905 $Y=2.035
+ $X2=0 $Y2=0
cc_594 N_RESET_B_c_651_n N_A_1440_304#_c_1083_n 0.00688117f $X=8.055 $Y=2.035
+ $X2=0 $Y2=0
cc_595 N_RESET_B_M1017_g N_A_1440_304#_c_1084_n 0.00225081f $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_596 RESET_B N_A_1440_304#_c_1084_n 0.00127868f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_597 N_RESET_B_c_650_n N_A_1440_304#_c_1084_n 0.00198806f $X=7.905 $Y=2.035
+ $X2=0 $Y2=0
cc_598 N_RESET_B_c_651_n N_A_1440_304#_c_1084_n 0.00224579f $X=8.055 $Y=2.035
+ $X2=0 $Y2=0
cc_599 N_RESET_B_c_644_n N_A_1245_128#_M1029_d 0.00125515f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_600 N_RESET_B_M1017_g N_A_1245_128#_c_1173_n 0.0602547f $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_601 N_RESET_B_M1017_g N_A_1245_128#_M1006_g 0.00762272f $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_602 N_RESET_B_c_650_n N_A_1245_128#_M1006_g 2.32179e-19 $X=7.905 $Y=2.035
+ $X2=0 $Y2=0
cc_603 N_RESET_B_c_651_n N_A_1245_128#_M1006_g 0.0271766f $X=8.055 $Y=2.035
+ $X2=0 $Y2=0
cc_604 N_RESET_B_c_644_n N_A_1245_128#_c_1205_n 0.0243493f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_605 N_RESET_B_M1017_g N_A_1245_128#_c_1179_n 0.0121174f $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_606 N_RESET_B_c_644_n N_A_1245_128#_c_1179_n 0.0129123f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_RESET_B_M1017_g N_A_1245_128#_c_1180_n 0.0121205f $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_608 N_RESET_B_M1017_g N_A_1245_128#_c_1182_n 3.53007e-19 $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_609 N_RESET_B_c_644_n N_A_1245_128#_c_1189_n 0.00985101f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_610 N_RESET_B_M1017_g N_A_1245_128#_c_1191_n 0.00372605f $X=7.815 $Y=0.85
+ $X2=0 $Y2=0
cc_611 N_RESET_B_c_651_n N_A_1245_128#_c_1198_n 8.89759e-19 $X=8.055 $Y=2.035
+ $X2=0 $Y2=0
cc_612 N_RESET_B_c_644_n N_VPWR_M1032_s 0.00202f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_613 N_RESET_B_M1025_g N_VPWR_c_1459_n 0.00255809f $X=1.86 $Y=2.525 $X2=0
+ $Y2=0
cc_614 N_RESET_B_M1015_g N_VPWR_c_1460_n 0.00429952f $X=4.78 $Y=2.525 $X2=0
+ $Y2=0
cc_615 N_RESET_B_M1015_g N_VPWR_c_1461_n 0.00600604f $X=4.78 $Y=2.525 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_644_n N_VPWR_c_1461_n 0.00882035f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_617 N_RESET_B_M1016_g N_VPWR_c_1462_n 0.00961768f $X=8.055 $Y=2.57 $X2=0
+ $Y2=0
cc_618 N_RESET_B_c_644_n N_VPWR_c_1462_n 0.0078155f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_619 RESET_B N_VPWR_c_1462_n 0.00162874f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_620 N_RESET_B_c_650_n N_VPWR_c_1462_n 0.013972f $X=7.905 $Y=2.035 $X2=0 $Y2=0
cc_621 N_RESET_B_c_651_n N_VPWR_c_1462_n 0.00586827f $X=8.055 $Y=2.035 $X2=0
+ $Y2=0
cc_622 N_RESET_B_M1016_g N_VPWR_c_1466_n 0.00410383f $X=8.055 $Y=2.57 $X2=0
+ $Y2=0
cc_623 N_RESET_B_M1025_g N_VPWR_c_1457_n 9.39239e-19 $X=1.86 $Y=2.525 $X2=0
+ $Y2=0
cc_624 N_RESET_B_M1015_g N_VPWR_c_1457_n 9.39239e-19 $X=4.78 $Y=2.525 $X2=0
+ $Y2=0
cc_625 N_RESET_B_M1016_g N_VPWR_c_1457_n 0.00444863f $X=8.055 $Y=2.57 $X2=0
+ $Y2=0
cc_626 N_RESET_B_M1025_g N_A_304_463#_c_1603_n 0.0087158f $X=1.86 $Y=2.525 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_633_n N_A_304_463#_c_1603_n 0.00176715f $X=2.04 $Y=1.56 $X2=0
+ $Y2=0
cc_628 N_RESET_B_c_642_n N_A_304_463#_c_1603_n 0.0104099f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_629 N_RESET_B_c_643_n N_A_304_463#_c_1603_n 6.92429e-19 $X=1.825 $Y=2.035
+ $X2=0 $Y2=0
cc_630 N_RESET_B_c_635_n N_A_304_463#_c_1603_n 0.00750877f $X=1.775 $Y=1.65
+ $X2=0 $Y2=0
cc_631 N_RESET_B_c_642_n N_A_304_463#_c_1599_n 0.0257982f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_632 N_RESET_B_c_641_n N_A_304_463#_c_1601_n 8.85503e-19 $X=1.775 $Y=2.155
+ $X2=0 $Y2=0
cc_633 N_RESET_B_c_643_n N_A_304_463#_c_1601_n 0.00423535f $X=1.825 $Y=2.035
+ $X2=0 $Y2=0
cc_634 N_RESET_B_c_635_n N_A_304_463#_c_1601_n 0.0102278f $X=1.775 $Y=1.65 $X2=0
+ $Y2=0
cc_635 N_RESET_B_c_642_n N_A_304_463#_c_1602_n 0.0254977f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_636 N_RESET_B_c_630_n N_VGND_c_1704_n 0.00934919f $X=2.115 $Y=0.54 $X2=0
+ $Y2=0
cc_637 N_RESET_B_c_629_n N_VGND_c_1705_n 0.00262778f $X=4.56 $Y=0.54 $X2=0 $Y2=0
cc_638 N_RESET_B_M1017_g N_VGND_c_1706_n 9.5404e-19 $X=7.815 $Y=0.85 $X2=0 $Y2=0
cc_639 N_RESET_B_M1017_g N_VGND_c_1714_n 0.00372577f $X=7.815 $Y=0.85 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_630_n N_VGND_c_1717_n 0.0150436f $X=2.115 $Y=0.54 $X2=0 $Y2=0
cc_641 N_RESET_B_M1017_g N_VGND_c_1717_n 0.00418775f $X=7.815 $Y=0.85 $X2=0
+ $Y2=0
cc_642 N_A_603_191#_c_827_n N_A_28_108#_c_928_n 0.00788265f $X=5.72 $Y=1.39
+ $X2=0 $Y2=0
cc_643 N_A_603_191#_c_834_n N_A_28_108#_c_943_n 0.00337372f $X=3.965 $Y=2.385
+ $X2=0 $Y2=0
cc_644 N_A_603_191#_c_828_n N_A_28_108#_M1011_g 0.0044787f $X=3.77 $Y=2.3 $X2=0
+ $Y2=0
cc_645 N_A_603_191#_c_834_n N_A_28_108#_M1011_g 0.012949f $X=3.965 $Y=2.385
+ $X2=0 $Y2=0
cc_646 N_A_603_191#_M1032_g N_A_28_108#_c_945_n 0.0103107f $X=5.73 $Y=2.315
+ $X2=0 $Y2=0
cc_647 N_A_603_191#_c_833_n N_A_28_108#_c_945_n 0.00817682f $X=4.85 $Y=2.385
+ $X2=0 $Y2=0
cc_648 N_A_603_191#_M1032_g N_A_28_108#_M1029_g 0.0146248f $X=5.73 $Y=2.315
+ $X2=0 $Y2=0
cc_649 N_A_603_191#_c_833_n N_VPWR_M1009_d 0.00315285f $X=4.85 $Y=2.385 $X2=0
+ $Y2=0
cc_650 N_A_603_191#_c_833_n N_VPWR_c_1460_n 0.0207882f $X=4.85 $Y=2.385 $X2=0
+ $Y2=0
cc_651 N_A_603_191#_M1032_g N_VPWR_c_1461_n 0.0136231f $X=5.73 $Y=2.315 $X2=0
+ $Y2=0
cc_652 N_A_603_191#_c_833_n N_VPWR_c_1461_n 0.0260566f $X=4.85 $Y=2.385 $X2=0
+ $Y2=0
cc_653 N_A_603_191#_c_834_n N_VPWR_c_1474_n 0.0077644f $X=3.965 $Y=2.385 $X2=0
+ $Y2=0
cc_654 N_A_603_191#_c_833_n N_VPWR_c_1475_n 0.00441176f $X=4.85 $Y=2.385 $X2=0
+ $Y2=0
cc_655 N_A_603_191#_M1032_g N_VPWR_c_1457_n 7.88961e-19 $X=5.73 $Y=2.315 $X2=0
+ $Y2=0
cc_656 N_A_603_191#_c_833_n N_VPWR_c_1457_n 0.0233341f $X=4.85 $Y=2.385 $X2=0
+ $Y2=0
cc_657 N_A_603_191#_c_834_n N_VPWR_c_1457_n 0.0118674f $X=3.965 $Y=2.385 $X2=0
+ $Y2=0
cc_658 N_A_603_191#_c_828_n N_A_304_463#_c_1602_n 0.00673626f $X=3.77 $Y=2.3
+ $X2=0 $Y2=0
cc_659 N_A_603_191#_c_834_n N_A_304_463#_c_1602_n 0.00233325f $X=3.965 $Y=2.385
+ $X2=0 $Y2=0
cc_660 N_A_603_191#_c_833_n A_789_463# 0.00124295f $X=4.85 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_661 N_A_603_191#_c_846_n N_VGND_M1026_d 0.0234753f $X=5.41 $Y=1.16 $X2=0
+ $Y2=0
cc_662 N_A_603_191#_c_829_n N_VGND_M1026_d 7.34787e-19 $X=5.505 $Y=1.555 $X2=0
+ $Y2=0
cc_663 N_A_603_191#_c_827_n N_VGND_c_1705_n 0.00161872f $X=5.72 $Y=1.39 $X2=0
+ $Y2=0
cc_664 N_A_603_191#_c_827_n N_VGND_c_1717_n 9.54497e-19 $X=5.72 $Y=1.39 $X2=0
+ $Y2=0
cc_665 N_A_603_191#_c_866_n A_762_191# 0.00793613f $X=4.07 $Y=1.115 $X2=-0.19
+ $Y2=-0.245
cc_666 N_A_603_191#_c_846_n A_848_191# 0.00452789f $X=5.41 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_667 N_A_28_108#_M1005_g N_A_1440_304#_M1033_g 0.0412786f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_668 N_A_28_108#_M1029_g N_A_1245_128#_c_1205_n 0.00151796f $X=6.39 $Y=2.48
+ $X2=0 $Y2=0
cc_669 N_A_28_108#_c_928_n N_A_1245_128#_c_1178_n 0.00385409f $X=6.95 $Y=0.18
+ $X2=0 $Y2=0
cc_670 N_A_28_108#_M1005_g N_A_1245_128#_c_1178_n 0.0169529f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_671 N_A_28_108#_M1005_g N_A_1245_128#_c_1179_n 0.00627841f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_672 N_A_28_108#_M1029_g N_A_1245_128#_c_1189_n 9.60337e-19 $X=6.39 $Y=2.48
+ $X2=0 $Y2=0
cc_673 N_A_28_108#_M1028_g N_VPWR_c_1458_n 0.0107891f $X=0.91 $Y=2.68 $X2=0
+ $Y2=0
cc_674 N_A_28_108#_c_940_n N_VPWR_c_1458_n 0.0071807f $X=0.985 $Y=3.15 $X2=0
+ $Y2=0
cc_675 N_A_28_108#_c_934_n N_VPWR_c_1458_n 0.0262636f $X=0.265 $Y=2.515 $X2=0
+ $Y2=0
cc_676 N_A_28_108#_c_939_n N_VPWR_c_1459_n 0.0264276f $X=2.865 $Y=3.15 $X2=0
+ $Y2=0
cc_677 N_A_28_108#_M1003_g N_VPWR_c_1459_n 0.00557219f $X=2.94 $Y=1.165 $X2=0
+ $Y2=0
cc_678 N_A_28_108#_M1011_g N_VPWR_c_1460_n 0.0063441f $X=3.87 $Y=2.525 $X2=0
+ $Y2=0
cc_679 N_A_28_108#_c_945_n N_VPWR_c_1460_n 0.0254009f $X=6.315 $Y=3.15 $X2=0
+ $Y2=0
cc_680 N_A_28_108#_c_945_n N_VPWR_c_1461_n 0.025796f $X=6.315 $Y=3.15 $X2=0
+ $Y2=0
cc_681 N_A_28_108#_M1029_g N_VPWR_c_1461_n 0.00384505f $X=6.39 $Y=2.48 $X2=0
+ $Y2=0
cc_682 N_A_28_108#_c_934_n N_VPWR_c_1472_n 0.0137031f $X=0.265 $Y=2.515 $X2=0
+ $Y2=0
cc_683 N_A_28_108#_c_940_n N_VPWR_c_1473_n 0.0330288f $X=0.985 $Y=3.15 $X2=0
+ $Y2=0
cc_684 N_A_28_108#_c_939_n N_VPWR_c_1474_n 0.0597153f $X=2.865 $Y=3.15 $X2=0
+ $Y2=0
cc_685 N_A_28_108#_c_945_n N_VPWR_c_1475_n 0.0212709f $X=6.315 $Y=3.15 $X2=0
+ $Y2=0
cc_686 N_A_28_108#_c_945_n N_VPWR_c_1476_n 0.0257875f $X=6.315 $Y=3.15 $X2=0
+ $Y2=0
cc_687 N_A_28_108#_c_939_n N_VPWR_c_1457_n 0.0467732f $X=2.865 $Y=3.15 $X2=0
+ $Y2=0
cc_688 N_A_28_108#_c_940_n N_VPWR_c_1457_n 0.00749832f $X=0.985 $Y=3.15 $X2=0
+ $Y2=0
cc_689 N_A_28_108#_c_943_n N_VPWR_c_1457_n 0.0222444f $X=3.795 $Y=3.15 $X2=0
+ $Y2=0
cc_690 N_A_28_108#_c_945_n N_VPWR_c_1457_n 0.0742071f $X=6.315 $Y=3.15 $X2=0
+ $Y2=0
cc_691 N_A_28_108#_c_948_n N_VPWR_c_1457_n 0.00421372f $X=2.94 $Y=3.15 $X2=0
+ $Y2=0
cc_692 N_A_28_108#_c_949_n N_VPWR_c_1457_n 0.00421372f $X=3.87 $Y=3.15 $X2=0
+ $Y2=0
cc_693 N_A_28_108#_c_934_n N_VPWR_c_1457_n 0.00975165f $X=0.265 $Y=2.515 $X2=0
+ $Y2=0
cc_694 N_A_28_108#_c_939_n N_A_304_463#_c_1603_n 0.00199547f $X=2.865 $Y=3.15
+ $X2=0 $Y2=0
cc_695 N_A_28_108#_M1003_g N_A_304_463#_c_1599_n 0.0177275f $X=2.94 $Y=1.165
+ $X2=0 $Y2=0
cc_696 N_A_28_108#_c_939_n N_A_304_463#_c_1601_n 0.00400794f $X=2.865 $Y=3.15
+ $X2=0 $Y2=0
cc_697 N_A_28_108#_M1003_g N_A_304_463#_c_1608_n 0.00380809f $X=2.94 $Y=1.165
+ $X2=0 $Y2=0
cc_698 N_A_28_108#_c_939_n N_A_304_463#_c_1602_n 0.00443431f $X=2.865 $Y=3.15
+ $X2=0 $Y2=0
cc_699 N_A_28_108#_M1003_g N_A_304_463#_c_1602_n 0.0274549f $X=2.94 $Y=1.165
+ $X2=0 $Y2=0
cc_700 N_A_28_108#_c_943_n N_A_304_463#_c_1602_n 0.00447307f $X=3.795 $Y=3.15
+ $X2=0 $Y2=0
cc_701 N_A_28_108#_c_929_n N_VGND_c_1703_n 0.0156678f $X=0.985 $Y=0.18 $X2=0
+ $Y2=0
cc_702 N_A_28_108#_c_935_n N_VGND_c_1703_n 0.0159659f $X=0.93 $Y=1.235 $X2=0
+ $Y2=0
cc_703 N_A_28_108#_c_936_n N_VGND_c_1703_n 9.30549e-19 $X=0.93 $Y=1.235 $X2=0
+ $Y2=0
cc_704 N_A_28_108#_M1014_g N_VGND_c_1704_n 0.00780385f $X=0.91 $Y=0.75 $X2=0
+ $Y2=0
cc_705 N_A_28_108#_c_928_n N_VGND_c_1704_n 0.0254714f $X=6.95 $Y=0.18 $X2=0
+ $Y2=0
cc_706 N_A_28_108#_c_928_n N_VGND_c_1705_n 0.0248335f $X=6.95 $Y=0.18 $X2=0
+ $Y2=0
cc_707 N_A_28_108#_c_928_n N_VGND_c_1706_n 0.0108684f $X=6.95 $Y=0.18 $X2=0
+ $Y2=0
cc_708 N_A_28_108#_c_928_n N_VGND_c_1709_n 0.0444293f $X=6.95 $Y=0.18 $X2=0
+ $Y2=0
cc_709 N_A_28_108#_c_933_n N_VGND_c_1711_n 0.00647699f $X=0.265 $Y=0.75 $X2=0
+ $Y2=0
cc_710 N_A_28_108#_c_929_n N_VGND_c_1712_n 0.0214934f $X=0.985 $Y=0.18 $X2=0
+ $Y2=0
cc_711 N_A_28_108#_c_928_n N_VGND_c_1713_n 0.0845253f $X=6.95 $Y=0.18 $X2=0
+ $Y2=0
cc_712 N_A_28_108#_c_928_n N_VGND_c_1717_n 0.170212f $X=6.95 $Y=0.18 $X2=0 $Y2=0
cc_713 N_A_28_108#_c_929_n N_VGND_c_1717_n 0.0112325f $X=0.985 $Y=0.18 $X2=0
+ $Y2=0
cc_714 N_A_28_108#_c_933_n N_VGND_c_1717_n 0.0102835f $X=0.265 $Y=0.75 $X2=0
+ $Y2=0
cc_715 N_A_1440_304#_c_1079_n N_A_1245_128#_c_1173_n 0.00403917f $X=8.61 $Y=0.85
+ $X2=0 $Y2=0
cc_716 N_A_1440_304#_c_1080_n N_A_1245_128#_c_1173_n 0.00240528f $X=8.7 $Y=1.6
+ $X2=0 $Y2=0
cc_717 N_A_1440_304#_c_1090_n N_A_1245_128#_M1006_g 0.00475915f $X=8.27 $Y=2.57
+ $X2=0 $Y2=0
cc_718 N_A_1440_304#_c_1091_n N_A_1245_128#_M1006_g 0.0101656f $X=8.292 $Y=2.345
+ $X2=0 $Y2=0
cc_719 N_A_1440_304#_c_1084_n N_A_1245_128#_M1006_g 0.0262074f $X=8.7 $Y=1.785
+ $X2=0 $Y2=0
cc_720 N_A_1440_304#_c_1079_n N_A_1245_128#_M1031_g 0.00272324f $X=8.61 $Y=0.85
+ $X2=0 $Y2=0
cc_721 N_A_1440_304#_M1033_g N_A_1245_128#_c_1178_n 0.00228324f $X=7.385 $Y=0.85
+ $X2=0 $Y2=0
cc_722 N_A_1440_304#_M1033_g N_A_1245_128#_c_1179_n 0.0175403f $X=7.385 $Y=0.85
+ $X2=0 $Y2=0
cc_723 N_A_1440_304#_c_1081_n N_A_1245_128#_c_1179_n 0.0248829f $X=7.365
+ $Y=1.685 $X2=0 $Y2=0
cc_724 N_A_1440_304#_c_1082_n N_A_1245_128#_c_1179_n 0.00518373f $X=7.365
+ $Y=1.685 $X2=0 $Y2=0
cc_725 N_A_1440_304#_c_1083_n N_A_1245_128#_c_1179_n 0.0241816f $X=8.25 $Y=1.785
+ $X2=0 $Y2=0
cc_726 N_A_1440_304#_M1033_g N_A_1245_128#_c_1180_n 0.00122798f $X=7.385 $Y=0.85
+ $X2=0 $Y2=0
cc_727 N_A_1440_304#_c_1080_n N_A_1245_128#_c_1180_n 0.00492208f $X=8.7 $Y=1.6
+ $X2=0 $Y2=0
cc_728 N_A_1440_304#_c_1079_n N_A_1245_128#_c_1181_n 0.0408812f $X=8.61 $Y=0.85
+ $X2=0 $Y2=0
cc_729 N_A_1440_304#_c_1079_n N_A_1245_128#_c_1183_n 0.0128645f $X=8.61 $Y=0.85
+ $X2=0 $Y2=0
cc_730 N_A_1440_304#_c_1080_n N_A_1245_128#_c_1183_n 0.0182108f $X=8.7 $Y=1.6
+ $X2=0 $Y2=0
cc_731 N_A_1440_304#_c_1083_n N_A_1245_128#_c_1183_n 0.0290943f $X=8.25 $Y=1.785
+ $X2=0 $Y2=0
cc_732 N_A_1440_304#_M1033_g N_A_1245_128#_c_1189_n 0.00221992f $X=7.385 $Y=0.85
+ $X2=0 $Y2=0
cc_733 N_A_1440_304#_c_1081_n N_A_1245_128#_c_1189_n 0.0227178f $X=7.365
+ $Y=1.685 $X2=0 $Y2=0
cc_734 N_A_1440_304#_c_1082_n N_A_1245_128#_c_1189_n 0.00127577f $X=7.365
+ $Y=1.685 $X2=0 $Y2=0
cc_735 N_A_1440_304#_M1033_g N_A_1245_128#_c_1191_n 2.85608e-19 $X=7.385 $Y=0.85
+ $X2=0 $Y2=0
cc_736 N_A_1440_304#_c_1083_n N_A_1245_128#_c_1191_n 0.0136635f $X=8.25 $Y=1.785
+ $X2=0 $Y2=0
cc_737 N_A_1440_304#_c_1079_n N_A_1245_128#_c_1192_n 0.00915093f $X=8.61 $Y=0.85
+ $X2=0 $Y2=0
cc_738 N_A_1440_304#_c_1079_n N_A_1245_128#_c_1193_n 0.0047842f $X=8.61 $Y=0.85
+ $X2=0 $Y2=0
cc_739 N_A_1440_304#_c_1079_n N_A_1245_128#_c_1198_n 0.00830453f $X=8.61 $Y=0.85
+ $X2=0 $Y2=0
cc_740 N_A_1440_304#_c_1080_n N_A_1245_128#_c_1198_n 0.0110879f $X=8.7 $Y=1.6
+ $X2=0 $Y2=0
cc_741 N_A_1440_304#_c_1083_n N_A_1245_128#_c_1198_n 0.0076918f $X=8.25 $Y=1.785
+ $X2=0 $Y2=0
cc_742 N_A_1440_304#_c_1079_n N_A_1796_139#_c_1376_n 0.00438052f $X=8.61 $Y=0.85
+ $X2=0 $Y2=0
cc_743 N_A_1440_304#_c_1080_n N_A_1796_139#_c_1376_n 0.0184546f $X=8.7 $Y=1.6
+ $X2=0 $Y2=0
cc_744 N_A_1440_304#_c_1080_n N_A_1796_139#_c_1377_n 0.0231793f $X=8.7 $Y=1.6
+ $X2=0 $Y2=0
cc_745 N_A_1440_304#_c_1091_n N_A_1796_139#_c_1377_n 0.0055477f $X=8.292
+ $Y=2.345 $X2=0 $Y2=0
cc_746 N_A_1440_304#_c_1084_n N_A_1796_139#_c_1377_n 0.0269579f $X=8.7 $Y=1.785
+ $X2=0 $Y2=0
cc_747 N_A_1440_304#_c_1091_n N_A_1796_139#_c_1383_n 0.00213431f $X=8.292
+ $Y=2.345 $X2=0 $Y2=0
cc_748 N_A_1440_304#_c_1091_n N_A_1796_139#_c_1386_n 0.00549902f $X=8.292
+ $Y=2.345 $X2=0 $Y2=0
cc_749 N_A_1440_304#_M1001_g N_VPWR_c_1462_n 0.0122105f $X=7.275 $Y=2.57 $X2=0
+ $Y2=0
cc_750 N_A_1440_304#_c_1087_n N_VPWR_c_1462_n 0.00116525f $X=7.365 $Y=2.19 $X2=0
+ $Y2=0
cc_751 N_A_1440_304#_c_1081_n N_VPWR_c_1462_n 0.0112645f $X=7.365 $Y=1.685 $X2=0
+ $Y2=0
cc_752 N_A_1440_304#_c_1083_n N_VPWR_c_1462_n 0.00261904f $X=8.25 $Y=1.785 $X2=0
+ $Y2=0
cc_753 N_A_1440_304#_c_1084_n N_VPWR_c_1463_n 0.00828564f $X=8.7 $Y=1.785 $X2=0
+ $Y2=0
cc_754 N_A_1440_304#_c_1090_n N_VPWR_c_1466_n 0.00446578f $X=8.27 $Y=2.57 $X2=0
+ $Y2=0
cc_755 N_A_1440_304#_M1001_g N_VPWR_c_1476_n 0.00379909f $X=7.275 $Y=2.57 $X2=0
+ $Y2=0
cc_756 N_A_1440_304#_M1001_g N_VPWR_c_1457_n 0.00412152f $X=7.275 $Y=2.57 $X2=0
+ $Y2=0
cc_757 N_A_1440_304#_c_1090_n N_VPWR_c_1457_n 0.00781865f $X=8.27 $Y=2.57 $X2=0
+ $Y2=0
cc_758 N_A_1440_304#_M1033_g N_VGND_c_1706_n 0.00312951f $X=7.385 $Y=0.85 $X2=0
+ $Y2=0
cc_759 N_A_1440_304#_M1033_g N_VGND_c_1709_n 0.00407505f $X=7.385 $Y=0.85 $X2=0
+ $Y2=0
cc_760 N_A_1440_304#_M1033_g N_VGND_c_1717_n 0.00465306f $X=7.385 $Y=0.85 $X2=0
+ $Y2=0
cc_761 N_A_1245_128#_c_1184_n N_A_1796_139#_M1031_s 0.00287157f $X=9.46 $Y=0.71
+ $X2=-0.19 $Y2=-0.245
cc_762 N_A_1245_128#_c_1192_n N_A_1796_139#_M1031_s 0.00269874f $X=9.045 $Y=0.43
+ $X2=-0.19 $Y2=-0.245
cc_763 N_A_1245_128#_M1031_g N_A_1796_139#_M1007_g 0.0180882f $X=9.455 $Y=0.905
+ $X2=0 $Y2=0
cc_764 N_A_1245_128#_c_1187_n N_A_1796_139#_M1007_g 5.62484e-19 $X=9.43 $Y=1.49
+ $X2=0 $Y2=0
cc_765 N_A_1245_128#_c_1188_n N_A_1796_139#_M1007_g 0.016611f $X=10.825 $Y=0.71
+ $X2=0 $Y2=0
cc_766 N_A_1245_128#_c_1193_n N_A_1796_139#_M1007_g 0.00623321f $X=9.492
+ $Y=1.325 $X2=0 $Y2=0
cc_767 N_A_1245_128#_c_1196_n N_A_1796_139#_M1007_g 0.00174094f $X=10.93 $Y=1.35
+ $X2=0 $Y2=0
cc_768 N_A_1245_128#_M1023_g N_A_1796_139#_c_1375_n 0.0214619f $X=10.965
+ $Y=2.465 $X2=0 $Y2=0
cc_769 N_A_1245_128#_M1031_g N_A_1796_139#_c_1376_n 0.00591751f $X=9.455
+ $Y=0.905 $X2=0 $Y2=0
cc_770 N_A_1245_128#_c_1184_n N_A_1796_139#_c_1376_n 0.0120136f $X=9.46 $Y=0.71
+ $X2=0 $Y2=0
cc_771 N_A_1245_128#_c_1187_n N_A_1796_139#_c_1376_n 0.00102469f $X=9.43 $Y=1.49
+ $X2=0 $Y2=0
cc_772 N_A_1245_128#_c_1192_n N_A_1796_139#_c_1376_n 0.0145709f $X=9.045 $Y=0.43
+ $X2=0 $Y2=0
cc_773 N_A_1245_128#_c_1193_n N_A_1796_139#_c_1376_n 0.0185241f $X=9.492
+ $Y=1.325 $X2=0 $Y2=0
cc_774 N_A_1245_128#_M1006_g N_A_1796_139#_c_1377_n 0.00457096f $X=8.485 $Y=2.57
+ $X2=0 $Y2=0
cc_775 N_A_1245_128#_M1031_g N_A_1796_139#_c_1377_n 0.00143634f $X=9.455
+ $Y=0.905 $X2=0 $Y2=0
cc_776 N_A_1245_128#_M1030_g N_A_1796_139#_c_1377_n 0.00382328f $X=9.455
+ $Y=2.755 $X2=0 $Y2=0
cc_777 N_A_1245_128#_c_1185_n N_A_1796_139#_c_1377_n 0.0477121f $X=9.492
+ $Y=1.472 $X2=0 $Y2=0
cc_778 N_A_1245_128#_c_1187_n N_A_1796_139#_c_1377_n 0.00832483f $X=9.43 $Y=1.49
+ $X2=0 $Y2=0
cc_779 N_A_1245_128#_c_1193_n N_A_1796_139#_c_1377_n 0.00352671f $X=9.492
+ $Y=1.325 $X2=0 $Y2=0
cc_780 N_A_1245_128#_M1006_g N_A_1796_139#_c_1383_n 0.00161561f $X=8.485 $Y=2.57
+ $X2=0 $Y2=0
cc_781 N_A_1245_128#_M1030_g N_A_1796_139#_c_1383_n 0.00415949f $X=9.455
+ $Y=2.755 $X2=0 $Y2=0
cc_782 N_A_1245_128#_M1030_g N_A_1796_139#_c_1384_n 0.0176375f $X=9.455 $Y=2.755
+ $X2=0 $Y2=0
cc_783 N_A_1245_128#_c_1204_n N_A_1796_139#_c_1384_n 0.00153546f $X=9.43
+ $Y=1.995 $X2=0 $Y2=0
cc_784 N_A_1245_128#_c_1186_n N_A_1796_139#_c_1384_n 0.0230434f $X=9.43 $Y=1.49
+ $X2=0 $Y2=0
cc_785 N_A_1245_128#_M1030_g N_A_1796_139#_c_1385_n 0.0034344f $X=9.455 $Y=2.755
+ $X2=0 $Y2=0
cc_786 N_A_1245_128#_c_1177_n N_A_1796_139#_c_1385_n 0.00195703f $X=9.43 $Y=1.83
+ $X2=0 $Y2=0
cc_787 N_A_1245_128#_c_1186_n N_A_1796_139#_c_1385_n 0.023172f $X=9.43 $Y=1.49
+ $X2=0 $Y2=0
cc_788 N_A_1245_128#_M1006_g N_A_1796_139#_c_1386_n 0.00311432f $X=8.485 $Y=2.57
+ $X2=0 $Y2=0
cc_789 N_A_1245_128#_c_1204_n N_A_1796_139#_c_1386_n 0.00287949f $X=9.43
+ $Y=1.995 $X2=0 $Y2=0
cc_790 N_A_1245_128#_c_1185_n N_A_1796_139#_c_1378_n 0.023172f $X=9.492 $Y=1.472
+ $X2=0 $Y2=0
cc_791 N_A_1245_128#_c_1187_n N_A_1796_139#_c_1378_n 3.67379e-19 $X=9.43 $Y=1.49
+ $X2=0 $Y2=0
cc_792 N_A_1245_128#_c_1188_n N_A_1796_139#_c_1378_n 0.00580242f $X=10.825
+ $Y=0.71 $X2=0 $Y2=0
cc_793 N_A_1245_128#_c_1185_n N_A_1796_139#_c_1379_n 0.00203396f $X=9.492
+ $Y=1.472 $X2=0 $Y2=0
cc_794 N_A_1245_128#_c_1187_n N_A_1796_139#_c_1379_n 0.0211439f $X=9.43 $Y=1.49
+ $X2=0 $Y2=0
cc_795 N_A_1245_128#_c_1188_n N_A_1796_139#_c_1379_n 0.00118075f $X=10.825
+ $Y=0.71 $X2=0 $Y2=0
cc_796 N_A_1245_128#_c_1196_n N_A_1796_139#_c_1379_n 0.00205542f $X=10.93
+ $Y=1.35 $X2=0 $Y2=0
cc_797 N_A_1245_128#_M1006_g N_VPWR_c_1462_n 4.52216e-19 $X=8.485 $Y=2.57 $X2=0
+ $Y2=0
cc_798 N_A_1245_128#_c_1206_n N_VPWR_c_1462_n 0.0113763f $X=6.605 $Y=2.205 $X2=0
+ $Y2=0
cc_799 N_A_1245_128#_M1006_g N_VPWR_c_1463_n 0.00403341f $X=8.485 $Y=2.57 $X2=0
+ $Y2=0
cc_800 N_A_1245_128#_M1030_g N_VPWR_c_1463_n 0.00282018f $X=9.455 $Y=2.755 $X2=0
+ $Y2=0
cc_801 N_A_1245_128#_M1030_g N_VPWR_c_1464_n 0.012947f $X=9.455 $Y=2.755 $X2=0
+ $Y2=0
cc_802 N_A_1245_128#_M1023_g N_VPWR_c_1465_n 0.00419321f $X=10.965 $Y=2.465
+ $X2=0 $Y2=0
cc_803 N_A_1245_128#_c_1195_n N_VPWR_c_1465_n 0.00218524f $X=10.93 $Y=1.35 $X2=0
+ $Y2=0
cc_804 N_A_1245_128#_c_1196_n N_VPWR_c_1465_n 0.00262673f $X=10.93 $Y=1.35 $X2=0
+ $Y2=0
cc_805 N_A_1245_128#_M1006_g N_VPWR_c_1466_n 0.00450619f $X=8.485 $Y=2.57 $X2=0
+ $Y2=0
cc_806 N_A_1245_128#_M1030_g N_VPWR_c_1468_n 0.00469214f $X=9.455 $Y=2.755 $X2=0
+ $Y2=0
cc_807 N_A_1245_128#_c_1206_n N_VPWR_c_1476_n 0.0112394f $X=6.605 $Y=2.205 $X2=0
+ $Y2=0
cc_808 N_A_1245_128#_M1023_g N_VPWR_c_1477_n 0.00579312f $X=10.965 $Y=2.465
+ $X2=0 $Y2=0
cc_809 N_A_1245_128#_M1006_g N_VPWR_c_1457_n 0.00490658f $X=8.485 $Y=2.57 $X2=0
+ $Y2=0
cc_810 N_A_1245_128#_M1030_g N_VPWR_c_1457_n 0.00945295f $X=9.455 $Y=2.755 $X2=0
+ $Y2=0
cc_811 N_A_1245_128#_M1023_g N_VPWR_c_1457_n 0.0115774f $X=10.965 $Y=2.465 $X2=0
+ $Y2=0
cc_812 N_A_1245_128#_c_1206_n N_VPWR_c_1457_n 0.0112734f $X=6.605 $Y=2.205 $X2=0
+ $Y2=0
cc_813 N_A_1245_128#_c_1188_n N_Q_M1007_d 0.0073298f $X=10.825 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_814 N_A_1245_128#_c_1188_n N_Q_c_1650_n 0.0207331f $X=10.825 $Y=0.71 $X2=0
+ $Y2=0
cc_815 N_A_1245_128#_c_1193_n N_Q_c_1650_n 0.00701341f $X=9.492 $Y=1.325 $X2=0
+ $Y2=0
cc_816 N_A_1245_128#_c_1197_n N_Q_c_1650_n 0.00864392f $X=10.92 $Y=1.185 $X2=0
+ $Y2=0
cc_817 N_A_1245_128#_c_1199_n N_Q_c_1650_n 9.91526e-19 $X=10.942 $Y=1.185 $X2=0
+ $Y2=0
cc_818 N_A_1245_128#_M1023_g Q 0.00196438f $X=10.965 $Y=2.465 $X2=0 $Y2=0
cc_819 N_A_1245_128#_c_1193_n Q 0.0057755f $X=9.492 $Y=1.325 $X2=0 $Y2=0
cc_820 N_A_1245_128#_c_1196_n Q 0.00318319f $X=10.93 $Y=1.35 $X2=0 $Y2=0
cc_821 N_A_1245_128#_c_1197_n Q 0.0137316f $X=10.92 $Y=1.185 $X2=0 $Y2=0
cc_822 N_A_1245_128#_M1030_g Q 0.00372326f $X=9.455 $Y=2.755 $X2=0 $Y2=0
cc_823 N_A_1245_128#_c_1197_n Q_N 0.0109f $X=10.92 $Y=1.185 $X2=0 $Y2=0
cc_824 N_A_1245_128#_c_1199_n Q_N 0.00277139f $X=10.942 $Y=1.185 $X2=0 $Y2=0
cc_825 N_A_1245_128#_M1023_g Q_N 0.0111967f $X=10.965 $Y=2.465 $X2=0 $Y2=0
cc_826 N_A_1245_128#_c_1195_n Q_N 0.0245418f $X=10.93 $Y=1.35 $X2=0 $Y2=0
cc_827 N_A_1245_128#_c_1197_n Q_N 0.00604183f $X=10.92 $Y=1.185 $X2=0 $Y2=0
cc_828 N_A_1245_128#_c_1199_n Q_N 0.0105699f $X=10.942 $Y=1.185 $X2=0 $Y2=0
cc_829 N_A_1245_128#_M1023_g Q_N 0.00206448f $X=10.965 $Y=2.465 $X2=0 $Y2=0
cc_830 N_A_1245_128#_c_1196_n Q_N 0.00335105f $X=10.93 $Y=1.35 $X2=0 $Y2=0
cc_831 N_A_1245_128#_M1023_g Q_N 0.0124115f $X=10.965 $Y=2.465 $X2=0 $Y2=0
cc_832 N_A_1245_128#_c_1188_n N_VGND_M1031_d 0.0113433f $X=10.825 $Y=0.71 $X2=0
+ $Y2=0
cc_833 N_A_1245_128#_c_1193_n N_VGND_M1031_d 0.00425849f $X=9.492 $Y=1.325 $X2=0
+ $Y2=0
cc_834 N_A_1245_128#_c_1188_n N_VGND_M1008_s 0.00720346f $X=10.825 $Y=0.71 $X2=0
+ $Y2=0
cc_835 N_A_1245_128#_c_1197_n N_VGND_M1008_s 0.00822136f $X=10.92 $Y=1.185 $X2=0
+ $Y2=0
cc_836 N_A_1245_128#_c_1178_n N_VGND_c_1706_n 0.00430849f $X=6.705 $Y=0.795
+ $X2=0 $Y2=0
cc_837 N_A_1245_128#_c_1179_n N_VGND_c_1706_n 0.00972448f $X=7.875 $Y=1.34 $X2=0
+ $Y2=0
cc_838 N_A_1245_128#_c_1180_n N_VGND_c_1706_n 0.0178415f $X=7.96 $Y=1.19 $X2=0
+ $Y2=0
cc_839 N_A_1245_128#_c_1182_n N_VGND_c_1706_n 0.0133497f $X=8.045 $Y=0.43 $X2=0
+ $Y2=0
cc_840 N_A_1245_128#_c_1188_n N_VGND_c_1707_n 0.0203332f $X=10.825 $Y=0.71 $X2=0
+ $Y2=0
cc_841 N_A_1245_128#_c_1192_n N_VGND_c_1707_n 0.00431819f $X=9.045 $Y=0.43 $X2=0
+ $Y2=0
cc_842 N_A_1245_128#_c_1194_n N_VGND_c_1707_n 0.00340062f $X=9.55 $Y=0.71 $X2=0
+ $Y2=0
cc_843 N_A_1245_128#_c_1188_n N_VGND_c_1708_n 0.0213396f $X=10.825 $Y=0.71 $X2=0
+ $Y2=0
cc_844 N_A_1245_128#_c_1199_n N_VGND_c_1708_n 0.00894929f $X=10.942 $Y=1.185
+ $X2=0 $Y2=0
cc_845 N_A_1245_128#_c_1178_n N_VGND_c_1709_n 0.00404505f $X=6.705 $Y=0.795
+ $X2=0 $Y2=0
cc_846 N_A_1245_128#_c_1173_n N_VGND_c_1714_n 5.82898e-19 $X=8.175 $Y=1.17 $X2=0
+ $Y2=0
cc_847 N_A_1245_128#_M1031_g N_VGND_c_1714_n 0.00294786f $X=9.455 $Y=0.905 $X2=0
+ $Y2=0
cc_848 N_A_1245_128#_c_1181_n N_VGND_c_1714_n 0.037645f $X=8.96 $Y=0.43 $X2=0
+ $Y2=0
cc_849 N_A_1245_128#_c_1182_n N_VGND_c_1714_n 0.00774075f $X=8.045 $Y=0.43 $X2=0
+ $Y2=0
cc_850 N_A_1245_128#_c_1184_n N_VGND_c_1714_n 0.00598765f $X=9.46 $Y=0.71 $X2=0
+ $Y2=0
cc_851 N_A_1245_128#_c_1192_n N_VGND_c_1714_n 0.00742542f $X=9.045 $Y=0.43 $X2=0
+ $Y2=0
cc_852 N_A_1245_128#_c_1194_n N_VGND_c_1714_n 0.00272132f $X=9.55 $Y=0.71 $X2=0
+ $Y2=0
cc_853 N_A_1245_128#_c_1188_n N_VGND_c_1715_n 0.0124196f $X=10.825 $Y=0.71 $X2=0
+ $Y2=0
cc_854 N_A_1245_128#_c_1199_n N_VGND_c_1716_n 0.00486043f $X=10.942 $Y=1.185
+ $X2=0 $Y2=0
cc_855 N_A_1245_128#_M1031_g N_VGND_c_1717_n 0.0045051f $X=9.455 $Y=0.905 $X2=0
+ $Y2=0
cc_856 N_A_1245_128#_c_1178_n N_VGND_c_1717_n 0.00525146f $X=6.705 $Y=0.795
+ $X2=0 $Y2=0
cc_857 N_A_1245_128#_c_1181_n N_VGND_c_1717_n 0.0324621f $X=8.96 $Y=0.43 $X2=0
+ $Y2=0
cc_858 N_A_1245_128#_c_1182_n N_VGND_c_1717_n 0.00629746f $X=8.045 $Y=0.43 $X2=0
+ $Y2=0
cc_859 N_A_1245_128#_c_1184_n N_VGND_c_1717_n 0.00941265f $X=9.46 $Y=0.71 $X2=0
+ $Y2=0
cc_860 N_A_1245_128#_c_1188_n N_VGND_c_1717_n 0.0234023f $X=10.825 $Y=0.71 $X2=0
+ $Y2=0
cc_861 N_A_1245_128#_c_1192_n N_VGND_c_1717_n 0.00613972f $X=9.045 $Y=0.43 $X2=0
+ $Y2=0
cc_862 N_A_1245_128#_c_1194_n N_VGND_c_1717_n 0.00444552f $X=9.55 $Y=0.71 $X2=0
+ $Y2=0
cc_863 N_A_1245_128#_c_1199_n N_VGND_c_1717_n 0.00917987f $X=10.942 $Y=1.185
+ $X2=0 $Y2=0
cc_864 N_A_1796_139#_c_1383_n N_VPWR_c_1463_n 0.0530452f $X=9.24 $Y=2.56 $X2=0
+ $Y2=0
cc_865 N_A_1796_139#_M1004_g N_VPWR_c_1464_n 0.00352559f $X=10.48 $Y=2.465 $X2=0
+ $Y2=0
cc_866 N_A_1796_139#_c_1384_n N_VPWR_c_1464_n 0.0240235f $X=9.83 $Y=2.25 $X2=0
+ $Y2=0
cc_867 N_A_1796_139#_M1004_g N_VPWR_c_1465_n 0.00403052f $X=10.48 $Y=2.465 $X2=0
+ $Y2=0
cc_868 N_A_1796_139#_c_1383_n N_VPWR_c_1468_n 0.0217713f $X=9.24 $Y=2.56 $X2=0
+ $Y2=0
cc_869 N_A_1796_139#_M1004_g N_VPWR_c_1470_n 0.0054895f $X=10.48 $Y=2.465 $X2=0
+ $Y2=0
cc_870 N_A_1796_139#_M1004_g N_VPWR_c_1457_n 0.0112178f $X=10.48 $Y=2.465 $X2=0
+ $Y2=0
cc_871 N_A_1796_139#_c_1383_n N_VPWR_c_1457_n 0.0126859f $X=9.24 $Y=2.56 $X2=0
+ $Y2=0
cc_872 N_A_1796_139#_M1007_g N_Q_c_1650_n 0.00465688f $X=10.04 $Y=0.765 $X2=0
+ $Y2=0
cc_873 N_A_1796_139#_c_1375_n N_Q_c_1650_n 0.00264885f $X=10.405 $Y=1.6 $X2=0
+ $Y2=0
cc_874 N_A_1796_139#_M1007_g Q 0.00254982f $X=10.04 $Y=0.765 $X2=0 $Y2=0
cc_875 N_A_1796_139#_c_1375_n Q 0.0157902f $X=10.405 $Y=1.6 $X2=0 $Y2=0
cc_876 N_A_1796_139#_M1004_g Q 0.0057137f $X=10.48 $Y=2.465 $X2=0 $Y2=0
cc_877 N_A_1796_139#_c_1385_n Q 0.0105985f $X=9.915 $Y=2.165 $X2=0 $Y2=0
cc_878 N_A_1796_139#_c_1378_n Q 0.0238766f $X=9.97 $Y=1.51 $X2=0 $Y2=0
cc_879 N_A_1796_139#_c_1379_n Q 0.00226557f $X=9.97 $Y=1.51 $X2=0 $Y2=0
cc_880 N_A_1796_139#_c_1375_n Q 0.00221984f $X=10.405 $Y=1.6 $X2=0 $Y2=0
cc_881 N_A_1796_139#_M1004_g Q 0.00132541f $X=10.48 $Y=2.465 $X2=0 $Y2=0
cc_882 N_A_1796_139#_c_1385_n Q 0.024356f $X=9.915 $Y=2.165 $X2=0 $Y2=0
cc_883 N_A_1796_139#_M1004_g Q 0.0135044f $X=10.48 $Y=2.465 $X2=0 $Y2=0
cc_884 N_A_1796_139#_c_1384_n Q 0.014539f $X=9.83 $Y=2.25 $X2=0 $Y2=0
cc_885 N_A_1796_139#_M1007_g N_VGND_c_1707_n 0.00750547f $X=10.04 $Y=0.765 $X2=0
+ $Y2=0
cc_886 N_A_1796_139#_M1007_g N_VGND_c_1708_n 0.00567452f $X=10.04 $Y=0.765 $X2=0
+ $Y2=0
cc_887 N_A_1796_139#_M1007_g N_VGND_c_1715_n 0.00341315f $X=10.04 $Y=0.765 $X2=0
+ $Y2=0
cc_888 N_A_1796_139#_M1007_g N_VGND_c_1717_n 0.00507883f $X=10.04 $Y=0.765 $X2=0
+ $Y2=0
cc_889 N_VPWR_M1025_d N_A_304_463#_c_1603_n 0.00627455f $X=1.935 $Y=2.315 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_1459_n N_A_304_463#_c_1603_n 0.0235704f $X=2.145 $Y=2.75 $X2=0
+ $Y2=0
cc_891 N_VPWR_c_1457_n N_A_304_463#_c_1603_n 0.0143212f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_892 N_VPWR_c_1473_n N_A_304_463#_c_1601_n 0.00421736f $X=1.97 $Y=3.33 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_1457_n N_A_304_463#_c_1601_n 0.00552714f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_894 N_VPWR_c_1474_n N_A_304_463#_c_1602_n 0.01602f $X=4.34 $Y=3.33 $X2=0
+ $Y2=0
cc_895 N_VPWR_c_1457_n N_A_304_463#_c_1602_n 0.0214601f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_896 N_VPWR_c_1457_n N_Q_M1004_s 0.00323f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_897 N_VPWR_c_1465_n Q 0.0458614f $X=10.73 $Y=1.985 $X2=0 $Y2=0
cc_898 N_VPWR_c_1464_n Q 0.0282409f $X=9.67 $Y=2.59 $X2=0 $Y2=0
cc_899 N_VPWR_c_1470_n Q 0.0160712f $X=10.6 $Y=3.33 $X2=0 $Y2=0
cc_900 N_VPWR_c_1457_n Q 0.00984745f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_901 N_VPWR_c_1457_n N_Q_N_M1023_d 0.00231914f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_902 N_VPWR_c_1465_n Q_N 0.0490221f $X=10.73 $Y=1.985 $X2=0 $Y2=0
cc_903 N_VPWR_c_1477_n Q_N 0.0261075f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_904 N_VPWR_c_1457_n Q_N 0.0153818f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_905 N_Q_N_c_1683_n N_VGND_c_1716_n 0.018528f $X=11.26 $Y=0.42 $X2=0 $Y2=0
cc_906 N_Q_N_M1008_d N_VGND_c_1717_n 0.00371702f $X=11.12 $Y=0.235 $X2=0 $Y2=0
cc_907 N_Q_N_c_1683_n N_VGND_c_1717_n 0.0104192f $X=11.26 $Y=0.42 $X2=0 $Y2=0
