* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor2_m A B VGND VNB VPB VPWR Y
X0 Y a_56_90# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 Y a_56_90# a_297_90# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR B a_56_90# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR A a_311_422# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_311_422# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_139_90# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_56_90# B a_139_90# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND A a_297_90# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_297_90# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_56_90# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
