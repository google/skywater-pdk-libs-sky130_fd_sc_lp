* File: sky130_fd_sc_lp__dlrtp_2.spice
* Created: Wed Sep  2 09:47:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrtp_2.pex.spice"
.subckt sky130_fd_sc_lp__dlrtp_2  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_D_M1011_g N_A_40_54#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.12705 AS=0.1113 PD=1.025 PS=1.37 NRD=89.988 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1019 N_A_251_475#_M1019_d N_GATE_M1019_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.12705 PD=1.41 PS=1.025 NRD=5.712 NRS=2.856 M=1 R=2.8
+ SA=75000.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_251_475#_M1021_g N_A_383_479#_M1021_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1004 A_574_47# N_A_40_54#_M1004_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_646_47#_M1007_d N_A_383_479#_M1007_g A_574_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1015 A_754_47# N_A_251_475#_M1015_g N_A_646_47#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_796_21#_M1005_g A_754_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1554 AS=0.0441 PD=1.58 PS=0.63 NRD=27.132 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1008 A_1043_73# N_A_646_47#_M1008_g N_A_796_21#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_RESET_B_M1002_g A_1043_73# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.0882 PD=1.23 PS=1.05 NRD=7.848 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1006 N_Q_M1006_d N_A_796_21#_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1659 AS=0.1638 PD=1.235 PS=1.23 NRD=9.996 NRS=7.848 M=1 R=5.6 SA=75001.1
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1016 N_Q_M1006_d N_A_796_21#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1659 AS=0.2478 PD=1.235 PS=2.27 NRD=6.42 NRS=2.856 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1017 N_VPWR_M1017_d N_D_M1017_g N_A_40_54#_M1017_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1568 AS=0.1696 PD=1.13 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1003 N_A_251_475#_M1003_d N_GATE_M1003_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.208 AS=0.1568 PD=1.93 PS=1.13 NRD=15.3857 NRS=64.6357 M=1
+ R=4.26667 SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 N_VPWR_M1020_d N_A_251_475#_M1020_g N_A_383_479#_M1020_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.184 AS=0.1696 PD=1.215 PS=1.81 NRD=83.0946 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1010 A_611_479# N_A_40_54#_M1010_g N_VPWR_M1020_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.184 PD=0.85 PS=1.215 NRD=15.3857 NRS=7.683 M=1 R=4.26667
+ SA=75000.9 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1013 N_A_646_47#_M1013_d N_A_251_475#_M1013_g A_611_479# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.124498 AS=0.0672 PD=1.20755 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.3 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1014 A_785_479# N_A_383_479#_M1014_g N_A_646_47#_M1013_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0817019 PD=0.66 PS=0.792453 NRD=30.4759 NRS=37.5088 M=1
+ R=2.8 SA=75001.8 SB=75003 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_796_21#_M1000_g A_785_479# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1344 AS=0.0504 PD=1.005 PS=0.66 NRD=111.384 NRS=30.4759 M=1 R=2.8
+ SA=75002.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_796_21#_M1012_d N_A_646_47#_M1012_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.4032 PD=1.54 PS=3.015 NRD=0 NRS=36.7405 M=1 R=8.4
+ SA=75001.2 SB=75001.7 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_RESET_B_M1018_g N_A_796_21#_M1012_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.34335 AS=0.1764 PD=1.805 PS=1.54 NRD=20.3107 NRS=0 M=1 R=8.4
+ SA=75001.6 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1018_d N_A_796_21#_M1001_g N_Q_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.34335 AS=0.1764 PD=1.805 PS=1.54 NRD=21.0987 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_796_21#_M1009_g N_Q_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX22_noxref VNB VPB NWDIODE A=14.1367 P=18.89
c_85 VNB 0 8.43473e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dlrtp_2.pxi.spice"
*
.ends
*
*
