* File: sky130_fd_sc_lp__a211oi_2.pxi.spice
* Created: Wed Sep  2 09:18:10 2020
* 
x_PM_SKY130_FD_SC_LP__A211OI_2%C1 N_C1_c_76_n N_C1_M1012_g N_C1_M1008_g
+ N_C1_c_78_n N_C1_M1013_g N_C1_M1014_g C1 C1 N_C1_c_81_n
+ PM_SKY130_FD_SC_LP__A211OI_2%C1
x_PM_SKY130_FD_SC_LP__A211OI_2%B1 N_B1_M1007_g N_B1_M1001_g N_B1_M1011_g
+ N_B1_M1009_g B1 B1 N_B1_c_120_n PM_SKY130_FD_SC_LP__A211OI_2%B1
x_PM_SKY130_FD_SC_LP__A211OI_2%A2 N_A2_M1004_g N_A2_M1000_g N_A2_M1005_g
+ N_A2_M1006_g N_A2_c_169_n N_A2_c_170_n N_A2_c_175_n A2 A2 N_A2_c_171_n
+ PM_SKY130_FD_SC_LP__A211OI_2%A2
x_PM_SKY130_FD_SC_LP__A211OI_2%A1 N_A1_c_223_n N_A1_M1002_g N_A1_M1003_g
+ N_A1_M1010_g N_A1_c_224_n N_A1_M1015_g N_A1_c_225_n A1 A1 N_A1_c_227_n
+ PM_SKY130_FD_SC_LP__A211OI_2%A1
x_PM_SKY130_FD_SC_LP__A211OI_2%A_41_367# N_A_41_367#_M1008_s N_A_41_367#_M1014_s
+ N_A_41_367#_M1009_d N_A_41_367#_c_271_n N_A_41_367#_c_272_n
+ N_A_41_367#_c_277_n N_A_41_367#_c_279_n N_A_41_367#_c_273_n
+ N_A_41_367#_c_274_n N_A_41_367#_c_295_p PM_SKY130_FD_SC_LP__A211OI_2%A_41_367#
x_PM_SKY130_FD_SC_LP__A211OI_2%Y N_Y_M1012_s N_Y_M1007_d N_Y_M1002_s N_Y_M1008_d
+ N_Y_c_306_n N_Y_c_307_n N_Y_c_303_n N_Y_c_304_n N_Y_c_338_n N_Y_c_313_n
+ N_Y_c_305_n Y Y N_Y_c_328_n PM_SKY130_FD_SC_LP__A211OI_2%Y
x_PM_SKY130_FD_SC_LP__A211OI_2%A_296_367# N_A_296_367#_M1001_s
+ N_A_296_367#_M1000_s N_A_296_367#_M1003_s N_A_296_367#_c_366_n
+ N_A_296_367#_c_363_n N_A_296_367#_c_370_n N_A_296_367#_c_397_p
+ N_A_296_367#_c_364_n N_A_296_367#_c_398_p N_A_296_367#_c_365_n
+ PM_SKY130_FD_SC_LP__A211OI_2%A_296_367#
x_PM_SKY130_FD_SC_LP__A211OI_2%VPWR N_VPWR_M1000_d N_VPWR_M1006_d N_VPWR_M1010_d
+ N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n VPWR
+ N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n N_VPWR_c_412_n N_VPWR_c_413_n
+ N_VPWR_c_404_n PM_SKY130_FD_SC_LP__A211OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A211OI_2%VGND N_VGND_M1012_d N_VGND_M1013_d N_VGND_M1011_s
+ N_VGND_M1004_d N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n
+ N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n VGND N_VGND_c_475_n
+ N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n N_VGND_c_479_n N_VGND_c_480_n
+ PM_SKY130_FD_SC_LP__A211OI_2%VGND
x_PM_SKY130_FD_SC_LP__A211OI_2%A_489_65# N_A_489_65#_M1004_s N_A_489_65#_M1005_s
+ N_A_489_65#_M1015_d N_A_489_65#_c_534_n N_A_489_65#_c_541_n
+ N_A_489_65#_c_535_n N_A_489_65#_c_544_n N_A_489_65#_c_536_n
+ N_A_489_65#_c_537_n N_A_489_65#_c_538_n PM_SKY130_FD_SC_LP__A211OI_2%A_489_65#
cc_1 VNB N_C1_c_76_n 0.022754f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.21
cc_2 VNB N_C1_M1008_g 0.00575006f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_3 VNB N_C1_c_78_n 0.0157081f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.21
cc_4 VNB N_C1_M1014_g 0.00547576f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_5 VNB C1 0.0228943f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_C1_c_81_n 0.0710597f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.375
cc_7 VNB N_B1_M1007_g 0.0224265f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.665
cc_8 VNB N_B1_M1011_g 0.0304927f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.54
cc_9 VNB B1 0.00373879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_c_120_n 0.0346084f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.295
cc_11 VNB N_A2_M1004_g 0.0274365f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.665
cc_12 VNB N_A2_M1005_g 0.0213363f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.54
cc_13 VNB N_A2_c_169_n 0.00136716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_170_n 0.00766091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_171_n 0.057952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_223_n 0.0163458f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.21
cc_17 VNB N_A1_c_224_n 0.0205698f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_18 VNB N_A1_c_225_n 0.00136843f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB A1 0.0202756f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_20 VNB N_A1_c_227_n 0.0789025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_303_n 0.004326f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_22 VNB N_Y_c_304_n 0.0270375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_305_n 0.00190113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_404_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_468_n 0.0124619f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_26 VNB N_VGND_c_469_n 0.035072f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_VGND_c_470_n 5.0291e-19 $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_28 VNB N_VGND_c_471_n 0.0115983f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_29 VNB N_VGND_c_472_n 0.00820588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_473_n 0.015042f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_31 VNB N_VGND_c_474_n 0.0053824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_475_n 0.0154973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_476_n 0.0187491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_477_n 0.0386225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_478_n 0.268867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_479_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_480_n 0.00632006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_489_65#_c_534_n 0.00630303f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_39 VNB N_A_489_65#_c_535_n 0.00189184f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_40 VNB N_A_489_65#_c_536_n 0.0121645f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_41 VNB N_A_489_65#_c_537_n 0.00203674f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_42 VNB N_A_489_65#_c_538_n 0.0233564f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.375
cc_43 VPB N_C1_M1008_g 0.0245703f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_44 VPB N_C1_M1014_g 0.0193745f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_45 VPB C1 0.0100517f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_46 VPB N_B1_M1001_g 0.0183355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B1_M1009_g 0.0239332f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_48 VPB B1 0.00657294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B1_c_120_n 0.00490112f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_50 VPB N_A2_M1000_g 0.0238526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A2_M1006_g 0.0180916f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_52 VPB N_A2_c_170_n 0.00810075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A2_c_175_n 0.00131986f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_54 VPB N_A2_c_171_n 0.0175458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A1_M1003_g 0.0180952f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_56 VPB N_A1_M1010_g 0.0233518f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=0.665
cc_57 VPB A1 0.00992715f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.375
cc_58 VPB N_A1_c_227_n 0.00450641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_41_367#_c_271_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=0.665
cc_60 VPB N_A_41_367#_c_272_n 0.0373257f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_61 VPB N_A_41_367#_c_273_n 0.00227906f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.375
cc_62 VPB N_A_41_367#_c_274_n 0.00776016f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.375
cc_63 VPB N_A_296_367#_c_363_n 0.0189431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_296_367#_c_364_n 0.00737761f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.375
cc_65 VPB N_A_296_367#_c_365_n 0.00218346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_405_n 0.0127427f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_67 VPB N_VPWR_c_406_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_68 VPB N_VPWR_c_407_n 0.0132106f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.375
cc_69 VPB N_VPWR_c_408_n 0.0482554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_409_n 0.0639702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_410_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_411_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_412_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_413_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_404_n 0.0658007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 N_C1_c_78_n N_B1_M1007_g 0.0185658f $X=0.975 $Y=1.21 $X2=0 $Y2=0
cc_77 N_C1_M1014_g N_B1_M1001_g 0.0185658f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_78 N_C1_c_81_n B1 0.00288466f $X=0.975 $Y=1.375 $X2=0 $Y2=0
cc_79 N_C1_c_81_n N_B1_c_120_n 0.0185658f $X=0.975 $Y=1.375 $X2=0 $Y2=0
cc_80 C1 N_A_41_367#_c_272_n 0.022879f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_C1_c_81_n N_A_41_367#_c_272_n 0.00119621f $X=0.975 $Y=1.375 $X2=0 $Y2=0
cc_82 N_C1_M1008_g N_A_41_367#_c_277_n 0.0115031f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_83 N_C1_M1014_g N_A_41_367#_c_277_n 0.0115031f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_84 N_C1_c_76_n N_Y_c_306_n 0.0109234f $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_85 N_C1_M1008_g N_Y_c_307_n 0.0221318f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_86 N_C1_M1014_g N_Y_c_307_n 0.0174077f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_87 C1 N_Y_c_307_n 0.0387702f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_88 N_C1_c_81_n N_Y_c_307_n 0.0195373f $X=0.975 $Y=1.375 $X2=0 $Y2=0
cc_89 N_C1_c_78_n N_Y_c_303_n 0.00785513f $X=0.975 $Y=1.21 $X2=0 $Y2=0
cc_90 N_C1_c_81_n N_Y_c_303_n 0.00628803f $X=0.975 $Y=1.375 $X2=0 $Y2=0
cc_91 N_C1_c_76_n N_Y_c_313_n 0.00778888f $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_92 N_C1_c_78_n N_Y_c_313_n 0.00302959f $X=0.975 $Y=1.21 $X2=0 $Y2=0
cc_93 C1 N_Y_c_313_n 0.00279991f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_94 N_C1_c_81_n N_Y_c_313_n 0.00405606f $X=0.975 $Y=1.375 $X2=0 $Y2=0
cc_95 N_C1_M1008_g N_VPWR_c_409_n 0.00357877f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_96 N_C1_M1014_g N_VPWR_c_409_n 0.00357877f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_97 N_C1_M1008_g N_VPWR_c_404_n 0.00634361f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_98 N_C1_M1014_g N_VPWR_c_404_n 0.00537654f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_99 N_C1_c_76_n N_VGND_c_469_n 0.00498793f $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_100 C1 N_VGND_c_469_n 0.021786f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_101 N_C1_c_81_n N_VGND_c_469_n 0.00193743f $X=0.975 $Y=1.375 $X2=0 $Y2=0
cc_102 N_C1_c_76_n N_VGND_c_470_n 6.87359e-19 $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_103 N_C1_c_78_n N_VGND_c_470_n 0.0113415f $X=0.975 $Y=1.21 $X2=0 $Y2=0
cc_104 N_C1_c_76_n N_VGND_c_475_n 0.00539298f $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_105 N_C1_c_78_n N_VGND_c_475_n 0.00477554f $X=0.975 $Y=1.21 $X2=0 $Y2=0
cc_106 N_C1_c_76_n N_VGND_c_478_n 0.0107711f $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_107 N_C1_c_78_n N_VGND_c_478_n 0.00825815f $X=0.975 $Y=1.21 $X2=0 $Y2=0
cc_108 B1 N_A2_c_170_n 0.0288708f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_109 N_B1_c_120_n N_A2_c_170_n 0.00508849f $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_110 N_B1_c_120_n N_A2_c_171_n 0.00688076f $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_111 B1 N_A_41_367#_c_279_n 0.0141407f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_112 N_B1_M1001_g N_A_41_367#_c_273_n 0.0115031f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B1_M1009_g N_A_41_367#_c_273_n 0.0115031f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_114 N_B1_M1007_g N_Y_c_307_n 9.40973e-19 $X=1.405 $Y=0.665 $X2=0 $Y2=0
cc_115 N_B1_M1001_g N_Y_c_307_n 9.99593e-19 $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_116 B1 N_Y_c_307_n 0.0251353f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_117 N_B1_c_120_n N_Y_c_307_n 2.43011e-19 $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_118 N_B1_M1007_g N_Y_c_303_n 0.01419f $X=1.405 $Y=0.665 $X2=0 $Y2=0
cc_119 B1 N_Y_c_303_n 0.0297732f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_120 N_B1_M1011_g N_Y_c_304_n 0.0158409f $X=1.835 $Y=0.665 $X2=0 $Y2=0
cc_121 B1 N_Y_c_304_n 0.00473669f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_122 N_B1_M1011_g N_Y_c_305_n 0.00205286f $X=1.835 $Y=0.665 $X2=0 $Y2=0
cc_123 B1 N_Y_c_305_n 0.0193461f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_124 N_B1_c_120_n N_Y_c_305_n 0.00255521f $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_125 N_B1_M1011_g N_Y_c_328_n 0.0140331f $X=1.835 $Y=0.665 $X2=0 $Y2=0
cc_126 N_B1_M1001_g N_A_296_367#_c_366_n 0.00840077f $X=1.405 $Y=2.465 $X2=0
+ $Y2=0
cc_127 N_B1_M1009_g N_A_296_367#_c_366_n 0.0142778f $X=1.835 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_B1_M1009_g N_A_296_367#_c_363_n 0.0143379f $X=1.835 $Y=2.465 $X2=0
+ $Y2=0
cc_129 B1 N_A_296_367#_c_363_n 0.00353236f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_130 N_B1_M1001_g N_A_296_367#_c_370_n 0.00207347f $X=1.405 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_B1_M1009_g N_A_296_367#_c_370_n 6.7411e-19 $X=1.835 $Y=2.465 $X2=0
+ $Y2=0
cc_132 B1 N_A_296_367#_c_370_n 0.0230324f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_133 N_B1_c_120_n N_A_296_367#_c_370_n 6.52992e-19 $X=1.835 $Y=1.51 $X2=0
+ $Y2=0
cc_134 N_B1_M1009_g N_VPWR_c_405_n 0.00175123f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_135 N_B1_M1001_g N_VPWR_c_409_n 0.00357877f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_136 N_B1_M1009_g N_VPWR_c_409_n 0.00357877f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_137 N_B1_M1001_g N_VPWR_c_404_n 0.00537654f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_138 N_B1_M1009_g N_VPWR_c_404_n 0.00665089f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_139 N_B1_M1007_g N_VGND_c_470_n 0.0113004f $X=1.405 $Y=0.665 $X2=0 $Y2=0
cc_140 N_B1_M1011_g N_VGND_c_470_n 6.93622e-19 $X=1.835 $Y=0.665 $X2=0 $Y2=0
cc_141 N_B1_M1011_g N_VGND_c_471_n 0.00326162f $X=1.835 $Y=0.665 $X2=0 $Y2=0
cc_142 N_B1_M1007_g N_VGND_c_473_n 0.00477554f $X=1.405 $Y=0.665 $X2=0 $Y2=0
cc_143 N_B1_M1011_g N_VGND_c_473_n 0.00569184f $X=1.835 $Y=0.665 $X2=0 $Y2=0
cc_144 N_B1_M1007_g N_VGND_c_478_n 0.00825815f $X=1.405 $Y=0.665 $X2=0 $Y2=0
cc_145 N_B1_M1011_g N_VGND_c_478_n 0.0117376f $X=1.835 $Y=0.665 $X2=0 $Y2=0
cc_146 N_A2_M1005_g N_A1_c_223_n 0.0201601f $X=3.375 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A2_M1006_g N_A1_M1003_g 0.0201601f $X=3.375 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A2_c_169_n N_A1_c_225_n 0.0101132f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A2_c_171_n N_A1_c_225_n 2.24742e-19 $X=3.375 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A2_c_169_n N_A1_c_227_n 2.24722e-19 $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A2_c_171_n N_A1_c_227_n 0.0201601f $X=3.375 $Y=1.51 $X2=0 $Y2=0
cc_152 N_A2_M1000_g N_A_41_367#_c_274_n 0.00160289f $X=2.945 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A2_M1004_g N_Y_c_304_n 0.0133336f $X=2.785 $Y=0.745 $X2=0 $Y2=0
cc_154 N_A2_M1005_g N_Y_c_304_n 0.0112465f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_155 N_A2_c_170_n N_Y_c_304_n 0.107433f $X=2.728 $Y=1.582 $X2=0 $Y2=0
cc_156 N_A2_c_171_n N_Y_c_304_n 0.0135879f $X=3.375 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A2_M1000_g N_A_296_367#_c_363_n 0.0149732f $X=2.945 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A2_c_169_n N_A_296_367#_c_363_n 0.0059402f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A2_c_170_n N_A_296_367#_c_363_n 0.0677577f $X=2.728 $Y=1.582 $X2=0
+ $Y2=0
cc_160 N_A2_c_171_n N_A_296_367#_c_363_n 0.00238517f $X=3.375 $Y=1.51 $X2=0
+ $Y2=0
cc_161 N_A2_M1006_g N_A_296_367#_c_364_n 0.0125328f $X=3.375 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A2_c_169_n N_A_296_367#_c_364_n 0.0134448f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_163 N_A2_M1000_g N_A_296_367#_c_365_n 0.00170776f $X=2.945 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A2_c_169_n N_A_296_367#_c_365_n 0.015226f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A2_c_171_n N_A_296_367#_c_365_n 0.00256759f $X=3.375 $Y=1.51 $X2=0
+ $Y2=0
cc_166 N_A2_M1000_g N_VPWR_c_405_n 0.0172659f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A2_M1006_g N_VPWR_c_405_n 6.80491e-19 $X=3.375 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A2_M1000_g N_VPWR_c_406_n 7.24342e-19 $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A2_M1006_g N_VPWR_c_406_n 0.0140821f $X=3.375 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A2_M1000_g N_VPWR_c_410_n 0.00486043f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A2_M1006_g N_VPWR_c_410_n 0.00486043f $X=3.375 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A2_M1000_g N_VPWR_c_404_n 0.00824727f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A2_M1006_g N_VPWR_c_404_n 0.00824727f $X=3.375 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A2_M1004_g N_VGND_c_471_n 0.00328393f $X=2.785 $Y=0.745 $X2=0 $Y2=0
cc_175 N_A2_M1004_g N_VGND_c_472_n 0.00459069f $X=2.785 $Y=0.745 $X2=0 $Y2=0
cc_176 N_A2_M1005_g N_VGND_c_472_n 0.00361512f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_177 N_A2_M1004_g N_VGND_c_476_n 0.00359326f $X=2.785 $Y=0.745 $X2=0 $Y2=0
cc_178 N_A2_M1005_g N_VGND_c_477_n 0.0035672f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_179 N_A2_M1004_g N_VGND_c_478_n 0.00558785f $X=2.785 $Y=0.745 $X2=0 $Y2=0
cc_180 N_A2_M1005_g N_VGND_c_478_n 0.00510388f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_181 N_A2_M1004_g N_A_489_65#_c_534_n 0.00683802f $X=2.785 $Y=0.745 $X2=0
+ $Y2=0
cc_182 N_A2_M1005_g N_A_489_65#_c_534_n 8.17594e-19 $X=3.375 $Y=0.745 $X2=0
+ $Y2=0
cc_183 N_A2_M1004_g N_A_489_65#_c_541_n 0.00956333f $X=2.785 $Y=0.745 $X2=0
+ $Y2=0
cc_184 N_A2_M1005_g N_A_489_65#_c_541_n 0.0102947f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_185 N_A2_M1004_g N_A_489_65#_c_535_n 7.15802e-19 $X=2.785 $Y=0.745 $X2=0
+ $Y2=0
cc_186 N_A2_M1004_g N_A_489_65#_c_544_n 7.93361e-19 $X=2.785 $Y=0.745 $X2=0
+ $Y2=0
cc_187 N_A2_M1005_g N_A_489_65#_c_544_n 0.00496189f $X=3.375 $Y=0.745 $X2=0
+ $Y2=0
cc_188 N_A2_M1005_g N_A_489_65#_c_537_n 0.0027743f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_189 N_A1_c_223_n N_Y_c_304_n 0.0127326f $X=3.805 $Y=1.275 $X2=0 $Y2=0
cc_190 N_A1_c_224_n N_Y_c_304_n 0.0082455f $X=4.315 $Y=1.275 $X2=0 $Y2=0
cc_191 N_A1_c_225_n N_Y_c_304_n 0.040635f $X=4.445 $Y=1.505 $X2=0 $Y2=0
cc_192 A1 N_Y_c_304_n 0.00276998f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_193 N_A1_c_227_n N_Y_c_304_n 0.00543694f $X=4.315 $Y=1.475 $X2=0 $Y2=0
cc_194 N_A1_c_224_n N_Y_c_338_n 0.00654168f $X=4.315 $Y=1.275 $X2=0 $Y2=0
cc_195 N_A1_M1003_g N_A_296_367#_c_364_n 0.0128633f $X=3.805 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A1_M1010_g N_A_296_367#_c_364_n 0.00221478f $X=4.235 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_A1_c_225_n N_A_296_367#_c_364_n 0.0287951f $X=4.445 $Y=1.505 $X2=0
+ $Y2=0
cc_198 N_A1_c_227_n N_A_296_367#_c_364_n 0.00266669f $X=4.315 $Y=1.475 $X2=0
+ $Y2=0
cc_199 N_A1_M1003_g N_VPWR_c_406_n 0.0140821f $X=3.805 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A1_M1010_g N_VPWR_c_406_n 7.24342e-19 $X=4.235 $Y=2.465 $X2=0 $Y2=0
cc_201 N_A1_M1003_g N_VPWR_c_408_n 7.72717e-19 $X=3.805 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A1_M1010_g N_VPWR_c_408_n 0.0205313f $X=4.235 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A1_c_225_n N_VPWR_c_408_n 0.00598826f $X=4.445 $Y=1.505 $X2=0 $Y2=0
cc_204 A1 N_VPWR_c_408_n 0.0152447f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_205 N_A1_c_227_n N_VPWR_c_408_n 0.00391249f $X=4.315 $Y=1.475 $X2=0 $Y2=0
cc_206 N_A1_M1003_g N_VPWR_c_411_n 0.00486043f $X=3.805 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A1_M1010_g N_VPWR_c_411_n 0.00486043f $X=4.235 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A1_M1003_g N_VPWR_c_404_n 0.00824727f $X=3.805 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A1_M1010_g N_VPWR_c_404_n 0.00824727f $X=4.235 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A1_c_223_n N_VGND_c_477_n 0.00302473f $X=3.805 $Y=1.275 $X2=0 $Y2=0
cc_211 N_A1_c_224_n N_VGND_c_477_n 0.00302501f $X=4.315 $Y=1.275 $X2=0 $Y2=0
cc_212 N_A1_c_223_n N_VGND_c_478_n 0.00443096f $X=3.805 $Y=1.275 $X2=0 $Y2=0
cc_213 N_A1_c_224_n N_VGND_c_478_n 0.00478352f $X=4.315 $Y=1.275 $X2=0 $Y2=0
cc_214 N_A1_c_223_n N_A_489_65#_c_541_n 0.0021345f $X=3.805 $Y=1.275 $X2=0 $Y2=0
cc_215 N_A1_c_223_n N_A_489_65#_c_544_n 0.00474233f $X=3.805 $Y=1.275 $X2=0
+ $Y2=0
cc_216 N_A1_c_224_n N_A_489_65#_c_544_n 5.37284e-19 $X=4.315 $Y=1.275 $X2=0
+ $Y2=0
cc_217 N_A1_c_223_n N_A_489_65#_c_536_n 0.00872289f $X=3.805 $Y=1.275 $X2=0
+ $Y2=0
cc_218 N_A1_c_224_n N_A_489_65#_c_536_n 0.0129928f $X=4.315 $Y=1.275 $X2=0 $Y2=0
cc_219 N_A1_c_223_n N_A_489_65#_c_537_n 0.00135267f $X=3.805 $Y=1.275 $X2=0
+ $Y2=0
cc_220 A1 N_A_489_65#_c_538_n 0.0224259f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_221 N_A1_c_227_n N_A_489_65#_c_538_n 0.00165222f $X=4.315 $Y=1.475 $X2=0
+ $Y2=0
cc_222 N_A_41_367#_c_277_n N_Y_M1008_d 0.00332344f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_223 N_A_41_367#_c_277_n N_Y_c_307_n 0.0159805f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_224 N_A_41_367#_c_279_n N_Y_c_303_n 3.99837e-19 $X=1.19 $Y=2.085 $X2=0 $Y2=0
cc_225 N_A_41_367#_c_273_n N_A_296_367#_M1001_s 0.00332344f $X=1.955 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_226 N_A_41_367#_c_273_n N_A_296_367#_c_366_n 0.0159805f $X=1.955 $Y=2.99
+ $X2=0 $Y2=0
cc_227 N_A_41_367#_M1009_d N_A_296_367#_c_363_n 0.00561813f $X=1.91 $Y=1.835
+ $X2=0 $Y2=0
cc_228 N_A_41_367#_c_274_n N_A_296_367#_c_363_n 0.0202165f $X=2.05 $Y=2.425
+ $X2=0 $Y2=0
cc_229 N_A_41_367#_c_273_n N_VPWR_c_405_n 0.00910673f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_230 N_A_41_367#_c_274_n N_VPWR_c_405_n 0.0319939f $X=2.05 $Y=2.425 $X2=0
+ $Y2=0
cc_231 N_A_41_367#_c_271_n N_VPWR_c_409_n 0.0179183f $X=0.295 $Y=2.905 $X2=0
+ $Y2=0
cc_232 N_A_41_367#_c_277_n N_VPWR_c_409_n 0.0361172f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_233 N_A_41_367#_c_273_n N_VPWR_c_409_n 0.0540354f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_234 N_A_41_367#_c_295_p N_VPWR_c_409_n 0.0125234f $X=1.19 $Y=2.91 $X2=0 $Y2=0
cc_235 N_A_41_367#_M1008_s N_VPWR_c_404_n 0.00215161f $X=0.205 $Y=1.835 $X2=0
+ $Y2=0
cc_236 N_A_41_367#_M1014_s N_VPWR_c_404_n 0.00223565f $X=1.05 $Y=1.835 $X2=0
+ $Y2=0
cc_237 N_A_41_367#_M1009_d N_VPWR_c_404_n 0.00215161f $X=1.91 $Y=1.835 $X2=0
+ $Y2=0
cc_238 N_A_41_367#_c_271_n N_VPWR_c_404_n 0.0101029f $X=0.295 $Y=2.905 $X2=0
+ $Y2=0
cc_239 N_A_41_367#_c_277_n N_VPWR_c_404_n 0.023676f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_240 N_A_41_367#_c_273_n N_VPWR_c_404_n 0.0337842f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_241 N_A_41_367#_c_295_p N_VPWR_c_404_n 0.00738676f $X=1.19 $Y=2.91 $X2=0
+ $Y2=0
cc_242 N_Y_c_304_n N_A_296_367#_c_363_n 0.00345671f $X=3.935 $Y=1.16 $X2=0 $Y2=0
cc_243 N_Y_c_304_n N_A_296_367#_c_364_n 0.00972247f $X=3.935 $Y=1.16 $X2=0 $Y2=0
cc_244 N_Y_M1008_d N_VPWR_c_404_n 0.00225186f $X=0.62 $Y=1.835 $X2=0 $Y2=0
cc_245 N_Y_c_303_n N_VGND_M1013_d 0.00176461f $X=1.525 $Y=1.16 $X2=0 $Y2=0
cc_246 N_Y_c_304_n N_VGND_M1011_s 0.00225342f $X=3.935 $Y=1.16 $X2=0 $Y2=0
cc_247 N_Y_c_304_n N_VGND_M1004_d 0.00386799f $X=3.935 $Y=1.16 $X2=0 $Y2=0
cc_248 N_Y_c_303_n N_VGND_c_470_n 0.0170777f $X=1.525 $Y=1.16 $X2=0 $Y2=0
cc_249 N_Y_c_304_n N_VGND_c_471_n 0.0202165f $X=3.935 $Y=1.16 $X2=0 $Y2=0
cc_250 N_Y_c_328_n N_VGND_c_473_n 0.0143246f $X=1.62 $Y=0.42 $X2=0 $Y2=0
cc_251 N_Y_c_306_n N_VGND_c_475_n 0.015688f $X=0.76 $Y=0.42 $X2=0 $Y2=0
cc_252 N_Y_M1012_s N_VGND_c_478_n 0.00380103f $X=0.62 $Y=0.245 $X2=0 $Y2=0
cc_253 N_Y_M1007_d N_VGND_c_478_n 0.00380103f $X=1.48 $Y=0.245 $X2=0 $Y2=0
cc_254 N_Y_c_306_n N_VGND_c_478_n 0.00984745f $X=0.76 $Y=0.42 $X2=0 $Y2=0
cc_255 N_Y_c_328_n N_VGND_c_478_n 0.00916141f $X=1.62 $Y=0.42 $X2=0 $Y2=0
cc_256 N_Y_c_304_n N_A_489_65#_M1004_s 0.00262981f $X=3.935 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_257 N_Y_c_304_n N_A_489_65#_M1005_s 0.00176461f $X=3.935 $Y=1.16 $X2=0 $Y2=0
cc_258 N_Y_c_304_n N_A_489_65#_c_541_n 0.0577223f $X=3.935 $Y=1.16 $X2=0 $Y2=0
cc_259 N_Y_c_304_n N_A_489_65#_c_535_n 0.0219393f $X=3.935 $Y=1.16 $X2=0 $Y2=0
cc_260 N_Y_M1002_s N_A_489_65#_c_536_n 0.00261503f $X=3.88 $Y=0.325 $X2=0 $Y2=0
cc_261 N_Y_c_304_n N_A_489_65#_c_536_n 0.00275981f $X=3.935 $Y=1.16 $X2=0 $Y2=0
cc_262 N_Y_c_338_n N_A_489_65#_c_536_n 0.0203258f $X=4.1 $Y=0.68 $X2=0 $Y2=0
cc_263 N_A_296_367#_c_363_n N_VPWR_M1000_d 0.00479121f $X=3.065 $Y=2.005
+ $X2=-0.19 $Y2=1.655
cc_264 N_A_296_367#_c_364_n N_VPWR_M1006_d 0.00176461f $X=3.925 $Y=1.85 $X2=0
+ $Y2=0
cc_265 N_A_296_367#_c_363_n N_VPWR_c_405_n 0.0220026f $X=3.065 $Y=2.005 $X2=0
+ $Y2=0
cc_266 N_A_296_367#_c_364_n N_VPWR_c_406_n 0.0170777f $X=3.925 $Y=1.85 $X2=0
+ $Y2=0
cc_267 N_A_296_367#_c_397_p N_VPWR_c_410_n 0.0124525f $X=3.16 $Y=2.455 $X2=0
+ $Y2=0
cc_268 N_A_296_367#_c_398_p N_VPWR_c_411_n 0.0124525f $X=4.02 $Y=1.98 $X2=0
+ $Y2=0
cc_269 N_A_296_367#_M1001_s N_VPWR_c_404_n 0.00225186f $X=1.48 $Y=1.835 $X2=0
+ $Y2=0
cc_270 N_A_296_367#_M1000_s N_VPWR_c_404_n 0.00536646f $X=3.02 $Y=1.835 $X2=0
+ $Y2=0
cc_271 N_A_296_367#_M1003_s N_VPWR_c_404_n 0.00536646f $X=3.88 $Y=1.835 $X2=0
+ $Y2=0
cc_272 N_A_296_367#_c_397_p N_VPWR_c_404_n 0.00730901f $X=3.16 $Y=2.455 $X2=0
+ $Y2=0
cc_273 N_A_296_367#_c_398_p N_VPWR_c_404_n 0.00730901f $X=4.02 $Y=1.98 $X2=0
+ $Y2=0
cc_274 N_VGND_c_471_n N_A_489_65#_c_534_n 0.0326659f $X=2.05 $Y=0.39 $X2=0 $Y2=0
cc_275 N_VGND_c_472_n N_A_489_65#_c_534_n 0.010078f $X=3.08 $Y=0.45 $X2=0 $Y2=0
cc_276 N_VGND_c_476_n N_A_489_65#_c_534_n 0.017603f $X=2.915 $Y=0 $X2=0 $Y2=0
cc_277 N_VGND_c_478_n N_A_489_65#_c_534_n 0.012271f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_M1004_d N_A_489_65#_c_541_n 0.00724401f $X=2.86 $Y=0.325 $X2=0
+ $Y2=0
cc_279 N_VGND_c_472_n N_A_489_65#_c_541_n 0.0255659f $X=3.08 $Y=0.45 $X2=0 $Y2=0
cc_280 N_VGND_c_476_n N_A_489_65#_c_541_n 0.00203769f $X=2.915 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_477_n N_A_489_65#_c_541_n 0.00203769f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_478_n N_A_489_65#_c_541_n 0.00957394f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_471_n N_A_489_65#_c_535_n 0.0137386f $X=2.05 $Y=0.39 $X2=0 $Y2=0
cc_284 N_VGND_c_477_n N_A_489_65#_c_536_n 0.0615871f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_478_n N_A_489_65#_c_536_n 0.0344158f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_472_n N_A_489_65#_c_537_n 0.00960644f $X=3.08 $Y=0.45 $X2=0
+ $Y2=0
cc_287 N_VGND_c_477_n N_A_489_65#_c_537_n 0.0234012f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_288 N_VGND_c_478_n N_A_489_65#_c_537_n 0.0125856f $X=4.56 $Y=0 $X2=0 $Y2=0
