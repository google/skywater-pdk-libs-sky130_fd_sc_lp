* File: sky130_fd_sc_lp__inputiso0p_lp.pex.spice
* Created: Wed Sep  2 09:55:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INPUTISO0P_LP%SLEEP 3 7 11 15 17 18 22
r34 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=1.465 $X2=0.71 $Y2=1.465
r35 18 23 6.14636 $w=3.73e-07 $l=2e-07 $layer=LI1_cond $X=0.732 $Y=1.665
+ $X2=0.732 $Y2=1.465
r36 17 23 5.22441 $w=3.73e-07 $l=1.7e-07 $layer=LI1_cond $X=0.732 $Y=1.295
+ $X2=0.732 $Y2=1.465
r37 13 22 100.035 $w=2.55e-07 $l=6.03324e-07 $layer=POLY_cond $X=0.845 $Y=1.985
+ $X2=0.665 $Y2=1.465
r38 13 15 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.845 $Y=1.985
+ $X2=0.845 $Y2=2.655
r39 9 22 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=0.845 $Y=1.3
+ $X2=0.665 $Y2=1.465
r40 9 11 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.845 $Y=1.3
+ $X2=0.845 $Y2=0.675
r41 5 22 100.035 $w=2.55e-07 $l=6.03324e-07 $layer=POLY_cond $X=0.485 $Y=1.985
+ $X2=0.665 $Y2=1.465
r42 5 7 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.485 $Y=1.985
+ $X2=0.485 $Y2=2.655
r43 1 22 32.933 $w=2.55e-07 $l=1.8e-07 $layer=POLY_cond $X=0.485 $Y=1.465
+ $X2=0.665 $Y2=1.465
r44 1 3 320.479 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.485 $Y=1.465
+ $X2=0.485 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0P_LP%A_27_93# 1 2 9 13 17 21 25 27 31 32 34
c55 27 0 7.5803e-20 $X=1.2 $Y=2.15
c56 13 0 4.20716e-20 $X=1.625 $Y=0.675
r57 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.43
+ $Y=1.475 $X2=1.43 $Y2=1.475
r58 29 31 17.2137 $w=3.93e-07 $l=5.9e-07 $layer=LI1_cond $X=1.397 $Y=2.065
+ $X2=1.397 $Y2=1.475
r59 28 34 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.375 $Y=2.15
+ $X2=0.265 $Y2=2.15
r60 27 29 8.32734 $w=1.7e-07 $l=2.35699e-07 $layer=LI1_cond $X=1.2 $Y=2.15
+ $X2=1.397 $Y2=2.065
r61 27 28 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.2 $Y=2.15
+ $X2=0.375 $Y2=2.15
r62 23 34 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.235
+ $X2=0.265 $Y2=2.15
r63 23 25 19.6439 $w=2.18e-07 $l=3.75e-07 $layer=LI1_cond $X=0.265 $Y=2.235
+ $X2=0.265 $Y2=2.61
r64 19 34 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.065
+ $X2=0.265 $Y2=2.15
r65 19 21 70.4562 $w=2.18e-07 $l=1.345e-06 $layer=LI1_cond $X=0.265 $Y=2.065
+ $X2=0.265 $Y2=0.72
r66 15 32 98.502 $w=2.54e-07 $l=5.93212e-07 $layer=POLY_cond $X=1.635 $Y=1.985
+ $X2=1.455 $Y2=1.475
r67 15 17 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.635 $Y=1.985
+ $X2=1.635 $Y2=2.655
r68 11 32 42.1589 $w=5.09e-07 $l=2.38642e-07 $layer=POLY_cond $X=1.625 $Y=1.31
+ $X2=1.455 $Y2=1.475
r69 11 13 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.625 $Y=1.31
+ $X2=1.625 $Y2=0.675
r70 7 32 98.502 $w=2.54e-07 $l=5.93212e-07 $layer=POLY_cond $X=1.275 $Y=1.985
+ $X2=1.455 $Y2=1.475
r71 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.275 $Y=1.985
+ $X2=1.275 $Y2=2.655
r72 2 25 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.445 $X2=0.27 $Y2=2.61
r73 1 21 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.27 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0P_LP%A 3 5 8 12 14 15 16 23 24
c46 24 0 1.49298e-19 $X=2.485 $Y=1.48
c47 8 0 7.5803e-20 $X=2.085 $Y=2.655
r48 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.485
+ $Y=1.48 $X2=2.485 $Y2=1.48
r49 21 23 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=2.445 $Y=1.48
+ $X2=2.485 $Y2=1.48
r50 20 21 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.085 $Y=1.48
+ $X2=2.445 $Y2=1.48
r51 18 20 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=2.055 $Y=1.48
+ $X2=2.085 $Y2=1.48
r52 16 24 3.3026 $w=6.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.315 $Y=1.665
+ $X2=2.315 $Y2=1.48
r53 14 15 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.02 $Y=0.995
+ $X2=2.02 $Y2=1.145
r54 10 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=1.645
+ $X2=2.445 $Y2=1.48
r55 10 12 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=2.445 $Y=1.645
+ $X2=2.445 $Y2=2.655
r56 6 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.085 $Y=1.645
+ $X2=2.085 $Y2=1.48
r57 6 8 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=2.085 $Y=1.645
+ $X2=2.085 $Y2=2.655
r58 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.055 $Y=1.315
+ $X2=2.055 $Y2=1.48
r59 5 15 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.055 $Y=1.315
+ $X2=2.055 $Y2=1.145
r60 3 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.985 $Y=0.675
+ $X2=1.985 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0P_LP%A_342_489# 1 2 7 9 12 14 16 19 23 25
+ 26 29 31 32 33 34 37
c68 29 0 4.20716e-20 $X=2.2 $Y=0.72
r69 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.06
+ $Y=1.17 $X2=3.06 $Y2=1.17
r70 33 36 2.67338 $w=4.1e-07 $l=1.1e-07 $layer=LI1_cond $X=3.025 $Y=1.225
+ $X2=3.025 $Y2=1.115
r71 33 34 20.5191 $w=4.08e-07 $l=7.3e-07 $layer=LI1_cond $X=3.025 $Y=1.225
+ $X2=3.025 $Y2=1.955
r72 31 36 4.98221 $w=2.2e-07 $l=2.05e-07 $layer=LI1_cond $X=2.82 $Y=1.115
+ $X2=3.025 $Y2=1.115
r73 31 32 26.9776 $w=2.18e-07 $l=5.15e-07 $layer=LI1_cond $X=2.82 $Y=1.115
+ $X2=2.305 $Y2=1.115
r74 27 32 6.82129 $w=2.2e-07 $l=1.53786e-07 $layer=LI1_cond $X=2.2 $Y=1.005
+ $X2=2.305 $Y2=1.115
r75 27 29 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.2 $Y=1.005
+ $X2=2.2 $Y2=0.72
r76 25 34 8.45803 $w=1.7e-07 $l=2.43824e-07 $layer=LI1_cond $X=2.82 $Y=2.04
+ $X2=3.025 $Y2=1.955
r77 25 26 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.82 $Y=2.04
+ $X2=1.975 $Y2=2.04
r78 21 26 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.87 $Y=2.125
+ $X2=1.975 $Y2=2.04
r79 21 23 25.6147 $w=2.08e-07 $l=4.85e-07 $layer=LI1_cond $X=1.87 $Y=2.125
+ $X2=1.87 $Y2=2.61
r80 17 37 99.0899 $w=2.55e-07 $l=5.98268e-07 $layer=POLY_cond $X=3.295 $Y=1.685
+ $X2=3.115 $Y2=1.17
r81 17 19 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.295 $Y=1.685
+ $X2=3.295 $Y2=2.465
r82 14 37 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=3.295 $Y=1.005
+ $X2=3.115 $Y2=1.17
r83 14 16 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.295 $Y=1.005
+ $X2=3.295 $Y2=0.675
r84 10 37 99.0899 $w=2.55e-07 $l=5.98268e-07 $layer=POLY_cond $X=2.935 $Y=1.685
+ $X2=3.115 $Y2=1.17
r85 10 12 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.935 $Y=1.685
+ $X2=2.935 $Y2=2.465
r86 7 37 32.933 $w=2.55e-07 $l=1.8e-07 $layer=POLY_cond $X=2.935 $Y=1.17
+ $X2=3.115 $Y2=1.17
r87 7 9 106.04 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.935 $Y=1.17
+ $X2=2.935 $Y2=0.675
r88 2 23 600 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.445 $X2=1.87 $Y2=2.61
r89 1 29 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.465 $X2=2.2 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0P_LP%VPWR 1 2 9 13 15 17 22 29 30 33 36
r44 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r48 27 36 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.91 $Y=3.33
+ $X2=2.717 $Y2=3.33
r49 27 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.91 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.06 $Y2=3.33
r53 23 25 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=1.225 $Y=3.33 $X2=2.16
+ $Y2=3.33
r54 22 36 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.717 $Y2=3.33
r55 22 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.06 $Y2=3.33
r59 17 19 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 11 36 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.717 $Y=3.245
+ $X2=2.717 $Y2=3.33
r63 11 13 25.8926 $w=3.83e-07 $l=8.65e-07 $layer=LI1_cond $X=2.717 $Y=3.245
+ $X2=2.717 $Y2=2.38
r64 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=3.245 $X2=1.06
+ $Y2=3.33
r65 7 9 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.06 $Y=3.245
+ $X2=1.06 $Y2=2.61
r66 2 13 300 $w=1.7e-07 $l=2.30217e-07 $layer=licon1_PDIFF $count=2 $X=2.52
+ $Y=2.445 $X2=2.72 $Y2=2.38
r67 1 9 600 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=0.92
+ $Y=2.445 $X2=1.06 $Y2=2.61
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0P_LP%X 1 2 7 8 9 10 11 18
r10 11 33 16.0693 $w=3.53e-07 $l=4.95e-07 $layer=LI1_cond $X=3.577 $Y=2.405
+ $X2=3.577 $Y2=2.9
r11 11 29 9.08969 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=3.577 $Y=2.405
+ $X2=3.577 $Y2=2.125
r12 10 29 2.92169 $w=3.53e-07 $l=9e-08 $layer=LI1_cond $X=3.577 $Y=2.035
+ $X2=3.577 $Y2=2.125
r13 9 10 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.577 $Y=1.665
+ $X2=3.577 $Y2=2.035
r14 8 9 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.577 $Y=1.295
+ $X2=3.577 $Y2=1.665
r15 7 8 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.577 $Y=0.925
+ $X2=3.577 $Y2=1.295
r16 7 18 6.65495 $w=3.53e-07 $l=2.05e-07 $layer=LI1_cond $X=3.577 $Y=0.925
+ $X2=3.577 $Y2=0.72
r17 2 33 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=1.835 $X2=3.51 $Y2=2.9
r18 2 29 400 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=1.835 $X2=3.51 $Y2=2.125
r19 1 18 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.465 $X2=3.51 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0P_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 27 36 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.717
+ $Y2=0
r46 27 29 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.6
+ $Y2=0
r47 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r49 23 33 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.235
+ $Y2=0
r50 23 25 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=2.16
+ $Y2=0
r51 22 36 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.717
+ $Y2=0
r52 22 25 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.16
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r54 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 17 33 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.235
+ $Y2=0
r56 17 19 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.72
+ $Y2=0
r57 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r58 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r59 11 36 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.717 $Y=0.085
+ $X2=2.717 $Y2=0
r60 11 13 21.8448 $w=3.33e-07 $l=6.35e-07 $layer=LI1_cond $X=2.717 $Y=0.085
+ $X2=2.717 $Y2=0.72
r61 7 33 2.80049 $w=6.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r62 7 9 10.3777 $w=6.78e-07 $l=5.9e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.675
r63 2 13 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.465 $X2=2.72 $Y2=0.72
r64 1 9 91 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=2 $X=0.92
+ $Y=0.465 $X2=1.41 $Y2=0.675
.ends

