* File: sky130_fd_sc_lp__dlrbp_1.pex.spice
* Created: Wed Sep  2 09:46:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRBP_1%GATE 3 5 8 10 11 12 16 17 18
c32 18 0 1.30066e-19 $X=0.697 $Y=0.995
r33 16 18 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.697 $Y=1.16
+ $X2=0.697 $Y2=0.995
r34 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.72
+ $Y=1.16 $X2=0.72 $Y2=1.16
r35 11 12 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.755 $Y=1.295
+ $X2=0.755 $Y2=1.665
r36 11 17 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.755 $Y=1.295
+ $X2=0.755 $Y2=1.16
r37 8 10 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=0.585 $Y=2.735
+ $X2=0.585 $Y2=1.665
r38 5 10 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.697 $Y=1.478
+ $X2=0.697 $Y2=1.665
r39 4 16 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.697 $Y=1.182
+ $X2=0.697 $Y2=1.16
r40 4 5 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.697 $Y=1.182
+ $X2=0.697 $Y2=1.478
r41 3 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.585 $Y=0.675
+ $X2=0.585 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%D 2 5 9 11 12 13 17
r48 17 19 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=2.167 $Y=1.615
+ $X2=2.167 $Y2=1.45
r49 12 13 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=2.205 $Y=1.615
+ $X2=2.205 $Y2=2.035
r50 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.16
+ $Y=1.615 $X2=2.16 $Y2=1.615
r51 9 19 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.265 $Y=0.805
+ $X2=2.265 $Y2=1.45
r52 5 11 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=2.205 $Y=2.725
+ $X2=2.205 $Y2=2.12
r53 2 11 40.4609 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=2.167 $Y=1.948
+ $X2=2.167 $Y2=2.12
r54 1 17 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=2.167 $Y=1.622
+ $X2=2.167 $Y2=1.615
r55 1 2 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=2.167 $Y=1.622
+ $X2=2.167 $Y2=1.948
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%A_373_481# 1 2 7 8 11 15 19 22 24 28 29 34
+ 38
r80 35 38 5.92685 $w=3.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.81 $Y=2.56
+ $X2=1.99 $Y2=2.56
r81 29 42 23.9404 $w=3.02e-07 $l=1.5e-07 $layer=POLY_cond $X=2.755 $Y=1.86
+ $X2=2.905 $Y2=1.86
r82 29 40 11.9702 $w=3.02e-07 $l=7.5e-08 $layer=POLY_cond $X=2.755 $Y=1.86
+ $X2=2.68 $Y2=1.86
r83 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.755
+ $Y=1.86 $X2=2.755 $Y2=1.86
r84 26 28 26.7367 $w=2.48e-07 $l=5.8e-07 $layer=LI1_cond $X=2.715 $Y=1.28
+ $X2=2.715 $Y2=1.86
r85 24 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.59 $Y=1.195
+ $X2=2.715 $Y2=1.28
r86 24 34 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.59 $Y=1.195
+ $X2=2.18 $Y2=1.195
r87 20 34 8.62937 $w=1.93e-07 $l=1.48e-07 $layer=LI1_cond $X=2.032 $Y=1.182
+ $X2=2.18 $Y2=1.182
r88 20 31 12.6266 $w=1.93e-07 $l=2.22e-07 $layer=LI1_cond $X=2.032 $Y=1.182
+ $X2=1.81 $Y2=1.182
r89 20 22 10.9384 $w=2.93e-07 $l=2.8e-07 $layer=LI1_cond $X=2.032 $Y=1.085
+ $X2=2.032 $Y2=0.805
r90 19 35 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.81 $Y=2.385 $X2=1.81
+ $Y2=2.56
r91 18 31 1.54022 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.81 $Y=1.28 $X2=1.81
+ $Y2=1.182
r92 18 19 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=1.81 $Y=1.28
+ $X2=1.81 $Y2=2.385
r93 13 42 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=2.025
+ $X2=2.905 $Y2=1.86
r94 13 15 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=2.905 $Y=2.025
+ $X2=2.905 $Y2=2.725
r95 11 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.695 $Y=0.805
+ $X2=2.695 $Y2=1.355
r96 8 40 14.8734 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.695
+ $X2=2.68 $Y2=1.86
r97 7 17 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.68 $Y=1.445 $X2=2.68
+ $Y2=1.355
r98 7 8 97.1774 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=2.68 $Y=1.445 $X2=2.68
+ $Y2=1.695
r99 2 38 600 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=2.405 $X2=1.99 $Y2=2.57
r100 1 22 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.595 $X2=2.05 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%A_218_483# 1 2 9 12 16 19 20 21 23 25 26 27
+ 30 31 34 35 39 43 44 47 49
c129 39 0 1.30066e-19 $X=1.385 $Y=0.675
c130 30 0 3.47362e-20 $X=3.93 $Y=2.3
c131 16 0 4.98098e-20 $X=2.255 $Y=2.99
c132 12 0 1.48731e-20 $X=3.79 $Y=2.835
r133 44 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.29
+ $X2=3.145 $Y2=1.125
r134 43 46 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=1.29
+ $X2=3.135 $Y2=1.455
r135 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.145
+ $Y=1.29 $X2=3.145 $Y2=1.29
r136 39 41 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0.675
+ $X2=1.385 $Y2=0.84
r137 35 41 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=1.46 $Y=2.425
+ $X2=1.46 $Y2=0.84
r138 34 36 10.7149 $w=4.78e-07 $l=4.3e-07 $layer=LI1_cond $X=1.305 $Y=2.56
+ $X2=1.305 $Y2=2.99
r139 34 35 8.64879 $w=4.78e-07 $l=1.35e-07 $layer=LI1_cond $X=1.305 $Y=2.56
+ $X2=1.305 $Y2=2.425
r140 31 51 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.93 $Y=2.3
+ $X2=3.79 $Y2=2.3
r141 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=2.3 $X2=3.93 $Y2=2.3
r142 28 30 26.8165 $w=2.58e-07 $l=6.05e-07 $layer=LI1_cond $X=3.885 $Y=2.905
+ $X2=3.885 $Y2=2.3
r143 26 28 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.755 $Y=2.99
+ $X2=3.885 $Y2=2.905
r144 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.755 $Y=2.99
+ $X2=3.195 $Y2=2.99
r145 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.11 $Y=2.905
+ $X2=3.195 $Y2=2.99
r146 24 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=2.46
+ $X2=3.11 $Y2=2.375
r147 24 25 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.11 $Y=2.46
+ $X2=3.11 $Y2=2.905
r148 23 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=2.29
+ $X2=3.11 $Y2=2.375
r149 23 46 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=3.11 $Y=2.29
+ $X2=3.11 $Y2=1.455
r150 20 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.025 $Y=2.375
+ $X2=3.11 $Y2=2.375
r151 20 21 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.025 $Y=2.375
+ $X2=2.425 $Y2=2.375
r152 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.34 $Y=2.46
+ $X2=2.425 $Y2=2.375
r153 18 19 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.34 $Y=2.46
+ $X2=2.34 $Y2=2.905
r154 17 36 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1.545 $Y=2.99
+ $X2=1.305 $Y2=2.99
r155 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.255 $Y=2.99
+ $X2=2.34 $Y2=2.905
r156 16 17 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.255 $Y=2.99
+ $X2=1.545 $Y2=2.99
r157 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=2.465
+ $X2=3.79 $Y2=2.3
r158 10 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.79 $Y=2.465
+ $X2=3.79 $Y2=2.835
r159 9 49 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.055 $Y=0.805
+ $X2=3.055 $Y2=1.125
r160 2 34 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.09
+ $Y=2.415 $X2=1.23 $Y2=2.56
r161 1 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.245
+ $Y=0.465 $X2=1.385 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%A_49_93# 1 2 9 11 13 15 16 19 20 21 24 26 27
+ 31 32 34 37 41 45 48 52
c113 24 0 1.74571e-19 $X=3.265 $Y=2.725
c114 9 0 4.98098e-20 $X=1.015 $Y=2.735
r115 45 47 5.94304 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.37 $Y=0.675
+ $X2=0.37 $Y2=0.825
r116 42 52 21.3331 $w=3.3e-07 $l=1.22e-07 $layer=POLY_cond $X=1.105 $Y=2.09
+ $X2=1.227 $Y2=2.09
r117 42 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.105 $Y=2.09
+ $X2=1.015 $Y2=2.09
r118 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=2.09 $X2=1.105 $Y2=2.09
r119 39 48 0.663103 $w=3.3e-07 $l=1.48e-07 $layer=LI1_cond $X=0.5 $Y=2.09
+ $X2=0.352 $Y2=2.09
r120 39 41 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=0.5 $Y=2.09
+ $X2=1.105 $Y2=2.09
r121 35 48 6.03966 $w=2.72e-07 $l=1.65e-07 $layer=LI1_cond $X=0.352 $Y=2.255
+ $X2=0.352 $Y2=2.09
r122 35 37 11.9151 $w=2.93e-07 $l=3.05e-07 $layer=LI1_cond $X=0.352 $Y=2.255
+ $X2=0.352 $Y2=2.56
r123 34 48 6.03966 $w=2.72e-07 $l=1.75656e-07 $layer=LI1_cond $X=0.33 $Y=1.925
+ $X2=0.352 $Y2=2.09
r124 34 47 50.7075 $w=2.48e-07 $l=1.1e-06 $layer=LI1_cond $X=0.33 $Y=1.925
+ $X2=0.33 $Y2=0.825
r125 29 31 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.595 $Y=1.745
+ $X2=3.595 $Y2=0.805
r126 28 31 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.595 $Y=0.255
+ $X2=3.595 $Y2=0.805
r127 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.52 $Y=1.82
+ $X2=3.595 $Y2=1.745
r128 26 27 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.52 $Y=1.82
+ $X2=3.34 $Y2=1.82
r129 22 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.265 $Y=1.895
+ $X2=3.34 $Y2=1.82
r130 22 24 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.265 $Y=1.895
+ $X2=3.265 $Y2=2.725
r131 20 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.52 $Y=0.18
+ $X2=3.595 $Y2=0.255
r132 20 21 856.319 $w=1.5e-07 $l=1.67e-06 $layer=POLY_cond $X=3.52 $Y=0.18
+ $X2=1.85 $Y2=0.18
r133 18 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.775 $Y=0.255
+ $X2=1.85 $Y2=0.18
r134 18 19 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.775 $Y=0.255
+ $X2=1.775 $Y2=0.995
r135 17 32 10.0082 $w=1.5e-07 $l=1.33e-07 $layer=POLY_cond $X=1.36 $Y=1.07
+ $X2=1.227 $Y2=1.07
r136 16 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.7 $Y=1.07
+ $X2=1.775 $Y2=0.995
r137 16 17 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.7 $Y=1.07 $X2=1.36
+ $Y2=1.07
r138 15 52 8.07087 $w=2.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.227 $Y=1.925
+ $X2=1.227 $Y2=2.09
r139 14 32 15.4588 $w=2.07e-07 $l=7.5e-08 $layer=POLY_cond $X=1.227 $Y=1.145
+ $X2=1.227 $Y2=1.07
r140 14 15 176.565 $w=2.65e-07 $l=7.8e-07 $layer=POLY_cond $X=1.227 $Y=1.145
+ $X2=1.227 $Y2=1.925
r141 11 32 15.4588 $w=2.07e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.17 $Y=0.995
+ $X2=1.227 $Y2=1.07
r142 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.17 $Y=0.995
+ $X2=1.17 $Y2=0.675
r143 7 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=2.255
+ $X2=1.015 $Y2=2.09
r144 7 9 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.015 $Y=2.255
+ $X2=1.015 $Y2=2.735
r145 2 37 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=2.415 $X2=0.37 $Y2=2.56
r146 1 45 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.465 $X2=0.37 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%A_776_93# 1 2 9 13 17 21 25 29 32 35 38 39
+ 42 43 44 47 49 50 53 56 58 59 62 63 65 69 70 72 76 77 84
c199 69 0 1.22982e-19 $X=5.945 $Y=1.46
c200 49 0 3.9997e-20 $X=5.64 $Y=0.74
c201 44 0 1.48731e-20 $X=4.355 $Y=2.385
c202 35 0 3.47362e-20 $X=4.22 $Y=1.925
c203 17 0 7.43952e-20 $X=5.86 $Y=0.865
r204 77 85 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=1.395
+ $X2=7.572 $Y2=1.56
r205 77 84 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=1.395
+ $X2=7.572 $Y2=1.23
r206 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.55
+ $Y=1.395 $X2=7.55 $Y2=1.395
r207 73 76 7.4385 $w=3.28e-07 $l=2.13e-07 $layer=LI1_cond $X=7.337 $Y=1.395
+ $X2=7.55 $Y2=1.395
r208 70 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.945 $Y=1.46
+ $X2=5.945 $Y2=1.625
r209 70 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.945 $Y=1.46
+ $X2=5.945 $Y2=1.295
r210 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.945
+ $Y=1.46 $X2=5.945 $Y2=1.46
r211 66 69 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=5.725 $Y=1.46
+ $X2=5.945 $Y2=1.46
r212 61 73 2.99809 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=7.337 $Y=1.56
+ $X2=7.337 $Y2=1.395
r213 61 62 39.1831 $w=2.23e-07 $l=7.65e-07 $layer=LI1_cond $X=7.337 $Y=1.56
+ $X2=7.337 $Y2=2.325
r214 60 72 4.86787 $w=1.82e-07 $l=9.12688e-08 $layer=LI1_cond $X=5.81 $Y=2.41
+ $X2=5.725 $Y2=2.397
r215 59 62 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=7.225 $Y=2.41
+ $X2=7.337 $Y2=2.325
r216 59 60 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=7.225 $Y=2.41
+ $X2=5.81 $Y2=2.41
r217 58 72 1.59926 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=5.725 $Y=2.3
+ $X2=5.725 $Y2=2.397
r218 57 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=1.625
+ $X2=5.725 $Y2=1.46
r219 57 58 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.725 $Y=1.625
+ $X2=5.725 $Y2=2.3
r220 56 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=1.295
+ $X2=5.725 $Y2=1.46
r221 55 56 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.725 $Y=0.825
+ $X2=5.725 $Y2=1.295
r222 54 65 6.0176 $w=1.82e-07 $l=1.1e-07 $layer=LI1_cond $X=5.215 $Y=2.397
+ $X2=5.105 $Y2=2.397
r223 53 72 4.86787 $w=1.82e-07 $l=8.5e-08 $layer=LI1_cond $X=5.64 $Y=2.397
+ $X2=5.725 $Y2=2.397
r224 53 54 24.1725 $w=1.93e-07 $l=4.25e-07 $layer=LI1_cond $X=5.64 $Y=2.397
+ $X2=5.215 $Y2=2.397
r225 49 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.64 $Y=0.74
+ $X2=5.725 $Y2=0.825
r226 49 50 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.64 $Y=0.74
+ $X2=4.875 $Y2=0.74
r227 45 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.71 $Y=0.655
+ $X2=4.875 $Y2=0.74
r228 45 47 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.71 $Y=0.655
+ $X2=4.71 $Y2=0.38
r229 43 65 6.0176 $w=1.82e-07 $l=1.15845e-07 $layer=LI1_cond $X=4.995 $Y=2.385
+ $X2=5.105 $Y2=2.397
r230 43 44 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.995 $Y=2.385
+ $X2=4.355 $Y2=2.385
r231 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.27 $Y=2.3
+ $X2=4.355 $Y2=2.385
r232 42 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.27 $Y=2.3
+ $X2=4.27 $Y2=1.925
r233 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.15
+ $Y=1.42 $X2=4.15 $Y2=1.42
r234 36 63 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.17 $Y=1.74
+ $X2=4.17 $Y2=1.925
r235 36 38 9.96707 $w=3.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.17 $Y=1.74
+ $X2=4.17 $Y2=1.42
r236 34 39 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.15 $Y=1.775
+ $X2=4.15 $Y2=1.42
r237 34 35 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.22 $Y=1.775
+ $X2=4.22 $Y2=1.925
r238 32 39 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.15 $Y=1.405
+ $X2=4.15 $Y2=1.42
r239 31 32 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.097 $Y=1.255
+ $X2=4.097 $Y2=1.405
r240 29 84 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.545 $Y=0.7
+ $X2=7.545 $Y2=1.23
r241 25 85 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=7.5 $Y=2.465
+ $X2=7.5 $Y2=1.56
r242 21 82 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.86 $Y=2.105
+ $X2=5.86 $Y2=1.625
r243 17 81 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.86 $Y=0.865
+ $X2=5.86 $Y2=1.295
r244 13 35 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.38 $Y=2.835
+ $X2=4.38 $Y2=1.925
r245 9 31 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.955 $Y=0.805
+ $X2=3.955 $Y2=1.255
r246 2 65 300 $w=1.7e-07 $l=7.46726e-07 $layer=licon1_PDIFF $count=2 $X=4.98
+ $Y=1.785 $X2=5.12 $Y2=2.465
r247 1 47 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.585
+ $Y=0.235 $X2=4.71 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%A_626_119# 1 2 9 11 13 14 16 20 27 28 31
c79 27 0 1.74571e-19 $X=3.48 $Y=2.57
c80 20 0 2.83637e-19 $X=4.69 $Y=1.35
r81 31 32 2.99379 $w=3.22e-07 $l=2e-08 $layer=POLY_cond $X=4.905 $Y=1.35
+ $X2=4.925 $Y2=1.35
r82 27 28 10.3163 $w=2.18e-07 $l=1.85e-07 $layer=LI1_cond $X=3.475 $Y=2.57
+ $X2=3.475 $Y2=2.385
r83 21 31 32.1832 $w=3.22e-07 $l=2.15e-07 $layer=POLY_cond $X=4.69 $Y=1.35
+ $X2=4.905 $Y2=1.35
r84 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.69
+ $Y=1.35 $X2=4.69 $Y2=1.35
r85 18 20 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=4.65 $Y=1.165
+ $X2=4.65 $Y2=1.35
r86 17 24 10.5759 $w=3.23e-07 $l=3.71537e-07 $layer=LI1_cond $X=3.585 $Y=1.08
+ $X2=3.372 $Y2=0.8
r87 16 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.525 $Y=1.08
+ $X2=4.65 $Y2=1.165
r88 16 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.525 $Y=1.08
+ $X2=3.585 $Y2=1.08
r89 14 17 5.9342 $w=3.23e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.5 $Y=1.165
+ $X2=3.585 $Y2=1.08
r90 14 28 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=3.5 $Y=1.165
+ $X2=3.5 $Y2=2.385
r91 11 32 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.925 $Y=1.185
+ $X2=4.925 $Y2=1.35
r92 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.925 $Y=1.185
+ $X2=4.925 $Y2=0.655
r93 7 31 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=1.515
+ $X2=4.905 $Y2=1.35
r94 7 9 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=4.905 $Y=1.515 $X2=4.905
+ $Y2=2.415
r95 2 27 600 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.405 $X2=3.48 $Y2=2.57
r96 1 24 182 $w=1.7e-07 $l=2.86356e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.595 $X2=3.325 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%RESET_B 3 7 9 10 11 16
c47 16 0 1.8139e-19 $X=5.375 $Y=1.375
c48 9 0 7.43952e-20 $X=5.04 $Y=1.295
c49 3 0 1.02248e-19 $X=5.285 $Y=0.655
r50 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.375 $Y=1.375
+ $X2=5.375 $Y2=1.54
r51 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.375 $Y=1.375
+ $X2=5.375 $Y2=1.21
r52 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.375
+ $Y=1.375 $X2=5.375 $Y2=1.375
r53 10 11 8.42951 $w=5.23e-07 $l=3.7e-07 $layer=LI1_cond $X=5.207 $Y=1.665
+ $X2=5.207 $Y2=2.035
r54 10 17 6.60691 $w=5.23e-07 $l=2.9e-07 $layer=LI1_cond $X=5.207 $Y=1.665
+ $X2=5.207 $Y2=1.375
r55 9 17 1.8226 $w=5.23e-07 $l=8e-08 $layer=LI1_cond $X=5.207 $Y=1.295 $X2=5.207
+ $Y2=1.375
r56 7 19 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=5.335 $Y=2.415
+ $X2=5.335 $Y2=1.54
r57 3 18 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.285 $Y=0.655
+ $X2=5.285 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%A_1187_131# 1 2 7 8 11 15 18 20 22 28 29 34
+ 36
c55 29 0 3.9997e-20 $X=6.485 $Y=0.93
c56 8 0 1.22982e-19 $X=6.65 $Y=1.36
r57 32 34 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.075 $Y=1.97
+ $X2=6.295 $Y2=1.97
r58 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.485
+ $Y=0.93 $X2=6.485 $Y2=0.93
r59 26 28 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.395 $Y=0.87
+ $X2=6.485 $Y2=0.87
r60 24 26 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6.075 $Y=0.87
+ $X2=6.395 $Y2=0.87
r61 22 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=1.805
+ $X2=6.295 $Y2=1.97
r62 22 36 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.295 $Y=1.805
+ $X2=6.295 $Y2=1.435
r63 20 36 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.395 $Y=1.25
+ $X2=6.395 $Y2=1.435
r64 19 26 0.0060886 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=1.035
+ $X2=6.395 $Y2=0.87
r65 19 20 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.395 $Y=1.035
+ $X2=6.395 $Y2=1.25
r66 17 29 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=6.485 $Y=1.285
+ $X2=6.485 $Y2=0.93
r67 13 18 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.1 $Y=1.285
+ $X2=7.085 $Y2=1.36
r68 13 15 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=7.1 $Y=1.285
+ $X2=7.1 $Y2=0.7
r69 9 18 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.07 $Y=1.435
+ $X2=7.085 $Y2=1.36
r70 9 11 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=7.07 $Y=1.435
+ $X2=7.07 $Y2=2.465
r71 8 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.65 $Y=1.36
+ $X2=6.485 $Y2=1.285
r72 7 18 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.995 $Y=1.36 $X2=7.085
+ $Y2=1.36
r73 7 8 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.995 $Y=1.36
+ $X2=6.65 $Y2=1.36
r74 2 32 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=5.935
+ $Y=1.785 $X2=6.075 $Y2=1.97
r75 1 24 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=5.935
+ $Y=0.655 $X2=6.075 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%VPWR 1 2 3 4 5 20 24 28 32 36 39 40 41 43 48
+ 53 66 67 70 73 76 79
r99 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r100 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r101 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r104 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r105 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r106 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r107 61 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r108 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r109 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r110 58 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.715 $Y=3.33
+ $X2=5.55 $Y2=3.33
r111 58 60 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.715 $Y=3.33
+ $X2=6 $Y2=3.33
r112 57 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r113 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r115 54 76 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.825 $Y=3.33
+ $X2=4.675 $Y2=3.33
r116 54 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.825 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.385 $Y=3.33
+ $X2=5.55 $Y2=3.33
r118 53 56 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.385 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r121 49 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.725 $Y2=3.33
r122 49 51 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.12 $Y2=3.33
r123 48 76 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.675 $Y2=3.33
r124 48 51 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 47 74 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r126 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 44 70 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.782 $Y2=3.33
r129 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 43 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=2.725 $Y2=3.33
r131 43 46 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 41 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r133 41 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r134 39 63 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.12 $Y=3.33
+ $X2=6.96 $Y2=3.33
r135 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.12 $Y=3.33
+ $X2=7.285 $Y2=3.33
r136 38 66 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=7.45 $Y=3.33
+ $X2=7.92 $Y2=3.33
r137 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=3.33
+ $X2=7.285 $Y2=3.33
r138 34 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.285 $Y=3.245
+ $X2=7.285 $Y2=3.33
r139 34 36 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=7.285 $Y=3.245
+ $X2=7.285 $Y2=2.79
r140 30 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=3.245
+ $X2=5.55 $Y2=3.33
r141 30 32 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.55 $Y=3.245
+ $X2=5.55 $Y2=2.75
r142 26 76 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.675 $Y=3.245
+ $X2=4.675 $Y2=3.33
r143 26 28 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=4.675 $Y=3.245
+ $X2=4.675 $Y2=2.805
r144 22 73 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=3.33
r145 22 24 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=2.795
r146 18 70 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.782 $Y=3.245
+ $X2=0.782 $Y2=3.33
r147 18 20 33.5489 $w=2.23e-07 $l=6.55e-07 $layer=LI1_cond $X=0.782 $Y=3.245
+ $X2=0.782 $Y2=2.59
r148 5 36 600 $w=1.7e-07 $l=1.02261e-06 $layer=licon1_PDIFF $count=1 $X=7.145
+ $Y=1.835 $X2=7.285 $Y2=2.79
r149 4 32 600 $w=1.7e-07 $l=1.03263e-06 $layer=licon1_PDIFF $count=1 $X=5.41
+ $Y=1.785 $X2=5.55 $Y2=2.75
r150 3 28 600 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=2.625 $X2=4.69 $Y2=2.805
r151 2 24 600 $w=1.7e-07 $l=5.72713e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=2.405 $X2=2.69 $Y2=2.795
r152 1 20 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=0.66
+ $Y=2.415 $X2=0.8 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%Q_N 1 2 7 8 9 10 11 18
r22 11 29 1.70033 $w=3.03e-07 $l=4.5e-08 $layer=LI1_cond $X=6.902 $Y=2.035
+ $X2=6.902 $Y2=1.99
r23 10 29 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=6.902 $Y=1.665
+ $X2=6.902 $Y2=1.99
r24 9 10 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=6.902 $Y=1.295
+ $X2=6.902 $Y2=1.665
r25 8 9 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=6.902 $Y=0.925
+ $X2=6.902 $Y2=1.295
r26 7 8 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=6.902 $Y=0.555
+ $X2=6.902 $Y2=0.925
r27 7 18 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=6.902 $Y=0.555
+ $X2=6.902 $Y2=0.425
r28 2 29 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.835 $X2=6.855 $Y2=1.99
r29 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.76
+ $Y=0.28 $X2=6.885 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%Q 1 2 7 8 9 10 11 12 13 25 35 38 40
r25 38 40 1.44581 $w=4.53e-07 $l=5.5e-08 $layer=LI1_cond $X=7.847 $Y=1.98
+ $X2=7.847 $Y2=2.035
r26 36 38 0.341737 $w=4.53e-07 $l=1.3e-08 $layer=LI1_cond $X=7.847 $Y=1.967
+ $X2=7.847 $Y2=1.98
r27 35 53 3.32435 $w=2.58e-07 $l=7.5e-08 $layer=LI1_cond $X=7.945 $Y=1.665
+ $X2=7.945 $Y2=1.74
r28 13 47 3.5488 $w=4.53e-07 $l=1.35e-07 $layer=LI1_cond $X=7.847 $Y=2.775
+ $X2=7.847 $Y2=2.91
r29 12 13 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=7.847 $Y=2.405
+ $X2=7.847 $Y2=2.775
r30 11 36 0.236587 $w=4.53e-07 $l=9e-09 $layer=LI1_cond $X=7.847 $Y=1.958
+ $X2=7.847 $Y2=1.967
r31 11 12 9.51605 $w=4.53e-07 $l=3.62e-07 $layer=LI1_cond $X=7.847 $Y=2.043
+ $X2=7.847 $Y2=2.405
r32 11 40 0.210299 $w=4.53e-07 $l=8e-09 $layer=LI1_cond $X=7.847 $Y=2.043
+ $X2=7.847 $Y2=2.035
r33 10 11 5.59922 $w=4.53e-07 $l=2.13e-07 $layer=LI1_cond $X=7.847 $Y=1.745
+ $X2=7.847 $Y2=1.958
r34 10 53 2.30998 $w=4.53e-07 $l=5e-09 $layer=LI1_cond $X=7.847 $Y=1.745
+ $X2=7.847 $Y2=1.74
r35 10 35 0.221624 $w=2.58e-07 $l=5e-09 $layer=LI1_cond $X=7.945 $Y=1.66
+ $X2=7.945 $Y2=1.665
r36 9 10 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=7.945 $Y=1.295
+ $X2=7.945 $Y2=1.66
r37 9 51 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=7.945 $Y=1.295
+ $X2=7.945 $Y2=1.06
r38 8 51 5.80516 $w=4.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.84 $Y=0.925
+ $X2=7.84 $Y2=1.06
r39 8 23 2.54485 $w=4.68e-07 $l=1e-07 $layer=LI1_cond $X=7.84 $Y=0.925 $X2=7.84
+ $Y2=0.825
r40 7 23 6.87109 $w=4.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.84 $Y=0.555
+ $X2=7.84 $Y2=0.825
r41 7 25 3.3083 $w=4.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.84 $Y=0.555 $X2=7.84
+ $Y2=0.425
r42 2 47 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.575
+ $Y=1.835 $X2=7.715 $Y2=2.91
r43 2 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.575
+ $Y=1.835 $X2=7.715 $Y2=1.98
r44 1 25 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=7.62
+ $Y=0.28 $X2=7.77 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_1%VGND 1 2 3 4 5 20 24 26 30 34 38 41 42 43 45
+ 53 66 67 70 73 76 79
r94 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r95 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r96 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r98 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r99 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r100 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r101 61 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r102 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r103 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r104 58 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=5.5
+ $Y2=0
r105 58 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=6
+ $Y2=0
r106 57 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r107 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r108 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.17
+ $Y2=0
r109 54 56 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=5.04 $Y2=0
r110 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.5
+ $Y2=0
r111 53 56 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.04
+ $Y2=0
r112 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r113 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r114 49 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r115 49 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r116 48 51 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r117 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r118 46 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.88
+ $Y2=0
r119 46 48 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.2
+ $Y2=0
r120 45 73 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.497
+ $Y2=0
r121 45 51 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.16
+ $Y2=0
r122 43 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r123 43 74 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r124 43 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r125 41 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.225 $Y=0
+ $X2=6.96 $Y2=0
r126 41 42 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.225 $Y=0 $X2=7.33
+ $Y2=0
r127 40 66 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=7.435 $Y=0
+ $X2=7.92 $Y2=0
r128 40 42 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.435 $Y=0 $X2=7.33
+ $Y2=0
r129 36 42 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=0.085
+ $X2=7.33 $Y2=0
r130 36 38 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=7.33 $Y=0.085
+ $X2=7.33 $Y2=0.425
r131 32 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=0.085 $X2=5.5
+ $Y2=0
r132 32 34 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.5 $Y=0.085
+ $X2=5.5 $Y2=0.4
r133 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0
r134 28 30 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0.74
r135 27 73 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.645 $Y=0
+ $X2=2.497 $Y2=0
r136 26 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.17
+ $Y2=0
r137 26 27 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.005 $Y=0
+ $X2=2.645 $Y2=0
r138 22 73 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.497 $Y=0.085
+ $X2=2.497 $Y2=0
r139 22 24 26.9554 $w=2.93e-07 $l=6.9e-07 $layer=LI1_cond $X=2.497 $Y=0.085
+ $X2=2.497 $Y2=0.775
r140 18 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=0.085
+ $X2=0.88 $Y2=0
r141 18 20 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.88 $Y=0.085
+ $X2=0.88 $Y2=0.675
r142 5 38 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=7.175
+ $Y=0.28 $X2=7.33 $Y2=0.425
r143 4 34 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.36
+ $Y=0.235 $X2=5.5 $Y2=0.4
r144 3 30 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.595 $X2=4.17 $Y2=0.74
r145 2 24 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.34
+ $Y=0.595 $X2=2.48 $Y2=0.775
r146 1 20 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.465 $X2=0.88 $Y2=0.675
.ends

