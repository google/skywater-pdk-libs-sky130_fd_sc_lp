* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4_lp A B C D VGND VNB VPB VPWR X
X0 a_720_55# a_186_485# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND D a_230_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_186_485# a_720_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_422_55# A a_186_485# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_114_485# D a_186_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_186_485# A a_588_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_430_485# B a_186_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR D a_114_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_230_55# C a_308_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_308_55# B a_422_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_186_485# C a_272_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_272_485# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VPWR a_186_485# a_746_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_588_485# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_746_485# a_186_485# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VPWR B a_430_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
