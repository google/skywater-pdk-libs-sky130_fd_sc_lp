* File: sky130_fd_sc_lp__a41oi_1.pex.spice
* Created: Wed Sep  2 09:29:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41OI_1%B1 1 3 6 8 9 10
c27 6 0 4.46493e-20 $X=0.565 $Y=2.465
c28 1 0 1.50396e-19 $X=0.565 $Y=1.185
r29 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.35 $X2=0.32 $Y2=1.35
r30 8 13 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.49 $Y=1.35 $X2=0.32
+ $Y2=1.35
r31 8 9 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.49 $Y=1.35 $X2=0.565
+ $Y2=1.35
r32 4 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.515
+ $X2=0.565 $Y2=1.35
r33 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.565 $Y=1.515
+ $X2=0.565 $Y2=2.465
r34 1 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.185
+ $X2=0.565 $Y2=1.35
r35 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.565 $Y=1.185
+ $X2=0.565 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_1%A4 3 7 9 10 18
c41 9 0 2.58448e-19 $X=1.2 $Y=1.295
r42 16 18 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=1.14 $Y=1.375
+ $X2=1.445 $Y2=1.375
r43 13 16 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.05 $Y=1.375 $X2=1.14
+ $Y2=1.375
r44 9 10 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.197 $Y=1.295
+ $X2=1.197 $Y2=1.665
r45 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.375 $X2=1.14 $Y2=1.375
r46 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.21
+ $X2=1.445 $Y2=1.375
r47 5 7 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.445 $Y=1.21
+ $X2=1.445 $Y2=0.655
r48 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.54
+ $X2=1.05 $Y2=1.375
r49 1 3 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.05 $Y=1.54 $X2=1.05
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_1%A3 3 7 9 10 14
c37 9 0 3.41837e-20 $X=1.68 $Y=1.295
c38 3 0 6.0165e-20 $X=1.875 $Y=0.655
r39 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.375
+ $X2=1.895 $Y2=1.54
r40 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.375
+ $X2=1.895 $Y2=1.21
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.895
+ $Y=1.375 $X2=1.895 $Y2=1.375
r42 10 15 6.48342 $w=5.33e-07 $l=2.9e-07 $layer=LI1_cond $X=1.792 $Y=1.665
+ $X2=1.792 $Y2=1.375
r43 9 15 1.78853 $w=5.33e-07 $l=8e-08 $layer=LI1_cond $X=1.792 $Y=1.295
+ $X2=1.792 $Y2=1.375
r44 7 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.985 $Y=2.465
+ $X2=1.985 $Y2=1.54
r45 3 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.875 $Y=0.655
+ $X2=1.875 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_1%A2 3 7 8 9 13 15
c34 15 0 3.41837e-20 $X=2.435 $Y=1.185
c35 8 0 6.0165e-20 $X=2.64 $Y=1.295
c36 3 0 1.74124e-19 $X=2.415 $Y=2.465
r37 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.35
+ $X2=2.435 $Y2=1.515
r38 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.35
+ $X2=2.435 $Y2=1.185
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=1.35 $X2=2.435 $Y2=1.35
r40 9 14 7.84926 $w=4.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.51 $Y=1.665
+ $X2=2.51 $Y2=1.35
r41 8 14 1.37051 $w=4.78e-07 $l=5.5e-08 $layer=LI1_cond $X=2.51 $Y=1.295
+ $X2=2.51 $Y2=1.35
r42 7 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.445 $Y=0.655
+ $X2=2.445 $Y2=1.185
r43 3 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.415 $Y=2.465
+ $X2=2.415 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_1%A1 3 6 8 9 13 15
c25 8 0 1.74124e-19 $X=3.12 $Y=1.295
r26 13 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.35
+ $X2=2.99 $Y2=1.515
r27 13 15 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.35
+ $X2=2.99 $Y2=1.185
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.005
+ $Y=1.35 $X2=3.005 $Y2=1.35
r29 9 14 10.2259 $w=3.53e-07 $l=3.15e-07 $layer=LI1_cond $X=3.097 $Y=1.665
+ $X2=3.097 $Y2=1.35
r30 8 14 1.78548 $w=3.53e-07 $l=5.5e-08 $layer=LI1_cond $X=3.097 $Y=1.295
+ $X2=3.097 $Y2=1.35
r31 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.885 $Y=2.465
+ $X2=2.885 $Y2=1.515
r32 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.885 $Y=0.655
+ $X2=2.885 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_1%Y 1 2 3 12 16 20 24 26 27 28 34 39 45
r58 34 39 1.17198 $w=2.93e-07 $l=3e-08 $layer=LI1_cond $X=0.722 $Y=1.695
+ $X2=0.722 $Y2=1.665
r59 33 45 9.16598 $w=1.78e-07 $l=1.48e-07 $layer=LI1_cond $X=0.722 $Y=0.925
+ $X2=0.87 $Y2=0.925
r60 28 34 0.130481 $w=1.68e-07 $l=2e-09 $layer=LI1_cond $X=0.72 $Y=1.78
+ $X2=0.722 $Y2=1.78
r61 28 39 1.09384 $w=2.93e-07 $l=2.8e-08 $layer=LI1_cond $X=0.722 $Y=1.637
+ $X2=0.722 $Y2=1.665
r62 27 28 13.3605 $w=2.93e-07 $l=3.42e-07 $layer=LI1_cond $X=0.722 $Y=1.295
+ $X2=0.722 $Y2=1.637
r63 27 33 10.9384 $w=2.93e-07 $l=2.8e-07 $layer=LI1_cond $X=0.722 $Y=1.295
+ $X2=0.722 $Y2=1.015
r64 26 33 0.123232 $w=1.78e-07 $l=2e-09 $layer=LI1_cond $X=0.72 $Y=0.925
+ $X2=0.722 $Y2=0.925
r65 22 24 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.1 $Y=0.835
+ $X2=3.1 $Y2=0.43
r66 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.935 $Y=0.92
+ $X2=3.1 $Y2=0.835
r67 20 45 134.722 $w=1.68e-07 $l=2.065e-06 $layer=LI1_cond $X=2.935 $Y=0.92
+ $X2=0.87 $Y2=0.92
r68 16 18 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.315 $Y=1.98
+ $X2=0.315 $Y2=2.91
r69 14 28 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.315 $Y=1.78
+ $X2=0.72 $Y2=1.78
r70 14 16 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=0.315 $Y=1.865
+ $X2=0.315 $Y2=1.98
r71 10 26 24.9545 $w=1.78e-07 $l=4.05e-07 $layer=LI1_cond $X=0.315 $Y=0.925
+ $X2=0.72 $Y2=0.925
r72 10 12 17.9515 $w=2.58e-07 $l=4.05e-07 $layer=LI1_cond $X=0.315 $Y=0.835
+ $X2=0.315 $Y2=0.43
r73 3 18 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.835 $X2=0.35 $Y2=2.91
r74 3 16 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.835 $X2=0.35 $Y2=1.98
r75 2 24 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.43
r76 1 12 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=0.225
+ $Y=0.235 $X2=0.35 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_1%A_128_367# 1 2 3 10 12 14 20 22 24 26 30 36
+ 38
r47 35 36 35.8078 $w=1.73e-07 $l=5.65e-07 $layer=LI1_cond $X=2.2 $Y=2.007
+ $X2=1.635 $Y2=2.007
r48 30 32 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.2 $Y=2.01 $X2=1.2
+ $Y2=2.12
r49 24 40 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=2.09
+ $X2=3.125 $Y2=2.005
r50 24 26 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.125 $Y=2.09
+ $X2=3.125 $Y2=2.46
r51 22 40 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.985 $Y=2.005
+ $X2=3.125 $Y2=2.005
r52 22 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.985 $Y=2.005
+ $X2=2.315 $Y2=2.005
r53 18 38 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.21 $Y=2.007
+ $X2=2.315 $Y2=2.007
r54 18 35 0.633766 $w=1.73e-07 $l=1e-08 $layer=LI1_cond $X=2.21 $Y=2.007 $X2=2.2
+ $Y2=2.007
r55 18 20 19.2771 $w=2.08e-07 $l=3.65e-07 $layer=LI1_cond $X=2.21 $Y=2.095
+ $X2=2.21 $Y2=2.46
r56 17 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.01
+ $X2=1.2 $Y2=2.01
r57 17 36 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.285 $Y=2.01
+ $X2=1.635 $Y2=2.01
r58 15 29 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.905 $Y=2.12
+ $X2=0.76 $Y2=2.12
r59 14 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.12
+ $X2=1.2 $Y2=2.12
r60 14 15 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.115 $Y=2.12
+ $X2=0.905 $Y2=2.12
r61 10 29 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=2.205
+ $X2=0.76 $Y2=2.12
r62 10 12 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=0.76 $Y=2.205
+ $X2=0.76 $Y2=2.525
r63 3 40 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.005
r64 3 26 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.46
r65 2 35 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.06
+ $Y=1.835 $X2=2.2 $Y2=2.005
r66 2 20 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=2.06
+ $Y=1.835 $X2=2.2 $Y2=2.46
r67 1 29 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.835 $X2=0.78 $Y2=2.12
r68 1 12 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.64
+ $Y=1.835 $X2=0.78 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_1%VPWR 1 2 7 10 13 17 19 24 31 32 35 38
c50 7 0 6.34028e-20 $X=1.505 $Y=2.805
r51 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.65 $Y2=3.33
r55 29 31 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 25 35 15.1677 $w=1.7e-07 $l=4.3e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=1.505 $Y2=3.33
r59 25 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.485 $Y=3.33
+ $X2=2.65 $Y2=3.33
r61 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 19 35 15.1677 $w=1.7e-07 $l=4.3e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=1.505 $Y2=3.33
r64 19 21 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 17 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 17 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 11 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=3.245
+ $X2=2.65 $Y2=3.33
r69 11 13 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=2.65 $Y=3.245
+ $X2=2.65 $Y2=2.375
r70 8 35 3.26792 $w=8.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=3.245
+ $X2=1.505 $Y2=3.33
r71 8 10 4.18488 $w=8.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.505 $Y=3.245
+ $X2=1.505 $Y2=2.95
r72 7 16 6.22459 $w=8.6e-07 $l=4.3e-07 $layer=LI1_cond $X=1.505 $Y=2.805
+ $X2=1.505 $Y2=2.375
r73 7 10 2.05698 $w=8.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.505 $Y=2.805
+ $X2=1.505 $Y2=2.95
r74 2 13 300 $w=1.7e-07 $l=6.14817e-07 $layer=licon1_PDIFF $count=2 $X=2.49
+ $Y=1.835 $X2=2.65 $Y2=2.375
r75 1 16 300 $w=1.7e-07 $l=8.74257e-07 $layer=licon1_PDIFF $count=2 $X=1.125
+ $Y=1.835 $X2=1.77 $Y2=2.375
r76 1 10 300 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=2 $X=1.125
+ $Y=1.835 $X2=1.265 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_1%VGND 1 4 16 17 22 28
r32 27 28 11.123 $w=7.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=0.29
+ $X2=1.395 $Y2=0.29
r33 24 27 0.478431 $w=7.48e-07 $l=3e-08 $layer=LI1_cond $X=1.2 $Y=0.29 $X2=1.23
+ $Y2=0.29
r34 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r36 20 24 7.6549 $w=7.48e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=0.29 $X2=1.2
+ $Y2=0.29
r37 20 22 10.1661 $w=7.48e-07 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=0.29
+ $X2=0.615 $Y2=0.29
r38 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 13 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r41 13 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.395
+ $Y2=0
r42 9 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r43 8 22 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.615
+ $Y2=0
r44 8 9 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r45 4 17 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r46 4 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r47 4 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r48 1 27 91 $w=1.7e-07 $l=7.2667e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.235 $X2=1.23 $Y2=0.54
.ends

