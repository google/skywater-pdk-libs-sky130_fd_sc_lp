# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a311o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a311o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.315000 1.210000 7.595000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.775000 1.345000 6.375000 1.750000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.895000 1.415000 5.605000 1.750000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.970000 1.415000 1.865000 1.750000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.430000 1.750000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.430400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 0.255000 2.560000 1.025000 ;
        RECT 2.375000 1.025000 4.230000 1.195000 ;
        RECT 2.990000 1.750000 4.395000 2.015000 ;
        RECT 3.230000 0.255000 3.420000 1.025000 ;
        RECT 4.060000 1.195000 4.230000 1.405000 ;
        RECT 4.060000 1.405000 4.725000 1.750000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.100000  0.085000 0.430000 1.040000 ;
      RECT 0.100000  1.920000 0.430000 2.905000 ;
      RECT 0.100000  2.905000 2.120000 3.075000 ;
      RECT 0.600000  0.255000 0.805000 1.075000 ;
      RECT 0.600000  1.075000 2.205000 1.245000 ;
      RECT 0.600000  1.245000 0.790000 2.735000 ;
      RECT 0.960000  1.920000 1.290000 2.905000 ;
      RECT 0.975000  0.085000 1.305000 0.905000 ;
      RECT 1.460000  1.920000 2.460000 2.090000 ;
      RECT 1.460000  2.090000 1.690000 2.735000 ;
      RECT 1.475000  0.255000 1.690000 1.075000 ;
      RECT 1.860000  0.085000 2.190000 0.905000 ;
      RECT 1.860000  2.260000 2.120000 2.905000 ;
      RECT 2.035000  1.245000 2.205000 1.365000 ;
      RECT 2.035000  1.365000 3.865000 1.535000 ;
      RECT 2.035000  1.535000 2.810000 1.585000 ;
      RECT 2.290000  2.090000 2.460000 2.525000 ;
      RECT 2.290000  2.525000 5.280000 2.695000 ;
      RECT 2.465000  2.865000 2.795000 3.245000 ;
      RECT 2.640000  1.585000 2.810000 2.185000 ;
      RECT 2.640000  2.185000 4.735000 2.355000 ;
      RECT 2.730000  0.085000 3.060000 0.855000 ;
      RECT 3.480000  2.865000 3.810000 3.245000 ;
      RECT 3.590000  0.085000 4.260000 0.855000 ;
      RECT 4.430000  0.255000 4.620000 1.065000 ;
      RECT 4.430000  1.065000 6.245000 1.175000 ;
      RECT 4.430000  1.175000 5.380000 1.235000 ;
      RECT 4.565000  1.920000 6.715000 2.090000 ;
      RECT 4.565000  2.090000 4.735000 2.185000 ;
      RECT 4.590000  2.865000 4.920000 3.245000 ;
      RECT 4.790000  0.085000 5.120000 0.845000 ;
      RECT 5.020000  2.260000 7.075000 2.430000 ;
      RECT 5.020000  2.430000 5.280000 2.525000 ;
      RECT 5.090000  2.695000 5.280000 3.075000 ;
      RECT 5.210000  1.005000 6.245000 1.065000 ;
      RECT 5.450000  0.255000 7.575000 0.425000 ;
      RECT 5.450000  0.425000 5.745000 0.835000 ;
      RECT 5.450000  2.600000 5.780000 3.245000 ;
      RECT 5.915000  0.595000 6.245000 1.005000 ;
      RECT 5.950000  2.430000 6.160000 3.075000 ;
      RECT 6.345000  2.600000 6.675000 3.245000 ;
      RECT 6.415000  0.425000 6.645000 1.175000 ;
      RECT 6.545000  1.345000 7.145000 1.645000 ;
      RECT 6.545000  1.645000 6.715000 1.920000 ;
      RECT 6.815000  0.595000 7.145000 1.345000 ;
      RECT 6.845000  2.430000 7.075000 3.075000 ;
      RECT 6.885000  1.815000 7.075000 2.260000 ;
      RECT 7.245000  1.920000 7.575000 3.245000 ;
      RECT 7.315000  0.425000 7.575000 1.040000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__a311o_4
END LIBRARY
