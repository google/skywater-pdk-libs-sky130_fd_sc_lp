* File: sky130_fd_sc_lp__or4bb_2.pex.spice
* Created: Wed Sep  2 10:33:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4BB_2%C_N 3 5 7 8 9 12 14 15 16 17 22 24
r46 22 24 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.652 $Y=0.93
+ $X2=0.652 $Y2=0.765
r47 16 17 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.697 $Y=0.925
+ $X2=0.697 $Y2=1.295
r48 16 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.675
+ $Y=0.93 $X2=0.675 $Y2=0.93
r49 15 16 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.697 $Y=0.555
+ $X2=0.697 $Y2=0.925
r50 10 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=0.875 $Y=1.835
+ $X2=0.875 $Y2=2.225
r51 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.8 $Y=1.76
+ $X2=0.875 $Y2=1.835
r52 8 9 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.8 $Y=1.76 $X2=0.615
+ $Y2=1.76
r53 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.54 $Y=1.685
+ $X2=0.615 $Y2=1.76
r54 7 14 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.54 $Y=1.685
+ $X2=0.54 $Y2=1.435
r55 5 14 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.652 $Y=1.248
+ $X2=0.652 $Y2=1.435
r56 4 22 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.652 $Y=0.952
+ $X2=0.652 $Y2=0.93
r57 4 5 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.652 $Y=0.952
+ $X2=0.652 $Y2=1.248
r58 3 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=0.445
+ $X2=0.54 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_2%A 3 6 9 10 11 12 13 17
c39 6 0 1.83188e-19 $X=1.305 $Y=2.225
r40 12 13 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.172 $Y=0.925
+ $X2=1.172 $Y2=1.295
r41 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.215
+ $Y=0.94 $X2=1.215 $Y2=0.94
r42 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.215 $Y=1.28
+ $X2=1.215 $Y2=0.94
r43 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=1.28
+ $X2=1.215 $Y2=1.445
r44 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=0.775
+ $X2=1.215 $Y2=0.94
r45 6 11 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.305 $Y=2.225
+ $X2=1.305 $Y2=1.445
r46 3 9 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.305 $Y=0.445
+ $X2=1.305 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_2%B 3 7 9 12 13
r37 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.02
+ $X2=1.755 $Y2=1.185
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.02
+ $X2=1.755 $Y2=0.855
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.755
+ $Y=1.02 $X2=1.755 $Y2=1.02
r40 9 13 7.54576 $w=4.18e-07 $l=2.75e-07 $layer=LI1_cond $X=1.71 $Y=1.295
+ $X2=1.71 $Y2=1.02
r41 7 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.735 $Y=0.445
+ $X2=1.735 $Y2=0.855
r42 3 15 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.665 $Y=2.225
+ $X2=1.665 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_2%A_40_47# 1 2 9 13 18 24 28 30 31 34 35
c74 28 0 1.83188e-19 $X=0.66 $Y=2.225
c75 18 0 1.79926e-19 $X=2.295 $Y=1.395
r76 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.295
+ $Y=1.04 $X2=2.295 $Y2=1.04
r77 32 34 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=2.295 $Y=1.625
+ $X2=2.295 $Y2=1.04
r78 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.13 $Y=1.71
+ $X2=2.295 $Y2=1.625
r79 30 31 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=2.13 $Y=1.71
+ $X2=0.79 $Y2=1.71
r80 26 31 9.65561 $w=1.68e-07 $l=1.48e-07 $layer=LI1_cond $X=0.642 $Y=1.71
+ $X2=0.79 $Y2=1.71
r81 26 28 16.7983 $w=2.93e-07 $l=4.3e-07 $layer=LI1_cond $X=0.642 $Y=1.795
+ $X2=0.642 $Y2=2.225
r82 22 26 23.2909 $w=1.68e-07 $l=3.57e-07 $layer=LI1_cond $X=0.285 $Y=1.71
+ $X2=0.642 $Y2=1.71
r83 22 24 54.3953 $w=2.48e-07 $l=1.18e-06 $layer=LI1_cond $X=0.285 $Y=1.625
+ $X2=0.285 $Y2=0.445
r84 21 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=0.875
+ $X2=2.295 $Y2=1.04
r85 18 35 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.295 $Y=1.395
+ $X2=2.295 $Y2=1.04
r86 15 18 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.025 $Y=1.47
+ $X2=2.295 $Y2=1.47
r87 13 21 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.385 $Y=0.445
+ $X2=2.385 $Y2=0.875
r88 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.025 $Y=1.545
+ $X2=2.025 $Y2=1.47
r89 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.025 $Y=1.545
+ $X2=2.025 $Y2=2.225
r90 2 28 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.535
+ $Y=2.015 $X2=0.66 $Y2=2.225
r91 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.235 $X2=0.325 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_2%A_462_351# 1 2 7 9 10 11 13 16 19 21 23 27
+ 30 31 33 35 36 37 40 44 46 49
c109 35 0 1.71309e-19 $X=4.035 $Y=2.445
c110 16 0 6.95413e-20 $X=2.815 $Y=0.445
c111 13 0 5.454e-20 $X=2.745 $Y=1.755
r112 42 44 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=4.5 $Y=1.065 $X2=4.5
+ $Y2=0.865
r113 38 46 0.432806 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=4.205 $Y=2.095
+ $X2=4.035 $Y2=2.095
r114 38 40 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.205 $Y=2.095
+ $X2=4.535 $Y2=2.095
r115 36 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.335 $Y=1.15
+ $X2=4.5 $Y2=1.065
r116 36 37 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.335 $Y=1.15
+ $X2=4.035 $Y2=1.15
r117 34 46 6.36606 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=2.26
+ $X2=4.035 $Y2=2.095
r118 34 35 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=4.035 $Y=2.26
+ $X2=4.035 $Y2=2.445
r119 33 46 6.36606 $w=2.55e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.95 $Y=1.93
+ $X2=4.035 $Y2=2.095
r120 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.95 $Y=1.235
+ $X2=4.035 $Y2=1.15
r121 32 33 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.95 $Y=1.235
+ $X2=3.95 $Y2=1.93
r122 30 35 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.865 $Y=2.53
+ $X2=4.035 $Y2=2.445
r123 30 31 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.865 $Y=2.53
+ $X2=2.805 $Y2=2.53
r124 28 49 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=2.64 $Y=2.94
+ $X2=2.875 $Y2=2.94
r125 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.64
+ $Y=2.94 $X2=2.64 $Y2=2.94
r126 25 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.64 $Y=2.615
+ $X2=2.805 $Y2=2.53
r127 25 27 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.64 $Y=2.615
+ $X2=2.64 $Y2=2.94
r128 22 23 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=2.745 $Y=1.83
+ $X2=2.875 $Y2=1.83
r129 20 21 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.78 $Y=0.795
+ $X2=2.78 $Y2=0.945
r130 19 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=2.775
+ $X2=2.875 $Y2=2.94
r131 18 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=1.905
+ $X2=2.875 $Y2=1.83
r132 18 19 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=2.875 $Y=1.905
+ $X2=2.875 $Y2=2.775
r133 16 20 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.815 $Y=0.445
+ $X2=2.815 $Y2=0.795
r134 13 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.745 $Y=1.755
+ $X2=2.745 $Y2=1.83
r135 13 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.745 $Y=1.755
+ $X2=2.745 $Y2=0.945
r136 10 22 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.67 $Y=1.83
+ $X2=2.745 $Y2=1.83
r137 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.67 $Y=1.83
+ $X2=2.46 $Y2=1.83
r138 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.385 $Y=1.905
+ $X2=2.46 $Y2=1.83
r139 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.385 $Y=1.905
+ $X2=2.385 $Y2=2.225
r140 2 40 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.835 $X2=4.535 $Y2=2.055
r141 1 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.36
+ $Y=0.655 $X2=4.5 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_2%A_276_47# 1 2 3 10 12 13 15 16 18 20 23 25
+ 28 30 31 33 35 38 42 49 51
c119 49 0 1.41502e-20 $X=2.725 $Y=2.135
c120 35 0 1.65776e-19 $X=2.725 $Y=1.995
c121 30 0 6.95413e-20 $X=2.435 $Y=0.67
r122 47 49 5.14483 $w=2.78e-07 $l=1.25e-07 $layer=LI1_cond $X=2.6 $Y=2.135
+ $X2=2.725 $Y2=2.135
r123 39 52 14.6061 $w=2.97e-07 $l=9e-08 $layer=POLY_cond $X=3.235 $Y=1.35
+ $X2=3.235 $Y2=1.26
r124 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.195
+ $Y=1.35 $X2=3.195 $Y2=1.35
r125 36 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=1.35
+ $X2=2.725 $Y2=1.35
r126 36 38 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.81 $Y=1.35
+ $X2=3.195 $Y2=1.35
r127 35 49 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.725 $Y=1.995
+ $X2=2.725 $Y2=2.135
r128 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=1.515
+ $X2=2.725 $Y2=1.35
r129 34 35 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.725 $Y=1.515
+ $X2=2.725 $Y2=1.995
r130 33 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=1.185
+ $X2=2.725 $Y2=1.35
r131 33 45 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.725 $Y=1.185
+ $X2=2.725 $Y2=0.755
r132 30 45 6.09592 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=2.622 $Y=0.67
+ $X2=2.622 $Y2=0.755
r133 30 42 6.91466 $w=3.73e-07 $l=2.25e-07 $layer=LI1_cond $X=2.622 $Y=0.67
+ $X2=2.622 $Y2=0.445
r134 30 31 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.435 $Y=0.67
+ $X2=1.65 $Y2=0.67
r135 26 31 13.1706 $w=1.08e-07 $l=1.54771e-07 $layer=LI1_cond $X=1.532 $Y=0.585
+ $X2=1.65 $Y2=0.67
r136 26 28 7.60122 $w=2.33e-07 $l=1.55e-07 $layer=LI1_cond $X=1.532 $Y=0.585
+ $X2=1.532 $Y2=0.43
r137 21 25 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=3.795 $Y=1.335
+ $X2=3.777 $Y2=1.26
r138 21 23 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.795 $Y=1.335
+ $X2=3.795 $Y2=2.465
r139 18 25 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=3.76 $Y=1.185
+ $X2=3.777 $Y2=1.26
r140 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.76 $Y=1.185
+ $X2=3.76 $Y2=0.655
r141 17 52 18.7323 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.405 $Y=1.26
+ $X2=3.235 $Y2=1.26
r142 16 25 5.30422 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=3.685 $Y=1.26
+ $X2=3.777 $Y2=1.26
r143 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.685 $Y=1.26
+ $X2=3.405 $Y2=1.26
r144 13 39 72.647 $w=2.97e-07 $l=4.35172e-07 $layer=POLY_cond $X=3.365 $Y=1.725
+ $X2=3.235 $Y2=1.35
r145 13 15 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.365 $Y=1.725
+ $X2=3.365 $Y2=2.465
r146 10 52 23.9601 $w=2.97e-07 $l=1.27083e-07 $layer=POLY_cond $X=3.33 $Y=1.185
+ $X2=3.235 $Y2=1.26
r147 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.33 $Y=1.185
+ $X2=3.33 $Y2=0.655
r148 3 47 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=2.015 $X2=2.6 $Y2=2.16
r149 2 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.235 $X2=2.6 $Y2=0.445
r150 1 28 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.38
+ $Y=0.235 $X2=1.52 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_2%D_N 3 7 9 12
r26 12 15 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.377 $Y=1.51
+ $X2=4.377 $Y2=1.675
r27 12 14 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.377 $Y=1.51
+ $X2=4.377 $Y2=1.345
r28 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.38
+ $Y=1.51 $X2=4.38 $Y2=1.51
r29 9 13 5.84337 $w=3.53e-07 $l=1.8e-07 $layer=LI1_cond $X=4.56 $Y=1.582
+ $X2=4.38 $Y2=1.582
r30 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.32 $Y=2.045
+ $X2=4.32 $Y2=1.675
r31 3 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.285 $Y=0.865
+ $X2=4.285 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_2%VPWR 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
c51 3 0 1.71309e-19 $X=3.87 $Y=1.835
r52 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.175 $Y=3.33
+ $X2=4.01 $Y2=3.33
r58 39 41 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.175 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.15 $Y2=3.33
r63 35 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.6 $Y2=3.33
r64 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=4.01 $Y2=3.33
r65 34 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=3.6 $Y2=3.33
r66 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 30 45 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=1.107 $Y2=3.33
r69 30 32 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=2.64 $Y2=3.33
r70 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=3.33
+ $X2=3.15 $Y2=3.33
r71 29 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=3.33
+ $X2=2.64 $Y2=3.33
r72 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 24 45 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=1.107 $Y2=3.33
r75 24 26 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r77 22 46 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r78 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.01 $Y=3.245
+ $X2=4.01 $Y2=3.33
r79 18 20 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.01 $Y=3.245
+ $X2=4.01 $Y2=2.89
r80 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=3.245
+ $X2=3.15 $Y2=3.33
r81 14 16 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.15 $Y=3.245
+ $X2=3.15 $Y2=2.89
r82 10 45 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.107 $Y=3.245
+ $X2=1.107 $Y2=3.33
r83 10 12 39.8472 $w=2.93e-07 $l=1.02e-06 $layer=LI1_cond $X=1.107 $Y=3.245
+ $X2=1.107 $Y2=2.225
r84 3 20 600 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.835 $X2=4.01 $Y2=2.89
r85 2 16 600 $w=1.7e-07 $l=1.11575e-06 $layer=licon1_PDIFF $count=1 $X=3.025
+ $Y=1.835 $X2=3.15 $Y2=2.89
r86 1 12 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.95
+ $Y=2.015 $X2=1.09 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_2%X 1 2 7 8 9 10 11 18
c21 18 0 5.454e-20 $X=3.545 $Y=0.42
r22 10 11 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.572 $Y=1.665
+ $X2=3.572 $Y2=2.035
r23 9 10 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.572 $Y=1.295
+ $X2=3.572 $Y2=1.665
r24 8 9 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.572 $Y=0.925
+ $X2=3.572 $Y2=1.295
r25 7 8 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.572 $Y=0.555
+ $X2=3.572 $Y2=0.925
r26 7 18 6.3502 $w=2.43e-07 $l=1.35e-07 $layer=LI1_cond $X=3.572 $Y=0.555
+ $X2=3.572 $Y2=0.42
r27 2 11 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.835 $X2=3.58 $Y2=2.11
r28 1 18 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.235 $X2=3.545 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_2%VGND 1 2 3 4 15 19 25 28 29 30 31 38 39 40
+ 49 58 59 62
r78 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r79 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r80 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r81 56 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r82 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r83 53 62 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.28 $Y=0 $X2=3.13
+ $Y2=0
r84 53 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.28 $Y=0 $X2=3.6
+ $Y2=0
r85 52 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r86 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r87 49 62 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.98 $Y=0 $X2=3.13
+ $Y2=0
r88 49 51 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.98 $Y=0 $X2=2.64
+ $Y2=0
r89 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r90 44 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r91 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r92 40 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r93 40 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r94 38 55 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.865 $Y=0 $X2=3.6
+ $Y2=0
r95 38 39 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=3.865 $Y=0 $X2=4.002
+ $Y2=0
r96 37 58 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.56
+ $Y2=0
r97 37 39 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.002
+ $Y2=0
r98 33 51 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.64
+ $Y2=0
r99 31 47 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.68
+ $Y2=0
r100 30 35 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.03
+ $Y2=0.32
r101 30 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.195
+ $Y2=0
r102 30 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=1.865
+ $Y2=0
r103 28 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0
+ $X2=0.72 $Y2=0
r104 28 29 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.115
+ $Y2=0
r105 27 47 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.245 $Y=0
+ $X2=1.68 $Y2=0
r106 27 29 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.115
+ $Y2=0
r107 23 39 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.002 $Y=0.085
+ $X2=4.002 $Y2=0
r108 23 25 12.3626 $w=2.73e-07 $l=2.95e-07 $layer=LI1_cond $X=4.002 $Y=0.085
+ $X2=4.002 $Y2=0.38
r109 19 21 18.0549 $w=2.98e-07 $l=4.7e-07 $layer=LI1_cond $X=3.13 $Y=0.38
+ $X2=3.13 $Y2=0.85
r110 17 62 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0
r111 17 19 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0.38
r112 13 29 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0
r113 13 15 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.44
r114 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.835
+ $Y=0.235 $X2=3.975 $Y2=0.38
r115 3 21 182 $w=1.7e-07 $l=7.18749e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.235 $X2=3.115 $Y2=0.85
r116 3 19 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.235 $X2=3.115 $Y2=0.38
r117 2 35 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=1.81
+ $Y=0.235 $X2=2.03 $Y2=0.32
r118 1 15 182 $w=1.7e-07 $l=5.68331e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=1.09 $Y2=0.44
.ends

