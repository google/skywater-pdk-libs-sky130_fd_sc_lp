* File: sky130_fd_sc_lp__o311a_2.pxi.spice
* Created: Fri Aug 28 11:13:39 2020
* 
x_PM_SKY130_FD_SC_LP__O311A_2%A_85_21# N_A_85_21#_M1007_d N_A_85_21#_M1005_d
+ N_A_85_21#_M1001_d N_A_85_21#_c_72_n N_A_85_21#_M1012_g N_A_85_21#_M1003_g
+ N_A_85_21#_c_74_n N_A_85_21#_M1013_g N_A_85_21#_M1011_g N_A_85_21#_c_76_n
+ N_A_85_21#_c_77_n N_A_85_21#_c_78_n N_A_85_21#_c_161_p N_A_85_21#_c_104_p
+ N_A_85_21#_c_105_p N_A_85_21#_c_109_p N_A_85_21#_c_79_n N_A_85_21#_c_80_n
+ N_A_85_21#_c_85_n N_A_85_21#_c_81_n N_A_85_21#_c_86_n
+ PM_SKY130_FD_SC_LP__O311A_2%A_85_21#
x_PM_SKY130_FD_SC_LP__O311A_2%A1 N_A1_M1009_g N_A1_M1000_g A1 A1 A1 A1
+ N_A1_c_187_n N_A1_c_188_n PM_SKY130_FD_SC_LP__O311A_2%A1
x_PM_SKY130_FD_SC_LP__O311A_2%A2 N_A2_c_225_n N_A2_M1008_g N_A2_M1004_g A2 A2 A2
+ A2 N_A2_c_229_n PM_SKY130_FD_SC_LP__O311A_2%A2
x_PM_SKY130_FD_SC_LP__O311A_2%A3 N_A3_M1005_g N_A3_M1002_g A3 A3 A3 A3
+ N_A3_c_261_n N_A3_c_262_n A3 PM_SKY130_FD_SC_LP__O311A_2%A3
x_PM_SKY130_FD_SC_LP__O311A_2%B1 N_B1_M1006_g N_B1_M1010_g B1 N_B1_c_299_n
+ N_B1_c_300_n PM_SKY130_FD_SC_LP__O311A_2%B1
x_PM_SKY130_FD_SC_LP__O311A_2%C1 N_C1_M1007_g N_C1_M1001_g N_C1_c_336_n C1
+ N_C1_c_337_n N_C1_c_338_n PM_SKY130_FD_SC_LP__O311A_2%C1
x_PM_SKY130_FD_SC_LP__O311A_2%VPWR N_VPWR_M1003_d N_VPWR_M1011_d N_VPWR_M1006_d
+ N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n
+ N_VPWR_c_367_n N_VPWR_c_368_n VPWR N_VPWR_c_369_n N_VPWR_c_361_n
+ N_VPWR_c_371_n PM_SKY130_FD_SC_LP__O311A_2%VPWR
x_PM_SKY130_FD_SC_LP__O311A_2%X N_X_M1012_s N_X_M1003_s X X X X X X X
+ N_X_c_418_n X PM_SKY130_FD_SC_LP__O311A_2%X
x_PM_SKY130_FD_SC_LP__O311A_2%VGND N_VGND_M1012_d N_VGND_M1013_d N_VGND_M1004_d
+ N_VGND_c_445_n N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n VGND
+ N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n
+ N_VGND_c_454_n PM_SKY130_FD_SC_LP__O311A_2%VGND
x_PM_SKY130_FD_SC_LP__O311A_2%A_355_47# N_A_355_47#_M1009_d N_A_355_47#_M1002_d
+ N_A_355_47#_c_503_n N_A_355_47#_c_510_n N_A_355_47#_c_504_n
+ N_A_355_47#_c_505_n N_A_355_47#_c_517_n PM_SKY130_FD_SC_LP__O311A_2%A_355_47#
cc_1 VNB N_A_85_21#_c_72_n 0.021472f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_2 VNB N_A_85_21#_M1003_g 0.0106048f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.465
cc_3 VNB N_A_85_21#_c_74_n 0.0176818f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.185
cc_4 VNB N_A_85_21#_M1011_g 0.00784811f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.465
cc_5 VNB N_A_85_21#_c_76_n 0.00563066f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.35
cc_6 VNB N_A_85_21#_c_77_n 0.0730855f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.35
cc_7 VNB N_A_85_21#_c_78_n 0.0319241f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=1.09
cc_8 VNB N_A_85_21#_c_79_n 0.00338599f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.92
cc_9 VNB N_A_85_21#_c_80_n 0.0310117f $X=-0.19 $Y=-0.245 $X2=3.895 $Y2=0.42
cc_10 VNB N_A_85_21#_c_81_n 0.00928985f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=1.005
cc_11 VNB N_A1_M1009_g 0.0280369f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=1.835
cc_12 VNB N_A1_c_187_n 0.0225493f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.655
cc_13 VNB N_A1_c_188_n 0.00508996f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=2.01
cc_14 VNB N_A2_c_225_n 0.0275833f $X=-0.19 $Y=-0.245 $X2=3.755 $Y2=0.235
cc_15 VNB N_A2_M1004_g 0.0257473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A3_M1002_g 0.0273335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_c_261_n 0.0242707f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.655
cc_18 VNB N_A3_c_262_n 0.00402047f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.515
cc_19 VNB N_B1_M1010_g 0.0245109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_299_n 0.0243232f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_21 VNB N_B1_c_300_n 0.00430745f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.515
cc_22 VNB N_C1_M1007_g 0.0272802f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=1.835
cc_23 VNB N_C1_M1001_g 0.00138656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C1_c_336_n 0.00900014f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_25 VNB N_C1_c_337_n 0.0495368f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.465
cc_26 VNB N_C1_c_338_n 0.0146189f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.465
cc_27 VNB N_VPWR_c_361_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_418_n 0.00289552f $X=-0.19 $Y=-0.245 $X2=1.107 $Y2=1.175
cc_29 VNB N_VGND_c_445_n 0.0118954f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_30 VNB N_VGND_c_446_n 0.0502045f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_31 VNB N_VGND_c_447_n 0.00183778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_448_n 0.00561608f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.515
cc_33 VNB N_VGND_c_449_n 0.0145469f $X=-0.19 $Y=-0.245 $X2=1.107 $Y2=1.175
cc_34 VNB N_VGND_c_450_n 0.0170954f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=1.09
cc_35 VNB N_VGND_c_451_n 0.0452864f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=2.01
cc_36 VNB N_VGND_c_452_n 0.235754f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.175
cc_37 VNB N_VGND_c_453_n 0.010461f $X=-0.19 $Y=-0.245 $X2=3.935 $Y2=2.1
cc_38 VNB N_VGND_c_454_n 0.00631622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A_85_21#_M1003_g 0.0264965f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.465
cc_40 VPB N_A_85_21#_M1011_g 0.0223078f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.465
cc_41 VPB N_A_85_21#_c_79_n 0.00138441f $X=-0.19 $Y=1.655 $X2=3.58 $Y2=1.92
cc_42 VPB N_A_85_21#_c_85_n 0.0369431f $X=-0.19 $Y=1.655 $X2=3.9 $Y2=2.91
cc_43 VPB N_A_85_21#_c_86_n 0.00743827f $X=-0.19 $Y=1.655 $X2=3.9 $Y2=2.095
cc_44 VPB N_A1_M1000_g 0.0191378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB A1 0.00319098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A1_c_187_n 0.00640403f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.655
cc_47 VPB N_A1_c_188_n 0.00639023f $X=-0.19 $Y=1.655 $X2=3.135 $Y2=2.01
cc_48 VPB N_A2_c_225_n 0.00677426f $X=-0.19 $Y=1.655 $X2=3.755 $Y2=0.235
cc_49 VPB N_A2_M1008_g 0.018701f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=1.835
cc_50 VPB N_A2_c_229_n 9.94852e-19 $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.655
cc_51 VPB N_A3_M1005_g 0.0206316f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=1.835
cc_52 VPB A3 0.00184642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A3_c_261_n 0.0076032f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.655
cc_54 VPB N_A3_c_262_n 0.004117f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.515
cc_55 VPB N_B1_M1006_g 0.0207498f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=1.835
cc_56 VPB N_B1_c_299_n 0.00631139f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.655
cc_57 VPB N_B1_c_300_n 0.00247208f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.515
cc_58 VPB N_C1_M1001_g 0.0240952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_C1_c_338_n 0.0131508f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.465
cc_60 VPB N_VPWR_c_362_n 0.0123094f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.185
cc_61 VPB N_VPWR_c_363_n 0.064594f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.655
cc_62 VPB N_VPWR_c_364_n 0.0199524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_365_n 0.00530675f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.515
cc_64 VPB N_VPWR_c_366_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.35
cc_65 VPB N_VPWR_c_367_n 0.0505741f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=1.09
cc_66 VPB N_VPWR_c_368_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.235 $Y2=1.09
cc_67 VPB N_VPWR_c_369_n 0.0204674f $X=-0.19 $Y=1.655 $X2=3.895 $Y2=0.42
cc_68 VPB N_VPWR_c_361_n 0.0535861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_371_n 0.00516749f $X=-0.19 $Y=1.655 $X2=3 $Y2=2.085
cc_70 VPB X 0.0032582f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.185
cc_71 VPB N_X_c_418_n 3.67206e-19 $X=-0.19 $Y=1.655 $X2=1.107 $Y2=1.175
cc_72 N_A_85_21#_c_74_n N_A1_M1009_g 0.00539789f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_73 N_A_85_21#_c_76_n N_A1_M1009_g 0.00110519f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_74 N_A_85_21#_c_77_n N_A1_M1009_g 0.00583392f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_75 N_A_85_21#_c_78_n N_A1_M1009_g 0.0161259f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_76 N_A_85_21#_M1011_g N_A1_M1000_g 0.0210158f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A_85_21#_M1011_g A1 0.00240959f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_85_21#_M1011_g N_A1_c_187_n 0.0041151f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A_85_21#_c_76_n N_A1_c_187_n 2.1416e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_80 N_A_85_21#_c_77_n N_A1_c_187_n 0.0113541f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_81 N_A_85_21#_c_78_n N_A1_c_187_n 0.0040357f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_82 N_A_85_21#_M1011_g N_A1_c_188_n 7.10266e-19 $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A_85_21#_c_76_n N_A1_c_188_n 0.0106754f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_84 N_A_85_21#_c_77_n N_A1_c_188_n 6.82967e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_85 N_A_85_21#_c_78_n N_A1_c_188_n 0.0286679f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_86 N_A_85_21#_c_78_n N_A2_c_225_n 0.00509038f $X=3.485 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A_85_21#_c_78_n N_A2_M1004_g 0.011695f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_88 N_A_85_21#_c_78_n N_A2_c_229_n 0.0236755f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_89 N_A_85_21#_c_104_p N_A3_M1005_g 7.3896e-19 $X=3.015 $Y=2.1 $X2=0 $Y2=0
cc_90 N_A_85_21#_c_105_p N_A3_M1005_g 0.00562714f $X=3 $Y=2.91 $X2=0 $Y2=0
cc_91 N_A_85_21#_c_78_n N_A3_M1002_g 0.0128423f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_92 N_A_85_21#_c_78_n N_A3_c_261_n 0.00125478f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_93 N_A_85_21#_c_78_n N_A3_c_262_n 0.0261586f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_94 N_A_85_21#_c_109_p N_B1_M1006_g 0.0129999f $X=3.485 $Y=2.01 $X2=0 $Y2=0
cc_95 N_A_85_21#_c_79_n N_B1_M1006_g 0.00406893f $X=3.58 $Y=1.92 $X2=0 $Y2=0
cc_96 N_A_85_21#_c_78_n N_B1_M1010_g 0.0174034f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_97 N_A_85_21#_c_79_n N_B1_M1010_g 0.00587749f $X=3.58 $Y=1.92 $X2=0 $Y2=0
cc_98 N_A_85_21#_c_80_n N_B1_M1010_g 0.00919479f $X=3.895 $Y=0.42 $X2=0 $Y2=0
cc_99 N_A_85_21#_c_78_n N_B1_c_299_n 0.00126279f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_100 N_A_85_21#_c_104_p N_B1_c_299_n 4.24685e-19 $X=3.015 $Y=2.1 $X2=0 $Y2=0
cc_101 N_A_85_21#_c_109_p N_B1_c_299_n 0.00157899f $X=3.485 $Y=2.01 $X2=0 $Y2=0
cc_102 N_A_85_21#_c_78_n N_B1_c_300_n 0.0256465f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_103 N_A_85_21#_c_104_p N_B1_c_300_n 0.0130754f $X=3.015 $Y=2.1 $X2=0 $Y2=0
cc_104 N_A_85_21#_c_109_p N_B1_c_300_n 0.0117274f $X=3.485 $Y=2.01 $X2=0 $Y2=0
cc_105 N_A_85_21#_c_79_n N_B1_c_300_n 0.0306931f $X=3.58 $Y=1.92 $X2=0 $Y2=0
cc_106 N_A_85_21#_c_79_n N_C1_M1007_g 0.00582779f $X=3.58 $Y=1.92 $X2=0 $Y2=0
cc_107 N_A_85_21#_c_80_n N_C1_M1007_g 0.017127f $X=3.895 $Y=0.42 $X2=0 $Y2=0
cc_108 N_A_85_21#_c_81_n N_C1_M1007_g 0.0102351f $X=3.485 $Y=1.005 $X2=0 $Y2=0
cc_109 N_A_85_21#_c_79_n N_C1_M1001_g 0.0107163f $X=3.58 $Y=1.92 $X2=0 $Y2=0
cc_110 N_A_85_21#_c_86_n N_C1_M1001_g 0.0146759f $X=3.9 $Y=2.095 $X2=0 $Y2=0
cc_111 N_A_85_21#_c_79_n N_C1_c_336_n 0.00951201f $X=3.58 $Y=1.92 $X2=0 $Y2=0
cc_112 N_A_85_21#_c_81_n N_C1_c_336_n 0.00945109f $X=3.485 $Y=1.005 $X2=0 $Y2=0
cc_113 N_A_85_21#_c_86_n N_C1_c_337_n 0.003345f $X=3.9 $Y=2.095 $X2=0 $Y2=0
cc_114 N_A_85_21#_c_79_n N_C1_c_338_n 0.0315415f $X=3.58 $Y=1.92 $X2=0 $Y2=0
cc_115 N_A_85_21#_c_81_n N_C1_c_338_n 0.0184528f $X=3.485 $Y=1.005 $X2=0 $Y2=0
cc_116 N_A_85_21#_c_86_n N_C1_c_338_n 0.019503f $X=3.9 $Y=2.095 $X2=0 $Y2=0
cc_117 N_A_85_21#_c_109_p N_VPWR_M1006_d 0.00455122f $X=3.485 $Y=2.01 $X2=0
+ $Y2=0
cc_118 N_A_85_21#_c_79_n N_VPWR_M1006_d 9.78012e-19 $X=3.58 $Y=1.92 $X2=0 $Y2=0
cc_119 N_A_85_21#_c_86_n N_VPWR_M1006_d 7.41438e-19 $X=3.9 $Y=2.095 $X2=0 $Y2=0
cc_120 N_A_85_21#_M1003_g N_VPWR_c_363_n 0.00885808f $X=0.535 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_A_85_21#_M1003_g N_VPWR_c_364_n 0.00564131f $X=0.535 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_A_85_21#_M1011_g N_VPWR_c_364_n 0.0054895f $X=0.965 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_85_21#_M1011_g N_VPWR_c_365_n 0.0162794f $X=0.965 $Y=2.465 $X2=0
+ $Y2=0
cc_124 N_A_85_21#_c_76_n N_VPWR_c_365_n 0.00390745f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_125 N_A_85_21#_c_77_n N_VPWR_c_365_n 5.65397e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_126 N_A_85_21#_c_109_p N_VPWR_c_366_n 0.00976044f $X=3.485 $Y=2.01 $X2=0
+ $Y2=0
cc_127 N_A_85_21#_c_86_n N_VPWR_c_366_n 0.00807522f $X=3.9 $Y=2.095 $X2=0 $Y2=0
cc_128 N_A_85_21#_c_105_p N_VPWR_c_367_n 0.0163512f $X=3 $Y=2.91 $X2=0 $Y2=0
cc_129 N_A_85_21#_c_85_n N_VPWR_c_369_n 0.0178111f $X=3.9 $Y=2.91 $X2=0 $Y2=0
cc_130 N_A_85_21#_M1005_d N_VPWR_c_361_n 0.0116735f $X=2.675 $Y=1.835 $X2=0
+ $Y2=0
cc_131 N_A_85_21#_M1001_d N_VPWR_c_361_n 0.00371702f $X=3.76 $Y=1.835 $X2=0
+ $Y2=0
cc_132 N_A_85_21#_M1003_g N_VPWR_c_361_n 0.0110936f $X=0.535 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_85_21#_M1011_g N_VPWR_c_361_n 0.0106603f $X=0.965 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_85_21#_c_105_p N_VPWR_c_361_n 0.00925289f $X=3 $Y=2.91 $X2=0 $Y2=0
cc_135 N_A_85_21#_c_85_n N_VPWR_c_361_n 0.0100304f $X=3.9 $Y=2.91 $X2=0 $Y2=0
cc_136 N_A_85_21#_M1003_g X 0.00715749f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_85_21#_M1011_g X 0.00983015f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A_85_21#_M1003_g X 0.0140624f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_85_21#_M1011_g X 0.0172125f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A_85_21#_c_72_n N_X_c_418_n 0.00312861f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_141 N_A_85_21#_M1003_g N_X_c_418_n 0.00874843f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_85_21#_c_74_n N_X_c_418_n 0.00139492f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_143 N_A_85_21#_M1011_g N_X_c_418_n 0.00235775f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_85_21#_c_76_n N_X_c_418_n 0.0241762f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_145 N_A_85_21#_c_77_n N_X_c_418_n 0.0291805f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_146 N_A_85_21#_c_161_p N_X_c_418_n 0.0110373f $X=1.235 $Y=1.09 $X2=0 $Y2=0
cc_147 N_A_85_21#_c_78_n N_VGND_M1013_d 0.00364762f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_148 N_A_85_21#_c_161_p N_VGND_M1013_d 0.00188677f $X=1.235 $Y=1.09 $X2=0
+ $Y2=0
cc_149 N_A_85_21#_c_78_n N_VGND_M1004_d 0.00312804f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_150 N_A_85_21#_c_72_n N_VGND_c_446_n 0.0071233f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_151 N_A_85_21#_c_72_n N_VGND_c_447_n 6.38919e-19 $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_152 N_A_85_21#_c_74_n N_VGND_c_447_n 0.0112232f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A_85_21#_c_77_n N_VGND_c_447_n 0.00106436f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_154 N_A_85_21#_c_78_n N_VGND_c_447_n 0.028842f $X=3.485 $Y=1.09 $X2=0 $Y2=0
cc_155 N_A_85_21#_c_161_p N_VGND_c_447_n 0.0172198f $X=1.235 $Y=1.09 $X2=0 $Y2=0
cc_156 N_A_85_21#_c_72_n N_VGND_c_449_n 0.00583607f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_157 N_A_85_21#_c_74_n N_VGND_c_449_n 0.00486043f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_158 N_A_85_21#_c_80_n N_VGND_c_451_n 0.0335572f $X=3.895 $Y=0.42 $X2=0 $Y2=0
cc_159 N_A_85_21#_M1007_d N_VGND_c_452_n 0.00215158f $X=3.755 $Y=0.235 $X2=0
+ $Y2=0
cc_160 N_A_85_21#_c_72_n N_VGND_c_452_n 0.011437f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_161 N_A_85_21#_c_74_n N_VGND_c_452_n 0.00824727f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_162 N_A_85_21#_c_80_n N_VGND_c_452_n 0.0201567f $X=3.895 $Y=0.42 $X2=0 $Y2=0
cc_163 N_A_85_21#_c_78_n N_A_355_47#_M1009_d 0.00297626f $X=3.485 $Y=1.09
+ $X2=-0.19 $Y2=-0.245
cc_164 N_A_85_21#_c_78_n N_A_355_47#_M1002_d 0.00304851f $X=3.485 $Y=1.09 $X2=0
+ $Y2=0
cc_165 N_A_85_21#_c_78_n N_A_355_47#_c_503_n 0.0217646f $X=3.485 $Y=1.09 $X2=0
+ $Y2=0
cc_166 N_A_85_21#_c_78_n N_A_355_47#_c_504_n 0.0406763f $X=3.485 $Y=1.09 $X2=0
+ $Y2=0
cc_167 N_A_85_21#_c_78_n N_A_355_47#_c_505_n 0.0221661f $X=3.485 $Y=1.09 $X2=0
+ $Y2=0
cc_168 N_A_85_21#_c_78_n A_679_47# 0.00122098f $X=3.485 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_85_21#_c_80_n A_679_47# 0.00873102f $X=3.895 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A_85_21#_c_81_n A_679_47# 0.00157887f $X=3.485 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A1_M1009_g N_A2_c_225_n 0.0576808f $X=1.7 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_172 N_A1_c_188_n N_A2_c_225_n 0.00198717f $X=1.712 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_173 A1 N_A2_M1008_g 0.00374202f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_174 N_A1_c_187_n N_A2_M1008_g 0.0576808f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_175 N_A1_M1009_g N_A2_M1004_g 0.0260519f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_176 N_A1_M1000_g N_A2_c_229_n 0.00140689f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_177 A1 N_A2_c_229_n 0.0531571f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A1_c_187_n N_A2_c_229_n 3.67042e-19 $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A1_c_188_n N_A2_c_229_n 0.0270219f $X=1.712 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A1_M1000_g N_VPWR_c_365_n 0.00997066f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A1_M1000_g N_VPWR_c_367_n 0.00380566f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_182 A1 N_VPWR_c_367_n 0.0075296f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_183 N_A1_M1000_g N_VPWR_c_361_n 0.00597216f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_184 A1 N_VPWR_c_361_n 0.00777135f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A1_c_188_n N_X_c_418_n 0.0047978f $X=1.712 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A1_M1009_g N_VGND_c_447_n 0.0124669f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_187 N_A1_M1009_g N_VGND_c_450_n 0.00486043f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A1_M1009_g N_VGND_c_452_n 0.00863238f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A2_M1008_g N_A3_M1005_g 0.0464155f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A2_c_229_n N_A3_M1005_g 0.00430887f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A2_M1004_g N_A3_M1002_g 0.0332145f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A2_c_225_n N_A3_c_261_n 0.0205991f $X=2.06 $Y=1.675 $X2=0 $Y2=0
cc_193 N_A2_c_229_n N_A3_c_261_n 3.66933e-19 $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_194 N_A2_c_225_n N_A3_c_262_n 0.0018999f $X=2.06 $Y=1.675 $X2=0 $Y2=0
cc_195 N_A2_M1008_g N_A3_c_262_n 0.0012205f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A2_c_229_n N_A3_c_262_n 0.0835842f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_197 N_A2_M1008_g N_VPWR_c_367_n 0.00402414f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A2_c_229_n N_VPWR_c_367_n 0.010856f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_199 N_A2_M1008_g N_VPWR_c_361_n 0.00620519f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A2_c_229_n N_VPWR_c_361_n 0.0104031f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_201 N_A2_c_229_n A_427_367# 0.0111394f $X=2.15 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_202 N_A2_M1004_g N_VGND_c_447_n 0.00108039f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_203 N_A2_M1004_g N_VGND_c_448_n 0.00471922f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_204 N_A2_M1004_g N_VGND_c_450_n 0.00429465f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_205 N_A2_M1004_g N_VGND_c_452_n 0.00640365f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_206 N_A2_M1004_g N_A_355_47#_c_504_n 0.0104796f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_207 N_A3_M1005_g N_B1_M1006_g 0.0187188f $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_208 A3 N_B1_M1006_g 0.00168582f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_209 N_A3_M1002_g N_B1_M1010_g 0.017034f $X=2.78 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A3_c_261_n N_B1_c_299_n 0.0205033f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_211 N_A3_c_262_n N_B1_c_299_n 3.23552e-19 $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_212 N_A3_M1005_g N_B1_c_300_n 2.39865e-19 $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_213 A3 N_B1_c_300_n 8.93167e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_214 N_A3_c_261_n N_B1_c_300_n 0.00203862f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_215 N_A3_c_262_n N_B1_c_300_n 0.0311812f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_216 N_A3_M1005_g N_VPWR_c_366_n 8.52912e-19 $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A3_M1005_g N_VPWR_c_367_n 0.00380566f $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_218 A3 N_VPWR_c_367_n 0.0078493f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A3_M1005_g N_VPWR_c_361_n 0.00629888f $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_220 A3 N_VPWR_c_361_n 0.00831863f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_221 N_A3_M1002_g N_VGND_c_448_n 0.00322656f $X=2.78 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A3_M1002_g N_VGND_c_451_n 0.00429465f $X=2.78 $Y=0.655 $X2=0 $Y2=0
cc_223 N_A3_M1002_g N_VGND_c_452_n 0.00630384f $X=2.78 $Y=0.655 $X2=0 $Y2=0
cc_224 N_A3_M1002_g N_A_355_47#_c_504_n 0.0104796f $X=2.78 $Y=0.655 $X2=0 $Y2=0
cc_225 N_B1_M1010_g N_C1_M1007_g 0.0406408f $X=3.32 $Y=0.655 $X2=0 $Y2=0
cc_226 N_B1_M1006_g N_C1_M1001_g 0.0355299f $X=3.255 $Y=2.465 $X2=0 $Y2=0
cc_227 N_B1_c_299_n N_C1_c_336_n 0.0544415f $X=3.23 $Y=1.51 $X2=0 $Y2=0
cc_228 N_B1_c_300_n N_C1_c_336_n 3.61249e-19 $X=3.23 $Y=1.51 $X2=0 $Y2=0
cc_229 N_B1_M1006_g N_VPWR_c_366_n 0.0160595f $X=3.255 $Y=2.465 $X2=0 $Y2=0
cc_230 N_B1_M1006_g N_VPWR_c_367_n 0.00486043f $X=3.255 $Y=2.465 $X2=0 $Y2=0
cc_231 N_B1_M1006_g N_VPWR_c_361_n 0.00872112f $X=3.255 $Y=2.465 $X2=0 $Y2=0
cc_232 N_B1_M1010_g N_VGND_c_451_n 0.00585385f $X=3.32 $Y=0.655 $X2=0 $Y2=0
cc_233 N_B1_M1010_g N_VGND_c_452_n 0.0109726f $X=3.32 $Y=0.655 $X2=0 $Y2=0
cc_234 N_C1_M1001_g N_VPWR_c_366_n 0.016474f $X=3.685 $Y=2.465 $X2=0 $Y2=0
cc_235 N_C1_M1001_g N_VPWR_c_369_n 0.00486043f $X=3.685 $Y=2.465 $X2=0 $Y2=0
cc_236 N_C1_M1001_g N_VPWR_c_361_n 0.00930006f $X=3.685 $Y=2.465 $X2=0 $Y2=0
cc_237 N_C1_M1007_g N_VGND_c_451_n 0.00357668f $X=3.68 $Y=0.655 $X2=0 $Y2=0
cc_238 N_C1_M1007_g N_VGND_c_452_n 0.00623883f $X=3.68 $Y=0.655 $X2=0 $Y2=0
cc_239 N_VPWR_c_361_n N_X_M1003_s 0.00223559f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_240 N_VPWR_c_363_n X 0.0477854f $X=0.32 $Y=1.98 $X2=0 $Y2=0
cc_241 N_VPWR_c_364_n X 0.0182419f $X=1.155 $Y=3.33 $X2=0 $Y2=0
cc_242 N_VPWR_c_365_n X 0.0713718f $X=1.32 $Y=2.02 $X2=0 $Y2=0
cc_243 N_VPWR_c_361_n X 0.0120429f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_361_n A_355_367# 0.00714082f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_245 N_VPWR_c_361_n A_427_367# 0.00923159f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_246 N_X_c_418_n N_VGND_c_446_n 0.0286552f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_247 N_X_c_418_n N_VGND_c_449_n 0.0133395f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_248 N_X_M1012_s N_VGND_c_452_n 0.00449678f $X=0.575 $Y=0.235 $X2=0 $Y2=0
cc_249 N_X_c_418_n N_VGND_c_452_n 0.00828095f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_250 N_VGND_c_452_n N_A_355_47#_M1009_d 0.0047248f $X=4.08 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_251 N_VGND_c_452_n N_A_355_47#_M1002_d 0.0042825f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_252 N_VGND_c_450_n N_A_355_47#_c_510_n 0.020857f $X=2.345 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_452_n N_A_355_47#_c_510_n 0.0126991f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_M1004_d N_A_355_47#_c_504_n 0.00606424f $X=2.31 $Y=0.235 $X2=0
+ $Y2=0
cc_255 N_VGND_c_448_n N_A_355_47#_c_504_n 0.0216197f $X=2.51 $Y=0.37 $X2=0 $Y2=0
cc_256 N_VGND_c_450_n N_A_355_47#_c_504_n 0.00267881f $X=2.345 $Y=0 $X2=0 $Y2=0
cc_257 N_VGND_c_451_n N_A_355_47#_c_504_n 0.00281453f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_452_n N_A_355_47#_c_504_n 0.011034f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_259 N_VGND_c_451_n N_A_355_47#_c_517_n 0.0210271f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_260 N_VGND_c_452_n N_A_355_47#_c_517_n 0.0126991f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_261 N_VGND_c_452_n A_679_47# 0.00607198f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
