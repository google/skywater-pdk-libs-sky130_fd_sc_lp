* File: sky130_fd_sc_lp__a2bb2o_0.pex.spice
* Created: Fri Aug 28 09:55:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%A_59_194# 1 2 8 11 13 14 17 19 25 26 27 29
+ 35 37 38 42
c101 37 0 1.24193e-19 $X=2.34 $Y=2.075
r102 37 38 9.23804 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=2.34 $Y=2.075
+ $X2=2.34 $Y2=2.245
r103 33 35 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=0.445
+ $X2=2.41 $Y2=0.445
r104 30 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=0.61
+ $X2=2.41 $Y2=0.445
r105 30 37 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=2.41 $Y=0.61
+ $X2=2.41 $Y2=2.075
r106 29 40 2.96548 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.302 $Y=2.88
+ $X2=2.302 $Y2=2.965
r107 29 38 31.1405 $w=2.33e-07 $l=6.35e-07 $layer=LI1_cond $X=2.302 $Y=2.88
+ $X2=2.302 $Y2=2.245
r108 26 40 4.08189 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.185 $Y=2.965
+ $X2=2.302 $Y2=2.965
r109 26 27 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.185 $Y=2.965
+ $X2=1.31 $Y2=2.965
r110 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.225 $Y=2.88
+ $X2=1.31 $Y2=2.965
r111 24 25 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.225 $Y=2.26
+ $X2=1.225 $Y2=2.88
r112 22 42 16.2954 $w=2.81e-07 $l=9.5e-08 $layer=POLY_cond $X=0.59 $Y=2.095
+ $X2=0.495 $Y2=2.095
r113 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=2.095 $X2=0.59 $Y2=2.095
r114 19 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=2.095
+ $X2=1.225 $Y2=2.26
r115 19 21 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=1.14 $Y=2.095
+ $X2=0.59 $Y2=2.095
r116 15 17 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=0.68 $Y=0.97
+ $X2=0.68 $Y2=0.445
r117 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.605 $Y=1.045
+ $X2=0.68 $Y2=0.97
r118 13 14 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.605 $Y=1.045
+ $X2=0.445 $Y2=1.045
r119 9 42 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=2.26
+ $X2=0.495 $Y2=2.095
r120 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.495 $Y=2.26
+ $X2=0.495 $Y2=2.77
r121 8 42 21.4413 $w=2.81e-07 $l=2.18746e-07 $layer=POLY_cond $X=0.37 $Y=1.93
+ $X2=0.495 $Y2=2.095
r122 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.37 $Y=1.12
+ $X2=0.445 $Y2=1.045
r123 7 8 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.37 $Y=1.12 $X2=0.37
+ $Y2=1.93
r124 2 40 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=2.165
+ $Y=2.675 $X2=2.29 $Y2=2.885
r125 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.185
+ $Y=0.235 $X2=2.325 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%A1_N 2 5 9 10 11 12 13 14 22
c58 11 0 1.9296e-19 $X=1.075 $Y=0.915
r59 19 22 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.85 $Y=1.525
+ $X2=1.04 $Y2=1.525
r60 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.85
+ $Y=1.525 $X2=0.85 $Y2=1.525
r61 14 20 3.98375 $w=4.03e-07 $l=1.4e-07 $layer=LI1_cond $X=0.732 $Y=1.665
+ $X2=0.732 $Y2=1.525
r62 13 20 6.54474 $w=4.03e-07 $l=2.3e-07 $layer=LI1_cond $X=0.732 $Y=1.295
+ $X2=0.732 $Y2=1.525
r63 12 13 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.732 $Y=0.925
+ $X2=0.732 $Y2=1.295
r64 10 11 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.075 $Y=0.765
+ $X2=1.075 $Y2=0.915
r65 9 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.11 $Y=0.445
+ $X2=1.11 $Y2=0.765
r66 3 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.69
+ $X2=1.04 $Y2=1.525
r67 3 5 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=1.04 $Y=1.69 $X2=1.04
+ $Y2=2.66
r68 2 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.36
+ $X2=1.04 $Y2=1.525
r69 2 11 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.04 $Y=1.36
+ $X2=1.04 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%A2_N 3 7 11 12 13 14 18
c52 11 0 1.4009e-19 $X=1.49 $Y=1.66
r53 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.49
+ $Y=1.32 $X2=1.49 $Y2=1.32
r54 14 19 7.50267 $w=5.48e-07 $l=3.45e-07 $layer=LI1_cond $X=1.38 $Y=1.665
+ $X2=1.38 $Y2=1.32
r55 13 19 0.543672 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=1.38 $Y=1.295
+ $X2=1.38 $Y2=1.32
r56 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.49 $Y=1.66
+ $X2=1.49 $Y2=1.32
r57 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.66
+ $X2=1.49 $Y2=1.825
r58 10 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.155
+ $X2=1.49 $Y2=1.32
r59 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.55 $Y=0.445
+ $X2=1.55 $Y2=1.155
r60 3 12 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=1.43 $Y=2.66 $X2=1.43
+ $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%A_237_47# 1 2 9 12 13 14 17 21 22 25 27 28
+ 29 35 38 39 41 42 43
r84 41 43 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.92 $Y=2.43
+ $X2=1.92 $Y2=1.905
r85 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.06 $Y=1.4
+ $X2=2.06 $Y2=1.4
r86 36 43 8.28018 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=1.995 $Y=1.745
+ $X2=1.995 $Y2=1.905
r87 36 38 12.4248 $w=3.18e-07 $l=3.45e-07 $layer=LI1_cond $X=1.995 $Y=1.745
+ $X2=1.995 $Y2=1.4
r88 35 42 8.28018 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=1.995 $Y=1.395
+ $X2=1.995 $Y2=1.235
r89 35 38 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=1.995 $Y=1.395
+ $X2=1.995 $Y2=1.4
r90 33 42 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.92 $Y=0.975
+ $X2=1.92 $Y2=1.235
r91 29 41 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.835 $Y=2.57
+ $X2=1.92 $Y2=2.43
r92 29 31 7.82015 $w=2.78e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=2.57
+ $X2=1.645 $Y2=2.57
r93 27 33 6.85817 $w=1.95e-07 $l=1.33918e-07 $layer=LI1_cond $X=1.835 $Y=0.877
+ $X2=1.92 $Y2=0.975
r94 27 28 21.0443 $w=1.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.835 $Y=0.877
+ $X2=1.465 $Y2=0.877
r95 23 28 7.04969 $w=1.95e-07 $l=1.76975e-07 $layer=LI1_cond $X=1.33 $Y=0.78
+ $X2=1.465 $Y2=0.877
r96 23 25 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.33 $Y=0.78
+ $X2=1.33 $Y2=0.445
r97 21 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.06 $Y=1.74
+ $X2=2.06 $Y2=1.4
r98 21 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.74
+ $X2=2.06 $Y2=1.905
r99 20 39 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.235
+ $X2=2.06 $Y2=1.4
r100 15 17 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.505 $Y=2.215
+ $X2=2.505 $Y2=2.885
r101 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.43 $Y=2.14
+ $X2=2.505 $Y2=2.215
r102 13 14 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.43 $Y=2.14
+ $X2=2.225 $Y2=2.14
r103 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.15 $Y=2.065
+ $X2=2.225 $Y2=2.14
r104 12 22 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.15 $Y=2.065
+ $X2=2.15 $Y2=1.905
r105 9 20 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.11 $Y=0.445
+ $X2=2.11 $Y2=1.235
r106 2 31 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=2.45 $X2=1.645 $Y2=2.605
r107 1 25 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=1.185
+ $Y=0.235 $X2=1.335 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%B2 3 7 9 10 11 12 18
c42 18 0 1.22418e-19 $X=2.845 $Y=1.32
r43 18 21 81.2291 $w=5.45e-07 $l=5.05e-07 $layer=POLY_cond $X=2.737 $Y=1.32
+ $X2=2.737 $Y2=1.825
r44 18 20 47.8511 $w=5.45e-07 $l=1.65e-07 $layer=POLY_cond $X=2.737 $Y=1.32
+ $X2=2.737 $Y2=1.155
r45 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.845
+ $Y=1.32 $X2=2.845 $Y2=1.32
r46 11 12 9.03161 $w=4.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.005 $Y=1.665
+ $X2=3.005 $Y2=2.035
r47 11 19 8.42137 $w=4.88e-07 $l=3.45e-07 $layer=LI1_cond $X=3.005 $Y=1.665
+ $X2=3.005 $Y2=1.32
r48 10 19 0.610244 $w=4.88e-07 $l=2.5e-08 $layer=LI1_cond $X=3.005 $Y=1.295
+ $X2=3.005 $Y2=1.32
r49 9 10 9.03161 $w=4.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.005 $Y=0.925
+ $X2=3.005 $Y2=1.295
r50 7 21 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=2.935 $Y=2.885
+ $X2=2.935 $Y2=1.825
r51 3 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.54 $Y=0.445
+ $X2=2.54 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%B1 1 3 4 5 8 12 13 14 15 16 17 24
c36 5 0 1.24193e-19 $X=3.005 $Y=0.84
r37 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.515
+ $Y=1.12 $X2=3.515 $Y2=1.12
r38 16 17 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=1.665
+ $X2=3.587 $Y2=2.035
r39 15 16 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=1.295
+ $X2=3.587 $Y2=1.665
r40 15 25 6.02022 $w=3.33e-07 $l=1.75e-07 $layer=LI1_cond $X=3.587 $Y=1.295
+ $X2=3.587 $Y2=1.12
r41 14 25 6.70825 $w=3.33e-07 $l=1.95e-07 $layer=LI1_cond $X=3.587 $Y=0.925
+ $X2=3.587 $Y2=1.12
r42 13 14 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=0.555
+ $X2=3.587 $Y2=0.925
r43 11 24 44.2071 $w=3.9e-07 $l=3.1e-07 $layer=POLY_cond $X=3.485 $Y=1.43
+ $X2=3.485 $Y2=1.12
r44 11 12 49.7341 $w=3.9e-07 $l=1.95e-07 $layer=POLY_cond $X=3.485 $Y=1.43
+ $X2=3.485 $Y2=1.625
r45 10 24 29.2337 $w=3.9e-07 $l=2.05e-07 $layer=POLY_cond $X=3.485 $Y=0.915
+ $X2=3.485 $Y2=1.12
r46 8 12 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=3.365 $Y=2.885
+ $X2=3.365 $Y2=1.625
r47 4 10 34.5134 $w=1.5e-07 $l=2.29456e-07 $layer=POLY_cond $X=3.29 $Y=0.84
+ $X2=3.485 $Y2=0.915
r48 4 5 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.29 $Y=0.84
+ $X2=3.005 $Y2=0.84
r49 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.93 $Y=0.765
+ $X2=3.005 $Y2=0.84
r50 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.93 $Y=0.765 $X2=2.93
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%X 1 2 11 13 14 15 16 17 18 37
r27 38 45 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2.61
+ $X2=0.265 $Y2=2.595
r28 37 43 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=0.21 $Y=2.405
+ $X2=0.21 $Y2=2.43
r29 18 38 5.28203 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.775
+ $X2=0.265 $Y2=2.61
r30 17 45 4.32166 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.265 $Y=2.46
+ $X2=0.265 $Y2=2.595
r31 17 43 2.04773 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=0.265 $Y=2.46
+ $X2=0.265 $Y2=2.43
r32 17 37 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=0.21 $Y=2.375 $X2=0.21
+ $Y2=2.405
r33 16 17 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.21 $Y=2.035
+ $X2=0.21 $Y2=2.375
r34 15 16 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=2.035
r35 14 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.295
+ $X2=0.21 $Y2=1.665
r36 13 14 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=0.925
+ $X2=0.21 $Y2=1.295
r37 8 13 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.21 $Y=0.61
+ $X2=0.21 $Y2=0.925
r38 7 11 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.21 $Y=0.445
+ $X2=0.465 $Y2=0.445
r39 7 8 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.21 $Y=0.445 $X2=0.21
+ $Y2=0.61
r40 2 45 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=2.45 $X2=0.28 $Y2=2.595
r41 1 11 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.235 $X2=0.465 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%VPWR 1 2 9 13 15 17 22 32 33 36 39
r50 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r54 30 39 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.285 $Y=3.33
+ $X2=3.152 $Y2=3.33
r55 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.285 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 23 36 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.792 $Y2=3.33
r62 23 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33 $X2=1.2
+ $Y2=3.33
r63 22 39 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=3.152 $Y2=3.33
r64 22 28 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r67 17 36 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.792 $Y2=3.33
r68 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r70 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r71 11 39 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.152 $Y=3.245
+ $X2=3.152 $Y2=3.33
r72 11 13 14.1337 $w=2.63e-07 $l=3.25e-07 $layer=LI1_cond $X=3.152 $Y=3.245
+ $X2=3.152 $Y2=2.92
r73 7 36 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.792 $Y=3.245
+ $X2=0.792 $Y2=3.33
r74 7 9 21.1011 $w=3.53e-07 $l=6.5e-07 $layer=LI1_cond $X=0.792 $Y=3.245
+ $X2=0.792 $Y2=2.595
r75 2 13 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=2.675 $X2=3.15 $Y2=2.92
r76 1 9 300 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=2.45 $X2=0.825 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%A_516_535# 1 2 9 11 12 15
c26 11 0 1.11547e-19 $X=3.455 $Y=2.5
r27 13 15 11.9218 $w=2.88e-07 $l=3e-07 $layer=LI1_cond $X=3.6 $Y=2.585 $X2=3.6
+ $Y2=2.885
r28 11 13 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=3.455 $Y=2.5
+ $X2=3.6 $Y2=2.585
r29 11 12 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.455 $Y=2.5
+ $X2=2.825 $Y2=2.5
r30 7 12 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=2.707 $Y=2.585
+ $X2=2.825 $Y2=2.5
r31 7 9 14.712 $w=2.33e-07 $l=3e-07 $layer=LI1_cond $X=2.707 $Y=2.585 $X2=2.707
+ $Y2=2.885
r32 2 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=2.675 $X2=3.58 $Y2=2.885
r33 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=2.675 $X2=2.72 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_0%VGND 1 2 3 12 14 18 22 24 25 26 32 39 40 43
+ 46
c55 22 0 1.08719e-20 $X=3.145 $Y=0.445
c56 14 0 1.9296e-19 $X=1.66 $Y=0
r57 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r58 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r59 40 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r60 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r61 37 46 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.115
+ $Y2=0
r62 37 39 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.6
+ $Y2=0
r63 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r64 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r65 33 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=0 $X2=1.825
+ $Y2=0
r66 33 35 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.99 $Y=0 $X2=2.64
+ $Y2=0
r67 32 46 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.98 $Y=0 $X2=3.115
+ $Y2=0
r68 32 35 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.98 $Y=0 $X2=2.64
+ $Y2=0
r69 30 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r70 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r71 26 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r72 26 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r73 24 29 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.72
+ $Y2=0
r74 24 25 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.895
+ $Y2=0
r75 20 46 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0.085
+ $X2=3.115 $Y2=0
r76 20 22 15.3659 $w=2.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.115 $Y=0.085
+ $X2=3.115 $Y2=0.445
r77 16 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=0.085
+ $X2=1.825 $Y2=0
r78 16 18 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.825 $Y=0.085
+ $X2=1.825 $Y2=0.445
r79 15 25 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=0.895
+ $Y2=0
r80 14 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=0 $X2=1.825
+ $Y2=0
r81 14 15 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.66 $Y=0 $X2=1.025
+ $Y2=0
r82 10 25 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0
r83 10 12 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0.445
r84 3 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.005
+ $Y=0.235 $X2=3.145 $Y2=0.445
r85 2 18 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.235 $X2=1.825 $Y2=0.445
r86 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.755
+ $Y=0.235 $X2=0.895 $Y2=0.445
.ends

