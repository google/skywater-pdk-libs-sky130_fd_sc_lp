* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21o_lp A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR a_218_57# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_218_57# B1 a_332_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_490_57# a_218_57# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND A2 a_140_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_332_57# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR A1 a_33_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VGND a_218_57# a_490_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_140_57# A1 a_218_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_33_409# B1 a_218_57# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_33_409# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
