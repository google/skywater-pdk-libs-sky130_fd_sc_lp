* File: sky130_fd_sc_lp__nor2_2.pxi.spice
* Created: Wed Sep  2 10:07:30 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2_2%A N_A_c_42_n N_A_M1000_g N_A_M1003_g N_A_c_44_n
+ N_A_M1002_g N_A_M1006_g A A N_A_c_47_n PM_SKY130_FD_SC_LP__NOR2_2%A
x_PM_SKY130_FD_SC_LP__NOR2_2%B N_B_M1001_g N_B_M1005_g N_B_M1004_g N_B_M1007_g B
+ B N_B_c_87_n N_B_c_88_n PM_SKY130_FD_SC_LP__NOR2_2%B
x_PM_SKY130_FD_SC_LP__NOR2_2%A_28_367# N_A_28_367#_M1003_d N_A_28_367#_M1006_d
+ N_A_28_367#_M1007_d N_A_28_367#_c_135_n N_A_28_367#_c_136_n
+ N_A_28_367#_c_141_n N_A_28_367#_c_146_n N_A_28_367#_c_153_p
+ N_A_28_367#_c_147_n N_A_28_367#_c_137_n N_A_28_367#_c_138_n
+ PM_SKY130_FD_SC_LP__NOR2_2%A_28_367#
x_PM_SKY130_FD_SC_LP__NOR2_2%VPWR N_VPWR_M1003_s N_VPWR_c_168_n VPWR
+ N_VPWR_c_169_n N_VPWR_c_170_n N_VPWR_c_167_n N_VPWR_c_172_n
+ PM_SKY130_FD_SC_LP__NOR2_2%VPWR
x_PM_SKY130_FD_SC_LP__NOR2_2%Y N_Y_M1000_d N_Y_M1001_s N_Y_M1005_s N_Y_c_233_p
+ N_Y_c_198_n N_Y_c_199_n N_Y_c_212_n N_Y_c_200_n N_Y_c_201_n Y Y N_Y_c_225_n
+ PM_SKY130_FD_SC_LP__NOR2_2%Y
x_PM_SKY130_FD_SC_LP__NOR2_2%VGND N_VGND_M1000_s N_VGND_M1002_s N_VGND_M1004_d
+ N_VGND_c_239_n N_VGND_c_240_n N_VGND_c_241_n N_VGND_c_242_n N_VGND_c_243_n
+ VGND N_VGND_c_244_n N_VGND_c_245_n N_VGND_c_246_n N_VGND_c_247_n
+ PM_SKY130_FD_SC_LP__NOR2_2%VGND
cc_1 VNB N_A_c_42_n 0.022383f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.21
cc_2 VNB N_A_M1003_g 0.00703465f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_3 VNB N_A_c_44_n 0.015724f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.21
cc_4 VNB N_A_M1006_g 0.00449224f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_5 VNB A 0.0201069f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A_c_47_n 0.0611464f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.375
cc_7 VNB N_B_M1001_g 0.0223637f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.665
cc_8 VNB N_B_M1004_g 0.0285775f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.54
cc_9 VNB N_B_c_87_n 0.00263028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_88_n 0.0378989f $X=-0.19 $Y=-0.245 $X2=0.257 $Y2=1.295
cc_11 VNB N_VPWR_c_167_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.375
cc_12 VNB N_Y_c_198_n 0.00838219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_Y_c_199_n 0.00133475f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_Y_c_200_n 0.0141043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_201_n 0.00947429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_239_n 0.010601f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.665
cc_17 VNB N_VGND_c_240_n 0.0341382f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_18 VNB N_VGND_c_241_n 5.00113e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_VGND_c_242_n 0.0138645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_243_n 0.0312168f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.375
cc_21 VNB N_VGND_c_244_n 0.0131655f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.375
cc_22 VNB N_VGND_c_245_n 0.0164909f $X=-0.19 $Y=-0.245 $X2=0.257 $Y2=1.375
cc_23 VNB N_VGND_c_246_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_247_n 0.152471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VPB N_A_M1003_g 0.0258135f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_26 VPB N_A_M1006_g 0.018974f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_27 VPB A 0.00711651f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_28 VPB N_B_M1005_g 0.0183294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_B_M1007_g 0.0230923f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_30 VPB N_B_c_87_n 0.00838131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_B_c_88_n 0.00675374f $X=-0.19 $Y=1.655 $X2=0.257 $Y2=1.295
cc_32 VPB N_A_28_367#_c_135_n 0.00755006f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.665
cc_33 VPB N_A_28_367#_c_136_n 0.0373194f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_34 VPB N_A_28_367#_c_137_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=1.375
cc_35 VPB N_A_28_367#_c_138_n 0.0509193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_168_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_37 VPB N_VPWR_c_169_n 0.015535f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.665
cc_38 VPB N_VPWR_c_170_n 0.0379392f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=1.375
cc_39 VPB N_VPWR_c_167_n 0.0453153f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=1.375
cc_40 VPB N_VPWR_c_172_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.375
cc_41 VPB N_Y_c_200_n 0.00583711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 N_A_c_44_n N_B_M1001_g 0.0233981f $X=0.91 $Y=1.21 $X2=0 $Y2=0
cc_43 N_A_M1006_g N_B_M1005_g 0.0196332f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_44 N_A_M1003_g N_B_c_87_n 0.00171969f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_45 N_A_M1006_g N_B_c_87_n 0.00904129f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_46 A N_B_c_87_n 0.0267681f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_A_c_47_n N_B_c_87_n 0.0144365f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_48 N_A_c_47_n N_B_c_88_n 0.0228959f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_49 A N_A_28_367#_c_135_n 0.0230165f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_50 N_A_c_47_n N_A_28_367#_c_135_n 8.56496e-19 $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_51 N_A_M1003_g N_A_28_367#_c_141_n 0.0160602f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_52 N_A_M1006_g N_A_28_367#_c_141_n 0.0122595f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_53 A N_A_28_367#_c_141_n 0.00378716f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_A_c_47_n N_A_28_367#_c_141_n 4.32697e-19 $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_55 N_A_M1003_g N_VPWR_c_168_n 0.0165482f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_56 N_A_M1006_g N_VPWR_c_168_n 0.0158312f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_57 N_A_M1003_g N_VPWR_c_169_n 0.00486043f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_58 N_A_M1006_g N_VPWR_c_170_n 0.00486043f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A_M1003_g N_VPWR_c_167_n 0.00918457f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_60 N_A_M1006_g N_VPWR_c_167_n 0.0082726f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_61 N_A_c_44_n N_Y_c_198_n 0.0101987f $X=0.91 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A_c_47_n N_Y_c_198_n 0.00398544f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_63 N_A_c_42_n N_Y_c_199_n 0.0039238f $X=0.48 $Y=1.21 $X2=0 $Y2=0
cc_64 A N_Y_c_199_n 0.0034413f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_c_47_n N_Y_c_199_n 0.00650507f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_66 N_A_c_42_n N_VGND_c_240_n 0.0166113f $X=0.48 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A_c_44_n N_VGND_c_240_n 6.66143e-19 $X=0.91 $Y=1.21 $X2=0 $Y2=0
cc_68 A N_VGND_c_240_n 0.0259278f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_c_47_n N_VGND_c_240_n 0.00160808f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_70 N_A_c_42_n N_VGND_c_241_n 6.15775e-19 $X=0.48 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_c_44_n N_VGND_c_241_n 0.0112038f $X=0.91 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_c_42_n N_VGND_c_244_n 0.00477554f $X=0.48 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A_c_44_n N_VGND_c_244_n 0.00477554f $X=0.91 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_c_42_n N_VGND_c_247_n 0.00825815f $X=0.48 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_c_44_n N_VGND_c_247_n 0.00825815f $X=0.91 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B_c_87_n N_A_28_367#_c_141_n 0.0283243f $X=1.36 $Y=1.51 $X2=0 $Y2=0
cc_77 N_B_c_87_n N_A_28_367#_c_146_n 0.0149586f $X=1.36 $Y=1.51 $X2=0 $Y2=0
cc_78 N_B_M1005_g N_A_28_367#_c_147_n 0.0111972f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_79 N_B_M1007_g N_A_28_367#_c_147_n 0.0152065f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_80 N_B_M1007_g N_A_28_367#_c_138_n 0.0207522f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_81 N_B_M1005_g N_VPWR_c_168_n 0.00109252f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_82 N_B_M1005_g N_VPWR_c_170_n 0.00357877f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_83 N_B_M1007_g N_VPWR_c_170_n 0.00357877f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_84 N_B_M1005_g N_VPWR_c_167_n 0.00537654f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_85 N_B_M1007_g N_VPWR_c_167_n 0.00655255f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_86 N_B_M1001_g N_Y_c_198_n 0.0142565f $X=1.34 $Y=0.665 $X2=0 $Y2=0
cc_87 N_B_c_87_n N_Y_c_198_n 0.0497985f $X=1.36 $Y=1.51 $X2=0 $Y2=0
cc_88 N_B_c_88_n N_Y_c_198_n 0.0017253f $X=1.77 $Y=1.51 $X2=0 $Y2=0
cc_89 N_B_c_87_n N_Y_c_199_n 0.0143526f $X=1.36 $Y=1.51 $X2=0 $Y2=0
cc_90 N_B_M1005_g N_Y_c_212_n 0.0118179f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B_M1007_g N_Y_c_212_n 0.0233545f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_92 N_B_c_87_n N_Y_c_212_n 0.00963602f $X=1.36 $Y=1.51 $X2=0 $Y2=0
cc_93 N_B_c_88_n N_Y_c_212_n 0.00231438f $X=1.77 $Y=1.51 $X2=0 $Y2=0
cc_94 N_B_M1001_g N_Y_c_200_n 2.46562e-19 $X=1.34 $Y=0.665 $X2=0 $Y2=0
cc_95 N_B_M1005_g N_Y_c_200_n 7.16468e-19 $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_96 N_B_M1004_g N_Y_c_200_n 0.00301053f $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_97 N_B_M1007_g N_Y_c_200_n 0.0085414f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_98 N_B_c_87_n N_Y_c_200_n 0.0250011f $X=1.36 $Y=1.51 $X2=0 $Y2=0
cc_99 N_B_c_88_n N_Y_c_200_n 0.0162233f $X=1.77 $Y=1.51 $X2=0 $Y2=0
cc_100 N_B_M1004_g N_Y_c_201_n 0.011326f $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_101 N_B_c_87_n N_Y_c_201_n 0.00547665f $X=1.36 $Y=1.51 $X2=0 $Y2=0
cc_102 N_B_c_88_n N_Y_c_201_n 0.0031956f $X=1.77 $Y=1.51 $X2=0 $Y2=0
cc_103 N_B_M1004_g N_Y_c_225_n 0.0185464f $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_104 N_B_M1001_g N_VGND_c_241_n 0.0114405f $X=1.34 $Y=0.665 $X2=0 $Y2=0
cc_105 N_B_M1004_g N_VGND_c_241_n 7.172e-19 $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_106 N_B_M1004_g N_VGND_c_243_n 0.00484468f $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_107 N_B_M1001_g N_VGND_c_245_n 0.00477554f $X=1.34 $Y=0.665 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_VGND_c_245_n 0.00472057f $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_109 N_B_M1001_g N_VGND_c_247_n 0.00825815f $X=1.34 $Y=0.665 $X2=0 $Y2=0
cc_110 N_B_M1004_g N_VGND_c_247_n 0.0092838f $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_111 N_A_28_367#_c_141_n N_VPWR_M1003_s 0.00337584f $X=1.03 $Y=2.005 $X2=-0.19
+ $Y2=1.655
cc_112 N_A_28_367#_c_141_n N_VPWR_c_168_n 0.0170777f $X=1.03 $Y=2.005 $X2=0
+ $Y2=0
cc_113 N_A_28_367#_c_136_n N_VPWR_c_169_n 0.0178111f $X=0.265 $Y=2.91 $X2=0
+ $Y2=0
cc_114 N_A_28_367#_c_153_p N_VPWR_c_170_n 0.0121686f $X=1.12 $Y=2.905 $X2=0
+ $Y2=0
cc_115 N_A_28_367#_c_147_n N_VPWR_c_170_n 0.0459292f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_116 N_A_28_367#_c_137_n N_VPWR_c_170_n 0.0175983f $X=2.17 $Y=2.905 $X2=0
+ $Y2=0
cc_117 N_A_28_367#_M1003_d N_VPWR_c_167_n 0.00371702f $X=0.14 $Y=1.835 $X2=0
+ $Y2=0
cc_118 N_A_28_367#_M1006_d N_VPWR_c_167_n 0.00376627f $X=0.985 $Y=1.835 $X2=0
+ $Y2=0
cc_119 N_A_28_367#_M1007_d N_VPWR_c_167_n 0.00337455f $X=1.845 $Y=1.835 $X2=0
+ $Y2=0
cc_120 N_A_28_367#_c_136_n N_VPWR_c_167_n 0.0100304f $X=0.265 $Y=2.91 $X2=0
+ $Y2=0
cc_121 N_A_28_367#_c_153_p N_VPWR_c_167_n 0.00698742f $X=1.12 $Y=2.905 $X2=0
+ $Y2=0
cc_122 N_A_28_367#_c_147_n N_VPWR_c_167_n 0.0299468f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_123 N_A_28_367#_c_137_n N_VPWR_c_167_n 0.00971414f $X=2.17 $Y=2.905 $X2=0
+ $Y2=0
cc_124 N_A_28_367#_c_147_n N_Y_M1005_s 0.00332344f $X=2.045 $Y=2.99 $X2=0 $Y2=0
cc_125 N_A_28_367#_c_147_n N_Y_c_212_n 0.0166589f $X=2.045 $Y=2.99 $X2=0 $Y2=0
cc_126 N_A_28_367#_c_138_n N_Y_c_212_n 0.0293912f $X=2.13 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A_28_367#_c_138_n N_Y_c_200_n 0.0113262f $X=2.13 $Y=1.985 $X2=0 $Y2=0
cc_128 N_VPWR_c_167_n N_Y_M1005_s 0.00225186f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_129 N_Y_c_198_n N_VGND_c_241_n 0.0207154f $X=1.46 $Y=1.17 $X2=0 $Y2=0
cc_130 N_Y_c_225_n N_VGND_c_243_n 0.0491048f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_131 N_Y_c_233_p N_VGND_c_244_n 0.0120977f $X=0.695 $Y=0.42 $X2=0 $Y2=0
cc_132 N_Y_c_225_n N_VGND_c_245_n 0.0187558f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_133 N_Y_M1000_d N_VGND_c_247_n 0.00571434f $X=0.555 $Y=0.245 $X2=0 $Y2=0
cc_134 N_Y_M1001_s N_VGND_c_247_n 0.00380103f $X=1.415 $Y=0.245 $X2=0 $Y2=0
cc_135 N_Y_c_233_p N_VGND_c_247_n 0.00691495f $X=0.695 $Y=0.42 $X2=0 $Y2=0
cc_136 N_Y_c_225_n N_VGND_c_247_n 0.011391f $X=1.555 $Y=0.42 $X2=0 $Y2=0
