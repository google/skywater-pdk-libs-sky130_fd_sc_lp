* File: sky130_fd_sc_lp__o31a_0.pex.spice
* Created: Wed Sep  2 10:24:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31A_0%A_90_309# 1 2 9 13 17 18 21 22 24 25 28 30 33
+ 34 38
r74 36 38 9.84815 $w=3.28e-07 $l=2.82e-07 $layer=LI1_cond $X=2.9 $Y=0.485
+ $X2=3.182 $Y2=0.485
r75 32 38 4.14273 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=3.182 $Y=0.65
+ $X2=3.182 $Y2=0.485
r76 32 33 83.0319 $w=1.83e-07 $l=1.385e-06 $layer=LI1_cond $X=3.182 $Y=0.65
+ $X2=3.182 $Y2=2.035
r77 31 34 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=2.125
+ $X2=2.28 $Y2=2.125
r78 30 33 6.81816 $w=1.8e-07 $l=1.29399e-07 $layer=LI1_cond $X=3.09 $Y=2.125
+ $X2=3.182 $Y2=2.035
r79 30 31 39.7424 $w=1.78e-07 $l=6.45e-07 $layer=LI1_cond $X=3.09 $Y=2.125
+ $X2=2.445 $Y2=2.125
r80 26 34 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.28 $Y=2.215 $X2=2.28
+ $Y2=2.125
r81 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.28 $Y=2.215
+ $X2=2.28 $Y2=2.55
r82 24 34 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=2.125
+ $X2=2.28 $Y2=2.125
r83 24 25 78.2525 $w=1.78e-07 $l=1.27e-06 $layer=LI1_cond $X=2.115 $Y=2.125
+ $X2=0.845 $Y2=2.125
r84 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.615
+ $Y=1.71 $X2=0.615 $Y2=1.71
r85 19 25 7.49754 $w=1.8e-07 $l=1.97949e-07 $layer=LI1_cond $X=0.687 $Y=2.035
+ $X2=0.845 $Y2=2.125
r86 19 21 11.8903 $w=3.13e-07 $l=3.25e-07 $layer=LI1_cond $X=0.687 $Y=2.035
+ $X2=0.687 $Y2=1.71
r87 17 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.615 $Y=2.05
+ $X2=0.615 $Y2=1.71
r88 17 18 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=2.05
+ $X2=0.615 $Y2=2.215
r89 16 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=1.545
+ $X2=0.615 $Y2=1.71
r90 13 16 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.705 $Y=0.485
+ $X2=0.705 $Y2=1.545
r91 9 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.68 $Y=2.725
+ $X2=0.68 $Y2=2.215
r92 2 28 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.13
+ $Y=2.405 $X2=2.28 $Y2=2.55
r93 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.76
+ $Y=0.275 $X2=2.9 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_0%A1 3 7 11 12 13 14 15 21 23 25
c45 25 0 1.23193e-19 $X=1.2 $Y=1.295
c46 23 0 1.92229e-19 $X=1.182 $Y=1.247
r47 23 25 1.65126 $w=3.33e-07 $l=4.8e-08 $layer=LI1_cond $X=1.182 $Y=1.247
+ $X2=1.182 $Y2=1.295
r48 14 23 0.844561 $w=3.35e-07 $l=1.9e-08 $layer=LI1_cond $X=1.182 $Y=1.228
+ $X2=1.182 $Y2=1.247
r49 14 15 12.1093 $w=3.33e-07 $l=3.52e-07 $layer=LI1_cond $X=1.182 $Y=1.313
+ $X2=1.182 $Y2=1.665
r50 14 25 0.619223 $w=3.33e-07 $l=1.8e-08 $layer=LI1_cond $X=1.182 $Y=1.313
+ $X2=1.182 $Y2=1.295
r51 13 14 12.2811 $w=3.01e-07 $l=3.03e-07 $layer=LI1_cond $X=1.182 $Y=0.925
+ $X2=1.182 $Y2=1.228
r52 13 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.185
+ $Y=1.005 $X2=1.185 $Y2=1.005
r53 11 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.185 $Y=1.345
+ $X2=1.185 $Y2=1.005
r54 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.345
+ $X2=1.185 $Y2=1.51
r55 10 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=0.84
+ $X2=1.185 $Y2=1.005
r56 7 12 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=1.275 $Y=2.725
+ $X2=1.275 $Y2=1.51
r57 3 10 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=1.275 $Y=0.485
+ $X2=1.275 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_0%A2 3 7 11 12 13 14 18
c44 18 0 1.92229e-19 $X=1.725 $Y=1.245
c45 3 0 1.23193e-19 $X=1.695 $Y=2.725
r46 13 14 16.6906 $w=2.88e-07 $l=4.2e-07 $layer=LI1_cond $X=1.665 $Y=1.245
+ $X2=1.665 $Y2=1.665
r47 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.725
+ $Y=1.245 $X2=1.725 $Y2=1.245
r48 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.725 $Y=1.585
+ $X2=1.725 $Y2=1.245
r49 11 12 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.585
+ $X2=1.725 $Y2=1.75
r50 10 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.08
+ $X2=1.725 $Y2=1.245
r51 7 10 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=1.785 $Y=0.485
+ $X2=1.785 $Y2=1.08
r52 3 12 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=1.695 $Y=2.725
+ $X2=1.695 $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_0%A3 3 7 9 12 13 17
r45 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.265
+ $Y=1.36 $X2=2.265 $Y2=1.36
r46 13 18 9.49987 $w=3.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.165 $Y=1.665
+ $X2=2.165 $Y2=1.36
r47 12 18 2.02456 $w=3.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.165 $Y=1.295
+ $X2=2.165 $Y2=1.36
r48 11 17 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.195
+ $X2=2.265 $Y2=1.36
r49 9 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.265 $Y=1.7
+ $X2=2.265 $Y2=1.36
r50 7 11 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.255 $Y=0.485
+ $X2=2.255 $Y2=1.195
r51 1 9 82.2016 $w=2.58e-07 $l=5.3479e-07 $layer=POLY_cond $X=2.055 $Y=2.14
+ $X2=2.265 $Y2=1.7
r52 1 3 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=2.055 $Y=2.14
+ $X2=2.055 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_0%B1 3 7 9 12 15 16 18 19 20 24 25
r43 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.835
+ $Y=1.22 $X2=2.835 $Y2=1.22
r44 19 20 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.72 $Y=1.295
+ $X2=2.72 $Y2=1.665
r45 19 25 2.16083 $w=3.98e-07 $l=7.5e-08 $layer=LI1_cond $X=2.72 $Y=1.295
+ $X2=2.72 $Y2=1.22
r46 17 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.835 $Y=1.56
+ $X2=2.835 $Y2=1.22
r47 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.56
+ $X2=2.835 $Y2=1.725
r48 16 24 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=2.835 $Y=0.955
+ $X2=2.835 $Y2=1.22
r49 15 16 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.805 $Y=0.805
+ $X2=2.805 $Y2=0.955
r50 10 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.535 $Y=2.18
+ $X2=2.745 $Y2=2.18
r51 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.745 $Y=2.105
+ $X2=2.745 $Y2=2.18
r52 9 18 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.745 $Y=2.105
+ $X2=2.745 $Y2=1.725
r53 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.685 $Y=0.485
+ $X2=2.685 $Y2=0.805
r54 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.535 $Y=2.255
+ $X2=2.535 $Y2=2.18
r55 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.535 $Y=2.255 $X2=2.535
+ $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_0%X 1 2 7 8 9 10 11 12 13 38 41
r19 41 42 2.93672 $w=4.83e-07 $l=2e-08 $layer=LI1_cond $X=0.327 $Y=2.405
+ $X2=0.327 $Y2=2.385
r20 22 33 2.04284 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=0.217 $Y=0.65
+ $X2=0.217 $Y2=0.485
r21 13 45 5.54882 $w=4.83e-07 $l=2.25e-07 $layer=LI1_cond $X=0.327 $Y=2.775
+ $X2=0.327 $Y2=2.55
r22 12 45 2.78674 $w=4.83e-07 $l=1.13e-07 $layer=LI1_cond $X=0.327 $Y=2.437
+ $X2=0.327 $Y2=2.55
r23 12 41 0.789165 $w=4.83e-07 $l=3.2e-08 $layer=LI1_cond $X=0.327 $Y=2.437
+ $X2=0.327 $Y2=2.405
r24 12 42 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=0.217 $Y=2.352
+ $X2=0.217 $Y2=2.385
r25 11 12 13.7858 $w=2.63e-07 $l=3.17e-07 $layer=LI1_cond $X=0.217 $Y=2.035
+ $X2=0.217 $Y2=2.352
r26 10 11 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.217 $Y=1.665
+ $X2=0.217 $Y2=2.035
r27 9 10 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.217 $Y=1.295
+ $X2=0.217 $Y2=1.665
r28 8 9 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.217 $Y=0.925
+ $X2=0.217 $Y2=1.295
r29 8 22 11.9593 $w=2.63e-07 $l=2.75e-07 $layer=LI1_cond $X=0.217 $Y=0.925
+ $X2=0.217 $Y2=0.65
r30 7 38 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.24 $Y=0.485
+ $X2=0.49 $Y2=0.485
r31 7 33 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=0.24 $Y=0.485
+ $X2=0.217 $Y2=0.485
r32 2 45 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.34
+ $Y=2.405 $X2=0.465 $Y2=2.55
r33 1 38 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.365
+ $Y=0.275 $X2=0.49 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_0%VPWR 1 2 9 13 16 17 18 24 30 31 34
r32 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.78 $Y2=3.33
r36 28 30 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=2.78 $Y2=3.33
r39 24 26 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 18 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 16 21 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.98 $Y2=3.33
r46 15 26 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.145 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=3.33
+ $X2=0.98 $Y2=3.33
r48 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=3.245
+ $X2=2.78 $Y2=3.33
r49 11 13 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.78 $Y=3.245
+ $X2=2.78 $Y2=2.55
r50 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.98 $Y=3.245 $X2=0.98
+ $Y2=3.33
r51 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.98 $Y=3.245
+ $X2=0.98 $Y2=2.55
r52 2 13 300 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=2 $X=2.61
+ $Y=2.405 $X2=2.78 $Y2=2.55
r53 1 9 300 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=2 $X=0.755
+ $Y=2.405 $X2=0.98 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_0%VGND 1 2 9 13 16 17 18 24 30 31 34
r40 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r41 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r42 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.02
+ $Y2=0
r44 28 30 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=3.12
+ $Y2=0
r45 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.02
+ $Y2=0
r46 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.68
+ $Y2=0
r47 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r49 18 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r50 18 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 16 21 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.72
+ $Y2=0
r52 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.99
+ $Y2=0
r53 15 26 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.68
+ $Y2=0
r54 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=0.99
+ $Y2=0
r55 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r56 11 13 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.44
r57 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=0.085 $X2=0.99
+ $Y2=0
r58 7 9 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.99 $Y=0.085 $X2=0.99
+ $Y2=0.485
r59 2 13 182 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.275 $X2=2.02 $Y2=0.44
r60 1 9 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=0.78
+ $Y=0.275 $X2=0.99 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_0%A_270_55# 1 2 7 11 14
r28 14 15 13.8237 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.525 $Y=0.485
+ $X2=1.525 $Y2=0.8
r29 9 11 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=2.48 $Y=0.715
+ $X2=2.48 $Y2=0.485
r30 8 15 3.61456 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.685 $Y=0.8 $X2=1.525
+ $Y2=0.8
r31 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.355 $Y=0.8
+ $X2=2.48 $Y2=0.715
r32 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.355 $Y=0.8 $X2=1.685
+ $Y2=0.8
r33 2 11 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.33
+ $Y=0.275 $X2=2.47 $Y2=0.485
r34 1 14 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1.35
+ $Y=0.275 $X2=1.53 $Y2=0.485
.ends

