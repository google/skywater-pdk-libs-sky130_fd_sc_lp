* File: sky130_fd_sc_lp__and4bb_4.spice
* Created: Fri Aug 28 10:09:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4bb_4.pex.spice"
.subckt sky130_fd_sc_lp__and4bb_4  VNB VPB B_N D C A_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A_N	A_N
* C	C
* D	D
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_B_N_M1001_g N_A_49_131#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=0.953333 PS=1.41 NRD=90 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75004.3 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_254_21#_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=1.90667 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1006_d N_A_254_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001 SB=75003.1
+ A=0.126 P=1.98 MULT=1
MM1013 N_X_M1013_d N_A_254_21#_M1013_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1015 N_X_M1013_d N_A_254_21#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2079 PD=1.12 PS=1.335 NRD=0 NRS=15 M=1 R=5.6 SA=75001.9
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1003 A_671_47# N_D_M1003_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.2079 PD=1.05 PS=1.335 NRD=7.14 NRS=15.708 M=1 R=5.6 SA=75002.5 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1005 A_743_47# N_C_M1005_g A_671_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75002.9 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1010 A_851_47# N_A_49_131#_M1010_g A_743_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=19.992 NRS=19.992 M=1 R=5.6 SA=75003.4
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1019 N_A_254_21#_M1019_d N_A_929_21#_M1019_g A_851_47# VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6
+ SA=75003.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1016 N_A_929_21#_M1016_d N_A_N_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_B_N_M1012_g N_A_49_131#_M1012_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1176 AS=0.1197 PD=0.925 PS=1.41 NRD=105.533 NRS=9.3772 M=1 R=2.8
+ SA=75000.2 SB=75004.8 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_254_21#_M1004_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3528 PD=1.54 PS=2.775 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1009 N_X_M1004_d N_A_254_21#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75003.3 A=0.189 P=2.82 MULT=1
MM1014 N_X_M1014_d N_A_254_21#_M1014_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.3
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1017 N_X_M1014_d N_A_254_21#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.26775 PD=1.54 PS=1.685 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75001.7
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1011 N_A_254_21#_M1011_d N_D_M1011_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.26775 PD=1.54 PS=1.685 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75002.3
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_A_254_21#_M1011_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.1764 PD=1.65 PS=1.54 NRD=9.3772 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1008 N_A_254_21#_M1008_d N_A_49_131#_M1008_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=8.5892 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_A_929_21#_M1018_g N_A_254_21#_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2898 AS=0.2457 PD=2.475 PS=1.65 NRD=0 NRS=8.5892 M=1 R=8.4
+ SA=75003.8 SB=75000.4 A=0.189 P=2.82 MULT=1
MM1002 N_A_929_21#_M1002_d N_A_N_M1002_g N_VPWR_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0966 PD=1.37 PS=0.825 NRD=0 NRS=82.0702 M=1 R=2.8
+ SA=75004.9 SB=75000.2 A=0.063 P=1.14 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3463 P=16.97
c_59 VNB 0 5.82218e-20 $X=0 $Y=0
c_107 VPB 0 1.63555e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__and4bb_4.pxi.spice"
*
.ends
*
*
