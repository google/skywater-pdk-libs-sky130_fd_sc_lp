* NGSPICE file created from sky130_fd_sc_lp__dlxtp_lp2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlxtp_lp2 D GATE VGND VNB VPB VPWR Q
M1000 a_880_47# a_240_409# a_778_47# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.512e+11p ps=1.56e+06u
M1001 a_928_21# a_778_47# a_1207_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1002 VGND D a_114_57# VNB nshort w=420000u l=150000u
+  ad=8.148e+11p pd=7.24e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_766_419# a_27_57# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=1.8553e+12p ps=1.181e+07u
M1004 VPWR D a_27_57# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1005 VGND a_928_21# a_880_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1477_83# a_928_21# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 Q a_928_21# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1008 Q a_928_21# a_1477_83# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1009 a_114_57# D a_27_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1010 VGND a_240_409# a_542_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1011 a_272_57# GATE VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1012 a_240_409# GATE a_272_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1013 VPWR a_240_409# a_452_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1014 a_240_409# GATE VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1015 a_778_47# a_240_409# a_766_419# VPB phighvt w=1e+06u l=250000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1016 VPWR a_928_21# a_972_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1017 a_542_47# a_240_409# a_452_419# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1018 a_700_47# a_27_57# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1019 a_972_419# a_452_419# a_778_47# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_928_21# a_778_47# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1021 a_778_47# a_452_419# a_700_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1207_47# a_778_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

