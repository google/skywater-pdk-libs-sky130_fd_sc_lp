* File: sky130_fd_sc_lp__o32a_m.spice
* Created: Fri Aug 28 11:17:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32a_m.pex.spice"
.subckt sky130_fd_sc_lp__o32a_m  VNB VPB A1 A2 A3 B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_86_55#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.10815 AS=0.1113 PD=0.935 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1009 N_A_249_81#_M1009_d N_A1_M1009_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.10815 PD=0.7 PS=0.935 NRD=0 NRS=61.428 M=1 R=2.8 SA=75000.9
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_249_81#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.105 AS=0.0588 PD=0.92 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_249_81#_M1004_d N_A3_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.105 PD=0.7 PS=0.92 NRD=0 NRS=57.132 M=1 R=2.8 SA=75001.9
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_A_86_55#_M1008_d N_B2_M1008_g N_A_249_81#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_249_81#_M1007_d N_B1_M1007_g N_A_86_55#_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1281 AS=0.0672 PD=1.45 PS=0.74 NRD=11.424 NRS=11.424 M=1 R=2.8
+ SA=75002.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_86_55#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.10815 AS=0.1113 PD=0.935 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1000 A_249_403# N_A1_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.10815 PD=0.63 PS=0.935 NRD=23.443 NRS=100.844 M=1 R=2.8
+ SA=75000.9 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1006 A_321_403# N_A2_M1006_g A_249_403# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=65.6601 NRS=23.443 M=1 R=2.8 SA=75001.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 N_A_86_55#_M1001_d N_A3_M1001_g A_321_403# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.11235 AS=0.0819 PD=0.955 PS=0.81 NRD=114.91 NRS=65.6601 M=1 R=2.8
+ SA=75001.8 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1010 A_566_403# N_B2_M1010_g N_A_86_55#_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.05145 AS=0.11235 PD=0.665 PS=0.955 NRD=31.6579 NRS=4.6886 M=1 R=2.8
+ SA=75002.4 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g A_566_403# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.05145 PD=1.41 PS=0.665 NRD=0 NRS=31.6579 M=1 R=2.8 SA=75002.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_42 VNB 0 2.96683e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o32a_m.pxi.spice"
*
.ends
*
*
