* File: sky130_fd_sc_lp__mux2i_2.pxi.spice
* Created: Fri Aug 28 10:45:08 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2I_2%S N_S_M1006_g N_S_M1012_g N_S_M1003_g N_S_M1004_g
+ N_S_M1010_g N_S_M1014_g N_S_c_135_p N_S_c_91_n N_S_c_100_n N_S_c_92_n
+ N_S_c_93_n S S S N_S_c_94_n N_S_c_95_n PM_SKY130_FD_SC_LP__MUX2I_2%S
x_PM_SKY130_FD_SC_LP__MUX2I_2%A_44_367# N_A_44_367#_M1012_s N_A_44_367#_M1006_s
+ N_A_44_367#_M1009_g N_A_44_367#_M1002_g N_A_44_367#_M1017_g
+ N_A_44_367#_M1015_g N_A_44_367#_c_193_n N_A_44_367#_c_194_n
+ N_A_44_367#_c_195_n N_A_44_367#_c_196_n N_A_44_367#_c_197_n
+ N_A_44_367#_c_226_n N_A_44_367#_c_198_n N_A_44_367#_c_199_n
+ PM_SKY130_FD_SC_LP__MUX2I_2%A_44_367#
x_PM_SKY130_FD_SC_LP__MUX2I_2%A0 N_A0_M1001_g N_A0_M1005_g N_A0_M1013_g
+ N_A0_M1011_g A0 A0 N_A0_c_270_n PM_SKY130_FD_SC_LP__MUX2I_2%A0
x_PM_SKY130_FD_SC_LP__MUX2I_2%A1 N_A1_M1000_g N_A1_M1007_g N_A1_c_328_n
+ N_A1_M1016_g N_A1_M1008_g N_A1_c_330_n A1 A1 N_A1_c_332_n
+ PM_SKY130_FD_SC_LP__MUX2I_2%A1
x_PM_SKY130_FD_SC_LP__MUX2I_2%VPWR N_VPWR_M1006_d N_VPWR_M1015_s N_VPWR_M1014_s
+ N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n VPWR N_VPWR_c_379_n
+ N_VPWR_c_380_n N_VPWR_c_375_n N_VPWR_c_382_n N_VPWR_c_383_n
+ PM_SKY130_FD_SC_LP__MUX2I_2%VPWR
x_PM_SKY130_FD_SC_LP__MUX2I_2%A_251_367# N_A_251_367#_M1002_d
+ N_A_251_367#_M1000_s N_A_251_367#_c_445_n N_A_251_367#_c_458_n
+ N_A_251_367#_c_492_p N_A_251_367#_c_452_n N_A_251_367#_c_446_n
+ PM_SKY130_FD_SC_LP__MUX2I_2%A_251_367#
x_PM_SKY130_FD_SC_LP__MUX2I_2%A_455_367# N_A_455_367#_M1004_d
+ N_A_455_367#_M1005_s N_A_455_367#_c_495_n N_A_455_367#_c_494_n
+ N_A_455_367#_c_501_n N_A_455_367#_c_506_n
+ PM_SKY130_FD_SC_LP__MUX2I_2%A_455_367#
x_PM_SKY130_FD_SC_LP__MUX2I_2%Y N_Y_M1001_d N_Y_M1013_d N_Y_M1008_s N_Y_M1005_d
+ N_Y_M1011_d N_Y_M1016_d N_Y_c_524_n N_Y_c_541_n N_Y_c_560_n N_Y_c_545_n
+ N_Y_c_525_n N_Y_c_531_n N_Y_c_532_n N_Y_c_526_n N_Y_c_527_n N_Y_c_548_n
+ N_Y_c_528_n Y Y N_Y_c_530_n PM_SKY130_FD_SC_LP__MUX2I_2%Y
x_PM_SKY130_FD_SC_LP__MUX2I_2%VGND N_VGND_M1012_d N_VGND_M1017_d N_VGND_M1010_d
+ N_VGND_c_612_n N_VGND_c_613_n N_VGND_c_658_p N_VGND_c_614_n N_VGND_c_615_n
+ N_VGND_c_616_n N_VGND_c_617_n N_VGND_c_618_n VGND N_VGND_c_619_n
+ N_VGND_c_620_n PM_SKY130_FD_SC_LP__MUX2I_2%VGND
x_PM_SKY130_FD_SC_LP__MUX2I_2%A_251_47# N_A_251_47#_M1009_s N_A_251_47#_M1001_s
+ N_A_251_47#_c_703_n N_A_251_47#_c_671_n N_A_251_47#_c_672_n
+ N_A_251_47#_c_673_n N_A_251_47#_c_674_n N_A_251_47#_c_675_n
+ PM_SKY130_FD_SC_LP__MUX2I_2%A_251_47#
x_PM_SKY130_FD_SC_LP__MUX2I_2%A_423_47# N_A_423_47#_M1003_s N_A_423_47#_M1007_d
+ N_A_423_47#_c_716_n N_A_423_47#_c_724_n N_A_423_47#_c_718_n
+ PM_SKY130_FD_SC_LP__MUX2I_2%A_423_47#
cc_1 VNB N_S_M1012_g 0.0286203f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.655
cc_2 VNB N_S_M1003_g 0.0232219f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=0.655
cc_3 VNB N_S_M1010_g 0.0313016f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=0.655
cc_4 VNB N_S_M1014_g 0.00958183f $X=-0.19 $Y=-0.245 $X2=2.63 $Y2=2.465
cc_5 VNB N_S_c_91_n 6.24257e-19 $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.51
cc_6 VNB N_S_c_92_n 0.00155076f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.537
cc_7 VNB N_S_c_93_n 0.00268534f $X=-0.19 $Y=-0.245 $X2=2.11 $Y2=1.51
cc_8 VNB N_S_c_94_n 0.0311865f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.51
cc_9 VNB N_S_c_95_n 0.0396985f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=1.495
cc_10 VNB N_A_44_367#_M1009_g 0.0224994f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.345
cc_11 VNB N_A_44_367#_M1017_g 0.022689f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=1.345
cc_12 VNB N_A_44_367#_c_193_n 0.0360614f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.855
cc_13 VNB N_A_44_367#_c_194_n 0.0260191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_44_367#_c_195_n 0.00401721f $X=-0.19 $Y=-0.245 $X2=2.11 $Y2=1.537
cc_15 VNB N_A_44_367#_c_196_n 0.00186456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_44_367#_c_197_n 0.00261724f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_17 VNB N_A_44_367#_c_198_n 0.0120286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_44_367#_c_199_n 0.030739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A0_M1001_g 0.0225015f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.465
cc_20 VNB N_A0_M1013_g 0.0192661f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=0.655
cc_21 VNB A0 0.00366321f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=0.655
cc_22 VNB N_A0_c_270_n 0.0349039f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.51
cc_23 VNB N_A1_M1000_g 0.00663107f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.465
cc_24 VNB N_A1_M1007_g 0.020166f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.655
cc_25 VNB N_A1_c_328_n 0.0100574f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.345
cc_26 VNB N_A1_M1008_g 0.0265473f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=1.345
cc_27 VNB N_A1_c_330_n 0.0106818f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=0.655
cc_28 VNB A1 0.0179127f $X=-0.19 $Y=-0.245 $X2=2.63 $Y2=1.495
cc_29 VNB N_A1_c_332_n 0.0261046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_375_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_524_n 0.00336286f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=0.655
cc_32 VNB N_Y_c_525_n 0.0136102f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.855
cc_33 VNB N_Y_c_526_n 0.0303392f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.95
cc_34 VNB N_Y_c_527_n 0.0035578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_528_n 0.00262892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB Y 0.00988135f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.495
cc_37 VNB N_Y_c_530_n 0.0142643f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.987
cc_38 VNB N_VGND_c_612_n 4.06069e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_613_n 0.0043071f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=1.345
cc_40 VNB N_VGND_c_614_n 0.00311372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_615_n 0.0223395f $X=-0.19 $Y=-0.245 $X2=2.63 $Y2=2.465
cc_42 VNB N_VGND_c_616_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_617_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.51
cc_44 VNB N_VGND_c_618_n 0.00422832f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.51
cc_45 VNB N_VGND_c_619_n 0.091919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_620_n 0.314394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_251_47#_c_671_n 0.0241185f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=0.655
cc_48 VNB N_A_251_47#_c_672_n 0.00368988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_251_47#_c_673_n 0.00756793f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=2.465
cc_50 VNB N_A_251_47#_c_674_n 0.00482789f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=2.465
cc_51 VNB N_A_251_47#_c_675_n 0.00892567f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=1.345
cc_52 VNB N_A_423_47#_c_716_n 0.0243027f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.655
cc_53 VPB N_S_M1006_g 0.0231726f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.465
cc_54 VPB N_S_M1004_g 0.0205855f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=2.465
cc_55 VPB N_S_M1014_g 0.0233172f $X=-0.19 $Y=1.655 $X2=2.63 $Y2=2.465
cc_56 VPB N_S_c_91_n 0.00174179f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.51
cc_57 VPB N_S_c_100_n 0.0016686f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.855
cc_58 VPB N_S_c_93_n 0.00355511f $X=-0.19 $Y=1.655 $X2=2.11 $Y2=1.51
cc_59 VPB N_S_c_94_n 0.00779678f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.51
cc_60 VPB N_S_c_95_n 0.0110729f $X=-0.19 $Y=1.655 $X2=2.47 $Y2=1.495
cc_61 VPB N_A_44_367#_M1002_g 0.0212836f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=1.675
cc_62 VPB N_A_44_367#_M1015_g 0.0200478f $X=-0.19 $Y=1.655 $X2=2.63 $Y2=1.495
cc_63 VPB N_A_44_367#_c_194_n 0.0561703f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_44_367#_c_199_n 0.00336956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A0_M1005_g 0.0231192f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.655
cc_66 VPB N_A0_M1011_g 0.0183361f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=2.465
cc_67 VPB A0 0.00553878f $X=-0.19 $Y=1.655 $X2=2.47 $Y2=0.655
cc_68 VPB N_A0_c_270_n 0.0048949f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.51
cc_69 VPB N_A1_M1000_g 0.0192191f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.465
cc_70 VPB N_A1_M1016_g 0.0244533f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=1.675
cc_71 VPB A1 0.0177145f $X=-0.19 $Y=1.655 $X2=2.63 $Y2=1.495
cc_72 VPB N_A1_c_332_n 0.00665874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_376_n 0.00564356f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=2.465
cc_74 VPB N_VPWR_c_377_n 0.0109593f $X=-0.19 $Y=1.655 $X2=2.47 $Y2=1.345
cc_75 VPB N_VPWR_c_378_n 0.0187902f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_379_n 0.019333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_380_n 0.0663362f $X=-0.19 $Y=1.655 $X2=2.11 $Y2=1.51
cc_78 VPB N_VPWR_c_375_n 0.0612326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_382_n 0.0286313f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.95
cc_80 VPB N_VPWR_c_383_n 0.0125639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_251_367#_c_445_n 0.00568868f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.655
cc_82 VPB N_A_251_367#_c_446_n 0.00771723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A_455_367#_c_494_n 0.00773363f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=0.655
cc_84 VPB N_Y_c_531_n 0.00797287f $X=-0.19 $Y=1.655 $X2=2.11 $Y2=1.537
cc_85 VPB N_Y_c_532_n 0.0374933f $X=-0.19 $Y=1.655 $X2=2.11 $Y2=1.51
cc_86 VPB N_Y_c_530_n 0.0121441f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.987
cc_87 N_S_M1012_g N_A_44_367#_M1009_g 0.0236346f $X=0.75 $Y=0.655 $X2=0 $Y2=0
cc_88 N_S_M1006_g N_A_44_367#_M1002_g 0.0303514f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_89 N_S_c_91_n N_A_44_367#_M1002_g 0.00341483f $X=0.695 $Y=1.51 $X2=0 $Y2=0
cc_90 N_S_c_100_n N_A_44_367#_M1002_g 8.72188e-19 $X=1.765 $Y=1.855 $X2=0 $Y2=0
cc_91 S N_A_44_367#_M1002_g 0.0201256f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_92 N_S_M1003_g N_A_44_367#_M1017_g 0.0266864f $X=2.04 $Y=0.655 $X2=0 $Y2=0
cc_93 N_S_M1004_g N_A_44_367#_M1015_g 0.0384112f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_94 N_S_c_100_n N_A_44_367#_M1015_g 0.00798118f $X=1.765 $Y=1.855 $X2=0 $Y2=0
cc_95 S N_A_44_367#_M1015_g 0.0140634f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_96 N_S_M1012_g N_A_44_367#_c_194_n 0.00405742f $X=0.75 $Y=0.655 $X2=0 $Y2=0
cc_97 N_S_c_91_n N_A_44_367#_c_194_n 0.0369921f $X=0.695 $Y=1.51 $X2=0 $Y2=0
cc_98 N_S_c_94_n N_A_44_367#_c_194_n 0.015392f $X=0.75 $Y=1.51 $X2=0 $Y2=0
cc_99 N_S_M1012_g N_A_44_367#_c_195_n 0.0150916f $X=0.75 $Y=0.655 $X2=0 $Y2=0
cc_100 N_S_c_91_n N_A_44_367#_c_195_n 0.0112095f $X=0.695 $Y=1.51 $X2=0 $Y2=0
cc_101 N_S_c_94_n N_A_44_367#_c_195_n 0.00159369f $X=0.75 $Y=1.51 $X2=0 $Y2=0
cc_102 N_S_M1012_g N_A_44_367#_c_196_n 0.00185499f $X=0.75 $Y=0.655 $X2=0 $Y2=0
cc_103 N_S_c_91_n N_A_44_367#_c_196_n 0.00498957f $X=0.695 $Y=1.51 $X2=0 $Y2=0
cc_104 N_S_c_92_n N_A_44_367#_c_196_n 2.73765e-19 $X=1.85 $Y=1.537 $X2=0 $Y2=0
cc_105 N_S_c_94_n N_A_44_367#_c_196_n 4.68395e-19 $X=0.75 $Y=1.51 $X2=0 $Y2=0
cc_106 N_S_c_91_n N_A_44_367#_c_197_n 0.0133546f $X=0.695 $Y=1.51 $X2=0 $Y2=0
cc_107 S N_A_44_367#_c_197_n 0.00855441f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_108 N_S_c_94_n N_A_44_367#_c_197_n 0.00125897f $X=0.75 $Y=1.51 $X2=0 $Y2=0
cc_109 N_S_c_92_n N_A_44_367#_c_226_n 0.010201f $X=1.85 $Y=1.537 $X2=0 $Y2=0
cc_110 S N_A_44_367#_c_226_n 0.0136484f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_111 N_S_c_91_n N_A_44_367#_c_198_n 0.00155683f $X=0.695 $Y=1.51 $X2=0 $Y2=0
cc_112 N_S_c_94_n N_A_44_367#_c_198_n 0.006113f $X=0.75 $Y=1.51 $X2=0 $Y2=0
cc_113 N_S_c_91_n N_A_44_367#_c_199_n 7.76658e-19 $X=0.695 $Y=1.51 $X2=0 $Y2=0
cc_114 N_S_c_92_n N_A_44_367#_c_199_n 0.0101796f $X=1.85 $Y=1.537 $X2=0 $Y2=0
cc_115 S N_A_44_367#_c_199_n 0.00237122f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_116 N_S_c_94_n N_A_44_367#_c_199_n 0.0177754f $X=0.75 $Y=1.51 $X2=0 $Y2=0
cc_117 N_S_c_95_n N_A_44_367#_c_199_n 0.0175458f $X=2.47 $Y=1.495 $X2=0 $Y2=0
cc_118 N_S_c_135_p N_VPWR_M1006_d 0.00172027f $X=0.7 $Y=1.855 $X2=-0.19
+ $Y2=-0.245
cc_119 N_S_c_91_n N_VPWR_M1006_d 2.4934e-19 $X=0.695 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_120 S N_VPWR_M1006_d 0.0106825f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_121 N_S_c_100_n N_VPWR_M1015_s 0.00568046f $X=1.765 $Y=1.855 $X2=0 $Y2=0
cc_122 N_S_M1006_g N_VPWR_c_376_n 0.0121008f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_123 N_S_c_135_p N_VPWR_c_376_n 0.0070777f $X=0.7 $Y=1.855 $X2=0 $Y2=0
cc_124 S N_VPWR_c_376_n 0.0208436f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_125 N_S_c_94_n N_VPWR_c_376_n 3.62324e-19 $X=0.75 $Y=1.51 $X2=0 $Y2=0
cc_126 N_S_M1004_g N_VPWR_c_377_n 0.00408156f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_127 N_S_M1004_g N_VPWR_c_379_n 0.00413624f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_128 N_S_M1014_g N_VPWR_c_379_n 0.00413624f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_129 N_S_M1006_g N_VPWR_c_375_n 0.0122586f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_130 N_S_M1004_g N_VPWR_c_375_n 0.00611928f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_131 N_S_M1014_g N_VPWR_c_375_n 0.00722417f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_132 N_S_M1006_g N_VPWR_c_382_n 0.00585385f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_133 N_S_M1014_g N_VPWR_c_383_n 0.0104248f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_134 S N_A_251_367#_M1002_d 0.00398049f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_135 N_S_M1004_g N_A_251_367#_c_445_n 0.0160649f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_136 N_S_M1014_g N_A_251_367#_c_445_n 0.0134215f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_137 N_S_c_100_n N_A_251_367#_c_445_n 0.00422673f $X=1.765 $Y=1.855 $X2=0
+ $Y2=0
cc_138 S N_A_251_367#_c_445_n 0.00360474f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_139 N_S_M1004_g N_A_251_367#_c_452_n 0.00225973f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_140 S N_A_251_367#_c_452_n 0.0176092f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_141 N_S_M1014_g N_A_251_367#_c_446_n 0.00422161f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_142 N_S_M1004_g N_A_455_367#_c_495_n 0.00757486f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_143 N_S_M1014_g N_A_455_367#_c_495_n 0.0113577f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_144 N_S_c_100_n N_A_455_367#_c_495_n 0.0118692f $X=1.765 $Y=1.855 $X2=0 $Y2=0
cc_145 N_S_c_93_n N_A_455_367#_c_495_n 0.00182306f $X=2.11 $Y=1.51 $X2=0 $Y2=0
cc_146 N_S_c_95_n N_A_455_367#_c_495_n 0.00265022f $X=2.47 $Y=1.495 $X2=0 $Y2=0
cc_147 N_S_M1014_g N_A_455_367#_c_494_n 0.0131906f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_148 N_S_M1004_g N_A_455_367#_c_501_n 0.00413475f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_149 N_S_M1014_g N_A_455_367#_c_501_n 7.15561e-19 $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_150 N_S_c_95_n Y 0.00582038f $X=2.47 $Y=1.495 $X2=0 $Y2=0
cc_151 N_S_M1014_g N_Y_c_530_n 0.0148481f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_152 N_S_c_93_n N_Y_c_530_n 0.00297993f $X=2.11 $Y=1.51 $X2=0 $Y2=0
cc_153 N_S_M1012_g N_VGND_c_612_n 0.0116893f $X=0.75 $Y=0.655 $X2=0 $Y2=0
cc_154 N_S_M1003_g N_VGND_c_613_n 0.00284552f $X=2.04 $Y=0.655 $X2=0 $Y2=0
cc_155 N_S_M1003_g N_VGND_c_614_n 0.0110436f $X=2.04 $Y=0.655 $X2=0 $Y2=0
cc_156 N_S_M1010_g N_VGND_c_614_n 0.0100435f $X=2.47 $Y=0.655 $X2=0 $Y2=0
cc_157 N_S_M1012_g N_VGND_c_615_n 0.00486043f $X=0.75 $Y=0.655 $X2=0 $Y2=0
cc_158 N_S_M1003_g N_VGND_c_619_n 0.00418726f $X=2.04 $Y=0.655 $X2=0 $Y2=0
cc_159 N_S_M1010_g N_VGND_c_619_n 0.00357877f $X=2.47 $Y=0.655 $X2=0 $Y2=0
cc_160 N_S_M1012_g N_VGND_c_620_n 0.00935659f $X=0.75 $Y=0.655 $X2=0 $Y2=0
cc_161 N_S_M1003_g N_VGND_c_620_n 0.00573747f $X=2.04 $Y=0.655 $X2=0 $Y2=0
cc_162 N_S_M1010_g N_VGND_c_620_n 0.00675087f $X=2.47 $Y=0.655 $X2=0 $Y2=0
cc_163 N_S_M1003_g N_A_251_47#_c_671_n 0.010446f $X=2.04 $Y=0.655 $X2=0 $Y2=0
cc_164 N_S_M1010_g N_A_251_47#_c_671_n 0.0141073f $X=2.47 $Y=0.655 $X2=0 $Y2=0
cc_165 N_S_c_92_n N_A_251_47#_c_671_n 0.0143768f $X=1.85 $Y=1.537 $X2=0 $Y2=0
cc_166 N_S_c_93_n N_A_251_47#_c_671_n 0.0311944f $X=2.11 $Y=1.51 $X2=0 $Y2=0
cc_167 S N_A_251_47#_c_671_n 0.00352718f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_168 N_S_c_95_n N_A_251_47#_c_671_n 0.0101635f $X=2.47 $Y=1.495 $X2=0 $Y2=0
cc_169 S N_A_251_47#_c_672_n 0.00242518f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_170 N_S_M1010_g N_A_251_47#_c_673_n 0.00329846f $X=2.47 $Y=0.655 $X2=0 $Y2=0
cc_171 N_S_M1010_g N_A_423_47#_c_716_n 0.00947844f $X=2.47 $Y=0.655 $X2=0 $Y2=0
cc_172 N_S_M1003_g N_A_423_47#_c_718_n 0.00305805f $X=2.04 $Y=0.655 $X2=0 $Y2=0
cc_173 N_S_M1010_g N_A_423_47#_c_718_n 0.00394338f $X=2.47 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A_44_367#_M1002_g N_VPWR_c_376_n 0.0133354f $X=1.18 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A_44_367#_M1015_g N_VPWR_c_377_n 0.00408156f $X=1.61 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_44_367#_M1002_g N_VPWR_c_378_n 0.0055231f $X=1.18 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_44_367#_M1015_g N_VPWR_c_378_n 0.00409176f $X=1.61 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_44_367#_M1006_s N_VPWR_c_375_n 0.00371702f $X=0.22 $Y=1.835 $X2=0
+ $Y2=0
cc_179 N_A_44_367#_M1002_g N_VPWR_c_375_n 0.0104566f $X=1.18 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_44_367#_M1015_g N_VPWR_c_375_n 0.00604968f $X=1.61 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_44_367#_c_194_n N_VPWR_c_375_n 0.0100304f $X=0.345 $Y=1.98 $X2=0
+ $Y2=0
cc_182 N_A_44_367#_c_194_n N_VPWR_c_382_n 0.0178111f $X=0.345 $Y=1.98 $X2=0
+ $Y2=0
cc_183 N_A_44_367#_M1015_g N_A_251_367#_c_445_n 0.0112821f $X=1.61 $Y=2.465
+ $X2=0 $Y2=0
cc_184 N_A_44_367#_M1002_g N_A_251_367#_c_452_n 0.00946194f $X=1.18 $Y=2.465
+ $X2=0 $Y2=0
cc_185 N_A_44_367#_M1015_g N_A_251_367#_c_452_n 0.0132368f $X=1.61 $Y=2.465
+ $X2=0 $Y2=0
cc_186 N_A_44_367#_M1015_g N_A_455_367#_c_495_n 8.77182e-19 $X=1.61 $Y=2.465
+ $X2=0 $Y2=0
cc_187 N_A_44_367#_M1015_g N_A_455_367#_c_501_n 7.62044e-19 $X=1.61 $Y=2.465
+ $X2=0 $Y2=0
cc_188 N_A_44_367#_c_195_n N_VGND_M1012_d 0.00178864f $X=0.96 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_189 N_A_44_367#_M1009_g N_VGND_c_612_n 0.01003f $X=1.18 $Y=0.655 $X2=0 $Y2=0
cc_190 N_A_44_367#_M1017_g N_VGND_c_612_n 6.24575e-19 $X=1.61 $Y=0.655 $X2=0
+ $Y2=0
cc_191 N_A_44_367#_c_195_n N_VGND_c_612_n 0.017927f $X=0.96 $Y=1.07 $X2=0 $Y2=0
cc_192 N_A_44_367#_M1017_g N_VGND_c_613_n 0.00155004f $X=1.61 $Y=0.655 $X2=0
+ $Y2=0
cc_193 N_A_44_367#_c_193_n N_VGND_c_615_n 0.0314316f $X=0.535 $Y=0.42 $X2=0
+ $Y2=0
cc_194 N_A_44_367#_M1009_g N_VGND_c_617_n 0.00486043f $X=1.18 $Y=0.655 $X2=0
+ $Y2=0
cc_195 N_A_44_367#_M1017_g N_VGND_c_617_n 0.00585385f $X=1.61 $Y=0.655 $X2=0
+ $Y2=0
cc_196 N_A_44_367#_M1012_s N_VGND_c_620_n 0.00371702f $X=0.41 $Y=0.235 $X2=0
+ $Y2=0
cc_197 N_A_44_367#_M1009_g N_VGND_c_620_n 0.00824727f $X=1.18 $Y=0.655 $X2=0
+ $Y2=0
cc_198 N_A_44_367#_M1017_g N_VGND_c_620_n 0.0105614f $X=1.61 $Y=0.655 $X2=0
+ $Y2=0
cc_199 N_A_44_367#_c_193_n N_VGND_c_620_n 0.0174172f $X=0.535 $Y=0.42 $X2=0
+ $Y2=0
cc_200 N_A_44_367#_M1017_g N_A_251_47#_c_671_n 0.0164802f $X=1.61 $Y=0.655 $X2=0
+ $Y2=0
cc_201 N_A_44_367#_M1009_g N_A_251_47#_c_672_n 0.00131418f $X=1.18 $Y=0.655
+ $X2=0 $Y2=0
cc_202 N_A_44_367#_c_195_n N_A_251_47#_c_672_n 0.00750776f $X=0.96 $Y=1.07 $X2=0
+ $Y2=0
cc_203 N_A_44_367#_c_196_n N_A_251_47#_c_672_n 0.00641961f $X=1.045 $Y=1.415
+ $X2=0 $Y2=0
cc_204 N_A_44_367#_c_226_n N_A_251_47#_c_672_n 0.0104349f $X=1.27 $Y=1.5 $X2=0
+ $Y2=0
cc_205 N_A_44_367#_c_199_n N_A_251_47#_c_672_n 0.00262478f $X=1.61 $Y=1.5 $X2=0
+ $Y2=0
cc_206 N_A0_M1011_g N_A1_M1000_g 0.0264218f $X=4.19 $Y=2.465 $X2=0 $Y2=0
cc_207 A0 N_A1_M1000_g 0.00944728f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_208 N_A0_M1013_g N_A1_M1007_g 0.0250763f $X=4.19 $Y=0.765 $X2=0 $Y2=0
cc_209 A0 N_A1_M1016_g 2.39336e-19 $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_210 A0 N_A1_c_330_n 0.00521878f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_211 N_A0_c_270_n N_A1_c_330_n 0.0264218f $X=4.19 $Y=1.51 $X2=0 $Y2=0
cc_212 A0 A1 0.0296328f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_213 A0 N_A1_c_332_n 5.99532e-19 $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_214 N_A0_M1005_g N_VPWR_c_380_n 0.00357877f $X=3.76 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A0_M1011_g N_VPWR_c_380_n 0.00357877f $X=4.19 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A0_M1005_g N_VPWR_c_375_n 0.0068216f $X=3.76 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A0_M1011_g N_VPWR_c_375_n 0.00544922f $X=4.19 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A0_M1005_g N_VPWR_c_383_n 0.00225041f $X=3.76 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A0_M1005_g N_A_251_367#_c_458_n 0.0121293f $X=3.76 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A0_M1011_g N_A_251_367#_c_458_n 0.0134852f $X=4.19 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A0_M1005_g N_A_251_367#_c_446_n 0.00903418f $X=3.76 $Y=2.465 $X2=0
+ $Y2=0
cc_222 N_A0_M1005_g N_A_455_367#_c_494_n 0.0124953f $X=3.76 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A0_M1005_g N_A_455_367#_c_506_n 0.00945723f $X=3.76 $Y=2.465 $X2=0
+ $Y2=0
cc_224 N_A0_M1001_g N_Y_c_524_n 0.0118409f $X=3.76 $Y=0.765 $X2=0 $Y2=0
cc_225 N_A0_M1013_g N_Y_c_524_n 0.0169781f $X=4.19 $Y=0.765 $X2=0 $Y2=0
cc_226 A0 N_Y_c_524_n 0.0283626f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_227 N_A0_c_270_n N_Y_c_524_n 0.00254295f $X=4.19 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A0_M1005_g N_Y_c_541_n 0.00920433f $X=3.76 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A0_M1011_g N_Y_c_541_n 0.01115f $X=4.19 $Y=2.465 $X2=0 $Y2=0
cc_230 A0 N_Y_c_541_n 0.0208256f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_231 N_A0_c_270_n N_Y_c_541_n 7.6966e-19 $X=4.19 $Y=1.51 $X2=0 $Y2=0
cc_232 A0 N_Y_c_545_n 0.00974964f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_233 A0 N_Y_c_525_n 0.00439604f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_234 N_A0_M1001_g N_Y_c_527_n 0.0021624f $X=3.76 $Y=0.765 $X2=0 $Y2=0
cc_235 N_A0_M1005_g N_Y_c_548_n 9.63823e-19 $X=3.76 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A0_M1011_g N_Y_c_548_n 0.0107071f $X=4.19 $Y=2.465 $X2=0 $Y2=0
cc_237 A0 N_Y_c_548_n 0.0230325f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_238 A0 N_Y_c_528_n 0.0273184f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_239 N_A0_M1001_g Y 0.00377805f $X=3.76 $Y=0.765 $X2=0 $Y2=0
cc_240 N_A0_M1013_g Y 4.80034e-19 $X=4.19 $Y=0.765 $X2=0 $Y2=0
cc_241 A0 Y 0.00981379f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_242 N_A0_c_270_n Y 0.0115381f $X=4.19 $Y=1.51 $X2=0 $Y2=0
cc_243 N_A0_M1005_g N_Y_c_530_n 0.00876026f $X=3.76 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A0_M1011_g N_Y_c_530_n 8.85693e-19 $X=4.19 $Y=2.465 $X2=0 $Y2=0
cc_245 A0 N_Y_c_530_n 0.0116489f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A0_c_270_n N_Y_c_530_n 0.00422415f $X=4.19 $Y=1.51 $X2=0 $Y2=0
cc_247 N_A0_M1001_g N_VGND_c_619_n 0.0029147f $X=3.76 $Y=0.765 $X2=0 $Y2=0
cc_248 N_A0_M1013_g N_VGND_c_619_n 0.0029147f $X=4.19 $Y=0.765 $X2=0 $Y2=0
cc_249 N_A0_M1001_g N_VGND_c_620_n 0.00428625f $X=3.76 $Y=0.765 $X2=0 $Y2=0
cc_250 N_A0_M1013_g N_VGND_c_620_n 0.0040339f $X=4.19 $Y=0.765 $X2=0 $Y2=0
cc_251 N_A0_M1001_g N_A_251_47#_c_671_n 4.14017e-19 $X=3.76 $Y=0.765 $X2=0 $Y2=0
cc_252 N_A0_M1001_g N_A_251_47#_c_673_n 0.0030403f $X=3.76 $Y=0.765 $X2=0 $Y2=0
cc_253 N_A0_M1001_g N_A_251_47#_c_675_n 0.0111493f $X=3.76 $Y=0.765 $X2=0 $Y2=0
cc_254 N_A0_M1013_g N_A_251_47#_c_675_n 0.00263201f $X=4.19 $Y=0.765 $X2=0 $Y2=0
cc_255 N_A0_M1001_g N_A_423_47#_c_716_n 0.0118489f $X=3.76 $Y=0.765 $X2=0 $Y2=0
cc_256 N_A0_M1013_g N_A_423_47#_c_716_n 0.0115786f $X=4.19 $Y=0.765 $X2=0 $Y2=0
cc_257 N_A1_M1000_g N_VPWR_c_380_n 0.00357877f $X=4.62 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A1_M1016_g N_VPWR_c_380_n 0.00585385f $X=5.05 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A1_M1000_g N_VPWR_c_375_n 0.00537849f $X=4.62 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A1_M1016_g N_VPWR_c_375_n 0.0118571f $X=5.05 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A1_M1000_g N_A_251_367#_c_458_n 0.0114565f $X=4.62 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A1_M1007_g N_Y_c_560_n 0.00461595f $X=4.7 $Y=0.765 $X2=0 $Y2=0
cc_263 N_A1_M1000_g N_Y_c_545_n 0.0114269f $X=4.62 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A1_c_328_n N_Y_c_545_n 2.29319e-19 $X=4.955 $Y=1.42 $X2=0 $Y2=0
cc_265 N_A1_M1016_g N_Y_c_545_n 0.0133021f $X=5.05 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A1_c_330_n N_Y_c_545_n 0.00362828f $X=4.66 $Y=1.42 $X2=0 $Y2=0
cc_267 A1 N_Y_c_545_n 0.0160721f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_268 N_A1_M1007_g N_Y_c_525_n 0.0101809f $X=4.7 $Y=0.765 $X2=0 $Y2=0
cc_269 N_A1_c_328_n N_Y_c_525_n 0.00447387f $X=4.955 $Y=1.42 $X2=0 $Y2=0
cc_270 N_A1_M1008_g N_Y_c_525_n 0.0139555f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_271 A1 N_Y_c_525_n 0.0536089f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_272 A1 N_Y_c_531_n 0.0235066f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_273 N_A1_c_332_n N_Y_c_531_n 8.44519e-19 $X=5.12 $Y=1.42 $X2=0 $Y2=0
cc_274 N_A1_M1008_g N_Y_c_526_n 0.00333601f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_275 N_A1_M1000_g N_Y_c_548_n 0.0105899f $X=4.62 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A1_M1016_g N_Y_c_548_n 5.73632e-19 $X=5.05 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A1_M1007_g N_Y_c_528_n 0.00390216f $X=4.7 $Y=0.765 $X2=0 $Y2=0
cc_278 N_A1_M1008_g N_Y_c_528_n 3.94875e-19 $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_279 N_A1_c_330_n N_Y_c_528_n 0.00237679f $X=4.66 $Y=1.42 $X2=0 $Y2=0
cc_280 N_A1_M1007_g N_VGND_c_619_n 0.0029147f $X=4.7 $Y=0.765 $X2=0 $Y2=0
cc_281 N_A1_M1008_g N_VGND_c_619_n 0.00450424f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_282 N_A1_M1007_g N_VGND_c_620_n 0.00407861f $X=4.7 $Y=0.765 $X2=0 $Y2=0
cc_283 N_A1_M1008_g N_VGND_c_620_n 0.00889332f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_284 N_A1_M1007_g N_A_423_47#_c_716_n 0.0123674f $X=4.7 $Y=0.765 $X2=0 $Y2=0
cc_285 N_A1_M1008_g N_A_423_47#_c_716_n 0.00609688f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_286 N_A1_M1008_g N_A_423_47#_c_724_n 0.00532885f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_287 N_VPWR_c_375_n N_A_251_367#_M1002_d 0.00236284f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_288 N_VPWR_c_375_n N_A_251_367#_M1000_s 0.00254871f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_289 N_VPWR_M1015_s N_A_251_367#_c_445_n 0.0142273f $X=1.685 $Y=1.835 $X2=0
+ $Y2=0
cc_290 N_VPWR_M1014_s N_A_251_367#_c_445_n 0.00932999f $X=2.705 $Y=1.835 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_377_n N_A_251_367#_c_445_n 0.0242216f $X=1.905 $Y=3.045 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_378_n N_A_251_367#_c_445_n 0.00310672f $X=1.74 $Y=3.33 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_379_n N_A_251_367#_c_445_n 0.0127155f $X=2.795 $Y=3.33 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_380_n N_A_251_367#_c_445_n 0.00388164f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_375_n N_A_251_367#_c_445_n 0.0342103f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_383_n N_A_251_367#_c_445_n 0.0244235f $X=2.96 $Y=3.045 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_380_n N_A_251_367#_c_458_n 0.083799f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_298 N_VPWR_c_375_n N_A_251_367#_c_458_n 0.0541863f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_376_n N_A_251_367#_c_452_n 0.0484479f $X=0.875 $Y=2.375 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_378_n N_A_251_367#_c_452_n 0.0113252f $X=1.74 $Y=3.33 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_375_n N_A_251_367#_c_452_n 0.0117838f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_380_n N_A_251_367#_c_446_n 0.0116549f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_375_n N_A_251_367#_c_446_n 0.00647164f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_383_n N_A_251_367#_c_446_n 0.0102808f $X=2.96 $Y=3.045 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_375_n N_A_455_367#_M1004_d 0.00296296f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_306 N_VPWR_c_375_n N_A_455_367#_M1005_s 0.00225186f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_307 N_VPWR_M1014_s N_A_455_367#_c_494_n 0.0123258f $X=2.705 $Y=1.835 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_375_n N_Y_M1005_d 0.00215172f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_c_375_n N_Y_M1011_d 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_310 N_VPWR_c_375_n N_Y_M1016_d 0.00249946f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_311 N_VPWR_c_380_n N_Y_c_532_n 0.0190529f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_312 N_VPWR_c_375_n N_Y_c_532_n 0.0113912f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_313 N_VPWR_M1014_s N_Y_c_530_n 0.00865036f $X=2.705 $Y=1.835 $X2=0 $Y2=0
cc_314 N_A_251_367#_c_445_n N_A_455_367#_M1004_d 0.0043979f $X=3.305 $Y=2.685
+ $X2=-0.19 $Y2=1.655
cc_315 N_A_251_367#_c_458_n N_A_455_367#_M1005_s 0.00332344f $X=4.74 $Y=2.99
+ $X2=0 $Y2=0
cc_316 N_A_251_367#_c_445_n N_A_455_367#_c_494_n 0.0484121f $X=3.305 $Y=2.685
+ $X2=0 $Y2=0
cc_317 N_A_251_367#_c_458_n N_A_455_367#_c_494_n 0.00886059f $X=4.74 $Y=2.99
+ $X2=0 $Y2=0
cc_318 N_A_251_367#_c_446_n N_A_455_367#_c_494_n 0.013617f $X=3.39 $Y=2.685
+ $X2=0 $Y2=0
cc_319 N_A_251_367#_c_445_n N_A_455_367#_c_501_n 0.0170334f $X=3.305 $Y=2.685
+ $X2=0 $Y2=0
cc_320 N_A_251_367#_c_458_n N_A_455_367#_c_506_n 0.0139212f $X=4.74 $Y=2.99
+ $X2=0 $Y2=0
cc_321 N_A_251_367#_c_446_n N_A_455_367#_c_506_n 0.00581257f $X=3.39 $Y=2.685
+ $X2=0 $Y2=0
cc_322 N_A_251_367#_c_458_n N_Y_M1005_d 0.00490137f $X=4.74 $Y=2.99 $X2=0 $Y2=0
cc_323 N_A_251_367#_c_446_n N_Y_M1005_d 0.00650249f $X=3.39 $Y=2.685 $X2=0 $Y2=0
cc_324 N_A_251_367#_c_458_n N_Y_M1011_d 0.00332344f $X=4.74 $Y=2.99 $X2=0 $Y2=0
cc_325 N_A_251_367#_M1000_s N_Y_c_545_n 0.00419382f $X=4.695 $Y=1.835 $X2=0
+ $Y2=0
cc_326 N_A_251_367#_c_492_p N_Y_c_545_n 0.0135577f $X=4.835 $Y=2.435 $X2=0 $Y2=0
cc_327 N_A_251_367#_c_458_n N_Y_c_548_n 0.0159805f $X=4.74 $Y=2.99 $X2=0 $Y2=0
cc_328 N_A_455_367#_c_494_n N_Y_M1005_d 0.00626979f $X=3.81 $Y=2.345 $X2=0 $Y2=0
cc_329 N_A_455_367#_M1005_s N_Y_c_541_n 0.0037006f $X=3.835 $Y=1.835 $X2=0 $Y2=0
cc_330 N_A_455_367#_c_494_n N_Y_c_541_n 0.0149701f $X=3.81 $Y=2.345 $X2=0 $Y2=0
cc_331 N_A_455_367#_c_495_n N_Y_c_530_n 0.0136419f $X=2.415 $Y=2.005 $X2=0 $Y2=0
cc_332 N_A_455_367#_c_494_n N_Y_c_530_n 0.0694325f $X=3.81 $Y=2.345 $X2=0 $Y2=0
cc_333 N_A_455_367#_c_495_n N_A_251_47#_c_671_n 0.00730715f $X=2.415 $Y=2.005
+ $X2=0 $Y2=0
cc_334 N_Y_c_526_n N_VGND_c_619_n 0.0125145f $X=5.425 $Y=0.495 $X2=0 $Y2=0
cc_335 N_Y_c_526_n N_VGND_c_620_n 0.00964185f $X=5.425 $Y=0.495 $X2=0 $Y2=0
cc_336 N_Y_c_524_n N_A_251_47#_M1001_s 0.00179632f $X=4.32 $Y=1.105 $X2=0 $Y2=0
cc_337 N_Y_c_527_n N_A_251_47#_c_671_n 0.0159284f $X=3.545 $Y=1.245 $X2=0 $Y2=0
cc_338 N_Y_c_530_n N_A_251_47#_c_671_n 0.0180749f $X=3.71 $Y=1.835 $X2=0 $Y2=0
cc_339 N_Y_c_527_n N_A_251_47#_c_673_n 0.00847199f $X=3.545 $Y=1.245 $X2=0 $Y2=0
cc_340 N_Y_M1001_d N_A_251_47#_c_675_n 0.0058534f $X=3.4 $Y=0.345 $X2=0 $Y2=0
cc_341 N_Y_c_524_n N_A_251_47#_c_675_n 0.0231803f $X=4.32 $Y=1.105 $X2=0 $Y2=0
cc_342 N_Y_c_527_n N_A_251_47#_c_675_n 0.0220894f $X=3.545 $Y=1.245 $X2=0 $Y2=0
cc_343 N_Y_c_525_n N_A_423_47#_M1007_d 0.00261503f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_344 N_Y_M1001_d N_A_423_47#_c_716_n 0.00295113f $X=3.4 $Y=0.345 $X2=0 $Y2=0
cc_345 N_Y_M1013_d N_A_423_47#_c_716_n 0.00261964f $X=4.265 $Y=0.345 $X2=0 $Y2=0
cc_346 N_Y_c_524_n N_A_423_47#_c_716_n 0.00348752f $X=4.32 $Y=1.105 $X2=0 $Y2=0
cc_347 N_Y_c_560_n N_A_423_47#_c_716_n 0.0204295f $X=4.485 $Y=0.69 $X2=0 $Y2=0
cc_348 N_Y_c_525_n N_A_423_47#_c_716_n 0.00281285f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_349 N_Y_c_526_n N_A_423_47#_c_716_n 0.00498721f $X=5.425 $Y=0.495 $X2=0 $Y2=0
cc_350 N_Y_c_525_n N_A_423_47#_c_724_n 0.02172f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_351 N_VGND_c_620_n N_A_251_47#_M1009_s 0.00397496f $X=5.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_352 N_VGND_c_617_n N_A_251_47#_c_703_n 0.0138717f $X=1.7 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_620_n N_A_251_47#_c_703_n 0.00886411f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_M1017_d N_A_251_47#_c_671_n 0.00176461f $X=1.685 $Y=0.235 $X2=0
+ $Y2=0
cc_355 N_VGND_M1010_d N_A_251_47#_c_671_n 0.00225881f $X=2.545 $Y=0.235 $X2=0
+ $Y2=0
cc_356 N_VGND_c_658_p N_A_251_47#_c_671_n 0.0135055f $X=1.92 $Y=0.785 $X2=0
+ $Y2=0
cc_357 N_VGND_c_614_n N_A_251_47#_c_671_n 0.0514469f $X=2.685 $Y=0.78 $X2=0
+ $Y2=0
cc_358 N_VGND_c_614_n N_A_251_47#_c_673_n 0.00838689f $X=2.685 $Y=0.78 $X2=0
+ $Y2=0
cc_359 N_VGND_c_614_n N_A_251_47#_c_674_n 0.0111499f $X=2.685 $Y=0.78 $X2=0
+ $Y2=0
cc_360 N_VGND_c_614_n N_A_423_47#_M1003_s 0.00337359f $X=2.685 $Y=0.78 $X2=-0.19
+ $Y2=-0.245
cc_361 N_VGND_c_620_n N_A_423_47#_M1003_s 0.00223577f $X=5.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_362 N_VGND_M1010_d N_A_423_47#_c_716_n 0.00538092f $X=2.545 $Y=0.235 $X2=0
+ $Y2=0
cc_363 N_VGND_c_614_n N_A_423_47#_c_716_n 0.0190286f $X=2.685 $Y=0.78 $X2=0
+ $Y2=0
cc_364 N_VGND_c_619_n N_A_423_47#_c_716_n 0.023489f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_620_n N_A_423_47#_c_716_n 0.0127001f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_614_n N_A_423_47#_c_718_n 0.0154146f $X=2.685 $Y=0.78 $X2=0
+ $Y2=0
cc_367 N_VGND_c_619_n N_A_423_47#_c_718_n 0.170146f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_620_n N_A_423_47#_c_718_n 0.100237f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_369 N_A_251_47#_c_671_n N_A_423_47#_M1003_s 0.00176891f $X=3.02 $Y=1.15
+ $X2=-0.19 $Y2=-0.245
cc_370 N_A_251_47#_M1001_s N_A_423_47#_c_716_n 0.00177204f $X=3.835 $Y=0.345
+ $X2=0 $Y2=0
cc_371 N_A_251_47#_c_671_n N_A_423_47#_c_716_n 0.00514754f $X=3.02 $Y=1.15 $X2=0
+ $Y2=0
cc_372 N_A_251_47#_c_674_n N_A_423_47#_c_716_n 0.0150169f $X=3.21 $Y=0.7 $X2=0
+ $Y2=0
cc_373 N_A_251_47#_c_675_n N_A_423_47#_c_716_n 0.0522103f $X=3.975 $Y=0.71 $X2=0
+ $Y2=0
