# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux4_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__mux4_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.210000 9.475000 1.460000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.740000 1.080000 7.075000 1.410000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.770000 0.765000 6.085000 1.095000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.550000 4.350000 2.150000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  1.002000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.885000 1.045000 5.565000 1.275000 ;
        RECT 4.885000 1.275000 6.495000 1.375000 ;
        RECT 5.395000 1.375000 6.495000 1.445000 ;
        RECT 5.815000 1.445000 6.145000 1.760000 ;
        RECT 6.325000 1.445000 6.495000 1.590000 ;
        RECT 6.325000 1.590000 7.610000 1.760000 ;
        RECT 7.280000 1.080000 7.610000 1.590000 ;
        RECT 7.440000 1.760000 7.610000 2.545000 ;
        RECT 7.440000 2.545000 8.350000 2.715000 ;
        RECT 8.180000 1.640000 9.620000 2.150000 ;
        RECT 8.180000 2.150000 8.350000 2.545000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 1.470000 1.805000 1.800000 ;
        RECT 1.635000 1.800000 1.805000 2.545000 ;
        RECT 1.635000 2.545000 2.505000 2.715000 ;
        RECT 2.335000 1.550000 2.755000 1.890000 ;
        RECT 2.335000 1.890000 2.505000 2.545000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.265000 0.445000 3.065000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.625000  0.645000  1.795000 0.815000 ;
      RECT 0.625000  0.815000  0.795000 1.980000 ;
      RECT 0.625000  1.980000  1.455000 2.150000 ;
      RECT 0.645000  2.330000  0.975000 3.245000 ;
      RECT 0.905000  0.085000  1.235000 0.465000 ;
      RECT 0.975000  0.995000  2.155000 1.260000 ;
      RECT 1.205000  2.150000  1.455000 2.895000 ;
      RECT 1.205000  2.895000  3.285000 3.065000 ;
      RECT 1.465000  0.265000  1.795000 0.645000 ;
      RECT 1.975000  0.265000  2.145000 0.995000 ;
      RECT 1.985000  1.260000  2.155000 2.365000 ;
      RECT 2.325000  0.265000  3.565000 0.435000 ;
      RECT 2.325000  0.435000  2.655000 0.725000 ;
      RECT 2.335000  0.990000  3.215000 1.320000 ;
      RECT 2.685000  2.165000  3.765000 2.335000 ;
      RECT 2.685000  2.335000  2.935000 2.715000 ;
      RECT 2.885000  0.615000  3.215000 0.990000 ;
      RECT 3.045000  1.320000  3.215000 1.655000 ;
      RECT 3.045000  1.655000  3.415000 1.985000 ;
      RECT 3.115000  2.515000  5.285000 2.685000 ;
      RECT 3.115000  2.685000  3.285000 2.895000 ;
      RECT 3.395000  0.435000  3.565000 1.125000 ;
      RECT 3.395000  1.125000  4.355000 1.295000 ;
      RECT 3.595000  1.295000  3.765000 2.165000 ;
      RECT 3.755000  0.085000  4.005000 0.945000 ;
      RECT 3.855000  2.865000  4.185000 3.245000 ;
      RECT 4.185000  0.265000  6.435000 0.435000 ;
      RECT 4.185000  0.435000  4.355000 1.125000 ;
      RECT 4.535000  0.615000  5.355000 0.865000 ;
      RECT 4.535000  0.865000  4.705000 2.515000 ;
      RECT 4.885000  1.585000  5.215000 1.745000 ;
      RECT 4.885000  1.745000  5.635000 1.915000 ;
      RECT 4.955000  2.095000  5.285000 2.515000 ;
      RECT 4.955000  2.685000  5.285000 3.065000 ;
      RECT 5.465000  1.915000  5.635000 1.940000 ;
      RECT 5.465000  1.940000  7.260000 2.110000 ;
      RECT 6.265000  0.435000  6.435000 0.730000 ;
      RECT 6.265000  0.730000  7.960000 0.900000 ;
      RECT 6.580000  2.290000  6.910000 3.245000 ;
      RECT 6.615000  0.085000  6.865000 0.550000 ;
      RECT 7.090000  2.110000  7.260000 2.895000 ;
      RECT 7.090000  2.895000  8.805000 3.065000 ;
      RECT 7.545000  0.265000  7.960000 0.730000 ;
      RECT 7.790000  0.900000  7.960000 2.365000 ;
      RECT 8.140000  0.765000  8.470000 0.860000 ;
      RECT 8.140000  0.860000  9.970000 1.030000 ;
      RECT 8.635000  2.330000  9.970000 2.500000 ;
      RECT 8.635000  2.500000  8.805000 2.895000 ;
      RECT 8.845000  0.085000  9.175000 0.675000 ;
      RECT 8.985000  2.680000  9.315000 3.245000 ;
      RECT 9.515000  2.500000  9.970000 3.065000 ;
      RECT 9.635000  0.265000  9.970000 0.860000 ;
      RECT 9.800000  1.030000  9.970000 2.330000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__mux4_lp
END LIBRARY
