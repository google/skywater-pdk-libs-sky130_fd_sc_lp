* NGSPICE file created from sky130_fd_sc_lp__einvp_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__einvp_0 A TE VGND VNB VPB VPWR Z
M1000 VPWR TE a_32_70# VPB phighvt w=420000u l=150000u
+  ad=2.158e+11p pd=2.03e+06u as=1.113e+11p ps=1.37e+06u
M1001 Z A a_220_484# VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=1.536e+11p ps=1.76e+06u
M1002 a_220_484# a_32_70# VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND TE a_32_70# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.113e+11p ps=1.37e+06u
M1004 a_201_70# TE VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1005 Z A a_201_70# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

