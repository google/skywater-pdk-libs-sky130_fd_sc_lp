* File: sky130_fd_sc_lp__or3b_lp.spice
* Created: Fri Aug 28 11:24:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or3b_lp.pex.spice"
.subckt sky130_fd_sc_lp__or3b_lp  VNB VPB C_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1002 A_114_47# N_C_N_M1002_g N_A_27_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_C_N_M1014_g A_114_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1003 A_272_47# N_A_27_47#_M1003_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_350_47#_M1004_d N_A_27_47#_M1004_g A_272_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_466_185# N_B_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.5
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_350_47#_M1006_d N_B_M1006_g A_466_185# VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.0441 PD=1.2 PS=0.63 NRD=61.428 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 A_640_101# N_A_M1013_g N_A_350_47#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1134 PD=0.66 PS=1.2 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g A_640_101# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1007 A_804_101# N_A_350_47#_M1007_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_350_47#_M1000_g A_804_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_C_N_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1010 N_A_350_47#_M1010_d N_A_27_47#_M1010_g N_A_263_373#_M1010_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1008 A_628_419# N_B_M1008_g N_A_263_373#_M1008_s VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g A_628_419# VPB PHIGHVT L=0.25 W=1 AD=0.195
+ AS=0.12 PD=1.39 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1011 N_X_M1011_d N_A_350_47#_M1011_g N_VPWR_M1012_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.195 PD=2.57 PS=1.39 NRD=0 NRS=21.67 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX15_noxref VNB VPB NWDIODE A=9.60895 P=14.15
*
.include "sky130_fd_sc_lp__or3b_lp.pxi.spice"
*
.ends
*
*
