* NGSPICE file created from sky130_fd_sc_lp__fa_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 a_941_419# B VPWR VPB phighvt w=640000u l=150000u
+  ad=5.4185e+11p pd=4.39e+06u as=2.4209e+12p ps=1.786e+07u
M1001 VGND A a_309_131# VNB nshort w=420000u l=150000u
+  ad=1.7743e+12p pd=1.445e+07u as=3.5865e+11p ps=3.49e+06u
M1002 a_710_119# A VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1003 COUT a_395_398# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1004 COUT a_395_398# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1005 VPWR CIN a_941_419# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_395_398# B a_1653_137# VNB nshort w=420000u l=150000u
+  ad=2.625e+11p pd=2.93e+06u as=8.82e+10p ps=1.26e+06u
M1007 VGND a_84_21# SUM VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1008 SUM a_84_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1653_137# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_710_419# A VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1011 a_395_398# CIN a_309_398# VPB phighvt w=640000u l=150000u
+  ad=3.648e+11p pd=3.7e+06u as=3.488e+11p ps=3.65e+06u
M1012 VPWR A a_309_398# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_782_419# B a_710_419# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1014 a_395_398# B a_1653_367# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1015 VGND CIN a_940_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1016 VGND a_395_398# COUT VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_84_21# CIN a_782_419# VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1018 a_395_398# CIN a_309_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_84_21# CIN a_782_119# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1020 SUM a_84_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1021 VPWR A a_941_419# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_940_119# a_395_398# a_84_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_309_131# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_940_119# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1653_367# A VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND A a_940_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_309_398# B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_395_398# COUT VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_782_119# B a_710_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_84_21# SUM VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_941_419# a_395_398# a_84_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

