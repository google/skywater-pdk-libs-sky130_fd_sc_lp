* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 a_110_70# a_250_443# a_614_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND SCE a_110_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_700_133# a_742_107# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_614_133# a_250_443# a_746_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_110_468# GATE a_110_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_110_70# a_282_70# a_614_133# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_614_133# a_282_70# a_700_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_614_133# a_742_107# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR a_614_133# a_742_107# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 GCLK a_1235_429# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR a_1235_429# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VPWR SCE a_110_468# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_1174_74# a_742_107# a_1235_429# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1235_429# a_742_107# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_110_70# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_1235_429# GCLK VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_250_443# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 VGND a_250_443# a_282_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_746_457# a_742_107# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VPWR a_250_443# a_282_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_250_443# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR CLK a_1235_429# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 VGND CLK a_1174_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 GCLK a_1235_429# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
