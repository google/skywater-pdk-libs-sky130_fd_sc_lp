* File: sky130_fd_sc_lp__a31o_0.pxi.spice
* Created: Fri Aug 28 09:58:58 2020
* 
x_PM_SKY130_FD_SC_LP__A31O_0%A_86_241# N_A_86_241#_M1009_d N_A_86_241#_M1007_d
+ N_A_86_241#_M1005_g N_A_86_241#_M1004_g N_A_86_241#_c_70_n N_A_86_241#_c_78_n
+ N_A_86_241#_c_71_n N_A_86_241#_c_72_n N_A_86_241#_c_73_n N_A_86_241#_c_74_n
+ N_A_86_241#_c_79_n N_A_86_241#_c_133_p N_A_86_241#_c_75_n N_A_86_241#_c_107_p
+ N_A_86_241#_c_80_n N_A_86_241#_c_81_n N_A_86_241#_c_82_n
+ PM_SKY130_FD_SC_LP__A31O_0%A_86_241#
x_PM_SKY130_FD_SC_LP__A31O_0%A3 N_A3_c_166_n N_A3_M1001_g N_A3_M1006_g
+ N_A3_c_169_n A3 N_A3_c_171_n PM_SKY130_FD_SC_LP__A31O_0%A3
x_PM_SKY130_FD_SC_LP__A31O_0%A2 N_A2_M1008_g N_A2_M1000_g N_A2_c_215_n
+ N_A2_c_216_n A2 A2 N_A2_c_218_n PM_SKY130_FD_SC_LP__A31O_0%A2
x_PM_SKY130_FD_SC_LP__A31O_0%A1 N_A1_M1003_g N_A1_M1009_g N_A1_c_255_n
+ N_A1_c_262_n N_A1_c_256_n N_A1_c_257_n A1 A1 N_A1_c_259_n
+ PM_SKY130_FD_SC_LP__A31O_0%A1
x_PM_SKY130_FD_SC_LP__A31O_0%B1 N_B1_c_302_n N_B1_M1007_g N_B1_M1002_g
+ N_B1_c_299_n B1 B1 B1 N_B1_c_301_n PM_SKY130_FD_SC_LP__A31O_0%B1
x_PM_SKY130_FD_SC_LP__A31O_0%X N_X_M1005_s N_X_M1004_s X X X X X X X X
+ N_X_c_329_n X PM_SKY130_FD_SC_LP__A31O_0%X
x_PM_SKY130_FD_SC_LP__A31O_0%VPWR N_VPWR_M1004_d N_VPWR_M1008_d N_VPWR_c_350_n
+ N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_355_n
+ VPWR N_VPWR_c_356_n N_VPWR_c_349_n PM_SKY130_FD_SC_LP__A31O_0%VPWR
x_PM_SKY130_FD_SC_LP__A31O_0%A_266_483# N_A_266_483#_M1001_d
+ N_A_266_483#_M1003_d N_A_266_483#_c_386_n N_A_266_483#_c_387_n
+ N_A_266_483#_c_388_n N_A_266_483#_c_389_n
+ PM_SKY130_FD_SC_LP__A31O_0%A_266_483#
x_PM_SKY130_FD_SC_LP__A31O_0%VGND N_VGND_M1005_d N_VGND_M1002_d N_VGND_c_411_n
+ N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n VGND
+ N_VGND_c_416_n N_VGND_c_417_n PM_SKY130_FD_SC_LP__A31O_0%VGND
cc_1 VNB N_A_86_241#_M1005_g 0.0477412f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.46
cc_2 VNB N_A_86_241#_c_70_n 0.022014f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.84
cc_3 VNB N_A_86_241#_c_71_n 0.00672556f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.37
cc_4 VNB N_A_86_241#_c_72_n 0.0198396f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.37
cc_5 VNB N_A_86_241#_c_73_n 0.0149101f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=0.755
cc_6 VNB N_A_86_241#_c_74_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.755
cc_7 VNB N_A_86_241#_c_75_n 0.0032914f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=0.46
cc_8 VNB N_A3_c_166_n 0.0187814f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=2.415
cc_9 VNB N_A3_M1001_g 0.00318318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A3_M1006_g 0.0257481f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.46
cc_11 VNB N_A3_c_169_n 0.0172848f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.99
cc_12 VNB A3 0.00703561f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.735
cc_13 VNB N_A3_c_171_n 0.0176633f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.37
cc_14 VNB N_A2_M1008_g 0.00807618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_M1000_g 0.0198955f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.205
cc_16 VNB N_A2_c_215_n 0.0230412f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.99
cc_17 VNB N_A2_c_216_n 0.0162396f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.735
cc_18 VNB A2 0.00267291f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.735
cc_19 VNB N_A2_c_218_n 0.0162843f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.84
cc_20 VNB N_A1_M1009_g 0.0209435f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.205
cc_21 VNB N_A1_c_255_n 0.00909231f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.99
cc_22 VNB N_A1_c_256_n 0.0209278f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.37
cc_23 VNB N_A1_c_257_n 0.0143869f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.205
cc_24 VNB A1 0.00846892f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.84
cc_25 VNB N_A1_c_259_n 0.0152604f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.37
cc_26 VNB N_B1_M1002_g 0.0264939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B1_c_299_n 0.0096819f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.46
cc_28 VNB B1 0.0375842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B1_c_301_n 0.100972f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.705
cc_30 VNB X 0.0580371f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.755
cc_31 VNB N_X_c_329_n 0.0118563f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=0.755
cc_32 VNB N_VPWR_c_349_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.775 $Y2=2.545
cc_33 VNB N_VGND_c_411_n 0.00609423f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.46
cc_34 VNB N_VGND_c_412_n 0.0155587f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.99
cc_35 VNB N_VGND_c_413_n 0.0181839f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.735
cc_36 VNB N_VGND_c_414_n 0.0205f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.205
cc_37 VNB N_VGND_c_415_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.84
cc_38 VNB N_VGND_c_416_n 0.0407966f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.37
cc_39 VNB N_VGND_c_417_n 0.203059f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.875
cc_40 VPB N_A_86_241#_M1004_g 0.0393476f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=2.735
cc_41 VPB N_A_86_241#_c_70_n 0.0143915f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.84
cc_42 VPB N_A_86_241#_c_78_n 0.0279782f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.99
cc_43 VPB N_A_86_241#_c_79_n 0.0449902f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=1.79
cc_44 VPB N_A_86_241#_c_80_n 0.00873416f $X=-0.19 $Y=1.655 $X2=2.775 $Y2=2.545
cc_45 VPB N_A_86_241#_c_81_n 0.0227188f $X=-0.19 $Y=1.655 $X2=2.76 $Y2=2.56
cc_46 VPB N_A_86_241#_c_82_n 0.00700943f $X=-0.19 $Y=1.655 $X2=2.775 $Y2=2.395
cc_47 VPB N_A3_M1001_g 0.0510779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_M1008_g 0.0485231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A1_M1003_g 0.0382913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A1_c_255_n 0.00543051f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=1.99
cc_51 VPB N_A1_c_262_n 0.0133083f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=2.735
cc_52 VPB N_B1_c_302_n 0.0203239f $X=-0.19 $Y=1.655 $X2=2.26 $Y2=0.25
cc_53 VPB N_B1_c_299_n 0.067129f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.46
cc_54 VPB B1 0.020876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB X 0.0408825f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.755
cc_56 VPB X 0.0501435f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.37
cc_57 VPB N_VPWR_c_350_n 0.00997297f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.46
cc_58 VPB N_VPWR_c_351_n 0.00821482f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=2.735
cc_59 VPB N_VPWR_c_352_n 0.0249581f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.205
cc_60 VPB N_VPWR_c_353_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.84
cc_61 VPB N_VPWR_c_354_n 0.0167145f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.99
cc_62 VPB N_VPWR_c_355_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_63 VPB N_VPWR_c_356_n 0.039395f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=2.395
cc_64 VPB N_VPWR_c_349_n 0.0731763f $X=-0.19 $Y=1.655 $X2=2.775 $Y2=2.545
cc_65 VPB N_A_266_483#_c_386_n 0.0062013f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.46
cc_66 VPB N_A_266_483#_c_387_n 0.00910988f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=1.99
cc_67 VPB N_A_266_483#_c_388_n 0.00480673f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=2.735
cc_68 VPB N_A_266_483#_c_389_n 0.00544214f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.37
cc_69 N_A_86_241#_c_71_n N_A3_c_166_n 4.01275e-19 $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_70 N_A_86_241#_c_72_n N_A3_c_166_n 0.0107517f $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_71 N_A_86_241#_c_70_n N_A3_M1001_g 0.00675853f $X=0.665 $Y=1.84 $X2=0 $Y2=0
cc_72 N_A_86_241#_c_78_n N_A3_M1001_g 0.0336575f $X=0.665 $Y=1.99 $X2=0 $Y2=0
cc_73 N_A_86_241#_c_71_n N_A3_M1001_g 5.90881e-19 $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_74 N_A_86_241#_c_79_n N_A3_M1001_g 0.0156266f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_75 N_A_86_241#_M1005_g N_A3_M1006_g 0.0146818f $X=0.605 $Y=0.46 $X2=0 $Y2=0
cc_76 N_A_86_241#_c_71_n N_A3_M1006_g 0.00156821f $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_77 N_A_86_241#_c_73_n N_A3_M1006_g 0.00488757f $X=1.235 $Y=0.755 $X2=0 $Y2=0
cc_78 N_A_86_241#_c_75_n N_A3_M1006_g 0.0163633f $X=1.405 $Y=0.46 $X2=0 $Y2=0
cc_79 N_A_86_241#_c_70_n N_A3_c_169_n 0.0107517f $X=0.665 $Y=1.84 $X2=0 $Y2=0
cc_80 N_A_86_241#_c_71_n N_A3_c_169_n 5.72538e-19 $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_81 N_A_86_241#_c_79_n N_A3_c_169_n 0.0059382f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_82 N_A_86_241#_M1005_g A3 2.21539e-19 $X=0.605 $Y=0.46 $X2=0 $Y2=0
cc_83 N_A_86_241#_c_71_n A3 0.0293437f $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_84 N_A_86_241#_c_72_n A3 0.0011536f $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_85 N_A_86_241#_c_73_n A3 0.0181736f $X=1.235 $Y=0.755 $X2=0 $Y2=0
cc_86 N_A_86_241#_c_79_n A3 0.0256865f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_87 N_A_86_241#_c_75_n A3 0.0100471f $X=1.405 $Y=0.46 $X2=0 $Y2=0
cc_88 N_A_86_241#_M1005_g N_A3_c_171_n 0.0103047f $X=0.605 $Y=0.46 $X2=0 $Y2=0
cc_89 N_A_86_241#_c_71_n N_A3_c_171_n 0.00246279f $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_90 N_A_86_241#_c_73_n N_A3_c_171_n 0.00600124f $X=1.235 $Y=0.755 $X2=0 $Y2=0
cc_91 N_A_86_241#_c_79_n N_A2_M1008_g 0.010706f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_92 N_A_86_241#_c_75_n N_A2_M1000_g 0.0026044f $X=1.405 $Y=0.46 $X2=0 $Y2=0
cc_93 N_A_86_241#_c_107_p N_A2_M1000_g 0.0156065f $X=2.44 $Y=0.46 $X2=0 $Y2=0
cc_94 N_A_86_241#_c_79_n N_A2_c_216_n 0.00344545f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_95 N_A_86_241#_c_79_n A2 0.0184446f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_96 N_A_86_241#_c_75_n A2 0.00350567f $X=1.405 $Y=0.46 $X2=0 $Y2=0
cc_97 N_A_86_241#_c_107_p A2 0.0175408f $X=2.44 $Y=0.46 $X2=0 $Y2=0
cc_98 N_A_86_241#_c_107_p N_A2_c_218_n 0.00274298f $X=2.44 $Y=0.46 $X2=0 $Y2=0
cc_99 N_A_86_241#_c_82_n N_A1_M1003_g 0.00285314f $X=2.775 $Y=2.395 $X2=0 $Y2=0
cc_100 N_A_86_241#_c_107_p N_A1_M1009_g 0.0123051f $X=2.44 $Y=0.46 $X2=0 $Y2=0
cc_101 N_A_86_241#_c_79_n N_A1_c_255_n 0.00458119f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_102 N_A_86_241#_c_79_n N_A1_c_262_n 0.00989364f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_103 N_A_86_241#_c_82_n N_A1_c_262_n 4.48562e-19 $X=2.775 $Y=2.395 $X2=0 $Y2=0
cc_104 N_A_86_241#_c_79_n N_A1_c_257_n 0.00271078f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_105 N_A_86_241#_c_79_n A1 0.0271067f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_106 N_A_86_241#_c_107_p A1 0.0263003f $X=2.44 $Y=0.46 $X2=0 $Y2=0
cc_107 N_A_86_241#_c_107_p N_A1_c_259_n 0.00283928f $X=2.44 $Y=0.46 $X2=0 $Y2=0
cc_108 N_A_86_241#_c_82_n N_B1_c_302_n 0.00338303f $X=2.775 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_86_241#_c_79_n N_B1_c_299_n 0.0223921f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_110 N_A_86_241#_c_80_n N_B1_c_299_n 0.00180564f $X=2.775 $Y=2.545 $X2=0 $Y2=0
cc_111 N_A_86_241#_c_82_n N_B1_c_299_n 0.0312781f $X=2.775 $Y=2.395 $X2=0 $Y2=0
cc_112 N_A_86_241#_c_79_n B1 0.0111895f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_113 N_A_86_241#_c_74_n N_X_M1005_s 2.1455e-19 $X=0.76 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_86_241#_M1005_g X 0.00855134f $X=0.605 $Y=0.46 $X2=0 $Y2=0
cc_115 N_A_86_241#_M1004_g X 0.0112628f $X=0.825 $Y=2.735 $X2=0 $Y2=0
cc_116 N_A_86_241#_c_71_n X 0.0670563f $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_117 N_A_86_241#_c_72_n X 0.0218401f $X=0.595 $Y=1.37 $X2=0 $Y2=0
cc_118 N_A_86_241#_c_74_n X 0.0147638f $X=0.76 $Y=0.755 $X2=0 $Y2=0
cc_119 N_A_86_241#_c_133_p X 0.0139501f $X=0.76 $Y=1.79 $X2=0 $Y2=0
cc_120 N_A_86_241#_M1005_g N_X_c_329_n 0.00299046f $X=0.605 $Y=0.46 $X2=0 $Y2=0
cc_121 N_A_86_241#_c_74_n N_X_c_329_n 0.00262888f $X=0.76 $Y=0.755 $X2=0 $Y2=0
cc_122 N_A_86_241#_M1004_g X 9.63756e-19 $X=0.825 $Y=2.735 $X2=0 $Y2=0
cc_123 N_A_86_241#_c_78_n X 0.00852643f $X=0.665 $Y=1.99 $X2=0 $Y2=0
cc_124 N_A_86_241#_c_133_p X 0.00877031f $X=0.76 $Y=1.79 $X2=0 $Y2=0
cc_125 N_A_86_241#_M1004_g N_VPWR_c_350_n 0.00290389f $X=0.825 $Y=2.735 $X2=0
+ $Y2=0
cc_126 N_A_86_241#_c_79_n N_VPWR_c_350_n 0.0100201f $X=2.625 $Y=1.79 $X2=0 $Y2=0
cc_127 N_A_86_241#_M1004_g N_VPWR_c_352_n 0.00545548f $X=0.825 $Y=2.735 $X2=0
+ $Y2=0
cc_128 N_A_86_241#_c_81_n N_VPWR_c_356_n 0.0213627f $X=2.76 $Y=2.56 $X2=0 $Y2=0
cc_129 N_A_86_241#_M1004_g N_VPWR_c_349_n 0.0113151f $X=0.825 $Y=2.735 $X2=0
+ $Y2=0
cc_130 N_A_86_241#_c_81_n N_VPWR_c_349_n 0.0115856f $X=2.76 $Y=2.56 $X2=0 $Y2=0
cc_131 N_A_86_241#_c_79_n N_A_266_483#_c_387_n 0.0610318f $X=2.625 $Y=1.79 $X2=0
+ $Y2=0
cc_132 N_A_86_241#_c_82_n N_A_266_483#_c_387_n 0.0141882f $X=2.775 $Y=2.395
+ $X2=0 $Y2=0
cc_133 N_A_86_241#_c_79_n N_A_266_483#_c_388_n 0.0214928f $X=2.625 $Y=1.79 $X2=0
+ $Y2=0
cc_134 N_A_86_241#_c_82_n N_A_266_483#_c_389_n 0.0161343f $X=2.775 $Y=2.395
+ $X2=0 $Y2=0
cc_135 N_A_86_241#_c_74_n N_VGND_M1005_d 0.00130154f $X=0.76 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_86_241#_M1005_g N_VGND_c_411_n 0.00496169f $X=0.605 $Y=0.46 $X2=0
+ $Y2=0
cc_137 N_A_86_241#_c_73_n N_VGND_c_411_n 0.0237572f $X=1.235 $Y=0.755 $X2=0
+ $Y2=0
cc_138 N_A_86_241#_c_74_n N_VGND_c_411_n 0.00199859f $X=0.76 $Y=0.755 $X2=0
+ $Y2=0
cc_139 N_A_86_241#_c_75_n N_VGND_c_411_n 0.0151686f $X=1.405 $Y=0.46 $X2=0 $Y2=0
cc_140 N_A_86_241#_M1005_g N_VGND_c_414_n 0.00406355f $X=0.605 $Y=0.46 $X2=0
+ $Y2=0
cc_141 N_A_86_241#_c_74_n N_VGND_c_414_n 0.00304654f $X=0.76 $Y=0.755 $X2=0
+ $Y2=0
cc_142 N_A_86_241#_c_73_n N_VGND_c_416_n 0.0028261f $X=1.235 $Y=0.755 $X2=0
+ $Y2=0
cc_143 N_A_86_241#_c_75_n N_VGND_c_416_n 0.00784459f $X=1.405 $Y=0.46 $X2=0
+ $Y2=0
cc_144 N_A_86_241#_c_107_p N_VGND_c_416_n 0.0567171f $X=2.44 $Y=0.46 $X2=0 $Y2=0
cc_145 N_A_86_241#_M1005_g N_VGND_c_417_n 0.00719663f $X=0.605 $Y=0.46 $X2=0
+ $Y2=0
cc_146 N_A_86_241#_c_73_n N_VGND_c_417_n 0.00591918f $X=1.235 $Y=0.755 $X2=0
+ $Y2=0
cc_147 N_A_86_241#_c_74_n N_VGND_c_417_n 0.00493807f $X=0.76 $Y=0.755 $X2=0
+ $Y2=0
cc_148 N_A_86_241#_c_75_n N_VGND_c_417_n 0.00577896f $X=1.405 $Y=0.46 $X2=0
+ $Y2=0
cc_149 N_A_86_241#_c_107_p N_VGND_c_417_n 0.0433539f $X=2.44 $Y=0.46 $X2=0 $Y2=0
cc_150 N_A_86_241#_c_107_p A_272_50# 0.0084824f $X=2.44 $Y=0.46 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_86_241#_c_107_p A_361_50# 0.00753099f $X=2.44 $Y=0.46 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A3_M1001_g N_A2_M1008_g 0.04166f $X=1.255 $Y=2.735 $X2=0 $Y2=0
cc_153 N_A3_c_169_n N_A2_M1008_g 0.00529228f $X=1.18 $Y=1.6 $X2=0 $Y2=0
cc_154 N_A3_M1006_g N_A2_M1000_g 0.0304844f $X=1.285 $Y=0.46 $X2=0 $Y2=0
cc_155 A3 N_A2_c_215_n 0.00174257f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A3_c_171_n N_A2_c_215_n 0.01418f $X=1.165 $Y=1.095 $X2=0 $Y2=0
cc_157 N_A3_c_166_n N_A2_c_216_n 0.01418f $X=1.18 $Y=1.42 $X2=0 $Y2=0
cc_158 N_A3_M1006_g A2 0.00130376f $X=1.285 $Y=0.46 $X2=0 $Y2=0
cc_159 A3 A2 0.0307648f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A3_c_171_n A2 6.24433e-19 $X=1.165 $Y=1.095 $X2=0 $Y2=0
cc_161 N_A3_M1006_g N_A2_c_218_n 0.01418f $X=1.285 $Y=0.46 $X2=0 $Y2=0
cc_162 N_A3_M1001_g N_VPWR_c_350_n 0.00169173f $X=1.255 $Y=2.735 $X2=0 $Y2=0
cc_163 N_A3_M1001_g N_VPWR_c_354_n 0.00545548f $X=1.255 $Y=2.735 $X2=0 $Y2=0
cc_164 N_A3_M1001_g N_VPWR_c_349_n 0.0103349f $X=1.255 $Y=2.735 $X2=0 $Y2=0
cc_165 N_A3_M1001_g N_A_266_483#_c_386_n 0.00496711f $X=1.255 $Y=2.735 $X2=0
+ $Y2=0
cc_166 N_A3_M1001_g N_A_266_483#_c_388_n 0.00568793f $X=1.255 $Y=2.735 $X2=0
+ $Y2=0
cc_167 N_A3_M1006_g N_VGND_c_411_n 0.00567415f $X=1.285 $Y=0.46 $X2=0 $Y2=0
cc_168 N_A3_M1006_g N_VGND_c_416_n 0.0036741f $X=1.285 $Y=0.46 $X2=0 $Y2=0
cc_169 N_A3_M1006_g N_VGND_c_417_n 0.00592531f $X=1.285 $Y=0.46 $X2=0 $Y2=0
cc_170 N_A2_M1000_g N_A1_M1009_g 0.0311687f $X=1.73 $Y=0.46 $X2=0 $Y2=0
cc_171 N_A2_M1008_g N_A1_c_255_n 0.00967031f $X=1.685 $Y=2.735 $X2=0 $Y2=0
cc_172 N_A2_M1008_g N_A1_c_262_n 0.0362265f $X=1.685 $Y=2.735 $X2=0 $Y2=0
cc_173 N_A2_c_215_n N_A1_c_256_n 0.0138106f $X=1.735 $Y=1.345 $X2=0 $Y2=0
cc_174 N_A2_c_216_n N_A1_c_257_n 0.0138106f $X=1.735 $Y=1.51 $X2=0 $Y2=0
cc_175 A2 A1 0.056442f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_176 N_A2_c_218_n A1 0.00431759f $X=1.735 $Y=1.005 $X2=0 $Y2=0
cc_177 A2 N_A1_c_259_n 6.24336e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_178 N_A2_c_218_n N_A1_c_259_n 0.0138106f $X=1.735 $Y=1.005 $X2=0 $Y2=0
cc_179 N_A2_M1008_g N_VPWR_c_351_n 0.00166462f $X=1.685 $Y=2.735 $X2=0 $Y2=0
cc_180 N_A2_M1008_g N_VPWR_c_354_n 0.00545548f $X=1.685 $Y=2.735 $X2=0 $Y2=0
cc_181 N_A2_M1008_g N_VPWR_c_349_n 0.0103485f $X=1.685 $Y=2.735 $X2=0 $Y2=0
cc_182 N_A2_M1008_g N_A_266_483#_c_386_n 0.0027683f $X=1.685 $Y=2.735 $X2=0
+ $Y2=0
cc_183 N_A2_M1008_g N_A_266_483#_c_387_n 0.0147457f $X=1.685 $Y=2.735 $X2=0
+ $Y2=0
cc_184 N_A2_M1000_g N_VGND_c_416_n 0.00355856f $X=1.73 $Y=0.46 $X2=0 $Y2=0
cc_185 N_A2_M1000_g N_VGND_c_417_n 0.00541034f $X=1.73 $Y=0.46 $X2=0 $Y2=0
cc_186 N_A1_M1009_g N_B1_M1002_g 0.0160387f $X=2.185 $Y=0.46 $X2=0 $Y2=0
cc_187 A1 N_B1_M1002_g 4.6864e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_188 N_A1_M1003_g N_B1_c_299_n 0.021757f $X=2.115 $Y=2.735 $X2=0 $Y2=0
cc_189 N_A1_c_255_n N_B1_c_299_n 0.0144452f $X=2.165 $Y=1.75 $X2=0 $Y2=0
cc_190 A1 B1 0.0190377f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_191 N_A1_c_259_n B1 0.00143195f $X=2.275 $Y=1.005 $X2=0 $Y2=0
cc_192 A1 N_B1_c_301_n 0.0028745f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_193 N_A1_c_259_n N_B1_c_301_n 0.0455963f $X=2.275 $Y=1.005 $X2=0 $Y2=0
cc_194 N_A1_M1003_g N_VPWR_c_351_n 0.00286411f $X=2.115 $Y=2.735 $X2=0 $Y2=0
cc_195 N_A1_M1003_g N_VPWR_c_356_n 0.00545548f $X=2.115 $Y=2.735 $X2=0 $Y2=0
cc_196 N_A1_M1003_g N_VPWR_c_349_n 0.0103485f $X=2.115 $Y=2.735 $X2=0 $Y2=0
cc_197 N_A1_M1003_g N_A_266_483#_c_387_n 0.0150264f $X=2.115 $Y=2.735 $X2=0
+ $Y2=0
cc_198 N_A1_c_262_n N_A_266_483#_c_387_n 0.00278277f $X=2.165 $Y=1.9 $X2=0 $Y2=0
cc_199 N_A1_M1003_g N_A_266_483#_c_389_n 0.00276049f $X=2.115 $Y=2.735 $X2=0
+ $Y2=0
cc_200 N_A1_M1009_g N_VGND_c_413_n 9.92194e-19 $X=2.185 $Y=0.46 $X2=0 $Y2=0
cc_201 N_A1_M1009_g N_VGND_c_416_n 0.00355856f $X=2.185 $Y=0.46 $X2=0 $Y2=0
cc_202 N_A1_M1009_g N_VGND_c_417_n 0.00560863f $X=2.185 $Y=0.46 $X2=0 $Y2=0
cc_203 N_B1_c_302_n N_VPWR_c_356_n 0.00545548f $X=2.545 $Y=2.29 $X2=0 $Y2=0
cc_204 N_B1_c_302_n N_VPWR_c_349_n 0.0115584f $X=2.545 $Y=2.29 $X2=0 $Y2=0
cc_205 N_B1_c_299_n N_A_266_483#_c_387_n 0.00120257f $X=2.755 $Y=2.14 $X2=0
+ $Y2=0
cc_206 N_B1_c_299_n N_A_266_483#_c_389_n 0.00171997f $X=2.755 $Y=2.14 $X2=0
+ $Y2=0
cc_207 N_B1_M1002_g N_VGND_c_413_n 0.0116455f $X=2.725 $Y=0.46 $X2=0 $Y2=0
cc_208 B1 N_VGND_c_413_n 0.00973921f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_209 N_B1_c_301_n N_VGND_c_413_n 0.00840821f $X=3.09 $Y=1.005 $X2=0 $Y2=0
cc_210 N_B1_M1002_g N_VGND_c_416_n 0.00473366f $X=2.725 $Y=0.46 $X2=0 $Y2=0
cc_211 N_B1_M1002_g N_VGND_c_417_n 0.00853602f $X=2.725 $Y=0.46 $X2=0 $Y2=0
cc_212 B1 N_VGND_c_417_n 0.00739521f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_213 X N_VPWR_c_350_n 0.00327831f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_214 X N_VPWR_c_352_n 0.0468114f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_215 X N_VPWR_c_349_n 0.0253871f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_216 N_X_c_329_n N_VGND_c_414_n 0.0263427f $X=0.39 $Y=0.375 $X2=0 $Y2=0
cc_217 N_X_c_329_n N_VGND_c_417_n 0.0175101f $X=0.39 $Y=0.375 $X2=0 $Y2=0
cc_218 N_VPWR_c_350_n N_A_266_483#_c_386_n 0.00305423f $X=1.04 $Y=2.56 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_351_n N_A_266_483#_c_386_n 0.00304519f $X=1.9 $Y=2.56 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_354_n N_A_266_483#_c_386_n 0.0188536f $X=1.775 $Y=3.33 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_349_n N_A_266_483#_c_386_n 0.0102248f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_351_n N_A_266_483#_c_387_n 0.0209462f $X=1.9 $Y=2.56 $X2=0 $Y2=0
cc_223 N_VPWR_c_351_n N_A_266_483#_c_389_n 0.00304078f $X=1.9 $Y=2.56 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_356_n N_A_266_483#_c_389_n 0.0184952f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_349_n N_A_266_483#_c_389_n 0.0100304f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
