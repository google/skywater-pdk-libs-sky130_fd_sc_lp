# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o211a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o211a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 1.210000 2.320000 2.120000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 1.210000 1.815000 2.120000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.930000 1.210000 1.285000 1.470000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.210000 0.355000 1.575000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 0.255000 3.065000 0.955000 ;
        RECT 2.735000 0.955000 3.200000 1.125000 ;
        RECT 3.030000 1.125000 3.200000 1.190000 ;
        RECT 3.030000 1.190000 3.220000 1.250000 ;
        RECT 3.030000 1.250000 3.485000 2.120000 ;
        RECT 3.030000 2.120000 3.225000 2.460000 ;
        RECT 3.035000 2.460000 3.225000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.095000  0.255000 0.425000 0.860000 ;
      RECT 0.095000  0.860000 0.705000 1.040000 ;
      RECT 0.265000  1.745000 1.425000 1.915000 ;
      RECT 0.265000  1.915000 0.545000 3.075000 ;
      RECT 0.525000  1.040000 0.705000 1.640000 ;
      RECT 0.525000  1.640000 1.425000 1.745000 ;
      RECT 0.715000  2.085000 1.045000 3.245000 ;
      RECT 0.885000  0.270000 1.215000 0.870000 ;
      RECT 0.885000  0.870000 2.165000 1.040000 ;
      RECT 1.215000  1.915000 1.425000 2.290000 ;
      RECT 1.215000  2.290000 2.660000 2.460000 ;
      RECT 1.215000  2.460000 1.615000 3.075000 ;
      RECT 1.405000  0.085000 1.735000 0.700000 ;
      RECT 1.905000  0.270000 2.165000 0.870000 ;
      RECT 2.195000  2.630000 2.865000 3.245000 ;
      RECT 2.335000  0.085000 2.565000 1.040000 ;
      RECT 2.490000  1.295000 2.860000 1.625000 ;
      RECT 2.490000  1.625000 2.660000 2.290000 ;
      RECT 3.235000  0.085000 3.620000 0.785000 ;
      RECT 3.370000  0.785000 3.620000 1.055000 ;
      RECT 3.395000  2.290000 3.725000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__o211a_2
END LIBRARY
