# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__fa_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__fa_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.636000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.260000 1.405000 0.695000 1.930000 ;
        RECT 0.260000 1.930000 1.670000 2.010000 ;
        RECT 0.525000 2.010000 1.670000 2.100000 ;
        RECT 1.500000 2.100000 1.670000 2.895000 ;
        RECT 1.500000 2.895000 2.465000 3.075000 ;
        RECT 2.295000 1.265000 2.530000 1.385000 ;
        RECT 2.295000 1.385000 3.990000 1.745000 ;
        RECT 2.295000 1.745000 4.995000 1.915000 ;
        RECT 2.295000 1.915000 2.465000 2.895000 ;
        RECT 4.825000 1.345000 5.720000 1.675000 ;
        RECT 4.825000 1.675000 4.995000 1.745000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.636000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.875000 1.550000 1.775000 1.755000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.075000 0.265000 2.245000 0.640000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.950000 0.255000 8.140000 0.840000 ;
        RECT 7.950000 0.840000 9.510000 1.010000 ;
        RECT 7.950000 1.755000 9.510000 1.925000 ;
        RECT 7.950000 1.925000 8.140000 3.075000 ;
        RECT 8.810000 0.255000 9.000000 0.840000 ;
        RECT 8.810000 1.925000 9.000000 3.075000 ;
        RECT 9.265000 1.010000 9.510000 1.755000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.230000 0.255000 6.420000 1.045000 ;
        RECT 6.230000 1.045000 7.575000 1.225000 ;
        RECT 6.230000 1.735000 7.575000 1.925000 ;
        RECT 6.230000 1.925000 6.420000 3.075000 ;
        RECT 7.090000 0.255000 7.280000 1.045000 ;
        RECT 7.090000 1.925000 7.280000 3.075000 ;
        RECT 7.215000 1.225000 7.575000 1.735000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.095000  2.180000 0.355000 2.280000 ;
      RECT 0.095000  2.280000 1.320000 2.450000 ;
      RECT 0.095000  2.450000 0.345000 2.850000 ;
      RECT 0.205000  0.705000 0.405000 1.065000 ;
      RECT 0.205000  1.065000 1.415000 1.235000 ;
      RECT 0.525000  2.620000 0.855000 3.245000 ;
      RECT 0.575000  0.085000 0.905000 0.885000 ;
      RECT 1.085000  0.810000 1.415000 1.065000 ;
      RECT 1.110000  2.450000 1.320000 2.610000 ;
      RECT 1.595000  0.810000 1.945000 1.210000 ;
      RECT 1.595000  1.210000 2.115000 1.380000 ;
      RECT 1.840000  2.055000 2.115000 2.725000 ;
      RECT 1.945000  1.380000 2.115000 2.055000 ;
      RECT 2.425000  0.085000 2.755000 1.040000 ;
      RECT 2.635000  2.105000 2.855000 3.245000 ;
      RECT 3.025000  2.095000 4.260000 2.265000 ;
      RECT 3.025000  2.265000 3.275000 2.765000 ;
      RECT 3.055000  0.765000 3.265000 1.045000 ;
      RECT 3.055000  1.045000 4.235000 1.215000 ;
      RECT 3.445000  0.085000 3.775000 0.865000 ;
      RECT 3.480000  2.435000 3.810000 3.245000 ;
      RECT 3.980000  2.265000 4.260000 2.765000 ;
      RECT 4.025000  0.765000 4.235000 1.045000 ;
      RECT 4.200000  1.385000 4.655000 1.575000 ;
      RECT 4.430000  2.095000 6.060000 2.265000 ;
      RECT 4.430000  2.265000 4.745000 2.765000 ;
      RECT 4.475000  1.200000 4.655000 1.385000 ;
      RECT 4.495000  0.700000 6.060000 1.030000 ;
      RECT 5.710000  0.085000 6.040000 0.530000 ;
      RECT 5.730000  2.435000 6.060000 3.245000 ;
      RECT 5.890000  1.030000 6.060000 1.395000 ;
      RECT 5.890000  1.395000 7.045000 1.565000 ;
      RECT 5.890000  1.565000 6.060000 2.095000 ;
      RECT 6.590000  0.085000 6.920000 0.875000 ;
      RECT 6.590000  2.105000 6.920000 3.245000 ;
      RECT 7.450000  0.085000 7.780000 0.875000 ;
      RECT 7.450000  2.105000 7.780000 3.245000 ;
      RECT 7.745000  1.180000 9.095000 1.515000 ;
      RECT 8.310000  0.085000 8.640000 0.670000 ;
      RECT 8.310000  2.105000 8.640000 3.245000 ;
      RECT 9.170000  0.085000 9.500000 0.670000 ;
      RECT 9.170000  2.105000 9.500000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  1.210000 4.645000 1.380000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  1.210000 8.005000 1.380000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
    LAYER met1 ;
      RECT 1.535000 1.180000 1.825000 1.225000 ;
      RECT 1.535000 1.225000 8.065000 1.365000 ;
      RECT 1.535000 1.365000 1.825000 1.410000 ;
      RECT 4.415000 1.180000 4.705000 1.225000 ;
      RECT 4.415000 1.365000 4.705000 1.410000 ;
      RECT 7.775000 1.180000 8.065000 1.225000 ;
      RECT 7.775000 1.365000 8.065000 1.410000 ;
  END
END sky130_fd_sc_lp__fa_4
END LIBRARY
