* File: sky130_fd_sc_lp__a2bb2oi_lp.pxi.spice
* Created: Wed Sep  2 09:24:42 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%B1 N_B1_M1003_g N_B1_M1010_g B1 B1 N_B1_c_82_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_LP%B1
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%B2 N_B2_M1007_g N_B2_M1001_g B2 B2 B2
+ N_B2_c_110_n PM_SKY130_FD_SC_LP__A2BB2OI_LP%B2
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%A_296_146# N_A_296_146#_M1012_d
+ N_A_296_146#_M1008_d N_A_296_146#_c_144_n N_A_296_146#_c_158_n
+ N_A_296_146#_M1002_g N_A_296_146#_c_145_n N_A_296_146#_M1006_g
+ N_A_296_146#_c_146_n N_A_296_146#_c_147_n N_A_296_146#_c_148_n
+ N_A_296_146#_M1004_g N_A_296_146#_c_149_n N_A_296_146#_c_150_n
+ N_A_296_146#_c_151_n N_A_296_146#_c_152_n N_A_296_146#_c_153_n
+ N_A_296_146#_c_154_n N_A_296_146#_c_155_n N_A_296_146#_c_156_n
+ N_A_296_146#_c_168_p N_A_296_146#_c_157_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_LP%A_296_146#
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%A2_N N_A2_N_c_246_n N_A2_N_M1011_g
+ N_A2_N_M1008_g N_A2_N_c_248_n N_A2_N_M1012_g A2_N N_A2_N_c_250_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_LP%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%A1_N N_A1_N_M1005_g N_A1_N_c_294_n
+ N_A1_N_c_295_n N_A1_N_M1000_g N_A1_N_M1009_g N_A1_N_c_297_n N_A1_N_c_298_n
+ A1_N A1_N N_A1_N_c_300_n PM_SKY130_FD_SC_LP__A2BB2OI_LP%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%A_27_409# N_A_27_409#_M1003_s
+ N_A_27_409#_M1007_d N_A_27_409#_c_339_n N_A_27_409#_c_340_n
+ N_A_27_409#_c_341_n N_A_27_409#_c_342_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%VPWR N_VPWR_M1003_d N_VPWR_M1009_d
+ N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n VPWR N_VPWR_c_370_n
+ N_VPWR_c_371_n N_VPWR_c_366_n PM_SKY130_FD_SC_LP__A2BB2OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%Y N_Y_M1001_d N_Y_M1002_d N_Y_c_405_n
+ N_Y_c_406_n N_Y_c_409_n Y Y PM_SKY130_FD_SC_LP__A2BB2OI_LP%Y
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%A_456_339# N_A_456_339#_M1008_s
+ N_A_456_339#_M1009_s N_A_456_339#_c_454_n N_A_456_339#_c_455_n
+ N_A_456_339#_c_456_n N_A_456_339#_c_457_n N_A_456_339#_c_458_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_LP%A_456_339#
x_PM_SKY130_FD_SC_LP__A2BB2OI_LP%VGND N_VGND_M1010_s N_VGND_M1004_d
+ N_VGND_M1000_d N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n VGND
+ N_VGND_c_486_n N_VGND_c_487_n N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n
+ N_VGND_c_491_n N_VGND_c_492_n N_VGND_c_493_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_LP%VGND
cc_1 VNB N_B1_M1003_g 0.0447703f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_2 VNB N_B1_M1010_g 0.0246719f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.445
cc_3 VNB B1 0.0241347f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_4 VNB N_B1_c_82_n 0.0471191f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.975
cc_5 VNB N_B2_M1001_g 0.0539238f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.445
cc_6 VNB B2 0.0203127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B2_c_110_n 0.0216334f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.975
cc_8 VNB N_A_296_146#_c_144_n 0.0101466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_296_146#_c_145_n 0.0134068f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.975
cc_10 VNB N_A_296_146#_c_146_n 0.011638f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.975
cc_11 VNB N_A_296_146#_c_147_n 0.0150744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_296_146#_c_148_n 0.0136543f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.975
cc_13 VNB N_A_296_146#_c_149_n 0.00734276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_296_146#_c_150_n 0.00514495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_296_146#_c_151_n 0.0201264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_296_146#_c_152_n 0.0111006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_296_146#_c_153_n 7.81587e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_296_146#_c_154_n 0.00513625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_296_146#_c_155_n 0.0109461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_296_146#_c_156_n 0.0119867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_296_146#_c_157_n 0.0365812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_N_c_246_n 0.0138908f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.14
cc_23 VNB N_A2_N_M1008_g 0.0303939f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.445
cc_24 VNB N_A2_N_c_248_n 0.0142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB A2_N 0.0102919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_N_c_250_n 0.0399062f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.81
cc_27 VNB N_A1_N_M1005_g 0.0298311f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_28 VNB N_A1_N_c_294_n 0.0159748f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.81
cc_29 VNB N_A1_N_c_295_n 0.010519f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.445
cc_30 VNB N_A1_N_M1000_g 0.0466841f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_31 VNB N_A1_N_c_297_n 0.0154238f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.975
cc_32 VNB N_A1_N_c_298_n 0.00397041f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.81
cc_33 VNB A1_N 0.0392049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A1_N_c_300_n 0.0331233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_366_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_405_n 0.0162918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_406_n 0.00364697f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_38 VNB Y 0.0115211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_483_n 0.01772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_484_n 0.00436014f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.975
cc_41 VNB N_VGND_c_485_n 0.0228982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_486_n 0.014713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_487_n 0.0320375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_488_n 0.0343439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_489_n 0.014713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_490_n 0.244676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_491_n 0.00511011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_492_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_493_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_B1_M1003_g 0.050083f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_51 VPB N_B2_M1007_g 0.0318543f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_52 VPB B2 0.0123959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_B2_c_110_n 0.00931036f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.975
cc_54 VPB N_A_296_146#_c_158_n 0.0109417f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_296_146#_M1002_g 0.0347114f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_56 VPB N_A_296_146#_c_151_n 0.00241632f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_296_146#_c_153_n 0.0156301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A2_N_M1008_g 0.0339946f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.445
cc_59 VPB N_A1_N_M1009_g 0.0343561f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_60 VPB N_A1_N_c_298_n 0.0326668f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.81
cc_61 VPB A1_N 0.0101349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_27_409#_c_339_n 0.0368459f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_63 VPB N_A_27_409#_c_340_n 0.01035f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_64 VPB N_A_27_409#_c_341_n 0.0106495f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_65 VPB N_A_27_409#_c_342_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.81
cc_66 VPB N_VPWR_c_367_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_368_n 0.0111973f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_68 VPB N_VPWR_c_369_n 0.0480195f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_69 VPB N_VPWR_c_370_n 0.0717889f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_70 VPB N_VPWR_c_371_n 0.0239038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_366_n 0.072926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_Y_c_406_n 0.00290759f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_73 VPB N_Y_c_409_n 0.0156858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_456_339#_c_454_n 0.0171337f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_75 VPB N_A_456_339#_c_455_n 0.0221929f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_76 VPB N_A_456_339#_c_456_n 0.00507162f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_77 VPB N_A_456_339#_c_457_n 0.00246318f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.975
cc_78 VPB N_A_456_339#_c_458_n 0.0166591f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.81
cc_79 N_B1_M1003_g N_B2_M1007_g 0.0321211f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_80 N_B1_M1010_g N_B2_M1001_g 0.0458019f $X=0.775 $Y=0.445 $X2=0 $Y2=0
cc_81 B1 N_B2_M1001_g 0.00281036f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_82 N_B1_c_82_n N_B2_M1001_g 0.0155222f $X=0.545 $Y=0.975 $X2=0 $Y2=0
cc_83 N_B1_M1003_g B2 0.0264301f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_84 B1 B2 0.036521f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_85 N_B1_c_82_n B2 0.00292345f $X=0.545 $Y=0.975 $X2=0 $Y2=0
cc_86 N_B1_M1003_g N_B2_c_110_n 0.0181444f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_87 N_B1_M1003_g N_A_27_409#_c_339_n 0.0164265f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_88 N_B1_M1003_g N_A_27_409#_c_340_n 0.0180843f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_89 N_B1_M1003_g N_A_27_409#_c_341_n 0.00198183f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_90 N_B1_M1003_g N_A_27_409#_c_342_n 9.07377e-19 $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_91 N_B1_M1003_g N_VPWR_c_367_n 0.0181825f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_92 N_B1_M1003_g N_VPWR_c_371_n 0.00769046f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_93 N_B1_M1003_g N_VPWR_c_366_n 0.014085f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_94 B1 N_Y_c_405_n 0.00878947f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_95 N_B1_M1010_g Y 0.00145228f $X=0.775 $Y=0.445 $X2=0 $Y2=0
cc_96 N_B1_M1010_g N_VGND_c_483_n 0.0122416f $X=0.775 $Y=0.445 $X2=0 $Y2=0
cc_97 B1 N_VGND_c_483_n 0.0227569f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_98 N_B1_c_82_n N_VGND_c_483_n 0.00774273f $X=0.545 $Y=0.975 $X2=0 $Y2=0
cc_99 N_B1_M1010_g N_VGND_c_487_n 0.00486043f $X=0.775 $Y=0.445 $X2=0 $Y2=0
cc_100 N_B1_M1010_g N_VGND_c_490_n 0.00492742f $X=0.775 $Y=0.445 $X2=0 $Y2=0
cc_101 B1 N_VGND_c_490_n 0.0144431f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_102 N_B1_c_82_n N_VGND_c_490_n 0.00129259f $X=0.545 $Y=0.975 $X2=0 $Y2=0
cc_103 N_B2_M1007_g N_A_296_146#_c_158_n 0.0194371f $X=1.075 $Y=2.545 $X2=0
+ $Y2=0
cc_104 N_B2_M1001_g N_A_296_146#_c_145_n 0.0116714f $X=1.165 $Y=0.445 $X2=0
+ $Y2=0
cc_105 N_B2_M1001_g N_A_296_146#_c_149_n 0.0283127f $X=1.165 $Y=0.445 $X2=0
+ $Y2=0
cc_106 N_B2_c_110_n N_A_296_146#_c_150_n 0.0283127f $X=1.075 $Y=1.615 $X2=0
+ $Y2=0
cc_107 B2 N_A_296_146#_c_151_n 0.00207534f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_B2_M1007_g N_A_27_409#_c_339_n 9.07377e-19 $X=1.075 $Y=2.545 $X2=0
+ $Y2=0
cc_109 N_B2_M1007_g N_A_27_409#_c_340_n 0.0195681f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_110 B2 N_A_27_409#_c_340_n 0.0573679f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_B2_c_110_n N_A_27_409#_c_340_n 0.00194355f $X=1.075 $Y=1.615 $X2=0
+ $Y2=0
cc_112 B2 N_A_27_409#_c_341_n 0.0245844f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_113 N_B2_M1007_g N_A_27_409#_c_342_n 0.0162664f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_114 N_B2_M1007_g N_VPWR_c_367_n 0.0171432f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_115 N_B2_M1007_g N_VPWR_c_370_n 0.00769046f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_116 N_B2_M1007_g N_VPWR_c_366_n 0.0134474f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_117 N_B2_M1001_g N_Y_c_405_n 0.00479242f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_118 B2 N_Y_c_405_n 0.014222f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_119 B2 N_Y_c_406_n 0.0119684f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_120 N_B2_M1007_g N_Y_c_409_n 0.00107506f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_121 N_B2_M1001_g Y 0.0155719f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_122 N_B2_M1001_g N_VGND_c_483_n 0.00162891f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B2_M1001_g N_VGND_c_487_n 0.00359964f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_124 N_B2_M1001_g N_VGND_c_490_n 0.00536967f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_296_146#_c_148_n N_A2_N_c_246_n 0.00900085f $X=1.955 $Y=0.73
+ $X2=-0.19 $Y2=-0.245
cc_126 N_A_296_146#_c_168_p N_A2_N_c_246_n 8.98058e-19 $X=3.11 $Y=0.43 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_296_146#_c_152_n N_A2_N_M1008_g 0.01847f $X=2.79 $Y=1.37 $X2=0 $Y2=0
cc_128 N_A_296_146#_c_153_n N_A2_N_M1008_g 0.0324968f $X=2.955 $Y=1.84 $X2=0
+ $Y2=0
cc_129 N_A_296_146#_c_154_n N_A2_N_M1008_g 0.00371105f $X=3.11 $Y=1.285 $X2=0
+ $Y2=0
cc_130 N_A_296_146#_c_155_n N_A2_N_M1008_g 0.00109637f $X=2.01 $Y=1.29 $X2=0
+ $Y2=0
cc_131 N_A_296_146#_c_156_n N_A2_N_M1008_g 0.0037596f $X=2.992 $Y=1.37 $X2=0
+ $Y2=0
cc_132 N_A_296_146#_c_157_n N_A2_N_M1008_g 0.0108982f $X=2.01 $Y=1.2 $X2=0 $Y2=0
cc_133 N_A_296_146#_c_154_n N_A2_N_c_248_n 0.00270976f $X=3.11 $Y=1.285 $X2=0
+ $Y2=0
cc_134 N_A_296_146#_c_168_p N_A2_N_c_248_n 0.00586076f $X=3.11 $Y=0.43 $X2=0
+ $Y2=0
cc_135 N_A_296_146#_c_147_n A2_N 5.15974e-19 $X=1.88 $Y=0.805 $X2=0 $Y2=0
cc_136 N_A_296_146#_c_152_n A2_N 0.018915f $X=2.79 $Y=1.37 $X2=0 $Y2=0
cc_137 N_A_296_146#_c_154_n A2_N 0.0237223f $X=3.11 $Y=1.285 $X2=0 $Y2=0
cc_138 N_A_296_146#_c_156_n A2_N 0.0043291f $X=2.992 $Y=1.37 $X2=0 $Y2=0
cc_139 N_A_296_146#_c_168_p A2_N 0.00218802f $X=3.11 $Y=0.43 $X2=0 $Y2=0
cc_140 N_A_296_146#_c_147_n N_A2_N_c_250_n 0.00900085f $X=1.88 $Y=0.805 $X2=0
+ $Y2=0
cc_141 N_A_296_146#_c_152_n N_A2_N_c_250_n 0.00750785f $X=2.79 $Y=1.37 $X2=0
+ $Y2=0
cc_142 N_A_296_146#_c_154_n N_A2_N_c_250_n 0.00189998f $X=3.11 $Y=1.285 $X2=0
+ $Y2=0
cc_143 N_A_296_146#_c_156_n N_A2_N_c_250_n 7.61897e-19 $X=2.992 $Y=1.37 $X2=0
+ $Y2=0
cc_144 N_A_296_146#_c_154_n N_A1_N_M1005_g 0.0136714f $X=3.11 $Y=1.285 $X2=0
+ $Y2=0
cc_145 N_A_296_146#_c_168_p N_A1_N_M1005_g 0.00721986f $X=3.11 $Y=0.43 $X2=0
+ $Y2=0
cc_146 N_A_296_146#_c_154_n N_A1_N_c_295_n 0.00635144f $X=3.11 $Y=1.285 $X2=0
+ $Y2=0
cc_147 N_A_296_146#_c_154_n N_A1_N_M1000_g 0.00274269f $X=3.11 $Y=1.285 $X2=0
+ $Y2=0
cc_148 N_A_296_146#_c_168_p N_A1_N_M1000_g 9.83916e-19 $X=3.11 $Y=0.43 $X2=0
+ $Y2=0
cc_149 N_A_296_146#_c_153_n N_A1_N_M1009_g 0.00124092f $X=2.955 $Y=1.84 $X2=0
+ $Y2=0
cc_150 N_A_296_146#_c_153_n N_A1_N_c_298_n 0.00654303f $X=2.955 $Y=1.84 $X2=0
+ $Y2=0
cc_151 N_A_296_146#_c_153_n A1_N 0.0156747f $X=2.955 $Y=1.84 $X2=0 $Y2=0
cc_152 N_A_296_146#_c_154_n A1_N 0.00896332f $X=3.11 $Y=1.285 $X2=0 $Y2=0
cc_153 N_A_296_146#_c_156_n A1_N 0.0104612f $X=2.992 $Y=1.37 $X2=0 $Y2=0
cc_154 N_A_296_146#_c_153_n N_A1_N_c_300_n 0.0030844f $X=2.955 $Y=1.84 $X2=0
+ $Y2=0
cc_155 N_A_296_146#_c_154_n N_A1_N_c_300_n 2.30023e-19 $X=3.11 $Y=1.285 $X2=0
+ $Y2=0
cc_156 N_A_296_146#_c_156_n N_A1_N_c_300_n 0.00181882f $X=2.992 $Y=1.37 $X2=0
+ $Y2=0
cc_157 N_A_296_146#_M1002_g N_A_27_409#_c_340_n 0.00468091f $X=1.605 $Y=2.545
+ $X2=0 $Y2=0
cc_158 N_A_296_146#_M1002_g N_A_27_409#_c_342_n 0.0163245f $X=1.605 $Y=2.545
+ $X2=0 $Y2=0
cc_159 N_A_296_146#_M1002_g N_VPWR_c_367_n 8.59418e-19 $X=1.605 $Y=2.545 $X2=0
+ $Y2=0
cc_160 N_A_296_146#_M1002_g N_VPWR_c_370_n 0.00826654f $X=1.605 $Y=2.545 $X2=0
+ $Y2=0
cc_161 N_A_296_146#_M1002_g N_VPWR_c_366_n 0.0158042f $X=1.605 $Y=2.545 $X2=0
+ $Y2=0
cc_162 N_A_296_146#_c_144_n N_Y_c_405_n 0.00738118f $X=1.555 $Y=1.125 $X2=0
+ $Y2=0
cc_163 N_A_296_146#_c_145_n N_Y_c_405_n 0.00247249f $X=1.595 $Y=0.73 $X2=0 $Y2=0
cc_164 N_A_296_146#_c_146_n N_Y_c_405_n 0.00339705f $X=1.845 $Y=1.2 $X2=0 $Y2=0
cc_165 N_A_296_146#_c_148_n N_Y_c_405_n 3.59266e-19 $X=1.955 $Y=0.73 $X2=0 $Y2=0
cc_166 N_A_296_146#_c_149_n N_Y_c_405_n 0.00801054f $X=1.575 $Y=0.805 $X2=0
+ $Y2=0
cc_167 N_A_296_146#_c_150_n N_Y_c_405_n 0.00379508f $X=1.555 $Y=1.2 $X2=0 $Y2=0
cc_168 N_A_296_146#_c_151_n N_Y_c_405_n 0.0111246f $X=1.605 $Y=1.695 $X2=0 $Y2=0
cc_169 N_A_296_146#_c_155_n N_Y_c_405_n 0.0231899f $X=2.01 $Y=1.29 $X2=0 $Y2=0
cc_170 N_A_296_146#_c_157_n N_Y_c_405_n 9.63409e-19 $X=2.01 $Y=1.2 $X2=0 $Y2=0
cc_171 N_A_296_146#_c_158_n N_Y_c_406_n 0.0152611f $X=1.605 $Y=1.82 $X2=0 $Y2=0
cc_172 N_A_296_146#_c_146_n N_Y_c_406_n 0.00438503f $X=1.845 $Y=1.2 $X2=0 $Y2=0
cc_173 N_A_296_146#_c_151_n N_Y_c_406_n 0.002694f $X=1.605 $Y=1.695 $X2=0 $Y2=0
cc_174 N_A_296_146#_c_155_n N_Y_c_406_n 0.0136693f $X=2.01 $Y=1.29 $X2=0 $Y2=0
cc_175 N_A_296_146#_c_157_n N_Y_c_406_n 0.00131587f $X=2.01 $Y=1.2 $X2=0 $Y2=0
cc_176 N_A_296_146#_c_158_n N_Y_c_409_n 6.82003e-19 $X=1.605 $Y=1.82 $X2=0 $Y2=0
cc_177 N_A_296_146#_M1002_g N_Y_c_409_n 0.0265001f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_178 N_A_296_146#_c_145_n Y 0.0100082f $X=1.595 $Y=0.73 $X2=0 $Y2=0
cc_179 N_A_296_146#_c_146_n Y 0.00175965f $X=1.845 $Y=1.2 $X2=0 $Y2=0
cc_180 N_A_296_146#_c_147_n Y 0.00129665f $X=1.88 $Y=0.805 $X2=0 $Y2=0
cc_181 N_A_296_146#_c_148_n Y 0.00303749f $X=1.955 $Y=0.73 $X2=0 $Y2=0
cc_182 N_A_296_146#_c_149_n Y 0.00103017f $X=1.575 $Y=0.805 $X2=0 $Y2=0
cc_183 N_A_296_146#_c_158_n N_A_456_339#_c_454_n 0.00281234f $X=1.605 $Y=1.82
+ $X2=0 $Y2=0
cc_184 N_A_296_146#_c_152_n N_A_456_339#_c_454_n 0.0229029f $X=2.79 $Y=1.37
+ $X2=0 $Y2=0
cc_185 N_A_296_146#_c_153_n N_A_456_339#_c_454_n 0.0685263f $X=2.955 $Y=1.84
+ $X2=0 $Y2=0
cc_186 N_A_296_146#_c_153_n N_A_456_339#_c_455_n 0.0246854f $X=2.955 $Y=1.84
+ $X2=0 $Y2=0
cc_187 N_A_296_146#_M1002_g N_A_456_339#_c_456_n 3.91664e-19 $X=1.605 $Y=2.545
+ $X2=0 $Y2=0
cc_188 N_A_296_146#_c_153_n N_A_456_339#_c_458_n 0.0465187f $X=2.955 $Y=1.84
+ $X2=0 $Y2=0
cc_189 N_A_296_146#_c_145_n N_VGND_c_484_n 0.00163043f $X=1.595 $Y=0.73 $X2=0
+ $Y2=0
cc_190 N_A_296_146#_c_148_n N_VGND_c_484_n 0.0107871f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_191 N_A_296_146#_c_152_n N_VGND_c_484_n 0.00544038f $X=2.79 $Y=1.37 $X2=0
+ $Y2=0
cc_192 N_A_296_146#_c_155_n N_VGND_c_484_n 0.00675873f $X=2.01 $Y=1.29 $X2=0
+ $Y2=0
cc_193 N_A_296_146#_c_168_p N_VGND_c_484_n 0.0109367f $X=3.11 $Y=0.43 $X2=0
+ $Y2=0
cc_194 N_A_296_146#_c_157_n N_VGND_c_484_n 0.001012f $X=2.01 $Y=1.2 $X2=0 $Y2=0
cc_195 N_A_296_146#_c_154_n N_VGND_c_485_n 0.00286662f $X=3.11 $Y=1.285 $X2=0
+ $Y2=0
cc_196 N_A_296_146#_c_168_p N_VGND_c_485_n 0.0125419f $X=3.11 $Y=0.43 $X2=0
+ $Y2=0
cc_197 N_A_296_146#_c_145_n N_VGND_c_487_n 0.00359964f $X=1.595 $Y=0.73 $X2=0
+ $Y2=0
cc_198 N_A_296_146#_c_148_n N_VGND_c_487_n 0.00486043f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_199 N_A_296_146#_c_168_p N_VGND_c_488_n 0.0207374f $X=3.11 $Y=0.43 $X2=0
+ $Y2=0
cc_200 N_A_296_146#_M1012_d N_VGND_c_490_n 0.00223855f $X=2.83 $Y=0.235 $X2=0
+ $Y2=0
cc_201 N_A_296_146#_c_145_n N_VGND_c_490_n 0.0052401f $X=1.595 $Y=0.73 $X2=0
+ $Y2=0
cc_202 N_A_296_146#_c_148_n N_VGND_c_490_n 0.00814425f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_203 N_A_296_146#_c_168_p N_VGND_c_490_n 0.0141529f $X=3.11 $Y=0.43 $X2=0
+ $Y2=0
cc_204 N_A2_N_M1008_g N_A1_N_M1005_g 0.0061359f $X=2.69 $Y=2.195 $X2=0 $Y2=0
cc_205 N_A2_N_c_248_n N_A1_N_M1005_g 0.0110084f $X=2.755 $Y=0.735 $X2=0 $Y2=0
cc_206 A2_N N_A1_N_M1005_g 3.63641e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_207 N_A2_N_c_250_n N_A1_N_M1005_g 0.0179157f $X=2.69 $Y=0.92 $X2=0 $Y2=0
cc_208 N_A2_N_M1008_g A1_N 3.52984e-19 $X=2.69 $Y=2.195 $X2=0 $Y2=0
cc_209 N_A2_N_M1008_g N_A1_N_c_300_n 0.00556951f $X=2.69 $Y=2.195 $X2=0 $Y2=0
cc_210 N_A2_N_M1008_g N_VPWR_c_370_n 3.19122e-19 $X=2.69 $Y=2.195 $X2=0 $Y2=0
cc_211 N_A2_N_c_246_n N_Y_c_405_n 6.39726e-19 $X=2.395 $Y=0.735 $X2=0 $Y2=0
cc_212 N_A2_N_M1008_g N_Y_c_406_n 0.00140608f $X=2.69 $Y=2.195 $X2=0 $Y2=0
cc_213 N_A2_N_M1008_g N_Y_c_409_n 0.00203276f $X=2.69 $Y=2.195 $X2=0 $Y2=0
cc_214 N_A2_N_M1008_g N_A_456_339#_c_454_n 0.0269654f $X=2.69 $Y=2.195 $X2=0
+ $Y2=0
cc_215 N_A2_N_M1008_g N_A_456_339#_c_455_n 0.00999807f $X=2.69 $Y=2.195 $X2=0
+ $Y2=0
cc_216 N_A2_N_M1008_g N_A_456_339#_c_458_n 0.00418443f $X=2.69 $Y=2.195 $X2=0
+ $Y2=0
cc_217 N_A2_N_c_246_n N_VGND_c_484_n 0.0123438f $X=2.395 $Y=0.735 $X2=0 $Y2=0
cc_218 N_A2_N_c_248_n N_VGND_c_484_n 0.00253827f $X=2.755 $Y=0.735 $X2=0 $Y2=0
cc_219 N_A2_N_c_246_n N_VGND_c_488_n 0.00525069f $X=2.395 $Y=0.735 $X2=0 $Y2=0
cc_220 N_A2_N_c_248_n N_VGND_c_488_n 0.00547815f $X=2.755 $Y=0.735 $X2=0 $Y2=0
cc_221 N_A2_N_c_250_n N_VGND_c_488_n 6.06977e-19 $X=2.69 $Y=0.92 $X2=0 $Y2=0
cc_222 N_A2_N_c_246_n N_VGND_c_490_n 0.00876208f $X=2.395 $Y=0.735 $X2=0 $Y2=0
cc_223 N_A2_N_c_248_n N_VGND_c_490_n 0.00595696f $X=2.755 $Y=0.735 $X2=0 $Y2=0
cc_224 A2_N N_VGND_c_490_n 0.00978611f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_225 N_A2_N_c_250_n N_VGND_c_490_n 8.02422e-19 $X=2.69 $Y=0.92 $X2=0 $Y2=0
cc_226 N_A1_N_M1009_g N_VPWR_c_369_n 0.0249256f $X=3.78 $Y=2.545 $X2=0 $Y2=0
cc_227 A1_N N_VPWR_c_369_n 0.0225338f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A1_N_M1009_g N_VPWR_c_370_n 0.00767656f $X=3.78 $Y=2.545 $X2=0 $Y2=0
cc_229 N_A1_N_M1009_g N_VPWR_c_366_n 0.014306f $X=3.78 $Y=2.545 $X2=0 $Y2=0
cc_230 N_A1_N_M1009_g N_A_456_339#_c_457_n 0.00373023f $X=3.78 $Y=2.545 $X2=0
+ $Y2=0
cc_231 N_A1_N_M1009_g N_A_456_339#_c_458_n 0.0160196f $X=3.78 $Y=2.545 $X2=0
+ $Y2=0
cc_232 N_A1_N_c_298_n N_A_456_339#_c_458_n 0.00489149f $X=3.637 $Y=1.613 $X2=0
+ $Y2=0
cc_233 A1_N N_A_456_339#_c_458_n 0.0136403f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_234 N_A1_N_M1005_g N_VGND_c_485_n 0.00236318f $X=3.185 $Y=0.445 $X2=0 $Y2=0
cc_235 N_A1_N_M1000_g N_VGND_c_485_n 0.0140864f $X=3.545 $Y=0.445 $X2=0 $Y2=0
cc_236 N_A1_N_c_297_n N_VGND_c_485_n 0.00418063f $X=3.637 $Y=1.185 $X2=0 $Y2=0
cc_237 A1_N N_VGND_c_485_n 0.0148401f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_238 N_A1_N_M1005_g N_VGND_c_488_n 0.00457646f $X=3.185 $Y=0.445 $X2=0 $Y2=0
cc_239 N_A1_N_M1000_g N_VGND_c_488_n 0.00486043f $X=3.545 $Y=0.445 $X2=0 $Y2=0
cc_240 N_A1_N_M1005_g N_VGND_c_490_n 0.00756643f $X=3.185 $Y=0.445 $X2=0 $Y2=0
cc_241 N_A1_N_M1000_g N_VGND_c_490_n 0.00814425f $X=3.545 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A_27_409#_c_340_n N_VPWR_M1003_d 0.00180746f $X=1.175 $Y=2.07 $X2=-0.19
+ $Y2=1.655
cc_243 N_A_27_409#_c_339_n N_VPWR_c_367_n 0.0481002f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_244 N_A_27_409#_c_340_n N_VPWR_c_367_n 0.0163515f $X=1.175 $Y=2.07 $X2=0
+ $Y2=0
cc_245 N_A_27_409#_c_342_n N_VPWR_c_367_n 0.0481002f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_246 N_A_27_409#_c_342_n N_VPWR_c_370_n 0.021949f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_247 N_A_27_409#_c_339_n N_VPWR_c_371_n 0.0220321f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_248 N_A_27_409#_c_339_n N_VPWR_c_366_n 0.0125808f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_249 N_A_27_409#_c_342_n N_VPWR_c_366_n 0.0124703f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_250 N_A_27_409#_c_340_n N_Y_c_406_n 7.27426e-19 $X=1.175 $Y=2.07 $X2=0 $Y2=0
cc_251 N_A_27_409#_c_340_n N_Y_c_409_n 0.0119061f $X=1.175 $Y=2.07 $X2=0 $Y2=0
cc_252 N_A_27_409#_c_342_n N_Y_c_409_n 0.0599276f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_253 N_VPWR_c_370_n N_Y_c_409_n 0.0220321f $X=3.88 $Y=3.33 $X2=0 $Y2=0
cc_254 N_VPWR_c_366_n N_Y_c_409_n 0.0125808f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_255 N_VPWR_c_370_n N_A_456_339#_c_455_n 0.0460277f $X=3.88 $Y=3.33 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_366_n N_A_456_339#_c_455_n 0.0283953f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_370_n N_A_456_339#_c_456_n 0.0222501f $X=3.88 $Y=3.33 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_366_n N_A_456_339#_c_456_n 0.0127687f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_369_n N_A_456_339#_c_457_n 0.0119061f $X=4.045 $Y=2.19 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_370_n N_A_456_339#_c_457_n 0.0221635f $X=3.88 $Y=3.33 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_366_n N_A_456_339#_c_457_n 0.0126536f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_369_n N_A_456_339#_c_458_n 0.0572919f $X=4.045 $Y=2.19 $X2=0
+ $Y2=0
cc_263 N_Y_c_406_n N_A_456_339#_c_454_n 0.00920229f $X=1.87 $Y=1.805 $X2=0 $Y2=0
cc_264 N_Y_c_409_n N_A_456_339#_c_454_n 0.0745781f $X=1.87 $Y=2.19 $X2=0 $Y2=0
cc_265 N_Y_c_409_n N_A_456_339#_c_456_n 0.0123491f $X=1.87 $Y=2.19 $X2=0 $Y2=0
cc_266 Y N_VGND_c_484_n 0.0287576f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_267 Y N_VGND_c_487_n 0.0390692f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_268 N_Y_M1001_d N_VGND_c_490_n 0.00225465f $X=1.24 $Y=0.235 $X2=0 $Y2=0
cc_269 Y N_VGND_c_490_n 0.0257113f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_270 Y A_334_47# 0.00427107f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_271 N_VGND_c_490_n A_170_47# 0.0101051f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_272 N_VGND_c_490_n A_334_47# 0.00464702f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_273 N_VGND_c_490_n A_494_47# 0.00418789f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_274 N_VGND_c_490_n A_652_47# 0.00899413f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
