# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o221a_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o221a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.955000 1.185000 3.225000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.185000 2.775000 1.515000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 1.210000 1.385000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.195000 1.905000 1.525000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.325000 1.345000 ;
        RECT 0.085000 1.345000 0.565000 1.750000 ;
        RECT 0.085000 1.750000 0.325000 2.575000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.581700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.650000 0.255000 4.235000 1.015000 ;
        RECT 3.655000 2.025000 4.235000 3.075000 ;
        RECT 3.735000 1.695000 4.235000 2.025000 ;
        RECT 3.925000 1.015000 4.235000 1.695000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.495000  0.255000 0.730000 1.005000 ;
      RECT 0.495000  1.005000 0.935000 1.175000 ;
      RECT 0.495000  1.930000 2.630000 2.100000 ;
      RECT 0.495000  2.100000 0.755000 3.075000 ;
      RECT 0.765000  1.175000 0.935000 1.930000 ;
      RECT 0.900000  0.255000 2.100000 0.425000 ;
      RECT 0.900000  0.425000 1.230000 0.835000 ;
      RECT 0.925000  2.270000 1.255000 3.245000 ;
      RECT 1.400000  0.595000 1.600000 0.845000 ;
      RECT 1.400000  0.845000 2.980000 1.015000 ;
      RECT 1.770000  0.425000 2.100000 0.675000 ;
      RECT 1.800000  1.695000 3.565000 1.865000 ;
      RECT 1.800000  1.865000 2.630000 1.930000 ;
      RECT 1.800000  2.100000 2.630000 3.075000 ;
      RECT 2.290000  0.085000 2.620000 0.675000 ;
      RECT 2.790000  0.255000 2.980000 0.845000 ;
      RECT 3.140000  2.035000 3.470000 3.245000 ;
      RECT 3.150000  0.085000 3.480000 1.015000 ;
      RECT 3.395000  1.185000 3.755000 1.515000 ;
      RECT 3.395000  1.515000 3.565000 1.695000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__o221a_1
