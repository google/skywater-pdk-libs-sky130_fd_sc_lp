* File: sky130_fd_sc_lp__o31a_m.pex.spice
* Created: Fri Aug 28 11:16:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31A_M%A1 3 7 11 12 13 14 18
c38 11 0 1.4009e-19 $X=1.03 $Y=1.66
c39 7 0 4.4852e-21 $X=1.12 $Y=2.195
c40 3 0 1.19165e-19 $X=1.12 $Y=0.445
r41 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.03
+ $Y=1.32 $X2=1.03 $Y2=1.32
r42 14 19 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=1.115 $Y=1.665
+ $X2=1.115 $Y2=1.32
r43 13 19 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=1.115 $Y=1.295
+ $X2=1.115 $Y2=1.32
r44 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.03 $Y=1.66
+ $X2=1.03 $Y2=1.32
r45 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.66
+ $X2=1.03 $Y2=1.825
r46 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.155
+ $X2=1.03 $Y2=1.32
r47 7 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.12 $Y=2.195
+ $X2=1.12 $Y2=1.825
r48 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.12 $Y=0.445
+ $X2=1.12 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_M%A_95_153# 1 2 8 12 13 15 16 17 20 22 23 28 29
+ 30 33 35 41
r75 39 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.315 $Y=2.94
+ $X2=1.315 $Y2=2.85
r76 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.315
+ $Y=2.94 $X2=1.315 $Y2=2.94
r77 35 38 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.315 $Y=2.755
+ $X2=1.315 $Y2=2.94
r78 31 33 75.5933 $w=1.88e-07 $l=1.295e-06 $layer=LI1_cond $X=3.01 $Y=1.805
+ $X2=3.01 $Y2=0.51
r79 29 31 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.915 $Y=1.89
+ $X2=3.01 $Y2=1.805
r80 29 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.915 $Y=1.89
+ $X2=2.34 $Y2=1.89
r81 26 28 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=2.235 $Y=2.67
+ $X2=2.235 $Y2=2.26
r82 25 30 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.235 $Y=1.975
+ $X2=2.34 $Y2=1.89
r83 25 28 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.235 $Y=1.975
+ $X2=2.235 $Y2=2.26
r84 24 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=2.755
+ $X2=1.315 $Y2=2.755
r85 23 26 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.13 $Y=2.755
+ $X2=2.235 $Y2=2.67
r86 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.13 $Y=2.755
+ $X2=1.48 $Y2=2.755
r87 16 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=2.85
+ $X2=1.315 $Y2=2.85
r88 16 17 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.15 $Y=2.85
+ $X2=0.655 $Y2=2.85
r89 13 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.69 $Y=0.765
+ $X2=0.69 $Y2=0.84
r90 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.69 $Y=0.765
+ $X2=0.69 $Y2=0.445
r91 12 22 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=0.58 $Y=2.195
+ $X2=0.58 $Y2=1.155
r92 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.58 $Y=2.775
+ $X2=0.655 $Y2=2.85
r93 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.58 $Y=2.775
+ $X2=0.58 $Y2=2.195
r94 8 22 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.565 $Y=1.065
+ $X2=0.565 $Y2=1.155
r95 7 20 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.565 $Y=0.84
+ $X2=0.69 $Y2=0.84
r96 7 8 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.565 $Y=0.915
+ $X2=0.565 $Y2=1.065
r97 2 28 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.985 $X2=2.235 $Y2=2.26
r98 1 33 182 $w=1.7e-07 $l=4.83322e-07 $layer=licon1_NDIFF $count=1 $X=2.635
+ $Y=0.235 $X2=3 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_M%A2 3 7 11 12 13 14 15 16 22
c43 11 0 1.4009e-19 $X=1.57 $Y=1.66
c44 3 0 4.4852e-21 $X=1.48 $Y=2.195
r45 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.57
+ $Y=1.32 $X2=1.57 $Y2=1.32
r46 15 16 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.625 $Y=2.035
+ $X2=1.625 $Y2=2.405
r47 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.625 $Y=1.665
+ $X2=1.625 $Y2=2.035
r48 14 23 14.1997 $w=2.78e-07 $l=3.45e-07 $layer=LI1_cond $X=1.625 $Y=1.665
+ $X2=1.625 $Y2=1.32
r49 13 23 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=1.625 $Y=1.295
+ $X2=1.625 $Y2=1.32
r50 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.57 $Y=1.66
+ $X2=1.57 $Y2=1.32
r51 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.66
+ $X2=1.57 $Y2=1.825
r52 10 22 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.155
+ $X2=1.57 $Y2=1.32
r53 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.55 $Y=0.445
+ $X2=1.55 $Y2=1.155
r54 3 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.48 $Y=2.195
+ $X2=1.48 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_M%A3 3 7 11 12 13 16
r40 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.11 $Y=1.1
+ $X2=2.11 $Y2=1.1
r41 13 17 1.17263 $w=5.08e-07 $l=5e-08 $layer=LI1_cond $X=2.16 $Y=1.27 $X2=2.11
+ $Y2=1.27
r42 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.11 $Y=1.44
+ $X2=2.11 $Y2=1.1
r43 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.44
+ $X2=2.11 $Y2=1.605
r44 10 16 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=0.935
+ $X2=2.11 $Y2=1.1
r45 7 10 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.075 $Y=0.445
+ $X2=2.075 $Y2=0.935
r46 3 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.02 $Y=2.195
+ $X2=2.02 $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_M%B1 3 6 9 10 11 12 13 14 19
r37 13 14 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=0.925
+ $X2=2.645 $Y2=1.295
r38 13 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.65
+ $Y=0.93 $X2=2.65 $Y2=0.93
r39 12 13 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=0.555
+ $X2=2.645 $Y2=0.925
r40 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.65 $Y=1.27
+ $X2=2.65 $Y2=0.93
r41 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.27
+ $X2=2.65 $Y2=1.435
r42 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=0.765
+ $X2=2.65 $Y2=0.93
r43 6 11 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.56 $Y=2.195
+ $X2=2.56 $Y2=1.435
r44 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.56 $Y=0.445 $X2=2.56
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_M%X 1 2 9 11 16
r22 14 16 1.03042 $w=4.23e-07 $l=3.8e-08 $layer=LI1_cond $X=0.367 $Y=0.887
+ $X2=0.367 $Y2=0.925
r23 11 14 0.650791 $w=4.23e-07 $l=2.4e-08 $layer=LI1_cond $X=0.367 $Y=0.863
+ $X2=0.367 $Y2=0.887
r24 11 22 8.04877 $w=4.23e-07 $l=1.88e-07 $layer=LI1_cond $X=0.367 $Y=0.863
+ $X2=0.367 $Y2=0.675
r25 11 19 32.0515 $w=4.23e-07 $l=1.182e-06 $layer=LI1_cond $X=0.367 $Y=0.948
+ $X2=0.367 $Y2=2.13
r26 11 16 0.623675 $w=4.23e-07 $l=2.3e-08 $layer=LI1_cond $X=0.367 $Y=0.948
+ $X2=0.367 $Y2=0.925
r27 9 22 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.475 $Y=0.51
+ $X2=0.475 $Y2=0.675
r28 2 19 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.24
+ $Y=1.985 $X2=0.365 $Y2=2.13
r29 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.35
+ $Y=0.235 $X2=0.475 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_M%VPWR 1 2 9 13 16 17 18 24 30 31 34
c32 31 0 8.97039e-21 $X=3.12 $Y=3.33
r33 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.94 $Y=3.33
+ $X2=2.775 $Y2=3.33
r37 28 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.94 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r39 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=2.775 $Y2=3.33
r40 24 26 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 18 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 16 21 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.76 $Y=3.33 $X2=0.72
+ $Y2=3.33
r46 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.76 $Y=3.33
+ $X2=0.865 $Y2=3.33
r47 15 26 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.865 $Y2=3.33
r49 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=3.245
+ $X2=2.775 $Y2=3.33
r50 11 13 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=2.775 $Y=3.245
+ $X2=2.775 $Y2=2.26
r51 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=3.33
r52 7 9 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=2.26
r53 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.985 $X2=2.775 $Y2=2.26
r54 1 9 600 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=1.985 $X2=0.865 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_M%VGND 1 2 9 11 15 17 18 19 30 31 34
r49 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r51 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r52 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r53 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=1.785
+ $Y2=0
r54 25 27 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=2.16
+ $Y2=0
r55 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r56 19 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r57 19 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r58 19 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r59 17 22 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.8 $Y=0 $X2=0.72
+ $Y2=0
r60 17 18 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.8 $Y=0 $X2=0.905
+ $Y2=0
r61 13 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0
r62 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0.38
r63 12 18 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.905
+ $Y2=0
r64 11 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.785
+ $Y2=0
r65 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.01
+ $Y2=0
r66 7 18 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.905 $Y=0.085
+ $X2=0.905 $Y2=0
r67 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0.085
+ $X2=0.905 $Y2=0.38
r68 2 15 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.235 $X2=1.785 $Y2=0.38
r69 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.765
+ $Y=0.235 $X2=0.905 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_M%A_239_47# 1 2 9 11 12 15
c30 15 0 1.41827e-19 $X=2.29 $Y=0.51
c31 9 0 2.89257e-19 $X=1.335 $Y=0.51
r32 13 15 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.28 $Y=0.665
+ $X2=2.28 $Y2=0.51
r33 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.185 $Y=0.75
+ $X2=2.28 $Y2=0.665
r34 11 12 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.185 $Y=0.75
+ $X2=1.44 $Y2=0.75
r35 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.335 $Y=0.665
+ $X2=1.44 $Y2=0.75
r36 7 9 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.335 $Y=0.665
+ $X2=1.335 $Y2=0.51
r37 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.15
+ $Y=0.235 $X2=2.29 $Y2=0.51
r38 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.235 $X2=1.335 $Y2=0.51
.ends

