* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux4_m A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_345_126# a_59_463# a_431_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_647_463# a_59_463# a_688_126# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_1184_171# S1 a_345_126# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_59_463# S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_616_126# S0 a_688_126# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_774_126# A0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_688_126# S0 a_805_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_805_463# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_688_126# S1 a_1184_171# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1118_37# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_59_463# S0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND A1 a_616_126# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_273_126# a_59_463# a_345_126# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_688_126# a_59_463# a_774_126# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_431_463# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VPWR A1 a_647_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VGND A2 a_273_126# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1184_171# a_1118_37# a_345_126# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 VPWR a_1184_171# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_345_126# S0 a_453_126# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR A2 a_273_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_273_463# S0 a_345_126# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_1118_37# S1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_1184_171# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_688_126# a_1118_37# a_1184_171# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_453_126# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
