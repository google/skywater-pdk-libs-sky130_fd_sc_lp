* File: sky130_fd_sc_lp__dlxbp_1.pxi.spice
* Created: Wed Sep  2 09:48:04 2020
* 
x_PM_SKY130_FD_SC_LP__DLXBP_1%D N_D_M1021_g N_D_M1002_g N_D_c_152_n N_D_c_153_n
+ N_D_c_154_n D D N_D_c_156_n PM_SKY130_FD_SC_LP__DLXBP_1%D
x_PM_SKY130_FD_SC_LP__DLXBP_1%GATE N_GATE_M1020_g N_GATE_M1008_g N_GATE_c_188_n
+ N_GATE_c_189_n GATE GATE N_GATE_c_191_n PM_SKY130_FD_SC_LP__DLXBP_1%GATE
x_PM_SKY130_FD_SC_LP__DLXBP_1%A_215_62# N_A_215_62#_M1020_d N_A_215_62#_M1008_d
+ N_A_215_62#_c_232_n N_A_215_62#_c_245_n N_A_215_62#_M1010_g
+ N_A_215_62#_M1013_g N_A_215_62#_M1019_g N_A_215_62#_c_234_n
+ N_A_215_62#_M1015_g N_A_215_62#_c_247_n N_A_215_62#_c_236_n
+ N_A_215_62#_c_237_n N_A_215_62#_c_238_n N_A_215_62#_c_248_n
+ N_A_215_62#_c_239_n N_A_215_62#_c_240_n N_A_215_62#_c_249_n
+ N_A_215_62#_c_250_n N_A_215_62#_c_241_n N_A_215_62#_c_242_n
+ N_A_215_62#_c_243_n PM_SKY130_FD_SC_LP__DLXBP_1%A_215_62#
x_PM_SKY130_FD_SC_LP__DLXBP_1%A_46_62# N_A_46_62#_M1021_s N_A_46_62#_M1002_s
+ N_A_46_62#_M1005_g N_A_46_62#_M1007_g N_A_46_62#_c_361_n N_A_46_62#_c_362_n
+ N_A_46_62#_c_368_n N_A_46_62#_c_369_n N_A_46_62#_c_363_n N_A_46_62#_c_364_n
+ N_A_46_62#_c_371_n N_A_46_62#_c_365_n PM_SKY130_FD_SC_LP__DLXBP_1%A_46_62#
x_PM_SKY130_FD_SC_LP__DLXBP_1%A_367_491# N_A_367_491#_M1013_s
+ N_A_367_491#_M1010_s N_A_367_491#_M1003_g N_A_367_491#_M1011_g
+ N_A_367_491#_c_444_n N_A_367_491#_c_436_n N_A_367_491#_c_445_n
+ N_A_367_491#_c_446_n N_A_367_491#_c_437_n N_A_367_491#_c_438_n
+ N_A_367_491#_c_439_n N_A_367_491#_c_448_n N_A_367_491#_c_440_n
+ N_A_367_491#_c_441_n N_A_367_491#_c_442_n
+ PM_SKY130_FD_SC_LP__DLXBP_1%A_367_491#
x_PM_SKY130_FD_SC_LP__DLXBP_1%A_758_359# N_A_758_359#_M1018_d
+ N_A_758_359#_M1009_d N_A_758_359#_M1006_g N_A_758_359#_M1001_g
+ N_A_758_359#_c_541_n N_A_758_359#_c_542_n N_A_758_359#_M1004_g
+ N_A_758_359#_M1017_g N_A_758_359#_c_544_n N_A_758_359#_c_545_n
+ N_A_758_359#_M1016_g N_A_758_359#_M1012_g N_A_758_359#_c_560_n
+ N_A_758_359#_c_547_n N_A_758_359#_c_548_n N_A_758_359#_c_549_n
+ N_A_758_359#_c_576_p N_A_758_359#_c_550_n N_A_758_359#_c_562_n
+ N_A_758_359#_c_563_n N_A_758_359#_c_551_n N_A_758_359#_c_564_n
+ N_A_758_359#_c_552_n N_A_758_359#_c_553_n N_A_758_359#_c_554_n
+ N_A_758_359#_c_566_n N_A_758_359#_c_555_n N_A_758_359#_c_556_n
+ PM_SKY130_FD_SC_LP__DLXBP_1%A_758_359#
x_PM_SKY130_FD_SC_LP__DLXBP_1%A_608_491# N_A_608_491#_M1003_d
+ N_A_608_491#_M1019_d N_A_608_491#_c_669_n N_A_608_491#_M1018_g
+ N_A_608_491#_M1009_g N_A_608_491#_c_677_n N_A_608_491#_c_671_n
+ N_A_608_491#_c_672_n N_A_608_491#_c_673_n N_A_608_491#_c_674_n
+ N_A_608_491#_c_685_n N_A_608_491#_c_675_n
+ PM_SKY130_FD_SC_LP__DLXBP_1%A_608_491#
x_PM_SKY130_FD_SC_LP__DLXBP_1%A_1266_147# N_A_1266_147#_M1016_d
+ N_A_1266_147#_M1012_d N_A_1266_147#_M1014_g N_A_1266_147#_M1000_g
+ N_A_1266_147#_c_758_n N_A_1266_147#_c_764_n N_A_1266_147#_c_759_n
+ N_A_1266_147#_c_760_n N_A_1266_147#_c_761_n N_A_1266_147#_c_762_n
+ PM_SKY130_FD_SC_LP__DLXBP_1%A_1266_147#
x_PM_SKY130_FD_SC_LP__DLXBP_1%VPWR N_VPWR_M1002_d N_VPWR_M1010_d N_VPWR_M1006_d
+ N_VPWR_M1017_d N_VPWR_M1000_s N_VPWR_c_798_n N_VPWR_c_799_n N_VPWR_c_800_n
+ N_VPWR_c_801_n N_VPWR_c_802_n N_VPWR_c_803_n N_VPWR_c_804_n N_VPWR_c_805_n
+ N_VPWR_c_806_n N_VPWR_c_807_n VPWR N_VPWR_c_808_n N_VPWR_c_809_n
+ N_VPWR_c_810_n N_VPWR_c_811_n N_VPWR_c_797_n N_VPWR_c_813_n N_VPWR_c_814_n
+ N_VPWR_c_815_n PM_SKY130_FD_SC_LP__DLXBP_1%VPWR
x_PM_SKY130_FD_SC_LP__DLXBP_1%Q N_Q_M1004_s N_Q_M1017_s N_Q_c_902_n N_Q_c_903_n
+ N_Q_c_899_n Q Q Q PM_SKY130_FD_SC_LP__DLXBP_1%Q
x_PM_SKY130_FD_SC_LP__DLXBP_1%Q_N N_Q_N_M1014_d N_Q_N_M1000_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N PM_SKY130_FD_SC_LP__DLXBP_1%Q_N
x_PM_SKY130_FD_SC_LP__DLXBP_1%VGND N_VGND_M1021_d N_VGND_M1013_d N_VGND_M1001_d
+ N_VGND_M1004_d N_VGND_M1014_s N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n
+ N_VGND_c_952_n N_VGND_c_953_n N_VGND_c_954_n VGND N_VGND_c_955_n
+ N_VGND_c_956_n N_VGND_c_957_n N_VGND_c_958_n N_VGND_c_959_n N_VGND_c_960_n
+ N_VGND_c_961_n N_VGND_c_962_n N_VGND_c_963_n N_VGND_c_964_n
+ PM_SKY130_FD_SC_LP__DLXBP_1%VGND
cc_1 VNB N_D_M1002_g 0.00850434f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.415
cc_2 VNB N_D_c_152_n 0.0208589f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.84
cc_3 VNB N_D_c_153_n 0.0241894f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.345
cc_4 VNB N_D_c_154_n 0.0168165f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.51
cc_5 VNB D 0.0102277f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_D_c_156_n 0.0162693f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.005
cc_7 VNB N_GATE_M1020_g 0.0205852f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.52
cc_8 VNB N_GATE_M1008_g 0.0430587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_GATE_c_188_n 0.037184f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.84
cc_10 VNB N_GATE_c_189_n 0.0086593f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.51
cc_11 VNB GATE 0.00752784f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_GATE_c_191_n 0.0501923f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.005
cc_13 VNB N_A_215_62#_c_232_n 0.0176921f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.005
cc_14 VNB N_A_215_62#_M1013_g 0.0376638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_215_62#_c_234_n 0.0338755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_215_62#_M1015_g 0.0420153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_215_62#_c_236_n 0.00732178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_215_62#_c_237_n 0.019929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_215_62#_c_238_n 0.00234259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_215_62#_c_239_n 0.0093079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_215_62#_c_240_n 0.00285548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_215_62#_c_241_n 0.00340212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_215_62#_c_242_n 0.037061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_215_62#_c_243_n 0.0243771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_46_62#_M1007_g 0.0262004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_46_62#_c_361_n 0.0184625f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.925
cc_27 VNB N_A_46_62#_c_362_n 0.048313f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.005
cc_28 VNB N_A_46_62#_c_363_n 0.00424113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_46_62#_c_364_n 0.0159209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_46_62#_c_365_n 0.0283234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_367_491#_c_436_n 0.00145986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_367_491#_c_437_n 0.0136573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_367_491#_c_438_n 0.0026958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_367_491#_c_439_n 0.00545343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_367_491#_c_440_n 0.00936464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_367_491#_c_441_n 0.0289969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_367_491#_c_442_n 0.0166696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_758_359#_M1001_g 0.0421698f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_39 VNB N_A_758_359#_c_541_n 0.0179599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_758_359#_c_542_n 0.0219857f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.005
cc_41 VNB N_A_758_359#_M1017_g 0.012771f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.005
cc_42 VNB N_A_758_359#_c_544_n 0.0152478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_758_359#_c_545_n 0.0205592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_758_359#_M1012_g 0.0140507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_758_359#_c_547_n 0.0159452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_758_359#_c_548_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_758_359#_c_549_n 0.00616293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_758_359#_c_550_n 0.0117115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_758_359#_c_551_n 0.00925875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_758_359#_c_552_n 0.00485812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_758_359#_c_553_n 3.68315e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_758_359#_c_554_n 0.00278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_758_359#_c_555_n 0.00302413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_758_359#_c_556_n 0.036322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_608_491#_c_669_n 0.0199456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_608_491#_M1009_g 0.00442157f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_57 VNB N_A_608_491#_c_671_n 0.00127317f $X=-0.19 $Y=-0.245 $X2=0.685
+ $Y2=0.925
cc_58 VNB N_A_608_491#_c_672_n 0.00427391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_608_491#_c_673_n 0.0180662f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.005
cc_60 VNB N_A_608_491#_c_674_n 0.00572135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_608_491#_c_675_n 0.0336557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1266_147#_c_758_n 0.00737849f $X=-0.19 $Y=-0.245 $X2=0.55
+ $Y2=1.005
cc_63 VNB N_A_1266_147#_c_759_n 0.00883085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1266_147#_c_760_n 0.0317205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1266_147#_c_761_n 0.00143323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1266_147#_c_762_n 0.0224572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VPWR_c_797_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_Q_c_899_n 0.00285973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB Q 0.00945817f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.005
cc_70 VNB Q 0.00205349f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.005
cc_71 VNB Q_N 0.0576438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_949_n 0.00737862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_950_n 0.00561515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_951_n 0.0369381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_952_n 0.00174825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_953_n 0.0264308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_954_n 0.026597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_955_n 0.0385009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_956_n 0.03375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_957_n 0.0218935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_958_n 0.0168564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_959_n 0.423821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_960_n 0.0248257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_961_n 0.00632057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_962_n 0.00632549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_963_n 0.0057671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_964_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VPB N_D_M1002_g 0.0398397f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.415
cc_89 VPB N_GATE_M1008_g 0.0437122f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_215_62#_c_232_n 0.0364514f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.005
cc_91 VPB N_A_215_62#_c_245_n 0.020279f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.84
cc_92 VPB N_A_215_62#_M1019_g 0.0508034f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.005
cc_93 VPB N_A_215_62#_c_247_n 0.0170526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_215_62#_c_248_n 0.0329967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_215_62#_c_249_n 0.00287832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_215_62#_c_250_n 0.0136652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_215_62#_c_243_n 0.00996597f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_46_62#_M1005_g 0.0325242f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.51
cc_99 VPB N_A_46_62#_c_362_n 0.00258945f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.005
cc_100 VPB N_A_46_62#_c_368_n 0.0387151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_46_62#_c_369_n 0.0297393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_46_62#_c_363_n 0.0284195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_46_62#_c_371_n 0.0229864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_367_491#_M1011_g 0.0177426f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_105 VPB N_A_367_491#_c_444_n 0.0121322f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.005
cc_106 VPB N_A_367_491#_c_445_n 0.00934705f $X=-0.19 $Y=1.655 $X2=0.685
+ $Y2=1.005
cc_107 VPB N_A_367_491#_c_446_n 0.00450583f $X=-0.19 $Y=1.655 $X2=0.685
+ $Y2=1.295
cc_108 VPB N_A_367_491#_c_439_n 0.00600393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_367_491#_c_448_n 0.0344897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_758_359#_M1006_g 0.0375756f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.84
cc_111 VPB N_A_758_359#_M1017_g 0.0277025f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.005
cc_112 VPB N_A_758_359#_M1012_g 0.0254364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_758_359#_c_560_n 0.0358306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_758_359#_c_550_n 0.0164042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_758_359#_c_562_n 0.00421638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_758_359#_c_563_n 0.00241736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_758_359#_c_564_n 0.0120809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_758_359#_c_553_n 0.0037348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_758_359#_c_566_n 0.00277697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_758_359#_c_556_n 0.00988353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_608_491#_M1009_g 0.025854f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_122 VPB N_A_608_491#_c_677_n 0.00457101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_608_491#_c_672_n 0.00602291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_1266_147#_M1000_g 0.0254717f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_125 VPB N_A_1266_147#_c_764_n 0.0151316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_1266_147#_c_759_n 0.00787623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_1266_147#_c_760_n 0.00710996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_798_n 0.0299211f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.005
cc_129 VPB N_VPWR_c_799_n 0.00239898f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.005
cc_130 VPB N_VPWR_c_800_n 0.00947986f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_801_n 0.0111958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_802_n 0.0302483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_803_n 0.029411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_804_n 0.0237449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_805_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_806_n 0.0363161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_807_n 0.00375746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_808_n 0.0358678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_809_n 0.02905f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_810_n 0.0218935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_811_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_797_n 0.117952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_813_n 0.0128726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_814_n 0.00574121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_815_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_Q_c_902_n 0.00335953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_Q_c_903_n 0.0102055f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.84
cc_148 VPB N_Q_c_899_n 0.00106921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB Q_N 0.057609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 N_D_c_152_n N_GATE_M1020_g 0.0114982f $X=0.55 $Y=0.84 $X2=0 $Y2=0
cc_151 D N_GATE_M1020_g 0.00148992f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_152 N_D_c_156_n N_GATE_M1020_g 0.00545117f $X=0.55 $Y=1.005 $X2=0 $Y2=0
cc_153 N_D_c_153_n N_GATE_M1008_g 0.0518804f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_154 D N_GATE_M1008_g 0.00364773f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_155 N_D_c_153_n N_GATE_c_189_n 0.00545117f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_156 D N_A_215_62#_c_236_n 0.0357121f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_157 N_D_c_156_n N_A_215_62#_c_236_n 3.23173e-19 $X=0.55 $Y=1.005 $X2=0 $Y2=0
cc_158 D N_A_215_62#_c_238_n 0.0193628f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_159 N_D_M1002_g N_A_46_62#_c_362_n 0.00601841f $X=0.64 $Y=2.415 $X2=0 $Y2=0
cc_160 N_D_c_152_n N_A_46_62#_c_362_n 0.00518096f $X=0.55 $Y=0.84 $X2=0 $Y2=0
cc_161 D N_A_46_62#_c_362_n 0.0522122f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_162 N_D_c_156_n N_A_46_62#_c_362_n 0.0163384f $X=0.55 $Y=1.005 $X2=0 $Y2=0
cc_163 N_D_M1002_g N_A_46_62#_c_368_n 0.00832307f $X=0.64 $Y=2.415 $X2=0 $Y2=0
cc_164 N_D_M1002_g N_A_46_62#_c_369_n 0.0185053f $X=0.64 $Y=2.415 $X2=0 $Y2=0
cc_165 D N_A_46_62#_c_369_n 0.0264331f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_166 N_D_c_156_n N_A_46_62#_c_364_n 0.00275842f $X=0.55 $Y=1.005 $X2=0 $Y2=0
cc_167 N_D_c_154_n N_A_46_62#_c_371_n 0.00407845f $X=0.55 $Y=1.51 $X2=0 $Y2=0
cc_168 D N_A_46_62#_c_371_n 0.00794588f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_169 N_D_M1002_g N_VPWR_c_798_n 0.00332801f $X=0.64 $Y=2.415 $X2=0 $Y2=0
cc_170 N_D_M1002_g N_VPWR_c_804_n 0.00431487f $X=0.64 $Y=2.415 $X2=0 $Y2=0
cc_171 N_D_M1002_g N_VPWR_c_797_n 0.00477801f $X=0.64 $Y=2.415 $X2=0 $Y2=0
cc_172 N_D_c_152_n N_VGND_c_949_n 0.00322927f $X=0.55 $Y=0.84 $X2=0 $Y2=0
cc_173 D N_VGND_c_949_n 0.0185078f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_174 N_D_c_156_n N_VGND_c_949_n 2.98046e-19 $X=0.55 $Y=1.005 $X2=0 $Y2=0
cc_175 N_D_c_152_n N_VGND_c_959_n 0.00598694f $X=0.55 $Y=0.84 $X2=0 $Y2=0
cc_176 D N_VGND_c_959_n 0.00644658f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_177 N_D_c_152_n N_VGND_c_960_n 0.00512921f $X=0.55 $Y=0.84 $X2=0 $Y2=0
cc_178 GATE N_A_215_62#_M1013_g 0.00292554f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_179 N_GATE_c_191_n N_A_215_62#_M1013_g 0.0142814f $X=1.615 $Y=0.505 $X2=0
+ $Y2=0
cc_180 N_GATE_M1020_g N_A_215_62#_c_236_n 0.00337968f $X=1 $Y=0.52 $X2=0 $Y2=0
cc_181 N_GATE_M1008_g N_A_215_62#_c_236_n 0.00852229f $X=1.07 $Y=2.415 $X2=0
+ $Y2=0
cc_182 N_GATE_c_188_n N_A_215_62#_c_236_n 0.0143078f $X=1.45 $Y=0.935 $X2=0
+ $Y2=0
cc_183 N_GATE_c_189_n N_A_215_62#_c_236_n 0.00213406f $X=1.035 $Y=0.935 $X2=0
+ $Y2=0
cc_184 GATE N_A_215_62#_c_236_n 0.0570265f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_185 N_GATE_c_191_n N_A_215_62#_c_236_n 0.00441226f $X=1.615 $Y=0.505 $X2=0
+ $Y2=0
cc_186 N_GATE_c_188_n N_A_215_62#_c_237_n 0.00808348f $X=1.45 $Y=0.935 $X2=0
+ $Y2=0
cc_187 GATE N_A_215_62#_c_237_n 0.0210761f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_188 N_GATE_M1008_g N_A_215_62#_c_238_n 0.0102758f $X=1.07 $Y=2.415 $X2=0
+ $Y2=0
cc_189 N_GATE_M1008_g N_A_215_62#_c_250_n 9.52487e-19 $X=1.07 $Y=2.415 $X2=0
+ $Y2=0
cc_190 GATE N_A_215_62#_c_241_n 0.00194531f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_191 GATE N_A_215_62#_c_242_n 6.59416e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_192 N_GATE_M1008_g N_A_46_62#_c_369_n 0.0215043f $X=1.07 $Y=2.415 $X2=0 $Y2=0
cc_193 N_GATE_c_188_n N_A_46_62#_c_369_n 7.15406e-19 $X=1.45 $Y=0.935 $X2=0
+ $Y2=0
cc_194 N_GATE_c_189_n N_A_46_62#_c_369_n 0.00172094f $X=1.035 $Y=0.935 $X2=0
+ $Y2=0
cc_195 N_GATE_M1008_g N_A_367_491#_c_444_n 0.00281739f $X=1.07 $Y=2.415 $X2=0
+ $Y2=0
cc_196 GATE N_A_367_491#_c_436_n 0.0341602f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_197 N_GATE_c_191_n N_A_367_491#_c_436_n 0.00310317f $X=1.615 $Y=0.505 $X2=0
+ $Y2=0
cc_198 GATE N_A_367_491#_c_438_n 0.0140146f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_199 N_GATE_c_191_n N_A_367_491#_c_438_n 0.0014945f $X=1.615 $Y=0.505 $X2=0
+ $Y2=0
cc_200 N_GATE_M1008_g N_VPWR_c_798_n 0.00332767f $X=1.07 $Y=2.415 $X2=0 $Y2=0
cc_201 N_GATE_M1008_g N_VPWR_c_806_n 0.00431487f $X=1.07 $Y=2.415 $X2=0 $Y2=0
cc_202 N_GATE_M1008_g N_VPWR_c_797_n 0.00477801f $X=1.07 $Y=2.415 $X2=0 $Y2=0
cc_203 N_GATE_M1020_g N_VGND_c_949_n 0.00256592f $X=1 $Y=0.52 $X2=0 $Y2=0
cc_204 GATE N_VGND_c_949_n 0.0025549f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_205 N_GATE_M1020_g N_VGND_c_955_n 0.00512921f $X=1 $Y=0.52 $X2=0 $Y2=0
cc_206 GATE N_VGND_c_955_n 0.0174199f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_207 N_GATE_c_191_n N_VGND_c_955_n 0.00414766f $X=1.615 $Y=0.505 $X2=0 $Y2=0
cc_208 N_GATE_M1020_g N_VGND_c_959_n 0.0105675f $X=1 $Y=0.52 $X2=0 $Y2=0
cc_209 GATE N_VGND_c_959_n 0.00944728f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_210 N_GATE_c_191_n N_VGND_c_959_n 0.002949f $X=1.615 $Y=0.505 $X2=0 $Y2=0
cc_211 N_A_215_62#_c_232_n N_A_46_62#_M1005_g 0.00680994f $X=2.065 $Y=2.195
+ $X2=0 $Y2=0
cc_212 N_A_215_62#_c_247_n N_A_46_62#_M1005_g 0.0317737f $X=2.175 $Y=2.27 $X2=0
+ $Y2=0
cc_213 N_A_215_62#_c_248_n N_A_46_62#_M1005_g 0.0107034f $X=2.89 $Y=2.165 $X2=0
+ $Y2=0
cc_214 N_A_215_62#_M1013_g N_A_46_62#_M1007_g 0.0172805f $X=2.245 $Y=0.445 $X2=0
+ $Y2=0
cc_215 N_A_215_62#_M1013_g N_A_46_62#_c_361_n 0.0144739f $X=2.245 $Y=0.445 $X2=0
+ $Y2=0
cc_216 N_A_215_62#_c_239_n N_A_46_62#_c_361_n 0.00424753f $X=2.89 $Y=1.45 $X2=0
+ $Y2=0
cc_217 N_A_215_62#_c_241_n N_A_46_62#_c_361_n 0.00188813f $X=2.155 $Y=1.25 $X2=0
+ $Y2=0
cc_218 N_A_215_62#_c_232_n N_A_46_62#_c_369_n 0.013442f $X=2.065 $Y=2.195 $X2=0
+ $Y2=0
cc_219 N_A_215_62#_M1019_g N_A_46_62#_c_369_n 5.95211e-19 $X=2.965 $Y=2.775
+ $X2=0 $Y2=0
cc_220 N_A_215_62#_c_247_n N_A_46_62#_c_369_n 5.73331e-19 $X=2.175 $Y=2.27 $X2=0
+ $Y2=0
cc_221 N_A_215_62#_c_237_n N_A_46_62#_c_369_n 0.0494234f $X=1.99 $Y=1.41 $X2=0
+ $Y2=0
cc_222 N_A_215_62#_c_238_n N_A_46_62#_c_369_n 0.0229424f $X=1.36 $Y=1.41 $X2=0
+ $Y2=0
cc_223 N_A_215_62#_c_248_n N_A_46_62#_c_369_n 0.0910889f $X=2.89 $Y=2.165 $X2=0
+ $Y2=0
cc_224 N_A_215_62#_c_239_n N_A_46_62#_c_369_n 0.025611f $X=2.89 $Y=1.45 $X2=0
+ $Y2=0
cc_225 N_A_215_62#_c_249_n N_A_46_62#_c_369_n 0.0130725f $X=3.015 $Y=2.075 $X2=0
+ $Y2=0
cc_226 N_A_215_62#_c_250_n N_A_46_62#_c_369_n 0.0251948f $X=1.285 $Y=2.24 $X2=0
+ $Y2=0
cc_227 N_A_215_62#_c_241_n N_A_46_62#_c_369_n 0.0258803f $X=2.155 $Y=1.25 $X2=0
+ $Y2=0
cc_228 N_A_215_62#_c_242_n N_A_46_62#_c_369_n 9.33213e-19 $X=2.155 $Y=1.25 $X2=0
+ $Y2=0
cc_229 N_A_215_62#_c_232_n N_A_46_62#_c_363_n 0.0220528f $X=2.065 $Y=2.195 $X2=0
+ $Y2=0
cc_230 N_A_215_62#_M1019_g N_A_46_62#_c_363_n 0.0584054f $X=2.965 $Y=2.775 $X2=0
+ $Y2=0
cc_231 N_A_215_62#_c_248_n N_A_46_62#_c_363_n 0.00444267f $X=2.89 $Y=2.165 $X2=0
+ $Y2=0
cc_232 N_A_215_62#_c_239_n N_A_46_62#_c_363_n 0.00428061f $X=2.89 $Y=1.45 $X2=0
+ $Y2=0
cc_233 N_A_215_62#_c_249_n N_A_46_62#_c_363_n 0.00142742f $X=3.015 $Y=2.075
+ $X2=0 $Y2=0
cc_234 N_A_215_62#_c_232_n N_A_46_62#_c_365_n 0.00793463f $X=2.065 $Y=2.195
+ $X2=0 $Y2=0
cc_235 N_A_215_62#_c_239_n N_A_46_62#_c_365_n 0.0107395f $X=2.89 $Y=1.45 $X2=0
+ $Y2=0
cc_236 N_A_215_62#_c_249_n N_A_46_62#_c_365_n 0.00115807f $X=3.015 $Y=2.075
+ $X2=0 $Y2=0
cc_237 N_A_215_62#_c_242_n N_A_46_62#_c_365_n 0.0144739f $X=2.155 $Y=1.25 $X2=0
+ $Y2=0
cc_238 N_A_215_62#_c_243_n N_A_46_62#_c_365_n 0.0584054f $X=3.055 $Y=1.44 $X2=0
+ $Y2=0
cc_239 N_A_215_62#_M1019_g N_A_367_491#_M1011_g 0.0172636f $X=2.965 $Y=2.775
+ $X2=0 $Y2=0
cc_240 N_A_215_62#_c_245_n N_A_367_491#_c_444_n 0.006417f $X=2.175 $Y=2.345
+ $X2=0 $Y2=0
cc_241 N_A_215_62#_c_250_n N_A_367_491#_c_444_n 0.00807176f $X=1.285 $Y=2.24
+ $X2=0 $Y2=0
cc_242 N_A_215_62#_M1013_g N_A_367_491#_c_436_n 0.00242633f $X=2.245 $Y=0.445
+ $X2=0 $Y2=0
cc_243 N_A_215_62#_c_245_n N_A_367_491#_c_445_n 0.00879064f $X=2.175 $Y=2.345
+ $X2=0 $Y2=0
cc_244 N_A_215_62#_M1019_g N_A_367_491#_c_445_n 0.0118816f $X=2.965 $Y=2.775
+ $X2=0 $Y2=0
cc_245 N_A_215_62#_c_248_n N_A_367_491#_c_445_n 0.0755046f $X=2.89 $Y=2.165
+ $X2=0 $Y2=0
cc_246 N_A_215_62#_c_245_n N_A_367_491#_c_446_n 0.00132014f $X=2.175 $Y=2.345
+ $X2=0 $Y2=0
cc_247 N_A_215_62#_c_247_n N_A_367_491#_c_446_n 0.00332867f $X=2.175 $Y=2.27
+ $X2=0 $Y2=0
cc_248 N_A_215_62#_c_248_n N_A_367_491#_c_446_n 0.0272505f $X=2.89 $Y=2.165
+ $X2=0 $Y2=0
cc_249 N_A_215_62#_c_250_n N_A_367_491#_c_446_n 0.00912409f $X=1.285 $Y=2.24
+ $X2=0 $Y2=0
cc_250 N_A_215_62#_M1013_g N_A_367_491#_c_437_n 0.0126272f $X=2.245 $Y=0.445
+ $X2=0 $Y2=0
cc_251 N_A_215_62#_c_239_n N_A_367_491#_c_437_n 0.0207058f $X=2.89 $Y=1.45 $X2=0
+ $Y2=0
cc_252 N_A_215_62#_c_240_n N_A_367_491#_c_437_n 0.00611134f $X=3.015 $Y=1.535
+ $X2=0 $Y2=0
cc_253 N_A_215_62#_c_241_n N_A_367_491#_c_437_n 0.0136374f $X=2.155 $Y=1.25
+ $X2=0 $Y2=0
cc_254 N_A_215_62#_c_242_n N_A_367_491#_c_437_n 2.44079e-19 $X=2.155 $Y=1.25
+ $X2=0 $Y2=0
cc_255 N_A_215_62#_c_243_n N_A_367_491#_c_437_n 8.90601e-19 $X=3.055 $Y=1.44
+ $X2=0 $Y2=0
cc_256 N_A_215_62#_c_237_n N_A_367_491#_c_438_n 0.00226293f $X=1.99 $Y=1.41
+ $X2=0 $Y2=0
cc_257 N_A_215_62#_c_241_n N_A_367_491#_c_438_n 0.0123985f $X=2.155 $Y=1.25
+ $X2=0 $Y2=0
cc_258 N_A_215_62#_c_242_n N_A_367_491#_c_438_n 0.00111388f $X=2.155 $Y=1.25
+ $X2=0 $Y2=0
cc_259 N_A_215_62#_M1019_g N_A_367_491#_c_439_n 0.00456674f $X=2.965 $Y=2.775
+ $X2=0 $Y2=0
cc_260 N_A_215_62#_c_234_n N_A_367_491#_c_439_n 0.0134733f $X=3.59 $Y=1.44 $X2=0
+ $Y2=0
cc_261 N_A_215_62#_M1015_g N_A_367_491#_c_439_n 0.00382577f $X=3.665 $Y=0.445
+ $X2=0 $Y2=0
cc_262 N_A_215_62#_c_248_n N_A_367_491#_c_439_n 0.014677f $X=2.89 $Y=2.165 $X2=0
+ $Y2=0
cc_263 N_A_215_62#_c_240_n N_A_367_491#_c_439_n 0.0131727f $X=3.015 $Y=1.535
+ $X2=0 $Y2=0
cc_264 N_A_215_62#_c_249_n N_A_367_491#_c_439_n 0.041256f $X=3.015 $Y=2.075
+ $X2=0 $Y2=0
cc_265 N_A_215_62#_c_243_n N_A_367_491#_c_439_n 0.00445396f $X=3.055 $Y=1.44
+ $X2=0 $Y2=0
cc_266 N_A_215_62#_M1019_g N_A_367_491#_c_448_n 0.0204967f $X=2.965 $Y=2.775
+ $X2=0 $Y2=0
cc_267 N_A_215_62#_c_234_n N_A_367_491#_c_448_n 0.00934521f $X=3.59 $Y=1.44
+ $X2=0 $Y2=0
cc_268 N_A_215_62#_c_248_n N_A_367_491#_c_448_n 0.00124596f $X=2.89 $Y=2.165
+ $X2=0 $Y2=0
cc_269 N_A_215_62#_c_249_n N_A_367_491#_c_448_n 6.77238e-19 $X=3.015 $Y=2.075
+ $X2=0 $Y2=0
cc_270 N_A_215_62#_M1015_g N_A_367_491#_c_440_n 0.00313925f $X=3.665 $Y=0.445
+ $X2=0 $Y2=0
cc_271 N_A_215_62#_c_240_n N_A_367_491#_c_440_n 0.00742631f $X=3.015 $Y=1.535
+ $X2=0 $Y2=0
cc_272 N_A_215_62#_c_243_n N_A_367_491#_c_440_n 0.00455586f $X=3.055 $Y=1.44
+ $X2=0 $Y2=0
cc_273 N_A_215_62#_M1015_g N_A_367_491#_c_441_n 0.019659f $X=3.665 $Y=0.445
+ $X2=0 $Y2=0
cc_274 N_A_215_62#_c_243_n N_A_367_491#_c_441_n 0.0150774f $X=3.055 $Y=1.44
+ $X2=0 $Y2=0
cc_275 N_A_215_62#_M1015_g N_A_367_491#_c_442_n 0.0141906f $X=3.665 $Y=0.445
+ $X2=0 $Y2=0
cc_276 N_A_215_62#_M1015_g N_A_758_359#_M1001_g 0.0424425f $X=3.665 $Y=0.445
+ $X2=0 $Y2=0
cc_277 N_A_215_62#_c_234_n N_A_758_359#_c_547_n 0.0424425f $X=3.59 $Y=1.44 $X2=0
+ $Y2=0
cc_278 N_A_215_62#_M1019_g N_A_608_491#_c_677_n 0.00546259f $X=2.965 $Y=2.775
+ $X2=0 $Y2=0
cc_279 N_A_215_62#_M1015_g N_A_608_491#_c_671_n 0.00293759f $X=3.665 $Y=0.445
+ $X2=0 $Y2=0
cc_280 N_A_215_62#_c_234_n N_A_608_491#_c_672_n 0.0050591f $X=3.59 $Y=1.44 $X2=0
+ $Y2=0
cc_281 N_A_215_62#_M1015_g N_A_608_491#_c_672_n 0.00385884f $X=3.665 $Y=0.445
+ $X2=0 $Y2=0
cc_282 N_A_215_62#_c_234_n N_A_608_491#_c_674_n 0.00229393f $X=3.59 $Y=1.44
+ $X2=0 $Y2=0
cc_283 N_A_215_62#_M1015_g N_A_608_491#_c_674_n 0.0232764f $X=3.665 $Y=0.445
+ $X2=0 $Y2=0
cc_284 N_A_215_62#_M1015_g N_A_608_491#_c_685_n 0.003846f $X=3.665 $Y=0.445
+ $X2=0 $Y2=0
cc_285 N_A_215_62#_c_250_n N_VPWR_c_798_n 0.00319103f $X=1.285 $Y=2.24 $X2=0
+ $Y2=0
cc_286 N_A_215_62#_c_245_n N_VPWR_c_799_n 0.00289494f $X=2.175 $Y=2.345 $X2=0
+ $Y2=0
cc_287 N_A_215_62#_M1019_g N_VPWR_c_799_n 0.00206028f $X=2.965 $Y=2.775 $X2=0
+ $Y2=0
cc_288 N_A_215_62#_c_245_n N_VPWR_c_806_n 0.00427134f $X=2.175 $Y=2.345 $X2=0
+ $Y2=0
cc_289 N_A_215_62#_c_250_n N_VPWR_c_806_n 0.00675656f $X=1.285 $Y=2.24 $X2=0
+ $Y2=0
cc_290 N_A_215_62#_M1019_g N_VPWR_c_808_n 0.00425651f $X=2.965 $Y=2.775 $X2=0
+ $Y2=0
cc_291 N_A_215_62#_c_245_n N_VPWR_c_797_n 0.00715113f $X=2.175 $Y=2.345 $X2=0
+ $Y2=0
cc_292 N_A_215_62#_M1019_g N_VPWR_c_797_n 0.00735215f $X=2.965 $Y=2.775 $X2=0
+ $Y2=0
cc_293 N_A_215_62#_c_250_n N_VPWR_c_797_n 0.00929055f $X=1.285 $Y=2.24 $X2=0
+ $Y2=0
cc_294 N_A_215_62#_M1013_g N_VGND_c_950_n 0.00325355f $X=2.245 $Y=0.445 $X2=0
+ $Y2=0
cc_295 N_A_215_62#_M1015_g N_VGND_c_951_n 0.00402323f $X=3.665 $Y=0.445 $X2=0
+ $Y2=0
cc_296 N_A_215_62#_M1015_g N_VGND_c_952_n 0.00251916f $X=3.665 $Y=0.445 $X2=0
+ $Y2=0
cc_297 N_A_215_62#_M1013_g N_VGND_c_955_n 0.00440547f $X=2.245 $Y=0.445 $X2=0
+ $Y2=0
cc_298 N_A_215_62#_c_236_n N_VGND_c_955_n 0.0103069f $X=1.215 $Y=0.53 $X2=0
+ $Y2=0
cc_299 N_A_215_62#_M1013_g N_VGND_c_959_n 0.00763061f $X=2.245 $Y=0.445 $X2=0
+ $Y2=0
cc_300 N_A_215_62#_M1015_g N_VGND_c_959_n 0.00594764f $X=3.665 $Y=0.445 $X2=0
+ $Y2=0
cc_301 N_A_215_62#_c_236_n N_VGND_c_959_n 0.00999125f $X=1.215 $Y=0.53 $X2=0
+ $Y2=0
cc_302 N_A_46_62#_M1005_g N_A_367_491#_c_444_n 7.61432e-19 $X=2.605 $Y=2.775
+ $X2=0 $Y2=0
cc_303 N_A_46_62#_M1005_g N_A_367_491#_c_445_n 0.0114138f $X=2.605 $Y=2.775
+ $X2=0 $Y2=0
cc_304 N_A_46_62#_M1007_g N_A_367_491#_c_437_n 0.0128005f $X=2.765 $Y=0.445
+ $X2=0 $Y2=0
cc_305 N_A_46_62#_c_361_n N_A_367_491#_c_437_n 0.00530498f $X=2.765 $Y=1.05
+ $X2=0 $Y2=0
cc_306 N_A_46_62#_c_365_n N_A_367_491#_c_439_n 0.0039461f $X=2.515 $Y=1.655
+ $X2=0 $Y2=0
cc_307 N_A_46_62#_M1007_g N_A_367_491#_c_440_n 0.00125187f $X=2.765 $Y=0.445
+ $X2=0 $Y2=0
cc_308 N_A_46_62#_c_361_n N_A_367_491#_c_440_n 0.00120124f $X=2.765 $Y=1.05
+ $X2=0 $Y2=0
cc_309 N_A_46_62#_c_365_n N_A_367_491#_c_440_n 0.00186685f $X=2.515 $Y=1.655
+ $X2=0 $Y2=0
cc_310 N_A_46_62#_c_361_n N_A_367_491#_c_441_n 0.0308379f $X=2.765 $Y=1.05 $X2=0
+ $Y2=0
cc_311 N_A_46_62#_M1007_g N_A_367_491#_c_442_n 0.0308379f $X=2.765 $Y=0.445
+ $X2=0 $Y2=0
cc_312 N_A_46_62#_M1005_g N_A_608_491#_c_677_n 8.34593e-19 $X=2.605 $Y=2.775
+ $X2=0 $Y2=0
cc_313 N_A_46_62#_c_368_n N_VPWR_c_798_n 0.00307927f $X=0.425 $Y=2.24 $X2=0
+ $Y2=0
cc_314 N_A_46_62#_c_369_n N_VPWR_c_798_n 0.0220348f $X=2.515 $Y=1.82 $X2=0 $Y2=0
cc_315 N_A_46_62#_M1005_g N_VPWR_c_799_n 0.0100625f $X=2.605 $Y=2.775 $X2=0
+ $Y2=0
cc_316 N_A_46_62#_c_368_n N_VPWR_c_804_n 0.00675656f $X=0.425 $Y=2.24 $X2=0
+ $Y2=0
cc_317 N_A_46_62#_M1005_g N_VPWR_c_808_n 0.00365202f $X=2.605 $Y=2.775 $X2=0
+ $Y2=0
cc_318 N_A_46_62#_M1005_g N_VPWR_c_797_n 0.00423089f $X=2.605 $Y=2.775 $X2=0
+ $Y2=0
cc_319 N_A_46_62#_c_368_n N_VPWR_c_797_n 0.00929055f $X=0.425 $Y=2.24 $X2=0
+ $Y2=0
cc_320 N_A_46_62#_M1007_g N_VGND_c_950_n 0.00325355f $X=2.765 $Y=0.445 $X2=0
+ $Y2=0
cc_321 N_A_46_62#_M1007_g N_VGND_c_951_n 0.00440547f $X=2.765 $Y=0.445 $X2=0
+ $Y2=0
cc_322 N_A_46_62#_M1007_g N_VGND_c_959_n 0.006063f $X=2.765 $Y=0.445 $X2=0 $Y2=0
cc_323 N_A_46_62#_c_364_n N_VGND_c_959_n 0.0146949f $X=0.355 $Y=0.505 $X2=0
+ $Y2=0
cc_324 N_A_46_62#_c_364_n N_VGND_c_960_n 0.0165256f $X=0.355 $Y=0.505 $X2=0
+ $Y2=0
cc_325 N_A_367_491#_M1011_g N_A_758_359#_M1006_g 0.039312f $X=3.49 $Y=2.665
+ $X2=0 $Y2=0
cc_326 N_A_367_491#_c_439_n N_A_758_359#_c_560_n 0.00133632f $X=3.415 $Y=2.13
+ $X2=0 $Y2=0
cc_327 N_A_367_491#_c_448_n N_A_758_359#_c_560_n 0.0203356f $X=3.415 $Y=2.13
+ $X2=0 $Y2=0
cc_328 N_A_367_491#_c_445_n N_A_608_491#_M1019_d 0.00278247f $X=3.31 $Y=2.51
+ $X2=0 $Y2=0
cc_329 N_A_367_491#_M1011_g N_A_608_491#_c_677_n 0.0154127f $X=3.49 $Y=2.665
+ $X2=0 $Y2=0
cc_330 N_A_367_491#_c_445_n N_A_608_491#_c_677_n 0.0284078f $X=3.31 $Y=2.51
+ $X2=0 $Y2=0
cc_331 N_A_367_491#_c_448_n N_A_608_491#_c_677_n 4.20143e-19 $X=3.415 $Y=2.13
+ $X2=0 $Y2=0
cc_332 N_A_367_491#_c_440_n N_A_608_491#_c_671_n 0.00547421f $X=3.215 $Y=0.93
+ $X2=0 $Y2=0
cc_333 N_A_367_491#_c_441_n N_A_608_491#_c_671_n 4.44563e-19 $X=3.215 $Y=0.93
+ $X2=0 $Y2=0
cc_334 N_A_367_491#_M1011_g N_A_608_491#_c_672_n 0.00527879f $X=3.49 $Y=2.665
+ $X2=0 $Y2=0
cc_335 N_A_367_491#_c_445_n N_A_608_491#_c_672_n 0.0134011f $X=3.31 $Y=2.51
+ $X2=0 $Y2=0
cc_336 N_A_367_491#_c_439_n N_A_608_491#_c_672_n 0.0907965f $X=3.415 $Y=2.13
+ $X2=0 $Y2=0
cc_337 N_A_367_491#_c_448_n N_A_608_491#_c_672_n 0.00200461f $X=3.415 $Y=2.13
+ $X2=0 $Y2=0
cc_338 N_A_367_491#_c_440_n N_A_608_491#_c_672_n 0.00308645f $X=3.215 $Y=0.93
+ $X2=0 $Y2=0
cc_339 N_A_367_491#_c_440_n N_A_608_491#_c_674_n 0.0231207f $X=3.215 $Y=0.93
+ $X2=0 $Y2=0
cc_340 N_A_367_491#_c_441_n N_A_608_491#_c_674_n 0.00275195f $X=3.215 $Y=0.93
+ $X2=0 $Y2=0
cc_341 N_A_367_491#_c_442_n N_A_608_491#_c_674_n 0.00343889f $X=3.215 $Y=0.765
+ $X2=0 $Y2=0
cc_342 N_A_367_491#_c_440_n N_A_608_491#_c_685_n 0.012922f $X=3.215 $Y=0.93
+ $X2=0 $Y2=0
cc_343 N_A_367_491#_c_445_n N_VPWR_M1010_d 0.00172285f $X=3.31 $Y=2.51 $X2=0
+ $Y2=0
cc_344 N_A_367_491#_c_445_n N_VPWR_c_799_n 0.0147386f $X=3.31 $Y=2.51 $X2=0
+ $Y2=0
cc_345 N_A_367_491#_c_444_n N_VPWR_c_806_n 0.0209837f $X=1.96 $Y=2.6 $X2=0 $Y2=0
cc_346 N_A_367_491#_c_445_n N_VPWR_c_806_n 0.00196209f $X=3.31 $Y=2.51 $X2=0
+ $Y2=0
cc_347 N_A_367_491#_M1011_g N_VPWR_c_808_n 7.94855e-19 $X=3.49 $Y=2.665 $X2=0
+ $Y2=0
cc_348 N_A_367_491#_c_445_n N_VPWR_c_808_n 0.00547813f $X=3.31 $Y=2.51 $X2=0
+ $Y2=0
cc_349 N_A_367_491#_M1010_s N_VPWR_c_797_n 0.00215158f $X=1.835 $Y=2.455 $X2=0
+ $Y2=0
cc_350 N_A_367_491#_c_444_n N_VPWR_c_797_n 0.0125539f $X=1.96 $Y=2.6 $X2=0 $Y2=0
cc_351 N_A_367_491#_c_445_n N_VPWR_c_797_n 0.0162105f $X=3.31 $Y=2.51 $X2=0
+ $Y2=0
cc_352 N_A_367_491#_c_445_n A_536_491# 0.0018586f $X=3.31 $Y=2.51 $X2=-0.19
+ $Y2=-0.245
cc_353 N_A_367_491#_c_437_n N_VGND_c_950_n 0.0229757f $X=3.05 $Y=0.83 $X2=0
+ $Y2=0
cc_354 N_A_367_491#_c_437_n N_VGND_c_951_n 0.00527279f $X=3.05 $Y=0.83 $X2=0
+ $Y2=0
cc_355 N_A_367_491#_c_440_n N_VGND_c_951_n 0.00244865f $X=3.215 $Y=0.93 $X2=0
+ $Y2=0
cc_356 N_A_367_491#_c_442_n N_VGND_c_951_n 0.00440413f $X=3.215 $Y=0.765 $X2=0
+ $Y2=0
cc_357 N_A_367_491#_c_436_n N_VGND_c_955_n 0.0107122f $X=2.03 $Y=0.445 $X2=0
+ $Y2=0
cc_358 N_A_367_491#_c_437_n N_VGND_c_955_n 0.00271124f $X=3.05 $Y=0.83 $X2=0
+ $Y2=0
cc_359 N_A_367_491#_M1013_s N_VGND_c_959_n 0.00376679f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_360 N_A_367_491#_c_436_n N_VGND_c_959_n 0.00720611f $X=2.03 $Y=0.445 $X2=0
+ $Y2=0
cc_361 N_A_367_491#_c_437_n N_VGND_c_959_n 0.0149741f $X=3.05 $Y=0.83 $X2=0
+ $Y2=0
cc_362 N_A_367_491#_c_440_n N_VGND_c_959_n 0.00415557f $X=3.215 $Y=0.93 $X2=0
+ $Y2=0
cc_363 N_A_367_491#_c_442_n N_VGND_c_959_n 0.00631653f $X=3.215 $Y=0.765 $X2=0
+ $Y2=0
cc_364 N_A_758_359#_M1001_g N_A_608_491#_c_669_n 0.0215758f $X=4.025 $Y=0.445
+ $X2=0 $Y2=0
cc_365 N_A_758_359#_c_551_n N_A_608_491#_c_669_n 0.00663007f $X=4.815 $Y=0.42
+ $X2=0 $Y2=0
cc_366 N_A_758_359#_c_552_n N_A_608_491#_c_669_n 0.00289953f $X=5.02 $Y=1.265
+ $X2=0 $Y2=0
cc_367 N_A_758_359#_c_576_p N_A_608_491#_M1009_g 0.00130117f $X=4.115 $Y=1.48
+ $X2=0 $Y2=0
cc_368 N_A_758_359#_c_550_n N_A_608_491#_M1009_g 0.0123382f $X=4.115 $Y=1.48
+ $X2=0 $Y2=0
cc_369 N_A_758_359#_c_562_n N_A_608_491#_M1009_g 0.0159132f $X=4.9 $Y=1.86 $X2=0
+ $Y2=0
cc_370 N_A_758_359#_c_563_n N_A_608_491#_M1009_g 2.01271e-19 $X=4.21 $Y=1.86
+ $X2=0 $Y2=0
cc_371 N_A_758_359#_c_564_n N_A_608_491#_M1009_g 0.00373924f $X=4.995 $Y=2.89
+ $X2=0 $Y2=0
cc_372 N_A_758_359#_c_553_n N_A_608_491#_M1009_g 0.00698758f $X=5.047 $Y=1.775
+ $X2=0 $Y2=0
cc_373 N_A_758_359#_M1006_g N_A_608_491#_c_677_n 0.00638685f $X=3.865 $Y=2.665
+ $X2=0 $Y2=0
cc_374 N_A_758_359#_M1001_g N_A_608_491#_c_671_n 0.00299669f $X=4.025 $Y=0.445
+ $X2=0 $Y2=0
cc_375 N_A_758_359#_M1006_g N_A_608_491#_c_672_n 0.0200663f $X=3.865 $Y=2.665
+ $X2=0 $Y2=0
cc_376 N_A_758_359#_M1001_g N_A_608_491#_c_672_n 0.00967476f $X=4.025 $Y=0.445
+ $X2=0 $Y2=0
cc_377 N_A_758_359#_c_560_n N_A_608_491#_c_672_n 0.00802036f $X=4.035 $Y=1.985
+ $X2=0 $Y2=0
cc_378 N_A_758_359#_c_576_p N_A_608_491#_c_672_n 0.0330983f $X=4.115 $Y=1.48
+ $X2=0 $Y2=0
cc_379 N_A_758_359#_c_563_n N_A_608_491#_c_672_n 0.0157322f $X=4.21 $Y=1.86
+ $X2=0 $Y2=0
cc_380 N_A_758_359#_M1001_g N_A_608_491#_c_673_n 0.0177927f $X=4.025 $Y=0.445
+ $X2=0 $Y2=0
cc_381 N_A_758_359#_c_560_n N_A_608_491#_c_673_n 0.00247927f $X=4.035 $Y=1.985
+ $X2=0 $Y2=0
cc_382 N_A_758_359#_c_547_n N_A_608_491#_c_673_n 0.00715113f $X=4.115 $Y=1.44
+ $X2=0 $Y2=0
cc_383 N_A_758_359#_c_576_p N_A_608_491#_c_673_n 0.0301302f $X=4.115 $Y=1.48
+ $X2=0 $Y2=0
cc_384 N_A_758_359#_c_562_n N_A_608_491#_c_673_n 0.0242587f $X=4.9 $Y=1.86 $X2=0
+ $Y2=0
cc_385 N_A_758_359#_c_552_n N_A_608_491#_c_673_n 0.0133059f $X=5.02 $Y=1.265
+ $X2=0 $Y2=0
cc_386 N_A_758_359#_c_554_n N_A_608_491#_c_673_n 0.00519904f $X=4.912 $Y=1.005
+ $X2=0 $Y2=0
cc_387 N_A_758_359#_c_555_n N_A_608_491#_c_673_n 0.0194435f $X=5.23 $Y=1.43
+ $X2=0 $Y2=0
cc_388 N_A_758_359#_c_556_n N_A_608_491#_c_673_n 2.07344e-19 $X=5.23 $Y=1.34
+ $X2=0 $Y2=0
cc_389 N_A_758_359#_M1001_g N_A_608_491#_c_674_n 0.00284754f $X=4.025 $Y=0.445
+ $X2=0 $Y2=0
cc_390 N_A_758_359#_c_547_n N_A_608_491#_c_675_n 0.0135848f $X=4.115 $Y=1.44
+ $X2=0 $Y2=0
cc_391 N_A_758_359#_c_562_n N_A_608_491#_c_675_n 0.00112425f $X=4.9 $Y=1.86
+ $X2=0 $Y2=0
cc_392 N_A_758_359#_c_552_n N_A_608_491#_c_675_n 0.00202989f $X=5.02 $Y=1.265
+ $X2=0 $Y2=0
cc_393 N_A_758_359#_c_554_n N_A_608_491#_c_675_n 0.00505057f $X=4.912 $Y=1.005
+ $X2=0 $Y2=0
cc_394 N_A_758_359#_c_555_n N_A_608_491#_c_675_n 0.0038242f $X=5.23 $Y=1.43
+ $X2=0 $Y2=0
cc_395 N_A_758_359#_c_556_n N_A_608_491#_c_675_n 0.0202455f $X=5.23 $Y=1.34
+ $X2=0 $Y2=0
cc_396 N_A_758_359#_c_542_n N_A_1266_147#_c_758_n 3.76836e-19 $X=5.73 $Y=1.265
+ $X2=0 $Y2=0
cc_397 N_A_758_359#_c_545_n N_A_1266_147#_c_758_n 0.00860465f $X=6.255 $Y=1.265
+ $X2=0 $Y2=0
cc_398 N_A_758_359#_c_549_n N_A_1266_147#_c_758_n 0.00407259f $X=6.255 $Y=1.34
+ $X2=0 $Y2=0
cc_399 N_A_758_359#_M1017_g N_A_1266_147#_c_764_n 5.85795e-19 $X=5.73 $Y=2.465
+ $X2=0 $Y2=0
cc_400 N_A_758_359#_M1012_g N_A_1266_147#_c_764_n 0.0138779f $X=6.255 $Y=2.155
+ $X2=0 $Y2=0
cc_401 N_A_758_359#_c_549_n N_A_1266_147#_c_760_n 0.00491544f $X=6.255 $Y=1.34
+ $X2=0 $Y2=0
cc_402 N_A_758_359#_M1017_g N_A_1266_147#_c_761_n 8.03855e-19 $X=5.73 $Y=2.465
+ $X2=0 $Y2=0
cc_403 N_A_758_359#_M1012_g N_A_1266_147#_c_761_n 0.0100352f $X=6.255 $Y=2.155
+ $X2=0 $Y2=0
cc_404 N_A_758_359#_c_549_n N_A_1266_147#_c_761_n 0.00362929f $X=6.255 $Y=1.34
+ $X2=0 $Y2=0
cc_405 N_A_758_359#_c_562_n N_VPWR_M1006_d 0.00511906f $X=4.9 $Y=1.86 $X2=0
+ $Y2=0
cc_406 N_A_758_359#_M1006_g N_VPWR_c_800_n 0.00727313f $X=3.865 $Y=2.665 $X2=0
+ $Y2=0
cc_407 N_A_758_359#_c_560_n N_VPWR_c_800_n 0.00303738f $X=4.035 $Y=1.985 $X2=0
+ $Y2=0
cc_408 N_A_758_359#_c_562_n N_VPWR_c_800_n 0.0305901f $X=4.9 $Y=1.86 $X2=0 $Y2=0
cc_409 N_A_758_359#_c_563_n N_VPWR_c_800_n 0.00944578f $X=4.21 $Y=1.86 $X2=0
+ $Y2=0
cc_410 N_A_758_359#_M1006_g N_VPWR_c_801_n 0.00395991f $X=3.865 $Y=2.665 $X2=0
+ $Y2=0
cc_411 N_A_758_359#_c_564_n N_VPWR_c_801_n 0.0152735f $X=4.995 $Y=2.89 $X2=0
+ $Y2=0
cc_412 N_A_758_359#_M1017_g N_VPWR_c_802_n 0.00755798f $X=5.73 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_A_758_359#_c_544_n N_VPWR_c_802_n 0.00384035f $X=6.18 $Y=1.34 $X2=0
+ $Y2=0
cc_414 N_A_758_359#_M1012_g N_VPWR_c_802_n 0.00510139f $X=6.255 $Y=2.155 $X2=0
+ $Y2=0
cc_415 N_A_758_359#_M1012_g N_VPWR_c_803_n 0.00395948f $X=6.255 $Y=2.155 $X2=0
+ $Y2=0
cc_416 N_A_758_359#_M1006_g N_VPWR_c_808_n 0.00342046f $X=3.865 $Y=2.665 $X2=0
+ $Y2=0
cc_417 N_A_758_359#_M1017_g N_VPWR_c_809_n 0.00571722f $X=5.73 $Y=2.465 $X2=0
+ $Y2=0
cc_418 N_A_758_359#_c_564_n N_VPWR_c_809_n 0.0164167f $X=4.995 $Y=2.89 $X2=0
+ $Y2=0
cc_419 N_A_758_359#_M1012_g N_VPWR_c_810_n 0.00312414f $X=6.255 $Y=2.155 $X2=0
+ $Y2=0
cc_420 N_A_758_359#_M1006_g N_VPWR_c_797_n 0.00311419f $X=3.865 $Y=2.665 $X2=0
+ $Y2=0
cc_421 N_A_758_359#_M1017_g N_VPWR_c_797_n 0.01288f $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_422 N_A_758_359#_M1012_g N_VPWR_c_797_n 0.00410284f $X=6.255 $Y=2.155 $X2=0
+ $Y2=0
cc_423 N_A_758_359#_c_564_n N_VPWR_c_797_n 0.00993371f $X=4.995 $Y=2.89 $X2=0
+ $Y2=0
cc_424 N_A_758_359#_c_541_n N_Q_c_902_n 0.00320899f $X=5.655 $Y=1.34 $X2=0 $Y2=0
cc_425 N_A_758_359#_M1017_g N_Q_c_902_n 0.00183333f $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_426 N_A_758_359#_c_564_n N_Q_c_902_n 0.0835826f $X=4.995 $Y=2.89 $X2=0 $Y2=0
cc_427 N_A_758_359#_c_566_n N_Q_c_902_n 0.0105942f $X=4.995 $Y=1.94 $X2=0 $Y2=0
cc_428 N_A_758_359#_c_556_n N_Q_c_902_n 0.00185298f $X=5.23 $Y=1.34 $X2=0 $Y2=0
cc_429 N_A_758_359#_M1017_g N_Q_c_903_n 0.013459f $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_430 N_A_758_359#_c_541_n N_Q_c_899_n 0.0118785f $X=5.655 $Y=1.34 $X2=0 $Y2=0
cc_431 N_A_758_359#_c_542_n N_Q_c_899_n 0.00501999f $X=5.73 $Y=1.265 $X2=0 $Y2=0
cc_432 N_A_758_359#_M1017_g N_Q_c_899_n 0.0128984f $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_433 N_A_758_359#_M1012_g N_Q_c_899_n 0.00137985f $X=6.255 $Y=2.155 $X2=0
+ $Y2=0
cc_434 N_A_758_359#_c_548_n N_Q_c_899_n 0.00435802f $X=5.73 $Y=1.34 $X2=0 $Y2=0
cc_435 N_A_758_359#_c_552_n N_Q_c_899_n 0.00507586f $X=5.02 $Y=1.265 $X2=0 $Y2=0
cc_436 N_A_758_359#_c_553_n N_Q_c_899_n 0.00817916f $X=5.047 $Y=1.775 $X2=0
+ $Y2=0
cc_437 N_A_758_359#_c_555_n N_Q_c_899_n 0.0234152f $X=5.23 $Y=1.43 $X2=0 $Y2=0
cc_438 N_A_758_359#_c_556_n N_Q_c_899_n 0.00126753f $X=5.23 $Y=1.34 $X2=0 $Y2=0
cc_439 N_A_758_359#_c_542_n Q 0.00839311f $X=5.73 $Y=1.265 $X2=0 $Y2=0
cc_440 N_A_758_359#_c_545_n Q 4.06133e-19 $X=6.255 $Y=1.265 $X2=0 $Y2=0
cc_441 N_A_758_359#_c_551_n Q 0.0271119f $X=4.815 $Y=0.42 $X2=0 $Y2=0
cc_442 N_A_758_359#_c_542_n Q 0.00144787f $X=5.73 $Y=1.265 $X2=0 $Y2=0
cc_443 N_A_758_359#_c_554_n Q 0.0271119f $X=4.912 $Y=1.005 $X2=0 $Y2=0
cc_444 N_A_758_359#_c_556_n Q 0.00604931f $X=5.23 $Y=1.34 $X2=0 $Y2=0
cc_445 N_A_758_359#_M1001_g N_VGND_c_951_n 0.00486043f $X=4.025 $Y=0.445 $X2=0
+ $Y2=0
cc_446 N_A_758_359#_M1001_g N_VGND_c_952_n 0.0174216f $X=4.025 $Y=0.445 $X2=0
+ $Y2=0
cc_447 N_A_758_359#_c_551_n N_VGND_c_952_n 0.0406088f $X=4.815 $Y=0.42 $X2=0
+ $Y2=0
cc_448 N_A_758_359#_c_542_n N_VGND_c_953_n 0.00497865f $X=5.73 $Y=1.265 $X2=0
+ $Y2=0
cc_449 N_A_758_359#_c_544_n N_VGND_c_953_n 0.00573814f $X=6.18 $Y=1.34 $X2=0
+ $Y2=0
cc_450 N_A_758_359#_c_545_n N_VGND_c_953_n 0.00418301f $X=6.255 $Y=1.265 $X2=0
+ $Y2=0
cc_451 N_A_758_359#_c_545_n N_VGND_c_954_n 0.005177f $X=6.255 $Y=1.265 $X2=0
+ $Y2=0
cc_452 N_A_758_359#_c_542_n N_VGND_c_956_n 0.00496398f $X=5.73 $Y=1.265 $X2=0
+ $Y2=0
cc_453 N_A_758_359#_c_551_n N_VGND_c_956_n 0.0271551f $X=4.815 $Y=0.42 $X2=0
+ $Y2=0
cc_454 N_A_758_359#_c_545_n N_VGND_c_957_n 0.00361794f $X=6.255 $Y=1.265 $X2=0
+ $Y2=0
cc_455 N_A_758_359#_M1018_d N_VGND_c_959_n 0.00458033f $X=4.655 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_A_758_359#_M1001_g N_VGND_c_959_n 0.00818711f $X=4.025 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_A_758_359#_c_542_n N_VGND_c_959_n 0.0107661f $X=5.73 $Y=1.265 $X2=0
+ $Y2=0
cc_458 N_A_758_359#_c_545_n N_VGND_c_959_n 0.00440068f $X=6.255 $Y=1.265 $X2=0
+ $Y2=0
cc_459 N_A_758_359#_c_551_n N_VGND_c_959_n 0.0148902f $X=4.815 $Y=0.42 $X2=0
+ $Y2=0
cc_460 N_A_608_491#_c_677_n N_VPWR_c_799_n 0.0107446f $X=3.68 $Y=2.92 $X2=0
+ $Y2=0
cc_461 N_A_608_491#_M1009_g N_VPWR_c_800_n 0.00671172f $X=4.78 $Y=2.405 $X2=0
+ $Y2=0
cc_462 N_A_608_491#_c_672_n N_VPWR_c_800_n 0.0358343f $X=3.765 $Y=2.765 $X2=0
+ $Y2=0
cc_463 N_A_608_491#_M1009_g N_VPWR_c_801_n 0.00981735f $X=4.78 $Y=2.405 $X2=0
+ $Y2=0
cc_464 N_A_608_491#_c_677_n N_VPWR_c_801_n 0.0277251f $X=3.68 $Y=2.92 $X2=0
+ $Y2=0
cc_465 N_A_608_491#_c_672_n N_VPWR_c_801_n 0.00425737f $X=3.765 $Y=2.765 $X2=0
+ $Y2=0
cc_466 N_A_608_491#_c_677_n N_VPWR_c_808_n 0.0545993f $X=3.68 $Y=2.92 $X2=0
+ $Y2=0
cc_467 N_A_608_491#_M1009_g N_VPWR_c_809_n 0.00437283f $X=4.78 $Y=2.405 $X2=0
+ $Y2=0
cc_468 N_A_608_491#_M1019_d N_VPWR_c_797_n 0.00215176f $X=3.04 $Y=2.455 $X2=0
+ $Y2=0
cc_469 N_A_608_491#_M1009_g N_VPWR_c_797_n 0.00884586f $X=4.78 $Y=2.405 $X2=0
+ $Y2=0
cc_470 N_A_608_491#_c_677_n N_VPWR_c_797_n 0.0317468f $X=3.68 $Y=2.92 $X2=0
+ $Y2=0
cc_471 N_A_608_491#_c_677_n A_713_491# 0.00233862f $X=3.68 $Y=2.92 $X2=-0.19
+ $Y2=-0.245
cc_472 N_A_608_491#_c_672_n A_713_491# 0.00304046f $X=3.765 $Y=2.765 $X2=-0.19
+ $Y2=-0.245
cc_473 N_A_608_491#_M1009_g N_Q_c_902_n 0.00203647f $X=4.78 $Y=2.405 $X2=0 $Y2=0
cc_474 N_A_608_491#_M1009_g N_Q_c_899_n 3.02285e-19 $X=4.78 $Y=2.405 $X2=0 $Y2=0
cc_475 N_A_608_491#_c_673_n N_VGND_M1001_d 0.00247141f $X=4.38 $Y=1.06 $X2=0
+ $Y2=0
cc_476 N_A_608_491#_c_674_n N_VGND_c_951_n 0.0263166f $X=3.39 $Y=0.41 $X2=0
+ $Y2=0
cc_477 N_A_608_491#_c_669_n N_VGND_c_952_n 0.0168861f $X=4.58 $Y=1.185 $X2=0
+ $Y2=0
cc_478 N_A_608_491#_c_673_n N_VGND_c_952_n 0.0329885f $X=4.38 $Y=1.06 $X2=0
+ $Y2=0
cc_479 N_A_608_491#_c_674_n N_VGND_c_952_n 0.0237143f $X=3.39 $Y=0.41 $X2=0
+ $Y2=0
cc_480 N_A_608_491#_c_669_n N_VGND_c_956_n 0.00486043f $X=4.58 $Y=1.185 $X2=0
+ $Y2=0
cc_481 N_A_608_491#_M1003_d N_VGND_c_959_n 0.00327208f $X=3.2 $Y=0.235 $X2=0
+ $Y2=0
cc_482 N_A_608_491#_c_669_n N_VGND_c_959_n 0.00954696f $X=4.58 $Y=1.185 $X2=0
+ $Y2=0
cc_483 N_A_608_491#_c_674_n N_VGND_c_959_n 0.0212651f $X=3.39 $Y=0.41 $X2=0
+ $Y2=0
cc_484 N_A_1266_147#_c_764_n N_VPWR_c_802_n 0.0270736f $X=6.47 $Y=1.98 $X2=0
+ $Y2=0
cc_485 N_A_1266_147#_M1000_g N_VPWR_c_803_n 0.0237794f $X=7.205 $Y=2.465 $X2=0
+ $Y2=0
cc_486 N_A_1266_147#_c_764_n N_VPWR_c_803_n 0.0500515f $X=6.47 $Y=1.98 $X2=0
+ $Y2=0
cc_487 N_A_1266_147#_c_759_n N_VPWR_c_803_n 0.0248138f $X=7.07 $Y=1.51 $X2=0
+ $Y2=0
cc_488 N_A_1266_147#_c_760_n N_VPWR_c_803_n 0.00506784f $X=7.07 $Y=1.51 $X2=0
+ $Y2=0
cc_489 N_A_1266_147#_M1000_g N_VPWR_c_811_n 0.00486043f $X=7.205 $Y=2.465 $X2=0
+ $Y2=0
cc_490 N_A_1266_147#_M1000_g N_VPWR_c_797_n 0.00917987f $X=7.205 $Y=2.465 $X2=0
+ $Y2=0
cc_491 N_A_1266_147#_c_764_n N_VPWR_c_797_n 0.0128958f $X=6.47 $Y=1.98 $X2=0
+ $Y2=0
cc_492 N_A_1266_147#_c_758_n N_Q_c_899_n 0.00411004f $X=6.47 $Y=0.955 $X2=0
+ $Y2=0
cc_493 N_A_1266_147#_c_764_n N_Q_c_899_n 0.0034231f $X=6.47 $Y=1.98 $X2=0 $Y2=0
cc_494 N_A_1266_147#_c_761_n N_Q_c_899_n 0.00828655f $X=6.47 $Y=1.51 $X2=0 $Y2=0
cc_495 N_A_1266_147#_c_759_n Q_N 0.0271104f $X=7.07 $Y=1.51 $X2=0 $Y2=0
cc_496 N_A_1266_147#_c_762_n Q_N 0.0265179f $X=7.092 $Y=1.345 $X2=0 $Y2=0
cc_497 N_A_1266_147#_c_758_n N_VGND_c_953_n 0.0148326f $X=6.47 $Y=0.955 $X2=0
+ $Y2=0
cc_498 N_A_1266_147#_c_758_n N_VGND_c_954_n 0.0296459f $X=6.47 $Y=0.955 $X2=0
+ $Y2=0
cc_499 N_A_1266_147#_c_759_n N_VGND_c_954_n 0.0248138f $X=7.07 $Y=1.51 $X2=0
+ $Y2=0
cc_500 N_A_1266_147#_c_760_n N_VGND_c_954_n 0.00506784f $X=7.07 $Y=1.51 $X2=0
+ $Y2=0
cc_501 N_A_1266_147#_c_762_n N_VGND_c_954_n 0.0199851f $X=7.092 $Y=1.345 $X2=0
+ $Y2=0
cc_502 N_A_1266_147#_c_762_n N_VGND_c_958_n 0.00465077f $X=7.092 $Y=1.345 $X2=0
+ $Y2=0
cc_503 N_A_1266_147#_c_758_n N_VGND_c_959_n 0.0133834f $X=6.47 $Y=0.955 $X2=0
+ $Y2=0
cc_504 N_A_1266_147#_c_762_n N_VGND_c_959_n 0.00451796f $X=7.092 $Y=1.345 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_797_n A_536_491# 0.00275129f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_506 N_VPWR_c_797_n N_Q_M1017_s 0.00215158f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_507 N_VPWR_c_802_n N_Q_c_902_n 0.0476845f $X=5.995 $Y=1.98 $X2=0 $Y2=0
cc_508 N_VPWR_c_801_n N_Q_c_903_n 6.23601e-19 $X=4.565 $Y=2.89 $X2=0 $Y2=0
cc_509 N_VPWR_c_809_n N_Q_c_903_n 0.0200241f $X=5.835 $Y=3.33 $X2=0 $Y2=0
cc_510 N_VPWR_c_797_n N_Q_c_903_n 0.0120544f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_511 N_VPWR_c_797_n N_Q_N_M1000_d 0.00371702f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_512 N_VPWR_c_811_n Q_N 0.018528f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_513 N_VPWR_c_797_n Q_N 0.0104192f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_514 N_VPWR_c_802_n N_VGND_c_953_n 0.0108695f $X=5.995 $Y=1.98 $X2=0 $Y2=0
cc_515 Q N_VGND_c_953_n 0.037153f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_516 Q N_VGND_c_956_n 0.0224063f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_517 Q N_VGND_c_959_n 0.0121275f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_518 Q_N N_VGND_c_954_n 0.0307847f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_519 Q_N N_VGND_c_958_n 0.0108661f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_520 Q_N N_VGND_c_959_n 0.00974763f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_521 N_VGND_c_959_n A_568_47# 0.0027827f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
cc_522 N_VGND_c_959_n A_748_47# 0.0056084f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
