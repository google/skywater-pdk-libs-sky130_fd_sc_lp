# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.470000 0.775000 0.815000 1.445000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.385000 0.295000 5.675000 3.075000 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.775000 1.285000 1.105000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.085000  0.265000 0.535000 0.605000 ;
      RECT 0.085000  0.605000 0.300000 1.625000 ;
      RECT 0.085000  1.625000 1.155000 1.795000 ;
      RECT 0.085000  1.795000 0.365000 2.775000 ;
      RECT 0.585000  2.135000 0.795000 3.245000 ;
      RECT 0.705000  0.085000 0.950000 0.605000 ;
      RECT 0.985000  1.365000 2.480000 1.535000 ;
      RECT 0.985000  1.535000 1.155000 1.625000 ;
      RECT 1.015000  1.965000 1.690000 2.135000 ;
      RECT 1.015000  2.135000 1.335000 2.775000 ;
      RECT 1.120000  0.255000 2.220000 0.435000 ;
      RECT 1.120000  0.435000 1.425000 0.605000 ;
      RECT 1.335000  1.705000 1.690000 1.965000 ;
      RECT 1.545000  2.305000 2.820000 2.475000 ;
      RECT 1.545000  2.475000 1.875000 2.965000 ;
      RECT 1.765000  0.675000 2.025000 1.015000 ;
      RECT 1.765000  1.015000 2.820000 1.185000 ;
      RECT 2.070000  2.645000 2.400000 3.245000 ;
      RECT 2.195000  0.605000 2.570000 0.845000 ;
      RECT 2.220000  1.535000 2.480000 1.745000 ;
      RECT 2.400000  0.085000 2.570000 0.605000 ;
      RECT 2.650000  1.185000 2.820000 1.395000 ;
      RECT 2.650000  1.395000 3.120000 1.725000 ;
      RECT 2.650000  1.725000 2.820000 2.305000 ;
      RECT 3.000000  0.795000 4.465000 1.005000 ;
      RECT 3.015000  2.075000 3.460000 2.745000 ;
      RECT 3.290000  1.005000 3.460000 2.075000 ;
      RECT 3.665000  1.185000 3.995000 1.695000 ;
      RECT 3.665000  1.695000 4.805000 1.865000 ;
      RECT 3.900000  0.085000 4.230000 0.625000 ;
      RECT 3.955000  2.035000 4.285000 3.245000 ;
      RECT 4.205000  1.005000 4.465000 1.515000 ;
      RECT 4.400000  0.285000 4.805000 0.625000 ;
      RECT 4.455000  1.865000 4.715000 2.950000 ;
      RECT 4.635000  0.625000 4.805000 1.265000 ;
      RECT 4.635000  1.265000 5.215000 1.595000 ;
      RECT 4.635000  1.595000 4.805000 1.695000 ;
      RECT 4.905000  2.035000 5.215000 3.245000 ;
      RECT 4.975000  0.085000 5.215000 1.095000 ;
      RECT 4.975000  1.815000 5.215000 2.035000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__dlxtp_1
END LIBRARY
