* File: sky130_fd_sc_lp__srdlstp_1.pex.spice
* Created: Fri Aug 28 11:33:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%D 2 5 9 11 12 13 17 18
r34 17 19 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.342 $Y=1.12
+ $X2=0.342 $Y2=0.955
r35 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=1.12 $X2=0.29 $Y2=1.12
r36 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r37 12 18 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.12
r38 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.485 $Y=2.32
+ $X2=0.485 $Y2=1.625
r39 5 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.475 $Y=0.555
+ $X2=0.475 $Y2=0.955
r40 2 11 53.1843 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=0.342 $Y=1.408
+ $X2=0.342 $Y2=1.625
r41 1 17 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=0.342 $Y=1.172
+ $X2=0.342 $Y2=1.12
r42 1 2 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=0.342 $Y=1.172
+ $X2=0.342 $Y2=1.408
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%A_27_400# 1 2 9 11 15 19 22 24 26 28 34 37
r67 35 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.645
+ $X2=0.965 $Y2=1.81
r68 35 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.965 $Y=1.645
+ $X2=0.965 $Y2=1.555
r69 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.645 $X2=0.965 $Y2=1.645
r70 31 34 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.77 $Y=1.645
+ $X2=0.965 $Y2=1.645
r71 28 30 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.69 $Y=0.555
+ $X2=0.69 $Y2=0.785
r72 23 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.81
+ $X2=0.77 $Y2=1.645
r73 23 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.77 $Y=1.81
+ $X2=0.77 $Y2=1.98
r74 22 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.48
+ $X2=0.77 $Y2=1.645
r75 22 30 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.77 $Y=1.48
+ $X2=0.77 $Y2=0.785
r76 20 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=2.065
+ $X2=0.27 $Y2=2.065
r77 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=2.065
+ $X2=0.77 $Y2=1.98
r78 19 20 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.685 $Y=2.065
+ $X2=0.435 $Y2=2.065
r79 13 15 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.425 $Y=1.48
+ $X2=1.425 $Y2=0.97
r80 12 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.555
+ $X2=0.965 $Y2=1.555
r81 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=1.555
+ $X2=1.425 $Y2=1.48
r82 11 12 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.35 $Y=1.555
+ $X2=1.13 $Y2=1.555
r83 9 40 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.02 $Y=2.42 $X2=1.02
+ $Y2=1.81
r84 2 26 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2 $X2=0.27 $Y2=2.145
r85 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.345 $X2=0.69 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%SET_B 1 3 4 8 13 14 16 17 21 23 24 28
c88 17 0 1.42204e-19 $X=5.435 $Y=0.34
c89 1 0 1.36774e-19 $X=1.785 $Y=0.53
r90 32 34 2.27458 $w=2.95e-07 $l=5.5e-08 $layer=LI1_cond $X=5.6 $Y=0.395 $X2=5.6
+ $Y2=0.34
r91 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.6
+ $Y=0.395 $X2=5.6 $Y2=0.395
r92 28 31 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.6 $Y=0.305 $X2=5.6
+ $Y2=0.395
r93 24 32 6.61695 $w=2.95e-07 $l=1.6e-07 $layer=LI1_cond $X=5.6 $Y=0.555 $X2=5.6
+ $Y2=0.395
r94 20 23 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0.365
+ $X2=2.31 $Y2=0.365
r95 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.145
+ $Y=0.365 $X2=2.145 $Y2=0.365
r96 17 34 3.96227 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=0.34
+ $X2=5.6 $Y2=0.34
r97 17 23 203.877 $w=1.68e-07 $l=3.125e-06 $layer=LI1_cond $X=5.435 $Y=0.34
+ $X2=2.31 $Y2=0.34
r98 15 16 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.145 $Y=1.165
+ $X2=6.145 $Y2=1.315
r99 14 21 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.86 $Y=0.365
+ $X2=2.145 $Y2=0.365
r100 13 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.235 $Y=0.845
+ $X2=6.235 $Y2=1.165
r101 10 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.235 $Y=0.38
+ $X2=6.235 $Y2=0.845
r102 8 16 221.124 $w=2.5e-07 $l=8.9e-07 $layer=POLY_cond $X=6.105 $Y=2.205
+ $X2=6.105 $Y2=1.315
r103 5 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.765 $Y=0.305
+ $X2=5.6 $Y2=0.305
r104 4 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.16 $Y=0.305
+ $X2=6.235 $Y2=0.38
r105 4 5 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.16 $Y=0.305
+ $X2=5.765 $Y2=0.305
r106 1 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.785 $Y=0.53
+ $X2=1.86 $Y2=0.365
r107 1 3 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.785 $Y=0.53
+ $X2=1.785 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%A_404_353# 1 2 7 9 12 14 15 18 22 26 32 33
+ 34 36 38 39 42 44 45 49 52 53 57 58 61 64 65
c198 57 0 4.12437e-20 $X=4.235 $Y=1.29
c199 52 0 1.9477e-19 $X=3.19 $Y=1.93
c200 18 0 1.70449e-19 $X=3.065 $Y=2.675
c201 14 0 5.8124e-20 $X=2.99 $Y=1.84
r202 63 65 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=8.59 $Y=1.08
+ $X2=8.755 $Y2=1.08
r203 63 64 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=8.59 $Y=1.08
+ $X2=8.425 $Y2=1.08
r204 58 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.29
+ $X2=4.235 $Y2=1.125
r205 57 60 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.235 $Y=1.29
+ $X2=4.235 $Y2=1.455
r206 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.235
+ $Y=1.29 $X2=4.235 $Y2=1.29
r207 53 66 21.6727 $w=2.78e-07 $l=1.25e-07 $layer=POLY_cond $X=3.19 $Y=1.93
+ $X2=3.065 $Y2=1.93
r208 52 55 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.19 $Y=1.93
+ $X2=3.19 $Y2=2.095
r209 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.93 $X2=3.19 $Y2=1.93
r210 47 49 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.23 $Y=1.31
+ $X2=9.23 $Y2=1.985
r211 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.065 $Y=1.225
+ $X2=9.23 $Y2=1.31
r212 45 65 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=9.065 $Y=1.225
+ $X2=8.755 $Y2=1.225
r213 44 64 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.09 $Y=1.225
+ $X2=8.425 $Y2=1.225
r214 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.005 $Y=1.31
+ $X2=8.09 $Y2=1.225
r215 41 42 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=8.005 $Y=1.31
+ $X2=8.005 $Y2=2.315
r216 40 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.4 $Y=2.4 $X2=4.315
+ $Y2=2.4
r217 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.92 $Y=2.4
+ $X2=8.005 $Y2=2.315
r218 39 40 229.647 $w=1.68e-07 $l=3.52e-06 $layer=LI1_cond $X=7.92 $Y=2.4
+ $X2=4.4 $Y2=2.4
r219 37 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=2.485
+ $X2=4.315 $Y2=2.4
r220 37 38 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.315 $Y=2.485
+ $X2=4.315 $Y2=2.905
r221 36 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=2.315
+ $X2=4.315 $Y2=2.4
r222 36 60 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=4.315 $Y=2.315
+ $X2=4.315 $Y2=1.455
r223 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.23 $Y=2.99
+ $X2=4.315 $Y2=2.905
r224 33 34 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=4.23 $Y=2.99
+ $X2=3.355 $Y2=2.99
r225 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.27 $Y=2.905
+ $X2=3.355 $Y2=2.99
r226 32 55 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.27 $Y=2.905
+ $X2=3.27 $Y2=2.095
r227 28 30 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.095 $Y=1.84
+ $X2=2.31 $Y2=1.84
r228 26 70 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.145 $Y=0.445
+ $X2=4.145 $Y2=1.125
r229 20 53 40.7446 $w=2.78e-07 $l=3.06594e-07 $layer=POLY_cond $X=3.425 $Y=2.095
+ $X2=3.19 $Y2=1.93
r230 20 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.425 $Y=2.095
+ $X2=3.425 $Y2=2.675
r231 16 66 17.1848 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=2.095
+ $X2=3.065 $Y2=1.93
r232 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.065 $Y=2.095
+ $X2=3.065 $Y2=2.675
r233 15 30 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.385 $Y=1.84
+ $X2=2.31 $Y2=1.84
r234 14 66 23.1551 $w=2.78e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.99 $Y=1.84
+ $X2=3.065 $Y2=1.93
r235 14 15 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=2.99 $Y=1.84
+ $X2=2.385 $Y2=1.84
r236 10 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.31 $Y=1.765
+ $X2=2.31 $Y2=1.84
r237 10 12 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.31 $Y=1.765
+ $X2=2.31 $Y2=1.08
r238 7 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.095 $Y=1.915
+ $X2=2.095 $Y2=1.84
r239 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.095 $Y=1.915
+ $X2=2.095 $Y2=2.345
r240 2 49 600 $w=1.7e-07 $l=4.54973e-07 $layer=licon1_PDIFF $count=1 $X=8.975
+ $Y=2.33 $X2=9.23 $Y2=1.985
r241 1 63 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.45
+ $Y=0.87 $X2=8.59 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%A_434_405# 1 2 7 9 10 14 17 20 22 23 24 25
+ 27 29 35 38 43
c96 43 0 1.36774e-19 $X=2.69 $Y=1.052
c97 35 0 5.8124e-20 $X=2.995 $Y=1.15
c98 27 0 3.24855e-20 $X=2.33 $Y=1.665
c99 25 0 9.60127e-20 $X=3.67 $Y=1.695
c100 23 0 9.87575e-20 $X=3.26 $Y=1.15
c101 14 0 4.12437e-20 $X=3.62 $Y=0.555
r102 42 43 5.97863 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=1.052
+ $X2=2.69 $Y2=1.052
r103 39 42 2.70326 $w=4.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.43 $Y=1.052
+ $X2=2.525 $Y2=1.052
r104 35 43 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.995 $Y=1.12
+ $X2=2.69 $Y2=1.12
r105 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.995
+ $Y=1.15 $X2=2.995 $Y2=1.15
r106 31 39 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=2.43 $Y=1.255
+ $X2=2.43 $Y2=1.052
r107 31 38 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.43 $Y=1.255
+ $X2=2.43 $Y2=1.48
r108 27 38 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.33 $Y=1.665
+ $X2=2.33 $Y2=1.48
r109 27 29 15.7293 $w=3.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.33 $Y=1.665
+ $X2=2.33 $Y2=2.17
r110 22 36 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.185 $Y=1.15
+ $X2=2.995 $Y2=1.15
r111 22 23 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=3.185 $Y=1.15
+ $X2=3.26 $Y2=1.15
r112 18 25 90.0579 $w=1.9e-07 $l=3.55e-07 $layer=POLY_cond $X=4.025 $Y=1.695
+ $X2=3.67 $Y2=1.695
r113 18 20 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=4.025 $Y=1.845
+ $X2=4.025 $Y2=2.595
r114 17 25 8.39207 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.67 $Y=1.545
+ $X2=3.67 $Y2=1.695
r115 16 24 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=3.67 $Y=1.315
+ $X2=3.645 $Y2=1.24
r116 16 17 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.67 $Y=1.315
+ $X2=3.67 $Y2=1.545
r117 12 24 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=3.62 $Y=1.165
+ $X2=3.645 $Y2=1.24
r118 12 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.62 $Y=1.165
+ $X2=3.62 $Y2=0.555
r119 11 23 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.335 $Y=1.24
+ $X2=3.26 $Y2=1.15
r120 10 24 5.30422 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=3.545 $Y=1.24
+ $X2=3.645 $Y2=1.24
r121 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.545 $Y=1.24
+ $X2=3.335 $Y2=1.24
r122 7 23 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=0.985
+ $X2=3.26 $Y2=1.15
r123 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.26 $Y=0.985
+ $X2=3.26 $Y2=0.555
r124 2 29 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.17
+ $Y=2.025 $X2=2.31 $Y2=2.17
r125 1 42 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.87 $X2=2.525 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%A_878_357# 1 2 9 11 13 14 15 16 18 20 21
+ 24 25 27 28 31 33 36 37
c109 25 0 4.16224e-20 $X=4.805 $Y=1.77
c110 14 0 1.42204e-19 $X=4.79 $Y=0.84
r111 36 38 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=7.585 $Y=1.915
+ $X2=7.585 $Y2=2.06
r112 36 37 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=7.585 $Y=1.915
+ $X2=7.585 $Y2=1.685
r113 31 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.04 $Y=0.885
+ $X2=7.665 $Y2=0.885
r114 31 33 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.04 $Y=0.8
+ $X2=8.04 $Y2=0.655
r115 29 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=0.97
+ $X2=7.665 $Y2=0.885
r116 29 37 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=7.665 $Y=0.97
+ $X2=7.665 $Y2=1.685
r117 27 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.42 $Y=2.06
+ $X2=7.585 $Y2=2.06
r118 27 28 159.84 $w=1.68e-07 $l=2.45e-06 $layer=LI1_cond $X=7.42 $Y=2.06
+ $X2=4.97 $Y2=2.06
r119 25 46 11.4762 $w=2.52e-07 $l=6e-08 $layer=POLY_cond $X=4.805 $Y=1.77
+ $X2=4.865 $Y2=1.77
r120 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.805
+ $Y=1.77 $X2=4.805 $Y2=1.77
r121 22 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.805 $Y=1.975
+ $X2=4.97 $Y2=2.06
r122 22 24 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.805 $Y=1.975
+ $X2=4.805 $Y2=1.77
r123 20 46 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.865 $Y=1.605
+ $X2=4.865 $Y2=1.77
r124 19 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.865 $Y=0.915
+ $X2=4.865 $Y2=0.84
r125 19 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.865 $Y=0.915
+ $X2=4.865 $Y2=1.605
r126 16 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.865 $Y=0.765
+ $X2=4.865 $Y2=0.84
r127 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.865 $Y=0.765
+ $X2=4.865 $Y2=0.445
r128 14 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.79 $Y=0.84
+ $X2=4.865 $Y2=0.84
r129 14 15 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.79 $Y=0.84
+ $X2=4.58 $Y2=0.84
r130 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.505 $Y=0.765
+ $X2=4.58 $Y2=0.84
r131 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.505 $Y=0.765
+ $X2=4.505 $Y2=0.445
r132 7 25 55.4683 $w=2.52e-07 $l=3.63249e-07 $layer=POLY_cond $X=4.515 $Y=1.935
+ $X2=4.805 $Y2=1.77
r133 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.515 $Y=1.935
+ $X2=4.515 $Y2=2.595
r134 2 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.445
+ $Y=1.705 $X2=7.585 $Y2=1.915
r135 1 33 182 $w=1.7e-07 $l=2.64811e-07 $layer=licon1_NDIFF $count=1 $X=7.785
+ $Y=0.635 $X2=8.04 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%A_1294_315# 1 2 10 11 13 15 16 18 19 20 24
+ 27 31 33 36 39
c100 31 0 6.72782e-20 $X=8.215 $Y=2.91
r101 36 38 8.62598 $w=3.38e-07 $l=2.3e-07 $layer=LI1_cond $X=10.425 $Y=0.865
+ $X2=10.425 $Y2=1.095
r102 31 42 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=8.215 $Y=2.91
+ $X2=8.215 $Y2=3.15
r103 30 33 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.215 $Y=2.91
+ $X2=8.345 $Y2=2.91
r104 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.215
+ $Y=2.91 $X2=8.215 $Y2=2.91
r105 25 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.38 $Y=2.49
+ $X2=10.38 $Y2=2.405
r106 25 27 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=10.38 $Y=2.49
+ $X2=10.38 $Y2=2.695
r107 24 38 41.027 $w=2.48e-07 $l=8.9e-07 $layer=LI1_cond $X=10.38 $Y=1.985
+ $X2=10.38 $Y2=1.095
r108 22 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.38 $Y=2.32
+ $X2=10.38 $Y2=2.405
r109 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=10.38 $Y=2.32
+ $X2=10.38 $Y2=1.985
r110 19 39 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.255 $Y=2.405
+ $X2=10.38 $Y2=2.405
r111 19 20 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=10.255 $Y=2.405
+ $X2=8.43 $Y2=2.405
r112 18 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.345 $Y=2.745
+ $X2=8.345 $Y2=2.91
r113 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.345 $Y=2.49
+ $X2=8.43 $Y2=2.405
r114 17 18 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.345 $Y=2.49
+ $X2=8.345 $Y2=2.745
r115 15 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.05 $Y=3.15
+ $X2=8.215 $Y2=3.15
r116 15 16 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=8.05 $Y=3.15
+ $X2=6.72 $Y2=3.15
r117 11 13 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.77 $Y=1.345
+ $X2=6.77 $Y2=0.845
r118 8 16 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=6.595 $Y=3.075
+ $X2=6.72 $Y2=3.15
r119 8 10 216.155 $w=2.5e-07 $l=8.7e-07 $layer=POLY_cond $X=6.595 $Y=3.075
+ $X2=6.595 $Y2=2.205
r120 7 11 71.895 $w=2.38e-07 $l=4.33763e-07 $layer=POLY_cond $X=6.595 $Y=1.7
+ $X2=6.77 $Y2=1.345
r121 7 10 125.469 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.595 $Y=1.7
+ $X2=6.595 $Y2=2.205
r122 2 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=10.28
+ $Y=1.84 $X2=10.42 $Y2=2.695
r123 2 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.28
+ $Y=1.84 $X2=10.42 $Y2=1.985
r124 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.29
+ $Y=0.655 $X2=10.43 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%GATE 1 2 5 9 12 13 14 18
c44 13 0 1.63376e-19 $X=8.4 $Y=1.665
r45 13 14 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=8.45 $Y=1.645
+ $X2=8.45 $Y2=2.035
r46 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.45
+ $Y=1.645 $X2=8.45 $Y2=1.645
r47 11 18 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.45 $Y=1.63
+ $X2=8.45 $Y2=1.645
r48 7 12 20.4101 $w=1.5e-07 $l=7.88987e-08 $layer=POLY_cond $X=8.915 $Y=1.48
+ $X2=8.907 $Y2=1.555
r49 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=8.915 $Y=1.48 $X2=8.915
+ $Y2=1.08
r50 3 12 20.4101 $w=1.5e-07 $l=7.84219e-08 $layer=POLY_cond $X=8.9 $Y=1.63
+ $X2=8.907 $Y2=1.555
r51 3 5 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=8.9 $Y=1.63 $X2=8.9
+ $Y2=2.65
r52 2 11 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.615 $Y=1.555
+ $X2=8.45 $Y2=1.63
r53 1 12 5.30422 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=8.825 $Y=1.555
+ $X2=8.907 $Y2=1.555
r54 1 2 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.825 $Y=1.555
+ $X2=8.615 $Y2=1.555
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%SLEEP_B 3 7 11 13 14 17 19 23 27 33 37 39
+ 40 44 45
c71 44 0 1.67603e-19 $X=10.89 $Y=1.645
c72 14 0 9.60979e-20 $X=9.74 $Y=1.555
r73 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.89
+ $Y=1.645 $X2=10.89 $Y2=1.645
r74 39 40 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.87 $Y=1.665
+ $X2=10.87 $Y2=2.035
r75 39 45 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=10.87 $Y=1.665
+ $X2=10.87 $Y2=1.645
r76 36 44 2.58377 $w=3.35e-07 $l=1.5e-08 $layer=POLY_cond $X=10.887 $Y=1.63
+ $X2=10.887 $Y2=1.645
r77 36 37 60.5064 $w=1.5e-07 $l=1.18e-07 $layer=POLY_cond $X=10.887 $Y=1.555
+ $X2=11.005 $Y2=1.555
r78 34 36 124.089 $w=1.5e-07 $l=2.42e-07 $layer=POLY_cond $X=10.645 $Y=1.555
+ $X2=10.887 $Y2=1.555
r79 31 32 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=9.445 $Y=1.555
+ $X2=9.665 $Y2=1.555
r80 29 31 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=9.305 $Y=1.555
+ $X2=9.445 $Y2=1.555
r81 25 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.005 $Y=1.48
+ $X2=11.005 $Y2=1.555
r82 25 27 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=11.005 $Y=1.48
+ $X2=11.005 $Y2=0.865
r83 21 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.645 $Y=1.48
+ $X2=10.645 $Y2=1.555
r84 21 23 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=10.645 $Y=1.48
+ $X2=10.645 $Y2=0.865
r85 20 33 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=10.28 $Y=1.555
+ $X2=10.155 $Y2=1.555
r86 19 34 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.57 $Y=1.555
+ $X2=10.645 $Y2=1.555
r87 19 20 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=10.57 $Y=1.555
+ $X2=10.28 $Y2=1.555
r88 15 33 1.63566 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.155 $Y=1.63
+ $X2=10.155 $Y2=1.555
r89 15 17 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=10.155 $Y=1.63
+ $X2=10.155 $Y2=2.34
r90 14 32 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.74 $Y=1.555
+ $X2=9.665 $Y2=1.555
r91 13 33 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=10.03 $Y=1.555
+ $X2=10.155 $Y2=1.555
r92 13 14 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=10.03 $Y=1.555
+ $X2=9.74 $Y2=1.555
r93 9 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.665 $Y=1.48
+ $X2=9.665 $Y2=1.555
r94 9 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=9.665 $Y=1.48 $X2=9.665
+ $Y2=1.08
r95 5 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.445 $Y=1.63
+ $X2=9.445 $Y2=1.555
r96 5 7 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.445 $Y=1.63
+ $X2=9.445 $Y2=2.16
r97 1 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.305 $Y=1.48
+ $X2=9.305 $Y2=1.555
r98 1 3 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=9.305 $Y=1.48 $X2=9.305
+ $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%A_700_451# 1 2 3 13 16 18 19 20 24 29 32
+ 36 38 40 42 43 44 47 48 49 50 52 56 60 66 69
c183 43 0 4.16224e-20 $X=3.755 $Y=2.075
c184 40 0 1.01441e-19 $X=3.755 $Y=2.405
r185 69 70 32.1566 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=7.265 $Y=1.26
+ $X2=7.265 $Y2=1.185
r186 67 72 31.8923 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.265 $Y=1.35
+ $X2=7.265 $Y2=1.515
r187 67 69 14.4261 $w=3.6e-07 $l=9e-08 $layer=POLY_cond $X=7.265 $Y=1.35
+ $X2=7.265 $Y2=1.26
r188 66 68 7.9931 $w=2.9e-07 $l=1.9e-07 $layer=LI1_cond $X=7.245 $Y=1.35
+ $X2=7.245 $Y2=1.54
r189 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.25
+ $Y=1.35 $X2=7.25 $Y2=1.35
r190 60 63 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.725 $Y=1.54
+ $X2=5.725 $Y2=1.72
r191 56 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.225 $Y=1.37
+ $X2=5.225 $Y2=1.54
r192 53 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=1.54
+ $X2=5.725 $Y2=1.54
r193 52 68 3.86198 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.08 $Y=1.54
+ $X2=7.245 $Y2=1.54
r194 52 53 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=7.08 $Y=1.54
+ $X2=5.89 $Y2=1.54
r195 51 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=1.54
+ $X2=5.225 $Y2=1.54
r196 50 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.56 $Y=1.54
+ $X2=5.725 $Y2=1.54
r197 50 51 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.56 $Y=1.54
+ $X2=5.31 $Y2=1.54
r198 48 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=1.37
+ $X2=5.225 $Y2=1.37
r199 48 49 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.14 $Y=1.37 $X2=4.74
+ $Y2=1.37
r200 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.655 $Y=1.285
+ $X2=4.74 $Y2=1.37
r201 46 47 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.655 $Y=0.895
+ $X2=4.655 $Y2=1.285
r202 45 55 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=0.745
+ $X2=3.755 $Y2=0.745
r203 44 46 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=4.57 $Y=0.745
+ $X2=4.655 $Y2=0.895
r204 44 45 28.0428 $w=2.98e-07 $l=7.3e-07 $layer=LI1_cond $X=4.57 $Y=0.745
+ $X2=3.84 $Y2=0.745
r205 42 55 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.755 $Y=0.895
+ $X2=3.755 $Y2=0.745
r206 42 43 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=3.755 $Y=0.895
+ $X2=3.755 $Y2=2.075
r207 38 43 7.1122 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=2.24
+ $X2=3.755 $Y2=2.075
r208 38 40 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=2.24
+ $X2=3.755 $Y2=2.405
r209 34 36 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=11.435 $Y=1.26
+ $X2=11.69 $Y2=1.26
r210 30 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.69 $Y=1.335
+ $X2=11.69 $Y2=1.26
r211 30 32 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=11.69 $Y=1.335
+ $X2=11.69 $Y2=2.155
r212 27 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.435 $Y=1.185
+ $X2=11.435 $Y2=1.26
r213 27 29 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.435 $Y=1.185
+ $X2=11.435 $Y2=0.865
r214 26 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.435 $Y=0.285
+ $X2=11.435 $Y2=0.865
r215 22 24 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.71 $Y=1.185
+ $X2=7.71 $Y2=0.845
r216 21 69 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.445 $Y=1.26
+ $X2=7.265 $Y2=1.26
r217 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.635 $Y=1.26
+ $X2=7.71 $Y2=1.185
r218 20 21 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.635 $Y=1.26
+ $X2=7.445 $Y2=1.26
r219 18 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.36 $Y=0.21
+ $X2=11.435 $Y2=0.285
r220 18 19 2094.65 $w=1.5e-07 $l=4.085e-06 $layer=POLY_cond $X=11.36 $Y=0.21
+ $X2=7.275 $Y2=0.21
r221 16 72 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.32 $Y=2.205
+ $X2=7.32 $Y2=1.515
r222 13 70 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.2 $Y=0.845 $X2=7.2
+ $Y2=1.185
r223 10 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.2 $Y=0.285
+ $X2=7.275 $Y2=0.21
r224 10 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.2 $Y=0.285
+ $X2=7.2 $Y2=0.845
r225 3 63 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.58
+ $Y=1.575 $X2=5.725 $Y2=1.72
r226 2 40 600 $w=1.7e-07 $l=3.21364e-07 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=2.255 $X2=3.755 $Y2=2.405
r227 1 55 182 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.235 $X2=3.835 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%A_2266_367# 1 2 9 13 15 16 19 23 27 30
c43 30 0 1.43064e-19 $X=11.31 $Y=1.475
c44 19 0 1.06489e-19 $X=11.475 $Y=1.98
r45 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.17
+ $Y=1.48 $X2=12.17 $Y2=1.48
r46 25 30 1.34256 $w=3.3e-07 $l=5.07494e-07 $layer=LI1_cond $X=11.815 $Y=1.48
+ $X2=11.31 $Y2=1.475
r47 25 27 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=11.815 $Y=1.48
+ $X2=12.17 $Y2=1.48
r48 21 30 5.16603 $w=3.3e-07 $l=4.12311e-07 $layer=LI1_cond $X=11.65 $Y=1.315
+ $X2=11.31 $Y2=1.475
r49 21 23 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=11.65 $Y=1.315
+ $X2=11.65 $Y2=0.865
r50 17 30 5.16603 $w=3.3e-07 $l=2.38642e-07 $layer=LI1_cond $X=11.475 $Y=1.645
+ $X2=11.31 $Y2=1.475
r51 17 19 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.475 $Y=1.645
+ $X2=11.475 $Y2=1.98
r52 15 28 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=12.38 $Y=1.48
+ $X2=12.17 $Y2=1.48
r53 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=12.38 $Y=1.48
+ $X2=12.455 $Y2=1.48
r54 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.455 $Y=1.645
+ $X2=12.455 $Y2=1.48
r55 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=12.455 $Y=1.645
+ $X2=12.455 $Y2=2.465
r56 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.455 $Y=1.315
+ $X2=12.455 $Y2=1.48
r57 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=12.455 $Y=1.315
+ $X2=12.455 $Y2=0.705
r58 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=11.33
+ $Y=1.835 $X2=11.475 $Y2=1.98
r59 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.51
+ $Y=0.655 $X2=11.65 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%VPWR 1 2 3 14 16 20 24 28 30 40 41 44 47
+ 50
r98 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r99 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 41 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r103 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r104 38 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.335 $Y=3.33
+ $X2=12.17 $Y2=3.33
r105 38 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.335 $Y=3.33
+ $X2=12.72 $Y2=3.33
r106 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r107 36 37 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=11.76
+ $Y=3.33 $X2=11.76 $Y2=3.33
r108 34 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 33 36 626.31 $w=1.68e-07 $l=9.6e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=11.76 $Y2=3.33
r110 33 34 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=2.16
+ $Y=3.33 $X2=2.16 $Y2=3.33
r111 31 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.775 $Y2=3.33
r112 31 33 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=2.16 $Y2=3.33
r113 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.005 $Y=3.33
+ $X2=12.17 $Y2=3.33
r114 30 36 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=12.005 $Y=3.33
+ $X2=11.76 $Y2=3.33
r115 28 37 1.47172 $w=4.9e-07 $l=5.28e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=11.76 $Y2=3.33
r116 28 34 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 24 27 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=12.17 $Y=1.98
+ $X2=12.17 $Y2=2.465
r118 22 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.17 $Y=3.245
+ $X2=12.17 $Y2=3.33
r119 22 27 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=12.17 $Y=3.245
+ $X2=12.17 $Y2=2.465
r120 18 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=3.33
r121 18 20 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=3.01
r122 17 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.805 $Y2=3.33
r123 16 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.775 $Y2=3.33
r124 16 17 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=0.97 $Y2=3.33
r125 12 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.33
r126 12 14 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=2.59
r127 3 27 300 $w=1.7e-07 $l=8.07496e-07 $layer=licon1_PDIFF $count=2 $X=11.765
+ $Y=1.835 $X2=12.17 $Y2=2.465
r128 3 24 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=11.765
+ $Y=1.835 $X2=12.17 $Y2=1.98
r129 2 20 600 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=1.64
+ $Y=2.025 $X2=1.775 $Y2=3.01
r130 1 14 600 $w=1.7e-07 $l=7.0189e-07 $layer=licon1_PDIFF $count=1 $X=0.56 $Y=2
+ $X2=0.805 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%A_217_130# 1 2 3 4 15 17 20 23 24 29 30 31
+ 36 37 38 40 41 42
c108 23 0 1.70449e-19 $X=2.685 $Y=2.59
r109 40 42 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.85 $Y=2.43
+ $X2=2.85 $Y2=2.59
r110 40 41 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=2.43
+ $X2=2.85 $Y2=2.265
r111 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.385 $Y=1.31
+ $X2=1.385 $Y2=1.98
r112 35 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.415 $Y=0.815
+ $X2=3.415 $Y2=1.425
r113 31 35 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.33 $Y=0.705
+ $X2=3.415 $Y2=0.815
r114 31 33 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=3.33 $Y=0.705
+ $X2=3.045 $Y2=0.705
r115 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.33 $Y=1.51
+ $X2=3.415 $Y2=1.425
r116 29 30 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.33 $Y=1.51
+ $X2=2.855 $Y2=1.51
r117 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=1.595
+ $X2=2.855 $Y2=1.51
r118 25 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.77 $Y=1.595
+ $X2=2.77 $Y2=2.265
r119 23 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=2.59
+ $X2=2.85 $Y2=2.59
r120 23 24 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.685 $Y=2.59
+ $X2=1.47 $Y2=2.59
r121 18 24 7.81568 $w=2.4e-07 $l=1.9799e-07 $layer=LI1_cond $X=1.31 $Y=2.505
+ $X2=1.47 $Y2=2.59
r122 18 20 12.965 $w=3.18e-07 $l=3.6e-07 $layer=LI1_cond $X=1.31 $Y=2.505
+ $X2=1.31 $Y2=2.145
r123 17 38 8.28018 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=1.31 $Y=2.14
+ $X2=1.31 $Y2=1.98
r124 17 20 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=1.31 $Y=2.14
+ $X2=1.31 $Y2=2.145
r125 13 37 10.0349 $w=4.23e-07 $l=2.12e-07 $layer=LI1_cond $X=1.257 $Y=1.098
+ $X2=1.257 $Y2=1.31
r126 13 15 8.21624 $w=4.23e-07 $l=3.03e-07 $layer=LI1_cond $X=1.257 $Y=1.098
+ $X2=1.257 $Y2=0.795
r127 4 40 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=2.715
+ $Y=2.255 $X2=2.85 $Y2=2.43
r128 3 20 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=2 $X2=1.235 $Y2=2.145
r129 2 33 182 $w=1.7e-07 $l=5.28819e-07 $layer=licon1_NDIFF $count=1 $X=2.92
+ $Y=0.235 $X2=3.045 $Y2=0.705
r130 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.65 $X2=1.21 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%KAPWR 1 2 3 4 13 19 23 32 37 40
c94 37 0 2.4539e-20 $X=9.36 $Y=2.82
r95 36 40 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=9.36 $Y=2.825
+ $X2=9.775 $Y2=2.825
r96 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=2.82
+ $X2=9.36 $Y2=2.82
r97 33 37 0.262345 $w=2.7e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=2.81
+ $X2=9.36 $Y2=2.81
r98 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.82
+ $X2=8.88 $Y2=2.82
r99 29 32 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=8.685 $Y=2.825
+ $X2=8.88 $Y2=2.825
r100 24 33 1.04938 $w=2.7e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=2.81
+ $X2=8.88 $Y2=2.81
r101 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=2.82
+ $X2=6.96 $Y2=2.82
r102 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.82
+ $X2=5.04 $Y2=2.82
r103 16 19 7.13417 $w=4.18e-07 $l=2.6e-07 $layer=LI1_cond $X=4.78 $Y=2.865
+ $X2=5.04 $Y2=2.865
r104 13 24 0.262345 $w=2.7e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=2.81
+ $X2=6.96 $Y2=2.81
r105 13 20 0.787035 $w=2.7e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=2.81
+ $X2=5.04 $Y2=2.81
r106 4 40 600 $w=1.7e-07 $l=1.10517e-06 $layer=licon1_PDIFF $count=1 $X=9.52
+ $Y=1.84 $X2=9.775 $Y2=2.825
r107 3 29 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=8.54
+ $Y=2.33 $X2=8.685 $Y2=2.825
r108 2 23 600 $w=1.7e-07 $l=1.23594e-06 $layer=licon1_PDIFF $count=1 $X=6.72
+ $Y=1.705 $X2=6.975 $Y2=2.82
r109 1 16 600 $w=1.7e-07 $l=8.37078e-07 $layer=licon1_PDIFF $count=1 $X=4.64
+ $Y=2.095 $X2=4.78 $Y2=2.865
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%Q 1 2 7 8 9 10 11 18
r14 11 32 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=12.67 $Y=1.98
+ $X2=12.67 $Y2=2.91
r15 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=12.67 $Y=1.665
+ $X2=12.67 $Y2=1.98
r16 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.67 $Y=1.295
+ $X2=12.67 $Y2=1.665
r17 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.67 $Y=0.925
+ $X2=12.67 $Y2=1.295
r18 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.67 $Y=0.555
+ $X2=12.67 $Y2=0.925
r19 7 18 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=12.67 $Y=0.555
+ $X2=12.67 $Y2=0.43
r20 2 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.835 $X2=12.67 $Y2=2.91
r21 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.835 $X2=12.67 $Y2=1.98
r22 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.53
+ $Y=0.285 $X2=12.67 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%VGND 1 2 3 4 5 6 7 22 24 27 28 33 37 41 45
+ 49 56 57 58 60 65 70 75 87 93 94 100 103 106 109 112
c144 28 0 3.24855e-20 $X=2 $Y=0.815
r145 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r146 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r147 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r148 103 104 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=0 $X2=6
+ $Y2=0
r149 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r150 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r151 94 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r152 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r153 91 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.325 $Y=0
+ $X2=12.2 $Y2=0
r154 91 93 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.325 $Y=0
+ $X2=12.72 $Y2=0
r155 90 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r156 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r157 87 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=12.2 $Y2=0
r158 87 89 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=11.76 $Y2=0
r159 86 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r160 86 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=9.84 $Y2=0
r161 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r162 83 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.045 $Y=0
+ $X2=9.88 $Y2=0
r163 83 85 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=10.045 $Y=0
+ $X2=10.8 $Y2=0
r164 82 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r165 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r166 79 82 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=9.36 $Y2=0
r167 79 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r168 78 81 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.44 $Y=0 $X2=9.36
+ $Y2=0
r169 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r170 76 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.15 $Y=0
+ $X2=6.985 $Y2=0
r171 76 78 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.15 $Y=0 $X2=7.44
+ $Y2=0
r172 75 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.715 $Y=0
+ $X2=9.88 $Y2=0
r173 75 81 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.715 $Y=0
+ $X2=9.36 $Y2=0
r174 71 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.185 $Y=0
+ $X2=6.06 $Y2=0
r175 71 73 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.185 $Y=0 $X2=6.48
+ $Y2=0
r176 70 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.82 $Y=0
+ $X2=6.985 $Y2=0
r177 70 73 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.48
+ $Y2=0
r178 69 104 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=6
+ $Y2=0
r179 69 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r180 68 69 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r181 66 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.725
+ $Y2=0
r182 66 68 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=2.16
+ $Y2=0
r183 65 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.935 $Y=0
+ $X2=6.06 $Y2=0
r184 65 68 246.283 $w=1.68e-07 $l=3.775e-06 $layer=LI1_cond $X=5.935 $Y=0
+ $X2=2.16 $Y2=0
r185 64 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r186 64 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r187 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r188 61 97 4.03846 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r189 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.72 $Y2=0
r190 60 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0 $X2=1.725
+ $Y2=0
r191 60 63 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.64 $Y=0 $X2=0.72
+ $Y2=0
r192 58 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r193 58 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r194 58 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r195 56 85 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=10.8 $Y2=0
r196 56 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=11.18 $Y2=0
r197 55 89 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=11.305 $Y=0
+ $X2=11.76 $Y2=0
r198 55 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.305 $Y=0
+ $X2=11.18 $Y2=0
r199 47 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.2 $Y=0.085
+ $X2=12.2 $Y2=0
r200 47 49 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=12.2 $Y=0.085
+ $X2=12.2 $Y2=0.43
r201 43 57 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.18 $Y=0.085
+ $X2=11.18 $Y2=0
r202 43 45 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=11.18 $Y=0.085
+ $X2=11.18 $Y2=0.865
r203 39 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.88 $Y=0.085
+ $X2=9.88 $Y2=0
r204 39 41 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=9.88 $Y=0.085
+ $X2=9.88 $Y2=1.08
r205 35 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=0.085
+ $X2=6.985 $Y2=0
r206 35 37 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=6.985 $Y=0.085
+ $X2=6.985 $Y2=0.815
r207 31 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.06 $Y=0.085
+ $X2=6.06 $Y2=0
r208 31 33 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=6.06 $Y=0.085
+ $X2=6.06 $Y2=0.78
r209 28 51 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2 $Y=0.73
+ $X2=1.725 $Y2=0.73
r210 28 30 5.91515 $w=3.3e-07 $l=1.6e-07 $layer=LI1_cond $X=2 $Y=0.815 $X2=2
+ $Y2=0.975
r211 27 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=0.645
+ $X2=1.725 $Y2=0.73
r212 26 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=0.085
+ $X2=1.725 $Y2=0
r213 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.725 $Y=0.085
+ $X2=1.725 $Y2=0.645
r214 22 97 3.10471 $w=2.5e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.172 $Y2=0
r215 22 24 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.22 $Y2=0.555
r216 7 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.1
+ $Y=0.285 $X2=12.24 $Y2=0.43
r217 6 45 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.08
+ $Y=0.655 $X2=11.22 $Y2=0.865
r218 5 41 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.74
+ $Y=0.87 $X2=9.88 $Y2=1.08
r219 4 37 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.845
+ $Y=0.635 $X2=6.985 $Y2=0.815
r220 3 33 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.885
+ $Y=0.635 $X2=6.02 $Y2=0.78
r221 2 30 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.65 $X2=2 $Y2=0.975
r222 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.345 $X2=0.26 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLSTP_1%A_988_47# 1 2 7 9 13 16 20
r44 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.565 $Y=0.925
+ $X2=5.565 $Y2=1.2
r45 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.14 $Y=0.76
+ $X2=5.14 $Y2=0.925
r46 11 13 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=6.515 $Y=1.115
+ $X2=6.515 $Y2=0.845
r47 10 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.65 $Y=1.2
+ $X2=5.565 $Y2=1.2
r48 9 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.39 $Y=1.2
+ $X2=6.515 $Y2=1.115
r49 9 10 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.39 $Y=1.2 $X2=5.65
+ $Y2=1.2
r50 8 18 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.265 $Y=0.925
+ $X2=5.14 $Y2=0.925
r51 7 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.925
+ $X2=5.565 $Y2=0.925
r52 7 8 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.48 $Y=0.925
+ $X2=5.265 $Y2=0.925
r53 2 13 182 $w=1.7e-07 $l=3.33879e-07 $layer=licon1_NDIFF $count=1 $X=6.31
+ $Y=0.635 $X2=6.555 $Y2=0.845
r54 1 16 182 $w=1.7e-07 $l=6.33739e-07 $layer=licon1_NDIFF $count=1 $X=4.94
+ $Y=0.235 $X2=5.18 $Y2=0.76
.ends

