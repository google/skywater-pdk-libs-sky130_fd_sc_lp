* File: sky130_fd_sc_lp__fa_lp.pex.spice
* Created: Fri Aug 28 10:35:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__FA_LP%A_84_209# 1 2 9 13 17 21 23 25 29 30 32 33 35
+ 36 37 38 41 42 44 46 47 49 50 51 56 59 64 68 69
c196 35 0 1.32001e-19 $X=2.86 $Y=1.545
c197 25 0 1.17014e-19 $X=7.945 $Y=2.595
c198 21 0 8.44273e-20 $X=7.795 $Y=0.915
r199 68 69 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.26 $Y=1.417
+ $X2=7.43 $Y2=1.417
r200 64 66 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.535 $Y=1.285
+ $X2=6.535 $Y2=1.55
r201 59 60 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.86 $Y=1.63 $X2=2.86
+ $Y2=1.83
r202 56 69 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=7.845 $Y=1.47
+ $X2=7.43 $Y2=1.47
r203 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.845
+ $Y=1.47 $X2=7.845 $Y2=1.47
r204 53 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.62 $Y=1.285
+ $X2=6.535 $Y2=1.285
r205 53 68 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.62 $Y=1.285
+ $X2=7.26 $Y2=1.285
r206 50 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=1.55
+ $X2=6.535 $Y2=1.55
r207 50 51 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=6.45 $Y=1.55
+ $X2=5.06 $Y2=1.55
r208 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=1.465
+ $X2=5.06 $Y2=1.55
r209 48 49 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.975 $Y=1
+ $X2=4.975 $Y2=1.465
r210 47 63 9.85688 $w=3.59e-07 $l=2.11305e-07 $layer=LI1_cond $X=3.605 $Y=0.915
+ $X2=3.415 $Y2=0.87
r211 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.89 $Y=0.915
+ $X2=4.975 $Y2=1
r212 46 47 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=4.89 $Y=0.915
+ $X2=3.605 $Y2=0.915
r213 42 44 11.7419 $w=2.63e-07 $l=2.7e-07 $layer=LI1_cond $X=3.425 $Y=2.582
+ $X2=3.695 $Y2=2.582
r214 41 42 7.24806 $w=2.65e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.34 $Y=2.45
+ $X2=3.425 $Y2=2.582
r215 40 41 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.34 $Y=1.915
+ $X2=3.34 $Y2=2.45
r216 39 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=1.83
+ $X2=2.86 $Y2=1.83
r217 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.255 $Y=1.83
+ $X2=3.34 $Y2=1.915
r218 38 39 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.255 $Y=1.83
+ $X2=2.945 $Y2=1.83
r219 36 63 7.29808 $w=3.59e-07 $l=1.9775e-07 $layer=LI1_cond $X=3.25 $Y=0.942
+ $X2=3.415 $Y2=0.87
r220 36 37 15.622 $w=2.23e-07 $l=3.05e-07 $layer=LI1_cond $X=3.25 $Y=0.942
+ $X2=2.945 $Y2=0.942
r221 35 59 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=1.545
+ $X2=2.86 $Y2=1.63
r222 34 37 6.9898 $w=2.25e-07 $l=1.49579e-07 $layer=LI1_cond $X=2.86 $Y=1.055
+ $X2=2.945 $Y2=0.942
r223 34 35 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.86 $Y=1.055
+ $X2=2.86 $Y2=1.545
r224 32 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=1.63
+ $X2=2.86 $Y2=1.63
r225 32 33 113.845 $w=1.68e-07 $l=1.745e-06 $layer=LI1_cond $X=2.775 $Y=1.63
+ $X2=1.03 $Y2=1.63
r226 30 71 63.4589 $w=6.1e-07 $l=5.05e-07 $layer=POLY_cond $X=0.725 $Y=1.21
+ $X2=0.725 $Y2=1.715
r227 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.865
+ $Y=1.21 $X2=0.865 $Y2=1.21
r228 27 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.865 $Y=1.545
+ $X2=1.03 $Y2=1.63
r229 27 29 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=1.545
+ $X2=0.865 $Y2=1.21
r230 23 57 47.2339 $w=3.08e-07 $l=3.2311e-07 $layer=POLY_cond $X=7.945 $Y=1.76
+ $X2=7.875 $Y2=1.47
r231 23 25 207.459 $w=2.5e-07 $l=8.35e-07 $layer=POLY_cond $X=7.945 $Y=1.76
+ $X2=7.945 $Y2=2.595
r232 19 57 38.5326 $w=3.08e-07 $l=2.0106e-07 $layer=POLY_cond $X=7.795 $Y=1.305
+ $X2=7.875 $Y2=1.47
r233 19 21 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=7.795 $Y=1.305
+ $X2=7.795 $Y2=0.915
r234 15 30 28.9593 $w=3.05e-07 $l=3.01413e-07 $layer=POLY_cond $X=0.955 $Y=1.045
+ $X2=0.725 $Y2=1.21
r235 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.955 $Y=1.045
+ $X2=0.955 $Y2=0.635
r236 11 30 28.9593 $w=3.05e-07 $l=2.20624e-07 $layer=POLY_cond $X=0.595 $Y=1.045
+ $X2=0.725 $Y2=1.21
r237 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.595 $Y=1.045
+ $X2=0.595 $Y2=0.635
r238 9 71 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.545 $Y=2.415
+ $X2=0.545 $Y2=1.715
r239 2 44 600 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=1 $X=3.555
+ $Y=2.095 $X2=3.695 $Y2=2.54
r240 1 63 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.275
+ $Y=0.705 $X2=3.415 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%B 1 3 4 6 8 10 12 13 15 16 18 20 21 23 24 26
+ 29 33 36 38 44 45 48 49 53 54 56 57 58 59 65 69
c192 54 0 6.36405e-20 $X=8.985 $Y=1.77
c193 49 0 9.52729e-20 $X=8.82 $Y=2.25
c194 38 0 2.16033e-20 $X=3.605 $Y=1.4
c195 29 0 1.7061e-19 $X=8.965 $Y=2.595
c196 13 0 1.94713e-19 $X=4.59 $Y=2.02
r197 65 67 52.5545 $w=3.21e-07 $l=3.5e-07 $layer=POLY_cond $X=4.6 $Y=1.382
+ $X2=4.95 $Y2=1.382
r198 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.6
+ $Y=1.4 $X2=4.6 $Y2=1.4
r199 63 65 9.00935 $w=3.21e-07 $l=6e-08 $layer=POLY_cond $X=4.54 $Y=1.382
+ $X2=4.6 $Y2=1.382
r200 57 58 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.04 $Y=2.217
+ $X2=4.21 $Y2=2.217
r201 54 70 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.985 $Y=1.77
+ $X2=8.985 $Y2=1.935
r202 54 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.985 $Y=1.77
+ $X2=8.985 $Y2=1.605
r203 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.985
+ $Y=1.77 $X2=8.985 $Y2=1.77
r204 51 53 14.4513 $w=3.13e-07 $l=3.95e-07 $layer=LI1_cond $X=8.977 $Y=2.165
+ $X2=8.977 $Y2=1.77
r205 49 51 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=8.82 $Y=2.25
+ $X2=8.977 $Y2=2.165
r206 49 58 300.759 $w=1.68e-07 $l=4.61e-06 $layer=LI1_cond $X=8.82 $Y=2.25
+ $X2=4.21 $Y2=2.25
r207 48 57 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.775 $Y=2.185
+ $X2=4.04 $Y2=2.185
r208 46 56 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.775 $Y=1.32
+ $X2=3.69 $Y2=1.4
r209 45 66 3.35256 $w=2.73e-07 $l=8e-08 $layer=LI1_cond $X=4.572 $Y=1.32
+ $X2=4.572 $Y2=1.4
r210 45 59 1.04768 $w=2.73e-07 $l=2.5e-08 $layer=LI1_cond $X=4.572 $Y=1.32
+ $X2=4.572 $Y2=1.295
r211 45 46 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.435 $Y=1.32
+ $X2=3.775 $Y2=1.32
r212 44 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.69 $Y=2.1
+ $X2=3.775 $Y2=2.185
r213 43 56 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.69 $Y=1.565
+ $X2=3.69 $Y2=1.4
r214 43 44 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.69 $Y=1.565
+ $X2=3.69 $Y2=2.1
r215 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.29
+ $Y=1.4 $X2=3.29 $Y2=1.4
r216 38 56 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=1.4
+ $X2=3.69 $Y2=1.4
r217 38 40 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.605 $Y=1.4
+ $X2=3.29 $Y2=1.4
r218 34 36 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.745 $Y=1.29
+ $X2=8.925 $Y2=1.29
r219 31 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.925 $Y=1.365
+ $X2=8.925 $Y2=1.29
r220 31 69 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.925 $Y=1.365
+ $X2=8.925 $Y2=1.605
r221 29 70 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.965 $Y=2.595
+ $X2=8.965 $Y2=1.935
r222 24 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.745 $Y=1.215
+ $X2=8.745 $Y2=1.29
r223 24 26 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=8.745 $Y=1.215 $X2=8.745
+ $Y2=0.915
r224 21 23 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.12 $Y=2.02
+ $X2=5.12 $Y2=2.595
r225 18 67 20.5661 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=4.95 $Y=1.2
+ $X2=4.95 $Y2=1.382
r226 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.95 $Y=1.2 $X2=4.95
+ $Y2=0.915
r227 17 33 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.715 $Y=1.945
+ $X2=4.59 $Y2=1.945
r228 16 21 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=4.995 $Y=1.945
+ $X2=5.12 $Y2=2.02
r229 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.995 $Y=1.945
+ $X2=4.715 $Y2=1.945
r230 13 33 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=4.59 $Y=2.02 $X2=4.59
+ $Y2=1.945
r231 13 15 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.59 $Y=2.02
+ $X2=4.59 $Y2=2.595
r232 12 33 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=4.54 $Y=1.87
+ $X2=4.59 $Y2=1.945
r233 11 63 20.5661 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=4.54 $Y=1.565
+ $X2=4.54 $Y2=1.382
r234 11 12 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=4.54 $Y=1.565
+ $X2=4.54 $Y2=1.87
r235 8 63 27.028 $w=3.21e-07 $l=2.56679e-07 $layer=POLY_cond $X=4.36 $Y=1.2
+ $X2=4.54 $Y2=1.382
r236 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.36 $Y=1.2 $X2=4.36
+ $Y2=0.915
r237 4 41 52.2154 $w=2.99e-07 $l=3.57176e-07 $layer=POLY_cond $X=3.43 $Y=1.715
+ $X2=3.34 $Y2=1.4
r238 4 6 218.639 $w=2.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.43 $Y=1.715
+ $X2=3.43 $Y2=2.595
r239 1 41 38.5562 $w=2.99e-07 $l=2.24332e-07 $layer=POLY_cond $X=3.2 $Y=1.235
+ $X2=3.34 $Y2=1.4
r240 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.2 $Y=1.235 $X2=3.2
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%CIN 1 3 8 12 16 20 24 28 31 32 33 34 38 40 41
+ 45 48 52
c153 40 0 2.87623e-19 $X=8.445 $Y=1.77
c154 38 0 9.52729e-20 $X=4.06 $Y=1.755
c155 24 0 1.94494e-19 $X=8.475 $Y=2.595
c156 20 0 1.01679e-19 $X=8.355 $Y=0.915
r157 49 61 5.96801 $w=2.78e-07 $l=1.45e-07 $layer=LI1_cond $X=6.94 $Y=1.755
+ $X2=6.94 $Y2=1.9
r158 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.915
+ $Y=1.755 $X2=6.915 $Y2=1.755
r159 45 49 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=6.94 $Y=1.665
+ $X2=6.94 $Y2=1.755
r160 41 56 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.77
+ $X2=8.445 $Y2=1.935
r161 41 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.77
+ $X2=8.445 $Y2=1.605
r162 40 43 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.445 $Y=1.77
+ $X2=8.445 $Y2=1.9
r163 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.445
+ $Y=1.77 $X2=8.445 $Y2=1.77
r164 38 53 30.6744 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=4.03 $Y=1.755
+ $X2=4.03 $Y2=1.92
r165 38 52 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=4.03 $Y=1.755
+ $X2=4.03 $Y2=1.59
r166 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=1.755 $X2=4.06 $Y2=1.755
r167 35 61 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.08 $Y=1.9 $X2=6.94
+ $Y2=1.9
r168 34 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=1.9
+ $X2=8.445 $Y2=1.9
r169 34 35 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=8.28 $Y=1.9
+ $X2=7.08 $Y2=1.9
r170 33 37 24.9926 $w=2.59e-07 $l=5.53624e-07 $layer=LI1_cond $X=4.56 $Y=1.9
+ $X2=4.06 $Y2=1.787
r171 32 61 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.8 $Y=1.9 $X2=6.94
+ $Y2=1.9
r172 32 33 146.139 $w=1.68e-07 $l=2.24e-06 $layer=LI1_cond $X=6.8 $Y=1.9
+ $X2=4.56 $Y2=1.9
r173 30 48 199.342 $w=3.3e-07 $l=1.14e-06 $layer=POLY_cond $X=5.775 $Y=1.755
+ $X2=6.915 $Y2=1.755
r174 30 31 1.50692 $w=3.3e-07 $l=4.25852e-07 $layer=POLY_cond $X=5.775 $Y=1.755
+ $X2=5.465 $Y2=1.48
r175 26 28 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=3.77 $Y=1.275
+ $X2=3.91 $Y2=1.275
r176 24 56 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.475 $Y=2.595
+ $X2=8.475 $Y2=1.935
r177 20 55 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.355 $Y=0.915
+ $X2=8.355 $Y2=1.605
r178 14 31 30.2679 $w=2e-07 $l=5.24404e-07 $layer=POLY_cond $X=5.65 $Y=1.92
+ $X2=5.465 $Y2=1.48
r179 14 16 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=5.65 $Y=1.92
+ $X2=5.65 $Y2=2.595
r180 10 31 30.2679 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=5.54 $Y=1.48
+ $X2=5.465 $Y2=1.48
r181 10 12 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=5.54 $Y=1.48
+ $X2=5.54 $Y2=0.915
r182 8 53 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.96 $Y=2.595
+ $X2=3.96 $Y2=1.92
r183 4 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.91 $Y=1.35
+ $X2=3.91 $Y2=1.275
r184 4 52 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.91 $Y=1.35
+ $X2=3.91 $Y2=1.59
r185 1 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=1.2 $X2=3.77
+ $Y2=1.275
r186 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.77 $Y=1.2 $X2=3.77
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%A 2 5 7 8 9 13 17 21 28 29 31 32 37 42 44 45
+ 46 50 52 53 54 55 61 62 64 65
c167 61 0 8.44273e-20 $X=7.07 $Y=0.43
c168 53 0 1.65463e-19 $X=9.425 $Y=1.365
c169 50 0 6.36405e-20 $X=9.315 $Y=0.9
c170 29 0 1.94494e-19 $X=7.415 $Y=2
c171 21 0 2.16033e-20 $X=2.81 $Y=0.915
c172 17 0 1.32001e-19 $X=2.215 $Y=0.915
c173 5 0 1.98572e-19 $X=1.635 $Y=2.545
r174 63 64 36.4263 $w=4.9e-07 $l=7.5e-08 $layer=POLY_cond $X=7.365 $Y=0.35
+ $X2=7.44 $Y2=0.35
r175 60 63 32.211 $w=4.9e-07 $l=2.95e-07 $layer=POLY_cond $X=7.07 $Y=0.35
+ $X2=7.365 $Y2=0.35
r176 60 62 46.2534 $w=4.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.07 $Y=0.35
+ $X2=6.905 $Y2=0.35
r177 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.07
+ $Y=0.43 $X2=7.07 $Y2=0.43
r178 55 61 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=7.07 $Y=0.555
+ $X2=7.07 $Y2=0.43
r179 55 65 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.07 $Y=0.555
+ $X2=6.905 $Y2=0.555
r180 55 65 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.89 $Y=0.555
+ $X2=6.905 $Y2=0.555
r181 54 55 20.5435 $w=2.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.48 $Y=0.555
+ $X2=6.89 $Y2=0.555
r182 52 53 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=9.425 $Y=1.215
+ $X2=9.425 $Y2=1.365
r183 48 50 48.7128 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=9.22 $Y=0.9
+ $X2=9.315 $Y2=0.9
r184 42 53 305.598 $w=2.5e-07 $l=1.23e-06 $layer=POLY_cond $X=9.485 $Y=2.595
+ $X2=9.485 $Y2=1.365
r185 38 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.315 $Y=0.975
+ $X2=9.315 $Y2=0.9
r186 38 52 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.315 $Y=0.975
+ $X2=9.315 $Y2=1.215
r187 35 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.22 $Y=0.825
+ $X2=9.22 $Y2=0.9
r188 35 37 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.22 $Y=0.825
+ $X2=9.22 $Y2=0.54
r189 34 37 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.22 $Y=0.255
+ $X2=9.22 $Y2=0.54
r190 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.145 $Y=0.18
+ $X2=9.22 $Y2=0.255
r191 32 64 874.266 $w=1.5e-07 $l=1.705e-06 $layer=POLY_cond $X=9.145 $Y=0.18
+ $X2=7.44 $Y2=0.18
r192 29 47 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=7.415 $Y=2
+ $X2=7.415 $Y2=1.875
r193 29 31 114.716 $w=2.5e-07 $l=5.95e-07 $layer=POLY_cond $X=7.415 $Y=2
+ $X2=7.415 $Y2=2.595
r194 28 47 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=7.365 $Y=0.915
+ $X2=7.365 $Y2=1.875
r195 25 63 30.8984 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=7.365 $Y=0.595
+ $X2=7.365 $Y2=0.35
r196 25 28 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.365 $Y=0.595
+ $X2=7.365 $Y2=0.915
r197 24 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=0.18
+ $X2=2.81 $Y2=0.18
r198 24 62 2061.32 $w=1.5e-07 $l=4.02e-06 $layer=POLY_cond $X=2.885 $Y=0.18
+ $X2=6.905 $Y2=0.18
r199 19 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.81 $Y=0.255
+ $X2=2.81 $Y2=0.18
r200 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.81 $Y=0.255
+ $X2=2.81 $Y2=0.915
r201 15 45 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=2.215 $Y=1.255
+ $X2=2.165 $Y2=1.33
r202 15 17 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.215 $Y=1.255
+ $X2=2.215 $Y2=0.915
r203 11 45 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=2.165 $Y=1.405
+ $X2=2.165 $Y2=1.33
r204 11 13 283.237 $w=2.5e-07 $l=1.14e-06 $layer=POLY_cond $X=2.165 $Y=1.405
+ $X2=2.165 $Y2=2.545
r205 10 44 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.76 $Y=1.33
+ $X2=1.635 $Y2=1.33
r206 9 45 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.04 $Y=1.33
+ $X2=2.165 $Y2=1.33
r207 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.04 $Y=1.33
+ $X2=1.76 $Y2=1.33
r208 7 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.735 $Y=0.18
+ $X2=2.81 $Y2=0.18
r209 7 8 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=2.735 $Y=0.18
+ $X2=1.66 $Y2=0.18
r210 3 44 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=1.635 $Y=1.405
+ $X2=1.635 $Y2=1.33
r211 3 5 283.237 $w=2.5e-07 $l=1.14e-06 $layer=POLY_cond $X=1.635 $Y=1.405
+ $X2=1.635 $Y2=2.545
r212 2 44 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=1.585 $Y=1.255
+ $X2=1.635 $Y2=1.33
r213 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.585 $Y=0.255
+ $X2=1.66 $Y2=0.18
r214 1 2 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=1.585 $Y=0.255
+ $X2=1.585 $Y2=1.255
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%A_1574_141# 1 2 7 9 10 11 14 16 18 22 23 24 25
+ 28 30 32 33 35 36 41 43 45 46
c102 33 0 7.00777e-20 $X=8.375 $Y=2.6
c103 28 0 1.24416e-19 $X=8.21 $Y=2.79
c104 22 0 1.65463e-19 $X=9.985 $Y=1.22
r105 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.985
+ $Y=1.385 $X2=9.985 $Y2=1.385
r106 37 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.485 $Y=1.305
+ $X2=9.4 $Y2=1.305
r107 36 45 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=9.82 $Y=1.305
+ $X2=9.97 $Y2=1.305
r108 36 37 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.82 $Y=1.305
+ $X2=9.485 $Y2=1.305
r109 34 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.4 $Y=1.39 $X2=9.4
+ $Y2=1.305
r110 34 35 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=9.4 $Y=1.39
+ $X2=9.4 $Y2=2.515
r111 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.315 $Y=2.6
+ $X2=9.4 $Y2=2.515
r112 32 33 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=9.315 $Y=2.6
+ $X2=8.375 $Y2=2.6
r113 31 41 16.0526 $w=3.04e-07 $l=4.87032e-07 $layer=LI1_cond $X=8.36 $Y=1.305
+ $X2=8.167 $Y2=0.905
r114 30 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.315 $Y=1.305
+ $X2=9.4 $Y2=1.305
r115 30 31 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=9.315 $Y=1.305
+ $X2=8.36 $Y2=1.305
r116 26 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.21 $Y=2.685
+ $X2=8.375 $Y2=2.6
r117 26 28 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=8.21 $Y=2.685
+ $X2=8.21 $Y2=2.79
r118 23 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.985 $Y=1.725
+ $X2=9.985 $Y2=1.385
r119 23 24 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.985 $Y=1.725
+ $X2=9.985 $Y2=1.89
r120 22 46 44.4756 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.985 $Y=1.22
+ $X2=9.985 $Y2=1.385
r121 19 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.065 $Y=0.975
+ $X2=10.065 $Y2=0.9
r122 19 22 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=10.065 $Y=0.975
+ $X2=10.065 $Y2=1.22
r123 16 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.065 $Y=0.825
+ $X2=10.065 $Y2=0.9
r124 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.065 $Y=0.825
+ $X2=10.065 $Y2=0.54
r125 14 24 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=10.015 $Y=2.595
+ $X2=10.015 $Y2=1.89
r126 10 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.99 $Y=0.9
+ $X2=10.065 $Y2=0.9
r127 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.99 $Y=0.9
+ $X2=9.78 $Y2=0.9
r128 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.705 $Y=0.825
+ $X2=9.78 $Y2=0.9
r129 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.705 $Y=0.825
+ $X2=9.705 $Y2=0.54
r130 2 28 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=2.095 $X2=8.21 $Y2=2.79
r131 1 41 182 $w=1.7e-07 $l=3.5623e-07 $layer=licon1_NDIFF $count=1 $X=7.87
+ $Y=0.705 $X2=8.14 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%COUT 1 2 7 8 9 10 11 12 13 24
r17 24 45 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=0.28 $Y=0.925 $X2=0.28
+ $Y2=0.865
r18 12 13 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.28 $Y=2.405
+ $X2=0.28 $Y2=2.77
r19 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=2.035
+ $X2=0.28 $Y2=2.405
r20 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.665
+ $X2=0.28 $Y2=2.035
r21 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.295
+ $X2=0.28 $Y2=1.665
r22 8 45 1.00085 $w=4.28e-07 $l=1.3e-08 $layer=LI1_cond $X=0.33 $Y=0.852
+ $X2=0.33 $Y2=0.865
r23 8 43 5.81582 $w=4.28e-07 $l=2.17e-07 $layer=LI1_cond $X=0.33 $Y=0.852
+ $X2=0.33 $Y2=0.635
r24 8 9 12.5023 $w=3.28e-07 $l=3.58e-07 $layer=LI1_cond $X=0.28 $Y=0.937
+ $X2=0.28 $Y2=1.295
r25 8 24 0.41907 $w=3.28e-07 $l=1.2e-08 $layer=LI1_cond $X=0.28 $Y=0.937
+ $X2=0.28 $Y2=0.925
r26 7 43 2.14408 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=0.33 $Y=0.555 $X2=0.33
+ $Y2=0.635
r27 2 13 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.915 $X2=0.28 $Y2=2.77
r28 2 11 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.915 $X2=0.28 $Y2=2.06
r29 1 43 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.425 $X2=0.38 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%VPWR 1 2 3 4 5 20 26 30 34 38 43 44 46 47 49
+ 50 51 63 72 73 76 79
r112 79 80 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r113 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r114 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r115 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r116 70 80 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=6 $Y2=3.33
r117 69 70 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r118 67 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=3.33
+ $X2=5.915 $Y2=3.33
r119 67 69 213.989 $w=1.68e-07 $l=3.28e-06 $layer=LI1_cond $X=6.08 $Y=3.33
+ $X2=9.36 $Y2=3.33
r120 66 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r121 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r122 63 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=3.33
+ $X2=5.915 $Y2=3.33
r123 63 65 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.75 $Y=3.33
+ $X2=5.52 $Y2=3.33
r124 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 59 62 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.56 $Y2=3.33
r126 58 61 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r128 56 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 56 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r131 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r132 53 55 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.68 $Y2=3.33
r133 51 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r134 51 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.56 $Y2=3.33
r135 49 69 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.665 $Y=3.33
+ $X2=9.36 $Y2=3.33
r136 49 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.665 $Y=3.33
+ $X2=9.79 $Y2=3.33
r137 48 72 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=9.915 $Y=3.33
+ $X2=10.32 $Y2=3.33
r138 48 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.915 $Y=3.33
+ $X2=9.79 $Y2=3.33
r139 46 61 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.69 $Y=3.33
+ $X2=4.56 $Y2=3.33
r140 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.69 $Y=3.33
+ $X2=4.855 $Y2=3.33
r141 45 65 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=5.02 $Y=3.33 $X2=5.52
+ $Y2=3.33
r142 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=4.855 $Y2=3.33
r143 43 55 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.68 $Y2=3.33
r144 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.9 $Y2=3.33
r145 42 58 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.16 $Y2=3.33
r146 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.9 $Y2=3.33
r147 38 41 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=9.79 $Y=2.24
+ $X2=9.79 $Y2=2.95
r148 36 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.79 $Y=3.245
+ $X2=9.79 $Y2=3.33
r149 36 41 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=9.79 $Y=3.245
+ $X2=9.79 $Y2=2.95
r150 32 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.915 $Y=3.245
+ $X2=5.915 $Y2=3.33
r151 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.915 $Y=3.245
+ $X2=5.915 $Y2=2.95
r152 28 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=3.245
+ $X2=4.855 $Y2=3.33
r153 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.855 $Y=3.245
+ $X2=4.855 $Y2=2.815
r154 24 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.9 $Y=3.245 $X2=1.9
+ $Y2=3.33
r155 24 26 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=1.9 $Y=3.245
+ $X2=1.9 $Y2=2.41
r156 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.06
+ $X2=0.81 $Y2=2.77
r157 18 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r158 18 23 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.77
r159 5 41 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=9.61
+ $Y=2.095 $X2=9.75 $Y2=2.95
r160 5 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.61
+ $Y=2.095 $X2=9.75 $Y2=2.24
r161 4 34 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=5.775
+ $Y=2.095 $X2=5.915 $Y2=2.95
r162 3 30 600 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=1 $X=4.715
+ $Y=2.095 $X2=4.855 $Y2=2.815
r163 2 26 300 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=2 $X=1.76
+ $Y=2.045 $X2=1.9 $Y2=2.41
r164 1 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.915 $X2=0.81 $Y2=2.77
r165 1 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.915 $X2=0.81 $Y2=2.06
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%A_245_409# 1 2 9 13 14 15 19 21
r43 21 23 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.33 $Y=1.98 $X2=2.33
+ $Y2=2.18
r44 17 19 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=2.95 $Y=2.265
+ $X2=2.95 $Y2=2.405
r45 16 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=2.18
+ $X2=2.33 $Y2=2.18
r46 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.825 $Y=2.18
+ $X2=2.95 $Y2=2.265
r47 15 16 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.825 $Y=2.18
+ $X2=2.415 $Y2=2.18
r48 13 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=1.98
+ $X2=2.33 $Y2=1.98
r49 13 14 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.245 $Y=1.98
+ $X2=1.535 $Y2=1.98
r50 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.37 $Y=2.19 $X2=1.37
+ $Y2=2.9
r51 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.37 $Y=2.065
+ $X2=1.535 $Y2=1.98
r52 7 9 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.37 $Y=2.065
+ $X2=1.37 $Y2=2.19
r53 2 19 600 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=2.095 $X2=2.99 $Y2=2.405
r54 1 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.045 $X2=1.37 $Y2=2.9
r55 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.045 $X2=1.37 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%A_458_409# 1 2 9 11 12 15
c37 12 0 4.93603e-20 $X=2.595 $Y=2.98
c38 9 0 1.49212e-19 $X=2.43 $Y=2.755
r39 13 15 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.225 $Y=2.895
+ $X2=4.225 $Y2=2.79
r40 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.06 $Y=2.98
+ $X2=4.225 $Y2=2.895
r41 11 12 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=4.06 $Y=2.98
+ $X2=2.595 $Y2=2.98
r42 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.43 $Y=2.895
+ $X2=2.595 $Y2=2.98
r43 7 9 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.43 $Y=2.895 $X2=2.43
+ $Y2=2.755
r44 2 15 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=4.085
+ $Y=2.095 $X2=4.225 $Y2=2.79
r45 1 9 600 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=2.045 $X2=2.43 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%A_1049_419# 1 2 9 11 12 15
c29 15 0 1.24416e-19 $X=7.68 $Y=2.79
c30 12 0 7.89914e-20 $X=5.55 $Y=2.6
c31 11 0 7.00777e-20 $X=7.515 $Y=2.6
c32 9 0 1.15722e-19 $X=5.385 $Y=2.79
r33 13 15 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.68 $Y=2.685
+ $X2=7.68 $Y2=2.79
r34 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.515 $Y=2.6
+ $X2=7.68 $Y2=2.685
r35 11 12 128.198 $w=1.68e-07 $l=1.965e-06 $layer=LI1_cond $X=7.515 $Y=2.6
+ $X2=5.55 $Y2=2.6
r36 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.385 $Y=2.685
+ $X2=5.55 $Y2=2.6
r37 7 9 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=5.385 $Y=2.685
+ $X2=5.385 $Y2=2.79
r38 2 15 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=2.095 $X2=7.68 $Y2=2.79
r39 1 9 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=5.245
+ $Y=2.095 $X2=5.385 $Y2=2.79
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%SUM 1 2 12 13 14 15 26
r24 19 26 2.01272 $w=3.53e-07 $l=6.2e-08 $layer=LI1_cond $X=10.292 $Y=0.863
+ $X2=10.292 $Y2=0.925
r25 15 28 6.5188 $w=3.53e-07 $l=1.04e-07 $layer=LI1_cond $X=10.292 $Y=0.936
+ $X2=10.292 $Y2=1.04
r26 15 26 0.357095 $w=3.53e-07 $l=1.1e-08 $layer=LI1_cond $X=10.292 $Y=0.936
+ $X2=10.292 $Y2=0.925
r27 15 19 0.389558 $w=3.53e-07 $l=1.2e-08 $layer=LI1_cond $X=10.292 $Y=0.851
+ $X2=10.292 $Y2=0.863
r28 14 15 10.0961 $w=3.53e-07 $l=3.11e-07 $layer=LI1_cond $X=10.292 $Y=0.54
+ $X2=10.292 $Y2=0.851
r29 13 28 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=10.385 $Y=2.075
+ $X2=10.385 $Y2=1.04
r30 12 13 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=10.292 $Y=2.24
+ $X2=10.292 $Y2=2.075
r31 2 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=10.14
+ $Y=2.095 $X2=10.28 $Y2=2.24
r32 1 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.14
+ $Y=0.33 $X2=10.28 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%VGND 1 2 3 4 5 17 19 20 21 24 28 32 36 39 42
+ 43 44 46 51 60 69 70 73 76 79
r128 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r129 76 77 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r130 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r131 70 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.36 $Y2=0
r132 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r133 67 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.6 $Y=0 $X2=9.435
+ $Y2=0
r134 67 69 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=9.6 $Y=0 $X2=10.32
+ $Y2=0
r135 66 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r136 65 66 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r137 63 66 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=6 $Y=0 $X2=8.88
+ $Y2=0
r138 62 65 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.88
+ $Y2=0
r139 62 63 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6
+ $Y2=0
r140 60 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.27 $Y=0 $X2=9.435
+ $Y2=0
r141 60 65 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.27 $Y=0 $X2=8.88
+ $Y2=0
r142 59 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r143 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r144 56 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=4.655
+ $Y2=0
r145 56 58 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=5.52
+ $Y2=0
r146 55 77 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=4.56 $Y2=0
r147 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r148 54 55 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r149 52 73 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.29
+ $Y2=0
r150 52 54 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.575 $Y=0
+ $X2=1.68 $Y2=0
r151 51 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.49 $Y=0 $X2=4.655
+ $Y2=0
r152 51 54 183.326 $w=1.68e-07 $l=2.81e-06 $layer=LI1_cond $X=4.49 $Y=0 $X2=1.68
+ $Y2=0
r153 49 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r154 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r155 46 73 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.29
+ $Y2=0
r156 46 48 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=0
+ $X2=0.72 $Y2=0
r157 44 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.52 $Y2=0
r158 44 77 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=4.56
+ $Y2=0
r159 42 58 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.52
+ $Y2=0
r160 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.755
+ $Y2=0
r161 41 62 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=5.92 $Y=0 $X2=6 $Y2=0
r162 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.92 $Y=0 $X2=5.755
+ $Y2=0
r163 39 40 11.325 $w=5.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.29 $Y=0.635
+ $X2=1.29 $Y2=0.865
r164 34 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.435 $Y=0.085
+ $X2=9.435 $Y2=0
r165 34 36 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=9.435 $Y=0.085
+ $X2=9.435 $Y2=0.54
r166 30 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0
r167 30 32 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0.85
r168 26 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.655 $Y=0.085
+ $X2=4.655 $Y2=0
r169 26 28 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.655 $Y=0.085
+ $X2=4.655 $Y2=0.485
r170 22 24 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.43 $Y=1.195
+ $X2=2.43 $Y2=0.915
r171 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.265 $Y=1.28
+ $X2=2.43 $Y2=1.195
r172 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.265 $Y=1.28
+ $X2=1.575 $Y2=1.28
r173 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.49 $Y=1.195
+ $X2=1.575 $Y2=1.28
r174 19 40 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.49 $Y=1.195
+ $X2=1.49 $Y2=0.865
r175 17 39 1.15411 $w=5.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.29 $Y=0.58
+ $X2=1.29 $Y2=0.635
r176 16 73 2.39972 $w=5.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.29 $Y=0.085
+ $X2=1.29 $Y2=0
r177 16 17 10.387 $w=5.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.29 $Y=0.085
+ $X2=1.29 $Y2=0.58
r178 5 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.295
+ $Y=0.33 $X2=9.435 $Y2=0.54
r179 4 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.615
+ $Y=0.705 $X2=5.755 $Y2=0.85
r180 3 28 182 $w=1.7e-07 $l=3.11127e-07 $layer=licon1_NDIFF $count=1 $X=4.435
+ $Y=0.705 $X2=4.655 $Y2=0.485
r181 2 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.29
+ $Y=0.705 $X2=2.43 $Y2=0.915
r182 1 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.425 $X2=1.17 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%A_355_141# 1 2 9 11 12 13
r37 13 16 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.065 $Y=0.405
+ $X2=4.065 $Y2=0.485
r38 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.9 $Y=0.405
+ $X2=4.065 $Y2=0.405
r39 11 12 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=3.9 $Y=0.405
+ $X2=2.085 $Y2=0.405
r40 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.92 $Y=0.49
+ $X2=2.085 $Y2=0.405
r41 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.92 $Y=0.49 $X2=1.92
+ $Y2=0.85
r42 2 16 182 $w=1.7e-07 $l=3.11127e-07 $layer=licon1_NDIFF $count=1 $X=3.845
+ $Y=0.705 $X2=4.065 $Y2=0.485
r43 1 9 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.705 $X2=1.92 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__FA_LP%A_1005_141# 1 2 8 9 10 11 14 17 22
c49 22 0 1.01679e-19 $X=7.58 $Y=0.85
r50 22 24 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.58 $Y=0.85
+ $X2=7.58 $Y2=0.935
r51 17 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.185 $Y=0.935
+ $X2=6.185 $Y2=1.2
r52 14 16 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.245 $Y=0.485
+ $X2=5.245 $Y2=0.65
r53 12 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=0.935
+ $X2=6.185 $Y2=0.935
r54 11 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.415 $Y=0.935
+ $X2=7.58 $Y2=0.935
r55 11 12 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=7.415 $Y=0.935
+ $X2=6.27 $Y2=0.935
r56 9 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.1 $Y=1.2 $X2=6.185
+ $Y2=1.2
r57 9 10 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.1 $Y=1.2 $X2=5.41
+ $Y2=1.2
r58 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.325 $Y=1.115
+ $X2=5.41 $Y2=1.2
r59 8 16 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.325 $Y=1.115
+ $X2=5.325 $Y2=0.65
r60 2 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.44
+ $Y=0.705 $X2=7.58 $Y2=0.85
r61 1 14 182 $w=1.7e-07 $l=3.11127e-07 $layer=licon1_NDIFF $count=1 $X=5.025
+ $Y=0.705 $X2=5.245 $Y2=0.485
.ends

