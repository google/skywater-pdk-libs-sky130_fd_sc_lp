* File: sky130_fd_sc_lp__and4_m.pxi.spice
* Created: Wed Sep  2 09:33:19 2020
* 
x_PM_SKY130_FD_SC_LP__AND4_M%A N_A_c_70_n N_A_M1002_g N_A_M1001_g N_A_c_66_n
+ N_A_c_67_n A A A N_A_c_69_n PM_SKY130_FD_SC_LP__AND4_M%A
x_PM_SKY130_FD_SC_LP__AND4_M%B N_B_M1008_g N_B_M1007_g N_B_c_99_n N_B_c_100_n
+ N_B_c_101_n B B B N_B_c_103_n PM_SKY130_FD_SC_LP__AND4_M%B
x_PM_SKY130_FD_SC_LP__AND4_M%C N_C_M1000_g N_C_M1009_g C C C N_C_c_141_n
+ PM_SKY130_FD_SC_LP__AND4_M%C
x_PM_SKY130_FD_SC_LP__AND4_M%D N_D_c_176_n N_D_M1003_g N_D_M1006_g N_D_c_177_n
+ N_D_c_178_n N_D_c_183_n D D D N_D_c_180_n N_D_c_181_n
+ PM_SKY130_FD_SC_LP__AND4_M%D
x_PM_SKY130_FD_SC_LP__AND4_M%A_53_47# N_A_53_47#_M1002_s N_A_53_47#_M1001_d
+ N_A_53_47#_M1009_d N_A_53_47#_c_232_n N_A_53_47#_c_227_n N_A_53_47#_M1005_g
+ N_A_53_47#_M1004_g N_A_53_47#_c_228_n N_A_53_47#_c_229_n N_A_53_47#_c_235_n
+ N_A_53_47#_c_230_n N_A_53_47#_c_231_n N_A_53_47#_c_237_n N_A_53_47#_c_238_n
+ N_A_53_47#_c_239_n N_A_53_47#_c_240_n N_A_53_47#_c_241_n
+ PM_SKY130_FD_SC_LP__AND4_M%A_53_47#
x_PM_SKY130_FD_SC_LP__AND4_M%VPWR N_VPWR_M1001_s N_VPWR_M1007_d N_VPWR_M1006_d
+ N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n
+ N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n VPWR N_VPWR_c_320_n
+ N_VPWR_c_311_n N_VPWR_c_322_n PM_SKY130_FD_SC_LP__AND4_M%VPWR
x_PM_SKY130_FD_SC_LP__AND4_M%X N_X_M1005_d N_X_M1004_d X X X X X X X
+ PM_SKY130_FD_SC_LP__AND4_M%X
x_PM_SKY130_FD_SC_LP__AND4_M%VGND N_VGND_M1003_d N_VGND_c_375_n VGND
+ N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n
+ PM_SKY130_FD_SC_LP__AND4_M%VGND
cc_1 VNB N_A_M1002_g 0.0317775f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.445
cc_2 VNB N_A_c_66_n 0.0382204f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.03
cc_3 VNB N_A_c_67_n 0.0257713f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_4 VNB A 0.00914588f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_A_c_69_n 0.0374549f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_6 VNB N_B_M1007_g 0.013453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B_c_99_n 0.0162506f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.165
cc_8 VNB N_B_c_100_n 0.0220991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B_c_101_n 0.0166688f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.03
cc_10 VNB B 0.00697333f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_11 VNB N_B_c_103_n 0.0153238f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_12 VNB N_C_M1000_g 0.0343811f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.955
cc_13 VNB N_C_M1009_g 0.00957975f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.825
cc_14 VNB C 0.00794126f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.165
cc_15 VNB N_C_c_141_n 0.0306856f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_16 VNB N_D_c_176_n 0.0168984f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.75
cc_17 VNB N_D_c_177_n 0.024403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_D_c_178_n 0.0114724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB D 0.00552695f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=1.75
cc_20 VNB N_D_c_180_n 0.0344888f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_21 VNB N_D_c_181_n 0.0127279f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_22 VNB N_A_53_47#_c_227_n 0.0204314f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_23 VNB N_A_53_47#_c_228_n 0.0416582f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_53_47#_c_229_n 0.0293002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_53_47#_c_230_n 0.0024911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_53_47#_c_231_n 0.0126184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_311_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB X 0.0418979f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.825
cc_29 VNB N_VGND_c_375_n 0.00561589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_376_n 0.0563958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_377_n 0.0197547f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_VGND_c_378_n 0.173548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_379_n 0.00631563f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_34 VPB N_A_c_70_n 0.0205986f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.75
cc_35 VPB N_A_M1001_g 0.0238753f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.165
cc_36 VPB N_A_c_67_n 0.0157563f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_37 VPB A 0.00858336f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_38 VPB N_B_M1007_g 0.0276637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_C_M1009_g 0.0275157f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.825
cc_40 VPB N_D_c_178_n 0.00258518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_D_c_183_n 0.0314063f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_42 VPB D 0.00229287f $X=-0.19 $Y=1.655 $X2=0.285 $Y2=1.75
cc_43 VPB N_A_53_47#_c_232_n 0.0423589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_53_47#_M1004_g 0.0369125f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_45 VPB N_A_53_47#_c_228_n 0.00173387f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_46 VPB N_A_53_47#_c_235_n 0.0298574f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_47 VPB N_A_53_47#_c_231_n 9.11941e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_53_47#_c_237_n 0.00176211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_53_47#_c_238_n 0.0203614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_53_47#_c_239_n 0.00626031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_53_47#_c_240_n 0.00955773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_53_47#_c_241_n 0.0430678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_312_n 0.0449512f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.105
cc_54 VPB N_VPWR_c_313_n 0.0250293f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_55 VPB N_VPWR_c_314_n 0.0187753f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_56 VPB N_VPWR_c_315_n 0.0157197f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_316_n 0.0137583f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_58 VPB N_VPWR_c_317_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_59 VPB N_VPWR_c_318_n 0.0206207f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_60 VPB N_VPWR_c_319_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_320_n 0.0194756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_311_n 0.0943009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_322_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB X 0.0379663f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.825
cc_65 N_A_c_70_n N_B_M1007_g 0.0204996f $X=0.61 $Y=1.75 $X2=0 $Y2=0
cc_66 N_A_c_69_n N_B_M1007_g 0.00178674f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_67 N_A_M1002_g N_B_c_99_n 0.0308208f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_c_69_n N_B_c_100_n 0.00466214f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_69 N_A_M1002_g B 5.72162e-19 $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_c_66_n N_B_c_103_n 0.0308208f $X=0.605 $Y=1.03 $X2=0 $Y2=0
cc_71 N_A_M1002_g N_A_53_47#_c_230_n 0.0118151f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A_c_66_n N_A_53_47#_c_230_n 0.00660503f $X=0.605 $Y=1.03 $X2=0 $Y2=0
cc_73 A N_A_53_47#_c_230_n 0.00568174f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_74 N_A_c_70_n N_A_53_47#_c_231_n 0.00496269f $X=0.61 $Y=1.75 $X2=0 $Y2=0
cc_75 N_A_M1002_g N_A_53_47#_c_231_n 0.0108594f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A_c_66_n N_A_53_47#_c_231_n 0.0052689f $X=0.605 $Y=1.03 $X2=0 $Y2=0
cc_77 A N_A_53_47#_c_231_n 0.0447027f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_78 N_A_c_69_n N_A_53_47#_c_231_n 0.0037735f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_79 N_A_M1001_g N_A_53_47#_c_237_n 0.00178215f $X=0.685 $Y=2.165 $X2=0 $Y2=0
cc_80 N_A_c_70_n N_A_53_47#_c_239_n 0.00734226f $X=0.61 $Y=1.75 $X2=0 $Y2=0
cc_81 N_A_M1001_g N_A_53_47#_c_239_n 0.00990377f $X=0.685 $Y=2.165 $X2=0 $Y2=0
cc_82 A N_A_53_47#_c_239_n 0.00183402f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_83 N_A_M1001_g N_VPWR_c_312_n 0.0037597f $X=0.685 $Y=2.165 $X2=0 $Y2=0
cc_84 N_A_c_67_n N_VPWR_c_312_n 0.0079099f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_85 N_A_M1001_g N_VPWR_c_311_n 0.00387136f $X=0.685 $Y=2.165 $X2=0 $Y2=0
cc_86 N_A_M1002_g N_VGND_c_376_n 0.00372993f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_VGND_c_378_n 0.0064053f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_88 A N_VGND_c_378_n 0.00522088f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_B_c_99_n N_C_M1000_g 0.0201679f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_90 B N_C_M1000_g 0.00665318f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_91 N_B_c_103_n N_C_M1000_g 0.0201676f $X=1.055 $Y=0.93 $X2=0 $Y2=0
cc_92 N_B_M1007_g N_C_M1009_g 0.0294204f $X=1.115 $Y=2.165 $X2=0 $Y2=0
cc_93 N_B_M1007_g C 2.70255e-19 $X=1.115 $Y=2.165 $X2=0 $Y2=0
cc_94 N_B_c_99_n C 2.44242e-19 $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_95 B C 0.0602636f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_96 N_B_c_103_n C 6.64353e-19 $X=1.055 $Y=0.93 $X2=0 $Y2=0
cc_97 N_B_M1007_g N_C_c_141_n 0.00266356f $X=1.115 $Y=2.165 $X2=0 $Y2=0
cc_98 N_B_c_100_n N_C_c_141_n 0.0201676f $X=1.055 $Y=1.27 $X2=0 $Y2=0
cc_99 N_B_c_99_n N_A_53_47#_c_230_n 0.00500134f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_100 B N_A_53_47#_c_230_n 0.0146193f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_101 N_B_M1007_g N_A_53_47#_c_231_n 0.0067903f $X=1.115 $Y=2.165 $X2=0 $Y2=0
cc_102 N_B_c_99_n N_A_53_47#_c_231_n 0.00720069f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_103 B N_A_53_47#_c_231_n 0.0554444f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_104 N_B_M1007_g N_A_53_47#_c_237_n 9.6003e-19 $X=1.115 $Y=2.165 $X2=0 $Y2=0
cc_105 N_B_M1007_g N_A_53_47#_c_238_n 0.0153629f $X=1.115 $Y=2.165 $X2=0 $Y2=0
cc_106 N_B_c_101_n N_A_53_47#_c_239_n 0.00341896f $X=1.055 $Y=1.435 $X2=0 $Y2=0
cc_107 B N_A_53_47#_c_239_n 0.0168776f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_108 N_B_M1007_g N_VPWR_c_313_n 0.00178443f $X=1.115 $Y=2.165 $X2=0 $Y2=0
cc_109 N_B_M1007_g N_VPWR_c_311_n 0.00387136f $X=1.115 $Y=2.165 $X2=0 $Y2=0
cc_110 B A_208_47# 0.00487949f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_111 N_B_c_99_n N_VGND_c_376_n 0.00499463f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_112 B N_VGND_c_376_n 0.00818334f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_113 N_B_c_103_n N_VGND_c_376_n 4.83856e-19 $X=1.055 $Y=0.93 $X2=0 $Y2=0
cc_114 N_B_c_99_n N_VGND_c_378_n 0.00865283f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_115 B N_VGND_c_378_n 0.010346f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_116 N_C_M1000_g N_D_c_176_n 0.0498735f $X=1.505 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_117 C N_D_c_176_n 0.00613266f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_118 N_C_M1009_g N_D_c_178_n 0.00750558f $X=1.545 $Y=2.165 $X2=0 $Y2=0
cc_119 N_C_M1009_g N_D_c_183_n 0.0176165f $X=1.545 $Y=2.165 $X2=0 $Y2=0
cc_120 N_C_M1000_g D 2.67896e-19 $X=1.505 $Y=0.445 $X2=0 $Y2=0
cc_121 N_C_M1009_g D 0.00119756f $X=1.545 $Y=2.165 $X2=0 $Y2=0
cc_122 C D 0.0327199f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_123 N_C_c_141_n D 3.69411e-19 $X=1.595 $Y=1.32 $X2=0 $Y2=0
cc_124 N_C_c_141_n N_D_c_180_n 0.0206146f $X=1.595 $Y=1.32 $X2=0 $Y2=0
cc_125 N_C_M1000_g N_D_c_181_n 0.00616855f $X=1.505 $Y=0.445 $X2=0 $Y2=0
cc_126 C N_D_c_181_n 0.00399968f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_127 N_C_M1009_g N_A_53_47#_c_238_n 0.0158705f $X=1.545 $Y=2.165 $X2=0 $Y2=0
cc_128 C N_A_53_47#_c_238_n 0.0164637f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_129 N_C_c_141_n N_A_53_47#_c_238_n 0.00258624f $X=1.595 $Y=1.32 $X2=0 $Y2=0
cc_130 N_C_M1009_g N_A_53_47#_c_240_n 0.00236435f $X=1.545 $Y=2.165 $X2=0 $Y2=0
cc_131 N_C_M1009_g N_A_53_47#_c_241_n 3.89852e-19 $X=1.545 $Y=2.165 $X2=0 $Y2=0
cc_132 N_C_M1009_g N_VPWR_c_313_n 0.00106626f $X=1.545 $Y=2.165 $X2=0 $Y2=0
cc_133 N_C_M1009_g N_VPWR_c_311_n 0.00374993f $X=1.545 $Y=2.165 $X2=0 $Y2=0
cc_134 C A_316_47# 0.00139886f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_135 N_C_M1000_g N_VGND_c_376_n 0.00499463f $X=1.505 $Y=0.445 $X2=0 $Y2=0
cc_136 C N_VGND_c_376_n 0.00603051f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_137 N_C_M1000_g N_VGND_c_378_n 0.00865283f $X=1.505 $Y=0.445 $X2=0 $Y2=0
cc_138 C N_VGND_c_378_n 0.00829629f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_139 N_D_c_183_n N_A_53_47#_c_232_n 0.00412877f $X=2.01 $Y=1.845 $X2=0 $Y2=0
cc_140 N_D_c_176_n N_A_53_47#_c_227_n 0.0138055f $X=1.865 $Y=0.765 $X2=0 $Y2=0
cc_141 N_D_c_183_n N_A_53_47#_M1004_g 0.0123852f $X=2.01 $Y=1.845 $X2=0 $Y2=0
cc_142 N_D_c_178_n N_A_53_47#_c_228_n 0.00383748f $X=2.01 $Y=1.695 $X2=0 $Y2=0
cc_143 D N_A_53_47#_c_228_n 0.00135304f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_144 N_D_c_180_n N_A_53_47#_c_228_n 0.017457f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_145 N_D_c_181_n N_A_53_47#_c_228_n 0.00306742f $X=2.135 $Y=1.125 $X2=0 $Y2=0
cc_146 N_D_c_177_n N_A_53_47#_c_229_n 0.00971476f $X=2.045 $Y=0.84 $X2=0 $Y2=0
cc_147 D N_A_53_47#_c_229_n 5.8615e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_148 N_D_c_183_n N_A_53_47#_c_235_n 0.0095338f $X=2.01 $Y=1.845 $X2=0 $Y2=0
cc_149 D N_A_53_47#_c_235_n 4.29844e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_150 N_D_c_183_n N_A_53_47#_c_238_n 0.00263547f $X=2.01 $Y=1.845 $X2=0 $Y2=0
cc_151 D N_A_53_47#_c_238_n 0.00267358f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_152 N_D_c_183_n N_A_53_47#_c_240_n 0.00236435f $X=2.01 $Y=1.845 $X2=0 $Y2=0
cc_153 N_D_c_183_n N_A_53_47#_c_241_n 0.00350866f $X=2.01 $Y=1.845 $X2=0 $Y2=0
cc_154 N_D_c_183_n N_VPWR_c_315_n 0.00190847f $X=2.01 $Y=1.845 $X2=0 $Y2=0
cc_155 D N_VPWR_c_315_n 0.00855762f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_156 N_D_c_180_n N_VPWR_c_315_n 0.00162416f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_157 N_D_c_177_n X 4.21557e-19 $X=2.045 $Y=0.84 $X2=0 $Y2=0
cc_158 N_D_c_178_n X 9.04968e-19 $X=2.01 $Y=1.695 $X2=0 $Y2=0
cc_159 N_D_c_183_n X 3.1027e-19 $X=2.01 $Y=1.845 $X2=0 $Y2=0
cc_160 D X 0.0491651f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_161 N_D_c_180_n X 0.0021123f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_162 N_D_c_181_n X 8.15648e-19 $X=2.135 $Y=1.125 $X2=0 $Y2=0
cc_163 N_D_c_176_n N_VGND_c_375_n 0.0033813f $X=1.865 $Y=0.765 $X2=0 $Y2=0
cc_164 N_D_c_177_n N_VGND_c_375_n 0.0050014f $X=2.045 $Y=0.84 $X2=0 $Y2=0
cc_165 D N_VGND_c_375_n 0.00880495f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_166 N_D_c_180_n N_VGND_c_375_n 0.00131241f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_167 N_D_c_176_n N_VGND_c_376_n 0.00585385f $X=1.865 $Y=0.765 $X2=0 $Y2=0
cc_168 N_D_c_176_n N_VGND_c_378_n 0.0107161f $X=1.865 $Y=0.765 $X2=0 $Y2=0
cc_169 D N_VGND_c_378_n 0.00100324f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_170 N_A_53_47#_c_238_n N_VPWR_c_313_n 0.0146902f $X=1.655 $Y=1.8 $X2=0 $Y2=0
cc_171 N_A_53_47#_c_240_n N_VPWR_c_313_n 0.0421044f $X=1.76 $Y=2.23 $X2=0 $Y2=0
cc_172 N_A_53_47#_c_241_n N_VPWR_c_313_n 0.00813147f $X=1.78 $Y=2.88 $X2=0 $Y2=0
cc_173 N_A_53_47#_c_240_n N_VPWR_c_314_n 0.0118318f $X=1.76 $Y=2.23 $X2=0 $Y2=0
cc_174 N_A_53_47#_c_241_n N_VPWR_c_314_n 0.00934322f $X=1.78 $Y=2.88 $X2=0 $Y2=0
cc_175 N_A_53_47#_c_232_n N_VPWR_c_315_n 0.020683f $X=2.33 $Y=2.97 $X2=0 $Y2=0
cc_176 N_A_53_47#_M1004_g N_VPWR_c_315_n 0.00831371f $X=2.405 $Y=2.165 $X2=0
+ $Y2=0
cc_177 N_A_53_47#_c_240_n N_VPWR_c_315_n 0.0415105f $X=1.76 $Y=2.23 $X2=0 $Y2=0
cc_178 N_A_53_47#_c_241_n N_VPWR_c_315_n 0.00156514f $X=1.78 $Y=2.88 $X2=0 $Y2=0
cc_179 N_A_53_47#_c_232_n N_VPWR_c_320_n 0.00644723f $X=2.33 $Y=2.97 $X2=0 $Y2=0
cc_180 N_A_53_47#_c_240_n N_VPWR_c_311_n 0.00782891f $X=1.76 $Y=2.23 $X2=0 $Y2=0
cc_181 N_A_53_47#_c_241_n N_VPWR_c_311_n 0.0141207f $X=1.78 $Y=2.88 $X2=0 $Y2=0
cc_182 N_A_53_47#_c_227_n X 0.00443413f $X=2.405 $Y=0.765 $X2=0 $Y2=0
cc_183 N_A_53_47#_M1004_g X 0.0160841f $X=2.405 $Y=2.165 $X2=0 $Y2=0
cc_184 N_A_53_47#_c_228_n X 0.0250247f $X=2.615 $Y=1.695 $X2=0 $Y2=0
cc_185 N_A_53_47#_c_229_n X 0.0110274f $X=2.615 $Y=0.84 $X2=0 $Y2=0
cc_186 N_A_53_47#_c_235_n X 0.0119352f $X=2.615 $Y=1.77 $X2=0 $Y2=0
cc_187 N_A_53_47#_c_238_n X 0.00410016f $X=1.655 $Y=1.8 $X2=0 $Y2=0
cc_188 N_A_53_47#_c_240_n X 0.00204746f $X=1.76 $Y=2.23 $X2=0 $Y2=0
cc_189 N_A_53_47#_c_230_n A_136_47# 0.0039738f $X=0.62 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_190 N_A_53_47#_c_227_n N_VGND_c_375_n 0.00445728f $X=2.405 $Y=0.765 $X2=0
+ $Y2=0
cc_191 N_A_53_47#_c_230_n N_VGND_c_376_n 0.0203008f $X=0.62 $Y=0.495 $X2=0 $Y2=0
cc_192 N_A_53_47#_c_227_n N_VGND_c_377_n 0.00585385f $X=2.405 $Y=0.765 $X2=0
+ $Y2=0
cc_193 N_A_53_47#_c_229_n N_VGND_c_377_n 9.75559e-19 $X=2.615 $Y=0.84 $X2=0
+ $Y2=0
cc_194 N_A_53_47#_M1002_s N_VGND_c_378_n 0.00234684f $X=0.265 $Y=0.235 $X2=0
+ $Y2=0
cc_195 N_A_53_47#_c_227_n N_VGND_c_378_n 0.0121529f $X=2.405 $Y=0.765 $X2=0
+ $Y2=0
cc_196 N_A_53_47#_c_229_n N_VGND_c_378_n 7.6639e-19 $X=2.615 $Y=0.84 $X2=0 $Y2=0
cc_197 N_A_53_47#_c_230_n N_VGND_c_378_n 0.0178558f $X=0.62 $Y=0.495 $X2=0 $Y2=0
cc_198 N_VPWR_c_315_n X 0.0313828f $X=2.19 $Y=2.23 $X2=0 $Y2=0
cc_199 N_VPWR_c_320_n X 0.00623633f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_200 N_VPWR_c_311_n X 0.00710559f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_201 X N_VGND_c_377_n 0.00877924f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_202 N_X_M1005_d N_VGND_c_378_n 0.00337555f $X=2.48 $Y=0.235 $X2=0 $Y2=0
cc_203 X N_VGND_c_378_n 0.00770513f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_204 A_136_47# N_VGND_c_378_n 0.00519157f $X=0.68 $Y=0.235 $X2=2.405 $Y2=0.84
cc_205 A_208_47# N_VGND_c_378_n 0.00856878f $X=1.04 $Y=0.235 $X2=1.127 $Y2=0.555
cc_206 A_316_47# N_VGND_c_378_n 0.00285223f $X=1.58 $Y=0.235 $X2=0 $Y2=0
