* File: sky130_fd_sc_lp__clkbuflp_8.pex.spice
* Created: Fri Aug 28 10:16:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_8%A 3 7 11 15 19 23 27 31 33 34 42 48
c76 42 0 4.25933e-20 $X=0.565 $Y=1.4
r77 50 57 2.77751 $w=3e-07 $l=2.13e-07 $layer=LI1_cond $X=0.275 $Y=1.565
+ $X2=0.275 $Y2=1.352
r78 47 48 85.682 $w=3.3e-07 $l=4.9e-07 $layer=POLY_cond $X=1.625 $Y=1.4
+ $X2=2.115 $Y2=1.4
r79 46 47 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.585 $Y=1.4 $X2=1.625
+ $Y2=1.4
r80 45 46 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=1.265 $Y=1.4
+ $X2=1.585 $Y2=1.4
r81 44 45 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.055 $Y=1.4
+ $X2=1.265 $Y2=1.4
r82 43 44 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.835 $Y=1.4
+ $X2=1.055 $Y2=1.4
r83 42 57 7.86373 $w=4.23e-07 $l=2.9e-07 $layer=LI1_cond $X=0.565 $Y=1.352
+ $X2=0.275 $Y2=1.352
r84 41 43 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.565 $Y=1.4
+ $X2=0.835 $Y2=1.4
r85 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.565
+ $Y=1.4 $X2=0.565 $Y2=1.4
r86 39 41 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.525 $Y=1.4 $X2=0.565
+ $Y2=1.4
r87 37 39 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.475 $Y=1.4 $X2=0.525
+ $Y2=1.4
r88 34 50 3.84148 $w=2.98e-07 $l=1e-07 $layer=LI1_cond $X=0.275 $Y=1.665
+ $X2=0.275 $Y2=1.565
r89 33 57 0.949071 $w=4.23e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.352
+ $X2=0.275 $Y2=1.352
r90 29 48 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.115 $Y=1.565
+ $X2=2.115 $Y2=1.4
r91 29 31 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.115 $Y=1.565
+ $X2=2.115 $Y2=2.585
r92 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=1.4
r93 25 27 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=0.555
r94 21 46 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.565
+ $X2=1.585 $Y2=1.4
r95 21 23 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.585 $Y=1.565
+ $X2=1.585 $Y2=2.585
r96 17 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.235
+ $X2=1.265 $Y2=1.4
r97 17 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.265 $Y=1.235
+ $X2=1.265 $Y2=0.555
r98 13 44 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.565
+ $X2=1.055 $Y2=1.4
r99 13 15 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.055 $Y=1.565
+ $X2=1.055 $Y2=2.585
r100 9 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=1.4
r101 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=0.555
r102 5 39 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.565
+ $X2=0.525 $Y2=1.4
r103 5 7 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=0.525 $Y=1.565
+ $X2=0.525 $Y2=2.585
r104 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=1.4
r105 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_8%A_130_417# 1 2 3 12 16 20 24 28 32 36 40
+ 44 48 52 56 60 64 68 72 76 82 85 88 92 97 103 121
r192 120 121 89.9507 $w=3.4e-07 $l=5.3e-07 $layer=POLY_cond $X=5.825 $Y=1.375
+ $X2=6.355 $Y2=1.375
r193 119 120 84.8592 $w=3.4e-07 $l=5e-07 $layer=POLY_cond $X=5.325 $Y=1.375
+ $X2=5.825 $Y2=1.375
r194 118 119 5.09155 $w=3.4e-07 $l=3e-08 $layer=POLY_cond $X=5.295 $Y=1.375
+ $X2=5.325 $Y2=1.375
r195 117 118 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=4.965 $Y=1.375
+ $X2=5.295 $Y2=1.375
r196 116 117 33.9437 $w=3.4e-07 $l=2e-07 $layer=POLY_cond $X=4.765 $Y=1.375
+ $X2=4.965 $Y2=1.375
r197 115 116 39.0352 $w=3.4e-07 $l=2.3e-07 $layer=POLY_cond $X=4.535 $Y=1.375
+ $X2=4.765 $Y2=1.375
r198 114 115 50.9155 $w=3.4e-07 $l=3e-07 $layer=POLY_cond $X=4.235 $Y=1.375
+ $X2=4.535 $Y2=1.375
r199 113 114 10.1831 $w=3.4e-07 $l=6e-08 $layer=POLY_cond $X=4.175 $Y=1.375
+ $X2=4.235 $Y2=1.375
r200 112 113 72.9789 $w=3.4e-07 $l=4.3e-07 $layer=POLY_cond $X=3.745 $Y=1.375
+ $X2=4.175 $Y2=1.375
r201 109 110 35.6408 $w=3.4e-07 $l=2.1e-07 $layer=POLY_cond $X=3.175 $Y=1.375
+ $X2=3.385 $Y2=1.375
r202 108 109 37.338 $w=3.4e-07 $l=2.2e-07 $layer=POLY_cond $X=2.955 $Y=1.375
+ $X2=3.175 $Y2=1.375
r203 104 106 8.48592 $w=3.4e-07 $l=5e-08 $layer=POLY_cond $X=2.595 $Y=1.375
+ $X2=2.645 $Y2=1.375
r204 101 102 14.995 $w=5.98e-07 $l=7.35e-07 $layer=LI1_cond $X=1.092 $Y=1.572
+ $X2=1.827 $Y2=1.572
r205 98 112 6.78873 $w=3.4e-07 $l=4e-08 $layer=POLY_cond $X=3.705 $Y=1.375
+ $X2=3.745 $Y2=1.375
r206 98 110 54.3099 $w=3.4e-07 $l=3.2e-07 $layer=POLY_cond $X=3.705 $Y=1.375
+ $X2=3.385 $Y2=1.375
r207 97 98 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.705
+ $Y=1.37 $X2=3.705 $Y2=1.37
r208 95 108 45.8239 $w=3.4e-07 $l=2.7e-07 $layer=POLY_cond $X=2.685 $Y=1.375
+ $X2=2.955 $Y2=1.375
r209 95 106 6.78873 $w=3.4e-07 $l=4e-08 $layer=POLY_cond $X=2.685 $Y=1.375
+ $X2=2.645 $Y2=1.375
r210 94 97 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=2.685 $Y=1.37
+ $X2=3.705 $Y2=1.37
r211 94 95 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.685
+ $Y=1.37 $X2=2.685 $Y2=1.37
r212 92 102 5.8593 $w=5.98e-07 $l=2.73386e-07 $layer=LI1_cond $X=1.995 $Y=1.37
+ $X2=1.827 $Y2=1.572
r213 92 94 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=1.995 $Y=1.37
+ $X2=2.685 $Y2=1.37
r214 88 90 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=1.827 $Y=2.23
+ $X2=1.827 $Y2=2.91
r215 86 102 4.1387 $w=3.35e-07 $l=3.68e-07 $layer=LI1_cond $X=1.827 $Y=1.94
+ $X2=1.827 $Y2=1.572
r216 86 88 9.97637 $w=3.33e-07 $l=2.9e-07 $layer=LI1_cond $X=1.827 $Y=1.94
+ $X2=1.827 $Y2=2.23
r217 85 101 5.31194 $w=2.75e-07 $l=3.67e-07 $layer=LI1_cond $X=1.092 $Y=1.205
+ $X2=1.092 $Y2=1.572
r218 85 103 9.21954 $w=2.73e-07 $l=2.2e-07 $layer=LI1_cond $X=1.092 $Y=1.205
+ $X2=1.092 $Y2=0.985
r219 80 103 6.25289 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=1.057 $Y=0.813
+ $X2=1.057 $Y2=0.985
r220 80 82 14.297 $w=3.43e-07 $l=4.28e-07 $layer=LI1_cond $X=1.057 $Y=0.813
+ $X2=1.057 $Y2=0.385
r221 76 78 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.79 $Y=2.23
+ $X2=0.79 $Y2=2.91
r222 74 101 6.1612 $w=5.98e-07 $l=4.96548e-07 $layer=LI1_cond $X=0.79 $Y=1.94
+ $X2=1.092 $Y2=1.572
r223 74 76 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.79 $Y=1.94
+ $X2=0.79 $Y2=2.23
r224 70 121 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.355 $Y=1.545
+ $X2=6.355 $Y2=1.375
r225 70 72 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=6.355 $Y=1.545
+ $X2=6.355 $Y2=2.585
r226 66 120 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.825 $Y=1.545
+ $X2=5.825 $Y2=1.375
r227 66 68 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=5.825 $Y=1.545
+ $X2=5.825 $Y2=2.585
r228 62 119 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.325 $Y=1.205
+ $X2=5.325 $Y2=1.375
r229 62 64 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.325 $Y=1.205
+ $X2=5.325 $Y2=0.51
r230 58 118 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.295 $Y=1.545
+ $X2=5.295 $Y2=1.375
r231 58 60 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=5.295 $Y=1.545
+ $X2=5.295 $Y2=2.585
r232 54 117 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.965 $Y=1.205
+ $X2=4.965 $Y2=1.375
r233 54 56 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=4.965 $Y=1.205
+ $X2=4.965 $Y2=0.51
r234 50 116 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.765 $Y=1.545
+ $X2=4.765 $Y2=1.375
r235 50 52 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=4.765 $Y=1.545
+ $X2=4.765 $Y2=2.585
r236 46 115 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.535 $Y=1.205
+ $X2=4.535 $Y2=1.375
r237 46 48 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=4.535 $Y=1.205
+ $X2=4.535 $Y2=0.51
r238 42 114 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.235 $Y=1.545
+ $X2=4.235 $Y2=1.375
r239 42 44 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=4.235 $Y=1.545
+ $X2=4.235 $Y2=2.585
r240 38 113 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.175 $Y=1.205
+ $X2=4.175 $Y2=1.375
r241 38 40 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=4.175 $Y=1.205
+ $X2=4.175 $Y2=0.51
r242 34 112 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.745 $Y=1.205
+ $X2=3.745 $Y2=1.375
r243 34 36 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.745 $Y=1.205
+ $X2=3.745 $Y2=0.51
r244 30 98 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.705 $Y=1.545
+ $X2=3.705 $Y2=1.375
r245 30 32 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=3.705 $Y=1.545
+ $X2=3.705 $Y2=2.585
r246 26 110 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.385 $Y=1.205
+ $X2=3.385 $Y2=1.375
r247 26 28 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.385 $Y=1.205
+ $X2=3.385 $Y2=0.51
r248 22 109 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.175 $Y=1.545
+ $X2=3.175 $Y2=1.375
r249 22 24 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=3.175 $Y=1.545
+ $X2=3.175 $Y2=2.585
r250 18 108 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.955 $Y=1.205
+ $X2=2.955 $Y2=1.375
r251 18 20 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.955 $Y=1.205
+ $X2=2.955 $Y2=0.51
r252 14 106 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.645 $Y=1.545
+ $X2=2.645 $Y2=1.375
r253 14 16 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.645 $Y=1.545
+ $X2=2.645 $Y2=2.585
r254 10 104 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.595 $Y=1.205
+ $X2=2.595 $Y2=1.375
r255 10 12 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.595 $Y=1.205
+ $X2=2.595 $Y2=0.51
r256 3 90 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.085 $X2=1.85 $Y2=2.91
r257 3 88 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.085 $X2=1.85 $Y2=2.23
r258 2 78 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.085 $X2=0.79 $Y2=2.91
r259 2 76 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.085 $X2=0.79 $Y2=2.23
r260 1 82 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.235 $X2=1.05 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_8%VPWR 1 2 3 4 5 6 7 22 24 28 32 38 44 50
+ 56 60 64 69 70 72 73 74 83 87 94 95 101 104 107 110
c111 24 0 4.25933e-20 $X=0.26 $Y=2.23
r112 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r113 108 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r115 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r117 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r119 95 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r120 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 92 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=3.33
+ $X2=6.62 $Y2=3.33
r122 92 94 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.785 $Y=3.33
+ $X2=6.96 $Y2=3.33
r123 91 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r124 91 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r126 88 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=4.5 $Y2=3.33
r127 88 90 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=5.04 $Y2=3.33
r128 87 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.56 $Y2=3.33
r129 87 90 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.04 $Y2=3.33
r130 86 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r131 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 83 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.5 $Y2=3.33
r133 83 85 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r135 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r136 79 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r137 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 76 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.32 $Y2=3.33
r139 76 78 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r140 74 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r141 74 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r142 72 81 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.12 $Y2=3.33
r143 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.44 $Y2=3.33
r144 71 85 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 71 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.44 $Y2=3.33
r146 69 78 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.16 $Y2=3.33
r147 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.38 $Y2=3.33
r148 68 81 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=3.12 $Y2=3.33
r149 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.38 $Y2=3.33
r150 64 67 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.62 $Y=2.23
+ $X2=6.62 $Y2=2.91
r151 62 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.62 $Y=3.245
+ $X2=6.62 $Y2=3.33
r152 62 67 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.62 $Y=3.245
+ $X2=6.62 $Y2=2.91
r153 61 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=3.33
+ $X2=5.56 $Y2=3.33
r154 60 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.455 $Y=3.33
+ $X2=6.62 $Y2=3.33
r155 60 61 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.455 $Y=3.33
+ $X2=5.725 $Y2=3.33
r156 56 59 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.56 $Y=2.23
+ $X2=5.56 $Y2=2.91
r157 54 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.56 $Y=3.245
+ $X2=5.56 $Y2=3.33
r158 54 59 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.56 $Y=3.245
+ $X2=5.56 $Y2=2.91
r159 50 53 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.5 $Y=2.23 $X2=4.5
+ $Y2=2.91
r160 48 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=3.245
+ $X2=4.5 $Y2=3.33
r161 48 53 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.5 $Y=3.245
+ $X2=4.5 $Y2=2.91
r162 44 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.44 $Y=2.23
+ $X2=3.44 $Y2=2.91
r163 42 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=3.33
r164 42 47 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=2.91
r165 38 41 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.38 $Y=2.23
+ $X2=2.38 $Y2=2.91
r166 36 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=3.33
r167 36 41 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=2.91
r168 32 35 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.32 $Y=2.23
+ $X2=1.32 $Y2=2.91
r169 30 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=3.245
+ $X2=1.32 $Y2=3.33
r170 30 35 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.32 $Y=3.245
+ $X2=1.32 $Y2=2.91
r171 29 98 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r172 28 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.32 $Y2=3.33
r173 28 29 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=0.425 $Y2=3.33
r174 24 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.23
+ $X2=0.26 $Y2=2.91
r175 22 98 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r176 22 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.91
r177 7 67 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=2.085 $X2=6.62 $Y2=2.91
r178 7 64 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=2.085 $X2=6.62 $Y2=2.23
r179 6 59 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=2.085 $X2=5.56 $Y2=2.91
r180 6 56 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=2.085 $X2=5.56 $Y2=2.23
r181 5 53 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.085 $X2=4.5 $Y2=2.91
r182 5 50 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.085 $X2=4.5 $Y2=2.23
r183 4 47 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=2.085 $X2=3.44 $Y2=2.91
r184 4 44 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=2.085 $X2=3.44 $Y2=2.23
r185 3 41 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=2.085 $X2=2.38 $Y2=2.91
r186 3 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=2.085 $X2=2.38 $Y2=2.23
r187 2 35 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=2.085 $X2=1.32 $Y2=2.91
r188 2 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=2.085 $X2=1.32 $Y2=2.23
r189 1 27 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.085 $X2=0.26 $Y2=2.91
r190 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.085 $X2=0.26 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_8%X 1 2 3 4 5 6 21 27 29 30 32 35 41 45 51
+ 55 57 59 60 61 79 80
r116 93 94 3.75609 $w=8.38e-07 $l=2.58e-07 $layer=LI1_cond $X=4.772 $Y=1.33
+ $X2=5.03 $Y2=1.33
r117 61 79 1.19478 $w=6.2e-07 $l=4.3e-07 $layer=LI1_cond $X=6.305 $Y=1.48
+ $X2=5.875 $Y2=1.48
r118 61 84 5.34532 $w=5.95e-07 $l=3.1e-07 $layer=LI1_cond $X=6.305 $Y=1.48
+ $X2=6.305 $Y2=1.17
r119 60 84 3.47558 $w=8.58e-07 $l=2.45e-07 $layer=LI1_cond $X=6.305 $Y=0.925
+ $X2=6.305 $Y2=1.17
r120 59 60 5.24884 $w=8.58e-07 $l=3.7e-07 $layer=LI1_cond $X=6.305 $Y=0.555
+ $X2=6.305 $Y2=0.925
r121 57 79 6.84851 $w=6.18e-07 $l=3.55e-07 $layer=LI1_cond $X=5.52 $Y=1.48
+ $X2=5.875 $Y2=1.48
r122 57 80 6.26977 $w=6.18e-07 $l=3.25e-07 $layer=LI1_cond $X=5.52 $Y=1.48
+ $X2=5.195 $Y2=1.48
r123 55 80 3.10719 $w=8.38e-07 $l=2.17428e-07 $layer=LI1_cond $X=5.04 $Y=1.33
+ $X2=5.195 $Y2=1.48
r124 55 94 0.145585 $w=8.38e-07 $l=1e-08 $layer=LI1_cond $X=5.04 $Y=1.33
+ $X2=5.03 $Y2=1.33
r125 51 53 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.09 $Y=2.23
+ $X2=6.09 $Y2=2.91
r126 49 61 5.34532 $w=5.95e-07 $l=4.03423e-07 $layer=LI1_cond $X=6.09 $Y=1.79
+ $X2=6.305 $Y2=1.48
r127 49 51 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=6.09 $Y=1.79
+ $X2=6.09 $Y2=2.23
r128 45 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.03 $Y=2.23
+ $X2=5.03 $Y2=2.91
r129 43 94 6.24443 $w=3.3e-07 $l=5.45e-07 $layer=LI1_cond $X=5.03 $Y=1.875
+ $X2=5.03 $Y2=1.33
r130 43 45 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.03 $Y=1.875
+ $X2=5.03 $Y2=2.23
r131 39 93 5.47333 $w=3.75e-07 $l=5.55e-07 $layer=LI1_cond $X=4.772 $Y=0.775
+ $X2=4.772 $Y2=1.33
r132 39 41 8.14393 $w=3.73e-07 $l=2.65e-07 $layer=LI1_cond $X=4.772 $Y=0.775
+ $X2=4.772 $Y2=0.51
r133 35 37 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.97 $Y=2.23
+ $X2=3.97 $Y2=2.91
r134 33 93 11.6759 $w=8.38e-07 $l=1.04322e-06 $layer=LI1_cond $X=3.97 $Y=1.885
+ $X2=4.772 $Y2=1.33
r135 33 35 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.97 $Y=1.885
+ $X2=3.97 $Y2=2.23
r136 29 33 8.23375 $w=8.38e-07 $l=1.04298e-06 $layer=LI1_cond $X=4.1 $Y=0.905
+ $X2=3.97 $Y2=1.885
r137 29 32 33.9084 $w=2.58e-07 $l=7.65e-07 $layer=LI1_cond $X=4.1 $Y=0.905
+ $X2=3.335 $Y2=0.905
r138 29 30 44.9798 $w=1.78e-07 $l=7.3e-07 $layer=LI1_cond $X=3.805 $Y=1.795
+ $X2=3.075 $Y2=1.795
r139 25 32 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=3.17 $Y=0.775
+ $X2=3.335 $Y2=0.905
r140 25 27 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.17 $Y=0.775
+ $X2=3.17 $Y2=0.51
r141 21 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.91 $Y=2.23
+ $X2=2.91 $Y2=2.91
r142 19 30 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.91 $Y=1.885
+ $X2=3.075 $Y2=1.795
r143 19 21 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.91 $Y=1.885
+ $X2=2.91 $Y2=2.23
r144 6 53 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=5.95
+ $Y=2.085 $X2=6.09 $Y2=2.91
r145 6 51 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.95
+ $Y=2.085 $X2=6.09 $Y2=2.23
r146 5 47 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.085 $X2=5.03 $Y2=2.91
r147 5 45 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.085 $X2=5.03 $Y2=2.23
r148 4 37 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=2.085 $X2=3.97 $Y2=2.91
r149 4 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=2.085 $X2=3.97 $Y2=2.23
r150 3 23 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=2.085 $X2=2.91 $Y2=2.91
r151 3 21 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=2.085 $X2=2.91 $Y2=2.23
r152 2 41 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.61
+ $Y=0.235 $X2=4.75 $Y2=0.51
r153 1 27 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.03
+ $Y=0.235 $X2=3.17 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_8%VGND 1 2 3 4 13 15 19 23 25 27 32 40 50
+ 51 68 71
r80 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r81 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r82 63 65 1.74286 $w=8.73e-07 $l=1.25e-07 $layer=LI1_cond $X=2.112 $Y=0.385
+ $X2=2.112 $Y2=0.51
r83 59 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r84 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r85 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r86 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r87 48 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r88 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=0 $X2=6.96 $Y2=0
r89 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r90 45 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.705 $Y=0 $X2=5.54
+ $Y2=0
r91 45 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.705 $Y=0 $X2=6
+ $Y2=0
r92 44 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r93 44 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r94 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r95 41 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.125 $Y=0 $X2=3.96
+ $Y2=0
r96 41 43 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=4.125 $Y=0 $X2=5.04
+ $Y2=0
r97 40 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=0 $X2=5.54
+ $Y2=0
r98 40 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.375 $Y=0 $X2=5.04
+ $Y2=0
r99 36 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r100 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r101 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r102 33 35 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.64
+ $Y2=0
r103 32 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.96
+ $Y2=0
r104 32 38 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.6
+ $Y2=0
r105 31 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r106 31 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r107 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r108 28 54 4.43563 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r109 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r110 27 63 5.368 $w=8.73e-07 $l=3.85e-07 $layer=LI1_cond $X=2.112 $Y=0 $X2=2.112
+ $Y2=0.385
r111 27 33 10.8128 $w=1.7e-07 $l=4.38e-07 $layer=LI1_cond $X=2.112 $Y=0 $X2=2.55
+ $Y2=0
r112 27 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r113 27 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r114 27 30 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.675 $Y=0
+ $X2=0.72 $Y2=0
r115 25 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r116 25 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r117 25 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r118 21 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.54 $Y=0.085
+ $X2=5.54 $Y2=0
r119 21 23 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=5.54 $Y=0.085
+ $X2=5.54 $Y2=0.51
r120 17 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0
r121 17 19 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0.44
r122 13 54 3.08204 $w=3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.212 $Y2=0
r123 13 15 11.5244 $w=2.98e-07 $l=3e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.385
r124 4 23 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.235 $X2=5.54 $Y2=0.51
r125 3 19 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.82
+ $Y=0.235 $X2=3.96 $Y2=0.44
r126 2 65 182 $w=1.7e-07 $l=8.05854e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.235 $X2=2.38 $Y2=0.51
r127 2 63 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=1.7
+ $Y=0.235 $X2=1.84 $Y2=0.385
r128 1 15 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.385
.ends

