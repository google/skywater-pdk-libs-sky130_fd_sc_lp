* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor2_2 A B VGND VNB VPB VPWR X
M1000 a_149_367# B a_149_65# VPB phighvt w=1.26e+06u l=150000u
+  ad=8.19e+11p pd=6.34e+06u as=3.528e+11p ps=3.08e+06u
M1001 a_149_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.8758e+12p ps=1.335e+07u
M1002 X a_149_65# a_532_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.3734e+12p ps=1.226e+07u
M1003 VGND A a_149_65# VNB nshort w=840000u l=150000u
+  ad=1.8502e+12p pd=1.342e+07u as=6.636e+11p ps=4.94e+06u
M1004 a_149_65# A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B a_532_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_532_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_149_65# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.914e+11p ps=4.53e+06u
M1008 a_814_65# A VGND VNB nshort w=840000u l=150000u
+  ad=7.77e+11p pd=5.21e+06u as=0p ps=0u
M1009 VGND B a_149_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A a_814_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_149_65# B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_814_65# B X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_532_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_149_65# B a_149_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A a_149_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_532_367# a_149_65# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_532_367# B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X B a_814_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_149_65# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
