* NGSPICE file created from sky130_fd_sc_lp__mux2i_lp2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__mux2i_lp2 A0 A1 S VGND VNB VPB VPWR Y
M1000 a_609_47# S VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=4.431e+11p ps=3.79e+06u
M1001 VPWR a_490_21# a_410_419# VPB phighvt w=1e+06u l=250000u
+  ad=6.15e+11p pd=5.23e+06u as=4.3e+11p ps=2.86e+06u
M1002 VGND a_490_21# a_422_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.428e+11p ps=1.52e+06u
M1003 a_490_21# S VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1004 Y A1 a_256_47# VNB nshort w=420000u l=150000u
+  ad=1.218e+11p pd=1.42e+06u as=1.008e+11p ps=1.32e+06u
M1005 a_256_47# S VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_148_419# S VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 Y A0 a_148_419# VPB phighvt w=1e+06u l=250000u
+  ad=5.7e+11p pd=3.14e+06u as=0p ps=0u
M1008 a_410_419# A1 Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_490_21# S a_609_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1010 a_422_47# A0 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

