* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 VGND CLK a_110_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_440_413# a_110_70# a_526_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_668_137# a_110_70# a_957_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 VPWR D a_440_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_626_163# a_668_137# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_957_379# a_1158_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 VPWR CLK a_110_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_217_413# a_110_70# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_1116_119# a_1158_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_526_413# a_217_413# a_626_163# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_217_413# a_110_70# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_526_413# a_110_70# a_666_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_957_379# a_110_70# a_1116_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_666_413# a_668_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 VGND a_1158_93# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR a_957_379# a_1158_93# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 VGND a_526_413# a_668_137# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 a_440_413# a_217_413# a_526_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_957_379# a_217_413# a_1116_379# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_1116_379# a_1158_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VPWR a_1158_93# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_668_137# a_217_413# a_957_379# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR a_526_413# a_668_137# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 VGND D a_440_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
