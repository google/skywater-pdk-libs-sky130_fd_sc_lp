* File: sky130_fd_sc_lp__o41a_m.spice
* Created: Fri Aug 28 11:19:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41a_m.pex.spice"
.subckt sky130_fd_sc_lp__o41a_m  VNB VPB B1 A4 A3 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_80_21#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_300_51#_M1009_d N_B1_M1009_g N_A_80_21#_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A4_M1001_g N_A_300_51#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_300_51#_M1008_d N_A3_M1008_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_300_51#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_300_51#_M1005_d N_A1_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_80_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06195 AS=0.1113 PD=0.715 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1007 N_A_80_21#_M1007_d N_B1_M1007_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06405 AS=0.06195 PD=0.725 PS=0.715 NRD=0 NRS=7.0329 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1003 A_329_535# N_A4_M1003_g N_A_80_21#_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.08925 AS=0.06405 PD=0.845 PS=0.725 NRD=73.875 NRS=11.7215 M=1 R=2.8
+ SA=75001.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1004 A_444_535# N_A3_M1004_g A_329_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.08925 PD=0.63 PS=0.845 NRD=23.443 NRS=73.875 M=1 R=2.8 SA=75001.7
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1010 A_516_535# N_A2_M1010_g A_444_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75002 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A1_M1011_g A_516_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_91 VPB 0 1.38473e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o41a_m.pxi.spice"
*
.ends
*
*
