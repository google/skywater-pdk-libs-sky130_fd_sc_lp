# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__edfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__edfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.180000 2.835000 1.510000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.285000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.920000 1.310000 2.735000 ;
        RECT 1.085000 2.735000 1.415000 3.065000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.571200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.045000 0.265000 14.300000 2.150000 ;
        RECT 14.050000 2.150000 14.300000 3.065000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.583800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.605000 1.835000 13.360000 2.165000 ;
        RECT 12.880000 0.895000 13.360000 1.145000 ;
        RECT 13.190000 1.145000 13.360000 1.835000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.840000 1.100000 7.170000 1.430000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.145000  0.085000  0.395000 1.335000 ;
      RECT  0.145000  2.385000  0.395000 3.245000 ;
      RECT  0.575000  0.875000  0.905000 1.235000 ;
      RECT  0.575000  1.235000  2.200000 1.565000 ;
      RECT  0.575000  1.565000  0.905000 3.065000 ;
      RECT  1.135000  0.265000  1.385000 0.885000 ;
      RECT  1.135000  0.885000  2.805000 1.000000 ;
      RECT  1.135000  1.000000  2.165000 1.055000 ;
      RECT  1.490000  1.745000  2.440000 1.915000 ;
      RECT  1.490000  1.915000  1.740000 2.555000 ;
      RECT  1.565000  0.085000  1.815000 0.705000 ;
      RECT  1.920000  2.095000  2.090000 3.245000 ;
      RECT  1.995000  0.265000  3.825000 0.435000 ;
      RECT  1.995000  0.435000  2.325000 0.650000 ;
      RECT  1.995000  0.830000  2.805000 0.885000 ;
      RECT  2.270000  1.915000  2.440000 2.735000 ;
      RECT  2.270000  2.735000  3.310000 2.905000 ;
      RECT  2.555000  0.615000  2.805000 0.830000 ;
      RECT  2.630000  1.745000  3.310000 1.915000 ;
      RECT  2.630000  1.915000  2.880000 2.555000 ;
      RECT  2.985000  0.615000  3.315000 1.000000 ;
      RECT  3.060000  2.095000  3.310000 2.735000 ;
      RECT  3.140000  1.000000  3.315000 1.100000 ;
      RECT  3.140000  1.100000  4.385000 1.270000 ;
      RECT  3.140000  1.270000  3.310000 1.745000 ;
      RECT  3.490000  1.450000  3.820000 1.780000 ;
      RECT  3.490000  1.780000  3.685000 2.150000 ;
      RECT  3.495000  0.435000  3.825000 0.920000 ;
      RECT  3.865000  1.960000  4.035000 2.895000 ;
      RECT  3.865000  2.895000  5.775000 3.065000 ;
      RECT  4.055000  0.435000  4.385000 1.100000 ;
      RECT  4.215000  1.270000  4.385000 2.545000 ;
      RECT  4.215000  2.545000  5.245000 2.715000 ;
      RECT  4.565000  0.435000  4.895000 1.075000 ;
      RECT  4.565000  1.075000  6.300000 1.245000 ;
      RECT  4.565000  1.245000  4.735000 2.365000 ;
      RECT  4.915000  1.450000  5.245000 1.780000 ;
      RECT  4.915000  1.960000  5.245000 2.545000 ;
      RECT  5.445000  2.265000  5.775000 2.895000 ;
      RECT  5.460000  0.085000  5.790000 0.895000 ;
      RECT  5.520000  1.555000  6.660000 1.885000 ;
      RECT  5.970000  0.985000  6.300000 1.075000 ;
      RECT  5.970000  1.245000  6.300000 1.315000 ;
      RECT  5.980000  2.065000  6.230000 3.245000 ;
      RECT  6.085000  0.265000  6.660000 0.805000 ;
      RECT  6.410000  1.885000  6.660000 2.820000 ;
      RECT  6.410000  2.820000  7.540000 2.990000 ;
      RECT  6.490000  0.805000  6.660000 1.555000 ;
      RECT  6.940000  1.610000  7.520000 1.780000 ;
      RECT  6.940000  1.780000  7.190000 2.640000 ;
      RECT  6.965000  0.540000  7.295000 0.750000 ;
      RECT  6.965000  0.750000  7.520000 0.920000 ;
      RECT  7.350000  0.920000  7.520000 1.100000 ;
      RECT  7.350000  1.100000  8.105000 1.270000 ;
      RECT  7.350000  1.270000  7.520000 1.610000 ;
      RECT  7.370000  1.960000  8.240000 2.130000 ;
      RECT  7.370000  2.130000  7.540000 2.820000 ;
      RECT  7.700000  0.085000  8.030000 0.920000 ;
      RECT  7.720000  2.310000  7.890000 3.245000 ;
      RECT  7.775000  1.270000  8.105000 1.770000 ;
      RECT  8.070000  2.130000  8.240000 2.515000 ;
      RECT  8.070000  2.515000  9.120000 2.685000 ;
      RECT  8.210000  0.460000  8.540000 0.920000 ;
      RECT  8.285000  0.920000  8.540000 1.385000 ;
      RECT  8.285000  1.385000  9.950000 1.555000 ;
      RECT  8.285000  1.555000  8.670000 1.780000 ;
      RECT  8.420000  1.780000  8.670000 2.335000 ;
      RECT  8.870000  2.865000 10.690000 3.065000 ;
      RECT  8.925000  0.685000  9.255000 0.895000 ;
      RECT  8.925000  0.895000 11.620000 1.065000 ;
      RECT  8.925000  1.065000  9.255000 1.145000 ;
      RECT  8.950000  1.735000 10.520000 1.905000 ;
      RECT  8.950000  1.905000  9.120000 2.515000 ;
      RECT  9.300000  2.085000  9.630000 2.435000 ;
      RECT  9.300000  2.435000 11.390000 2.605000 ;
      RECT  9.300000  2.605000  9.630000 2.685000 ;
      RECT  9.470000  0.265000  9.800000 0.545000 ;
      RECT  9.470000  0.545000 13.865000 0.595000 ;
      RECT  9.470000  0.595000 11.110000 0.715000 ;
      RECT  9.620000  1.245000  9.950000 1.385000 ;
      RECT  9.830000  2.085000 11.820000 2.255000 ;
      RECT 10.190000  1.345000 10.520000 1.735000 ;
      RECT 10.360000  2.785000 10.690000 2.865000 ;
      RECT 10.430000  0.085000 10.760000 0.365000 ;
      RECT 10.870000  2.785000 11.040000 3.245000 ;
      RECT 10.940000  0.265000 11.970000 0.545000 ;
      RECT 11.220000  2.605000 11.390000 2.705000 ;
      RECT 11.220000  2.705000 12.380000 2.875000 ;
      RECT 11.290000  0.775000 11.620000 0.895000 ;
      RECT 11.290000  1.065000 11.620000 1.145000 ;
      RECT 11.565000  1.595000 13.010000 1.655000 ;
      RECT 11.565000  1.655000 12.355000 1.905000 ;
      RECT 11.570000  2.255000 11.820000 2.525000 ;
      RECT 11.800000  0.595000 13.865000 0.715000 ;
      RECT 11.860000  0.895000 12.190000 1.325000 ;
      RECT 11.860000  1.325000 13.010000 1.595000 ;
      RECT 12.020000  1.905000 12.355000 2.165000 ;
      RECT 12.210000  2.345000 13.865000 2.515000 ;
      RECT 12.210000  2.515000 12.380000 2.705000 ;
      RECT 12.370000  0.085000 12.700000 0.365000 ;
      RECT 12.560000  2.695000 12.890000 3.245000 ;
      RECT 13.420000  0.085000 13.750000 0.365000 ;
      RECT 13.540000  0.715000 13.865000 2.345000 ;
      RECT 13.540000  2.695000 13.870000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  1.950000  3.685000 2.120000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.580000  5.125000 1.750000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.580000  8.485000 1.750000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  1.950000 12.325000 2.120000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
    LAYER met1 ;
      RECT  3.455000 1.920000  3.745000 1.965000 ;
      RECT  3.455000 1.965000 12.385000 2.105000 ;
      RECT  3.455000 2.105000  3.745000 2.150000 ;
      RECT  4.895000 1.550000  5.185000 1.595000 ;
      RECT  4.895000 1.595000  8.545000 1.735000 ;
      RECT  4.895000 1.735000  5.185000 1.780000 ;
      RECT  8.255000 1.550000  8.545000 1.595000 ;
      RECT  8.255000 1.735000  8.545000 1.780000 ;
      RECT 12.095000 1.920000 12.385000 1.965000 ;
      RECT 12.095000 2.105000 12.385000 2.150000 ;
  END
END sky130_fd_sc_lp__edfxbp_1
END LIBRARY
