* File: sky130_fd_sc_lp__nor4b_1.pxi.spice
* Created: Wed Sep  2 10:10:55 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4B_1%D_N N_D_N_M1005_g N_D_N_M1009_g N_D_N_c_63_n
+ N_D_N_c_64_n D_N N_D_N_c_65_n PM_SKY130_FD_SC_LP__NOR4B_1%D_N
x_PM_SKY130_FD_SC_LP__NOR4B_1%A N_A_M1006_g N_A_M1001_g A A N_A_c_93_n
+ N_A_c_94_n PM_SKY130_FD_SC_LP__NOR4B_1%A
x_PM_SKY130_FD_SC_LP__NOR4B_1%B N_B_M1003_g N_B_M1002_g B N_B_c_130_n
+ N_B_c_131_n N_B_c_132_n PM_SKY130_FD_SC_LP__NOR4B_1%B
x_PM_SKY130_FD_SC_LP__NOR4B_1%C N_C_M1007_g N_C_M1008_g C N_C_c_168_n
+ N_C_c_169_n N_C_c_172_n PM_SKY130_FD_SC_LP__NOR4B_1%C
x_PM_SKY130_FD_SC_LP__NOR4B_1%A_80_131# N_A_80_131#_M1005_s N_A_80_131#_M1009_s
+ N_A_80_131#_M1004_g N_A_80_131#_M1000_g N_A_80_131#_c_208_n
+ N_A_80_131#_c_214_n N_A_80_131#_c_209_n N_A_80_131#_c_234_n
+ N_A_80_131#_c_216_n N_A_80_131#_c_210_n N_A_80_131#_c_230_n
+ N_A_80_131#_c_211_n N_A_80_131#_c_212_n PM_SKY130_FD_SC_LP__NOR4B_1%A_80_131#
x_PM_SKY130_FD_SC_LP__NOR4B_1%VPWR N_VPWR_M1009_d N_VPWR_c_290_n VPWR
+ N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_289_n N_VPWR_c_294_n
+ PM_SKY130_FD_SC_LP__NOR4B_1%VPWR
x_PM_SKY130_FD_SC_LP__NOR4B_1%Y N_Y_M1006_d N_Y_M1008_d N_Y_M1000_d N_Y_c_331_n
+ N_Y_c_324_n N_Y_c_325_n N_Y_c_341_n N_Y_c_326_n N_Y_c_327_n Y Y Y N_Y_c_328_n
+ Y PM_SKY130_FD_SC_LP__NOR4B_1%Y
x_PM_SKY130_FD_SC_LP__NOR4B_1%VGND N_VGND_M1005_d N_VGND_M1002_d N_VGND_M1004_d
+ N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n
+ N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n VGND N_VGND_c_386_n
+ N_VGND_c_387_n PM_SKY130_FD_SC_LP__NOR4B_1%VGND
cc_1 VNB N_D_N_M1005_g 0.0321907f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=0.865
cc_2 VNB N_D_N_c_63_n 0.0376205f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.51
cc_3 VNB N_D_N_c_64_n 0.00907398f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.51
cc_4 VNB N_D_N_c_65_n 0.0149796f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_5 VNB N_A_M1001_g 0.00687248f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.045
cc_6 VNB A 0.00241781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_c_93_n 0.0326458f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_8 VNB N_A_c_94_n 0.0186054f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_9 VNB N_B_M1003_g 0.00341416f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=0.865
cc_10 VNB N_B_c_130_n 0.0374802f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB N_B_c_131_n 4.33617e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_c_132_n 0.0169076f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_13 VNB N_C_M1008_g 0.0254197f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.045
cc_14 VNB N_C_c_168_n 0.0244806f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_C_c_169_n 0.00333947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_80_131#_M1004_g 0.0281716f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.51
cc_17 VNB N_A_80_131#_c_208_n 0.0156811f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.592
cc_18 VNB N_A_80_131#_c_209_n 0.00274179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_80_131#_c_210_n 0.0142587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_80_131#_c_211_n 0.00295904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_80_131#_c_212_n 0.0255954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_289_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_324_n 0.00735546f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_24 VNB N_Y_c_325_n 0.00587681f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_25 VNB N_Y_c_326_n 0.0214066f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.592
cc_26 VNB N_Y_c_327_n 0.0051755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_328_n 0.0245542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_378_n 0.0149551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_379_n 0.00430889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_380_n 0.0156289f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.592
cc_31 VNB N_VGND_c_381_n 0.0253393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_382_n 0.0262736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_383_n 0.0073833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_384_n 0.0161841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_385_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_386_n 0.0151002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_387_n 0.212499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_D_N_M1009_g 0.0300424f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.045
cc_39 VPB N_D_N_c_63_n 0.0132284f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.51
cc_40 VPB N_D_N_c_64_n 6.62969e-19 $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.51
cc_41 VPB N_D_N_c_65_n 0.0170379f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=1.51
cc_42 VPB N_A_M1001_g 0.0212018f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.045
cc_43 VPB A 0.00185829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_B_M1003_g 0.0200051f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=0.865
cc_45 VPB N_B_c_131_n 0.00256202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_C_c_168_n 0.00972833f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_47 VPB N_C_c_169_n 0.00273901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_C_c_172_n 0.0176926f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=1.51
cc_49 VPB N_A_80_131#_M1000_g 0.0225724f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=1.51
cc_50 VPB N_A_80_131#_c_214_n 0.010409f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_80_131#_c_209_n 0.00128026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_80_131#_c_216_n 0.0014691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_80_131#_c_211_n 4.51888e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_80_131#_c_212_n 0.00761581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_290_n 0.0312828f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.045
cc_56 VPB N_VPWR_c_291_n 0.0307831f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.51
cc_57 VPB N_VPWR_c_292_n 0.065039f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.592
cc_58 VPB N_VPWR_c_289_n 0.0784897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_294_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB Y 0.0564761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_Y_c_328_n 0.00949208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 N_D_N_c_64_n N_A_M1001_g 0.0232239f $X=0.74 $Y=1.51 $X2=0 $Y2=0
cc_63 N_D_N_M1005_g A 5.23459e-19 $X=0.74 $Y=0.865 $X2=0 $Y2=0
cc_64 N_D_N_c_64_n A 7.39329e-19 $X=0.74 $Y=1.51 $X2=0 $Y2=0
cc_65 N_D_N_M1005_g N_A_c_93_n 0.0203917f $X=0.74 $Y=0.865 $X2=0 $Y2=0
cc_66 N_D_N_M1005_g N_A_c_94_n 0.0129476f $X=0.74 $Y=0.865 $X2=0 $Y2=0
cc_67 N_D_N_M1005_g N_A_80_131#_c_208_n 6.81439e-19 $X=0.74 $Y=0.865 $X2=0 $Y2=0
cc_68 N_D_N_M1009_g N_A_80_131#_c_214_n 0.00868156f $X=0.74 $Y=2.045 $X2=0 $Y2=0
cc_69 N_D_N_c_63_n N_A_80_131#_c_214_n 0.00270669f $X=0.665 $Y=1.51 $X2=0 $Y2=0
cc_70 N_D_N_c_65_n N_A_80_131#_c_214_n 0.0186708f $X=0.43 $Y=1.51 $X2=0 $Y2=0
cc_71 N_D_N_M1005_g N_A_80_131#_c_209_n 0.00436146f $X=0.74 $Y=0.865 $X2=0 $Y2=0
cc_72 N_D_N_M1009_g N_A_80_131#_c_209_n 0.010497f $X=0.74 $Y=2.045 $X2=0 $Y2=0
cc_73 N_D_N_c_64_n N_A_80_131#_c_209_n 0.0105715f $X=0.74 $Y=1.51 $X2=0 $Y2=0
cc_74 N_D_N_c_65_n N_A_80_131#_c_209_n 0.025095f $X=0.43 $Y=1.51 $X2=0 $Y2=0
cc_75 N_D_N_M1005_g N_A_80_131#_c_210_n 0.0156449f $X=0.74 $Y=0.865 $X2=0 $Y2=0
cc_76 N_D_N_c_63_n N_A_80_131#_c_210_n 0.00789557f $X=0.665 $Y=1.51 $X2=0 $Y2=0
cc_77 N_D_N_c_65_n N_A_80_131#_c_210_n 0.0176803f $X=0.43 $Y=1.51 $X2=0 $Y2=0
cc_78 N_D_N_M1009_g N_A_80_131#_c_230_n 0.00617411f $X=0.74 $Y=2.045 $X2=0 $Y2=0
cc_79 N_D_N_M1009_g N_VPWR_c_290_n 0.0020569f $X=0.74 $Y=2.045 $X2=0 $Y2=0
cc_80 N_D_N_M1005_g N_VGND_c_378_n 0.0129869f $X=0.74 $Y=0.865 $X2=0 $Y2=0
cc_81 N_D_N_M1005_g N_VGND_c_382_n 0.00332367f $X=0.74 $Y=0.865 $X2=0 $Y2=0
cc_82 N_D_N_M1005_g N_VGND_c_387_n 0.00387424f $X=0.74 $Y=0.865 $X2=0 $Y2=0
cc_83 N_A_M1001_g N_B_M1003_g 0.0636834f $X=1.28 $Y=2.465 $X2=0 $Y2=0
cc_84 A N_B_c_130_n 0.00228807f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A_c_93_n N_B_c_130_n 0.0636834f $X=1.19 $Y=1.35 $X2=0 $Y2=0
cc_86 A N_B_c_131_n 0.022331f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A_c_93_n N_B_c_131_n 0.00157042f $X=1.19 $Y=1.35 $X2=0 $Y2=0
cc_88 N_A_c_94_n N_B_c_132_n 0.0131577f $X=1.19 $Y=1.185 $X2=0 $Y2=0
cc_89 N_A_M1001_g N_A_80_131#_c_209_n 0.00326293f $X=1.28 $Y=2.465 $X2=0 $Y2=0
cc_90 A N_A_80_131#_c_209_n 0.0402227f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A_c_93_n N_A_80_131#_c_209_n 0.00161233f $X=1.19 $Y=1.35 $X2=0 $Y2=0
cc_92 N_A_M1001_g N_A_80_131#_c_234_n 0.0165233f $X=1.28 $Y=2.465 $X2=0 $Y2=0
cc_93 A N_A_80_131#_c_234_n 0.012212f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A_c_93_n N_A_80_131#_c_234_n 0.00255229f $X=1.19 $Y=1.35 $X2=0 $Y2=0
cc_95 A N_A_80_131#_c_210_n 0.0130324f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A_c_93_n N_A_80_131#_c_210_n 4.85341e-19 $X=1.19 $Y=1.35 $X2=0 $Y2=0
cc_97 N_A_c_94_n N_A_80_131#_c_210_n 3.86628e-19 $X=1.19 $Y=1.185 $X2=0 $Y2=0
cc_98 N_A_M1001_g N_A_80_131#_c_230_n 9.75296e-19 $X=1.28 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_M1001_g N_VPWR_c_290_n 0.0225272f $X=1.28 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_M1001_g N_VPWR_c_292_n 0.00486043f $X=1.28 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A_M1001_g N_VPWR_c_289_n 0.00818711f $X=1.28 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_c_94_n N_Y_c_331_n 0.004326f $X=1.19 $Y=1.185 $X2=0 $Y2=0
cc_103 A N_Y_c_325_n 0.00566835f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_A_c_94_n N_Y_c_325_n 0.00309955f $X=1.19 $Y=1.185 $X2=0 $Y2=0
cc_105 A N_VGND_c_378_n 0.00904577f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_106 N_A_c_93_n N_VGND_c_378_n 0.00370647f $X=1.19 $Y=1.35 $X2=0 $Y2=0
cc_107 N_A_c_94_n N_VGND_c_378_n 0.0192313f $X=1.19 $Y=1.185 $X2=0 $Y2=0
cc_108 N_A_c_94_n N_VGND_c_384_n 0.00447018f $X=1.19 $Y=1.185 $X2=0 $Y2=0
cc_109 N_A_c_94_n N_VGND_c_387_n 0.00775973f $X=1.19 $Y=1.185 $X2=0 $Y2=0
cc_110 N_B_c_130_n N_C_M1008_g 0.00758075f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_111 N_B_c_132_n N_C_M1008_g 0.011976f $X=1.73 $Y=1.185 $X2=0 $Y2=0
cc_112 N_B_M1003_g N_C_c_168_n 0.0578639f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B_c_130_n N_C_c_168_n 0.0150032f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_114 N_B_c_131_n N_C_c_168_n 0.00102077f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_115 N_B_M1003_g N_C_c_169_n 5.30471e-19 $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B_c_130_n N_C_c_169_n 0.00133446f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_117 N_B_c_131_n N_C_c_169_n 0.036526f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_118 N_B_M1003_g N_A_80_131#_c_234_n 0.015028f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B_c_130_n N_A_80_131#_c_234_n 6.75677e-19 $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_120 N_B_c_131_n N_A_80_131#_c_234_n 0.0233346f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_121 N_B_M1003_g N_VPWR_c_290_n 0.00506879f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_122 N_B_M1003_g N_VPWR_c_292_n 0.00585385f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B_M1003_g N_VPWR_c_289_n 0.011101f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B_c_132_n N_Y_c_331_n 0.00946463f $X=1.73 $Y=1.185 $X2=0 $Y2=0
cc_125 N_B_c_130_n N_Y_c_324_n 0.00182968f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_126 N_B_c_131_n N_Y_c_324_n 0.0156305f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_127 N_B_c_132_n N_Y_c_324_n 0.0131165f $X=1.73 $Y=1.185 $X2=0 $Y2=0
cc_128 N_B_c_130_n N_Y_c_325_n 0.00377847f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_129 N_B_c_131_n N_Y_c_325_n 0.0103022f $X=1.73 $Y=1.42 $X2=0 $Y2=0
cc_130 N_B_c_132_n N_Y_c_325_n 0.0010422f $X=1.73 $Y=1.185 $X2=0 $Y2=0
cc_131 N_B_c_132_n N_Y_c_341_n 3.50616e-19 $X=1.73 $Y=1.185 $X2=0 $Y2=0
cc_132 N_B_c_132_n N_VGND_c_378_n 7.43856e-19 $X=1.73 $Y=1.185 $X2=0 $Y2=0
cc_133 N_B_c_132_n N_VGND_c_379_n 0.0017823f $X=1.73 $Y=1.185 $X2=0 $Y2=0
cc_134 N_B_c_132_n N_VGND_c_384_n 0.00579312f $X=1.73 $Y=1.185 $X2=0 $Y2=0
cc_135 N_B_c_132_n N_VGND_c_387_n 0.0108127f $X=1.73 $Y=1.185 $X2=0 $Y2=0
cc_136 N_C_M1008_g N_A_80_131#_M1004_g 0.024485f $X=2.29 $Y=0.655 $X2=0 $Y2=0
cc_137 N_C_c_169_n N_A_80_131#_M1000_g 2.55025e-19 $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_138 N_C_c_172_n N_A_80_131#_M1000_g 0.0477046f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_139 N_C_c_168_n N_A_80_131#_c_234_n 0.00334683f $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_140 N_C_c_169_n N_A_80_131#_c_234_n 0.0186442f $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_141 N_C_c_172_n N_A_80_131#_c_234_n 0.0161077f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_142 N_C_c_168_n N_A_80_131#_c_216_n 3.10063e-19 $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_143 N_C_c_169_n N_A_80_131#_c_216_n 0.00960555f $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_144 N_C_c_172_n N_A_80_131#_c_216_n 0.00346437f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_145 N_C_c_168_n N_A_80_131#_c_211_n 0.00220021f $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_146 N_C_c_169_n N_A_80_131#_c_211_n 0.0260787f $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_147 N_C_c_168_n N_A_80_131#_c_212_n 0.0234944f $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_148 N_C_c_169_n N_A_80_131#_c_212_n 2.86228e-19 $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_149 N_C_c_172_n N_VPWR_c_292_n 0.00585385f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_150 N_C_c_172_n N_VPWR_c_289_n 0.011557f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_151 N_C_M1008_g N_Y_c_331_n 3.77632e-19 $X=2.29 $Y=0.655 $X2=0 $Y2=0
cc_152 N_C_M1008_g N_Y_c_324_n 0.0128049f $X=2.29 $Y=0.655 $X2=0 $Y2=0
cc_153 N_C_c_168_n N_Y_c_324_n 7.55836e-19 $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_154 N_C_c_169_n N_Y_c_324_n 0.0209945f $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_155 N_C_M1008_g N_Y_c_341_n 0.00949957f $X=2.29 $Y=0.655 $X2=0 $Y2=0
cc_156 N_C_M1008_g N_Y_c_327_n 0.00187559f $X=2.29 $Y=0.655 $X2=0 $Y2=0
cc_157 N_C_c_168_n N_Y_c_327_n 0.00312334f $X=2.27 $Y=1.51 $X2=0 $Y2=0
cc_158 N_C_M1008_g N_VGND_c_379_n 0.0017186f $X=2.29 $Y=0.655 $X2=0 $Y2=0
cc_159 N_C_M1008_g N_VGND_c_381_n 6.85043e-19 $X=2.29 $Y=0.655 $X2=0 $Y2=0
cc_160 N_C_M1008_g N_VGND_c_386_n 0.00571722f $X=2.29 $Y=0.655 $X2=0 $Y2=0
cc_161 N_C_M1008_g N_VGND_c_387_n 0.0105634f $X=2.29 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A_80_131#_c_209_n N_VPWR_M1009_d 0.00117769f $X=0.85 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_80_131#_c_234_n N_VPWR_M1009_d 0.00747572f $X=2.525 $Y=2.055
+ $X2=-0.19 $Y2=-0.245
cc_164 N_A_80_131#_c_230_n N_VPWR_M1009_d 0.0022391f $X=0.85 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A_80_131#_c_234_n N_VPWR_c_290_n 0.0190878f $X=2.525 $Y=2.055 $X2=0
+ $Y2=0
cc_166 N_A_80_131#_c_230_n N_VPWR_c_290_n 0.00308053f $X=0.85 $Y=2.035 $X2=0
+ $Y2=0
cc_167 N_A_80_131#_M1000_g N_VPWR_c_292_n 0.00585385f $X=2.72 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_80_131#_M1000_g N_VPWR_c_289_n 0.0122168f $X=2.72 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_80_131#_c_234_n A_271_367# 0.00732587f $X=2.525 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A_80_131#_c_234_n A_343_367# 0.0177931f $X=2.525 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_80_131#_c_234_n A_451_367# 0.0157906f $X=2.525 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_172 N_A_80_131#_c_216_n A_451_367# 0.00167884f $X=2.61 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_80_131#_c_210_n N_Y_c_325_n 3.78847e-19 $X=0.85 $Y=1.17 $X2=0 $Y2=0
cc_174 N_A_80_131#_M1004_g N_Y_c_326_n 0.0155226f $X=2.72 $Y=0.655 $X2=0 $Y2=0
cc_175 N_A_80_131#_c_211_n N_Y_c_326_n 0.02091f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A_80_131#_c_212_n N_Y_c_326_n 0.00522192f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A_80_131#_c_211_n N_Y_c_327_n 0.00637106f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_178 N_A_80_131#_M1000_g Y 0.0253614f $X=2.72 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A_80_131#_c_234_n Y 0.0141922f $X=2.525 $Y=2.055 $X2=0 $Y2=0
cc_180 N_A_80_131#_c_216_n Y 0.00938007f $X=2.61 $Y=1.97 $X2=0 $Y2=0
cc_181 N_A_80_131#_c_211_n Y 0.00239484f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A_80_131#_c_212_n Y 0.00423088f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A_80_131#_M1004_g N_Y_c_328_n 0.00564501f $X=2.72 $Y=0.655 $X2=0 $Y2=0
cc_184 N_A_80_131#_M1000_g N_Y_c_328_n 0.00306041f $X=2.72 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_80_131#_c_216_n N_Y_c_328_n 0.00688405f $X=2.61 $Y=1.97 $X2=0 $Y2=0
cc_186 N_A_80_131#_c_211_n N_Y_c_328_n 0.0253922f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_187 N_A_80_131#_c_212_n N_Y_c_328_n 0.00820562f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_188 N_A_80_131#_c_210_n N_VGND_c_378_n 0.00915057f $X=0.85 $Y=1.17 $X2=0
+ $Y2=0
cc_189 N_A_80_131#_M1004_g N_VGND_c_381_n 0.0111637f $X=2.72 $Y=0.655 $X2=0
+ $Y2=0
cc_190 N_A_80_131#_c_208_n N_VGND_c_382_n 0.0041128f $X=0.525 $Y=0.865 $X2=0
+ $Y2=0
cc_191 N_A_80_131#_M1004_g N_VGND_c_386_n 0.00486043f $X=2.72 $Y=0.655 $X2=0
+ $Y2=0
cc_192 N_A_80_131#_M1004_g N_VGND_c_387_n 0.0082726f $X=2.72 $Y=0.655 $X2=0
+ $Y2=0
cc_193 N_A_80_131#_c_208_n N_VGND_c_387_n 0.00726513f $X=0.525 $Y=0.865 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_289_n A_271_367# 0.00899413f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_195 N_VPWR_c_289_n A_343_367# 0.0167135f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_196 N_VPWR_c_289_n A_451_367# 0.0167135f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_197 N_VPWR_c_289_n N_Y_M1000_d 0.00487993f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_198 N_VPWR_c_292_n Y 0.0289335f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_289_n Y 0.0158621f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_200 N_Y_c_324_n N_VGND_M1002_d 0.0029901f $X=2.355 $Y=1.08 $X2=0 $Y2=0
cc_201 N_Y_c_326_n N_VGND_M1004_d 0.00263371f $X=3.065 $Y=1.075 $X2=0 $Y2=0
cc_202 N_Y_c_331_n N_VGND_c_378_n 0.0425995f $X=1.54 $Y=0.42 $X2=0 $Y2=0
cc_203 N_Y_c_324_n N_VGND_c_379_n 0.0220482f $X=2.355 $Y=1.08 $X2=0 $Y2=0
cc_204 N_Y_c_326_n N_VGND_c_381_n 0.0223528f $X=3.065 $Y=1.075 $X2=0 $Y2=0
cc_205 N_Y_c_331_n N_VGND_c_384_n 0.0140046f $X=1.54 $Y=0.42 $X2=0 $Y2=0
cc_206 N_Y_c_341_n N_VGND_c_386_n 0.0146655f $X=2.505 $Y=0.42 $X2=0 $Y2=0
cc_207 N_Y_M1006_d N_VGND_c_387_n 0.00607622f $X=1.355 $Y=0.235 $X2=0 $Y2=0
cc_208 N_Y_M1008_d N_VGND_c_387_n 0.00380103f $X=2.365 $Y=0.235 $X2=0 $Y2=0
cc_209 N_Y_c_331_n N_VGND_c_387_n 0.00877263f $X=1.54 $Y=0.42 $X2=0 $Y2=0
cc_210 N_Y_c_341_n N_VGND_c_387_n 0.00933292f $X=2.505 $Y=0.42 $X2=0 $Y2=0
