* File: sky130_fd_sc_lp__dlclkp_2.pxi.spice
* Created: Wed Sep  2 09:45:47 2020
* 
x_PM_SKY130_FD_SC_LP__DLCLKP_2%A_78_269# N_A_78_269#_M1015_d N_A_78_269#_M1004_d
+ N_A_78_269#_M1009_g N_A_78_269#_M1005_g N_A_78_269#_c_150_n
+ N_A_78_269#_c_158_n N_A_78_269#_c_151_n N_A_78_269#_c_160_n
+ N_A_78_269#_c_166_p N_A_78_269#_c_152_n N_A_78_269#_c_168_p
+ N_A_78_269#_c_153_n N_A_78_269#_c_154_n N_A_78_269#_c_171_p
+ N_A_78_269#_c_155_n PM_SKY130_FD_SC_LP__DLCLKP_2%A_78_269#
x_PM_SKY130_FD_SC_LP__DLCLKP_2%GATE N_GATE_M1011_g N_GATE_M1020_g GATE
+ N_GATE_c_257_n PM_SKY130_FD_SC_LP__DLCLKP_2%GATE
x_PM_SKY130_FD_SC_LP__DLCLKP_2%A_284_367# N_A_284_367#_M1019_d
+ N_A_284_367#_M1001_d N_A_284_367#_M1004_g N_A_284_367#_M1021_g
+ N_A_284_367#_c_314_n N_A_284_367#_c_315_n N_A_284_367#_c_306_n
+ N_A_284_367#_c_307_n N_A_284_367#_c_317_n N_A_284_367#_c_308_n
+ N_A_284_367#_c_309_n N_A_284_367#_c_310_n N_A_284_367#_c_319_n
+ N_A_284_367#_c_311_n N_A_284_367#_c_320_n N_A_284_367#_c_321_n
+ N_A_284_367#_c_312_n PM_SKY130_FD_SC_LP__DLCLKP_2%A_284_367#
x_PM_SKY130_FD_SC_LP__DLCLKP_2%A_300_55# N_A_300_55#_M1007_s N_A_300_55#_M1008_s
+ N_A_300_55#_M1015_g N_A_300_55#_c_427_n N_A_300_55#_c_428_n
+ N_A_300_55#_M1012_g N_A_300_55#_M1019_g N_A_300_55#_M1001_g
+ N_A_300_55#_c_430_n N_A_300_55#_c_431_n N_A_300_55#_c_432_n
+ N_A_300_55#_c_433_n N_A_300_55#_c_434_n N_A_300_55#_c_435_n
+ N_A_300_55#_c_507_p N_A_300_55#_c_436_n N_A_300_55#_c_437_n
+ N_A_300_55#_c_438_n N_A_300_55#_c_439_n PM_SKY130_FD_SC_LP__DLCLKP_2%A_300_55#
x_PM_SKY130_FD_SC_LP__DLCLKP_2%A_33_47# N_A_33_47#_M1005_s N_A_33_47#_M1009_s
+ N_A_33_47#_M1014_g N_A_33_47#_M1013_g N_A_33_47#_c_555_n N_A_33_47#_c_556_n
+ N_A_33_47#_M1002_g N_A_33_47#_M1016_g N_A_33_47#_c_540_n N_A_33_47#_c_558_n
+ N_A_33_47#_c_541_n N_A_33_47#_c_575_n N_A_33_47#_c_577_n N_A_33_47#_c_542_n
+ N_A_33_47#_c_543_n N_A_33_47#_c_559_n N_A_33_47#_c_560_n N_A_33_47#_c_618_n
+ N_A_33_47#_c_585_n N_A_33_47#_c_544_n N_A_33_47#_c_561_n N_A_33_47#_c_562_n
+ N_A_33_47#_c_563_n N_A_33_47#_c_545_n N_A_33_47#_c_546_n N_A_33_47#_c_547_n
+ N_A_33_47#_c_548_n N_A_33_47#_c_549_n N_A_33_47#_c_565_n N_A_33_47#_c_550_n
+ N_A_33_47#_c_567_n N_A_33_47#_c_551_n N_A_33_47#_c_552_n N_A_33_47#_c_568_n
+ N_A_33_47#_c_553_n PM_SKY130_FD_SC_LP__DLCLKP_2%A_33_47#
x_PM_SKY130_FD_SC_LP__DLCLKP_2%CLK N_CLK_c_768_n N_CLK_M1007_g N_CLK_c_775_n
+ N_CLK_M1008_g N_CLK_M1006_g N_CLK_c_776_n N_CLK_M1000_g N_CLK_c_771_n CLK
+ N_CLK_c_772_n N_CLK_c_773_n PM_SKY130_FD_SC_LP__DLCLKP_2%CLK
x_PM_SKY130_FD_SC_LP__DLCLKP_2%A_1039_367# N_A_1039_367#_M1002_d
+ N_A_1039_367#_M1000_d N_A_1039_367#_M1003_g N_A_1039_367#_M1010_g
+ N_A_1039_367#_c_832_n N_A_1039_367#_M1017_g N_A_1039_367#_M1018_g
+ N_A_1039_367#_c_835_n N_A_1039_367#_c_842_n N_A_1039_367#_c_843_n
+ N_A_1039_367#_c_844_n N_A_1039_367#_c_836_n N_A_1039_367#_c_837_n
+ N_A_1039_367#_c_838_n N_A_1039_367#_c_839_n
+ PM_SKY130_FD_SC_LP__DLCLKP_2%A_1039_367#
x_PM_SKY130_FD_SC_LP__DLCLKP_2%VPWR N_VPWR_M1009_d N_VPWR_M1014_d N_VPWR_M1008_d
+ N_VPWR_M1016_d N_VPWR_M1018_d N_VPWR_c_907_n N_VPWR_c_908_n N_VPWR_c_909_n
+ N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_913_n VPWR
+ N_VPWR_c_914_n N_VPWR_c_915_n N_VPWR_c_916_n N_VPWR_c_917_n N_VPWR_c_918_n
+ N_VPWR_c_919_n N_VPWR_c_920_n N_VPWR_c_906_n PM_SKY130_FD_SC_LP__DLCLKP_2%VPWR
x_PM_SKY130_FD_SC_LP__DLCLKP_2%GCLK N_GCLK_M1003_s N_GCLK_M1010_s GCLK GCLK GCLK
+ GCLK GCLK GCLK GCLK N_GCLK_c_996_n PM_SKY130_FD_SC_LP__DLCLKP_2%GCLK
x_PM_SKY130_FD_SC_LP__DLCLKP_2%VGND N_VGND_M1005_d N_VGND_M1013_d N_VGND_M1007_d
+ N_VGND_M1003_d N_VGND_M1017_d N_VGND_c_1014_n N_VGND_c_1015_n N_VGND_c_1016_n
+ N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n N_VGND_c_1020_n VGND
+ N_VGND_c_1021_n N_VGND_c_1022_n N_VGND_c_1023_n N_VGND_c_1024_n
+ N_VGND_c_1025_n N_VGND_c_1026_n N_VGND_c_1027_n N_VGND_c_1028_n
+ PM_SKY130_FD_SC_LP__DLCLKP_2%VGND
cc_1 VNB N_A_78_269#_M1005_g 0.0326355f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_2 VNB N_A_78_269#_c_150_n 0.00882991f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.645
cc_3 VNB N_A_78_269#_c_151_n 0.00656732f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.645
cc_4 VNB N_A_78_269#_c_152_n 0.00526455f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.56
cc_5 VNB N_A_78_269#_c_153_n 0.00177148f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.51
cc_6 VNB N_A_78_269#_c_154_n 0.0288009f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.51
cc_7 VNB N_A_78_269#_c_155_n 0.00317836f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.69
cc_8 VNB N_GATE_M1011_g 0.0103506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_GATE_M1020_g 0.0256842f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.675
cc_10 VNB GATE 0.00634567f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.465
cc_11 VNB N_GATE_c_257_n 0.0331671f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_12 VNB N_A_284_367#_c_306_n 0.00875212f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.645
cc_13 VNB N_A_284_367#_c_307_n 0.0190734f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=0.845
cc_14 VNB N_A_284_367#_c_308_n 0.00510953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_284_367#_c_309_n 0.00313307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_284_367#_c_310_n 0.0287171f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.645
cc_17 VNB N_A_284_367#_c_311_n 0.00255704f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.69
cc_18 VNB N_A_284_367#_c_312_n 0.0158728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_300_55#_M1015_g 0.0410981f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.465
cc_20 VNB N_A_300_55#_c_427_n 0.0189375f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.345
cc_21 VNB N_A_300_55#_c_428_n 0.0064959f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_22 VNB N_A_300_55#_M1001_g 0.00254669f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=2.365
cc_23 VNB N_A_300_55#_c_430_n 0.00583111f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=2.45
cc_24 VNB N_A_300_55#_c_431_n 0.0233917f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=2.57
cc_25 VNB N_A_300_55#_c_432_n 0.0387593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_300_55#_c_433_n 0.017963f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.51
cc_27 VNB N_A_300_55#_c_434_n 0.00983025f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.51
cc_28 VNB N_A_300_55#_c_435_n 0.0244949f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.645
cc_29 VNB N_A_300_55#_c_436_n 0.0191703f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.69
cc_30 VNB N_A_300_55#_c_437_n 0.0176933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_300_55#_c_438_n 0.00134058f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.51
cc_32 VNB N_A_300_55#_c_439_n 0.011075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_33_47#_M1002_g 0.020487f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=2.28
cc_34 VNB N_A_33_47#_M1016_g 0.00270855f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=2.365
cc_35 VNB N_A_33_47#_c_540_n 0.0159574f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=2.57
cc_36 VNB N_A_33_47#_c_541_n 0.00465245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_33_47#_c_542_n 0.00932976f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.725
cc_38 VNB N_A_33_47#_c_543_n 0.002342f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.69
cc_39 VNB N_A_33_47#_c_544_n 0.00119954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_33_47#_c_545_n 4.39498e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_33_47#_c_546_n 0.00142546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_33_47#_c_547_n 0.0111269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_33_47#_c_548_n 0.0479434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_33_47#_c_549_n 0.0216011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_33_47#_c_550_n 0.0265343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_33_47#_c_551_n 0.00517695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_33_47#_c_552_n 0.0338703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_33_47#_c_553_n 0.0170289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_CLK_c_768_n 0.0121762f $X=-0.19 $Y=-0.245 $X2=1.65 $Y2=0.405
cc_50 VNB N_CLK_M1007_g 0.0326072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_CLK_M1006_g 0.0284363f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_52 VNB N_CLK_c_771_n 0.0372985f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.645
cc_53 VNB N_CLK_c_772_n 0.0185797f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=0.845
cc_54 VNB N_CLK_c_773_n 0.0023078f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=2.57
cc_55 VNB N_A_1039_367#_M1003_g 0.027658f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.465
cc_56 VNB N_A_1039_367#_c_832_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.645
cc_57 VNB N_A_1039_367#_M1017_g 0.0343508f $X=-0.19 $Y=-0.245 $X2=1.505
+ $Y2=1.645
cc_58 VNB N_A_1039_367#_M1018_g 0.0127435f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=0.845
cc_59 VNB N_A_1039_367#_c_835_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=2.45
cc_60 VNB N_A_1039_367#_c_836_n 0.0119835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1039_367#_c_837_n 0.00190724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1039_367#_c_838_n 0.00693069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1039_367#_c_839_n 0.0267273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VPWR_c_906_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_GCLK_c_996_n 0.00713842f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=2.365
cc_66 VNB N_VGND_c_1014_n 0.00487234f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=2.28
cc_67 VNB N_VGND_c_1015_n 0.00998567f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=2.365
cc_68 VNB N_VGND_c_1016_n 0.0182909f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=2.57
cc_69 VNB N_VGND_c_1017_n 0.0125005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1018_n 0.0496258f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.51
cc_71 VNB N_VGND_c_1019_n 0.0429461f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.645
cc_72 VNB N_VGND_c_1020_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1021_n 0.0159682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1022_n 0.0415728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1023_n 0.0335558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1024_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1025_n 0.00510306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1026_n 0.0197062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1027_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1028_n 0.419211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VPB N_A_78_269#_M1009_g 0.02571f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.465
cc_82 VPB N_A_78_269#_c_150_n 0.0117834f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.645
cc_83 VPB N_A_78_269#_c_158_n 0.0052162f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=2.28
cc_84 VPB N_A_78_269#_c_151_n 0.00440583f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=1.645
cc_85 VPB N_A_78_269#_c_160_n 0.00463408f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=2.365
cc_86 VPB N_A_78_269#_c_153_n 0.00520645f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.51
cc_87 VPB N_A_78_269#_c_154_n 0.0064426f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.51
cc_88 VPB N_GATE_M1011_g 0.0491489f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_284_367#_M1004_g 0.0206495f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.465
cc_90 VPB N_A_284_367#_c_314_n 0.00414998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_284_367#_c_315_n 0.03026f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=1.73
cc_92 VPB N_A_284_367#_c_306_n 0.00249812f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=1.645
cc_93 VPB N_A_284_367#_c_317_n 0.0169305f $X=-0.19 $Y=1.655 $X2=1.685 $Y2=2.45
cc_94 VPB N_A_284_367#_c_308_n 7.23502e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_284_367#_c_319_n 0.00423566f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=1.645
cc_96 VPB N_A_284_367#_c_320_n 0.012536f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.345
cc_97 VPB N_A_284_367#_c_321_n 0.00848808f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.675
cc_98 VPB N_A_300_55#_M1012_g 0.0441087f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.645
cc_99 VPB N_A_300_55#_M1001_g 0.036642f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=2.365
cc_100 VPB N_A_300_55#_c_430_n 0.0066709f $X=-0.19 $Y=1.655 $X2=1.685 $Y2=2.45
cc_101 VPB N_A_300_55#_c_434_n 0.00618043f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.51
cc_102 VPB N_A_300_55#_c_435_n 0.0195645f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.645
cc_103 VPB N_A_300_55#_c_439_n 0.00582619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_33_47#_M1014_g 0.0242294f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.465
cc_105 VPB N_A_33_47#_c_555_n 0.0589721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_33_47#_c_556_n 0.0120388f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.645
cc_107 VPB N_A_33_47#_M1016_g 0.0232235f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=2.365
cc_108 VPB N_A_33_47#_c_558_n 0.0292908f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.51
cc_109 VPB N_A_33_47#_c_559_n 0.0116915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_33_47#_c_560_n 0.00156976f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.675
cc_111 VPB N_A_33_47#_c_561_n 0.0125202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_33_47#_c_562_n 0.0568279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_33_47#_c_563_n 0.0218301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_33_47#_c_545_n 0.00132227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_33_47#_c_565_n 0.00666696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_33_47#_c_550_n 0.0115702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_33_47#_c_567_n 9.93719e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_33_47#_c_568_n 0.00422587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_CLK_c_768_n 0.0151888f $X=-0.19 $Y=1.655 $X2=1.65 $Y2=0.405
cc_120 VPB N_CLK_c_775_n 0.0223224f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=1.675
cc_121 VPB N_CLK_c_776_n 0.0198424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_CLK_c_771_n 0.0316106f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=1.645
cc_123 VPB N_CLK_c_772_n 0.0211415f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=0.845
cc_124 VPB N_CLK_c_773_n 0.00531213f $X=-0.19 $Y=1.655 $X2=1.71 $Y2=2.57
cc_125 VPB N_A_1039_367#_M1010_g 0.0206806f $X=-0.19 $Y=1.655 $X2=0.525
+ $Y2=0.655
cc_126 VPB N_A_1039_367#_M1018_g 0.0272186f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=0.845
cc_127 VPB N_A_1039_367#_c_842_n 0.0072437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_1039_367#_c_843_n 0.00293302f $X=-0.19 $Y=1.655 $X2=0.555
+ $Y2=1.51
cc_129 VPB N_A_1039_367#_c_844_n 0.00365976f $X=-0.19 $Y=1.655 $X2=0.555
+ $Y2=1.51
cc_130 VPB N_A_1039_367#_c_837_n 3.04024e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_1039_367#_c_839_n 0.00789152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_907_n 0.0081699f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=1.645
cc_133 VPB N_VPWR_c_908_n 0.0386802f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.56
cc_134 VPB N_VPWR_c_909_n 0.026016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_910_n 0.0119938f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_911_n 0.0640295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_912_n 0.0525124f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=0.69
cc_138 VPB N_VPWR_c_913_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_914_n 0.0393665f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.675
cc_140 VPB N_VPWR_c_915_n 0.0249166f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_916_n 0.0155666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_917_n 0.0120814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_918_n 0.0196842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_919_n 0.00552821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_920_n 0.00683954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_906_n 0.0854426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_GCLK_c_996_n 0.00390539f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=2.365
cc_148 N_A_78_269#_M1009_g N_GATE_M1011_g 0.0319981f $X=0.51 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_78_269#_c_150_n N_GATE_M1011_g 0.00301404f $X=1.07 $Y=1.645 $X2=0
+ $Y2=0
cc_150 N_A_78_269#_c_158_n N_GATE_M1011_g 0.0175921f $X=1.155 $Y=2.28 $X2=0
+ $Y2=0
cc_151 N_A_78_269#_c_166_p N_GATE_M1011_g 0.00823722f $X=1.24 $Y=2.365 $X2=0
+ $Y2=0
cc_152 N_A_78_269#_c_152_n N_GATE_M1011_g 6.11349e-19 $X=1.59 $Y=1.56 $X2=0
+ $Y2=0
cc_153 N_A_78_269#_c_168_p N_GATE_M1011_g 9.93658e-19 $X=1.71 $Y=2.57 $X2=0
+ $Y2=0
cc_154 N_A_78_269#_c_153_n N_GATE_M1011_g 7.25759e-19 $X=0.555 $Y=1.51 $X2=0
+ $Y2=0
cc_155 N_A_78_269#_c_154_n N_GATE_M1011_g 0.00791881f $X=0.555 $Y=1.51 $X2=0
+ $Y2=0
cc_156 N_A_78_269#_c_171_p N_GATE_M1011_g 0.00738208f $X=1.155 $Y=1.645 $X2=0
+ $Y2=0
cc_157 N_A_78_269#_M1005_g N_GATE_M1020_g 0.0125959f $X=0.525 $Y=0.655 $X2=0
+ $Y2=0
cc_158 N_A_78_269#_c_152_n N_GATE_M1020_g 0.00192177f $X=1.59 $Y=1.56 $X2=0
+ $Y2=0
cc_159 N_A_78_269#_c_155_n N_GATE_M1020_g 7.65149e-19 $X=1.79 $Y=0.69 $X2=0
+ $Y2=0
cc_160 N_A_78_269#_M1005_g GATE 8.80968e-19 $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_161 N_A_78_269#_c_150_n GATE 0.00804716f $X=1.07 $Y=1.645 $X2=0 $Y2=0
cc_162 N_A_78_269#_c_151_n GATE 0.00715399f $X=1.505 $Y=1.645 $X2=0 $Y2=0
cc_163 N_A_78_269#_c_152_n GATE 0.0197864f $X=1.59 $Y=1.56 $X2=0 $Y2=0
cc_164 N_A_78_269#_c_153_n GATE 0.00249585f $X=0.555 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A_78_269#_c_171_p GATE 0.0134753f $X=1.155 $Y=1.645 $X2=0 $Y2=0
cc_166 N_A_78_269#_M1005_g N_GATE_c_257_n 0.00837596f $X=0.525 $Y=0.655 $X2=0
+ $Y2=0
cc_167 N_A_78_269#_c_150_n N_GATE_c_257_n 0.0025f $X=1.07 $Y=1.645 $X2=0 $Y2=0
cc_168 N_A_78_269#_c_151_n N_GATE_c_257_n 0.00142775f $X=1.505 $Y=1.645 $X2=0
+ $Y2=0
cc_169 N_A_78_269#_c_152_n N_GATE_c_257_n 7.98859e-19 $X=1.59 $Y=1.56 $X2=0
+ $Y2=0
cc_170 N_A_78_269#_c_153_n N_GATE_c_257_n 5.53693e-19 $X=0.555 $Y=1.51 $X2=0
+ $Y2=0
cc_171 N_A_78_269#_c_154_n N_GATE_c_257_n 0.00652232f $X=0.555 $Y=1.51 $X2=0
+ $Y2=0
cc_172 N_A_78_269#_c_171_p N_GATE_c_257_n 8.88538e-19 $X=1.155 $Y=1.645 $X2=0
+ $Y2=0
cc_173 N_A_78_269#_c_160_n N_A_284_367#_M1004_g 0.00992484f $X=1.545 $Y=2.365
+ $X2=0 $Y2=0
cc_174 N_A_78_269#_c_168_p N_A_284_367#_M1004_g 0.00453378f $X=1.71 $Y=2.57
+ $X2=0 $Y2=0
cc_175 N_A_78_269#_c_158_n N_A_284_367#_c_314_n 0.0158946f $X=1.155 $Y=2.28
+ $X2=0 $Y2=0
cc_176 N_A_78_269#_c_151_n N_A_284_367#_c_314_n 0.0200427f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_177 N_A_78_269#_c_160_n N_A_284_367#_c_314_n 0.0309082f $X=1.545 $Y=2.365
+ $X2=0 $Y2=0
cc_178 N_A_78_269#_c_158_n N_A_284_367#_c_315_n 0.00463139f $X=1.155 $Y=2.28
+ $X2=0 $Y2=0
cc_179 N_A_78_269#_c_151_n N_A_284_367#_c_315_n 0.00353938f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_180 N_A_78_269#_c_160_n N_A_284_367#_c_315_n 0.00442109f $X=1.545 $Y=2.365
+ $X2=0 $Y2=0
cc_181 N_A_78_269#_c_158_n N_A_284_367#_c_306_n 0.00517133f $X=1.155 $Y=2.28
+ $X2=0 $Y2=0
cc_182 N_A_78_269#_c_151_n N_A_284_367#_c_306_n 0.0132434f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_183 N_A_78_269#_c_152_n N_A_284_367#_c_306_n 0.0206567f $X=1.59 $Y=1.56 $X2=0
+ $Y2=0
cc_184 N_A_78_269#_c_152_n N_A_284_367#_c_309_n 0.0189844f $X=1.59 $Y=1.56 $X2=0
+ $Y2=0
cc_185 N_A_78_269#_c_155_n N_A_284_367#_c_309_n 0.00748297f $X=1.79 $Y=0.69
+ $X2=0 $Y2=0
cc_186 N_A_78_269#_c_152_n N_A_284_367#_c_310_n 0.00235048f $X=1.59 $Y=1.56
+ $X2=0 $Y2=0
cc_187 N_A_78_269#_c_155_n N_A_284_367#_c_310_n 0.00174025f $X=1.79 $Y=0.69
+ $X2=0 $Y2=0
cc_188 N_A_78_269#_c_152_n N_A_284_367#_c_312_n 0.00167714f $X=1.59 $Y=1.56
+ $X2=0 $Y2=0
cc_189 N_A_78_269#_c_155_n N_A_284_367#_c_312_n 0.00454344f $X=1.79 $Y=0.69
+ $X2=0 $Y2=0
cc_190 N_A_78_269#_c_152_n N_A_300_55#_M1015_g 0.0185933f $X=1.59 $Y=1.56 $X2=0
+ $Y2=0
cc_191 N_A_78_269#_c_155_n N_A_300_55#_M1015_g 0.00738586f $X=1.79 $Y=0.69 $X2=0
+ $Y2=0
cc_192 N_A_78_269#_c_151_n N_A_300_55#_c_427_n 0.00122514f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_193 N_A_78_269#_c_152_n N_A_300_55#_c_427_n 0.00189129f $X=1.59 $Y=1.56 $X2=0
+ $Y2=0
cc_194 N_A_78_269#_c_155_n N_A_300_55#_c_427_n 0.00407754f $X=1.79 $Y=0.69 $X2=0
+ $Y2=0
cc_195 N_A_78_269#_c_151_n N_A_300_55#_c_428_n 0.00235018f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_196 N_A_78_269#_c_152_n N_A_300_55#_c_428_n 0.00222637f $X=1.59 $Y=1.56 $X2=0
+ $Y2=0
cc_197 N_A_78_269#_c_160_n N_A_300_55#_M1012_g 0.00278815f $X=1.545 $Y=2.365
+ $X2=0 $Y2=0
cc_198 N_A_78_269#_c_168_p N_A_300_55#_M1012_g 0.00210996f $X=1.71 $Y=2.57 $X2=0
+ $Y2=0
cc_199 N_A_78_269#_c_151_n N_A_300_55#_c_430_n 6.34935e-19 $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_200 N_A_78_269#_M1009_g N_A_33_47#_c_558_n 0.0119166f $X=0.51 $Y=2.465 $X2=0
+ $Y2=0
cc_201 N_A_78_269#_c_166_p N_A_33_47#_c_558_n 0.00470316f $X=1.24 $Y=2.365 $X2=0
+ $Y2=0
cc_202 N_A_78_269#_M1005_g N_A_33_47#_c_541_n 0.0128135f $X=0.525 $Y=0.655 $X2=0
+ $Y2=0
cc_203 N_A_78_269#_c_153_n N_A_33_47#_c_541_n 0.00697521f $X=0.555 $Y=1.51 $X2=0
+ $Y2=0
cc_204 N_A_78_269#_c_154_n N_A_33_47#_c_541_n 4.62581e-19 $X=0.555 $Y=1.51 $X2=0
+ $Y2=0
cc_205 N_A_78_269#_c_155_n N_A_33_47#_c_541_n 0.0102209f $X=1.79 $Y=0.69 $X2=0
+ $Y2=0
cc_206 N_A_78_269#_M1009_g N_A_33_47#_c_575_n 0.0127343f $X=0.51 $Y=2.465 $X2=0
+ $Y2=0
cc_207 N_A_78_269#_c_166_p N_A_33_47#_c_575_n 0.0058194f $X=1.24 $Y=2.365 $X2=0
+ $Y2=0
cc_208 N_A_78_269#_M1005_g N_A_33_47#_c_577_n 9.94468e-19 $X=0.525 $Y=0.655
+ $X2=0 $Y2=0
cc_209 N_A_78_269#_c_155_n N_A_33_47#_c_577_n 0.00317423f $X=1.79 $Y=0.69 $X2=0
+ $Y2=0
cc_210 N_A_78_269#_M1015_d N_A_33_47#_c_542_n 0.0017535f $X=1.65 $Y=0.405 $X2=0
+ $Y2=0
cc_211 N_A_78_269#_c_155_n N_A_33_47#_c_542_n 0.0227298f $X=1.79 $Y=0.69 $X2=0
+ $Y2=0
cc_212 N_A_78_269#_M1004_d N_A_33_47#_c_559_n 0.00269124f $X=1.57 $Y=2.325 $X2=0
+ $Y2=0
cc_213 N_A_78_269#_c_160_n N_A_33_47#_c_559_n 0.00530888f $X=1.545 $Y=2.365
+ $X2=0 $Y2=0
cc_214 N_A_78_269#_c_168_p N_A_33_47#_c_559_n 0.0161646f $X=1.71 $Y=2.57 $X2=0
+ $Y2=0
cc_215 N_A_78_269#_c_168_p N_A_33_47#_c_560_n 0.0160308f $X=1.71 $Y=2.57 $X2=0
+ $Y2=0
cc_216 N_A_78_269#_c_160_n N_A_33_47#_c_585_n 0.00917741f $X=1.545 $Y=2.365
+ $X2=0 $Y2=0
cc_217 N_A_78_269#_c_168_p N_A_33_47#_c_585_n 0.00525351f $X=1.71 $Y=2.57 $X2=0
+ $Y2=0
cc_218 N_A_78_269#_c_155_n N_A_33_47#_c_544_n 0.00503556f $X=1.79 $Y=0.69 $X2=0
+ $Y2=0
cc_219 N_A_78_269#_M1005_g N_A_33_47#_c_549_n 0.00777492f $X=0.525 $Y=0.655
+ $X2=0 $Y2=0
cc_220 N_A_78_269#_c_154_n N_A_33_47#_c_549_n 0.00239053f $X=0.555 $Y=1.51 $X2=0
+ $Y2=0
cc_221 N_A_78_269#_M1009_g N_A_33_47#_c_565_n 0.00450317f $X=0.51 $Y=2.465 $X2=0
+ $Y2=0
cc_222 N_A_78_269#_c_158_n N_A_33_47#_c_565_n 0.00916461f $X=1.155 $Y=2.28 $X2=0
+ $Y2=0
cc_223 N_A_78_269#_M1009_g N_A_33_47#_c_550_n 0.00520322f $X=0.51 $Y=2.465 $X2=0
+ $Y2=0
cc_224 N_A_78_269#_M1005_g N_A_33_47#_c_550_n 0.00484732f $X=0.525 $Y=0.655
+ $X2=0 $Y2=0
cc_225 N_A_78_269#_c_153_n N_A_33_47#_c_550_n 0.0283785f $X=0.555 $Y=1.51 $X2=0
+ $Y2=0
cc_226 N_A_78_269#_c_154_n N_A_33_47#_c_550_n 0.00803689f $X=0.555 $Y=1.51 $X2=0
+ $Y2=0
cc_227 N_A_78_269#_M1009_g N_A_33_47#_c_567_n 9.11509e-19 $X=0.51 $Y=2.465 $X2=0
+ $Y2=0
cc_228 N_A_78_269#_c_160_n N_A_33_47#_c_567_n 0.00391728f $X=1.545 $Y=2.365
+ $X2=0 $Y2=0
cc_229 N_A_78_269#_c_166_p N_A_33_47#_c_567_n 0.00461904f $X=1.24 $Y=2.365 $X2=0
+ $Y2=0
cc_230 N_A_78_269#_c_168_p N_A_33_47#_c_567_n 0.00617018f $X=1.71 $Y=2.57 $X2=0
+ $Y2=0
cc_231 N_A_78_269#_c_155_n N_A_33_47#_c_553_n 2.42734e-19 $X=1.79 $Y=0.69 $X2=0
+ $Y2=0
cc_232 N_A_78_269#_M1009_g N_VPWR_c_917_n 0.00539556f $X=0.51 $Y=2.465 $X2=0
+ $Y2=0
cc_233 N_A_78_269#_M1009_g N_VPWR_c_918_n 0.00408781f $X=0.51 $Y=2.465 $X2=0
+ $Y2=0
cc_234 N_A_78_269#_M1009_g N_VPWR_c_906_n 0.00803284f $X=0.51 $Y=2.465 $X2=0
+ $Y2=0
cc_235 N_A_78_269#_c_160_n A_242_465# 0.00130477f $X=1.545 $Y=2.365 $X2=-0.19
+ $Y2=-0.245
cc_236 N_A_78_269#_M1005_g N_VGND_c_1014_n 0.00937741f $X=0.525 $Y=0.655 $X2=0
+ $Y2=0
cc_237 N_A_78_269#_M1005_g N_VGND_c_1021_n 0.00358185f $X=0.525 $Y=0.655 $X2=0
+ $Y2=0
cc_238 N_A_78_269#_M1005_g N_VGND_c_1028_n 0.00510012f $X=0.525 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_GATE_M1011_g N_A_284_367#_c_314_n 2.46657e-19 $X=1.135 $Y=2.645 $X2=0
+ $Y2=0
cc_240 N_GATE_M1011_g N_A_284_367#_c_315_n 0.0780801f $X=1.135 $Y=2.645 $X2=0
+ $Y2=0
cc_241 N_GATE_M1011_g N_A_284_367#_c_306_n 8.51654e-19 $X=1.135 $Y=2.645 $X2=0
+ $Y2=0
cc_242 N_GATE_M1011_g N_A_300_55#_M1015_g 0.00763377f $X=1.135 $Y=2.645 $X2=0
+ $Y2=0
cc_243 N_GATE_M1020_g N_A_300_55#_M1015_g 0.0707602f $X=1.215 $Y=0.615 $X2=0
+ $Y2=0
cc_244 GATE N_A_300_55#_M1015_g 0.00135589f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_245 N_GATE_M1020_g N_A_33_47#_c_541_n 0.00838281f $X=1.215 $Y=0.615 $X2=0
+ $Y2=0
cc_246 GATE N_A_33_47#_c_541_n 0.0148434f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_247 N_GATE_c_257_n N_A_33_47#_c_541_n 0.00430629f $X=1.125 $Y=1.295 $X2=0
+ $Y2=0
cc_248 N_GATE_M1011_g N_A_33_47#_c_575_n 0.00795544f $X=1.135 $Y=2.645 $X2=0
+ $Y2=0
cc_249 N_GATE_M1020_g N_A_33_47#_c_577_n 0.0072344f $X=1.215 $Y=0.615 $X2=0
+ $Y2=0
cc_250 N_GATE_M1020_g N_A_33_47#_c_542_n 0.00391181f $X=1.215 $Y=0.615 $X2=0
+ $Y2=0
cc_251 N_GATE_M1020_g N_A_33_47#_c_543_n 0.00490977f $X=1.215 $Y=0.615 $X2=0
+ $Y2=0
cc_252 N_GATE_M1020_g N_A_33_47#_c_549_n 0.0011073f $X=1.215 $Y=0.615 $X2=0
+ $Y2=0
cc_253 N_GATE_M1011_g N_A_33_47#_c_565_n 0.00244404f $X=1.135 $Y=2.645 $X2=0
+ $Y2=0
cc_254 GATE N_A_33_47#_c_550_n 0.00527494f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_255 N_GATE_M1011_g N_A_33_47#_c_567_n 0.009875f $X=1.135 $Y=2.645 $X2=0 $Y2=0
cc_256 N_GATE_M1011_g N_VPWR_c_914_n 0.00303969f $X=1.135 $Y=2.645 $X2=0 $Y2=0
cc_257 N_GATE_M1011_g N_VPWR_c_917_n 0.00148161f $X=1.135 $Y=2.645 $X2=0 $Y2=0
cc_258 N_GATE_M1011_g N_VPWR_c_906_n 0.00384886f $X=1.135 $Y=2.645 $X2=0 $Y2=0
cc_259 N_GATE_M1020_g N_VGND_c_1014_n 7.91923e-19 $X=1.215 $Y=0.615 $X2=0 $Y2=0
cc_260 N_GATE_M1020_g N_VGND_c_1019_n 9.47364e-19 $X=1.215 $Y=0.615 $X2=0 $Y2=0
cc_261 N_A_284_367#_c_307_n N_A_300_55#_M1007_s 0.00382602f $X=4.535 $Y=0.61
+ $X2=-0.19 $Y2=-0.245
cc_262 N_A_284_367#_c_317_n N_A_300_55#_M1008_s 0.00935352f $X=4.535 $Y=2.08
+ $X2=0 $Y2=0
cc_263 N_A_284_367#_c_306_n N_A_300_55#_M1015_g 0.00138091f $X=1.94 $Y=1.9 $X2=0
+ $Y2=0
cc_264 N_A_284_367#_c_309_n N_A_300_55#_M1015_g 7.87633e-19 $X=2.025 $Y=1.1
+ $X2=0 $Y2=0
cc_265 N_A_284_367#_c_310_n N_A_300_55#_M1015_g 0.0211502f $X=2.025 $Y=1.1 $X2=0
+ $Y2=0
cc_266 N_A_284_367#_c_312_n N_A_300_55#_M1015_g 0.0146829f $X=2.025 $Y=0.935
+ $X2=0 $Y2=0
cc_267 N_A_284_367#_c_314_n N_A_300_55#_c_427_n 0.00370836f $X=1.855 $Y=2.005
+ $X2=0 $Y2=0
cc_268 N_A_284_367#_c_306_n N_A_300_55#_c_427_n 0.00656077f $X=1.94 $Y=1.9 $X2=0
+ $Y2=0
cc_269 N_A_284_367#_c_310_n N_A_300_55#_c_427_n 0.0220347f $X=2.025 $Y=1.1 $X2=0
+ $Y2=0
cc_270 N_A_284_367#_c_315_n N_A_300_55#_c_428_n 0.0159721f $X=1.585 $Y=2 $X2=0
+ $Y2=0
cc_271 N_A_284_367#_M1004_g N_A_300_55#_M1012_g 0.0141137f $X=1.495 $Y=2.645
+ $X2=0 $Y2=0
cc_272 N_A_284_367#_c_315_n N_A_300_55#_M1012_g 0.0214509f $X=1.585 $Y=2 $X2=0
+ $Y2=0
cc_273 N_A_284_367#_c_306_n N_A_300_55#_M1012_g 0.00481585f $X=1.94 $Y=1.9 $X2=0
+ $Y2=0
cc_274 N_A_284_367#_c_319_n N_A_300_55#_M1012_g 0.00674783f $X=1.94 $Y=2.005
+ $X2=0 $Y2=0
cc_275 N_A_284_367#_c_320_n N_A_300_55#_M1012_g 0.00904413f $X=3.07 $Y=2.052
+ $X2=0 $Y2=0
cc_276 N_A_284_367#_c_320_n N_A_300_55#_M1001_g 0.0100869f $X=3.07 $Y=2.052
+ $X2=0 $Y2=0
cc_277 N_A_284_367#_c_321_n N_A_300_55#_M1001_g 0.00456473f $X=3.4 $Y=2.052
+ $X2=0 $Y2=0
cc_278 N_A_284_367#_c_306_n N_A_300_55#_c_430_n 0.0114196f $X=1.94 $Y=1.9 $X2=0
+ $Y2=0
cc_279 N_A_284_367#_c_309_n N_A_300_55#_c_430_n 8.0425e-19 $X=2.025 $Y=1.1 $X2=0
+ $Y2=0
cc_280 N_A_284_367#_c_311_n N_A_300_55#_c_431_n 0.00290535f $X=3.4 $Y=0.59 $X2=0
+ $Y2=0
cc_281 N_A_284_367#_c_321_n N_A_300_55#_c_433_n 0.00213336f $X=3.4 $Y=2.052
+ $X2=0 $Y2=0
cc_282 N_A_284_367#_c_306_n N_A_300_55#_c_434_n 0.0205861f $X=1.94 $Y=1.9 $X2=0
+ $Y2=0
cc_283 N_A_284_367#_c_320_n N_A_300_55#_c_434_n 0.080021f $X=3.07 $Y=2.052 $X2=0
+ $Y2=0
cc_284 N_A_284_367#_c_320_n N_A_300_55#_c_435_n 0.00839692f $X=3.07 $Y=2.052
+ $X2=0 $Y2=0
cc_285 N_A_284_367#_c_311_n N_A_300_55#_c_436_n 9.74602e-19 $X=3.4 $Y=0.59 $X2=0
+ $Y2=0
cc_286 N_A_284_367#_c_307_n N_A_300_55#_c_437_n 0.0206039f $X=4.535 $Y=0.61
+ $X2=0 $Y2=0
cc_287 N_A_284_367#_c_308_n N_A_300_55#_c_437_n 0.0149338f $X=4.62 $Y=1.985
+ $X2=0 $Y2=0
cc_288 N_A_284_367#_c_311_n N_A_300_55#_c_437_n 0.0577152f $X=3.4 $Y=0.59 $X2=0
+ $Y2=0
cc_289 N_A_284_367#_c_311_n N_A_300_55#_c_438_n 0.0110779f $X=3.4 $Y=0.59 $X2=0
+ $Y2=0
cc_290 N_A_284_367#_c_317_n N_A_300_55#_c_439_n 0.02698f $X=4.535 $Y=2.08 $X2=0
+ $Y2=0
cc_291 N_A_284_367#_c_308_n N_A_300_55#_c_439_n 0.0557675f $X=4.62 $Y=1.985
+ $X2=0 $Y2=0
cc_292 N_A_284_367#_c_320_n N_A_33_47#_M1014_g 0.00166227f $X=3.07 $Y=2.052
+ $X2=0 $Y2=0
cc_293 N_A_284_367#_c_309_n N_A_33_47#_c_542_n 0.00538167f $X=2.025 $Y=1.1 $X2=0
+ $Y2=0
cc_294 N_A_284_367#_c_310_n N_A_33_47#_c_542_n 0.00176436f $X=2.025 $Y=1.1 $X2=0
+ $Y2=0
cc_295 N_A_284_367#_c_312_n N_A_33_47#_c_542_n 0.0119571f $X=2.025 $Y=0.935
+ $X2=0 $Y2=0
cc_296 N_A_284_367#_M1004_g N_A_33_47#_c_559_n 0.0110279f $X=1.495 $Y=2.645
+ $X2=0 $Y2=0
cc_297 N_A_284_367#_M1004_g N_A_33_47#_c_560_n 9.58749e-19 $X=1.495 $Y=2.645
+ $X2=0 $Y2=0
cc_298 N_A_284_367#_M1001_d N_A_33_47#_c_618_n 0.00495522f $X=3.095 $Y=1.955
+ $X2=0 $Y2=0
cc_299 N_A_284_367#_c_320_n N_A_33_47#_c_618_n 0.0449883f $X=3.07 $Y=2.052 $X2=0
+ $Y2=0
cc_300 N_A_284_367#_c_321_n N_A_33_47#_c_618_n 0.0153371f $X=3.4 $Y=2.052 $X2=0
+ $Y2=0
cc_301 N_A_284_367#_c_319_n N_A_33_47#_c_585_n 0.00192273f $X=1.94 $Y=2.005
+ $X2=0 $Y2=0
cc_302 N_A_284_367#_c_320_n N_A_33_47#_c_585_n 0.00665659f $X=3.07 $Y=2.052
+ $X2=0 $Y2=0
cc_303 N_A_284_367#_c_312_n N_A_33_47#_c_544_n 0.00299571f $X=2.025 $Y=0.935
+ $X2=0 $Y2=0
cc_304 N_A_284_367#_M1001_d N_A_33_47#_c_561_n 0.00123821f $X=3.095 $Y=1.955
+ $X2=0 $Y2=0
cc_305 N_A_284_367#_c_321_n N_A_33_47#_c_562_n 9.71528e-19 $X=3.4 $Y=2.052 $X2=0
+ $Y2=0
cc_306 N_A_284_367#_c_317_n N_A_33_47#_c_563_n 0.0688814f $X=4.535 $Y=2.08 $X2=0
+ $Y2=0
cc_307 N_A_284_367#_c_317_n N_A_33_47#_c_545_n 0.015458f $X=4.535 $Y=2.08 $X2=0
+ $Y2=0
cc_308 N_A_284_367#_c_308_n N_A_33_47#_c_545_n 0.0319848f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_309 N_A_284_367#_c_308_n N_A_33_47#_c_546_n 0.014562f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_310 N_A_284_367#_M1004_g N_A_33_47#_c_567_n 0.00274753f $X=1.495 $Y=2.645
+ $X2=0 $Y2=0
cc_311 N_A_284_367#_c_309_n N_A_33_47#_c_551_n 0.0200227f $X=2.025 $Y=1.1 $X2=0
+ $Y2=0
cc_312 N_A_284_367#_c_310_n N_A_33_47#_c_551_n 0.00273979f $X=2.025 $Y=1.1 $X2=0
+ $Y2=0
cc_313 N_A_284_367#_c_309_n N_A_33_47#_c_552_n 2.85696e-19 $X=2.025 $Y=1.1 $X2=0
+ $Y2=0
cc_314 N_A_284_367#_c_310_n N_A_33_47#_c_552_n 0.0212408f $X=2.025 $Y=1.1 $X2=0
+ $Y2=0
cc_315 N_A_284_367#_M1001_d N_A_33_47#_c_568_n 9.22636e-19 $X=3.095 $Y=1.955
+ $X2=0 $Y2=0
cc_316 N_A_284_367#_c_321_n N_A_33_47#_c_568_n 0.0280002f $X=3.4 $Y=2.052 $X2=0
+ $Y2=0
cc_317 N_A_284_367#_c_312_n N_A_33_47#_c_553_n 0.0233881f $X=2.025 $Y=0.935
+ $X2=0 $Y2=0
cc_318 N_A_284_367#_c_307_n N_CLK_c_768_n 9.64994e-19 $X=4.535 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_319 N_A_284_367#_c_317_n N_CLK_c_768_n 0.00613778f $X=4.535 $Y=2.08 $X2=-0.19
+ $Y2=-0.245
cc_320 N_A_284_367#_c_307_n N_CLK_M1007_g 0.0131825f $X=4.535 $Y=0.61 $X2=0
+ $Y2=0
cc_321 N_A_284_367#_c_308_n N_CLK_M1007_g 0.00806457f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_322 N_A_284_367#_c_317_n N_CLK_c_775_n 0.0144663f $X=4.535 $Y=2.08 $X2=0
+ $Y2=0
cc_323 N_A_284_367#_c_308_n N_CLK_c_775_n 0.011056f $X=4.62 $Y=1.985 $X2=0 $Y2=0
cc_324 N_A_284_367#_c_307_n N_CLK_M1006_g 0.00480287f $X=4.535 $Y=0.61 $X2=0
+ $Y2=0
cc_325 N_A_284_367#_c_308_n N_CLK_M1006_g 0.0103138f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_326 N_A_284_367#_c_307_n N_CLK_c_771_n 0.00145588f $X=4.535 $Y=0.61 $X2=0
+ $Y2=0
cc_327 N_A_284_367#_c_317_n N_CLK_c_771_n 0.00207697f $X=4.535 $Y=2.08 $X2=0
+ $Y2=0
cc_328 N_A_284_367#_c_308_n N_CLK_c_771_n 0.0180321f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_329 N_A_284_367#_c_317_n N_CLK_c_772_n 0.00196379f $X=4.535 $Y=2.08 $X2=0
+ $Y2=0
cc_330 N_A_284_367#_c_317_n N_CLK_c_773_n 0.0266999f $X=4.535 $Y=2.08 $X2=0
+ $Y2=0
cc_331 N_A_284_367#_c_308_n N_A_1039_367#_c_838_n 0.0120944f $X=4.62 $Y=1.985
+ $X2=0 $Y2=0
cc_332 N_A_284_367#_c_320_n N_VPWR_M1014_d 0.00530608f $X=3.07 $Y=2.052 $X2=0
+ $Y2=0
cc_333 N_A_284_367#_c_317_n N_VPWR_M1008_d 0.00223357f $X=4.535 $Y=2.08 $X2=0
+ $Y2=0
cc_334 N_A_284_367#_c_308_n N_VPWR_M1008_d 0.00133183f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A_284_367#_M1004_g N_VPWR_c_914_n 0.0028086f $X=1.495 $Y=2.645 $X2=0
+ $Y2=0
cc_336 N_A_284_367#_M1004_g N_VPWR_c_906_n 0.0037128f $X=1.495 $Y=2.645 $X2=0
+ $Y2=0
cc_337 N_A_284_367#_c_307_n N_VGND_M1007_d 0.00881317f $X=4.535 $Y=0.61 $X2=0
+ $Y2=0
cc_338 N_A_284_367#_c_308_n N_VGND_M1007_d 0.0125912f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_A_284_367#_c_312_n N_VGND_c_1019_n 9.29198e-19 $X=2.025 $Y=0.935 $X2=0
+ $Y2=0
cc_340 N_A_284_367#_c_307_n N_VGND_c_1022_n 0.0244094f $X=4.535 $Y=0.61 $X2=0
+ $Y2=0
cc_341 N_A_284_367#_c_311_n N_VGND_c_1022_n 0.00781724f $X=3.4 $Y=0.59 $X2=0
+ $Y2=0
cc_342 N_A_284_367#_c_307_n N_VGND_c_1026_n 0.0195949f $X=4.535 $Y=0.61 $X2=0
+ $Y2=0
cc_343 N_A_284_367#_c_307_n N_VGND_c_1028_n 0.0340238f $X=4.535 $Y=0.61 $X2=0
+ $Y2=0
cc_344 N_A_284_367#_c_311_n N_VGND_c_1028_n 0.0106224f $X=3.4 $Y=0.59 $X2=0
+ $Y2=0
cc_345 N_A_300_55#_M1012_g N_A_33_47#_M1014_g 0.0417764f $X=2.035 $Y=2.535 $X2=0
+ $Y2=0
cc_346 N_A_300_55#_M1001_g N_A_33_47#_M1014_g 0.0142716f $X=3.02 $Y=2.275 $X2=0
+ $Y2=0
cc_347 N_A_300_55#_c_435_n N_A_33_47#_M1014_g 0.00388244f $X=2.37 $Y=1.64 $X2=0
+ $Y2=0
cc_348 N_A_300_55#_M1001_g N_A_33_47#_c_555_n 0.00804766f $X=3.02 $Y=2.275 $X2=0
+ $Y2=0
cc_349 N_A_300_55#_M1015_g N_A_33_47#_c_541_n 4.87617e-19 $X=1.575 $Y=0.615
+ $X2=0 $Y2=0
cc_350 N_A_300_55#_M1015_g N_A_33_47#_c_577_n 0.00122125f $X=1.575 $Y=0.615
+ $X2=0 $Y2=0
cc_351 N_A_300_55#_M1015_g N_A_33_47#_c_542_n 0.00981172f $X=1.575 $Y=0.615
+ $X2=0 $Y2=0
cc_352 N_A_300_55#_M1012_g N_A_33_47#_c_559_n 0.00167267f $X=2.035 $Y=2.535
+ $X2=0 $Y2=0
cc_353 N_A_300_55#_M1012_g N_A_33_47#_c_560_n 0.0104034f $X=2.035 $Y=2.535 $X2=0
+ $Y2=0
cc_354 N_A_300_55#_M1001_g N_A_33_47#_c_618_n 0.0129483f $X=3.02 $Y=2.275 $X2=0
+ $Y2=0
cc_355 N_A_300_55#_M1012_g N_A_33_47#_c_585_n 0.00626149f $X=2.035 $Y=2.535
+ $X2=0 $Y2=0
cc_356 N_A_300_55#_c_431_n N_A_33_47#_c_544_n 8.35117e-19 $X=3.11 $Y=0.935 $X2=0
+ $Y2=0
cc_357 N_A_300_55#_c_438_n N_A_33_47#_c_544_n 0.00187538f $X=3.235 $Y=0.97 $X2=0
+ $Y2=0
cc_358 N_A_300_55#_M1001_g N_A_33_47#_c_561_n 0.00666784f $X=3.02 $Y=2.275 $X2=0
+ $Y2=0
cc_359 N_A_300_55#_M1008_s N_A_33_47#_c_563_n 0.00522589f $X=4.055 $Y=1.605
+ $X2=0 $Y2=0
cc_360 N_A_300_55#_c_434_n N_A_33_47#_c_551_n 0.0241582f $X=3.025 $Y=1.617 $X2=0
+ $Y2=0
cc_361 N_A_300_55#_c_435_n N_A_33_47#_c_551_n 0.00135988f $X=2.37 $Y=1.64 $X2=0
+ $Y2=0
cc_362 N_A_300_55#_c_507_p N_A_33_47#_c_551_n 0.00935852f $X=3.11 $Y=1.1 $X2=0
+ $Y2=0
cc_363 N_A_300_55#_c_436_n N_A_33_47#_c_551_n 0.00122103f $X=3.11 $Y=1.1 $X2=0
+ $Y2=0
cc_364 N_A_300_55#_c_438_n N_A_33_47#_c_551_n 0.00668987f $X=3.235 $Y=0.97 $X2=0
+ $Y2=0
cc_365 N_A_300_55#_c_434_n N_A_33_47#_c_552_n 0.00492068f $X=3.025 $Y=1.617
+ $X2=0 $Y2=0
cc_366 N_A_300_55#_c_435_n N_A_33_47#_c_552_n 0.00874203f $X=2.37 $Y=1.64 $X2=0
+ $Y2=0
cc_367 N_A_300_55#_c_507_p N_A_33_47#_c_552_n 2.23733e-19 $X=3.11 $Y=1.1 $X2=0
+ $Y2=0
cc_368 N_A_300_55#_c_436_n N_A_33_47#_c_552_n 0.0201592f $X=3.11 $Y=1.1 $X2=0
+ $Y2=0
cc_369 N_A_300_55#_c_431_n N_A_33_47#_c_553_n 0.011225f $X=3.11 $Y=0.935 $X2=0
+ $Y2=0
cc_370 N_A_300_55#_c_439_n N_CLK_c_768_n 0.0158584f $X=4.2 $Y=1.73 $X2=-0.19
+ $Y2=-0.245
cc_371 N_A_300_55#_c_437_n N_CLK_M1007_g 0.00981749f $X=4.035 $Y=0.97 $X2=0
+ $Y2=0
cc_372 N_A_300_55#_c_439_n N_CLK_M1007_g 0.0111709f $X=4.2 $Y=1.73 $X2=0 $Y2=0
cc_373 N_A_300_55#_c_439_n N_CLK_c_771_n 0.0112921f $X=4.2 $Y=1.73 $X2=0 $Y2=0
cc_374 N_A_300_55#_M1001_g N_CLK_c_772_n 0.00269336f $X=3.02 $Y=2.275 $X2=0
+ $Y2=0
cc_375 N_A_300_55#_c_432_n N_CLK_c_772_n 0.0126117f $X=3.11 $Y=1.44 $X2=0 $Y2=0
cc_376 N_A_300_55#_c_434_n N_CLK_c_772_n 5.29933e-19 $X=3.025 $Y=1.617 $X2=0
+ $Y2=0
cc_377 N_A_300_55#_c_507_p N_CLK_c_772_n 5.68609e-19 $X=3.11 $Y=1.1 $X2=0 $Y2=0
cc_378 N_A_300_55#_c_437_n N_CLK_c_772_n 0.0125466f $X=4.035 $Y=0.97 $X2=0 $Y2=0
cc_379 N_A_300_55#_c_439_n N_CLK_c_772_n 0.00182721f $X=4.2 $Y=1.73 $X2=0 $Y2=0
cc_380 N_A_300_55#_M1001_g N_CLK_c_773_n 5.87481e-19 $X=3.02 $Y=2.275 $X2=0
+ $Y2=0
cc_381 N_A_300_55#_c_433_n N_CLK_c_773_n 9.73903e-19 $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_382 N_A_300_55#_c_434_n N_CLK_c_773_n 0.0222245f $X=3.025 $Y=1.617 $X2=0
+ $Y2=0
cc_383 N_A_300_55#_c_507_p N_CLK_c_773_n 0.00100574f $X=3.11 $Y=1.1 $X2=0 $Y2=0
cc_384 N_A_300_55#_c_437_n N_CLK_c_773_n 0.0167215f $X=4.035 $Y=0.97 $X2=0 $Y2=0
cc_385 N_A_300_55#_c_439_n N_CLK_c_773_n 0.0221147f $X=4.2 $Y=1.73 $X2=0 $Y2=0
cc_386 N_A_300_55#_M1001_g N_VPWR_c_907_n 5.6275e-19 $X=3.02 $Y=2.275 $X2=0
+ $Y2=0
cc_387 N_A_300_55#_M1012_g N_VPWR_c_914_n 4.98428e-19 $X=2.035 $Y=2.535 $X2=0
+ $Y2=0
cc_388 N_A_300_55#_M1001_g N_VPWR_c_906_n 8.50993e-19 $X=3.02 $Y=2.275 $X2=0
+ $Y2=0
cc_389 N_A_300_55#_c_431_n N_VGND_c_1015_n 0.00333698f $X=3.11 $Y=0.935 $X2=0
+ $Y2=0
cc_390 N_A_300_55#_M1015_g N_VGND_c_1019_n 9.29198e-19 $X=1.575 $Y=0.615 $X2=0
+ $Y2=0
cc_391 N_A_300_55#_c_431_n N_VGND_c_1022_n 0.00528195f $X=3.11 $Y=0.935 $X2=0
+ $Y2=0
cc_392 N_A_300_55#_c_431_n N_VGND_c_1028_n 0.00534666f $X=3.11 $Y=0.935 $X2=0
+ $Y2=0
cc_393 N_A_33_47#_c_563_n N_CLK_c_775_n 0.0142003f $X=4.875 $Y=2.43 $X2=0 $Y2=0
cc_394 N_A_33_47#_c_545_n N_CLK_c_775_n 0.00459604f $X=4.96 $Y=2.345 $X2=0 $Y2=0
cc_395 N_A_33_47#_M1002_g N_CLK_M1006_g 0.0509103f $X=5.295 $Y=0.875 $X2=0 $Y2=0
cc_396 N_A_33_47#_c_546_n N_CLK_M1006_g 0.008001f $X=5.045 $Y=1.44 $X2=0 $Y2=0
cc_397 N_A_33_47#_c_548_n N_CLK_M1006_g 0.00596905f $X=5.57 $Y=1.44 $X2=0 $Y2=0
cc_398 N_A_33_47#_c_563_n N_CLK_c_776_n 0.00241254f $X=4.875 $Y=2.43 $X2=0 $Y2=0
cc_399 N_A_33_47#_c_545_n N_CLK_c_776_n 0.00461878f $X=4.96 $Y=2.345 $X2=0 $Y2=0
cc_400 N_A_33_47#_M1016_g N_CLK_c_771_n 0.0115388f $X=5.645 $Y=2.155 $X2=0 $Y2=0
cc_401 N_A_33_47#_c_563_n N_CLK_c_771_n 0.00430323f $X=4.875 $Y=2.43 $X2=0 $Y2=0
cc_402 N_A_33_47#_c_545_n N_CLK_c_771_n 0.0105997f $X=4.96 $Y=2.345 $X2=0 $Y2=0
cc_403 N_A_33_47#_c_546_n N_CLK_c_771_n 0.00662821f $X=5.045 $Y=1.44 $X2=0 $Y2=0
cc_404 N_A_33_47#_c_547_n N_CLK_c_771_n 0.00723293f $X=5.57 $Y=1.44 $X2=0 $Y2=0
cc_405 N_A_33_47#_c_548_n N_CLK_c_771_n 0.00221954f $X=5.57 $Y=1.44 $X2=0 $Y2=0
cc_406 N_A_33_47#_c_548_n N_A_1039_367#_M1003_g 0.00306925f $X=5.57 $Y=1.44
+ $X2=0 $Y2=0
cc_407 N_A_33_47#_M1016_g N_A_1039_367#_M1010_g 0.0167919f $X=5.645 $Y=2.155
+ $X2=0 $Y2=0
cc_408 N_A_33_47#_M1016_g N_A_1039_367#_c_842_n 2.02e-19 $X=5.645 $Y=2.155 $X2=0
+ $Y2=0
cc_409 N_A_33_47#_c_563_n N_A_1039_367#_c_842_n 0.00711422f $X=4.875 $Y=2.43
+ $X2=0 $Y2=0
cc_410 N_A_33_47#_M1016_g N_A_1039_367#_c_843_n 0.0154684f $X=5.645 $Y=2.155
+ $X2=0 $Y2=0
cc_411 N_A_33_47#_c_547_n N_A_1039_367#_c_843_n 0.0127408f $X=5.57 $Y=1.44 $X2=0
+ $Y2=0
cc_412 N_A_33_47#_c_548_n N_A_1039_367#_c_843_n 8.79541e-19 $X=5.57 $Y=1.44
+ $X2=0 $Y2=0
cc_413 N_A_33_47#_c_545_n N_A_1039_367#_c_844_n 0.0108128f $X=4.96 $Y=2.345
+ $X2=0 $Y2=0
cc_414 N_A_33_47#_c_547_n N_A_1039_367#_c_844_n 0.0279523f $X=5.57 $Y=1.44 $X2=0
+ $Y2=0
cc_415 N_A_33_47#_c_548_n N_A_1039_367#_c_844_n 0.00477596f $X=5.57 $Y=1.44
+ $X2=0 $Y2=0
cc_416 N_A_33_47#_M1002_g N_A_1039_367#_c_836_n 3.58849e-19 $X=5.295 $Y=0.875
+ $X2=0 $Y2=0
cc_417 N_A_33_47#_c_547_n N_A_1039_367#_c_836_n 0.00432592f $X=5.57 $Y=1.44
+ $X2=0 $Y2=0
cc_418 N_A_33_47#_c_548_n N_A_1039_367#_c_836_n 0.00178875f $X=5.57 $Y=1.44
+ $X2=0 $Y2=0
cc_419 N_A_33_47#_M1002_g N_A_1039_367#_c_837_n 9.17231e-19 $X=5.295 $Y=0.875
+ $X2=0 $Y2=0
cc_420 N_A_33_47#_M1016_g N_A_1039_367#_c_837_n 0.00111372f $X=5.645 $Y=2.155
+ $X2=0 $Y2=0
cc_421 N_A_33_47#_c_547_n N_A_1039_367#_c_837_n 0.0124122f $X=5.57 $Y=1.44 $X2=0
+ $Y2=0
cc_422 N_A_33_47#_c_548_n N_A_1039_367#_c_837_n 0.00388871f $X=5.57 $Y=1.44
+ $X2=0 $Y2=0
cc_423 N_A_33_47#_M1002_g N_A_1039_367#_c_838_n 0.0115925f $X=5.295 $Y=0.875
+ $X2=0 $Y2=0
cc_424 N_A_33_47#_c_547_n N_A_1039_367#_c_838_n 0.0257009f $X=5.57 $Y=1.44 $X2=0
+ $Y2=0
cc_425 N_A_33_47#_c_548_n N_A_1039_367#_c_838_n 0.00867898f $X=5.57 $Y=1.44
+ $X2=0 $Y2=0
cc_426 N_A_33_47#_M1016_g N_A_1039_367#_c_839_n 0.00420555f $X=5.645 $Y=2.155
+ $X2=0 $Y2=0
cc_427 N_A_33_47#_c_547_n N_A_1039_367#_c_839_n 7.39521e-19 $X=5.57 $Y=1.44
+ $X2=0 $Y2=0
cc_428 N_A_33_47#_c_548_n N_A_1039_367#_c_839_n 0.0173543f $X=5.57 $Y=1.44 $X2=0
+ $Y2=0
cc_429 N_A_33_47#_c_575_n N_VPWR_M1009_d 0.0186075f $X=1.15 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_430 N_A_33_47#_c_618_n N_VPWR_M1014_d 0.00917229f $X=3.335 $Y=2.43 $X2=0
+ $Y2=0
cc_431 N_A_33_47#_c_563_n N_VPWR_M1008_d 0.00822345f $X=4.875 $Y=2.43 $X2=0
+ $Y2=0
cc_432 N_A_33_47#_c_545_n N_VPWR_M1008_d 0.00778991f $X=4.96 $Y=2.345 $X2=0
+ $Y2=0
cc_433 N_A_33_47#_M1014_g N_VPWR_c_907_n 0.0067943f $X=2.395 $Y=2.535 $X2=0
+ $Y2=0
cc_434 N_A_33_47#_c_555_n N_VPWR_c_907_n 0.024517f $X=3.335 $Y=3.055 $X2=0 $Y2=0
cc_435 N_A_33_47#_c_559_n N_VPWR_c_907_n 0.00795027f $X=1.995 $Y=2.99 $X2=0
+ $Y2=0
cc_436 N_A_33_47#_c_560_n N_VPWR_c_907_n 0.00830158f $X=2.08 $Y=2.905 $X2=0
+ $Y2=0
cc_437 N_A_33_47#_c_618_n N_VPWR_c_907_n 0.0260418f $X=3.335 $Y=2.43 $X2=0 $Y2=0
cc_438 N_A_33_47#_c_561_n N_VPWR_c_907_n 0.0150306f $X=3.5 $Y=2.94 $X2=0 $Y2=0
cc_439 N_A_33_47#_c_562_n N_VPWR_c_907_n 0.0038529f $X=3.5 $Y=2.94 $X2=0 $Y2=0
cc_440 N_A_33_47#_c_563_n N_VPWR_c_908_n 0.0270429f $X=4.875 $Y=2.43 $X2=0 $Y2=0
cc_441 N_A_33_47#_M1016_g N_VPWR_c_909_n 0.00627301f $X=5.645 $Y=2.155 $X2=0
+ $Y2=0
cc_442 N_A_33_47#_c_555_n N_VPWR_c_912_n 0.0196597f $X=3.335 $Y=3.055 $X2=0
+ $Y2=0
cc_443 N_A_33_47#_c_561_n N_VPWR_c_912_n 0.0223605f $X=3.5 $Y=2.94 $X2=0 $Y2=0
cc_444 N_A_33_47#_c_556_n N_VPWR_c_914_n 0.00788956f $X=2.47 $Y=3.055 $X2=0
+ $Y2=0
cc_445 N_A_33_47#_c_575_n N_VPWR_c_914_n 0.00338574f $X=1.15 $Y=2.715 $X2=0
+ $Y2=0
cc_446 N_A_33_47#_c_559_n N_VPWR_c_914_n 0.0552033f $X=1.995 $Y=2.99 $X2=0 $Y2=0
cc_447 N_A_33_47#_c_567_n N_VPWR_c_914_n 0.0114718f $X=1.235 $Y=2.715 $X2=0
+ $Y2=0
cc_448 N_A_33_47#_M1016_g N_VPWR_c_915_n 0.00312414f $X=5.645 $Y=2.155 $X2=0
+ $Y2=0
cc_449 N_A_33_47#_c_575_n N_VPWR_c_917_n 0.0240513f $X=1.15 $Y=2.715 $X2=0 $Y2=0
cc_450 N_A_33_47#_c_567_n N_VPWR_c_917_n 0.00759507f $X=1.235 $Y=2.715 $X2=0
+ $Y2=0
cc_451 N_A_33_47#_c_558_n N_VPWR_c_918_n 0.00770305f $X=0.29 $Y=2.63 $X2=0 $Y2=0
cc_452 N_A_33_47#_c_575_n N_VPWR_c_918_n 0.00335382f $X=1.15 $Y=2.715 $X2=0
+ $Y2=0
cc_453 N_A_33_47#_M1009_s N_VPWR_c_906_n 0.00272491f $X=0.17 $Y=1.835 $X2=0
+ $Y2=0
cc_454 N_A_33_47#_c_555_n N_VPWR_c_906_n 0.0156986f $X=3.335 $Y=3.055 $X2=0
+ $Y2=0
cc_455 N_A_33_47#_c_556_n N_VPWR_c_906_n 0.00548813f $X=2.47 $Y=3.055 $X2=0
+ $Y2=0
cc_456 N_A_33_47#_M1016_g N_VPWR_c_906_n 0.00410284f $X=5.645 $Y=2.155 $X2=0
+ $Y2=0
cc_457 N_A_33_47#_c_558_n N_VPWR_c_906_n 0.0109878f $X=0.29 $Y=2.63 $X2=0 $Y2=0
cc_458 N_A_33_47#_c_575_n N_VPWR_c_906_n 0.0119321f $X=1.15 $Y=2.715 $X2=0 $Y2=0
cc_459 N_A_33_47#_c_559_n N_VPWR_c_906_n 0.0313011f $X=1.995 $Y=2.99 $X2=0 $Y2=0
cc_460 N_A_33_47#_c_618_n N_VPWR_c_906_n 0.0271182f $X=3.335 $Y=2.43 $X2=0 $Y2=0
cc_461 N_A_33_47#_c_561_n N_VPWR_c_906_n 0.0112511f $X=3.5 $Y=2.94 $X2=0 $Y2=0
cc_462 N_A_33_47#_c_562_n N_VPWR_c_906_n 0.00851462f $X=3.5 $Y=2.94 $X2=0 $Y2=0
cc_463 N_A_33_47#_c_563_n N_VPWR_c_906_n 0.0380529f $X=4.875 $Y=2.43 $X2=0 $Y2=0
cc_464 N_A_33_47#_c_567_n N_VPWR_c_906_n 0.00619154f $X=1.235 $Y=2.715 $X2=0
+ $Y2=0
cc_465 N_A_33_47#_c_559_n A_242_465# 8.78902e-19 $X=1.995 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_466 N_A_33_47#_c_567_n A_242_465# 0.00401868f $X=1.235 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_467 N_A_33_47#_c_618_n A_422_465# 0.00294039f $X=3.335 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_468 N_A_33_47#_c_541_n N_VGND_M1005_d 0.0137346f $X=1.075 $Y=0.75 $X2=-0.19
+ $Y2=-0.245
cc_469 N_A_33_47#_c_577_n N_VGND_M1005_d 0.0033033f $X=1.165 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_470 N_A_33_47#_c_543_n N_VGND_M1005_d 2.93339e-19 $X=1.255 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_471 N_A_33_47#_c_541_n N_VGND_c_1014_n 0.0206911f $X=1.075 $Y=0.75 $X2=0
+ $Y2=0
cc_472 N_A_33_47#_c_577_n N_VGND_c_1014_n 0.00456739f $X=1.165 $Y=0.665 $X2=0
+ $Y2=0
cc_473 N_A_33_47#_c_543_n N_VGND_c_1014_n 0.0149379f $X=1.255 $Y=0.35 $X2=0
+ $Y2=0
cc_474 N_A_33_47#_c_542_n N_VGND_c_1015_n 0.0137f $X=2.36 $Y=0.35 $X2=0 $Y2=0
cc_475 N_A_33_47#_c_544_n N_VGND_c_1015_n 0.0233354f $X=2.445 $Y=0.935 $X2=0
+ $Y2=0
cc_476 N_A_33_47#_c_551_n N_VGND_c_1015_n 0.00239484f $X=2.565 $Y=1.1 $X2=0
+ $Y2=0
cc_477 N_A_33_47#_c_552_n N_VGND_c_1015_n 6.75574e-19 $X=2.565 $Y=1.1 $X2=0
+ $Y2=0
cc_478 N_A_33_47#_c_553_n N_VGND_c_1015_n 0.0034436f $X=2.565 $Y=0.935 $X2=0
+ $Y2=0
cc_479 N_A_33_47#_M1002_g N_VGND_c_1016_n 0.00425581f $X=5.295 $Y=0.875 $X2=0
+ $Y2=0
cc_480 N_A_33_47#_c_541_n N_VGND_c_1019_n 0.00276529f $X=1.075 $Y=0.75 $X2=0
+ $Y2=0
cc_481 N_A_33_47#_c_542_n N_VGND_c_1019_n 0.0783961f $X=2.36 $Y=0.35 $X2=0 $Y2=0
cc_482 N_A_33_47#_c_543_n N_VGND_c_1019_n 0.0119765f $X=1.255 $Y=0.35 $X2=0
+ $Y2=0
cc_483 N_A_33_47#_c_553_n N_VGND_c_1019_n 0.00154062f $X=2.565 $Y=0.935 $X2=0
+ $Y2=0
cc_484 N_A_33_47#_c_540_n N_VGND_c_1021_n 0.0195758f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_485 N_A_33_47#_c_541_n N_VGND_c_1021_n 0.00182048f $X=1.075 $Y=0.75 $X2=0
+ $Y2=0
cc_486 N_A_33_47#_c_549_n N_VGND_c_1021_n 4.73146e-19 $X=0.287 $Y=0.75 $X2=0
+ $Y2=0
cc_487 N_A_33_47#_M1002_g N_VGND_c_1023_n 0.00381268f $X=5.295 $Y=0.875 $X2=0
+ $Y2=0
cc_488 N_A_33_47#_M1005_s N_VGND_c_1028_n 0.00248746f $X=0.165 $Y=0.235 $X2=0
+ $Y2=0
cc_489 N_A_33_47#_M1002_g N_VGND_c_1028_n 0.00458517f $X=5.295 $Y=0.875 $X2=0
+ $Y2=0
cc_490 N_A_33_47#_c_540_n N_VGND_c_1028_n 0.0110024f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_491 N_A_33_47#_c_541_n N_VGND_c_1028_n 0.00894579f $X=1.075 $Y=0.75 $X2=0
+ $Y2=0
cc_492 N_A_33_47#_c_542_n N_VGND_c_1028_n 0.0478642f $X=2.36 $Y=0.35 $X2=0 $Y2=0
cc_493 N_A_33_47#_c_543_n N_VGND_c_1028_n 0.00693168f $X=1.255 $Y=0.35 $X2=0
+ $Y2=0
cc_494 N_A_33_47#_c_549_n N_VGND_c_1028_n 0.00136257f $X=0.287 $Y=0.75 $X2=0
+ $Y2=0
cc_495 N_A_33_47#_c_553_n N_VGND_c_1028_n 7.12888e-19 $X=2.565 $Y=0.935 $X2=0
+ $Y2=0
cc_496 N_A_33_47#_c_542_n A_258_81# 0.00366293f $X=2.36 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_497 N_A_33_47#_c_542_n A_416_81# 0.00670061f $X=2.36 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_498 N_CLK_c_771_n N_A_1039_367#_c_844_n 0.00133887f $X=4.935 $Y=1.552 $X2=0
+ $Y2=0
cc_499 N_CLK_M1006_g N_A_1039_367#_c_838_n 0.00138807f $X=4.935 $Y=0.875 $X2=0
+ $Y2=0
cc_500 N_CLK_c_775_n N_VPWR_c_912_n 0.00312414f $X=4.53 $Y=1.725 $X2=0 $Y2=0
cc_501 N_CLK_c_776_n N_VPWR_c_915_n 0.00312414f $X=5.12 $Y=1.725 $X2=0 $Y2=0
cc_502 N_CLK_c_775_n N_VPWR_c_906_n 0.00410284f $X=4.53 $Y=1.725 $X2=0 $Y2=0
cc_503 N_CLK_c_776_n N_VPWR_c_906_n 0.00410284f $X=5.12 $Y=1.725 $X2=0 $Y2=0
cc_504 N_CLK_M1007_g N_VGND_c_1022_n 6.65218e-19 $X=4.31 $Y=0.875 $X2=0 $Y2=0
cc_505 N_CLK_M1006_g N_VGND_c_1023_n 0.00394852f $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_506 N_CLK_M1006_g N_VGND_c_1028_n 0.00458517f $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_507 N_A_1039_367#_c_843_n N_VPWR_M1016_d 0.00373046f $X=5.945 $Y=1.79 $X2=0
+ $Y2=0
cc_508 N_A_1039_367#_M1010_g N_VPWR_c_909_n 0.02108f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_509 N_A_1039_367#_M1018_g N_VPWR_c_909_n 7.69857e-19 $X=6.675 $Y=2.465 $X2=0
+ $Y2=0
cc_510 N_A_1039_367#_c_842_n N_VPWR_c_909_n 0.00132442f $X=5.385 $Y=1.98 $X2=0
+ $Y2=0
cc_511 N_A_1039_367#_c_843_n N_VPWR_c_909_n 0.0308105f $X=5.945 $Y=1.79 $X2=0
+ $Y2=0
cc_512 N_A_1039_367#_c_839_n N_VPWR_c_909_n 9.997e-19 $X=6.132 $Y=1.42 $X2=0
+ $Y2=0
cc_513 N_A_1039_367#_M1018_g N_VPWR_c_911_n 0.00742417f $X=6.675 $Y=2.465 $X2=0
+ $Y2=0
cc_514 N_A_1039_367#_M1010_g N_VPWR_c_916_n 0.00486043f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_515 N_A_1039_367#_M1018_g N_VPWR_c_916_n 0.00585385f $X=6.675 $Y=2.465 $X2=0
+ $Y2=0
cc_516 N_A_1039_367#_M1010_g N_VPWR_c_906_n 0.00824727f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_517 N_A_1039_367#_M1018_g N_VPWR_c_906_n 0.0115673f $X=6.675 $Y=2.465 $X2=0
+ $Y2=0
cc_518 N_A_1039_367#_c_842_n N_VPWR_c_906_n 0.0131878f $X=5.385 $Y=1.98 $X2=0
+ $Y2=0
cc_519 N_A_1039_367#_M1003_g N_GCLK_c_996_n 0.00248435f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_520 N_A_1039_367#_c_832_n N_GCLK_c_996_n 0.0159431f $X=6.6 $Y=1.42 $X2=0
+ $Y2=0
cc_521 N_A_1039_367#_M1017_g N_GCLK_c_996_n 0.00737032f $X=6.675 $Y=0.655 $X2=0
+ $Y2=0
cc_522 N_A_1039_367#_M1018_g N_GCLK_c_996_n 0.00938361f $X=6.675 $Y=2.465 $X2=0
+ $Y2=0
cc_523 N_A_1039_367#_c_843_n N_GCLK_c_996_n 0.0122469f $X=5.945 $Y=1.79 $X2=0
+ $Y2=0
cc_524 N_A_1039_367#_c_836_n N_GCLK_c_996_n 0.0107811f $X=5.945 $Y=1.09 $X2=0
+ $Y2=0
cc_525 N_A_1039_367#_c_837_n N_GCLK_c_996_n 0.039141f $X=6.11 $Y=1.51 $X2=0
+ $Y2=0
cc_526 N_A_1039_367#_c_839_n N_GCLK_c_996_n 0.0033053f $X=6.132 $Y=1.42 $X2=0
+ $Y2=0
cc_527 N_A_1039_367#_c_836_n N_VGND_M1003_d 0.00259701f $X=5.945 $Y=1.09 $X2=0
+ $Y2=0
cc_528 N_A_1039_367#_M1003_g N_VGND_c_1016_n 0.0113201f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_529 N_A_1039_367#_M1017_g N_VGND_c_1016_n 6.28227e-19 $X=6.675 $Y=0.655 $X2=0
+ $Y2=0
cc_530 N_A_1039_367#_c_836_n N_VGND_c_1016_n 0.0236483f $X=5.945 $Y=1.09 $X2=0
+ $Y2=0
cc_531 N_A_1039_367#_c_838_n N_VGND_c_1016_n 0.0096253f $X=5.51 $Y=0.875 $X2=0
+ $Y2=0
cc_532 N_A_1039_367#_c_839_n N_VGND_c_1016_n 7.7289e-19 $X=6.132 $Y=1.42 $X2=0
+ $Y2=0
cc_533 N_A_1039_367#_M1017_g N_VGND_c_1018_n 0.00707803f $X=6.675 $Y=0.655 $X2=0
+ $Y2=0
cc_534 N_A_1039_367#_c_838_n N_VGND_c_1023_n 0.00480601f $X=5.51 $Y=0.875 $X2=0
+ $Y2=0
cc_535 N_A_1039_367#_M1003_g N_VGND_c_1024_n 0.00486043f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_536 N_A_1039_367#_M1017_g N_VGND_c_1024_n 0.00585385f $X=6.675 $Y=0.655 $X2=0
+ $Y2=0
cc_537 N_A_1039_367#_M1003_g N_VGND_c_1028_n 0.00824727f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_538 N_A_1039_367#_M1017_g N_VGND_c_1028_n 0.011499f $X=6.675 $Y=0.655 $X2=0
+ $Y2=0
cc_539 N_A_1039_367#_c_838_n N_VGND_c_1028_n 0.0092047f $X=5.51 $Y=0.875 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_906_n N_GCLK_M1010_s 0.0041489f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_541 N_VPWR_c_911_n N_GCLK_c_996_n 0.00137338f $X=6.89 $Y=1.98 $X2=0 $Y2=0
cc_542 N_VPWR_c_916_n N_GCLK_c_996_n 0.0136943f $X=6.785 $Y=3.33 $X2=0 $Y2=0
cc_543 N_VPWR_c_906_n N_GCLK_c_996_n 0.00866972f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_544 N_GCLK_c_996_n N_VGND_c_1018_n 0.0015231f $X=6.46 $Y=0.42 $X2=0 $Y2=0
cc_545 N_GCLK_c_996_n N_VGND_c_1024_n 0.0136943f $X=6.46 $Y=0.42 $X2=0 $Y2=0
cc_546 N_GCLK_M1003_s N_VGND_c_1028_n 0.0041489f $X=6.32 $Y=0.235 $X2=0 $Y2=0
cc_547 N_GCLK_c_996_n N_VGND_c_1028_n 0.00866972f $X=6.46 $Y=0.42 $X2=0 $Y2=0
