* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_508_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND a_304_153# a_22_259# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_22_259# A1 a_594_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND B1_N a_304_153# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR B1_N a_304_153# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 X a_22_259# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 X a_22_259# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VPWR a_22_259# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR A2 a_508_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_22_259# a_304_153# a_508_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND a_22_259# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_594_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
