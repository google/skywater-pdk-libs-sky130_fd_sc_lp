* File: sky130_fd_sc_lp__o31a_0.pxi.spice
* Created: Fri Aug 28 11:15:16 2020
* 
x_PM_SKY130_FD_SC_LP__O31A_0%A_90_309# N_A_90_309#_M1007_d N_A_90_309#_M1009_d
+ N_A_90_309#_M1001_g N_A_90_309#_M1008_g N_A_90_309#_c_81_n N_A_90_309#_c_82_n
+ N_A_90_309#_c_76_n N_A_90_309#_c_77_n N_A_90_309#_c_85_n N_A_90_309#_c_86_n
+ N_A_90_309#_c_87_n N_A_90_309#_c_88_n N_A_90_309#_c_78_n N_A_90_309#_c_90_n
+ N_A_90_309#_c_79_n PM_SKY130_FD_SC_LP__O31A_0%A_90_309#
x_PM_SKY130_FD_SC_LP__O31A_0%A1 N_A1_M1000_g N_A1_M1004_g N_A1_c_151_n
+ N_A1_c_152_n A1 A1 A1 N_A1_c_153_n N_A1_c_154_n A1
+ PM_SKY130_FD_SC_LP__O31A_0%A1
x_PM_SKY130_FD_SC_LP__O31A_0%A2 N_A2_M1002_g N_A2_M1005_g N_A2_c_195_n
+ N_A2_c_196_n A2 A2 N_A2_c_198_n PM_SKY130_FD_SC_LP__O31A_0%A2
x_PM_SKY130_FD_SC_LP__O31A_0%A3 N_A3_M1009_g N_A3_M1003_g N_A3_c_239_n A3 A3
+ N_A3_c_241_n PM_SKY130_FD_SC_LP__O31A_0%A3
x_PM_SKY130_FD_SC_LP__O31A_0%B1 N_B1_M1006_g N_B1_M1007_g N_B1_c_289_n
+ N_B1_c_290_n N_B1_c_283_n N_B1_c_284_n N_B1_c_285_n B1 B1 N_B1_c_286_n
+ N_B1_c_287_n PM_SKY130_FD_SC_LP__O31A_0%B1
x_PM_SKY130_FD_SC_LP__O31A_0%X N_X_M1008_s N_X_M1001_s X X X X X X X N_X_c_327_n
+ X PM_SKY130_FD_SC_LP__O31A_0%X
x_PM_SKY130_FD_SC_LP__O31A_0%VPWR N_VPWR_M1001_d N_VPWR_M1006_d N_VPWR_c_346_n
+ N_VPWR_c_347_n N_VPWR_c_348_n N_VPWR_c_349_n VPWR N_VPWR_c_350_n
+ N_VPWR_c_351_n N_VPWR_c_345_n N_VPWR_c_353_n PM_SKY130_FD_SC_LP__O31A_0%VPWR
x_PM_SKY130_FD_SC_LP__O31A_0%VGND N_VGND_M1008_d N_VGND_M1005_d N_VGND_c_377_n
+ N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n VGND N_VGND_c_381_n
+ N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n PM_SKY130_FD_SC_LP__O31A_0%VGND
x_PM_SKY130_FD_SC_LP__O31A_0%A_270_55# N_A_270_55#_M1000_d N_A_270_55#_M1003_d
+ N_A_270_55#_c_417_n N_A_270_55#_c_418_n N_A_270_55#_c_419_n
+ PM_SKY130_FD_SC_LP__O31A_0%A_270_55#
cc_1 VNB N_A_90_309#_M1008_g 0.0643805f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.485
cc_2 VNB N_A_90_309#_c_76_n 0.00736408f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.71
cc_3 VNB N_A_90_309#_c_77_n 0.0156885f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.71
cc_4 VNB N_A_90_309#_c_78_n 0.0491882f $X=-0.19 $Y=-0.245 $X2=3.182 $Y2=2.035
cc_5 VNB N_A_90_309#_c_79_n 0.0208973f $X=-0.19 $Y=-0.245 $X2=3.182 $Y2=0.485
cc_6 VNB N_A1_M1000_g 0.0208315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A1_M1004_g 0.00724415f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.215
cc_8 VNB N_A1_c_151_n 0.0207254f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.545
cc_9 VNB N_A1_c_152_n 0.0155656f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.485
cc_10 VNB N_A1_c_153_n 0.0165343f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.71
cc_11 VNB N_A1_c_154_n 0.00761178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A1 0.00377826f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.125
cc_13 VNB N_A2_M1005_g 0.0317751f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.215
cc_14 VNB N_A2_c_195_n 0.0208556f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.545
cc_15 VNB N_A2_c_196_n 0.00432132f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.485
cc_16 VNB A2 0.0053436f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.485
cc_17 VNB N_A2_c_198_n 0.0156542f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.215
cc_18 VNB N_A3_M1003_g 0.037052f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.215
cc_19 VNB N_A3_c_239_n 0.0185053f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.725
cc_20 VNB A3 0.00530849f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.485
cc_21 VNB N_A3_c_241_n 0.0155242f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.05
cc_22 VNB N_B1_c_283_n 0.020419f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.71
cc_23 VNB N_B1_c_284_n 0.0206773f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.545
cc_24 VNB N_B1_c_285_n 0.00664129f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.215
cc_25 VNB N_B1_c_286_n 0.0437335f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.125
cc_26 VNB N_B1_c_287_n 0.00588385f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.125
cc_27 VNB X 0.0571722f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.725
cc_28 VNB N_X_c_327_n 0.019899f $X=-0.19 $Y=-0.245 $X2=3.182 $Y2=0.485
cc_29 VNB N_VPWR_c_345_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=2.125
cc_30 VNB N_VGND_c_377_n 0.00695557f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.725
cc_31 VNB N_VGND_c_378_n 0.00151893f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.485
cc_32 VNB N_VGND_c_379_n 0.0241749f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.545
cc_33 VNB N_VGND_c_380_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.05
cc_34 VNB N_VGND_c_381_n 0.018137f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.125
cc_35 VNB N_VGND_c_382_n 0.0319043f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=2.125
cc_36 VNB N_VGND_c_383_n 0.204498f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=2.125
cc_37 VNB N_VGND_c_384_n 0.00485433f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=2.125
cc_38 VNB N_A_270_55#_c_417_n 0.0165133f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.215
cc_39 VNB N_A_270_55#_c_418_n 3.69861e-19 $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.545
cc_40 VNB N_A_270_55#_c_419_n 0.00570532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_A_90_309#_M1001_g 0.0261238f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.725
cc_42 VPB N_A_90_309#_c_81_n 0.0258499f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.05
cc_43 VPB N_A_90_309#_c_82_n 0.0175594f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.215
cc_44 VPB N_A_90_309#_c_76_n 0.00345269f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.71
cc_45 VPB N_A_90_309#_c_77_n 0.0042093f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.71
cc_46 VPB N_A_90_309#_c_85_n 0.0397359f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.125
cc_47 VPB N_A_90_309#_c_86_n 0.00456184f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.125
cc_48 VPB N_A_90_309#_c_87_n 0.00428585f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=2.55
cc_49 VPB N_A_90_309#_c_88_n 0.0317992f $X=-0.19 $Y=1.655 $X2=3.09 $Y2=2.125
cc_50 VPB N_A_90_309#_c_78_n 0.0187162f $X=-0.19 $Y=1.655 $X2=3.182 $Y2=2.035
cc_51 VPB N_A_90_309#_c_90_n 0.00213872f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=2.125
cc_52 VPB N_A1_M1004_g 0.0523549f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.215
cc_53 VPB A1 0.00307191f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.125
cc_54 VPB N_A2_M1002_g 0.0417852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A2_c_196_n 0.0109731f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.485
cc_56 VPB A2 0.00331136f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.485
cc_57 VPB N_A3_M1009_g 0.0230588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A3_c_239_n 0.0416112f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.725
cc_59 VPB A3 0.00292035f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.485
cc_60 VPB N_B1_M1006_g 0.0252387f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_B1_c_289_n 0.0229608f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.725
cc_62 VPB N_B1_c_290_n 0.0245882f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.485
cc_63 VPB N_B1_c_285_n 0.0100508f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.215
cc_64 VPB N_B1_c_287_n 0.00442535f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.125
cc_65 VPB X 0.0387255f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.725
cc_66 VPB X 0.0428359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_346_n 0.0107254f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.725
cc_68 VPB N_VPWR_c_347_n 0.0363106f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.485
cc_69 VPB N_VPWR_c_348_n 0.0235343f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.545
cc_70 VPB N_VPWR_c_349_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.05
cc_71 VPB N_VPWR_c_350_n 0.0436832f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.125
cc_72 VPB N_VPWR_c_351_n 0.0153494f $X=-0.19 $Y=1.655 $X2=3.09 $Y2=2.125
cc_73 VPB N_VPWR_c_345_n 0.0888678f $X=-0.19 $Y=1.655 $X2=2.445 $Y2=2.125
cc_74 VPB N_VPWR_c_353_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=2.125
cc_75 N_A_90_309#_M1008_g N_A1_M1000_g 0.0165609f $X=0.705 $Y=0.485 $X2=0 $Y2=0
cc_76 N_A_90_309#_M1001_g N_A1_M1004_g 0.0204319f $X=0.68 $Y=2.725 $X2=0 $Y2=0
cc_77 N_A_90_309#_M1008_g N_A1_M1004_g 0.0177526f $X=0.705 $Y=0.485 $X2=0 $Y2=0
cc_78 N_A_90_309#_c_76_n N_A1_M1004_g 0.00415805f $X=0.615 $Y=1.71 $X2=0 $Y2=0
cc_79 N_A_90_309#_c_85_n N_A1_M1004_g 0.0160127f $X=2.115 $Y=2.125 $X2=0 $Y2=0
cc_80 N_A_90_309#_c_85_n N_A1_c_152_n 5.93261e-19 $X=2.115 $Y=2.125 $X2=0 $Y2=0
cc_81 N_A_90_309#_M1008_g N_A1_c_153_n 0.033731f $X=0.705 $Y=0.485 $X2=0 $Y2=0
cc_82 N_A_90_309#_M1008_g N_A1_c_154_n 0.00420105f $X=0.705 $Y=0.485 $X2=0 $Y2=0
cc_83 N_A_90_309#_M1008_g A1 0.0030027f $X=0.705 $Y=0.485 $X2=0 $Y2=0
cc_84 N_A_90_309#_c_76_n A1 0.0265785f $X=0.615 $Y=1.71 $X2=0 $Y2=0
cc_85 N_A_90_309#_c_77_n A1 0.00106262f $X=0.615 $Y=1.71 $X2=0 $Y2=0
cc_86 N_A_90_309#_c_85_n A1 0.0269963f $X=2.115 $Y=2.125 $X2=0 $Y2=0
cc_87 N_A_90_309#_c_85_n N_A2_M1002_g 0.0148524f $X=2.115 $Y=2.125 $X2=0 $Y2=0
cc_88 N_A_90_309#_c_87_n N_A2_M1002_g 0.00412521f $X=2.28 $Y=2.55 $X2=0 $Y2=0
cc_89 N_A_90_309#_c_85_n N_A2_c_196_n 0.00349567f $X=2.115 $Y=2.125 $X2=0 $Y2=0
cc_90 N_A_90_309#_c_85_n A2 0.0231719f $X=2.115 $Y=2.125 $X2=0 $Y2=0
cc_91 N_A_90_309#_c_85_n N_A3_M1009_g 0.00754116f $X=2.115 $Y=2.125 $X2=0 $Y2=0
cc_92 N_A_90_309#_c_87_n N_A3_M1009_g 0.0163184f $X=2.28 $Y=2.55 $X2=0 $Y2=0
cc_93 N_A_90_309#_c_90_n N_A3_M1009_g 0.00109023f $X=2.28 $Y=2.125 $X2=0 $Y2=0
cc_94 N_A_90_309#_c_85_n N_A3_c_239_n 0.00318276f $X=2.115 $Y=2.125 $X2=0 $Y2=0
cc_95 N_A_90_309#_c_90_n N_A3_c_239_n 0.0123971f $X=2.28 $Y=2.125 $X2=0 $Y2=0
cc_96 N_A_90_309#_c_85_n A3 0.0107356f $X=2.115 $Y=2.125 $X2=0 $Y2=0
cc_97 N_A_90_309#_c_90_n A3 0.0202319f $X=2.28 $Y=2.125 $X2=0 $Y2=0
cc_98 N_A_90_309#_c_88_n N_B1_c_289_n 0.00558978f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_99 N_A_90_309#_c_78_n N_B1_c_289_n 0.00604011f $X=3.182 $Y=2.035 $X2=0 $Y2=0
cc_100 N_A_90_309#_c_87_n N_B1_c_290_n 0.00523965f $X=2.28 $Y=2.55 $X2=0 $Y2=0
cc_101 N_A_90_309#_c_88_n N_B1_c_290_n 0.0188127f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_102 N_A_90_309#_c_78_n N_B1_c_283_n 0.00241777f $X=3.182 $Y=2.035 $X2=0 $Y2=0
cc_103 N_A_90_309#_c_78_n N_B1_c_284_n 0.0259513f $X=3.182 $Y=2.035 $X2=0 $Y2=0
cc_104 N_A_90_309#_c_79_n N_B1_c_284_n 0.0077689f $X=3.182 $Y=0.485 $X2=0 $Y2=0
cc_105 N_A_90_309#_c_88_n N_B1_c_285_n 0.0034004f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_106 N_A_90_309#_c_88_n N_B1_c_287_n 0.0324972f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_107 N_A_90_309#_c_78_n N_B1_c_287_n 0.0627276f $X=3.182 $Y=2.035 $X2=0 $Y2=0
cc_108 N_A_90_309#_c_79_n N_B1_c_287_n 0.00516447f $X=3.182 $Y=0.485 $X2=0 $Y2=0
cc_109 N_A_90_309#_M1001_g X 0.00556974f $X=0.68 $Y=2.725 $X2=0 $Y2=0
cc_110 N_A_90_309#_M1008_g X 0.0205467f $X=0.705 $Y=0.485 $X2=0 $Y2=0
cc_111 N_A_90_309#_c_76_n X 0.0363088f $X=0.615 $Y=1.71 $X2=0 $Y2=0
cc_112 N_A_90_309#_c_77_n X 0.0165543f $X=0.615 $Y=1.71 $X2=0 $Y2=0
cc_113 N_A_90_309#_c_86_n X 0.0141862f $X=0.845 $Y=2.125 $X2=0 $Y2=0
cc_114 N_A_90_309#_M1001_g X 0.00122519f $X=0.68 $Y=2.725 $X2=0 $Y2=0
cc_115 N_A_90_309#_c_82_n X 0.00412481f $X=0.615 $Y=2.215 $X2=0 $Y2=0
cc_116 N_A_90_309#_c_86_n X 0.00347742f $X=0.845 $Y=2.125 $X2=0 $Y2=0
cc_117 N_A_90_309#_M1001_g N_VPWR_c_346_n 0.00972211f $X=0.68 $Y=2.725 $X2=0
+ $Y2=0
cc_118 N_A_90_309#_c_85_n N_VPWR_c_346_n 0.0253142f $X=2.115 $Y=2.125 $X2=0
+ $Y2=0
cc_119 N_A_90_309#_c_86_n N_VPWR_c_346_n 0.00266746f $X=0.845 $Y=2.125 $X2=0
+ $Y2=0
cc_120 N_A_90_309#_c_87_n N_VPWR_c_347_n 0.00232983f $X=2.28 $Y=2.55 $X2=0 $Y2=0
cc_121 N_A_90_309#_c_88_n N_VPWR_c_347_n 0.0270339f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_122 N_A_90_309#_M1001_g N_VPWR_c_348_n 0.0053602f $X=0.68 $Y=2.725 $X2=0
+ $Y2=0
cc_123 N_A_90_309#_c_87_n N_VPWR_c_350_n 0.0208231f $X=2.28 $Y=2.55 $X2=0 $Y2=0
cc_124 N_A_90_309#_M1001_g N_VPWR_c_345_n 0.0113243f $X=0.68 $Y=2.725 $X2=0
+ $Y2=0
cc_125 N_A_90_309#_c_87_n N_VPWR_c_345_n 0.012564f $X=2.28 $Y=2.55 $X2=0 $Y2=0
cc_126 N_A_90_309#_M1008_g N_VGND_c_377_n 0.00550347f $X=0.705 $Y=0.485 $X2=0
+ $Y2=0
cc_127 N_A_90_309#_M1008_g N_VGND_c_379_n 0.00545548f $X=0.705 $Y=0.485 $X2=0
+ $Y2=0
cc_128 N_A_90_309#_c_79_n N_VGND_c_382_n 0.0227914f $X=3.182 $Y=0.485 $X2=0
+ $Y2=0
cc_129 N_A_90_309#_M1008_g N_VGND_c_383_n 0.0114801f $X=0.705 $Y=0.485 $X2=0
+ $Y2=0
cc_130 N_A_90_309#_c_79_n N_VGND_c_383_n 0.018372f $X=3.182 $Y=0.485 $X2=0 $Y2=0
cc_131 N_A_90_309#_c_78_n N_A_270_55#_c_417_n 0.0069197f $X=3.182 $Y=2.035 $X2=0
+ $Y2=0
cc_132 N_A_90_309#_c_78_n N_A_270_55#_c_418_n 0.0015417f $X=3.182 $Y=2.035 $X2=0
+ $Y2=0
cc_133 N_A1_M1004_g N_A2_M1002_g 0.0696047f $X=1.275 $Y=2.725 $X2=0 $Y2=0
cc_134 N_A1_M1000_g N_A2_M1005_g 0.018134f $X=1.275 $Y=0.485 $X2=0 $Y2=0
cc_135 N_A1_c_154_n N_A2_M1005_g 0.00109318f $X=1.182 $Y=1.247 $X2=0 $Y2=0
cc_136 N_A1_c_152_n N_A2_c_195_n 0.0137825f $X=1.185 $Y=1.51 $X2=0 $Y2=0
cc_137 A1 N_A2_c_195_n 5.77951e-19 $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_138 N_A1_M1004_g N_A2_c_196_n 0.0137825f $X=1.275 $Y=2.725 $X2=0 $Y2=0
cc_139 N_A1_c_151_n A2 0.00386238f $X=1.185 $Y=1.345 $X2=0 $Y2=0
cc_140 N_A1_c_154_n A2 0.0131602f $X=1.182 $Y=1.247 $X2=0 $Y2=0
cc_141 A1 A2 0.0483507f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_142 N_A1_c_151_n N_A2_c_198_n 0.0137825f $X=1.185 $Y=1.345 $X2=0 $Y2=0
cc_143 N_A1_c_154_n X 0.013264f $X=1.182 $Y=1.247 $X2=0 $Y2=0
cc_144 A1 X 0.00930291f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_145 N_A1_M1004_g N_VPWR_c_346_n 0.00781315f $X=1.275 $Y=2.725 $X2=0 $Y2=0
cc_146 N_A1_M1004_g N_VPWR_c_350_n 0.0053602f $X=1.275 $Y=2.725 $X2=0 $Y2=0
cc_147 N_A1_M1004_g N_VPWR_c_345_n 0.0105654f $X=1.275 $Y=2.725 $X2=0 $Y2=0
cc_148 N_A1_M1000_g N_VGND_c_377_n 0.00550347f $X=1.275 $Y=0.485 $X2=0 $Y2=0
cc_149 N_A1_c_153_n N_VGND_c_377_n 9.60108e-19 $X=1.185 $Y=1.005 $X2=0 $Y2=0
cc_150 N_A1_c_154_n N_VGND_c_377_n 0.0119434f $X=1.182 $Y=1.247 $X2=0 $Y2=0
cc_151 N_A1_M1000_g N_VGND_c_378_n 9.87958e-19 $X=1.275 $Y=0.485 $X2=0 $Y2=0
cc_152 N_A1_M1000_g N_VGND_c_381_n 0.00545548f $X=1.275 $Y=0.485 $X2=0 $Y2=0
cc_153 N_A1_M1000_g N_VGND_c_383_n 0.00795079f $X=1.275 $Y=0.485 $X2=0 $Y2=0
cc_154 N_A1_c_154_n N_VGND_c_383_n 0.00544454f $X=1.182 $Y=1.247 $X2=0 $Y2=0
cc_155 N_A1_M1000_g N_A_270_55#_c_419_n 0.00517971f $X=1.275 $Y=0.485 $X2=0
+ $Y2=0
cc_156 N_A1_c_154_n N_A_270_55#_c_419_n 0.00541015f $X=1.182 $Y=1.247 $X2=0
+ $Y2=0
cc_157 N_A2_M1005_g N_A3_M1003_g 0.0228814f $X=1.785 $Y=0.485 $X2=0 $Y2=0
cc_158 A2 N_A3_M1003_g 6.06643e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A2_c_198_n N_A3_M1003_g 0.00491066f $X=1.725 $Y=1.245 $X2=0 $Y2=0
cc_160 N_A2_M1002_g N_A3_c_239_n 0.0841119f $X=1.695 $Y=2.725 $X2=0 $Y2=0
cc_161 N_A2_c_195_n N_A3_c_239_n 0.017115f $X=1.725 $Y=1.585 $X2=0 $Y2=0
cc_162 A2 N_A3_c_239_n 3.08978e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A2_M1002_g A3 3.89002e-19 $X=1.695 $Y=2.725 $X2=0 $Y2=0
cc_164 A2 A3 0.0534035f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A2_c_198_n A3 0.00371512f $X=1.725 $Y=1.245 $X2=0 $Y2=0
cc_166 A2 N_A3_c_241_n 4.83776e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_167 N_A2_c_198_n N_A3_c_241_n 0.017115f $X=1.725 $Y=1.245 $X2=0 $Y2=0
cc_168 N_A2_M1002_g N_VPWR_c_350_n 0.0053602f $X=1.695 $Y=2.725 $X2=0 $Y2=0
cc_169 N_A2_M1002_g N_VPWR_c_345_n 0.0103205f $X=1.695 $Y=2.725 $X2=0 $Y2=0
cc_170 N_A2_M1005_g N_VGND_c_378_n 0.00701578f $X=1.785 $Y=0.485 $X2=0 $Y2=0
cc_171 N_A2_M1005_g N_VGND_c_381_n 0.0038905f $X=1.785 $Y=0.485 $X2=0 $Y2=0
cc_172 N_A2_M1005_g N_VGND_c_383_n 0.00491812f $X=1.785 $Y=0.485 $X2=0 $Y2=0
cc_173 N_A2_M1005_g N_A_270_55#_c_417_n 0.0135642f $X=1.785 $Y=0.485 $X2=0 $Y2=0
cc_174 A2 N_A_270_55#_c_417_n 0.00851851f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A2_c_198_n N_A_270_55#_c_417_n 0.00136716f $X=1.725 $Y=1.245 $X2=0
+ $Y2=0
cc_176 N_A2_M1005_g N_A_270_55#_c_419_n 3.84036e-19 $X=1.785 $Y=0.485 $X2=0
+ $Y2=0
cc_177 A2 N_A_270_55#_c_419_n 0.0131665f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A2_c_198_n N_A_270_55#_c_419_n 9.39773e-19 $X=1.725 $Y=1.245 $X2=0
+ $Y2=0
cc_179 N_A3_c_239_n N_B1_c_289_n 0.00784798f $X=2.265 $Y=1.7 $X2=0 $Y2=0
cc_180 N_A3_M1009_g N_B1_c_290_n 0.0141021f $X=2.055 $Y=2.725 $X2=0 $Y2=0
cc_181 N_A3_c_239_n N_B1_c_290_n 0.0022697f $X=2.265 $Y=1.7 $X2=0 $Y2=0
cc_182 N_A3_M1003_g N_B1_c_283_n 0.0191335f $X=2.255 $Y=0.485 $X2=0 $Y2=0
cc_183 N_A3_c_239_n N_B1_c_285_n 0.0173878f $X=2.265 $Y=1.7 $X2=0 $Y2=0
cc_184 N_A3_M1003_g N_B1_c_286_n 0.00888797f $X=2.255 $Y=0.485 $X2=0 $Y2=0
cc_185 A3 N_B1_c_286_n 5.70358e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A3_c_241_n N_B1_c_286_n 0.0173878f $X=2.265 $Y=1.36 $X2=0 $Y2=0
cc_187 N_A3_M1003_g N_B1_c_287_n 0.00342259f $X=2.255 $Y=0.485 $X2=0 $Y2=0
cc_188 A3 N_B1_c_287_n 0.0542081f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A3_c_241_n N_B1_c_287_n 0.00483511f $X=2.265 $Y=1.36 $X2=0 $Y2=0
cc_190 N_A3_M1009_g N_VPWR_c_350_n 0.00516731f $X=2.055 $Y=2.725 $X2=0 $Y2=0
cc_191 N_A3_M1009_g N_VPWR_c_345_n 0.00989939f $X=2.055 $Y=2.725 $X2=0 $Y2=0
cc_192 N_A3_M1003_g N_VGND_c_378_n 0.00689355f $X=2.255 $Y=0.485 $X2=0 $Y2=0
cc_193 N_A3_M1003_g N_VGND_c_382_n 0.0038905f $X=2.255 $Y=0.485 $X2=0 $Y2=0
cc_194 N_A3_M1003_g N_VGND_c_383_n 0.004779f $X=2.255 $Y=0.485 $X2=0 $Y2=0
cc_195 N_A3_M1003_g N_A_270_55#_c_417_n 0.0125961f $X=2.255 $Y=0.485 $X2=0 $Y2=0
cc_196 A3 N_A_270_55#_c_417_n 0.0186789f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A3_c_241_n N_A_270_55#_c_417_n 0.00382239f $X=2.265 $Y=1.36 $X2=0 $Y2=0
cc_198 N_A3_M1003_g N_A_270_55#_c_418_n 3.40397e-19 $X=2.255 $Y=0.485 $X2=0
+ $Y2=0
cc_199 N_B1_M1006_g N_VPWR_c_347_n 0.00544417f $X=2.535 $Y=2.725 $X2=0 $Y2=0
cc_200 N_B1_c_290_n N_VPWR_c_347_n 0.00541747f $X=2.745 $Y=2.18 $X2=0 $Y2=0
cc_201 N_B1_M1006_g N_VPWR_c_350_n 0.0053602f $X=2.535 $Y=2.725 $X2=0 $Y2=0
cc_202 N_B1_M1006_g N_VPWR_c_345_n 0.0111686f $X=2.535 $Y=2.725 $X2=0 $Y2=0
cc_203 N_B1_c_283_n N_VGND_c_378_n 0.00109223f $X=2.805 $Y=0.805 $X2=0 $Y2=0
cc_204 N_B1_c_283_n N_VGND_c_382_n 0.00545548f $X=2.805 $Y=0.805 $X2=0 $Y2=0
cc_205 N_B1_c_283_n N_VGND_c_383_n 0.0113854f $X=2.805 $Y=0.805 $X2=0 $Y2=0
cc_206 N_B1_c_284_n N_VGND_c_383_n 3.91649e-19 $X=2.805 $Y=0.955 $X2=0 $Y2=0
cc_207 N_B1_c_283_n N_A_270_55#_c_417_n 0.00268795f $X=2.805 $Y=0.805 $X2=0
+ $Y2=0
cc_208 N_B1_c_287_n N_A_270_55#_c_417_n 0.00776378f $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_209 N_B1_c_283_n N_A_270_55#_c_418_n 3.1341e-19 $X=2.805 $Y=0.805 $X2=0 $Y2=0
cc_210 X N_VPWR_c_346_n 0.0228483f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_211 X N_VPWR_c_348_n 0.0346421f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_212 X N_VPWR_c_345_n 0.0187812f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_213 N_X_c_327_n N_VGND_c_379_n 0.0237149f $X=0.49 $Y=0.485 $X2=0 $Y2=0
cc_214 N_X_c_327_n N_VGND_c_383_n 0.0187395f $X=0.49 $Y=0.485 $X2=0 $Y2=0
cc_215 N_VGND_c_378_n N_A_270_55#_c_417_n 0.0208016f $X=2.02 $Y=0.44 $X2=0 $Y2=0
cc_216 N_VGND_c_381_n N_A_270_55#_c_417_n 0.00235166f $X=1.855 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_382_n N_A_270_55#_c_417_n 0.00235166f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_383_n N_A_270_55#_c_417_n 0.00900713f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_382_n N_A_270_55#_c_418_n 0.0102172f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_383_n N_A_270_55#_c_418_n 0.00926695f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_c_381_n N_A_270_55#_c_419_n 0.0138134f $X=1.855 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_383_n N_A_270_55#_c_419_n 0.011898f $X=3.12 $Y=0 $X2=0 $Y2=0
