* File: sky130_fd_sc_lp__or4bb_4.spice
* Created: Wed Sep  2 10:33:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4bb_4.pex.spice"
.subckt sky130_fd_sc_lp__or4bb_4  VNB VPB C_N A B D_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D_N	D_N
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_C_N_M1011_g N_A_79_137#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0917 AS=0.1113 PD=0.82 PS=1.37 NRD=2.856 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1001 N_A_270_53#_M1001_d N_A_M1001_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1428 AS=0.1834 PD=1.18 PS=1.64 NRD=5.352 NRS=7.14 M=1 R=5.6 SA=75000.5
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_B_M1015_g N_A_270_53#_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1554 AS=0.1428 PD=1.21 PS=1.18 NRD=7.14 NRS=3.204 M=1 R=5.6 SA=75000.9
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1007 N_A_270_53#_M1007_d N_A_79_137#_M1007_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1554 PD=1.12 PS=1.21 NRD=0 NRS=5.712 M=1 R=5.6
+ SA=75001.5 SB=75003.1 A=0.126 P=1.98 MULT=1
MM1018 N_VGND_M1018_d N_A_528_27#_M1018_g N_A_270_53#_M1007_d VNB NSHORT L=0.15
+ W=0.84 AD=0.24695 AS=0.1176 PD=1.5 PS=1.12 NRD=17.136 NRS=0 M=1 R=5.6
+ SA=75001.9 SB=75002.7 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1018_d N_A_270_53#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.24695 AS=0.1176 PD=1.5 PS=1.12 NRD=22.848 NRS=0 M=1 R=5.6 SA=75002.6
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A_270_53#_M1006_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.18425 AS=0.1176 PD=1.37 PS=1.12 NRD=9.276 NRS=0 M=1 R=5.6 SA=75003
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1006_d N_A_270_53#_M1016_g N_X_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.18425 AS=0.1176 PD=1.37 PS=1.12 NRD=9.276 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1017_d N_A_270_53#_M1017_g N_X_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.276067 AS=0.1176 PD=1.94667 PS=1.12 NRD=17.136 NRS=0 M=1 R=5.6 SA=75004
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1012 N_A_528_27#_M1012_d N_D_N_M1012_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.138033 PD=1.37 PS=0.973333 NRD=0 NRS=34.284 M=1 R=2.8
+ SA=75004.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_C_N_M1014_g N_A_79_137#_M1014_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0966 AS=0.1113 PD=0.825 PS=1.37 NRD=82.0702 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 A_270_367# N_A_M1004_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=1.26 AD=0.189
+ AS=0.2898 PD=1.56 PS=2.475 NRD=14.8341 NRS=0 M=1 R=8.4 SA=75000.4 SB=75001.6
+ A=0.189 P=2.82 MULT=1
MM1009 A_360_367# N_B_M1009_g A_270_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.189
+ AS=0.189 PD=1.56 PS=1.56 NRD=14.8341 NRS=14.8341 M=1 R=8.4 SA=75000.8
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1013 A_450_367# N_A_79_137#_M1013_g A_360_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.189 PD=1.65 PS=1.56 NRD=21.8867 NRS=14.8341 M=1 R=8.4
+ SA=75001.3 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1002 N_A_270_53#_M1002_d N_A_528_27#_M1002_g A_450_367# VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4
+ SA=75001.8 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A_270_53#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_270_53#_M1005_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1005_d N_A_270_53#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1019_d N_A_270_53#_M1019_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.4 A=0.189 P=2.82 MULT=1
MM1008 N_A_528_27#_M1008_d N_D_N_M1008_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.095025 PD=1.37 PS=0.8175 NRD=0 NRS=46.886 M=1 R=2.8
+ SA=75002 SB=75000.2 A=0.063 P=1.14 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3463 P=16.97
*
.include "sky130_fd_sc_lp__or4bb_4.pxi.spice"
*
.ends
*
*
