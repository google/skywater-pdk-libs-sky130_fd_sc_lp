* NGSPICE file created from sky130_fd_sc_lp__a31o_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a31o_m A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 VPWR a_86_172# X VPB phighvt w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=1.113e+11p ps=1.37e+06u
M1001 a_86_172# A1 a_354_66# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1002 VPWR A2 a_274_512# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1003 a_282_66# A3 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.583e+11p ps=2.91e+06u
M1004 a_354_66# A2 a_282_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_86_172# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 VGND B1 a_86_172# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_86_172# B1 a_274_512# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 a_274_512# A3 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_274_512# A1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

