* File: sky130_fd_sc_lp__a221oi_lp.pxi.spice
* Created: Wed Sep  2 09:22:08 2020
* 
x_PM_SKY130_FD_SC_LP__A221OI_LP%B2 N_B2_M1010_g N_B2_M1008_g N_B2_c_68_n
+ N_B2_c_69_n B2 B2 N_B2_c_71_n PM_SKY130_FD_SC_LP__A221OI_LP%B2
x_PM_SKY130_FD_SC_LP__A221OI_LP%B1 N_B1_M1009_g N_B1_M1007_g N_B1_c_104_n
+ N_B1_c_105_n N_B1_c_106_n B1 B1 B1 N_B1_c_108_n
+ PM_SKY130_FD_SC_LP__A221OI_LP%B1
x_PM_SKY130_FD_SC_LP__A221OI_LP%A1 N_A1_M1005_g N_A1_M1001_g A1 N_A1_c_168_n
+ PM_SKY130_FD_SC_LP__A221OI_LP%A1
x_PM_SKY130_FD_SC_LP__A221OI_LP%A2 N_A2_c_209_n N_A2_M1002_g N_A2_M1000_g
+ N_A2_c_211_n A2 A2 N_A2_c_213_n PM_SKY130_FD_SC_LP__A221OI_LP%A2
x_PM_SKY130_FD_SC_LP__A221OI_LP%C1 N_C1_M1006_g N_C1_M1004_g N_C1_M1003_g
+ N_C1_c_254_n N_C1_c_255_n C1 C1 N_C1_c_257_n PM_SKY130_FD_SC_LP__A221OI_LP%C1
x_PM_SKY130_FD_SC_LP__A221OI_LP%A_56_412# N_A_56_412#_M1010_s
+ N_A_56_412#_M1007_d N_A_56_412#_c_296_n N_A_56_412#_c_297_n
+ N_A_56_412#_c_303_n N_A_56_412#_c_298_n
+ PM_SKY130_FD_SC_LP__A221OI_LP%A_56_412#
x_PM_SKY130_FD_SC_LP__A221OI_LP%A_163_412# N_A_163_412#_M1010_d
+ N_A_163_412#_M1002_d N_A_163_412#_c_333_n N_A_163_412#_c_337_n
+ N_A_163_412#_c_336_n N_A_163_412#_c_334_n
+ PM_SKY130_FD_SC_LP__A221OI_LP%A_163_412#
x_PM_SKY130_FD_SC_LP__A221OI_LP%VPWR N_VPWR_M1005_d N_VPWR_c_364_n
+ N_VPWR_c_365_n N_VPWR_c_366_n VPWR N_VPWR_c_367_n N_VPWR_c_363_n
+ PM_SKY130_FD_SC_LP__A221OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A221OI_LP%Y N_Y_M1009_d N_Y_M1003_d N_Y_M1004_d
+ N_Y_c_407_n N_Y_c_400_n N_Y_c_404_n N_Y_c_405_n N_Y_c_401_n Y Y N_Y_c_402_n
+ N_Y_c_403_n PM_SKY130_FD_SC_LP__A221OI_LP%Y
x_PM_SKY130_FD_SC_LP__A221OI_LP%VGND N_VGND_M1008_s N_VGND_M1000_d
+ N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n VGND
+ N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n
+ PM_SKY130_FD_SC_LP__A221OI_LP%VGND
cc_1 VNB N_B2_M1008_g 0.04805f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.45
cc_2 VNB N_B2_c_68_n 0.020707f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.26
cc_3 VNB N_B2_c_69_n 0.00428462f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.78
cc_4 VNB B2 0.0463736f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_B2_c_71_n 0.0321522f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.275
cc_6 VNB N_B1_M1009_g 0.0301514f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.56
cc_7 VNB N_B1_c_104_n 0.00936181f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.26
cc_8 VNB N_B1_c_105_n 0.0329278f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.63
cc_9 VNB N_B1_c_106_n 0.00227887f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB B1 0.00933509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_c_108_n 0.0133316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_M1001_g 0.058862f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.45
cc_13 VNB A1 0.00261592f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.26
cc_14 VNB N_A1_c_168_n 0.0172805f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_A2_c_209_n 0.00671617f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.78
cc_16 VNB N_A2_M1000_g 0.0314777f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.45
cc_17 VNB N_A2_c_211_n 0.0183849f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.26
cc_18 VNB A2 0.0193677f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.63
cc_19 VNB N_A2_c_213_n 0.0308198f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_C1_M1006_g 0.0369418f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.56
cc_21 VNB N_C1_M1003_g 0.0370668f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.26
cc_22 VNB N_C1_c_254_n 0.0269099f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_23 VNB N_C1_c_255_n 0.00314574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB C1 3.45983e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C1_c_257_n 0.0349901f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.445
cc_26 VNB N_VPWR_c_363_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.275
cc_27 VNB N_Y_c_400_n 0.00504209f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_28 VNB N_Y_c_401_n 0.0412667f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.275
cc_29 VNB N_Y_c_402_n 0.0171207f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.445
cc_30 VNB N_Y_c_403_n 0.0383677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_453_n 0.0229342f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.26
cc_32 VNB N_VGND_c_454_n 0.00299757f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.63
cc_33 VNB N_VGND_c_455_n 0.0123263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_456_n 0.00517222f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_35 VNB N_VGND_c_457_n 0.0379483f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.275
cc_36 VNB N_VGND_c_458_n 0.0388249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_459_n 0.219373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_460_n 0.00513949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_B2_M1010_g 0.044347f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.56
cc_40 VPB N_B2_c_69_n 0.0156398f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.78
cc_41 VPB B2 0.0133884f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_42 VPB N_B1_M1007_g 0.0260322f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.45
cc_43 VPB N_B1_c_106_n 0.00162785f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_44 VPB B1 0.00636365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_B1_c_108_n 0.0159943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A1_M1005_g 0.028318f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.56
cc_47 VPB A1 7.38393e-19 $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.26
cc_48 VPB N_A1_c_168_n 0.0345081f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_49 VPB N_A2_c_209_n 0.00187595f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.78
cc_50 VPB N_A2_M1002_g 0.0383918f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.56
cc_51 VPB N_C1_M1004_g 0.0383593f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.45
cc_52 VPB N_C1_c_255_n 0.0120565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB C1 8.77644e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_56_412#_c_296_n 0.0113575f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.45
cc_55 VPB N_A_56_412#_c_297_n 0.0331804f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.26
cc_56 VPB N_A_56_412#_c_298_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_163_412#_c_333_n 0.00207208f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.45
cc_58 VPB N_A_163_412#_c_334_n 0.00207208f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.63
cc_59 VPB N_VPWR_c_364_n 0.00385686f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.45
cc_60 VPB N_VPWR_c_365_n 0.0365356f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.26
cc_61 VPB N_VPWR_c_366_n 0.00537149f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.11
cc_62 VPB N_VPWR_c_367_n 0.0592382f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.275
cc_63 VPB N_VPWR_c_363_n 0.0671335f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.275
cc_64 VPB N_Y_c_404_n 0.0396141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_Y_c_405_n 0.02353f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.275
cc_66 VPB N_Y_c_401_n 0.0193114f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.275
cc_67 N_B2_M1008_g N_B1_M1009_g 0.03079f $X=0.7 $Y=0.45 $X2=0 $Y2=0
cc_68 N_B2_M1008_g N_B1_c_104_n 7.04063e-19 $X=0.7 $Y=0.45 $X2=0 $Y2=0
cc_69 B2 N_B1_c_104_n 0.0187499f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_B2_c_68_n N_B1_c_105_n 0.03079f $X=0.58 $Y=1.26 $X2=0 $Y2=0
cc_71 B2 N_B1_c_105_n 8.6896e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_B2_c_71_n N_B1_c_105_n 0.00289389f $X=0.55 $Y=1.275 $X2=0 $Y2=0
cc_73 N_B2_M1010_g N_A1_M1005_g 0.0438884f $X=0.69 $Y=2.56 $X2=0 $Y2=0
cc_74 N_B2_c_69_n A1 0.00100215f $X=0.6 $Y=1.78 $X2=0 $Y2=0
cc_75 B2 A1 0.0160664f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B2_c_69_n N_A1_c_168_n 0.0157367f $X=0.6 $Y=1.78 $X2=0 $Y2=0
cc_77 B2 N_A1_c_168_n 0.00158274f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_78 N_B2_c_71_n N_A1_c_168_n 0.00208594f $X=0.55 $Y=1.275 $X2=0 $Y2=0
cc_79 N_B2_M1010_g N_A_56_412#_c_296_n 0.00204008f $X=0.69 $Y=2.56 $X2=0 $Y2=0
cc_80 N_B2_c_69_n N_A_56_412#_c_296_n 0.00457009f $X=0.6 $Y=1.78 $X2=0 $Y2=0
cc_81 B2 N_A_56_412#_c_296_n 0.0217593f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_82 N_B2_M1010_g N_A_56_412#_c_297_n 0.0144532f $X=0.69 $Y=2.56 $X2=0 $Y2=0
cc_83 N_B2_M1010_g N_A_56_412#_c_303_n 0.0188427f $X=0.69 $Y=2.56 $X2=0 $Y2=0
cc_84 B2 N_A_56_412#_c_303_n 0.0114186f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_B2_M1010_g N_A_163_412#_c_333_n 0.00975364f $X=0.69 $Y=2.56 $X2=0 $Y2=0
cc_86 N_B2_M1010_g N_A_163_412#_c_336_n 0.00484817f $X=0.69 $Y=2.56 $X2=0 $Y2=0
cc_87 N_B2_M1010_g N_VPWR_c_364_n 8.79243e-19 $X=0.69 $Y=2.56 $X2=0 $Y2=0
cc_88 N_B2_M1010_g N_VPWR_c_365_n 0.00848972f $X=0.69 $Y=2.56 $X2=0 $Y2=0
cc_89 N_B2_M1010_g N_VPWR_c_363_n 0.0158996f $X=0.69 $Y=2.56 $X2=0 $Y2=0
cc_90 N_B2_M1008_g N_VGND_c_453_n 0.0155213f $X=0.7 $Y=0.45 $X2=0 $Y2=0
cc_91 N_B2_c_68_n N_VGND_c_453_n 0.00540422f $X=0.58 $Y=1.26 $X2=0 $Y2=0
cc_92 B2 N_VGND_c_453_n 0.0147104f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_93 N_B2_M1008_g N_VGND_c_457_n 0.0048178f $X=0.7 $Y=0.45 $X2=0 $Y2=0
cc_94 N_B2_M1008_g N_VGND_c_459_n 0.00825139f $X=0.7 $Y=0.45 $X2=0 $Y2=0
cc_95 N_B1_M1009_g N_A1_M1001_g 0.0205716f $X=1.09 $Y=0.45 $X2=0 $Y2=0
cc_96 N_B1_c_104_n N_A1_M1001_g 0.0111587f $X=1.565 $Y=1.165 $X2=0 $Y2=0
cc_97 N_B1_c_105_n N_A1_M1001_g 0.021337f $X=1.18 $Y=1.165 $X2=0 $Y2=0
cc_98 N_B1_c_106_n N_A1_M1001_g 0.0123073f $X=1.65 $Y=1.57 $X2=0 $Y2=0
cc_99 N_B1_c_104_n A1 0.0217603f $X=1.565 $Y=1.165 $X2=0 $Y2=0
cc_100 N_B1_c_105_n A1 0.00184024f $X=1.18 $Y=1.165 $X2=0 $Y2=0
cc_101 N_B1_c_106_n A1 0.0265696f $X=1.65 $Y=1.57 $X2=0 $Y2=0
cc_102 N_B1_c_104_n N_A1_c_168_n 0.00702782f $X=1.565 $Y=1.165 $X2=0 $Y2=0
cc_103 N_B1_c_105_n N_A1_c_168_n 0.0158398f $X=1.18 $Y=1.165 $X2=0 $Y2=0
cc_104 N_B1_c_106_n N_A1_c_168_n 0.012315f $X=1.65 $Y=1.57 $X2=0 $Y2=0
cc_105 B1 N_A2_c_209_n 0.00883257f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_106 N_B1_c_108_n N_A2_c_209_n 0.0213656f $X=2.54 $Y=1.735 $X2=-0.19
+ $Y2=-0.245
cc_107 N_B1_M1007_g N_A2_M1002_g 0.0441653f $X=2.57 $Y=2.56 $X2=0 $Y2=0
cc_108 B1 N_A2_M1002_g 0.0120723f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_109 N_B1_c_106_n N_A2_c_211_n 0.0034747f $X=1.65 $Y=1.57 $X2=0 $Y2=0
cc_110 N_B1_c_104_n A2 0.0251137f $X=1.565 $Y=1.165 $X2=0 $Y2=0
cc_111 N_B1_c_106_n A2 0.00425947f $X=1.65 $Y=1.57 $X2=0 $Y2=0
cc_112 B1 A2 0.0626861f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_113 N_B1_c_108_n A2 0.00848307f $X=2.54 $Y=1.735 $X2=0 $Y2=0
cc_114 N_B1_c_104_n N_A2_c_213_n 0.00135657f $X=1.565 $Y=1.165 $X2=0 $Y2=0
cc_115 B1 N_A2_c_213_n 7.70312e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_116 N_B1_M1007_g N_C1_M1004_g 0.0273452f $X=2.57 $Y=2.56 $X2=0 $Y2=0
cc_117 B1 N_C1_M1004_g 0.00311796f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_118 N_B1_c_108_n N_C1_M1004_g 0.00535983f $X=2.54 $Y=1.735 $X2=0 $Y2=0
cc_119 B1 C1 0.0161775f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_120 N_B1_c_108_n C1 2.40913e-19 $X=2.54 $Y=1.735 $X2=0 $Y2=0
cc_121 B1 N_C1_c_257_n 0.00137574f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_122 N_B1_c_108_n N_C1_c_257_n 0.0110891f $X=2.54 $Y=1.735 $X2=0 $Y2=0
cc_123 N_B1_M1007_g N_A_56_412#_c_303_n 0.0178302f $X=2.57 $Y=2.56 $X2=0 $Y2=0
cc_124 N_B1_c_106_n N_A_56_412#_c_303_n 0.0129169f $X=1.65 $Y=1.57 $X2=0 $Y2=0
cc_125 B1 N_A_56_412#_c_303_n 0.0604931f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_126 N_B1_c_108_n N_A_56_412#_c_303_n 0.00143014f $X=2.54 $Y=1.735 $X2=0 $Y2=0
cc_127 N_B1_M1007_g N_A_56_412#_c_298_n 0.0183374f $X=2.57 $Y=2.56 $X2=0 $Y2=0
cc_128 B1 N_A_56_412#_c_298_n 0.00436189f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_129 N_B1_M1007_g N_A_163_412#_c_337_n 0.00471531f $X=2.57 $Y=2.56 $X2=0 $Y2=0
cc_130 N_B1_M1007_g N_A_163_412#_c_334_n 0.00940176f $X=2.57 $Y=2.56 $X2=0 $Y2=0
cc_131 N_B1_M1007_g N_VPWR_c_367_n 0.00848972f $X=2.57 $Y=2.56 $X2=0 $Y2=0
cc_132 N_B1_M1007_g N_VPWR_c_363_n 0.015071f $X=2.57 $Y=2.56 $X2=0 $Y2=0
cc_133 N_B1_M1009_g N_Y_c_407_n 0.00546004f $X=1.09 $Y=0.45 $X2=0 $Y2=0
cc_134 N_B1_M1009_g N_Y_c_400_n 0.00493377f $X=1.09 $Y=0.45 $X2=0 $Y2=0
cc_135 N_B1_c_104_n N_Y_c_400_n 0.0270125f $X=1.565 $Y=1.165 $X2=0 $Y2=0
cc_136 N_B1_c_105_n N_Y_c_400_n 0.00218511f $X=1.18 $Y=1.165 $X2=0 $Y2=0
cc_137 N_B1_M1007_g N_Y_c_405_n 4.71925e-19 $X=2.57 $Y=2.56 $X2=0 $Y2=0
cc_138 N_B1_c_104_n N_Y_c_402_n 0.0114935f $X=1.565 $Y=1.165 $X2=0 $Y2=0
cc_139 N_B1_M1009_g N_VGND_c_453_n 0.00243235f $X=1.09 $Y=0.45 $X2=0 $Y2=0
cc_140 N_B1_M1009_g N_VGND_c_457_n 0.0058025f $X=1.09 $Y=0.45 $X2=0 $Y2=0
cc_141 N_B1_M1009_g N_VGND_c_459_n 0.0111254f $X=1.09 $Y=0.45 $X2=0 $Y2=0
cc_142 N_A1_c_168_n N_A2_c_209_n 0.0214311f $X=1.63 $Y=1.735 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A1_M1005_g N_A2_M1002_g 0.0236254f $X=1.22 $Y=2.56 $X2=0 $Y2=0
cc_144 N_A1_M1001_g N_A2_M1000_g 0.0665213f $X=1.63 $Y=0.45 $X2=0 $Y2=0
cc_145 N_A1_M1001_g N_A2_c_211_n 0.00883233f $X=1.63 $Y=0.45 $X2=0 $Y2=0
cc_146 N_A1_M1001_g A2 6.3923e-19 $X=1.63 $Y=0.45 $X2=0 $Y2=0
cc_147 N_A1_M1005_g N_A_56_412#_c_297_n 0.00101902f $X=1.22 $Y=2.56 $X2=0 $Y2=0
cc_148 N_A1_M1005_g N_A_56_412#_c_303_n 0.0161597f $X=1.22 $Y=2.56 $X2=0 $Y2=0
cc_149 A1 N_A_56_412#_c_303_n 0.0200549f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A1_c_168_n N_A_56_412#_c_303_n 0.00741867f $X=1.63 $Y=1.735 $X2=0 $Y2=0
cc_151 N_A1_M1005_g N_A_163_412#_c_333_n 0.0145964f $X=1.22 $Y=2.56 $X2=0 $Y2=0
cc_152 N_A1_M1005_g N_A_163_412#_c_337_n 0.0152493f $X=1.22 $Y=2.56 $X2=0 $Y2=0
cc_153 N_A1_M1005_g N_A_163_412#_c_336_n 0.00216412f $X=1.22 $Y=2.56 $X2=0 $Y2=0
cc_154 N_A1_M1005_g N_VPWR_c_364_n 0.0103965f $X=1.22 $Y=2.56 $X2=0 $Y2=0
cc_155 N_A1_M1005_g N_VPWR_c_365_n 0.006023f $X=1.22 $Y=2.56 $X2=0 $Y2=0
cc_156 N_A1_M1005_g N_VPWR_c_363_n 0.00714345f $X=1.22 $Y=2.56 $X2=0 $Y2=0
cc_157 N_A1_M1001_g N_Y_c_407_n 0.0069097f $X=1.63 $Y=0.45 $X2=0 $Y2=0
cc_158 N_A1_M1001_g N_Y_c_400_n 0.0027886f $X=1.63 $Y=0.45 $X2=0 $Y2=0
cc_159 N_A1_M1001_g N_Y_c_402_n 0.00829842f $X=1.63 $Y=0.45 $X2=0 $Y2=0
cc_160 N_A1_M1001_g N_VGND_c_454_n 0.00177613f $X=1.63 $Y=0.45 $X2=0 $Y2=0
cc_161 N_A1_M1001_g N_VGND_c_457_n 0.00413457f $X=1.63 $Y=0.45 $X2=0 $Y2=0
cc_162 N_A1_M1001_g N_VGND_c_459_n 0.0060902f $X=1.63 $Y=0.45 $X2=0 $Y2=0
cc_163 N_A2_M1000_g N_C1_M1006_g 0.0110388f $X=2.02 $Y=0.45 $X2=0 $Y2=0
cc_164 A2 N_C1_M1006_g 0.0059368f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A2_c_213_n N_C1_M1006_g 0.00430305f $X=2.11 $Y=1.165 $X2=0 $Y2=0
cc_166 A2 C1 0.0216047f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_167 A2 N_C1_c_257_n 0.00214021f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_168 N_A2_c_213_n N_C1_c_257_n 7.37406e-19 $X=2.11 $Y=1.165 $X2=0 $Y2=0
cc_169 N_A2_M1002_g N_A_56_412#_c_303_n 0.0161698f $X=2.04 $Y=2.56 $X2=0 $Y2=0
cc_170 N_A2_M1002_g N_A_56_412#_c_298_n 0.00101902f $X=2.04 $Y=2.56 $X2=0 $Y2=0
cc_171 N_A2_M1002_g N_A_163_412#_c_337_n 0.0177091f $X=2.04 $Y=2.56 $X2=0 $Y2=0
cc_172 N_A2_M1002_g N_A_163_412#_c_334_n 0.0155289f $X=2.04 $Y=2.56 $X2=0 $Y2=0
cc_173 N_A2_M1002_g N_VPWR_c_364_n 0.00541898f $X=2.04 $Y=2.56 $X2=0 $Y2=0
cc_174 N_A2_M1002_g N_VPWR_c_367_n 0.00671212f $X=2.04 $Y=2.56 $X2=0 $Y2=0
cc_175 N_A2_M1002_g N_VPWR_c_363_n 0.00927607f $X=2.04 $Y=2.56 $X2=0 $Y2=0
cc_176 N_A2_M1000_g N_Y_c_407_n 0.00146956f $X=2.02 $Y=0.45 $X2=0 $Y2=0
cc_177 N_A2_M1000_g N_Y_c_402_n 0.0129088f $X=2.02 $Y=0.45 $X2=0 $Y2=0
cc_178 A2 N_Y_c_402_n 0.0605415f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A2_c_213_n N_Y_c_402_n 0.00428262f $X=2.11 $Y=1.165 $X2=0 $Y2=0
cc_180 N_A2_M1000_g N_VGND_c_454_n 0.00962855f $X=2.02 $Y=0.45 $X2=0 $Y2=0
cc_181 N_A2_M1000_g N_VGND_c_457_n 0.00351853f $X=2.02 $Y=0.45 $X2=0 $Y2=0
cc_182 N_A2_M1000_g N_VGND_c_459_n 0.00411872f $X=2.02 $Y=0.45 $X2=0 $Y2=0
cc_183 N_C1_M1004_g N_A_56_412#_c_298_n 0.0211288f $X=3.1 $Y=2.56 $X2=0 $Y2=0
cc_184 C1 N_A_56_412#_c_298_n 0.00208435f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_185 N_C1_M1004_g N_VPWR_c_367_n 0.00848972f $X=3.1 $Y=2.56 $X2=0 $Y2=0
cc_186 N_C1_M1004_g N_VPWR_c_363_n 0.0159211f $X=3.1 $Y=2.56 $X2=0 $Y2=0
cc_187 N_C1_M1004_g N_Y_c_404_n 0.0132603f $X=3.1 $Y=2.56 $X2=0 $Y2=0
cc_188 N_C1_M1004_g N_Y_c_405_n 0.00540303f $X=3.1 $Y=2.56 $X2=0 $Y2=0
cc_189 N_C1_c_255_n N_Y_c_405_n 3.64752e-19 $X=3.11 $Y=1.78 $X2=0 $Y2=0
cc_190 C1 N_Y_c_405_n 0.00461083f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_191 N_C1_M1004_g N_Y_c_401_n 0.00801731f $X=3.1 $Y=2.56 $X2=0 $Y2=0
cc_192 N_C1_M1003_g N_Y_c_401_n 0.0127397f $X=3.23 $Y=0.45 $X2=0 $Y2=0
cc_193 C1 N_Y_c_401_n 0.0355945f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_194 N_C1_c_257_n N_Y_c_401_n 0.0108474f $X=3.11 $Y=1.275 $X2=0 $Y2=0
cc_195 N_C1_M1006_g N_Y_c_402_n 0.0170597f $X=2.87 $Y=0.45 $X2=0 $Y2=0
cc_196 C1 N_Y_c_402_n 0.0183259f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_197 N_C1_M1006_g N_Y_c_403_n 0.00842918f $X=2.87 $Y=0.45 $X2=0 $Y2=0
cc_198 N_C1_M1003_g N_Y_c_403_n 0.0201421f $X=3.23 $Y=0.45 $X2=0 $Y2=0
cc_199 N_C1_c_254_n N_Y_c_403_n 2.1341e-19 $X=3.23 $Y=1.185 $X2=0 $Y2=0
cc_200 N_C1_M1006_g N_VGND_c_454_n 0.00426152f $X=2.87 $Y=0.45 $X2=0 $Y2=0
cc_201 N_C1_M1006_g N_VGND_c_458_n 0.0042308f $X=2.87 $Y=0.45 $X2=0 $Y2=0
cc_202 N_C1_M1003_g N_VGND_c_458_n 0.00356594f $X=3.23 $Y=0.45 $X2=0 $Y2=0
cc_203 N_C1_M1006_g N_VGND_c_459_n 0.00656972f $X=2.87 $Y=0.45 $X2=0 $Y2=0
cc_204 N_C1_M1003_g N_VGND_c_459_n 0.00624301f $X=3.23 $Y=0.45 $X2=0 $Y2=0
cc_205 N_A_56_412#_c_303_n N_A_163_412#_M1010_d 0.00814128f $X=2.67 $Y=2.165
+ $X2=-0.19 $Y2=1.655
cc_206 N_A_56_412#_c_303_n N_A_163_412#_M1002_d 0.00358885f $X=2.67 $Y=2.165
+ $X2=0 $Y2=0
cc_207 N_A_56_412#_c_297_n N_A_163_412#_c_333_n 0.0306062f $X=0.425 $Y=2.9 $X2=0
+ $Y2=0
cc_208 N_A_56_412#_c_303_n N_A_163_412#_c_337_n 0.0772981f $X=2.67 $Y=2.165
+ $X2=0 $Y2=0
cc_209 N_A_56_412#_c_298_n N_A_163_412#_c_337_n 0.0119061f $X=2.835 $Y=2.245
+ $X2=0 $Y2=0
cc_210 N_A_56_412#_c_297_n N_A_163_412#_c_336_n 0.0119061f $X=0.425 $Y=2.9 $X2=0
+ $Y2=0
cc_211 N_A_56_412#_c_303_n N_A_163_412#_c_336_n 0.0164853f $X=2.67 $Y=2.165
+ $X2=0 $Y2=0
cc_212 N_A_56_412#_c_298_n N_A_163_412#_c_334_n 0.0306062f $X=2.835 $Y=2.245
+ $X2=0 $Y2=0
cc_213 N_A_56_412#_c_303_n N_VPWR_M1005_d 0.0117008f $X=2.67 $Y=2.165 $X2=-0.19
+ $Y2=1.655
cc_214 N_A_56_412#_c_297_n N_VPWR_c_365_n 0.0220321f $X=0.425 $Y=2.9 $X2=0 $Y2=0
cc_215 N_A_56_412#_c_298_n N_VPWR_c_367_n 0.021949f $X=2.835 $Y=2.245 $X2=0
+ $Y2=0
cc_216 N_A_56_412#_c_297_n N_VPWR_c_363_n 0.0125808f $X=0.425 $Y=2.9 $X2=0 $Y2=0
cc_217 N_A_56_412#_c_298_n N_VPWR_c_363_n 0.0124703f $X=2.835 $Y=2.245 $X2=0
+ $Y2=0
cc_218 N_A_56_412#_c_298_n N_Y_c_405_n 0.067826f $X=2.835 $Y=2.245 $X2=0 $Y2=0
cc_219 N_A_163_412#_c_337_n N_VPWR_M1005_d 0.013214f $X=2.14 $Y=2.515 $X2=-0.19
+ $Y2=1.655
cc_220 N_A_163_412#_c_333_n N_VPWR_c_364_n 0.0187788f $X=0.955 $Y=2.6 $X2=0
+ $Y2=0
cc_221 N_A_163_412#_c_337_n N_VPWR_c_364_n 0.0200431f $X=2.14 $Y=2.515 $X2=0
+ $Y2=0
cc_222 N_A_163_412#_c_334_n N_VPWR_c_364_n 0.00973677f $X=2.305 $Y=2.6 $X2=0
+ $Y2=0
cc_223 N_A_163_412#_c_333_n N_VPWR_c_365_n 0.0218366f $X=0.955 $Y=2.6 $X2=0
+ $Y2=0
cc_224 N_A_163_412#_c_337_n N_VPWR_c_365_n 0.00263072f $X=2.14 $Y=2.515 $X2=0
+ $Y2=0
cc_225 N_A_163_412#_c_337_n N_VPWR_c_367_n 0.00637271f $X=2.14 $Y=2.515 $X2=0
+ $Y2=0
cc_226 N_A_163_412#_c_334_n N_VPWR_c_367_n 0.0218366f $X=2.305 $Y=2.6 $X2=0
+ $Y2=0
cc_227 N_A_163_412#_c_333_n N_VPWR_c_363_n 0.0124467f $X=0.955 $Y=2.6 $X2=0
+ $Y2=0
cc_228 N_A_163_412#_c_337_n N_VPWR_c_363_n 0.0175205f $X=2.14 $Y=2.515 $X2=0
+ $Y2=0
cc_229 N_A_163_412#_c_334_n N_VPWR_c_363_n 0.0124467f $X=2.305 $Y=2.6 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_367_n N_Y_c_404_n 0.0345056f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_231 N_VPWR_c_363_n N_Y_c_404_n 0.019739f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_232 N_Y_c_402_n N_VGND_M1000_d 0.00874616f $X=3.005 $Y=0.542 $X2=0 $Y2=0
cc_233 N_Y_c_407_n N_VGND_c_453_n 0.0110342f $X=1.415 $Y=0.47 $X2=0 $Y2=0
cc_234 N_Y_c_400_n N_VGND_c_453_n 9.50772e-19 $X=1.58 $Y=0.735 $X2=0 $Y2=0
cc_235 N_Y_c_407_n N_VGND_c_454_n 0.00649454f $X=1.415 $Y=0.47 $X2=0 $Y2=0
cc_236 N_Y_c_402_n N_VGND_c_454_n 0.0195747f $X=3.005 $Y=0.542 $X2=0 $Y2=0
cc_237 N_Y_c_403_n N_VGND_c_454_n 0.00668766f $X=3.63 $Y=0.542 $X2=0 $Y2=0
cc_238 N_Y_c_407_n N_VGND_c_457_n 0.0195017f $X=1.415 $Y=0.47 $X2=0 $Y2=0
cc_239 N_Y_c_402_n N_VGND_c_457_n 0.00712994f $X=3.005 $Y=0.542 $X2=0 $Y2=0
cc_240 N_Y_c_402_n N_VGND_c_458_n 0.00916988f $X=3.005 $Y=0.542 $X2=0 $Y2=0
cc_241 N_Y_c_403_n N_VGND_c_458_n 0.0422076f $X=3.63 $Y=0.542 $X2=0 $Y2=0
cc_242 N_Y_M1009_d N_VGND_c_459_n 0.00613083f $X=1.165 $Y=0.24 $X2=0 $Y2=0
cc_243 N_Y_M1003_d N_VGND_c_459_n 0.00231257f $X=3.305 $Y=0.24 $X2=0 $Y2=0
cc_244 N_Y_c_407_n N_VGND_c_459_n 0.0125116f $X=1.415 $Y=0.47 $X2=0 $Y2=0
cc_245 N_Y_c_402_n N_VGND_c_459_n 0.030431f $X=3.005 $Y=0.542 $X2=0 $Y2=0
cc_246 N_Y_c_403_n N_VGND_c_459_n 0.0266149f $X=3.63 $Y=0.542 $X2=0 $Y2=0
cc_247 N_Y_c_402_n A_341_48# 0.00223195f $X=3.005 $Y=0.542 $X2=-0.19 $Y2=-0.245
cc_248 N_Y_c_403_n A_589_48# 0.00622478f $X=3.63 $Y=0.542 $X2=-0.19 $Y2=-0.245
cc_249 N_VGND_c_459_n A_155_48# 0.010279f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_250 N_VGND_c_459_n A_341_48# 0.00284298f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_251 N_VGND_c_459_n A_589_48# 0.0019186f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
