* File: sky130_fd_sc_lp__srsdfrtp_1.pxi.spice
* Created: Wed Sep  2 10:39:14 2020
* 
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%SCE N_SCE_M1003_g N_SCE_M1034_g N_SCE_c_360_n
+ N_SCE_c_365_n N_SCE_M1017_g N_SCE_M1040_g N_SCE_c_362_n N_SCE_c_367_n SCE SCE
+ N_SCE_c_363_n PM_SKY130_FD_SC_LP__SRSDFRTP_1%SCE
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%D N_D_M1039_g N_D_M1021_g D N_D_c_421_n
+ N_D_c_422_n PM_SKY130_FD_SC_LP__SRSDFRTP_1%D
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_27_110# N_A_27_110#_M1003_s
+ N_A_27_110#_M1034_s N_A_27_110#_M1010_g N_A_27_110#_M1008_g
+ N_A_27_110#_c_457_n N_A_27_110#_c_458_n N_A_27_110#_c_459_n
+ N_A_27_110#_c_460_n N_A_27_110#_c_461_n N_A_27_110#_c_462_n
+ N_A_27_110#_c_463_n N_A_27_110#_c_464_n N_A_27_110#_c_465_n
+ N_A_27_110#_c_466_n PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_27_110#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%SCD N_SCD_c_542_n N_SCD_M1019_g N_SCD_c_543_n
+ N_SCD_M1009_g N_SCD_c_544_n SCD N_SCD_c_546_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%SCD
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_969_318# N_A_969_318#_M1029_d
+ N_A_969_318#_M1013_d N_A_969_318#_M1000_g N_A_969_318#_M1033_g
+ N_A_969_318#_c_580_n N_A_969_318#_M1035_g N_A_969_318#_c_581_n
+ N_A_969_318#_c_582_n N_A_969_318#_c_583_n N_A_969_318#_M1026_g
+ N_A_969_318#_c_592_n N_A_969_318#_c_593_n N_A_969_318#_M1005_g
+ N_A_969_318#_c_594_n N_A_969_318#_c_595_n N_A_969_318#_c_596_n
+ N_A_969_318#_c_597_n N_A_969_318#_c_612_p N_A_969_318#_c_584_n
+ N_A_969_318#_c_599_n N_A_969_318#_c_600_n N_A_969_318#_c_585_n
+ N_A_969_318#_c_586_n N_A_969_318#_c_602_n N_A_969_318#_c_608_p
+ N_A_969_318#_c_587_n N_A_969_318#_c_603_n N_A_969_318#_c_588_n
+ N_A_969_318#_c_604_n N_A_969_318#_c_605_n N_A_969_318#_c_589_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_969_318#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_1176_349# N_A_1176_349#_M1046_s
+ N_A_1176_349#_M1035_s N_A_1176_349#_M1001_s N_A_1176_349#_M1038_d
+ N_A_1176_349#_M1020_g N_A_1176_349#_M1050_g N_A_1176_349#_c_770_n
+ N_A_1176_349#_c_785_n N_A_1176_349#_c_771_n N_A_1176_349#_c_772_n
+ N_A_1176_349#_c_773_n N_A_1176_349#_c_787_n N_A_1176_349#_c_774_n
+ N_A_1176_349#_c_775_n N_A_1176_349#_c_776_n N_A_1176_349#_c_777_n
+ N_A_1176_349#_c_778_n N_A_1176_349#_c_779_n N_A_1176_349#_c_780_n
+ N_A_1176_349#_c_781_n N_A_1176_349#_c_782_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_1176_349#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_999_424# N_A_999_424#_M1033_d
+ N_A_999_424#_M1000_d N_A_999_424#_M1043_d N_A_999_424#_M1001_g
+ N_A_999_424#_c_925_n N_A_999_424#_M1046_g N_A_999_424#_c_926_n
+ N_A_999_424#_c_933_n N_A_999_424#_c_934_n N_A_999_424#_c_927_n
+ N_A_999_424#_c_928_n N_A_999_424#_c_937_n N_A_999_424#_c_929_n
+ N_A_999_424#_c_930_n PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_999_424#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_2176_99# N_A_2176_99#_M1006_s
+ N_A_2176_99#_M1041_d N_A_2176_99#_c_1020_n N_A_2176_99#_M1011_g
+ N_A_2176_99#_c_1021_n N_A_2176_99#_M1002_g N_A_2176_99#_M1022_g
+ N_A_2176_99#_c_1023_n N_A_2176_99#_c_1024_n N_A_2176_99#_c_1034_n
+ N_A_2176_99#_c_1025_n N_A_2176_99#_c_1035_n N_A_2176_99#_c_1036_n
+ N_A_2176_99#_c_1026_n N_A_2176_99#_c_1027_n N_A_2176_99#_c_1028_n
+ N_A_2176_99#_c_1029_n N_A_2176_99#_c_1030_n N_A_2176_99#_c_1031_n
+ N_A_2176_99#_c_1032_n N_A_2176_99#_c_1040_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_2176_99#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_1098_271# N_A_1098_271#_M1048_s
+ N_A_1098_271#_M1024_d N_A_1098_271#_M1004_g N_A_1098_271#_c_1144_n
+ N_A_1098_271#_M1032_g N_A_1098_271#_c_1159_n N_A_1098_271#_c_1160_n
+ N_A_1098_271#_M1013_g N_A_1098_271#_c_1162_n N_A_1098_271#_M1029_g
+ N_A_1098_271#_M1037_g N_A_1098_271#_c_1164_n N_A_1098_271#_c_1165_n
+ N_A_1098_271#_c_1166_n N_A_1098_271#_M1018_g N_A_1098_271#_M1038_g
+ N_A_1098_271#_c_1169_n N_A_1098_271#_c_1170_n N_A_1098_271#_c_1147_n
+ N_A_1098_271#_c_1148_n N_A_1098_271#_c_1172_n N_A_1098_271#_c_1173_n
+ N_A_1098_271#_c_1174_n N_A_1098_271#_c_1175_n N_A_1098_271#_c_1176_n
+ N_A_1098_271#_c_1149_n N_A_1098_271#_c_1150_n N_A_1098_271#_c_1151_n
+ N_A_1098_271#_c_1152_n N_A_1098_271#_c_1153_n N_A_1098_271#_c_1154_n
+ N_A_1098_271#_c_1280_p N_A_1098_271#_c_1155_n N_A_1098_271#_c_1156_n
+ N_A_1098_271#_c_1157_n PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_1098_271#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_1982_397# N_A_1982_397#_M1026_d
+ N_A_1982_397#_M1037_s N_A_1982_397#_M1005_s N_A_1982_397#_M1006_g
+ N_A_1982_397#_M1044_g N_A_1982_397#_M1015_g N_A_1982_397#_M1051_g
+ N_A_1982_397#_M1031_g N_A_1982_397#_c_1374_n N_A_1982_397#_c_1384_n
+ N_A_1982_397#_c_1385_n N_A_1982_397#_c_1386_n N_A_1982_397#_c_1408_n
+ N_A_1982_397#_c_1387_n N_A_1982_397#_c_1388_n N_A_1982_397#_c_1389_n
+ N_A_1982_397#_c_1390_n N_A_1982_397#_c_1391_n N_A_1982_397#_c_1392_n
+ N_A_1982_397#_c_1393_n N_A_1982_397#_c_1375_n N_A_1982_397#_c_1376_n
+ N_A_1982_397#_c_1536_p N_A_1982_397#_c_1377_n N_A_1982_397#_c_1378_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_1982_397#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_2586_249# N_A_2586_249#_M1012_s
+ N_A_2586_249#_M1025_d N_A_2586_249#_M1047_g N_A_2586_249#_c_1585_n
+ N_A_2586_249#_M1036_g N_A_2586_249#_c_1569_n N_A_2586_249#_c_1570_n
+ N_A_2586_249#_c_1571_n N_A_2586_249#_c_1572_n N_A_2586_249#_c_1573_n
+ N_A_2586_249#_c_1574_n N_A_2586_249#_c_1575_n N_A_2586_249#_c_1576_n
+ N_A_2586_249#_c_1577_n N_A_2586_249#_c_1578_n N_A_2586_249#_c_1579_n
+ N_A_2586_249#_c_1580_n N_A_2586_249#_c_1581_n N_A_2586_249#_c_1582_n
+ N_A_2586_249#_c_1583_n N_A_2586_249#_c_1584_n N_A_2586_249#_c_1588_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_2586_249#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%RESET_B N_RESET_B_M1023_g N_RESET_B_M1045_g
+ N_RESET_B_c_1721_n N_RESET_B_c_1722_n N_RESET_B_c_1723_n N_RESET_B_M1043_g
+ N_RESET_B_c_1739_n N_RESET_B_c_1740_n N_RESET_B_M1042_g N_RESET_B_c_1725_n
+ N_RESET_B_c_1726_n N_RESET_B_M1007_g N_RESET_B_c_1728_n N_RESET_B_c_1729_n
+ N_RESET_B_M1041_g N_RESET_B_c_1731_n N_RESET_B_c_1732_n N_RESET_B_c_1733_n
+ N_RESET_B_c_1734_n RESET_B N_RESET_B_c_1736_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%RESET_B
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%CLK N_CLK_M1048_g N_CLK_M1024_g CLK
+ N_CLK_c_1889_n PM_SKY130_FD_SC_LP__SRSDFRTP_1%CLK
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%SLEEP_B N_SLEEP_B_c_1931_n N_SLEEP_B_M1028_g
+ N_SLEEP_B_M1027_g N_SLEEP_B_c_1933_n N_SLEEP_B_M1030_g N_SLEEP_B_c_1934_n
+ N_SLEEP_B_c_1935_n N_SLEEP_B_c_1944_n N_SLEEP_B_M1025_g N_SLEEP_B_c_1936_n
+ N_SLEEP_B_M1012_g N_SLEEP_B_M1014_g N_SLEEP_B_c_1939_n N_SLEEP_B_c_1940_n
+ SLEEP_B N_SLEEP_B_c_1942_n PM_SKY130_FD_SC_LP__SRSDFRTP_1%SLEEP_B
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_3751_367# N_A_3751_367#_M1031_d
+ N_A_3751_367#_M1051_s N_A_3751_367#_M1016_g N_A_3751_367#_M1049_g
+ N_A_3751_367#_c_2023_n N_A_3751_367#_c_2024_n N_A_3751_367#_c_2025_n
+ N_A_3751_367#_c_2026_n N_A_3751_367#_c_2032_n N_A_3751_367#_c_2027_n
+ N_A_3751_367#_c_2028_n N_A_3751_367#_c_2029_n N_A_3751_367#_c_2030_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_3751_367#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%VPWR N_VPWR_M1034_d N_VPWR_M1009_d
+ N_VPWR_M1020_d N_VPWR_M1001_d N_VPWR_M1051_d N_VPWR_c_2094_n N_VPWR_c_2095_n
+ N_VPWR_c_2096_n N_VPWR_c_2097_n N_VPWR_c_2098_n N_VPWR_c_2099_n
+ N_VPWR_c_2100_n N_VPWR_c_2101_n N_VPWR_c_2102_n N_VPWR_c_2103_n
+ N_VPWR_c_2104_n VPWR N_VPWR_c_2105_n N_VPWR_c_2106_n N_VPWR_c_2107_n
+ N_VPWR_c_2093_n N_VPWR_c_2109_n N_VPWR_c_2110_n VPWR
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%VPWR
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_332_136# N_A_332_136#_M1040_d
+ N_A_332_136#_M1032_d N_A_332_136#_M1039_d N_A_332_136#_M1045_d
+ N_A_332_136#_c_2249_n N_A_332_136#_c_2239_n N_A_332_136#_c_2240_n
+ N_A_332_136#_c_2266_n N_A_332_136#_c_2267_n N_A_332_136#_c_2241_n
+ N_A_332_136#_c_2251_n N_A_332_136#_c_2252_n N_A_332_136#_c_2242_n
+ N_A_332_136#_c_2243_n N_A_332_136#_c_2244_n N_A_332_136#_c_2245_n
+ N_A_332_136#_c_2246_n N_A_332_136#_c_2247_n N_A_332_136#_c_2248_n
+ N_A_332_136#_c_2254_n N_A_332_136#_c_2255_n N_A_332_136#_c_2256_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_332_136#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%KAPWR N_KAPWR_M1022_d N_KAPWR_M1015_d
+ N_KAPWR_M1027_d KAPWR N_KAPWR_c_2379_n N_KAPWR_c_2380_n N_KAPWR_c_2381_n
+ N_KAPWR_c_2382_n KAPWR PM_SKY130_FD_SC_LP__SRSDFRTP_1%KAPWR
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%Q N_Q_M1049_d N_Q_M1016_d N_Q_c_2504_n Q Q Q Q
+ Q N_Q_c_2503_n PM_SKY130_FD_SC_LP__SRSDFRTP_1%Q
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%VGND N_VGND_M1003_d N_VGND_M1023_s
+ N_VGND_M1042_d N_VGND_M1046_d N_VGND_M1002_d N_VGND_M1047_d N_VGND_M1030_d
+ N_VGND_M1014_d N_VGND_M1049_s N_VGND_c_2525_n N_VGND_c_2526_n N_VGND_c_2527_n
+ N_VGND_c_2528_n N_VGND_c_2529_n N_VGND_c_2530_n N_VGND_c_2531_n
+ N_VGND_c_2532_n N_VGND_c_2533_n N_VGND_c_2534_n N_VGND_c_2535_n
+ N_VGND_c_2536_n N_VGND_c_2537_n N_VGND_c_2538_n N_VGND_c_2539_n
+ N_VGND_c_2540_n N_VGND_c_2541_n N_VGND_c_2542_n VGND N_VGND_c_2543_n
+ N_VGND_c_2544_n N_VGND_c_2545_n N_VGND_c_2546_n N_VGND_c_2547_n
+ N_VGND_c_2548_n N_VGND_c_2549_n N_VGND_c_2550_n N_VGND_c_2551_n
+ N_VGND_c_2552_n N_VGND_c_2553_n VGND PM_SKY130_FD_SC_LP__SRSDFRTP_1%VGND
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%noxref_29 N_noxref_29_M1040_s
+ N_noxref_29_M1019_d N_noxref_29_c_2697_n N_noxref_29_c_2698_n
+ N_noxref_29_c_2699_n N_noxref_29_c_2700_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%noxref_29
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%noxref_31 N_noxref_31_M1010_d
+ N_noxref_31_M1023_d N_noxref_31_c_2726_n N_noxref_31_c_2723_n
+ N_noxref_31_c_2724_n N_noxref_31_c_2725_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%noxref_31
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_929_152# N_A_929_152#_M1033_s
+ N_A_929_152#_M1050_s N_A_929_152#_c_2755_n N_A_929_152#_c_2756_n
+ N_A_929_152#_c_2757_n N_A_929_152#_c_2758_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_929_152#
x_PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_2544_119# N_A_2544_119#_M1044_d
+ N_A_2544_119#_M1007_d N_A_2544_119#_c_2791_n N_A_2544_119#_c_2792_n
+ N_A_2544_119#_c_2793_n N_A_2544_119#_c_2794_n
+ PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_2544_119#
cc_1 VNB N_SCE_M1003_g 0.0546885f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.76
cc_2 VNB N_SCE_c_360_n 0.0398906f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.525
cc_3 VNB N_SCE_M1040_g 0.0378673f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.89
cc_4 VNB N_SCE_c_362_n 0.0243125f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.525
cc_5 VNB N_SCE_c_363_n 0.00398477f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.665
cc_6 VNB N_D_M1021_g 0.0387357f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.65
cc_7 VNB N_A_27_110#_M1010_g 0.0358051f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.525
cc_8 VNB N_A_27_110#_c_457_n 0.028881f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=1.45
cc_9 VNB N_A_27_110#_c_458_n 0.013883f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.6
cc_10 VNB N_A_27_110#_c_459_n 0.03092f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.02
cc_11 VNB N_A_27_110#_c_460_n 0.00199251f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_12 VNB N_A_27_110#_c_461_n 0.00675089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_110#_c_462_n 9.54542e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_110#_c_463_n 0.00406647f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.665
cc_15 VNB N_A_27_110#_c_464_n 0.00994965f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.665
cc_16 VNB N_A_27_110#_c_465_n 0.00267785f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.035
cc_17 VNB N_A_27_110#_c_466_n 0.00869422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SCD_c_542_n 0.0194666f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.45
cc_19 VNB N_SCD_c_543_n 0.0131567f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.17
cc_20 VNB N_SCD_c_544_n 0.0212656f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.095
cc_21 VNB SCD 0.00100628f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.65
cc_22 VNB N_SCD_c_546_n 0.0196288f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.89
cc_23 VNB N_A_969_318#_M1033_g 0.0298781f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.17
cc_24 VNB N_A_969_318#_c_580_n 0.016926f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.65
cc_25 VNB N_A_969_318#_c_581_n 0.0279899f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.89
cc_26 VNB N_A_969_318#_c_582_n 0.0559694f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.89
cc_27 VNB N_A_969_318#_c_583_n 0.015643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_969_318#_c_584_n 0.0100194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_969_318#_c_585_n 0.0103595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_969_318#_c_586_n 0.00200328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_969_318#_c_587_n 0.0176683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_969_318#_c_588_n 0.0151666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_969_318#_c_589_n 0.0123912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_1176_349#_M1050_g 0.017829f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.6
cc_35 VNB N_A_1176_349#_c_770_n 0.0122779f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.02
cc_36 VNB N_A_1176_349#_c_771_n 0.00761172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1176_349#_c_772_n 0.065245f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.665
cc_38 VNB N_A_1176_349#_c_773_n 0.00147945f $X=-0.19 $Y=-0.245 $X2=0.77
+ $Y2=1.665
cc_39 VNB N_A_1176_349#_c_774_n 0.00698728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1176_349#_c_775_n 0.00438058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1176_349#_c_776_n 0.0167696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1176_349#_c_777_n 0.0175119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1176_349#_c_778_n 0.0366016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1176_349#_c_779_n 0.00961883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1176_349#_c_780_n 0.0109112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1176_349#_c_781_n 0.015236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1176_349#_c_782_n 5.9046e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_999_424#_c_925_n 0.0204098f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.65
cc_49 VNB N_A_999_424#_c_926_n 0.00377347f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.89
cc_50 VNB N_A_999_424#_c_927_n 0.00383185f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.02
cc_51 VNB N_A_999_424#_c_928_n 0.0045334f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_52 VNB N_A_999_424#_c_929_n 5.63519e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_999_424#_c_930_n 0.0434417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_2176_99#_c_1020_n 0.0120728f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.65
cc_55 VNB N_A_2176_99#_c_1021_n 0.0166105f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.525
cc_56 VNB N_A_2176_99#_M1022_g 0.00355372f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.65
cc_57 VNB N_A_2176_99#_c_1023_n 0.0274109f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.6
cc_58 VNB N_A_2176_99#_c_1024_n 0.00173091f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.02
cc_59 VNB N_A_2176_99#_c_1025_n 0.0244793f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_60 VNB N_A_2176_99#_c_1026_n 0.00924148f $X=-0.19 $Y=-0.245 $X2=0.77
+ $Y2=1.665
cc_61 VNB N_A_2176_99#_c_1027_n 0.00410747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_2176_99#_c_1028_n 7.13627e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_2176_99#_c_1029_n 0.018051f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.035
cc_64 VNB N_A_2176_99#_c_1030_n 2.63885e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_2176_99#_c_1031_n 0.0329838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_2176_99#_c_1032_n 0.0544015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1098_271#_M1004_g 0.00715535f $X=-0.19 $Y=-0.245 $X2=0.95
+ $Y2=1.525
cc_68 VNB N_A_1098_271#_c_1144_n 0.0175583f $X=-0.19 $Y=-0.245 $X2=1.415
+ $Y2=2.095
cc_69 VNB N_A_1098_271#_M1029_g 0.0559454f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.095
cc_70 VNB N_A_1098_271#_M1018_g 0.0474129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1098_271#_c_1147_n 0.0156692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1098_271#_c_1148_n 0.00839164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1098_271#_c_1149_n 0.0113398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1098_271#_c_1150_n 0.0323877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1098_271#_c_1151_n 0.00394924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1098_271#_c_1152_n 0.00505936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1098_271#_c_1153_n 0.0107567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1098_271#_c_1154_n 0.0133001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1098_271#_c_1155_n 0.00329003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1098_271#_c_1156_n 0.00313042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1098_271#_c_1157_n 0.0194646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1982_397#_M1006_g 0.0496585f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.095
cc_83 VNB N_A_1982_397#_M1044_g 0.0410131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1982_397#_M1051_g 5.51943e-19 $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=2.095
cc_85 VNB N_A_1982_397#_M1031_g 0.0470731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1982_397#_c_1374_n 0.0142089f $X=-0.19 $Y=-0.245 $X2=0.77
+ $Y2=1.665
cc_87 VNB N_A_1982_397#_c_1375_n 0.0227518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1982_397#_c_1376_n 0.00450723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1982_397#_c_1377_n 0.00180903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1982_397#_c_1378_n 0.037577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2586_249#_M1047_g 0.0224774f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.525
cc_92 VNB N_A_2586_249#_c_1569_n 0.0489631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2586_249#_c_1570_n 0.0266813f $X=-0.19 $Y=-0.245 $X2=1.585
+ $Y2=1.45
cc_94 VNB N_A_2586_249#_c_1571_n 0.0409455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2586_249#_c_1572_n 0.0209528f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.02
cc_96 VNB N_A_2586_249#_c_1573_n 0.0209568f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=2.095
cc_97 VNB N_A_2586_249#_c_1574_n 0.0036935f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_98 VNB N_A_2586_249#_c_1575_n 0.00407549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2586_249#_c_1576_n 0.0344644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2586_249#_c_1577_n 0.00728984f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.665
cc_101 VNB N_A_2586_249#_c_1578_n 4.61089e-19 $X=-0.19 $Y=-0.245 $X2=0.77
+ $Y2=1.665
cc_102 VNB N_A_2586_249#_c_1579_n 0.00911265f $X=-0.19 $Y=-0.245 $X2=0.77
+ $Y2=1.665
cc_103 VNB N_A_2586_249#_c_1580_n 6.1061e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2586_249#_c_1581_n 0.0111868f $X=-0.19 $Y=-0.245 $X2=0.77
+ $Y2=2.035
cc_105 VNB N_A_2586_249#_c_1582_n 0.00791577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2586_249#_c_1583_n 0.0379986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2586_249#_c_1584_n 0.00655103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_RESET_B_M1023_g 0.0469365f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.76
cc_109 VNB N_RESET_B_c_1721_n 0.0784575f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.525
cc_110 VNB N_RESET_B_c_1722_n 0.16983f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=2.095
cc_111 VNB N_RESET_B_c_1723_n 0.0125974f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.095
cc_112 VNB N_RESET_B_M1042_g 0.0283265f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.525
cc_113 VNB N_RESET_B_c_1725_n 0.0211407f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.095
cc_114 VNB N_RESET_B_c_1726_n 0.490328f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_115 VNB N_RESET_B_M1007_g 0.0398434f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.665
cc_116 VNB N_RESET_B_c_1728_n 0.156211f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.665
cc_117 VNB N_RESET_B_c_1729_n 0.0121341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_RESET_B_M1041_g 0.0352041f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.035
cc_119 VNB N_RESET_B_c_1731_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_RESET_B_c_1732_n 0.0127943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_RESET_B_c_1733_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_RESET_B_c_1734_n 0.0532521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB RESET_B 8.23858e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_RESET_B_c_1736_n 0.015378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_CLK_M1048_g 0.0517621f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.76
cc_126 VNB CLK 0.00298781f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.525
cc_127 VNB N_CLK_c_1889_n 0.0197363f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.095
cc_128 VNB N_SLEEP_B_c_1931_n 0.0141606f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.45
cc_129 VNB N_SLEEP_B_M1027_g 0.0118485f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.65
cc_130 VNB N_SLEEP_B_c_1933_n 0.0170161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_SLEEP_B_c_1934_n 0.031836f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=2.095
cc_132 VNB N_SLEEP_B_c_1935_n 0.0407409f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.095
cc_133 VNB N_SLEEP_B_c_1936_n 0.0165884f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.89
cc_134 VNB N_SLEEP_B_M1012_g 0.0209001f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.02
cc_135 VNB N_SLEEP_B_M1014_g 0.0172948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_SLEEP_B_c_1939_n 0.00672496f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.665
cc_137 VNB N_SLEEP_B_c_1940_n 0.0142212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB SLEEP_B 0.00404315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_SLEEP_B_c_1942_n 0.0685871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_3751_367#_M1016_g 6.21878e-19 $X=-0.19 $Y=-0.245 $X2=1.51
+ $Y2=1.525
cc_141 VNB N_A_3751_367#_M1049_g 0.0288233f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.17
cc_142 VNB N_A_3751_367#_c_2023_n 0.00693876f $X=-0.19 $Y=-0.245 $X2=1.585
+ $Y2=1.45
cc_143 VNB N_A_3751_367#_c_2024_n 0.00132024f $X=-0.19 $Y=-0.245 $X2=1.585
+ $Y2=0.89
cc_144 VNB N_A_3751_367#_c_2025_n 0.0121458f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.6
cc_145 VNB N_A_3751_367#_c_2026_n 0.00372455f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=2.095
cc_146 VNB N_A_3751_367#_c_2027_n 0.0109992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_3751_367#_c_2028_n 0.00875879f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.665
cc_148 VNB N_A_3751_367#_c_2029_n 0.00602645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_A_3751_367#_c_2030_n 0.056016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VPWR_c_2093_n 0.860265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_A_332_136#_c_2239_n 0.00818265f $X=-0.19 $Y=-0.245 $X2=1.49
+ $Y2=2.65
cc_152 VNB N_A_332_136#_c_2240_n 6.34478e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_A_332_136#_c_2241_n 0.00716785f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.6
cc_154 VNB N_A_332_136#_c_2242_n 0.00228882f $X=-0.19 $Y=-0.245 $X2=0.77
+ $Y2=1.665
cc_155 VNB N_A_332_136#_c_2243_n 0.0143079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_A_332_136#_c_2244_n 0.00280128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_A_332_136#_c_2245_n 4.15415e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_A_332_136#_c_2246_n 0.0135566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_A_332_136#_c_2247_n 0.00223139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_A_332_136#_c_2248_n 0.0127454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_Q_c_2503_n 0.0587923f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.02
cc_162 VNB N_VGND_c_2525_n 0.0238155f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.665
cc_163 VNB N_VGND_c_2526_n 0.0231485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2527_n 0.00799757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2528_n 0.0218039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2529_n 0.018072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2530_n 0.0123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2531_n 0.0132895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2532_n 0.0076789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2533_n 0.0218598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2534_n 0.00749576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2535_n 0.0655137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2536_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2537_n 0.0800561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2538_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2539_n 0.0169652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2540_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2541_n 0.0778393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2542_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2543_n 0.0178086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2544_n 0.0404597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2545_n 0.101325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2546_n 0.0289799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2547_n 0.0186878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2548_n 1.00794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_VGND_c_2549_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2550_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_VGND_c_2551_n 0.00632231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_189 VNB N_VGND_c_2552_n 0.00458122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_190 VNB N_VGND_c_2553_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_191 VNB N_noxref_29_c_2697_n 0.0126552f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.525
cc_192 VNB N_noxref_29_c_2698_n 0.0524472f $X=-0.19 $Y=-0.245 $X2=1.415
+ $Y2=2.095
cc_193 VNB N_noxref_29_c_2699_n 0.00508641f $X=-0.19 $Y=-0.245 $X2=0.95
+ $Y2=2.095
cc_194 VNB N_noxref_29_c_2700_n 0.0134866f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.65
cc_195 VNB N_noxref_31_c_2723_n 0.0354663f $X=-0.19 $Y=-0.245 $X2=1.415
+ $Y2=2.095
cc_196 VNB N_noxref_31_c_2724_n 0.00523306f $X=-0.19 $Y=-0.245 $X2=0.95
+ $Y2=2.095
cc_197 VNB N_noxref_31_c_2725_n 0.00960466f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.65
cc_198 VNB N_A_929_152#_c_2755_n 0.0157943f $X=-0.19 $Y=-0.245 $X2=1.51
+ $Y2=1.525
cc_199 VNB N_A_929_152#_c_2756_n 0.0388478f $X=-0.19 $Y=-0.245 $X2=1.415
+ $Y2=2.095
cc_200 VNB N_A_929_152#_c_2757_n 0.00339766f $X=-0.19 $Y=-0.245 $X2=0.95
+ $Y2=2.095
cc_201 VNB N_A_929_152#_c_2758_n 0.0100666f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.65
cc_202 VNB N_A_2544_119#_c_2791_n 0.00196087f $X=-0.19 $Y=-0.245 $X2=1.51
+ $Y2=1.525
cc_203 VNB N_A_2544_119#_c_2792_n 0.00782682f $X=-0.19 $Y=-0.245 $X2=1.415
+ $Y2=2.095
cc_204 VNB N_A_2544_119#_c_2793_n 0.00326783f $X=-0.19 $Y=-0.245 $X2=0.95
+ $Y2=2.095
cc_205 VNB N_A_2544_119#_c_2794_n 0.00243084f $X=-0.19 $Y=-0.245 $X2=1.49
+ $Y2=2.65
cc_206 VPB N_SCE_M1034_g 0.0267996f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.65
cc_207 VPB N_SCE_c_365_n 0.0371548f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=2.095
cc_208 VPB N_SCE_M1017_g 0.0217466f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_209 VPB N_SCE_c_367_n 0.0172831f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.095
cc_210 VPB SCE 0.00177942f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_211 VPB N_SCE_c_363_n 0.0330238f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.665
cc_212 VPB N_D_M1039_g 0.0232681f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.76
cc_213 VPB N_D_M1021_g 0.0130845f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.65
cc_214 VPB N_D_c_421_n 0.0473027f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.17
cc_215 VPB N_D_c_422_n 0.00824147f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_216 VPB N_A_27_110#_M1008_g 0.0368628f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.17
cc_217 VPB N_A_27_110#_c_458_n 0.0602976f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.6
cc_218 VPB N_A_27_110#_c_465_n 0.00458927f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.035
cc_219 VPB N_A_27_110#_c_466_n 0.0217254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_SCD_M1009_g 0.0473738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB SCD 0.0018235f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_222 VPB N_SCD_c_546_n 0.030263f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.89
cc_223 VPB N_A_969_318#_M1000_g 0.0239899f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.525
cc_224 VPB N_A_969_318#_c_582_n 0.00839388f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.89
cc_225 VPB N_A_969_318#_c_592_n 0.047852f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.02
cc_226 VPB N_A_969_318#_c_593_n 0.02621f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_227 VPB N_A_969_318#_c_594_n 0.00225747f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.665
cc_228 VPB N_A_969_318#_c_595_n 0.0116391f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.665
cc_229 VPB N_A_969_318#_c_596_n 0.00166874f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.665
cc_230 VPB N_A_969_318#_c_597_n 0.0176381f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.665
cc_231 VPB N_A_969_318#_c_584_n 0.0104183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_969_318#_c_599_n 0.0162341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_969_318#_c_600_n 0.0662637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_969_318#_c_586_n 0.00443824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_969_318#_c_602_n 0.00339229f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_969_318#_c_603_n 0.00704942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_969_318#_c_604_n 0.0014329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_969_318#_c_605_n 0.0588135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_969_318#_c_589_n 0.0297187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_1176_349#_M1020_g 0.022919f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_241 VPB N_A_1176_349#_c_770_n 0.00629987f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.02
cc_242 VPB N_A_1176_349#_c_785_n 0.020837f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.095
cc_243 VPB N_A_1176_349#_c_771_n 0.00253208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_1176_349#_c_787_n 0.00671003f $X=-0.19 $Y=1.655 $X2=0.77
+ $Y2=1.665
cc_245 VPB N_A_1176_349#_c_775_n 0.00412551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_1176_349#_c_780_n 0.0033602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_999_424#_M1001_g 0.0241858f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.095
cc_248 VPB N_A_999_424#_c_926_n 0.00323319f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.89
cc_249 VPB N_A_999_424#_c_933_n 0.0116415f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.89
cc_250 VPB N_A_999_424#_c_934_n 0.00999679f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.525
cc_251 VPB N_A_999_424#_c_927_n 2.17225e-19 $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.02
cc_252 VPB N_A_999_424#_c_928_n 0.00983599f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_253 VPB N_A_999_424#_c_937_n 0.00504361f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.665
cc_254 VPB N_A_999_424#_c_930_n 0.00577049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_2176_99#_M1022_g 0.0371328f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_256 VPB N_A_2176_99#_c_1034_n 0.00321512f $X=-0.19 $Y=1.655 $X2=0.72
+ $Y2=2.095
cc_257 VPB N_A_2176_99#_c_1035_n 0.0415974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_2176_99#_c_1036_n 0.00716964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_2176_99#_c_1028_n 0.00592672f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_2176_99#_c_1030_n 0.00226568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_2176_99#_c_1031_n 0.0221631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_2176_99#_c_1040_n 0.00671308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_1098_271#_M1004_g 0.0631692f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=1.525
cc_264 VPB N_A_1098_271#_c_1159_n 0.192443f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_265 VPB N_A_1098_271#_c_1160_n 0.012806f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_266 VPB N_A_1098_271#_M1013_g 0.0263966f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.89
cc_267 VPB N_A_1098_271#_c_1162_n 0.123276f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_1098_271#_M1037_g 0.0181293f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.665
cc_269 VPB N_A_1098_271#_c_1164_n 0.00908813f $X=-0.19 $Y=1.655 $X2=0.77
+ $Y2=1.665
cc_270 VPB N_A_1098_271#_c_1165_n 0.0102011f $X=-0.19 $Y=1.655 $X2=0.77
+ $Y2=1.665
cc_271 VPB N_A_1098_271#_c_1166_n 0.0110145f $X=-0.19 $Y=1.655 $X2=0.77
+ $Y2=1.665
cc_272 VPB N_A_1098_271#_M1018_g 0.00418321f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_1098_271#_M1038_g 0.0182365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_A_1098_271#_c_1169_n 0.0751883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_1098_271#_c_1170_n 0.0926124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_1098_271#_c_1148_n 0.0171496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_A_1098_271#_c_1172_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_A_1098_271#_c_1173_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_1098_271#_c_1174_n 0.0074047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_A_1098_271#_c_1175_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_A_1098_271#_c_1176_n 0.0516669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_A_1098_271#_c_1149_n 4.8095e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_A_1098_271#_c_1155_n 0.00591357f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_1098_271#_c_1156_n 0.00166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_A_1098_271#_c_1157_n 0.0170267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_A_1982_397#_M1006_g 0.0330847f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.095
cc_287 VPB N_A_1982_397#_M1044_g 0.0460584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_A_1982_397#_M1015_g 0.0302591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_289 VPB N_A_1982_397#_M1051_g 0.0273611f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.095
cc_290 VPB N_A_1982_397#_c_1374_n 0.0093581f $X=-0.19 $Y=1.655 $X2=0.77
+ $Y2=1.665
cc_291 VPB N_A_1982_397#_c_1384_n 0.0229935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB N_A_1982_397#_c_1385_n 0.0216238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 VPB N_A_1982_397#_c_1386_n 0.00969107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_A_1982_397#_c_1387_n 0.00225951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_295 VPB N_A_1982_397#_c_1388_n 0.0189972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_296 VPB N_A_1982_397#_c_1389_n 0.00227551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_A_1982_397#_c_1390_n 0.0271375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_A_1982_397#_c_1391_n 0.00210493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_A_1982_397#_c_1392_n 0.0501477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_300 VPB N_A_1982_397#_c_1393_n 3.03892e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_301 VPB N_A_1982_397#_c_1375_n 0.00668398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_302 VPB N_A_1982_397#_c_1376_n 0.00131699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_303 VPB N_A_2586_249#_c_1585_n 0.0262148f $X=-0.19 $Y=1.655 $X2=1.415
+ $Y2=2.095
cc_304 VPB N_A_2586_249#_c_1569_n 0.0094597f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_A_2586_249#_c_1581_n 5.8786e-19 $X=-0.19 $Y=1.655 $X2=0.77
+ $Y2=2.035
cc_306 VPB N_A_2586_249#_c_1588_n 0.00782847f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 VPB N_RESET_B_M1045_g 0.0527304f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.65
cc_308 VPB N_RESET_B_M1043_g 0.0292594f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_309 VPB N_RESET_B_c_1739_n 0.0280314f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=1.45
cc_310 VPB N_RESET_B_c_1740_n 0.00791731f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.89
cc_311 VPB N_RESET_B_c_1725_n 0.00402206f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.095
cc_312 VPB N_RESET_B_M1041_g 0.0309975f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.035
cc_313 VPB RESET_B 0.00333667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_314 VPB N_RESET_B_c_1736_n 0.0363398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_315 VPB N_CLK_M1024_g 0.0217441f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.65
cc_316 VPB CLK 0.00345374f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.525
cc_317 VPB N_CLK_c_1889_n 0.0172173f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.095
cc_318 VPB N_SLEEP_B_M1027_g 0.0293271f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.65
cc_319 VPB N_SLEEP_B_c_1944_n 0.011773f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_320 VPB N_SLEEP_B_M1025_g 0.0317441f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=1.45
cc_321 VPB N_SLEEP_B_c_1940_n 0.00237021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_322 VPB N_A_3751_367#_M1016_g 0.0284242f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.525
cc_323 VPB N_A_3751_367#_c_2032_n 0.0052024f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.95
cc_324 VPB N_A_3751_367#_c_2027_n 0.00422431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_2094_n 0.00675797f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.89
cc_326 VPB N_VPWR_c_2095_n 0.00944286f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.525
cc_327 VPB N_VPWR_c_2096_n 0.011888f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_328 VPB N_VPWR_c_2097_n 0.0104615f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.665
cc_329 VPB N_VPWR_c_2098_n 0.0218838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_2099_n 0.070131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2100_n 0.0060562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_2101_n 0.0713389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_2102_n 0.0043669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_2103_n 0.295548f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_2104_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_336 VPB N_VPWR_c_2105_n 0.0190361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_337 VPB N_VPWR_c_2106_n 0.037869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_338 VPB N_VPWR_c_2107_n 0.0248683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_339 VPB N_VPWR_c_2093_n 0.106326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_340 VPB N_VPWR_c_2109_n 0.00606267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_341 VPB N_VPWR_c_2110_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_342 VPB N_A_332_136#_c_2249_n 0.0141282f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_343 VPB N_A_332_136#_c_2239_n 0.00572084f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_344 VPB N_A_332_136#_c_2251_n 0.0442811f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_345 VPB N_A_332_136#_c_2252_n 0.00792057f $X=-0.19 $Y=1.655 $X2=0.72
+ $Y2=1.665
cc_346 VPB N_A_332_136#_c_2242_n 0.00670783f $X=-0.19 $Y=1.655 $X2=0.77
+ $Y2=1.665
cc_347 VPB N_A_332_136#_c_2254_n 0.00585867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_348 VPB N_A_332_136#_c_2255_n 0.00289772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_349 VPB N_A_332_136#_c_2256_n 0.00315052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_350 VPB N_KAPWR_c_2379_n 0.0029065f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.17
cc_351 VPB N_KAPWR_c_2380_n 0.0057423f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.89
cc_352 VPB N_KAPWR_c_2381_n 0.143878f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_353 VPB N_KAPWR_c_2382_n 0.0134841f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.665
cc_354 VPB N_Q_c_2504_n 0.028729f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.525
cc_355 VPB Q 0.0229617f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=2.65
cc_356 VPB N_Q_c_2503_n 0.0105239f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.02
cc_357 N_SCE_M1017_g N_D_M1039_g 0.0307482f $X=1.49 $Y=2.65 $X2=0 $Y2=0
cc_358 N_SCE_M1040_g N_D_M1021_g 0.0184568f $X=1.585 $Y=0.89 $X2=0 $Y2=0
cc_359 N_SCE_c_365_n N_D_c_421_n 0.0307482f $X=1.415 $Y=2.095 $X2=0 $Y2=0
cc_360 N_SCE_c_360_n N_D_c_422_n 5.78814e-19 $X=1.51 $Y=1.525 $X2=0 $Y2=0
cc_361 N_SCE_c_365_n N_D_c_422_n 0.00149452f $X=1.415 $Y=2.095 $X2=0 $Y2=0
cc_362 N_SCE_M1003_g N_A_27_110#_c_457_n 0.00834942f $X=0.485 $Y=0.76 $X2=0
+ $Y2=0
cc_363 N_SCE_M1003_g N_A_27_110#_c_458_n 0.00750747f $X=0.485 $Y=0.76 $X2=0
+ $Y2=0
cc_364 N_SCE_c_362_n N_A_27_110#_c_458_n 0.00776714f $X=0.68 $Y=1.525 $X2=0
+ $Y2=0
cc_365 SCE N_A_27_110#_c_458_n 0.0525325f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_366 N_SCE_c_363_n N_A_27_110#_c_458_n 0.024277f $X=0.77 $Y=1.665 $X2=0 $Y2=0
cc_367 N_SCE_M1003_g N_A_27_110#_c_459_n 0.0160015f $X=0.485 $Y=0.76 $X2=0 $Y2=0
cc_368 N_SCE_M1040_g N_A_27_110#_c_459_n 0.00865253f $X=1.585 $Y=0.89 $X2=0
+ $Y2=0
cc_369 N_SCE_c_362_n N_A_27_110#_c_459_n 0.0225043f $X=0.68 $Y=1.525 $X2=0 $Y2=0
cc_370 SCE N_A_27_110#_c_459_n 0.0261806f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_371 N_SCE_M1040_g N_A_27_110#_c_460_n 0.0145781f $X=1.585 $Y=0.89 $X2=0 $Y2=0
cc_372 N_SCE_M1040_g N_A_27_110#_c_462_n 0.0087237f $X=1.585 $Y=0.89 $X2=0 $Y2=0
cc_373 N_SCE_M1040_g N_A_27_110#_c_463_n 5.51941e-19 $X=1.585 $Y=0.89 $X2=0
+ $Y2=0
cc_374 N_SCE_M1003_g N_A_27_110#_c_464_n 0.00513266f $X=0.485 $Y=0.76 $X2=0
+ $Y2=0
cc_375 N_SCE_M1034_g N_VPWR_c_2094_n 0.0184915f $X=0.565 $Y=2.65 $X2=0 $Y2=0
cc_376 N_SCE_M1017_g N_VPWR_c_2094_n 0.0139024f $X=1.49 $Y=2.65 $X2=0 $Y2=0
cc_377 N_SCE_c_367_n N_VPWR_c_2094_n 0.00232112f $X=0.72 $Y=2.095 $X2=0 $Y2=0
cc_378 SCE N_VPWR_c_2094_n 0.0238123f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_379 N_SCE_M1017_g N_VPWR_c_2099_n 0.00469667f $X=1.49 $Y=2.65 $X2=0 $Y2=0
cc_380 N_SCE_M1034_g N_VPWR_c_2105_n 0.00405619f $X=0.565 $Y=2.65 $X2=0 $Y2=0
cc_381 N_SCE_M1034_g N_VPWR_c_2093_n 0.00318651f $X=0.565 $Y=2.65 $X2=0 $Y2=0
cc_382 N_SCE_M1017_g N_VPWR_c_2093_n 0.00357541f $X=1.49 $Y=2.65 $X2=0 $Y2=0
cc_383 N_SCE_M1034_g N_A_332_136#_c_2249_n 0.0037584f $X=0.565 $Y=2.65 $X2=0
+ $Y2=0
cc_384 N_SCE_c_365_n N_A_332_136#_c_2249_n 0.0117939f $X=1.415 $Y=2.095 $X2=0
+ $Y2=0
cc_385 N_SCE_M1017_g N_A_332_136#_c_2249_n 0.00661315f $X=1.49 $Y=2.65 $X2=0
+ $Y2=0
cc_386 SCE N_A_332_136#_c_2249_n 0.0246f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_387 N_SCE_c_363_n N_A_332_136#_c_2249_n 0.00537887f $X=0.77 $Y=1.665 $X2=0
+ $Y2=0
cc_388 N_SCE_c_360_n N_A_332_136#_c_2239_n 0.0102906f $X=1.51 $Y=1.525 $X2=0
+ $Y2=0
cc_389 N_SCE_c_365_n N_A_332_136#_c_2239_n 0.00170197f $X=1.415 $Y=2.095 $X2=0
+ $Y2=0
cc_390 N_SCE_c_360_n N_A_332_136#_c_2240_n 0.00737398f $X=1.51 $Y=1.525 $X2=0
+ $Y2=0
cc_391 SCE N_A_332_136#_c_2240_n 0.00914283f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_392 N_SCE_M1017_g N_A_332_136#_c_2266_n 0.0129464f $X=1.49 $Y=2.65 $X2=0
+ $Y2=0
cc_393 N_SCE_M1034_g N_A_332_136#_c_2267_n 6.44824e-19 $X=0.565 $Y=2.65 $X2=0
+ $Y2=0
cc_394 N_SCE_M1040_g N_A_332_136#_c_2241_n 0.00670467f $X=1.585 $Y=0.89 $X2=0
+ $Y2=0
cc_395 N_SCE_M1034_g N_KAPWR_c_2381_n 0.00600451f $X=0.565 $Y=2.65 $X2=0 $Y2=0
cc_396 N_SCE_M1017_g N_KAPWR_c_2381_n 0.00997536f $X=1.49 $Y=2.65 $X2=0 $Y2=0
cc_397 N_SCE_c_367_n N_KAPWR_c_2381_n 0.00534433f $X=0.72 $Y=2.095 $X2=0 $Y2=0
cc_398 SCE N_KAPWR_c_2381_n 0.00170664f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_399 N_SCE_M1003_g N_VGND_c_2525_n 0.0143268f $X=0.485 $Y=0.76 $X2=0 $Y2=0
cc_400 N_SCE_M1003_g N_VGND_c_2543_n 0.00379909f $X=0.485 $Y=0.76 $X2=0 $Y2=0
cc_401 N_SCE_M1003_g N_VGND_c_2548_n 0.00412152f $X=0.485 $Y=0.76 $X2=0 $Y2=0
cc_402 N_SCE_M1003_g N_noxref_29_c_2697_n 0.00126079f $X=0.485 $Y=0.76 $X2=0
+ $Y2=0
cc_403 N_SCE_M1040_g N_noxref_29_c_2697_n 0.00433482f $X=1.585 $Y=0.89 $X2=0
+ $Y2=0
cc_404 N_SCE_M1040_g N_noxref_29_c_2698_n 0.00416468f $X=1.585 $Y=0.89 $X2=0
+ $Y2=0
cc_405 N_D_M1021_g N_A_27_110#_M1010_g 0.0413666f $X=2.235 $Y=0.89 $X2=0 $Y2=0
cc_406 N_D_M1039_g N_A_27_110#_M1008_g 0.0087396f $X=1.88 $Y=2.65 $X2=0 $Y2=0
cc_407 N_D_c_421_n N_A_27_110#_M1008_g 0.00659623f $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_408 N_D_c_422_n N_A_27_110#_M1008_g 9.16554e-19 $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_409 N_D_M1021_g N_A_27_110#_c_460_n 6.9832e-19 $X=2.235 $Y=0.89 $X2=0 $Y2=0
cc_410 N_D_M1021_g N_A_27_110#_c_461_n 0.0136156f $X=2.235 $Y=0.89 $X2=0 $Y2=0
cc_411 N_D_M1021_g N_A_27_110#_c_463_n 0.0151652f $X=2.235 $Y=0.89 $X2=0 $Y2=0
cc_412 N_D_M1021_g N_A_27_110#_c_465_n 0.0104295f $X=2.235 $Y=0.89 $X2=0 $Y2=0
cc_413 N_D_c_421_n N_A_27_110#_c_465_n 0.00211691f $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_414 N_D_c_422_n N_A_27_110#_c_465_n 0.00725673f $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_415 N_D_c_421_n N_A_27_110#_c_466_n 0.0413666f $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_416 N_D_M1039_g N_VPWR_c_2099_n 0.00469667f $X=1.88 $Y=2.65 $X2=0 $Y2=0
cc_417 N_D_M1039_g N_VPWR_c_2093_n 0.00350455f $X=1.88 $Y=2.65 $X2=0 $Y2=0
cc_418 N_D_c_421_n N_A_332_136#_c_2249_n 8.2448e-19 $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_419 N_D_c_422_n N_A_332_136#_c_2249_n 0.0260833f $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_420 N_D_M1021_g N_A_332_136#_c_2239_n 0.0027846f $X=2.235 $Y=0.89 $X2=0 $Y2=0
cc_421 N_D_c_421_n N_A_332_136#_c_2239_n 0.00697375f $X=1.97 $Y=2.005 $X2=0
+ $Y2=0
cc_422 N_D_c_422_n N_A_332_136#_c_2239_n 0.0419521f $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_423 N_D_M1039_g N_A_332_136#_c_2266_n 0.0112569f $X=1.88 $Y=2.65 $X2=0 $Y2=0
cc_424 N_D_c_421_n N_A_332_136#_c_2266_n 0.0095872f $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_425 N_D_c_422_n N_A_332_136#_c_2266_n 0.0349457f $X=1.97 $Y=2.005 $X2=0 $Y2=0
cc_426 N_D_M1021_g N_A_332_136#_c_2241_n 0.00578359f $X=2.235 $Y=0.89 $X2=0
+ $Y2=0
cc_427 N_D_M1039_g N_A_332_136#_c_2254_n 0.0122783f $X=1.88 $Y=2.65 $X2=0 $Y2=0
cc_428 N_D_c_421_n N_A_332_136#_c_2254_n 2.80077e-19 $X=1.97 $Y=2.005 $X2=0
+ $Y2=0
cc_429 N_D_c_422_n N_A_332_136#_c_2254_n 0.00571315f $X=1.97 $Y=2.005 $X2=0
+ $Y2=0
cc_430 N_D_M1039_g N_KAPWR_c_2381_n 0.00869977f $X=1.88 $Y=2.65 $X2=0 $Y2=0
cc_431 N_D_M1021_g N_noxref_29_c_2698_n 0.00416656f $X=2.235 $Y=0.89 $X2=0 $Y2=0
cc_432 N_D_M1021_g N_noxref_31_c_2726_n 3.62467e-19 $X=2.235 $Y=0.89 $X2=0 $Y2=0
cc_433 N_A_27_110#_M1010_g N_SCD_c_542_n 0.0186544f $X=2.595 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_434 N_A_27_110#_M1010_g N_SCD_c_543_n 0.00661786f $X=2.595 $Y=0.89 $X2=0
+ $Y2=0
cc_435 N_A_27_110#_M1008_g N_SCD_M1009_g 0.0409224f $X=2.685 $Y=2.65 $X2=0 $Y2=0
cc_436 N_A_27_110#_c_465_n SCD 0.00964703f $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_437 N_A_27_110#_c_466_n SCD 2.56902e-19 $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_438 N_A_27_110#_c_465_n N_SCD_c_546_n 0.00159221f $X=2.715 $Y=1.765 $X2=0
+ $Y2=0
cc_439 N_A_27_110#_c_466_n N_SCD_c_546_n 0.0180819f $X=2.715 $Y=1.765 $X2=0
+ $Y2=0
cc_440 N_A_27_110#_c_458_n N_VPWR_c_2094_n 0.026558f $X=0.35 $Y=2.475 $X2=0
+ $Y2=0
cc_441 N_A_27_110#_M1008_g N_VPWR_c_2095_n 0.00227081f $X=2.685 $Y=2.65 $X2=0
+ $Y2=0
cc_442 N_A_27_110#_M1008_g N_VPWR_c_2099_n 0.00441827f $X=2.685 $Y=2.65 $X2=0
+ $Y2=0
cc_443 N_A_27_110#_c_458_n N_VPWR_c_2105_n 0.0152467f $X=0.35 $Y=2.475 $X2=0
+ $Y2=0
cc_444 N_A_27_110#_M1008_g N_VPWR_c_2093_n 0.00370097f $X=2.685 $Y=2.65 $X2=0
+ $Y2=0
cc_445 N_A_27_110#_c_458_n N_VPWR_c_2093_n 0.00323204f $X=0.35 $Y=2.475 $X2=0
+ $Y2=0
cc_446 N_A_27_110#_c_461_n N_A_332_136#_M1040_d 0.00855267f $X=2.305 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_447 N_A_27_110#_c_459_n N_A_332_136#_c_2239_n 0.0197306f $X=1.49 $Y=1.245
+ $X2=0 $Y2=0
cc_448 N_A_27_110#_c_463_n N_A_332_136#_c_2239_n 0.00654459f $X=2.39 $Y=1.6
+ $X2=0 $Y2=0
cc_449 N_A_27_110#_c_465_n N_A_332_136#_c_2239_n 0.00491831f $X=2.715 $Y=1.765
+ $X2=0 $Y2=0
cc_450 N_A_27_110#_c_459_n N_A_332_136#_c_2240_n 0.0135849f $X=1.49 $Y=1.245
+ $X2=0 $Y2=0
cc_451 N_A_27_110#_c_459_n N_A_332_136#_c_2241_n 0.0138519f $X=1.49 $Y=1.245
+ $X2=0 $Y2=0
cc_452 N_A_27_110#_c_460_n N_A_332_136#_c_2241_n 0.0162482f $X=1.575 $Y=1.16
+ $X2=0 $Y2=0
cc_453 N_A_27_110#_c_461_n N_A_332_136#_c_2241_n 0.0201769f $X=2.305 $Y=0.68
+ $X2=0 $Y2=0
cc_454 N_A_27_110#_c_463_n N_A_332_136#_c_2241_n 0.0335423f $X=2.39 $Y=1.6 $X2=0
+ $Y2=0
cc_455 N_A_27_110#_M1008_g N_A_332_136#_c_2251_n 0.00910492f $X=2.685 $Y=2.65
+ $X2=0 $Y2=0
cc_456 N_A_27_110#_c_465_n N_A_332_136#_c_2251_n 0.0179454f $X=2.715 $Y=1.765
+ $X2=0 $Y2=0
cc_457 N_A_27_110#_c_466_n N_A_332_136#_c_2251_n 0.00269047f $X=2.715 $Y=1.765
+ $X2=0 $Y2=0
cc_458 N_A_27_110#_M1008_g N_A_332_136#_c_2254_n 0.00952129f $X=2.685 $Y=2.65
+ $X2=0 $Y2=0
cc_459 N_A_27_110#_c_465_n N_A_332_136#_c_2254_n 0.0284201f $X=2.715 $Y=1.765
+ $X2=0 $Y2=0
cc_460 N_A_27_110#_c_466_n N_A_332_136#_c_2254_n 0.00245159f $X=2.715 $Y=1.765
+ $X2=0 $Y2=0
cc_461 N_A_27_110#_M1008_g N_A_332_136#_c_2255_n 0.00837722f $X=2.685 $Y=2.65
+ $X2=0 $Y2=0
cc_462 N_A_27_110#_M1034_s N_KAPWR_c_2381_n 0.00240507f $X=0.205 $Y=2.33 $X2=0
+ $Y2=0
cc_463 N_A_27_110#_M1008_g N_KAPWR_c_2381_n 0.00472621f $X=2.685 $Y=2.65 $X2=0
+ $Y2=0
cc_464 N_A_27_110#_c_458_n N_KAPWR_c_2381_n 0.0384907f $X=0.35 $Y=2.475 $X2=0
+ $Y2=0
cc_465 N_A_27_110#_c_457_n N_VGND_c_2525_n 0.0179429f $X=0.27 $Y=0.76 $X2=0
+ $Y2=0
cc_466 N_A_27_110#_c_459_n N_VGND_c_2525_n 0.0275039f $X=1.49 $Y=1.245 $X2=0
+ $Y2=0
cc_467 N_A_27_110#_c_457_n N_VGND_c_2543_n 0.00635816f $X=0.27 $Y=0.76 $X2=0
+ $Y2=0
cc_468 N_A_27_110#_c_457_n N_VGND_c_2548_n 0.00812262f $X=0.27 $Y=0.76 $X2=0
+ $Y2=0
cc_469 N_A_27_110#_c_459_n N_noxref_29_c_2697_n 0.0205583f $X=1.49 $Y=1.245
+ $X2=0 $Y2=0
cc_470 N_A_27_110#_c_462_n N_noxref_29_c_2697_n 0.0106098f $X=1.66 $Y=0.68 $X2=0
+ $Y2=0
cc_471 N_A_27_110#_M1010_g N_noxref_29_c_2698_n 0.00620038f $X=2.595 $Y=0.89
+ $X2=0 $Y2=0
cc_472 N_A_27_110#_c_461_n N_noxref_29_c_2698_n 0.0585685f $X=2.305 $Y=0.68
+ $X2=0 $Y2=0
cc_473 N_A_27_110#_c_462_n N_noxref_29_c_2698_n 0.0128284f $X=1.66 $Y=0.68 $X2=0
+ $Y2=0
cc_474 N_A_27_110#_M1010_g N_noxref_31_c_2726_n 0.0064482f $X=2.595 $Y=0.89
+ $X2=0 $Y2=0
cc_475 N_A_27_110#_c_463_n N_noxref_31_c_2726_n 0.0207609f $X=2.39 $Y=1.6 $X2=0
+ $Y2=0
cc_476 N_A_27_110#_M1010_g N_noxref_31_c_2724_n 0.00419787f $X=2.595 $Y=0.89
+ $X2=0 $Y2=0
cc_477 N_A_27_110#_c_463_n N_noxref_31_c_2724_n 0.0135839f $X=2.39 $Y=1.6 $X2=0
+ $Y2=0
cc_478 N_A_27_110#_c_465_n N_noxref_31_c_2724_n 0.0161428f $X=2.715 $Y=1.765
+ $X2=0 $Y2=0
cc_479 N_A_27_110#_c_466_n N_noxref_31_c_2724_n 0.00508216f $X=2.715 $Y=1.765
+ $X2=0 $Y2=0
cc_480 N_SCD_c_544_n N_RESET_B_M1023_g 0.00591069f $X=3.195 $Y=1.285 $X2=0 $Y2=0
cc_481 SCD RESET_B 0.0228415f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_482 N_SCD_c_546_n RESET_B 3.88475e-19 $X=3.515 $Y=1.715 $X2=0 $Y2=0
cc_483 SCD N_RESET_B_c_1736_n 0.00216533f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_484 N_SCD_c_546_n N_RESET_B_c_1736_n 0.0183293f $X=3.515 $Y=1.715 $X2=0 $Y2=0
cc_485 N_SCD_M1009_g N_VPWR_c_2095_n 0.0176721f $X=3.195 $Y=2.65 $X2=0 $Y2=0
cc_486 N_SCD_M1009_g N_VPWR_c_2099_n 0.00389963f $X=3.195 $Y=2.65 $X2=0 $Y2=0
cc_487 N_SCD_M1009_g N_VPWR_c_2093_n 0.0029773f $X=3.195 $Y=2.65 $X2=0 $Y2=0
cc_488 N_SCD_M1009_g N_A_332_136#_c_2251_n 0.0182992f $X=3.195 $Y=2.65 $X2=0
+ $Y2=0
cc_489 SCD N_A_332_136#_c_2251_n 0.0227609f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_490 N_SCD_c_546_n N_A_332_136#_c_2251_n 0.0100046f $X=3.515 $Y=1.715 $X2=0
+ $Y2=0
cc_491 N_SCD_M1009_g N_A_332_136#_c_2254_n 0.00260193f $X=3.195 $Y=2.65 $X2=0
+ $Y2=0
cc_492 N_SCD_M1009_g N_KAPWR_c_2381_n 0.00473287f $X=3.195 $Y=2.65 $X2=0 $Y2=0
cc_493 N_SCD_c_542_n N_noxref_29_c_2698_n 0.00620038f $X=3.025 $Y=1.21 $X2=0
+ $Y2=0
cc_494 N_SCD_c_542_n N_noxref_29_c_2700_n 0.00526146f $X=3.025 $Y=1.21 $X2=0
+ $Y2=0
cc_495 N_SCD_c_544_n N_noxref_29_c_2700_n 0.00310229f $X=3.195 $Y=1.285 $X2=0
+ $Y2=0
cc_496 N_SCD_c_542_n N_noxref_31_c_2726_n 0.0123681f $X=3.025 $Y=1.21 $X2=0
+ $Y2=0
cc_497 N_SCD_c_543_n N_noxref_31_c_2723_n 0.0075464f $X=3.195 $Y=1.55 $X2=0
+ $Y2=0
cc_498 N_SCD_c_544_n N_noxref_31_c_2723_n 0.0170881f $X=3.195 $Y=1.285 $X2=0
+ $Y2=0
cc_499 SCD N_noxref_31_c_2723_n 0.0275767f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_500 N_SCD_c_546_n N_noxref_31_c_2723_n 0.0104041f $X=3.515 $Y=1.715 $X2=0
+ $Y2=0
cc_501 N_SCD_c_544_n N_noxref_31_c_2724_n 0.00248047f $X=3.195 $Y=1.285 $X2=0
+ $Y2=0
cc_502 N_A_969_318#_c_597_n N_A_1176_349#_M1001_s 0.0055776f $X=7.51 $Y=2.515
+ $X2=0 $Y2=0
cc_503 N_A_969_318#_c_608_p N_A_1176_349#_M1001_s 0.00864623f $X=7.595 $Y=2.35
+ $X2=0 $Y2=0
cc_504 N_A_969_318#_c_597_n N_A_1176_349#_M1020_g 0.00695713f $X=7.51 $Y=2.515
+ $X2=0 $Y2=0
cc_505 N_A_969_318#_c_602_n N_A_1176_349#_M1020_g 0.00609327f $X=5.865 $Y=2.515
+ $X2=0 $Y2=0
cc_506 N_A_969_318#_c_597_n N_A_1176_349#_c_787_n 0.00689371f $X=7.51 $Y=2.515
+ $X2=0 $Y2=0
cc_507 N_A_969_318#_c_612_p N_A_1176_349#_c_787_n 0.029436f $X=8.395 $Y=2.35
+ $X2=0 $Y2=0
cc_508 N_A_969_318#_c_584_n N_A_1176_349#_c_787_n 0.0151578f $X=8.56 $Y=2.265
+ $X2=0 $Y2=0
cc_509 N_A_969_318#_c_608_p N_A_1176_349#_c_787_n 0.00834973f $X=7.595 $Y=2.35
+ $X2=0 $Y2=0
cc_510 N_A_969_318#_c_584_n N_A_1176_349#_c_775_n 0.0105878f $X=8.56 $Y=2.265
+ $X2=0 $Y2=0
cc_511 N_A_969_318#_c_587_n N_A_1176_349#_c_775_n 0.0204648f $X=8.99 $Y=1.5
+ $X2=0 $Y2=0
cc_512 N_A_969_318#_M1029_d N_A_1176_349#_c_776_n 0.0176259f $X=8.58 $Y=0.815
+ $X2=0 $Y2=0
cc_513 N_A_969_318#_c_580_n N_A_1176_349#_c_776_n 0.00628581f $X=9.58 $Y=1.365
+ $X2=0 $Y2=0
cc_514 N_A_969_318#_c_582_n N_A_1176_349#_c_776_n 0.00226637f $X=9.655 $Y=1.44
+ $X2=0 $Y2=0
cc_515 N_A_969_318#_c_583_n N_A_1176_349#_c_776_n 8.71358e-19 $X=9.94 $Y=1.365
+ $X2=0 $Y2=0
cc_516 N_A_969_318#_c_585_n N_A_1176_349#_c_776_n 0.0106724f $X=9.21 $Y=1.58
+ $X2=0 $Y2=0
cc_517 N_A_969_318#_c_587_n N_A_1176_349#_c_776_n 0.0416862f $X=8.99 $Y=1.5
+ $X2=0 $Y2=0
cc_518 N_A_969_318#_c_588_n N_A_1176_349#_c_776_n 0.0229025f $X=9.375 $Y=1.58
+ $X2=0 $Y2=0
cc_519 N_A_969_318#_c_580_n N_A_1176_349#_c_777_n 0.0120872f $X=9.58 $Y=1.365
+ $X2=0 $Y2=0
cc_520 N_A_969_318#_c_583_n N_A_1176_349#_c_777_n 0.00172543f $X=9.94 $Y=1.365
+ $X2=0 $Y2=0
cc_521 N_A_969_318#_c_580_n N_A_1176_349#_c_778_n 0.00307326f $X=9.58 $Y=1.365
+ $X2=0 $Y2=0
cc_522 N_A_969_318#_c_583_n N_A_1176_349#_c_778_n 0.00371137f $X=9.94 $Y=1.365
+ $X2=0 $Y2=0
cc_523 N_A_969_318#_c_594_n N_A_999_424#_M1000_d 0.00437086f $X=5.01 $Y=2.6
+ $X2=0 $Y2=0
cc_524 N_A_969_318#_c_597_n N_A_999_424#_M1043_d 0.00461301f $X=7.51 $Y=2.515
+ $X2=0 $Y2=0
cc_525 N_A_969_318#_c_597_n N_A_999_424#_M1001_g 9.57796e-19 $X=7.51 $Y=2.515
+ $X2=0 $Y2=0
cc_526 N_A_969_318#_c_612_p N_A_999_424#_M1001_g 0.0076404f $X=8.395 $Y=2.35
+ $X2=0 $Y2=0
cc_527 N_A_969_318#_c_584_n N_A_999_424#_M1001_g 0.00132904f $X=8.56 $Y=2.265
+ $X2=0 $Y2=0
cc_528 N_A_969_318#_c_599_n N_A_999_424#_M1001_g 7.62832e-19 $X=8.56 $Y=2.66
+ $X2=0 $Y2=0
cc_529 N_A_969_318#_c_608_p N_A_999_424#_M1001_g 0.0112091f $X=7.595 $Y=2.35
+ $X2=0 $Y2=0
cc_530 N_A_969_318#_c_587_n N_A_999_424#_c_925_n 5.95371e-19 $X=8.99 $Y=1.5
+ $X2=0 $Y2=0
cc_531 N_A_969_318#_M1000_g N_A_999_424#_c_926_n 5.34274e-19 $X=4.92 $Y=2.33
+ $X2=0 $Y2=0
cc_532 N_A_969_318#_M1033_g N_A_999_424#_c_926_n 0.00485762f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_533 N_A_969_318#_c_594_n N_A_999_424#_c_926_n 0.00880832f $X=5.01 $Y=2.6
+ $X2=0 $Y2=0
cc_534 N_A_969_318#_c_586_n N_A_999_424#_c_926_n 0.0248005f $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_535 N_A_969_318#_c_595_n N_A_999_424#_c_933_n 0.00730406f $X=5.78 $Y=2.685
+ $X2=0 $Y2=0
cc_536 N_A_969_318#_c_597_n N_A_999_424#_c_933_n 0.0444868f $X=7.51 $Y=2.515
+ $X2=0 $Y2=0
cc_537 N_A_969_318#_c_602_n N_A_999_424#_c_933_n 0.00783284f $X=5.865 $Y=2.515
+ $X2=0 $Y2=0
cc_538 N_A_969_318#_c_597_n N_A_999_424#_c_934_n 0.0255088f $X=7.51 $Y=2.515
+ $X2=0 $Y2=0
cc_539 N_A_969_318#_M1000_g N_A_999_424#_c_937_n 0.00114497f $X=4.92 $Y=2.33
+ $X2=0 $Y2=0
cc_540 N_A_969_318#_c_594_n N_A_999_424#_c_937_n 0.026688f $X=5.01 $Y=2.6 $X2=0
+ $Y2=0
cc_541 N_A_969_318#_c_595_n N_A_999_424#_c_937_n 0.0183581f $X=5.78 $Y=2.685
+ $X2=0 $Y2=0
cc_542 N_A_969_318#_M1033_g N_A_999_424#_c_929_n 0.00226788f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_543 N_A_969_318#_c_593_n N_A_2176_99#_M1022_g 0.0743973f $X=14.055 $Y=3.06
+ $X2=0 $Y2=0
cc_544 N_A_969_318#_c_593_n N_A_2176_99#_c_1035_n 0.016592f $X=14.055 $Y=3.06
+ $X2=0 $Y2=0
cc_545 N_A_969_318#_M1000_g N_A_1098_271#_M1004_g 0.0112284f $X=4.92 $Y=2.33
+ $X2=0 $Y2=0
cc_546 N_A_969_318#_c_594_n N_A_1098_271#_M1004_g 0.00386382f $X=5.01 $Y=2.6
+ $X2=0 $Y2=0
cc_547 N_A_969_318#_c_595_n N_A_1098_271#_M1004_g 0.0130855f $X=5.78 $Y=2.685
+ $X2=0 $Y2=0
cc_548 N_A_969_318#_c_586_n N_A_1098_271#_M1004_g 3.28011e-19 $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_549 N_A_969_318#_c_602_n N_A_1098_271#_M1004_g 0.00420918f $X=5.865 $Y=2.515
+ $X2=0 $Y2=0
cc_550 N_A_969_318#_c_589_n N_A_1098_271#_M1004_g 0.0145273f $X=5.175 $Y=1.755
+ $X2=0 $Y2=0
cc_551 N_A_969_318#_M1033_g N_A_1098_271#_c_1144_n 0.0138395f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_552 N_A_969_318#_c_595_n N_A_1098_271#_c_1159_n 8.83139e-19 $X=5.78 $Y=2.685
+ $X2=0 $Y2=0
cc_553 N_A_969_318#_c_597_n N_A_1098_271#_c_1159_n 0.0183907f $X=7.51 $Y=2.515
+ $X2=0 $Y2=0
cc_554 N_A_969_318#_c_612_p N_A_1098_271#_c_1159_n 0.00126921f $X=8.395 $Y=2.35
+ $X2=0 $Y2=0
cc_555 N_A_969_318#_c_602_n N_A_1098_271#_c_1159_n 0.00225407f $X=5.865 $Y=2.515
+ $X2=0 $Y2=0
cc_556 N_A_969_318#_c_608_p N_A_1098_271#_c_1159_n 0.00209562f $X=7.595 $Y=2.35
+ $X2=0 $Y2=0
cc_557 N_A_969_318#_c_612_p N_A_1098_271#_M1013_g 0.0119437f $X=8.395 $Y=2.35
+ $X2=0 $Y2=0
cc_558 N_A_969_318#_c_584_n N_A_1098_271#_M1013_g 0.00625005f $X=8.56 $Y=2.265
+ $X2=0 $Y2=0
cc_559 N_A_969_318#_c_599_n N_A_1098_271#_M1013_g 0.0116148f $X=8.56 $Y=2.66
+ $X2=0 $Y2=0
cc_560 N_A_969_318#_c_608_p N_A_1098_271#_M1013_g 8.30929e-19 $X=7.595 $Y=2.35
+ $X2=0 $Y2=0
cc_561 N_A_969_318#_c_603_n N_A_1098_271#_M1013_g 3.84191e-19 $X=8.56 $Y=2.31
+ $X2=0 $Y2=0
cc_562 N_A_969_318#_c_599_n N_A_1098_271#_c_1162_n 0.00507066f $X=8.56 $Y=2.66
+ $X2=0 $Y2=0
cc_563 N_A_969_318#_c_600_n N_A_1098_271#_c_1162_n 0.032404f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_564 N_A_969_318#_c_582_n N_A_1098_271#_M1029_g 0.00431482f $X=9.655 $Y=1.44
+ $X2=0 $Y2=0
cc_565 N_A_969_318#_c_584_n N_A_1098_271#_M1029_g 0.00970863f $X=8.56 $Y=2.265
+ $X2=0 $Y2=0
cc_566 N_A_969_318#_c_587_n N_A_1098_271#_M1029_g 0.0166739f $X=8.99 $Y=1.5
+ $X2=0 $Y2=0
cc_567 N_A_969_318#_c_588_n N_A_1098_271#_M1029_g 2.48905e-19 $X=9.375 $Y=1.58
+ $X2=0 $Y2=0
cc_568 N_A_969_318#_c_600_n N_A_1098_271#_M1037_g 0.00963104f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_569 N_A_969_318#_c_582_n N_A_1098_271#_c_1165_n 0.00185692f $X=9.655 $Y=1.44
+ $X2=0 $Y2=0
cc_570 N_A_969_318#_c_600_n N_A_1098_271#_c_1166_n 7.04503e-19 $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_571 N_A_969_318#_c_583_n N_A_1098_271#_M1018_g 0.0161251f $X=9.94 $Y=1.365
+ $X2=0 $Y2=0
cc_572 N_A_969_318#_c_600_n N_A_1098_271#_M1038_g 0.00963813f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_573 N_A_969_318#_c_600_n N_A_1098_271#_c_1169_n 0.01773f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_574 N_A_969_318#_c_600_n N_A_1098_271#_c_1170_n 0.0128925f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_575 N_A_969_318#_M1033_g N_A_1098_271#_c_1147_n 0.0145273f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_576 N_A_969_318#_c_584_n N_A_1098_271#_c_1148_n 0.0114009f $X=8.56 $Y=2.265
+ $X2=0 $Y2=0
cc_577 N_A_969_318#_c_593_n N_A_1098_271#_c_1176_n 0.00886372f $X=14.055 $Y=3.06
+ $X2=0 $Y2=0
cc_578 N_A_969_318#_c_582_n N_A_1982_397#_c_1374_n 0.00482965f $X=9.655 $Y=1.44
+ $X2=0 $Y2=0
cc_579 N_A_969_318#_c_583_n N_A_1982_397#_c_1374_n 0.0150241f $X=9.94 $Y=1.365
+ $X2=0 $Y2=0
cc_580 N_A_969_318#_c_588_n N_A_1982_397#_c_1374_n 0.00937484f $X=9.375 $Y=1.58
+ $X2=0 $Y2=0
cc_581 N_A_969_318#_c_600_n N_A_1982_397#_c_1384_n 0.116771f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_582 N_A_969_318#_c_592_n N_A_1982_397#_c_1385_n 0.00184928f $X=13.93 $Y=3.135
+ $X2=0 $Y2=0
cc_583 N_A_969_318#_c_600_n N_A_1982_397#_c_1385_n 0.0154973f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_584 N_A_969_318#_c_604_n N_A_1982_397#_c_1385_n 0.015121f $X=13.29 $Y=2.91
+ $X2=0 $Y2=0
cc_585 N_A_969_318#_c_605_n N_A_1982_397#_c_1385_n 0.00216756f $X=13.29 $Y=2.91
+ $X2=0 $Y2=0
cc_586 N_A_969_318#_c_592_n N_A_1982_397#_c_1386_n 0.00509533f $X=13.93 $Y=3.135
+ $X2=0 $Y2=0
cc_587 N_A_969_318#_c_593_n N_A_1982_397#_c_1386_n 0.00983975f $X=14.055 $Y=3.06
+ $X2=0 $Y2=0
cc_588 N_A_969_318#_c_604_n N_A_1982_397#_c_1386_n 0.0157068f $X=13.29 $Y=2.91
+ $X2=0 $Y2=0
cc_589 N_A_969_318#_c_605_n N_A_1982_397#_c_1386_n 0.00152069f $X=13.29 $Y=2.91
+ $X2=0 $Y2=0
cc_590 N_A_969_318#_c_593_n N_A_1982_397#_c_1408_n 0.0117837f $X=14.055 $Y=3.06
+ $X2=0 $Y2=0
cc_591 N_A_969_318#_c_581_n N_A_1982_397#_c_1390_n 0.00412192f $X=9.865 $Y=1.44
+ $X2=0 $Y2=0
cc_592 N_A_969_318#_c_600_n N_A_1982_397#_c_1390_n 0.0405383f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_593 N_A_969_318#_c_600_n N_A_1982_397#_c_1391_n 0.0235808f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_594 N_A_969_318#_c_600_n N_A_1982_397#_c_1392_n 0.00264527f $X=13.125 $Y=2.99
+ $X2=0 $Y2=0
cc_595 N_A_969_318#_c_593_n N_A_1982_397#_c_1393_n 0.00355057f $X=14.055 $Y=3.06
+ $X2=0 $Y2=0
cc_596 N_A_969_318#_c_593_n N_A_2586_249#_c_1570_n 0.00131263f $X=14.055 $Y=3.06
+ $X2=0 $Y2=0
cc_597 N_A_969_318#_M1000_g N_RESET_B_M1045_g 0.00925773f $X=4.92 $Y=2.33 $X2=0
+ $Y2=0
cc_598 N_A_969_318#_c_594_n N_RESET_B_M1045_g 2.40451e-19 $X=5.01 $Y=2.6 $X2=0
+ $Y2=0
cc_599 N_A_969_318#_M1033_g N_RESET_B_c_1721_n 0.014487f $X=5.175 $Y=1.035 $X2=0
+ $Y2=0
cc_600 N_A_969_318#_M1033_g N_RESET_B_c_1722_n 0.0031339f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_601 N_A_969_318#_c_597_n N_RESET_B_M1043_g 0.0135457f $X=7.51 $Y=2.515 $X2=0
+ $Y2=0
cc_602 N_A_969_318#_c_602_n N_RESET_B_M1043_g 4.16687e-19 $X=5.865 $Y=2.515
+ $X2=0 $Y2=0
cc_603 N_A_969_318#_c_597_n N_RESET_B_c_1739_n 0.00106966f $X=7.51 $Y=2.515
+ $X2=0 $Y2=0
cc_604 N_A_969_318#_c_580_n N_RESET_B_c_1726_n 0.00738071f $X=9.58 $Y=1.365
+ $X2=0 $Y2=0
cc_605 N_A_969_318#_c_583_n N_RESET_B_c_1726_n 0.00737233f $X=9.94 $Y=1.365
+ $X2=0 $Y2=0
cc_606 N_A_969_318#_c_589_n N_RESET_B_c_1736_n 0.0141642f $X=5.175 $Y=1.755
+ $X2=0 $Y2=0
cc_607 N_A_969_318#_c_597_n N_VPWR_M1020_d 0.00780659f $X=7.51 $Y=2.515 $X2=0
+ $Y2=0
cc_608 N_A_969_318#_c_612_p N_VPWR_M1001_d 0.0105049f $X=8.395 $Y=2.35 $X2=0
+ $Y2=0
cc_609 N_A_969_318#_c_597_n N_VPWR_c_2096_n 0.0211232f $X=7.51 $Y=2.515 $X2=0
+ $Y2=0
cc_610 N_A_969_318#_c_612_p N_VPWR_c_2097_n 0.0246974f $X=8.395 $Y=2.35 $X2=0
+ $Y2=0
cc_611 N_A_969_318#_c_599_n N_VPWR_c_2097_n 0.0229563f $X=8.56 $Y=2.66 $X2=0
+ $Y2=0
cc_612 N_A_969_318#_M1000_g N_VPWR_c_2101_n 0.00205103f $X=4.92 $Y=2.33 $X2=0
+ $Y2=0
cc_613 N_A_969_318#_c_595_n N_VPWR_c_2101_n 0.0158514f $X=5.78 $Y=2.685 $X2=0
+ $Y2=0
cc_614 N_A_969_318#_c_596_n N_VPWR_c_2101_n 0.00416831f $X=5.095 $Y=2.685 $X2=0
+ $Y2=0
cc_615 N_A_969_318#_c_597_n N_VPWR_c_2101_n 0.00203541f $X=7.51 $Y=2.515 $X2=0
+ $Y2=0
cc_616 N_A_969_318#_c_602_n N_VPWR_c_2101_n 0.00407423f $X=5.865 $Y=2.515 $X2=0
+ $Y2=0
cc_617 N_A_969_318#_c_599_n N_VPWR_c_2103_n 0.0160672f $X=8.56 $Y=2.66 $X2=0
+ $Y2=0
cc_618 N_A_969_318#_c_600_n N_VPWR_c_2103_n 0.282055f $X=13.125 $Y=2.99 $X2=0
+ $Y2=0
cc_619 N_A_969_318#_c_604_n N_VPWR_c_2103_n 0.0212434f $X=13.29 $Y=2.91 $X2=0
+ $Y2=0
cc_620 N_A_969_318#_c_605_n N_VPWR_c_2103_n 0.0293449f $X=13.29 $Y=2.91 $X2=0
+ $Y2=0
cc_621 N_A_969_318#_c_597_n N_VPWR_c_2106_n 0.0130818f $X=7.51 $Y=2.515 $X2=0
+ $Y2=0
cc_622 N_A_969_318#_c_608_p N_VPWR_c_2106_n 0.00180956f $X=7.595 $Y=2.35 $X2=0
+ $Y2=0
cc_623 N_A_969_318#_c_592_n N_VPWR_c_2093_n 0.0170595f $X=13.93 $Y=3.135 $X2=0
+ $Y2=0
cc_624 N_A_969_318#_c_595_n N_VPWR_c_2093_n 0.00233353f $X=5.78 $Y=2.685 $X2=0
+ $Y2=0
cc_625 N_A_969_318#_c_596_n N_VPWR_c_2093_n 5.23798e-19 $X=5.095 $Y=2.685 $X2=0
+ $Y2=0
cc_626 N_A_969_318#_c_599_n N_VPWR_c_2093_n 0.00195531f $X=8.56 $Y=2.66 $X2=0
+ $Y2=0
cc_627 N_A_969_318#_c_600_n N_VPWR_c_2093_n 0.0340616f $X=13.125 $Y=2.99 $X2=0
+ $Y2=0
cc_628 N_A_969_318#_c_602_n N_VPWR_c_2093_n 4.63082e-19 $X=5.865 $Y=2.515 $X2=0
+ $Y2=0
cc_629 N_A_969_318#_c_604_n N_VPWR_c_2093_n 0.00250438f $X=13.29 $Y=2.91 $X2=0
+ $Y2=0
cc_630 N_A_969_318#_c_605_n N_VPWR_c_2093_n 0.00895349f $X=13.29 $Y=2.91 $X2=0
+ $Y2=0
cc_631 N_A_969_318#_M1000_g N_A_332_136#_c_2252_n 0.0033083f $X=4.92 $Y=2.33
+ $X2=0 $Y2=0
cc_632 N_A_969_318#_c_594_n N_A_332_136#_c_2252_n 0.0244339f $X=5.01 $Y=2.6
+ $X2=0 $Y2=0
cc_633 N_A_969_318#_c_596_n N_A_332_136#_c_2252_n 0.0132787f $X=5.095 $Y=2.685
+ $X2=0 $Y2=0
cc_634 N_A_969_318#_M1033_g N_A_332_136#_c_2242_n 0.00148812f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_635 N_A_969_318#_c_594_n N_A_332_136#_c_2242_n 0.0109297f $X=5.01 $Y=2.6
+ $X2=0 $Y2=0
cc_636 N_A_969_318#_c_586_n N_A_332_136#_c_2242_n 0.0248004f $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_637 N_A_969_318#_c_589_n N_A_332_136#_c_2242_n 0.00400938f $X=5.175 $Y=1.755
+ $X2=0 $Y2=0
cc_638 N_A_969_318#_M1033_g N_A_332_136#_c_2243_n 0.00728806f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_639 N_A_969_318#_c_586_n N_A_332_136#_c_2243_n 0.0258968f $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_640 N_A_969_318#_c_589_n N_A_332_136#_c_2243_n 0.00325414f $X=5.175 $Y=1.755
+ $X2=0 $Y2=0
cc_641 N_A_969_318#_M1033_g N_A_332_136#_c_2245_n 0.013407f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_642 N_A_969_318#_M1033_g N_A_332_136#_c_2246_n 0.00360028f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_643 N_A_969_318#_M1033_g N_A_332_136#_c_2247_n 0.00234388f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_644 N_A_969_318#_M1033_g N_A_332_136#_c_2248_n 5.85323e-19 $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_645 N_A_969_318#_M1000_g N_A_332_136#_c_2256_n 0.00150797f $X=4.92 $Y=2.33
+ $X2=0 $Y2=0
cc_646 N_A_969_318#_c_594_n N_A_332_136#_c_2256_n 0.013453f $X=5.01 $Y=2.6 $X2=0
+ $Y2=0
cc_647 N_A_969_318#_c_602_n A_1128_424# 0.0017085f $X=5.865 $Y=2.515 $X2=-0.19
+ $Y2=-0.245
cc_648 N_A_969_318#_c_593_n N_KAPWR_c_2379_n 0.00106116f $X=14.055 $Y=3.06 $X2=0
+ $Y2=0
cc_649 N_A_969_318#_M1000_g N_KAPWR_c_2381_n 0.00266541f $X=4.92 $Y=2.33 $X2=0
+ $Y2=0
cc_650 N_A_969_318#_c_592_n N_KAPWR_c_2381_n 0.0010139f $X=13.93 $Y=3.135 $X2=0
+ $Y2=0
cc_651 N_A_969_318#_c_593_n N_KAPWR_c_2381_n 0.00648301f $X=14.055 $Y=3.06 $X2=0
+ $Y2=0
cc_652 N_A_969_318#_c_595_n N_KAPWR_c_2381_n 0.0317647f $X=5.78 $Y=2.685 $X2=0
+ $Y2=0
cc_653 N_A_969_318#_c_596_n N_KAPWR_c_2381_n 0.0127471f $X=5.095 $Y=2.685 $X2=0
+ $Y2=0
cc_654 N_A_969_318#_c_597_n N_KAPWR_c_2381_n 0.0578372f $X=7.51 $Y=2.515 $X2=0
+ $Y2=0
cc_655 N_A_969_318#_c_612_p N_KAPWR_c_2381_n 0.0176757f $X=8.395 $Y=2.35 $X2=0
+ $Y2=0
cc_656 N_A_969_318#_c_599_n N_KAPWR_c_2381_n 0.0374685f $X=8.56 $Y=2.66 $X2=0
+ $Y2=0
cc_657 N_A_969_318#_c_600_n N_KAPWR_c_2381_n 0.122376f $X=13.125 $Y=2.99 $X2=0
+ $Y2=0
cc_658 N_A_969_318#_c_602_n N_KAPWR_c_2381_n 0.0101588f $X=5.865 $Y=2.515 $X2=0
+ $Y2=0
cc_659 N_A_969_318#_c_608_p N_KAPWR_c_2381_n 0.00660814f $X=7.595 $Y=2.35 $X2=0
+ $Y2=0
cc_660 N_A_969_318#_c_604_n N_KAPWR_c_2381_n 0.0179696f $X=13.29 $Y=2.91 $X2=0
+ $Y2=0
cc_661 N_A_969_318#_c_605_n N_KAPWR_c_2381_n 0.00753265f $X=13.29 $Y=2.91 $X2=0
+ $Y2=0
cc_662 N_A_969_318#_M1033_g N_A_929_152#_c_2755_n 0.00132423f $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_663 N_A_969_318#_M1033_g N_A_929_152#_c_2756_n 4.19837e-19 $X=5.175 $Y=1.035
+ $X2=0 $Y2=0
cc_664 N_A_1176_349#_c_787_n N_A_999_424#_M1001_g 0.0116772f $X=7.965 $Y=1.97
+ $X2=0 $Y2=0
cc_665 N_A_1176_349#_c_774_n N_A_999_424#_c_925_n 0.00207207f $X=7.715 $Y=0.995
+ $X2=0 $Y2=0
cc_666 N_A_1176_349#_c_775_n N_A_999_424#_c_925_n 0.00917691f $X=8.05 $Y=1.845
+ $X2=0 $Y2=0
cc_667 N_A_1176_349#_c_782_n N_A_999_424#_c_925_n 0.0151309f $X=8.135 $Y=1.085
+ $X2=0 $Y2=0
cc_668 N_A_1176_349#_c_785_n N_A_999_424#_c_926_n 0.00175588f $X=6.085 $Y=1.895
+ $X2=0 $Y2=0
cc_669 N_A_1176_349#_c_771_n N_A_999_424#_c_926_n 0.0141554f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_670 N_A_1176_349#_c_772_n N_A_999_424#_c_926_n 7.48899e-19 $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_671 N_A_1176_349#_M1020_g N_A_999_424#_c_933_n 0.0135355f $X=5.955 $Y=2.33
+ $X2=0 $Y2=0
cc_672 N_A_1176_349#_c_785_n N_A_999_424#_c_933_n 0.00659912f $X=6.085 $Y=1.895
+ $X2=0 $Y2=0
cc_673 N_A_1176_349#_c_771_n N_A_999_424#_c_933_n 0.0304767f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_674 N_A_1176_349#_c_772_n N_A_999_424#_c_933_n 0.0014843f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_675 N_A_1176_349#_c_770_n N_A_999_424#_c_934_n 3.09302e-19 $X=6.085 $Y=1.745
+ $X2=0 $Y2=0
cc_676 N_A_1176_349#_c_785_n N_A_999_424#_c_934_n 2.21635e-19 $X=6.085 $Y=1.895
+ $X2=0 $Y2=0
cc_677 N_A_1176_349#_c_771_n N_A_999_424#_c_934_n 0.00493477f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_678 N_A_1176_349#_c_787_n N_A_999_424#_c_934_n 0.0174213f $X=7.965 $Y=1.97
+ $X2=0 $Y2=0
cc_679 N_A_1176_349#_c_770_n N_A_999_424#_c_927_n 6.53549e-19 $X=6.085 $Y=1.745
+ $X2=0 $Y2=0
cc_680 N_A_1176_349#_c_771_n N_A_999_424#_c_927_n 0.0258801f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_681 N_A_1176_349#_c_772_n N_A_999_424#_c_927_n 0.00124913f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_682 N_A_1176_349#_c_781_n N_A_999_424#_c_927_n 0.0265155f $X=7.59 $Y=1.085
+ $X2=0 $Y2=0
cc_683 N_A_1176_349#_c_787_n N_A_999_424#_c_928_n 0.0351535f $X=7.965 $Y=1.97
+ $X2=0 $Y2=0
cc_684 N_A_1176_349#_c_775_n N_A_999_424#_c_928_n 0.0256551f $X=8.05 $Y=1.845
+ $X2=0 $Y2=0
cc_685 N_A_1176_349#_c_781_n N_A_999_424#_c_928_n 0.0527025f $X=7.59 $Y=1.085
+ $X2=0 $Y2=0
cc_686 N_A_1176_349#_M1020_g N_A_999_424#_c_937_n 9.11387e-19 $X=5.955 $Y=2.33
+ $X2=0 $Y2=0
cc_687 N_A_1176_349#_c_787_n N_A_999_424#_c_930_n 0.00782202f $X=7.965 $Y=1.97
+ $X2=0 $Y2=0
cc_688 N_A_1176_349#_c_775_n N_A_999_424#_c_930_n 0.0109974f $X=8.05 $Y=1.845
+ $X2=0 $Y2=0
cc_689 N_A_1176_349#_c_781_n N_A_999_424#_c_930_n 0.0099934f $X=7.59 $Y=1.085
+ $X2=0 $Y2=0
cc_690 N_A_1176_349#_c_780_n N_A_2176_99#_c_1020_n 0.0164963f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_691 N_A_1176_349#_c_780_n N_A_2176_99#_c_1021_n 0.00228801f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_692 N_A_1176_349#_c_780_n N_A_2176_99#_c_1023_n 0.00502026f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_693 N_A_1176_349#_c_780_n N_A_2176_99#_c_1024_n 0.0133399f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_694 N_A_1176_349#_c_780_n N_A_2176_99#_c_1034_n 0.0536853f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_695 N_A_1176_349#_c_780_n N_A_2176_99#_c_1036_n 0.0145003f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_696 N_A_1176_349#_c_780_n N_A_2176_99#_c_1031_n 0.00413472f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_697 N_A_1176_349#_c_770_n N_A_1098_271#_M1004_g 0.00841712f $X=6.085 $Y=1.745
+ $X2=0 $Y2=0
cc_698 N_A_1176_349#_c_785_n N_A_1098_271#_M1004_g 0.0489374f $X=6.085 $Y=1.895
+ $X2=0 $Y2=0
cc_699 N_A_1176_349#_c_771_n N_A_1098_271#_M1004_g 0.00110539f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_700 N_A_1176_349#_c_771_n N_A_1098_271#_c_1144_n 7.71827e-19 $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_701 N_A_1176_349#_c_772_n N_A_1098_271#_c_1144_n 0.00859516f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_702 N_A_1176_349#_M1020_g N_A_1098_271#_c_1159_n 0.00413813f $X=5.955 $Y=2.33
+ $X2=0 $Y2=0
cc_703 N_A_1176_349#_c_787_n N_A_1098_271#_M1029_g 2.86902e-19 $X=7.965 $Y=1.97
+ $X2=0 $Y2=0
cc_704 N_A_1176_349#_c_775_n N_A_1098_271#_M1029_g 0.0048634f $X=8.05 $Y=1.845
+ $X2=0 $Y2=0
cc_705 N_A_1176_349#_c_776_n N_A_1098_271#_M1029_g 0.019797f $X=9.2 $Y=1.08
+ $X2=0 $Y2=0
cc_706 N_A_1176_349#_c_777_n N_A_1098_271#_M1029_g 0.00720239f $X=9.365 $Y=0.77
+ $X2=0 $Y2=0
cc_707 N_A_1176_349#_c_782_n N_A_1098_271#_M1029_g 2.22021e-19 $X=8.135 $Y=1.085
+ $X2=0 $Y2=0
cc_708 N_A_1176_349#_c_780_n N_A_1098_271#_M1037_g 3.41303e-19 $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_709 N_A_1176_349#_c_778_n N_A_1098_271#_M1018_g 0.00371137f $X=10.68 $Y=0.35
+ $X2=0 $Y2=0
cc_710 N_A_1176_349#_c_780_n N_A_1098_271#_M1018_g 0.0106277f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_711 N_A_1176_349#_c_780_n N_A_1098_271#_M1038_g 0.00861789f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_712 N_A_1176_349#_c_770_n N_A_1098_271#_c_1147_n 0.00558875f $X=6.085
+ $Y=1.745 $X2=0 $Y2=0
cc_713 N_A_1176_349#_c_771_n N_A_1098_271#_c_1147_n 2.66364e-19 $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_714 N_A_1176_349#_c_787_n N_A_1098_271#_c_1148_n 0.00213342f $X=7.965 $Y=1.97
+ $X2=0 $Y2=0
cc_715 N_A_1176_349#_c_780_n N_A_1098_271#_c_1174_n 0.00517966f $X=10.845
+ $Y=2.18 $X2=0 $Y2=0
cc_716 N_A_1176_349#_c_776_n N_A_1982_397#_c_1374_n 0.0078998f $X=9.2 $Y=1.08
+ $X2=0 $Y2=0
cc_717 N_A_1176_349#_c_777_n N_A_1982_397#_c_1374_n 0.0102611f $X=9.365 $Y=0.77
+ $X2=0 $Y2=0
cc_718 N_A_1176_349#_c_778_n N_A_1982_397#_c_1374_n 0.0243858f $X=10.68 $Y=0.35
+ $X2=0 $Y2=0
cc_719 N_A_1176_349#_c_780_n N_A_1982_397#_c_1374_n 0.0869913f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_720 N_A_1176_349#_M1038_d N_A_1982_397#_c_1384_n 0.00616004f $X=10.705
+ $Y=1.985 $X2=0 $Y2=0
cc_721 N_A_1176_349#_c_780_n N_A_1982_397#_c_1384_n 0.0141899f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_722 N_A_1176_349#_M1050_g N_RESET_B_c_1722_n 0.0103062f $X=6.64 $Y=0.805
+ $X2=0 $Y2=0
cc_723 N_A_1176_349#_M1020_g N_RESET_B_M1043_g 0.0187702f $X=5.955 $Y=2.33 $X2=0
+ $Y2=0
cc_724 N_A_1176_349#_c_785_n N_RESET_B_M1043_g 0.00474432f $X=6.085 $Y=1.895
+ $X2=0 $Y2=0
cc_725 N_A_1176_349#_c_787_n N_RESET_B_M1043_g 3.93817e-19 $X=7.965 $Y=1.97
+ $X2=0 $Y2=0
cc_726 N_A_1176_349#_c_781_n N_RESET_B_c_1739_n 0.00199369f $X=7.59 $Y=1.085
+ $X2=0 $Y2=0
cc_727 N_A_1176_349#_c_770_n N_RESET_B_c_1740_n 0.00474432f $X=6.085 $Y=1.745
+ $X2=0 $Y2=0
cc_728 N_A_1176_349#_c_771_n N_RESET_B_c_1740_n 0.00135542f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_729 N_A_1176_349#_c_772_n N_RESET_B_c_1740_n 0.0106489f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_730 N_A_1176_349#_c_781_n N_RESET_B_c_1740_n 4.2362e-19 $X=7.59 $Y=1.085
+ $X2=0 $Y2=0
cc_731 N_A_1176_349#_M1050_g N_RESET_B_M1042_g 0.0249094f $X=6.64 $Y=0.805 $X2=0
+ $Y2=0
cc_732 N_A_1176_349#_c_774_n N_RESET_B_M1042_g 0.00320825f $X=7.715 $Y=0.995
+ $X2=0 $Y2=0
cc_733 N_A_1176_349#_c_781_n N_RESET_B_M1042_g 0.0114668f $X=7.59 $Y=1.085 $X2=0
+ $Y2=0
cc_734 N_A_1176_349#_c_782_n N_RESET_B_M1042_g 2.5779e-19 $X=8.135 $Y=1.085
+ $X2=0 $Y2=0
cc_735 N_A_1176_349#_c_770_n N_RESET_B_c_1725_n 0.00260496f $X=6.085 $Y=1.745
+ $X2=0 $Y2=0
cc_736 N_A_1176_349#_c_771_n N_RESET_B_c_1725_n 9.73449e-19 $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_737 N_A_1176_349#_c_772_n N_RESET_B_c_1725_n 0.0117623f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_738 N_A_1176_349#_c_774_n N_RESET_B_c_1726_n 0.00486845f $X=7.715 $Y=0.995
+ $X2=0 $Y2=0
cc_739 N_A_1176_349#_c_778_n N_RESET_B_c_1726_n 0.025364f $X=10.68 $Y=0.35 $X2=0
+ $Y2=0
cc_740 N_A_1176_349#_c_779_n N_RESET_B_c_1726_n 0.00772631f $X=9.53 $Y=0.35
+ $X2=0 $Y2=0
cc_741 N_A_1176_349#_c_771_n N_RESET_B_c_1732_n 5.27831e-19 $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_742 N_A_1176_349#_c_772_n N_RESET_B_c_1732_n 0.0249094f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_743 N_A_1176_349#_c_781_n N_RESET_B_c_1732_n 0.00522933f $X=7.59 $Y=1.085
+ $X2=0 $Y2=0
cc_744 N_A_1176_349#_c_787_n N_VPWR_M1001_d 0.00744027f $X=7.965 $Y=1.97 $X2=0
+ $Y2=0
cc_745 N_A_1176_349#_M1050_g N_A_332_136#_c_2248_n 0.00377949f $X=6.64 $Y=0.805
+ $X2=0 $Y2=0
cc_746 N_A_1176_349#_c_785_n N_A_332_136#_c_2248_n 0.00277194f $X=6.085 $Y=1.895
+ $X2=0 $Y2=0
cc_747 N_A_1176_349#_c_771_n N_A_332_136#_c_2248_n 0.0137946f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_748 N_A_1176_349#_c_772_n N_A_332_136#_c_2248_n 0.00379357f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_749 N_A_1176_349#_c_773_n N_A_332_136#_c_2248_n 0.0122549f $X=6.61 $Y=1.09
+ $X2=0 $Y2=0
cc_750 N_A_1176_349#_M1001_s N_KAPWR_c_2381_n 0.00231069f $X=7.36 $Y=1.865 $X2=0
+ $Y2=0
cc_751 N_A_1176_349#_M1020_g N_KAPWR_c_2381_n 0.00163747f $X=5.955 $Y=2.33 $X2=0
+ $Y2=0
cc_752 N_A_1176_349#_c_787_n N_KAPWR_c_2381_n 0.00103274f $X=7.965 $Y=1.97 $X2=0
+ $Y2=0
cc_753 N_A_1176_349#_c_780_n N_KAPWR_c_2381_n 0.00159441f $X=10.845 $Y=2.18
+ $X2=0 $Y2=0
cc_754 N_A_1176_349#_c_781_n N_VGND_M1042_d 0.00234976f $X=7.59 $Y=1.085 $X2=0
+ $Y2=0
cc_755 N_A_1176_349#_c_775_n N_VGND_M1046_d 8.62822e-19 $X=8.05 $Y=1.845 $X2=0
+ $Y2=0
cc_756 N_A_1176_349#_c_776_n N_VGND_M1046_d 0.0124553f $X=9.2 $Y=1.08 $X2=0
+ $Y2=0
cc_757 N_A_1176_349#_c_782_n N_VGND_M1046_d 5.82151e-19 $X=8.135 $Y=1.085 $X2=0
+ $Y2=0
cc_758 N_A_1176_349#_M1050_g N_VGND_c_2527_n 0.00100708f $X=6.64 $Y=0.805 $X2=0
+ $Y2=0
cc_759 N_A_1176_349#_c_774_n N_VGND_c_2527_n 0.0182858f $X=7.715 $Y=0.995 $X2=0
+ $Y2=0
cc_760 N_A_1176_349#_c_781_n N_VGND_c_2527_n 0.0219716f $X=7.59 $Y=1.085 $X2=0
+ $Y2=0
cc_761 N_A_1176_349#_c_774_n N_VGND_c_2528_n 0.0096883f $X=7.715 $Y=0.995 $X2=0
+ $Y2=0
cc_762 N_A_1176_349#_c_782_n N_VGND_c_2528_n 0.0218628f $X=8.135 $Y=1.085 $X2=0
+ $Y2=0
cc_763 N_A_1176_349#_c_778_n N_VGND_c_2529_n 0.00783795f $X=10.68 $Y=0.35 $X2=0
+ $Y2=0
cc_764 N_A_1176_349#_c_780_n N_VGND_c_2529_n 0.0193724f $X=10.845 $Y=2.18 $X2=0
+ $Y2=0
cc_765 N_A_1176_349#_c_774_n N_VGND_c_2539_n 0.00551001f $X=7.715 $Y=0.995 $X2=0
+ $Y2=0
cc_766 N_A_1176_349#_c_778_n N_VGND_c_2541_n 0.0864978f $X=10.68 $Y=0.35 $X2=0
+ $Y2=0
cc_767 N_A_1176_349#_c_779_n N_VGND_c_2541_n 0.0222408f $X=9.53 $Y=0.35 $X2=0
+ $Y2=0
cc_768 N_A_1176_349#_M1050_g N_VGND_c_2548_n 7.85159e-19 $X=6.64 $Y=0.805 $X2=0
+ $Y2=0
cc_769 N_A_1176_349#_c_774_n N_VGND_c_2548_n 0.00671715f $X=7.715 $Y=0.995 $X2=0
+ $Y2=0
cc_770 N_A_1176_349#_c_778_n N_VGND_c_2548_n 0.0470596f $X=10.68 $Y=0.35 $X2=0
+ $Y2=0
cc_771 N_A_1176_349#_c_779_n N_VGND_c_2548_n 0.0114525f $X=9.53 $Y=0.35 $X2=0
+ $Y2=0
cc_772 N_A_1176_349#_c_773_n N_A_929_152#_M1050_s 0.00240325f $X=6.61 $Y=1.09
+ $X2=0 $Y2=0
cc_773 N_A_1176_349#_M1050_g N_A_929_152#_c_2758_n 0.00905702f $X=6.64 $Y=0.805
+ $X2=0 $Y2=0
cc_774 N_A_1176_349#_c_771_n N_A_929_152#_c_2758_n 6.17554e-19 $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_775 N_A_1176_349#_c_772_n N_A_929_152#_c_2758_n 0.00181816f $X=6.445 $Y=1.32
+ $X2=0 $Y2=0
cc_776 N_A_1176_349#_c_773_n N_A_929_152#_c_2758_n 0.022118f $X=6.61 $Y=1.09
+ $X2=0 $Y2=0
cc_777 N_A_1176_349#_c_781_n A_1343_119# 0.00366293f $X=7.59 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_778 N_A_999_424#_c_926_n N_A_1098_271#_M1004_g 0.015096f $X=5.47 $Y=2.09
+ $X2=0 $Y2=0
cc_779 N_A_999_424#_c_933_n N_A_1098_271#_M1004_g 0.00839717f $X=6.78 $Y=2.175
+ $X2=0 $Y2=0
cc_780 N_A_999_424#_c_937_n N_A_1098_271#_M1004_g 0.00593509f $X=5.555 $Y=2.26
+ $X2=0 $Y2=0
cc_781 N_A_999_424#_c_929_n N_A_1098_271#_c_1144_n 0.00239168f $X=5.46 $Y=1.1
+ $X2=0 $Y2=0
cc_782 N_A_999_424#_M1001_g N_A_1098_271#_c_1159_n 0.00863957f $X=7.72 $Y=2.285
+ $X2=0 $Y2=0
cc_783 N_A_999_424#_c_925_n N_A_1098_271#_M1029_g 0.0193918f $X=7.97 $Y=1.345
+ $X2=0 $Y2=0
cc_784 N_A_999_424#_c_930_n N_A_1098_271#_M1029_g 0.00476652f $X=7.72 $Y=1.51
+ $X2=0 $Y2=0
cc_785 N_A_999_424#_c_926_n N_A_1098_271#_c_1147_n 0.00531138f $X=5.47 $Y=2.09
+ $X2=0 $Y2=0
cc_786 N_A_999_424#_c_933_n N_A_1098_271#_c_1147_n 0.00296572f $X=6.78 $Y=2.175
+ $X2=0 $Y2=0
cc_787 N_A_999_424#_M1001_g N_A_1098_271#_c_1148_n 0.0208534f $X=7.72 $Y=2.285
+ $X2=0 $Y2=0
cc_788 N_A_999_424#_c_933_n N_RESET_B_M1043_g 0.0139104f $X=6.78 $Y=2.175 $X2=0
+ $Y2=0
cc_789 N_A_999_424#_c_934_n N_RESET_B_M1043_g 0.00866015f $X=6.945 $Y=2.09 $X2=0
+ $Y2=0
cc_790 N_A_999_424#_c_933_n N_RESET_B_c_1739_n 0.00290299f $X=6.78 $Y=2.175
+ $X2=0 $Y2=0
cc_791 N_A_999_424#_c_934_n N_RESET_B_c_1739_n 0.0187143f $X=6.945 $Y=2.09 $X2=0
+ $Y2=0
cc_792 N_A_999_424#_M1001_g N_RESET_B_c_1725_n 0.00330135f $X=7.72 $Y=2.285
+ $X2=0 $Y2=0
cc_793 N_A_999_424#_c_934_n N_RESET_B_c_1725_n 0.00173144f $X=6.945 $Y=2.09
+ $X2=0 $Y2=0
cc_794 N_A_999_424#_c_927_n N_RESET_B_c_1725_n 0.0152159f $X=7.11 $Y=1.51 $X2=0
+ $Y2=0
cc_795 N_A_999_424#_c_930_n N_RESET_B_c_1725_n 0.0107124f $X=7.72 $Y=1.51 $X2=0
+ $Y2=0
cc_796 N_A_999_424#_c_925_n N_RESET_B_c_1726_n 0.0103107f $X=7.97 $Y=1.345 $X2=0
+ $Y2=0
cc_797 N_A_999_424#_c_927_n N_RESET_B_c_1732_n 3.75015e-19 $X=7.11 $Y=1.51 $X2=0
+ $Y2=0
cc_798 N_A_999_424#_c_933_n N_VPWR_M1020_d 0.00522803f $X=6.78 $Y=2.175 $X2=0
+ $Y2=0
cc_799 N_A_999_424#_M1001_g N_VPWR_c_2097_n 0.0039878f $X=7.72 $Y=2.285 $X2=0
+ $Y2=0
cc_800 N_A_999_424#_c_926_n N_A_332_136#_c_2242_n 0.00483676f $X=5.47 $Y=2.09
+ $X2=0 $Y2=0
cc_801 N_A_999_424#_c_926_n N_A_332_136#_c_2243_n 0.0117946f $X=5.47 $Y=2.09
+ $X2=0 $Y2=0
cc_802 N_A_999_424#_c_929_n N_A_332_136#_c_2243_n 0.00120076f $X=5.46 $Y=1.1
+ $X2=0 $Y2=0
cc_803 N_A_999_424#_c_929_n N_A_332_136#_c_2245_n 0.0221858f $X=5.46 $Y=1.1
+ $X2=0 $Y2=0
cc_804 N_A_999_424#_c_929_n N_A_332_136#_c_2246_n 0.014184f $X=5.46 $Y=1.1 $X2=0
+ $Y2=0
cc_805 N_A_999_424#_c_929_n N_A_332_136#_c_2248_n 0.0131035f $X=5.46 $Y=1.1
+ $X2=0 $Y2=0
cc_806 N_A_999_424#_c_933_n A_1128_424# 0.00159108f $X=6.78 $Y=2.175 $X2=-0.19
+ $Y2=-0.245
cc_807 N_A_999_424#_M1001_g N_KAPWR_c_2381_n 0.00644124f $X=7.72 $Y=2.285 $X2=0
+ $Y2=0
cc_808 N_A_999_424#_c_933_n N_KAPWR_c_2381_n 0.00352645f $X=6.78 $Y=2.175 $X2=0
+ $Y2=0
cc_809 N_A_999_424#_c_937_n N_KAPWR_c_2381_n 0.00187211f $X=5.555 $Y=2.26 $X2=0
+ $Y2=0
cc_810 N_A_999_424#_c_925_n N_VGND_c_2527_n 0.00221113f $X=7.97 $Y=1.345 $X2=0
+ $Y2=0
cc_811 N_A_999_424#_c_925_n N_VGND_c_2528_n 0.00829167f $X=7.97 $Y=1.345 $X2=0
+ $Y2=0
cc_812 N_A_999_424#_c_925_n N_VGND_c_2548_n 7.88961e-19 $X=7.97 $Y=1.345 $X2=0
+ $Y2=0
cc_813 N_A_2176_99#_c_1020_n N_A_1098_271#_M1018_g 0.0470877f $X=10.955 $Y=1.155
+ $X2=0 $Y2=0
cc_814 N_A_2176_99#_c_1031_n N_A_1098_271#_M1018_g 0.00835505f $X=11.265 $Y=1.32
+ $X2=0 $Y2=0
cc_815 N_A_2176_99#_c_1035_n N_A_1098_271#_c_1170_n 0.0140633f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_816 N_A_2176_99#_c_1034_n N_A_1098_271#_c_1174_n 8.35275e-19 $X=11.265
+ $Y=2.01 $X2=0 $Y2=0
cc_817 N_A_2176_99#_c_1031_n N_A_1098_271#_c_1174_n 0.00265453f $X=11.265
+ $Y=1.32 $X2=0 $Y2=0
cc_818 N_A_2176_99#_M1022_g N_A_1098_271#_c_1176_n 0.0085318f $X=14.545 $Y=2.45
+ $X2=0 $Y2=0
cc_819 N_A_2176_99#_c_1025_n N_A_1098_271#_c_1176_n 0.0134748f $X=11.905 $Y=1.24
+ $X2=0 $Y2=0
cc_820 N_A_2176_99#_c_1035_n N_A_1098_271#_c_1176_n 0.181899f $X=14.695 $Y=2.095
+ $X2=0 $Y2=0
cc_821 N_A_2176_99#_c_1028_n N_A_1098_271#_c_1176_n 0.0140117f $X=14.825 $Y=2.01
+ $X2=0 $Y2=0
cc_822 N_A_2176_99#_M1022_g N_A_1098_271#_c_1149_n 0.00196646f $X=14.545 $Y=2.45
+ $X2=0 $Y2=0
cc_823 N_A_2176_99#_c_1027_n N_A_1098_271#_c_1149_n 0.0242205f $X=14.825 $Y=1.61
+ $X2=0 $Y2=0
cc_824 N_A_2176_99#_c_1028_n N_A_1098_271#_c_1149_n 0.00433327f $X=14.825
+ $Y=2.01 $X2=0 $Y2=0
cc_825 N_A_2176_99#_c_1032_n N_A_1098_271#_c_1149_n 0.0148252f $X=14.79 $Y=1.445
+ $X2=0 $Y2=0
cc_826 N_A_2176_99#_c_1027_n N_A_1098_271#_c_1150_n 0.0207781f $X=14.825 $Y=1.61
+ $X2=0 $Y2=0
cc_827 N_A_2176_99#_c_1029_n N_A_1098_271#_c_1150_n 0.038427f $X=15.645 $Y=1.525
+ $X2=0 $Y2=0
cc_828 N_A_2176_99#_c_1032_n N_A_1098_271#_c_1150_n 0.00877308f $X=14.79
+ $Y=1.445 $X2=0 $Y2=0
cc_829 N_A_2176_99#_c_1034_n N_A_1098_271#_c_1156_n 0.0209762f $X=11.265 $Y=2.01
+ $X2=0 $Y2=0
cc_830 N_A_2176_99#_c_1025_n N_A_1098_271#_c_1156_n 0.023754f $X=11.905 $Y=1.24
+ $X2=0 $Y2=0
cc_831 N_A_2176_99#_c_1035_n N_A_1098_271#_c_1156_n 0.0242156f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_832 N_A_2176_99#_c_1031_n N_A_1098_271#_c_1156_n 0.00109712f $X=11.265
+ $Y=1.32 $X2=0 $Y2=0
cc_833 N_A_2176_99#_c_1034_n N_A_1098_271#_c_1157_n 0.00743562f $X=11.265
+ $Y=2.01 $X2=0 $Y2=0
cc_834 N_A_2176_99#_c_1025_n N_A_1098_271#_c_1157_n 0.00231265f $X=11.905
+ $Y=1.24 $X2=0 $Y2=0
cc_835 N_A_2176_99#_c_1035_n N_A_1098_271#_c_1157_n 0.00126186f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_836 N_A_2176_99#_c_1031_n N_A_1098_271#_c_1157_n 0.0191963f $X=11.265 $Y=1.32
+ $X2=0 $Y2=0
cc_837 N_A_2176_99#_c_1035_n N_A_1982_397#_M1005_s 0.00577375f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_838 N_A_2176_99#_c_1025_n N_A_1982_397#_M1006_g 0.00776047f $X=11.905 $Y=1.24
+ $X2=0 $Y2=0
cc_839 N_A_2176_99#_c_1035_n N_A_1982_397#_M1006_g 0.0106348f $X=14.695 $Y=2.095
+ $X2=0 $Y2=0
cc_840 N_A_2176_99#_c_1026_n N_A_1982_397#_M1006_g 0.0133078f $X=12.07 $Y=0.805
+ $X2=0 $Y2=0
cc_841 N_A_2176_99#_c_1025_n N_A_1982_397#_M1044_g 8.4399e-19 $X=11.905 $Y=1.24
+ $X2=0 $Y2=0
cc_842 N_A_2176_99#_c_1035_n N_A_1982_397#_M1044_g 0.0120466f $X=14.695 $Y=2.095
+ $X2=0 $Y2=0
cc_843 N_A_2176_99#_c_1026_n N_A_1982_397#_M1044_g 0.00158673f $X=12.07 $Y=0.805
+ $X2=0 $Y2=0
cc_844 N_A_2176_99#_c_1030_n N_A_1982_397#_M1015_g 0.00146054f $X=15.73 $Y=1.93
+ $X2=0 $Y2=0
cc_845 N_A_2176_99#_c_1040_n N_A_1982_397#_M1015_g 0.00489453f $X=15.915
+ $Y=2.095 $X2=0 $Y2=0
cc_846 N_A_2176_99#_c_1035_n N_A_1982_397#_c_1384_n 0.0272138f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_847 N_A_2176_99#_c_1036_n N_A_1982_397#_c_1384_n 0.0130984f $X=11.43 $Y=2.095
+ $X2=0 $Y2=0
cc_848 N_A_2176_99#_c_1035_n N_A_1982_397#_c_1385_n 0.0775194f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_849 N_A_2176_99#_M1022_g N_A_1982_397#_c_1386_n 0.00155797f $X=14.545 $Y=2.45
+ $X2=0 $Y2=0
cc_850 N_A_2176_99#_M1041_d N_A_1982_397#_c_1408_n 0.00387959f $X=15.775 $Y=1.95
+ $X2=0 $Y2=0
cc_851 N_A_2176_99#_M1022_g N_A_1982_397#_c_1408_n 0.0150892f $X=14.545 $Y=2.45
+ $X2=0 $Y2=0
cc_852 N_A_2176_99#_c_1035_n N_A_1982_397#_c_1408_n 0.0576028f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_853 N_A_2176_99#_c_1040_n N_A_1982_397#_c_1408_n 0.0223136f $X=15.915
+ $Y=2.095 $X2=0 $Y2=0
cc_854 N_A_2176_99#_c_1030_n N_A_1982_397#_c_1387_n 0.00671998f $X=15.73 $Y=1.93
+ $X2=0 $Y2=0
cc_855 N_A_2176_99#_c_1040_n N_A_1982_397#_c_1387_n 0.0182049f $X=15.915
+ $Y=2.095 $X2=0 $Y2=0
cc_856 N_A_2176_99#_c_1035_n N_A_1982_397#_c_1391_n 0.0236714f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_857 N_A_2176_99#_c_1035_n N_A_1982_397#_c_1392_n 2.11484e-19 $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_858 N_A_2176_99#_c_1035_n N_A_1982_397#_c_1393_n 0.0212734f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_859 N_A_2176_99#_c_1029_n N_A_1982_397#_c_1375_n 6.41702e-19 $X=15.645
+ $Y=1.525 $X2=0 $Y2=0
cc_860 N_A_2176_99#_c_1030_n N_A_1982_397#_c_1375_n 3.74884e-19 $X=15.73 $Y=1.93
+ $X2=0 $Y2=0
cc_861 N_A_2176_99#_c_1040_n N_A_1982_397#_c_1375_n 0.00156437f $X=15.915
+ $Y=2.095 $X2=0 $Y2=0
cc_862 N_A_2176_99#_c_1029_n N_A_1982_397#_c_1376_n 0.0146833f $X=15.645
+ $Y=1.525 $X2=0 $Y2=0
cc_863 N_A_2176_99#_c_1030_n N_A_1982_397#_c_1376_n 0.0099142f $X=15.73 $Y=1.93
+ $X2=0 $Y2=0
cc_864 N_A_2176_99#_c_1040_n N_A_1982_397#_c_1376_n 0.00666601f $X=15.915
+ $Y=2.095 $X2=0 $Y2=0
cc_865 N_A_2176_99#_M1022_g N_A_2586_249#_c_1585_n 0.0346351f $X=14.545 $Y=2.45
+ $X2=0 $Y2=0
cc_866 N_A_2176_99#_c_1035_n N_A_2586_249#_c_1585_n 0.00535987f $X=14.695
+ $Y=2.095 $X2=0 $Y2=0
cc_867 N_A_2176_99#_c_1028_n N_A_2586_249#_c_1585_n 0.00493391f $X=14.825
+ $Y=2.01 $X2=0 $Y2=0
cc_868 N_A_2176_99#_c_1029_n N_A_2586_249#_c_1585_n 0.00397563f $X=15.645
+ $Y=1.525 $X2=0 $Y2=0
cc_869 N_A_2176_99#_c_1040_n N_A_2586_249#_c_1585_n 0.00130986f $X=15.915
+ $Y=2.095 $X2=0 $Y2=0
cc_870 N_A_2176_99#_M1022_g N_A_2586_249#_c_1569_n 0.00327278f $X=14.545 $Y=2.45
+ $X2=0 $Y2=0
cc_871 N_A_2176_99#_c_1027_n N_A_2586_249#_c_1569_n 0.00107347f $X=14.825
+ $Y=1.61 $X2=0 $Y2=0
cc_872 N_A_2176_99#_c_1028_n N_A_2586_249#_c_1569_n 0.00488505f $X=14.825
+ $Y=2.01 $X2=0 $Y2=0
cc_873 N_A_2176_99#_c_1029_n N_A_2586_249#_c_1569_n 0.0149634f $X=15.645
+ $Y=1.525 $X2=0 $Y2=0
cc_874 N_A_2176_99#_c_1030_n N_A_2586_249#_c_1569_n 0.00165938f $X=15.73 $Y=1.93
+ $X2=0 $Y2=0
cc_875 N_A_2176_99#_c_1032_n N_A_2586_249#_c_1569_n 0.0205536f $X=14.79 $Y=1.445
+ $X2=0 $Y2=0
cc_876 N_A_2176_99#_c_1032_n N_A_2586_249#_c_1570_n 0.00119511f $X=14.79
+ $Y=1.445 $X2=0 $Y2=0
cc_877 N_A_2176_99#_c_1032_n N_A_2586_249#_c_1572_n 2.33182e-19 $X=14.79
+ $Y=1.445 $X2=0 $Y2=0
cc_878 N_A_2176_99#_c_1032_n N_A_2586_249#_c_1573_n 5.67104e-19 $X=14.79
+ $Y=1.445 $X2=0 $Y2=0
cc_879 N_A_2176_99#_c_1020_n N_RESET_B_c_1726_n 0.00851956f $X=10.955 $Y=1.155
+ $X2=0 $Y2=0
cc_880 N_A_2176_99#_c_1021_n N_RESET_B_c_1726_n 0.00894529f $X=11.315 $Y=1.155
+ $X2=0 $Y2=0
cc_881 N_A_2176_99#_c_1026_n N_RESET_B_c_1726_n 0.00624358f $X=12.07 $Y=0.805
+ $X2=0 $Y2=0
cc_882 N_A_2176_99#_c_1029_n N_RESET_B_M1041_g 0.0161567f $X=15.645 $Y=1.525
+ $X2=0 $Y2=0
cc_883 N_A_2176_99#_c_1030_n N_RESET_B_M1041_g 0.00983261f $X=15.73 $Y=1.93
+ $X2=0 $Y2=0
cc_884 N_A_2176_99#_c_1040_n N_RESET_B_M1041_g 0.00926612f $X=15.915 $Y=2.095
+ $X2=0 $Y2=0
cc_885 N_A_2176_99#_M1022_g N_VPWR_c_2103_n 0.0079122f $X=14.545 $Y=2.45 $X2=0
+ $Y2=0
cc_886 N_A_2176_99#_M1022_g N_VPWR_c_2093_n 0.00531456f $X=14.545 $Y=2.45 $X2=0
+ $Y2=0
cc_887 N_A_2176_99#_c_1035_n A_2836_390# 0.00265407f $X=14.695 $Y=2.095
+ $X2=-0.19 $Y2=-0.245
cc_888 N_A_2176_99#_c_1035_n N_KAPWR_M1022_d 0.00566444f $X=14.695 $Y=2.095
+ $X2=-0.19 $Y2=-0.245
cc_889 N_A_2176_99#_c_1028_n N_KAPWR_M1022_d 0.00103572f $X=14.825 $Y=2.01
+ $X2=-0.19 $Y2=-0.245
cc_890 N_A_2176_99#_M1022_g N_KAPWR_c_2379_n 0.00970035f $X=14.545 $Y=2.45 $X2=0
+ $Y2=0
cc_891 N_A_2176_99#_M1041_d N_KAPWR_c_2381_n 0.00368941f $X=15.775 $Y=1.95 $X2=0
+ $Y2=0
cc_892 N_A_2176_99#_M1022_g N_KAPWR_c_2381_n 0.00424289f $X=14.545 $Y=2.45 $X2=0
+ $Y2=0
cc_893 N_A_2176_99#_c_1035_n N_KAPWR_c_2381_n 0.00962656f $X=14.695 $Y=2.095
+ $X2=0 $Y2=0
cc_894 N_A_2176_99#_c_1036_n N_KAPWR_c_2381_n 0.00223406f $X=11.43 $Y=2.095
+ $X2=0 $Y2=0
cc_895 N_A_2176_99#_c_1020_n N_VGND_c_2529_n 0.0013145f $X=10.955 $Y=1.155 $X2=0
+ $Y2=0
cc_896 N_A_2176_99#_c_1021_n N_VGND_c_2529_n 0.0107827f $X=11.315 $Y=1.155 $X2=0
+ $Y2=0
cc_897 N_A_2176_99#_c_1024_n N_VGND_c_2529_n 0.00368231f $X=11.265 $Y=1.325
+ $X2=0 $Y2=0
cc_898 N_A_2176_99#_c_1025_n N_VGND_c_2529_n 0.0210806f $X=11.905 $Y=1.24 $X2=0
+ $Y2=0
cc_899 N_A_2176_99#_c_1026_n N_VGND_c_2529_n 0.0294413f $X=12.07 $Y=0.805 $X2=0
+ $Y2=0
cc_900 N_A_2176_99#_c_1026_n N_VGND_c_2544_n 0.00749462f $X=12.07 $Y=0.805 $X2=0
+ $Y2=0
cc_901 N_A_2176_99#_c_1020_n N_VGND_c_2548_n 6.35988e-19 $X=10.955 $Y=1.155
+ $X2=0 $Y2=0
cc_902 N_A_2176_99#_c_1021_n N_VGND_c_2548_n 7.97988e-19 $X=11.315 $Y=1.155
+ $X2=0 $Y2=0
cc_903 N_A_2176_99#_c_1026_n N_VGND_c_2548_n 0.00907254f $X=12.07 $Y=0.805 $X2=0
+ $Y2=0
cc_904 N_A_2176_99#_c_1026_n N_A_2544_119#_c_2791_n 0.013252f $X=12.07 $Y=0.805
+ $X2=0 $Y2=0
cc_905 N_A_2176_99#_c_1026_n N_A_2544_119#_c_2793_n 0.00603269f $X=12.07
+ $Y=0.805 $X2=0 $Y2=0
cc_906 N_A_1098_271#_c_1170_n N_A_1982_397#_M1006_g 0.0262347f $X=11.715
+ $Y=3.075 $X2=0 $Y2=0
cc_907 N_A_1098_271#_c_1176_n N_A_1982_397#_M1006_g 0.013686f $X=14.355 $Y=1.755
+ $X2=0 $Y2=0
cc_908 N_A_1098_271#_c_1156_n N_A_1982_397#_M1006_g 0.00115306f $X=11.805
+ $Y=1.675 $X2=0 $Y2=0
cc_909 N_A_1098_271#_c_1157_n N_A_1982_397#_M1006_g 0.0182617f $X=11.805
+ $Y=1.675 $X2=0 $Y2=0
cc_910 N_A_1098_271#_c_1176_n N_A_1982_397#_M1044_g 0.0161386f $X=14.355
+ $Y=1.755 $X2=0 $Y2=0
cc_911 N_A_1098_271#_M1037_g N_A_1982_397#_c_1374_n 0.00421653f $X=10.27
+ $Y=2.405 $X2=0 $Y2=0
cc_912 N_A_1098_271#_c_1164_n N_A_1982_397#_c_1374_n 0.00882072f $X=10.52 $Y=1.8
+ $X2=0 $Y2=0
cc_913 N_A_1098_271#_c_1165_n N_A_1982_397#_c_1374_n 0.00735402f $X=10.345
+ $Y=1.8 $X2=0 $Y2=0
cc_914 N_A_1098_271#_M1018_g N_A_1982_397#_c_1374_n 0.0134313f $X=10.595
+ $Y=0.835 $X2=0 $Y2=0
cc_915 N_A_1098_271#_M1038_g N_A_1982_397#_c_1374_n 0.00201847f $X=10.63
+ $Y=2.405 $X2=0 $Y2=0
cc_916 N_A_1098_271#_M1038_g N_A_1982_397#_c_1384_n 0.0139556f $X=10.63 $Y=2.405
+ $X2=0 $Y2=0
cc_917 N_A_1098_271#_c_1170_n N_A_1982_397#_c_1384_n 0.0137416f $X=11.715
+ $Y=3.075 $X2=0 $Y2=0
cc_918 N_A_1098_271#_M1024_d N_A_1982_397#_c_1388_n 0.00402013f $X=16.85 $Y=1.95
+ $X2=0 $Y2=0
cc_919 N_A_1098_271#_c_1280_p N_A_1982_397#_c_1388_n 0.0334554f $X=17.325
+ $Y=2.095 $X2=0 $Y2=0
cc_920 N_A_1098_271#_M1037_g N_A_1982_397#_c_1390_n 0.0158707f $X=10.27 $Y=2.405
+ $X2=0 $Y2=0
cc_921 N_A_1098_271#_M1038_g N_A_1982_397#_c_1390_n 2.55458e-19 $X=10.63
+ $Y=2.405 $X2=0 $Y2=0
cc_922 N_A_1098_271#_c_1170_n N_A_1982_397#_c_1391_n 0.00144051f $X=11.715
+ $Y=3.075 $X2=0 $Y2=0
cc_923 N_A_1098_271#_c_1150_n N_A_1982_397#_c_1375_n 0.00262513f $X=16.105
+ $Y=1.025 $X2=0 $Y2=0
cc_924 N_A_1098_271#_c_1154_n N_A_1982_397#_c_1375_n 0.00520485f $X=16.76
+ $Y=1.205 $X2=0 $Y2=0
cc_925 N_A_1098_271#_c_1150_n N_A_1982_397#_c_1376_n 0.00587859f $X=16.105
+ $Y=1.025 $X2=0 $Y2=0
cc_926 N_A_1098_271#_c_1154_n N_A_1982_397#_c_1376_n 0.0179175f $X=16.76
+ $Y=1.205 $X2=0 $Y2=0
cc_927 N_A_1098_271#_c_1149_n N_A_2586_249#_c_1569_n 0.00366812f $X=14.44
+ $Y=1.67 $X2=0 $Y2=0
cc_928 N_A_1098_271#_c_1150_n N_A_2586_249#_c_1569_n 0.0132208f $X=16.105
+ $Y=1.025 $X2=0 $Y2=0
cc_929 N_A_1098_271#_c_1176_n N_A_2586_249#_c_1570_n 0.0951188f $X=14.355
+ $Y=1.755 $X2=0 $Y2=0
cc_930 N_A_1098_271#_c_1149_n N_A_2586_249#_c_1570_n 0.0152006f $X=14.44 $Y=1.67
+ $X2=0 $Y2=0
cc_931 N_A_1098_271#_c_1176_n N_A_2586_249#_c_1571_n 0.00872625f $X=14.355
+ $Y=1.755 $X2=0 $Y2=0
cc_932 N_A_1098_271#_c_1149_n N_A_2586_249#_c_1572_n 0.0157375f $X=14.44 $Y=1.67
+ $X2=0 $Y2=0
cc_933 N_A_1098_271#_c_1151_n N_A_2586_249#_c_1572_n 0.0143583f $X=14.525
+ $Y=1.025 $X2=0 $Y2=0
cc_934 N_A_1098_271#_c_1150_n N_A_2586_249#_c_1573_n 0.0345629f $X=16.105
+ $Y=1.025 $X2=0 $Y2=0
cc_935 N_A_1098_271#_c_1151_n N_A_2586_249#_c_1573_n 0.0143582f $X=14.525
+ $Y=1.025 $X2=0 $Y2=0
cc_936 N_A_1098_271#_c_1150_n N_A_2586_249#_c_1575_n 0.0251543f $X=16.105
+ $Y=1.025 $X2=0 $Y2=0
cc_937 N_A_1098_271#_c_1150_n N_A_2586_249#_c_1576_n 0.0264495f $X=16.105
+ $Y=1.025 $X2=0 $Y2=0
cc_938 N_A_1098_271#_c_1152_n N_A_2586_249#_c_1576_n 0.0249405f $X=16.27 $Y=0.76
+ $X2=0 $Y2=0
cc_939 N_A_1098_271#_c_1154_n N_A_2586_249#_c_1576_n 0.0103903f $X=16.76
+ $Y=1.205 $X2=0 $Y2=0
cc_940 N_A_1098_271#_c_1152_n N_A_2586_249#_c_1578_n 0.00595662f $X=16.27
+ $Y=0.76 $X2=0 $Y2=0
cc_941 N_A_1098_271#_c_1153_n N_A_2586_249#_c_1579_n 0.0295015f $X=17.325
+ $Y=1.205 $X2=0 $Y2=0
cc_942 N_A_1098_271#_c_1152_n N_A_2586_249#_c_1580_n 0.00574702f $X=16.27
+ $Y=0.76 $X2=0 $Y2=0
cc_943 N_A_1098_271#_c_1153_n N_A_2586_249#_c_1580_n 0.0132688f $X=17.325
+ $Y=1.205 $X2=0 $Y2=0
cc_944 N_A_1098_271#_c_1154_n N_A_2586_249#_c_1580_n 3.96313e-19 $X=16.76
+ $Y=1.205 $X2=0 $Y2=0
cc_945 N_A_1098_271#_c_1153_n N_A_2586_249#_c_1581_n 0.00792984f $X=17.325
+ $Y=1.205 $X2=0 $Y2=0
cc_946 N_A_1098_271#_c_1155_n N_A_2586_249#_c_1581_n 0.0205765f $X=17.41 $Y=2.01
+ $X2=0 $Y2=0
cc_947 N_A_1098_271#_c_1150_n N_A_2586_249#_c_1583_n 0.00415365f $X=16.105
+ $Y=1.025 $X2=0 $Y2=0
cc_948 N_A_1098_271#_c_1280_p N_A_2586_249#_c_1588_n 0.00749913f $X=17.325
+ $Y=2.095 $X2=0 $Y2=0
cc_949 N_A_1098_271#_c_1155_n N_A_2586_249#_c_1588_n 0.00649223f $X=17.41
+ $Y=2.01 $X2=0 $Y2=0
cc_950 N_A_1098_271#_c_1144_n N_RESET_B_c_1722_n 0.0031339f $X=5.675 $Y=1.355
+ $X2=0 $Y2=0
cc_951 N_A_1098_271#_c_1159_n N_RESET_B_M1043_g 0.00444656f $X=8.27 $Y=3.15
+ $X2=0 $Y2=0
cc_952 N_A_1098_271#_M1029_g N_RESET_B_c_1726_n 0.00495681f $X=8.505 $Y=1.025
+ $X2=0 $Y2=0
cc_953 N_A_1098_271#_M1018_g N_RESET_B_c_1726_n 0.00737233f $X=10.595 $Y=0.835
+ $X2=0 $Y2=0
cc_954 N_A_1098_271#_c_1150_n N_RESET_B_c_1729_n 0.0107342f $X=16.105 $Y=1.025
+ $X2=0 $Y2=0
cc_955 N_A_1098_271#_c_1154_n N_RESET_B_c_1729_n 3.59908e-19 $X=16.76 $Y=1.205
+ $X2=0 $Y2=0
cc_956 N_A_1098_271#_c_1150_n N_RESET_B_c_1734_n 0.00850394f $X=16.105 $Y=1.025
+ $X2=0 $Y2=0
cc_957 N_A_1098_271#_c_1152_n N_RESET_B_c_1734_n 0.010775f $X=16.27 $Y=0.76
+ $X2=0 $Y2=0
cc_958 N_A_1098_271#_c_1152_n N_CLK_M1048_g 0.00897709f $X=16.27 $Y=0.76 $X2=0
+ $Y2=0
cc_959 N_A_1098_271#_c_1154_n N_CLK_M1048_g 0.0266757f $X=16.76 $Y=1.205 $X2=0
+ $Y2=0
cc_960 N_A_1098_271#_c_1155_n N_CLK_M1048_g 6.64745e-19 $X=17.41 $Y=2.01 $X2=0
+ $Y2=0
cc_961 N_A_1098_271#_c_1153_n CLK 0.030618f $X=17.325 $Y=1.205 $X2=0 $Y2=0
cc_962 N_A_1098_271#_c_1154_n CLK 0.0132027f $X=16.76 $Y=1.205 $X2=0 $Y2=0
cc_963 N_A_1098_271#_c_1280_p CLK 0.0160371f $X=17.325 $Y=2.095 $X2=0 $Y2=0
cc_964 N_A_1098_271#_c_1155_n CLK 0.0272626f $X=17.41 $Y=2.01 $X2=0 $Y2=0
cc_965 N_A_1098_271#_c_1153_n N_CLK_c_1889_n 0.00337834f $X=17.325 $Y=1.205
+ $X2=0 $Y2=0
cc_966 N_A_1098_271#_c_1154_n N_CLK_c_1889_n 0.00217604f $X=16.76 $Y=1.205 $X2=0
+ $Y2=0
cc_967 N_A_1098_271#_c_1280_p N_CLK_c_1889_n 0.00127863f $X=17.325 $Y=2.095
+ $X2=0 $Y2=0
cc_968 N_A_1098_271#_c_1154_n N_SLEEP_B_c_1931_n 0.00488514f $X=16.76 $Y=1.205
+ $X2=-0.19 $Y2=-0.245
cc_969 N_A_1098_271#_c_1280_p N_SLEEP_B_M1027_g 0.0130773f $X=17.325 $Y=2.095
+ $X2=0 $Y2=0
cc_970 N_A_1098_271#_c_1155_n N_SLEEP_B_M1027_g 0.00871623f $X=17.41 $Y=2.01
+ $X2=0 $Y2=0
cc_971 N_A_1098_271#_c_1155_n N_SLEEP_B_c_1934_n 0.00862258f $X=17.41 $Y=2.01
+ $X2=0 $Y2=0
cc_972 N_A_1098_271#_c_1153_n N_SLEEP_B_c_1935_n 0.029926f $X=17.325 $Y=1.205
+ $X2=0 $Y2=0
cc_973 N_A_1098_271#_c_1155_n N_SLEEP_B_c_1935_n 0.00412588f $X=17.41 $Y=2.01
+ $X2=0 $Y2=0
cc_974 N_A_1098_271#_c_1280_p N_SLEEP_B_M1025_g 0.00163399f $X=17.325 $Y=2.095
+ $X2=0 $Y2=0
cc_975 N_A_1098_271#_c_1155_n N_SLEEP_B_c_1940_n 0.00449563f $X=17.41 $Y=2.01
+ $X2=0 $Y2=0
cc_976 N_A_1098_271#_M1004_g N_VPWR_c_2096_n 0.00633492f $X=5.565 $Y=2.33 $X2=0
+ $Y2=0
cc_977 N_A_1098_271#_c_1159_n N_VPWR_c_2096_n 0.0247934f $X=8.27 $Y=3.15 $X2=0
+ $Y2=0
cc_978 N_A_1098_271#_c_1159_n N_VPWR_c_2097_n 0.0255538f $X=8.27 $Y=3.15 $X2=0
+ $Y2=0
cc_979 N_A_1098_271#_M1013_g N_VPWR_c_2097_n 0.00737681f $X=8.345 $Y=2.485 $X2=0
+ $Y2=0
cc_980 N_A_1098_271#_c_1160_n N_VPWR_c_2101_n 0.0161929f $X=5.64 $Y=3.15 $X2=0
+ $Y2=0
cc_981 N_A_1098_271#_c_1159_n N_VPWR_c_2103_n 0.0808488f $X=8.27 $Y=3.15 $X2=0
+ $Y2=0
cc_982 N_A_1098_271#_c_1159_n N_VPWR_c_2106_n 0.0373685f $X=8.27 $Y=3.15 $X2=0
+ $Y2=0
cc_983 N_A_1098_271#_c_1159_n N_VPWR_c_2093_n 0.0361698f $X=8.27 $Y=3.15 $X2=0
+ $Y2=0
cc_984 N_A_1098_271#_c_1160_n N_VPWR_c_2093_n 0.00559617f $X=5.64 $Y=3.15 $X2=0
+ $Y2=0
cc_985 N_A_1098_271#_c_1162_n N_VPWR_c_2093_n 0.0320636f $X=10.195 $Y=3.15 $X2=0
+ $Y2=0
cc_986 N_A_1098_271#_c_1166_n N_VPWR_c_2093_n 0.00421462f $X=10.555 $Y=3.15
+ $X2=0 $Y2=0
cc_987 N_A_1098_271#_c_1169_n N_VPWR_c_2093_n 0.0225254f $X=11.64 $Y=3.15 $X2=0
+ $Y2=0
cc_988 N_A_1098_271#_c_1172_n N_VPWR_c_2093_n 0.00357864f $X=8.345 $Y=3.15 $X2=0
+ $Y2=0
cc_989 N_A_1098_271#_c_1173_n N_VPWR_c_2093_n 0.00310744f $X=10.27 $Y=3.15 $X2=0
+ $Y2=0
cc_990 N_A_1098_271#_c_1175_n N_VPWR_c_2093_n 0.00310744f $X=10.63 $Y=3.15 $X2=0
+ $Y2=0
cc_991 N_A_1098_271#_c_1144_n N_A_332_136#_c_2245_n 6.05373e-19 $X=5.675
+ $Y=1.355 $X2=0 $Y2=0
cc_992 N_A_1098_271#_c_1144_n N_A_332_136#_c_2246_n 0.0102108f $X=5.675 $Y=1.355
+ $X2=0 $Y2=0
cc_993 N_A_1098_271#_c_1147_n N_A_332_136#_c_2246_n 0.00142225f $X=5.675 $Y=1.43
+ $X2=0 $Y2=0
cc_994 N_A_1098_271#_c_1144_n N_A_332_136#_c_2248_n 0.00948707f $X=5.675
+ $Y=1.355 $X2=0 $Y2=0
cc_995 N_A_1098_271#_c_1280_p N_KAPWR_M1027_d 0.00365987f $X=17.325 $Y=2.095
+ $X2=0 $Y2=0
cc_996 N_A_1098_271#_c_1155_n N_KAPWR_M1027_d 7.52847e-19 $X=17.41 $Y=2.01 $X2=0
+ $Y2=0
cc_997 N_A_1098_271#_M1004_g N_KAPWR_c_2381_n 0.00706328f $X=5.565 $Y=2.33 $X2=0
+ $Y2=0
cc_998 N_A_1098_271#_c_1159_n N_KAPWR_c_2381_n 0.0185096f $X=8.27 $Y=3.15 $X2=0
+ $Y2=0
cc_999 N_A_1098_271#_M1013_g N_KAPWR_c_2381_n 0.00769535f $X=8.345 $Y=2.485
+ $X2=0 $Y2=0
cc_1000 N_A_1098_271#_c_1162_n N_KAPWR_c_2381_n 5.57362e-19 $X=10.195 $Y=3.15
+ $X2=0 $Y2=0
cc_1001 N_A_1098_271#_M1037_g N_KAPWR_c_2381_n 0.00305687f $X=10.27 $Y=2.405
+ $X2=0 $Y2=0
cc_1002 N_A_1098_271#_M1038_g N_KAPWR_c_2381_n 0.00352427f $X=10.63 $Y=2.405
+ $X2=0 $Y2=0
cc_1003 N_A_1098_271#_c_1170_n N_KAPWR_c_2381_n 0.00554431f $X=11.715 $Y=3.075
+ $X2=0 $Y2=0
cc_1004 N_A_1098_271#_M1029_g N_VGND_c_2528_n 0.00385594f $X=8.505 $Y=1.025
+ $X2=0 $Y2=0
cc_1005 N_A_1098_271#_M1029_g N_VGND_c_2548_n 9.72468e-19 $X=8.505 $Y=1.025
+ $X2=0 $Y2=0
cc_1006 N_A_1098_271#_c_1144_n N_A_929_152#_c_2756_n 4.20626e-19 $X=5.675
+ $Y=1.355 $X2=0 $Y2=0
cc_1007 N_A_1098_271#_c_1144_n N_A_929_152#_c_2758_n 5.56636e-19 $X=5.675
+ $Y=1.355 $X2=0 $Y2=0
cc_1008 N_A_1098_271#_c_1176_n N_A_2544_119#_c_2793_n 0.00879467f $X=14.355
+ $Y=1.755 $X2=0 $Y2=0
cc_1009 N_A_1982_397#_c_1388_n N_A_2586_249#_M1025_d 0.0100859f $X=19.155
+ $Y=2.435 $X2=0 $Y2=0
cc_1010 N_A_1982_397#_M1044_g N_A_2586_249#_M1047_g 0.0179736f $X=12.645
+ $Y=0.805 $X2=0 $Y2=0
cc_1011 N_A_1982_397#_c_1408_n N_A_2586_249#_c_1585_n 0.0225488f $X=16.25
+ $Y=2.435 $X2=0 $Y2=0
cc_1012 N_A_1982_397#_M1044_g N_A_2586_249#_c_1570_n 0.00117485f $X=12.645
+ $Y=0.805 $X2=0 $Y2=0
cc_1013 N_A_1982_397#_M1044_g N_A_2586_249#_c_1571_n 0.021096f $X=12.645
+ $Y=0.805 $X2=0 $Y2=0
cc_1014 N_A_1982_397#_c_1388_n N_A_2586_249#_c_1588_n 0.0387361f $X=19.155
+ $Y=2.435 $X2=0 $Y2=0
cc_1015 N_A_1982_397#_M1006_g N_RESET_B_c_1726_n 0.0103003f $X=12.285 $Y=0.805
+ $X2=0 $Y2=0
cc_1016 N_A_1982_397#_M1044_g N_RESET_B_c_1726_n 0.0103003f $X=12.645 $Y=0.805
+ $X2=0 $Y2=0
cc_1017 N_A_1982_397#_M1015_g N_RESET_B_M1041_g 0.0493387f $X=16.18 $Y=2.45
+ $X2=0 $Y2=0
cc_1018 N_A_1982_397#_c_1408_n N_RESET_B_M1041_g 0.0181948f $X=16.25 $Y=2.435
+ $X2=0 $Y2=0
cc_1019 N_A_1982_397#_c_1387_n N_RESET_B_M1041_g 7.84738e-19 $X=16.335 $Y=2.35
+ $X2=0 $Y2=0
cc_1020 N_A_1982_397#_c_1375_n N_RESET_B_M1041_g 0.0213004f $X=16.15 $Y=1.575
+ $X2=0 $Y2=0
cc_1021 N_A_1982_397#_c_1376_n N_RESET_B_M1041_g 5.48664e-19 $X=16.335 $Y=1.575
+ $X2=0 $Y2=0
cc_1022 N_A_1982_397#_c_1375_n N_CLK_M1048_g 0.0205145f $X=16.15 $Y=1.575 $X2=0
+ $Y2=0
cc_1023 N_A_1982_397#_c_1376_n N_CLK_M1048_g 0.00317733f $X=16.335 $Y=1.575
+ $X2=0 $Y2=0
cc_1024 N_A_1982_397#_M1015_g N_CLK_M1024_g 0.0243962f $X=16.18 $Y=2.45 $X2=0
+ $Y2=0
cc_1025 N_A_1982_397#_c_1387_n N_CLK_M1024_g 0.00877002f $X=16.335 $Y=2.35 $X2=0
+ $Y2=0
cc_1026 N_A_1982_397#_c_1388_n N_CLK_M1024_g 0.0130374f $X=19.155 $Y=2.435 $X2=0
+ $Y2=0
cc_1027 N_A_1982_397#_c_1387_n CLK 0.00385819f $X=16.335 $Y=2.35 $X2=0 $Y2=0
cc_1028 N_A_1982_397#_c_1388_n CLK 0.00643086f $X=19.155 $Y=2.435 $X2=0 $Y2=0
cc_1029 N_A_1982_397#_c_1375_n CLK 2.52952e-19 $X=16.15 $Y=1.575 $X2=0 $Y2=0
cc_1030 N_A_1982_397#_c_1376_n CLK 0.0236101f $X=16.335 $Y=1.575 $X2=0 $Y2=0
cc_1031 N_A_1982_397#_M1015_g N_CLK_c_1889_n 0.00292332f $X=16.18 $Y=2.45 $X2=0
+ $Y2=0
cc_1032 N_A_1982_397#_c_1387_n N_CLK_c_1889_n 3.31341e-19 $X=16.335 $Y=2.35
+ $X2=0 $Y2=0
cc_1033 N_A_1982_397#_c_1388_n N_CLK_c_1889_n 0.00375054f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1034 N_A_1982_397#_c_1388_n N_SLEEP_B_M1027_g 0.011591f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1035 N_A_1982_397#_c_1388_n N_SLEEP_B_M1025_g 0.0204954f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1036 N_A_1982_397#_M1031_g N_SLEEP_B_M1014_g 0.0197472f $X=19.185 $Y=0.575
+ $X2=0 $Y2=0
cc_1037 N_A_1982_397#_M1031_g N_SLEEP_B_c_1942_n 0.00362793f $X=19.185 $Y=0.575
+ $X2=0 $Y2=0
cc_1038 N_A_1982_397#_c_1378_n N_SLEEP_B_c_1942_n 0.00267244f $X=19.21 $Y=1.48
+ $X2=0 $Y2=0
cc_1039 N_A_1982_397#_c_1388_n N_A_3751_367#_M1051_s 0.00314434f $X=19.155
+ $Y=2.435 $X2=0 $Y2=0
cc_1040 N_A_1982_397#_M1051_g N_A_3751_367#_M1016_g 0.00928924f $X=19.115
+ $Y=2.155 $X2=0 $Y2=0
cc_1041 N_A_1982_397#_c_1389_n N_A_3751_367#_M1016_g 0.00319648f $X=19.24
+ $Y=2.35 $X2=0 $Y2=0
cc_1042 N_A_1982_397#_M1031_g N_A_3751_367#_c_2023_n 0.011413f $X=19.185
+ $Y=0.575 $X2=0 $Y2=0
cc_1043 N_A_1982_397#_c_1377_n N_A_3751_367#_c_2023_n 0.0118583f $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1044 N_A_1982_397#_c_1378_n N_A_3751_367#_c_2023_n 0.0017307f $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1045 N_A_1982_397#_M1031_g N_A_3751_367#_c_2025_n 0.0134005f $X=19.185
+ $Y=0.575 $X2=0 $Y2=0
cc_1046 N_A_1982_397#_M1031_g N_A_3751_367#_c_2026_n 0.00356655f $X=19.185
+ $Y=0.575 $X2=0 $Y2=0
cc_1047 N_A_1982_397#_M1051_g N_A_3751_367#_c_2032_n 4.40799e-19 $X=19.115
+ $Y=2.155 $X2=0 $Y2=0
cc_1048 N_A_1982_397#_c_1388_n N_A_3751_367#_c_2032_n 0.0190759f $X=19.155
+ $Y=2.435 $X2=0 $Y2=0
cc_1049 N_A_1982_397#_c_1389_n N_A_3751_367#_c_2032_n 0.0131279f $X=19.24
+ $Y=2.35 $X2=0 $Y2=0
cc_1050 N_A_1982_397#_M1031_g N_A_3751_367#_c_2027_n 0.00198316f $X=19.185
+ $Y=0.575 $X2=0 $Y2=0
cc_1051 N_A_1982_397#_c_1389_n N_A_3751_367#_c_2027_n 0.00906598f $X=19.24
+ $Y=2.35 $X2=0 $Y2=0
cc_1052 N_A_1982_397#_c_1377_n N_A_3751_367#_c_2027_n 0.0244257f $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1053 N_A_1982_397#_c_1378_n N_A_3751_367#_c_2027_n 0.00933109f $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1054 N_A_1982_397#_M1031_g N_A_3751_367#_c_2028_n 0.00446384f $X=19.185
+ $Y=0.575 $X2=0 $Y2=0
cc_1055 N_A_1982_397#_c_1377_n N_A_3751_367#_c_2028_n 0.00952147f $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1056 N_A_1982_397#_c_1378_n N_A_3751_367#_c_2028_n 0.00204252f $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1057 N_A_1982_397#_c_1377_n N_A_3751_367#_c_2029_n 0.0266166f $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1058 N_A_1982_397#_c_1378_n N_A_3751_367#_c_2029_n 0.00253121f $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1059 N_A_1982_397#_c_1377_n N_A_3751_367#_c_2030_n 3.00671e-19 $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1060 N_A_1982_397#_c_1378_n N_A_3751_367#_c_2030_n 0.0120985f $X=19.21
+ $Y=1.48 $X2=0 $Y2=0
cc_1061 N_A_1982_397#_c_1388_n N_VPWR_M1051_d 0.00124906f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1062 N_A_1982_397#_c_1389_n N_VPWR_M1051_d 0.00492477f $X=19.24 $Y=2.35 $X2=0
+ $Y2=0
cc_1063 N_A_1982_397#_M1051_g N_VPWR_c_2098_n 0.00425371f $X=19.115 $Y=2.155
+ $X2=0 $Y2=0
cc_1064 N_A_1982_397#_c_1388_n N_VPWR_c_2098_n 0.0146259f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1065 N_A_1982_397#_c_1389_n N_VPWR_c_2098_n 0.0409063f $X=19.24 $Y=2.35 $X2=0
+ $Y2=0
cc_1066 N_A_1982_397#_M1015_g N_VPWR_c_2103_n 0.00923926f $X=16.18 $Y=2.45 $X2=0
+ $Y2=0
cc_1067 N_A_1982_397#_M1051_g N_VPWR_c_2103_n 0.00312414f $X=19.115 $Y=2.155
+ $X2=0 $Y2=0
cc_1068 N_A_1982_397#_c_1386_n N_VPWR_c_2103_n 0.013898f $X=13.79 $Y=2.66 $X2=0
+ $Y2=0
cc_1069 N_A_1982_397#_M1015_g N_VPWR_c_2093_n 0.00531456f $X=16.18 $Y=2.45 $X2=0
+ $Y2=0
cc_1070 N_A_1982_397#_c_1386_n N_VPWR_c_2093_n 0.00304108f $X=13.79 $Y=2.66
+ $X2=0 $Y2=0
cc_1071 N_A_1982_397#_c_1390_n A_2069_397# 4.54001e-19 $X=10.055 $Y=2.13
+ $X2=-0.19 $Y2=-0.245
cc_1072 N_A_1982_397#_c_1408_n A_2836_390# 0.00295351f $X=16.25 $Y=2.435
+ $X2=-0.19 $Y2=-0.245
cc_1073 N_A_1982_397#_c_1408_n N_KAPWR_M1022_d 0.00757154f $X=16.25 $Y=2.435
+ $X2=-0.19 $Y2=-0.245
cc_1074 N_A_1982_397#_c_1387_n N_KAPWR_M1015_d 0.00509849f $X=16.335 $Y=2.35
+ $X2=0 $Y2=0
cc_1075 N_A_1982_397#_c_1388_n N_KAPWR_M1015_d 0.008356f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1076 N_A_1982_397#_c_1536_p N_KAPWR_M1015_d 5.71553e-19 $X=16.335 $Y=2.435
+ $X2=0 $Y2=0
cc_1077 N_A_1982_397#_c_1388_n N_KAPWR_M1027_d 0.0168891f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1078 N_A_1982_397#_c_1386_n N_KAPWR_c_2379_n 0.00374751f $X=13.79 $Y=2.66
+ $X2=0 $Y2=0
cc_1079 N_A_1982_397#_c_1408_n N_KAPWR_c_2379_n 0.025597f $X=16.25 $Y=2.435
+ $X2=0 $Y2=0
cc_1080 N_A_1982_397#_M1015_g N_KAPWR_c_2380_n 0.00715744f $X=16.18 $Y=2.45
+ $X2=0 $Y2=0
cc_1081 N_A_1982_397#_c_1388_n N_KAPWR_c_2380_n 0.0154471f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1082 N_A_1982_397#_c_1536_p N_KAPWR_c_2380_n 0.00681059f $X=16.335 $Y=2.435
+ $X2=0 $Y2=0
cc_1083 N_A_1982_397#_M1015_g N_KAPWR_c_2381_n 0.00630248f $X=16.18 $Y=2.45
+ $X2=0 $Y2=0
cc_1084 N_A_1982_397#_M1051_g N_KAPWR_c_2381_n 0.00480838f $X=19.115 $Y=2.155
+ $X2=0 $Y2=0
cc_1085 N_A_1982_397#_c_1384_n N_KAPWR_c_2381_n 0.0663534f $X=12.21 $Y=2.65
+ $X2=0 $Y2=0
cc_1086 N_A_1982_397#_c_1385_n N_KAPWR_c_2381_n 0.036846f $X=13.625 $Y=2.435
+ $X2=0 $Y2=0
cc_1087 N_A_1982_397#_c_1386_n N_KAPWR_c_2381_n 0.0278749f $X=13.79 $Y=2.66
+ $X2=0 $Y2=0
cc_1088 N_A_1982_397#_c_1408_n N_KAPWR_c_2381_n 0.0951609f $X=16.25 $Y=2.435
+ $X2=0 $Y2=0
cc_1089 N_A_1982_397#_c_1388_n N_KAPWR_c_2381_n 0.118149f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1090 N_A_1982_397#_c_1390_n N_KAPWR_c_2381_n 0.0461448f $X=10.055 $Y=2.13
+ $X2=0 $Y2=0
cc_1091 N_A_1982_397#_c_1391_n N_KAPWR_c_2381_n 0.0134907f $X=12.375 $Y=2.435
+ $X2=0 $Y2=0
cc_1092 N_A_1982_397#_c_1536_p N_KAPWR_c_2381_n 0.00542768f $X=16.335 $Y=2.435
+ $X2=0 $Y2=0
cc_1093 N_A_1982_397#_M1015_g N_KAPWR_c_2382_n 0.00178545f $X=16.18 $Y=2.45
+ $X2=0 $Y2=0
cc_1094 N_A_1982_397#_c_1388_n N_KAPWR_c_2382_n 0.0480512f $X=19.155 $Y=2.435
+ $X2=0 $Y2=0
cc_1095 N_A_1982_397#_c_1408_n A_3063_390# 0.00489024f $X=16.25 $Y=2.435
+ $X2=-0.19 $Y2=-0.245
cc_1096 N_A_1982_397#_M1006_g N_VGND_c_2529_n 0.00359922f $X=12.285 $Y=0.805
+ $X2=0 $Y2=0
cc_1097 N_A_1982_397#_M1044_g N_VGND_c_2530_n 6.2241e-19 $X=12.645 $Y=0.805
+ $X2=0 $Y2=0
cc_1098 N_A_1982_397#_M1031_g N_VGND_c_2532_n 0.00319684f $X=19.185 $Y=0.575
+ $X2=0 $Y2=0
cc_1099 N_A_1982_397#_M1031_g N_VGND_c_2533_n 0.00438034f $X=19.185 $Y=0.575
+ $X2=0 $Y2=0
cc_1100 N_A_1982_397#_M1031_g N_VGND_c_2534_n 0.00396391f $X=19.185 $Y=0.575
+ $X2=0 $Y2=0
cc_1101 N_A_1982_397#_M1006_g N_VGND_c_2548_n 9.39239e-19 $X=12.285 $Y=0.805
+ $X2=0 $Y2=0
cc_1102 N_A_1982_397#_M1044_g N_VGND_c_2548_n 9.39239e-19 $X=12.645 $Y=0.805
+ $X2=0 $Y2=0
cc_1103 N_A_1982_397#_M1031_g N_VGND_c_2548_n 0.00838463f $X=19.185 $Y=0.575
+ $X2=0 $Y2=0
cc_1104 N_A_1982_397#_M1006_g N_A_2544_119#_c_2791_n 0.00110389f $X=12.285
+ $Y=0.805 $X2=0 $Y2=0
cc_1105 N_A_1982_397#_M1044_g N_A_2544_119#_c_2791_n 0.00706674f $X=12.645
+ $Y=0.805 $X2=0 $Y2=0
cc_1106 N_A_1982_397#_M1006_g N_A_2544_119#_c_2793_n 4.60652e-19 $X=12.285
+ $Y=0.805 $X2=0 $Y2=0
cc_1107 N_A_1982_397#_M1044_g N_A_2544_119#_c_2793_n 0.00512038f $X=12.645
+ $Y=0.805 $X2=0 $Y2=0
cc_1108 N_A_2586_249#_M1047_g N_RESET_B_c_1726_n 0.0103107f $X=13.075 $Y=0.805
+ $X2=0 $Y2=0
cc_1109 N_A_2586_249#_M1047_g N_RESET_B_M1007_g 0.0127349f $X=13.075 $Y=0.805
+ $X2=0 $Y2=0
cc_1110 N_A_2586_249#_c_1570_n N_RESET_B_M1007_g 0.00103411f $X=14.015 $Y=1.41
+ $X2=0 $Y2=0
cc_1111 N_A_2586_249#_c_1572_n N_RESET_B_M1007_g 6.4344e-19 $X=14.1 $Y=1.32
+ $X2=0 $Y2=0
cc_1112 N_A_2586_249#_c_1573_n N_RESET_B_c_1728_n 0.0145904f $X=14.985 $Y=0.685
+ $X2=0 $Y2=0
cc_1113 N_A_2586_249#_c_1574_n N_RESET_B_c_1728_n 0.0033875f $X=14.185 $Y=0.685
+ $X2=0 $Y2=0
cc_1114 N_A_2586_249#_c_1576_n N_RESET_B_c_1728_n 0.00516323f $X=16.93 $Y=0.34
+ $X2=0 $Y2=0
cc_1115 N_A_2586_249#_c_1577_n N_RESET_B_c_1728_n 0.00253817f $X=15.315 $Y=0.34
+ $X2=0 $Y2=0
cc_1116 N_A_2586_249#_c_1583_n N_RESET_B_c_1728_n 0.0213759f $X=15.15 $Y=0.63
+ $X2=0 $Y2=0
cc_1117 N_A_2586_249#_c_1569_n N_RESET_B_c_1729_n 0.0681173f $X=15.19 $Y=1.82
+ $X2=0 $Y2=0
cc_1118 N_A_2586_249#_c_1576_n N_RESET_B_c_1729_n 4.57988e-19 $X=16.93 $Y=0.34
+ $X2=0 $Y2=0
cc_1119 N_A_2586_249#_c_1585_n N_RESET_B_M1041_g 0.0681173f $X=15.19 $Y=1.945
+ $X2=0 $Y2=0
cc_1120 N_A_2586_249#_c_1575_n N_RESET_B_c_1734_n 0.00311641f $X=15.15 $Y=0.6
+ $X2=0 $Y2=0
cc_1121 N_A_2586_249#_c_1576_n N_RESET_B_c_1734_n 0.015435f $X=16.93 $Y=0.34
+ $X2=0 $Y2=0
cc_1122 N_A_2586_249#_c_1583_n N_RESET_B_c_1734_n 0.0236901f $X=15.15 $Y=0.63
+ $X2=0 $Y2=0
cc_1123 N_A_2586_249#_c_1576_n N_CLK_M1048_g 0.00949795f $X=16.93 $Y=0.34 $X2=0
+ $Y2=0
cc_1124 N_A_2586_249#_c_1578_n N_CLK_M1048_g 0.00164034f $X=17.015 $Y=0.78 $X2=0
+ $Y2=0
cc_1125 N_A_2586_249#_c_1580_n N_CLK_M1048_g 5.63197e-19 $X=17.1 $Y=0.865 $X2=0
+ $Y2=0
cc_1126 N_A_2586_249#_c_1576_n N_SLEEP_B_c_1931_n 0.00619259f $X=16.93 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_1127 N_A_2586_249#_c_1578_n N_SLEEP_B_c_1931_n 0.00899233f $X=17.015 $Y=0.78
+ $X2=-0.19 $Y2=-0.245
cc_1128 N_A_2586_249#_c_1580_n N_SLEEP_B_c_1931_n 0.00680982f $X=17.1 $Y=0.865
+ $X2=-0.19 $Y2=-0.245
cc_1129 N_A_2586_249#_c_1588_n N_SLEEP_B_M1027_g 2.15381e-19 $X=18.325 $Y=2.015
+ $X2=0 $Y2=0
cc_1130 N_A_2586_249#_c_1576_n N_SLEEP_B_c_1933_n 6.45019e-19 $X=16.93 $Y=0.34
+ $X2=0 $Y2=0
cc_1131 N_A_2586_249#_c_1578_n N_SLEEP_B_c_1933_n 0.00482976f $X=17.015 $Y=0.78
+ $X2=0 $Y2=0
cc_1132 N_A_2586_249#_c_1579_n N_SLEEP_B_c_1933_n 0.0131919f $X=17.895 $Y=0.865
+ $X2=0 $Y2=0
cc_1133 N_A_2586_249#_c_1581_n N_SLEEP_B_c_1933_n 0.0044978f $X=17.98 $Y=1.85
+ $X2=0 $Y2=0
cc_1134 N_A_2586_249#_c_1582_n N_SLEEP_B_c_1933_n 0.00429736f $X=18.18 $Y=0.575
+ $X2=0 $Y2=0
cc_1135 N_A_2586_249#_c_1579_n N_SLEEP_B_c_1934_n 0.0127365f $X=17.895 $Y=0.865
+ $X2=0 $Y2=0
cc_1136 N_A_2586_249#_c_1579_n N_SLEEP_B_c_1935_n 6.49981e-19 $X=17.895 $Y=0.865
+ $X2=0 $Y2=0
cc_1137 N_A_2586_249#_c_1581_n N_SLEEP_B_c_1935_n 8.91232e-19 $X=17.98 $Y=1.85
+ $X2=0 $Y2=0
cc_1138 N_A_2586_249#_c_1581_n N_SLEEP_B_c_1944_n 0.00660493f $X=17.98 $Y=1.85
+ $X2=0 $Y2=0
cc_1139 N_A_2586_249#_c_1581_n N_SLEEP_B_M1025_g 0.00206039f $X=17.98 $Y=1.85
+ $X2=0 $Y2=0
cc_1140 N_A_2586_249#_c_1588_n N_SLEEP_B_M1025_g 0.0195752f $X=18.325 $Y=2.015
+ $X2=0 $Y2=0
cc_1141 N_A_2586_249#_c_1581_n N_SLEEP_B_c_1936_n 0.00649257f $X=17.98 $Y=1.85
+ $X2=0 $Y2=0
cc_1142 N_A_2586_249#_c_1584_n N_SLEEP_B_c_1936_n 0.0056244f $X=18.12 $Y=0.865
+ $X2=0 $Y2=0
cc_1143 N_A_2586_249#_c_1588_n N_SLEEP_B_c_1936_n 0.0103366f $X=18.325 $Y=2.015
+ $X2=0 $Y2=0
cc_1144 N_A_2586_249#_c_1582_n N_SLEEP_B_M1012_g 0.00803496f $X=18.18 $Y=0.575
+ $X2=0 $Y2=0
cc_1145 N_A_2586_249#_c_1584_n N_SLEEP_B_M1012_g 0.00610785f $X=18.12 $Y=0.865
+ $X2=0 $Y2=0
cc_1146 N_A_2586_249#_c_1582_n N_SLEEP_B_M1014_g 0.00118315f $X=18.18 $Y=0.575
+ $X2=0 $Y2=0
cc_1147 N_A_2586_249#_c_1584_n N_SLEEP_B_M1014_g 6.58536e-19 $X=18.12 $Y=0.865
+ $X2=0 $Y2=0
cc_1148 N_A_2586_249#_c_1581_n N_SLEEP_B_c_1939_n 0.0060075f $X=17.98 $Y=1.85
+ $X2=0 $Y2=0
cc_1149 N_A_2586_249#_c_1581_n N_SLEEP_B_c_1940_n 0.00841211f $X=17.98 $Y=1.85
+ $X2=0 $Y2=0
cc_1150 N_A_2586_249#_c_1581_n SLEEP_B 0.0242156f $X=17.98 $Y=1.85 $X2=0 $Y2=0
cc_1151 N_A_2586_249#_c_1584_n SLEEP_B 0.00907709f $X=18.12 $Y=0.865 $X2=0 $Y2=0
cc_1152 N_A_2586_249#_c_1588_n SLEEP_B 0.0106755f $X=18.325 $Y=2.015 $X2=0 $Y2=0
cc_1153 N_A_2586_249#_c_1581_n N_SLEEP_B_c_1942_n 0.00585222f $X=17.98 $Y=1.85
+ $X2=0 $Y2=0
cc_1154 N_A_2586_249#_c_1584_n N_SLEEP_B_c_1942_n 0.00421488f $X=18.12 $Y=0.865
+ $X2=0 $Y2=0
cc_1155 N_A_2586_249#_c_1581_n N_A_3751_367#_c_2024_n 0.00422769f $X=17.98
+ $Y=1.85 $X2=0 $Y2=0
cc_1156 N_A_2586_249#_c_1588_n N_A_3751_367#_c_2032_n 0.0217869f $X=18.325
+ $Y=2.015 $X2=0 $Y2=0
cc_1157 N_A_2586_249#_c_1581_n N_A_3751_367#_c_2027_n 0.010996f $X=17.98 $Y=1.85
+ $X2=0 $Y2=0
cc_1158 N_A_2586_249#_c_1585_n N_VPWR_c_2103_n 0.00951574f $X=15.19 $Y=1.945
+ $X2=0 $Y2=0
cc_1159 N_A_2586_249#_c_1585_n N_VPWR_c_2093_n 0.00531456f $X=15.19 $Y=1.945
+ $X2=0 $Y2=0
cc_1160 N_A_2586_249#_c_1585_n N_KAPWR_c_2379_n 0.00642552f $X=15.19 $Y=1.945
+ $X2=0 $Y2=0
cc_1161 N_A_2586_249#_M1025_d N_KAPWR_c_2381_n 0.00726763f $X=18.07 $Y=1.95
+ $X2=0 $Y2=0
cc_1162 N_A_2586_249#_c_1585_n N_KAPWR_c_2381_n 0.00964907f $X=15.19 $Y=1.945
+ $X2=0 $Y2=0
cc_1163 N_A_2586_249#_c_1579_n N_VGND_M1030_d 0.00494917f $X=17.895 $Y=0.865
+ $X2=0 $Y2=0
cc_1164 N_A_2586_249#_M1047_g N_VGND_c_2530_n 0.00647125f $X=13.075 $Y=0.805
+ $X2=0 $Y2=0
cc_1165 N_A_2586_249#_c_1576_n N_VGND_c_2531_n 0.00867005f $X=16.93 $Y=0.34
+ $X2=0 $Y2=0
cc_1166 N_A_2586_249#_c_1578_n N_VGND_c_2531_n 0.00805183f $X=17.015 $Y=0.78
+ $X2=0 $Y2=0
cc_1167 N_A_2586_249#_c_1579_n N_VGND_c_2531_n 0.026088f $X=17.895 $Y=0.865
+ $X2=0 $Y2=0
cc_1168 N_A_2586_249#_c_1582_n N_VGND_c_2531_n 0.0190293f $X=18.18 $Y=0.575
+ $X2=0 $Y2=0
cc_1169 N_A_2586_249#_c_1582_n N_VGND_c_2532_n 0.0142341f $X=18.18 $Y=0.575
+ $X2=0 $Y2=0
cc_1170 N_A_2586_249#_c_1584_n N_VGND_c_2532_n 8.69708e-19 $X=18.12 $Y=0.865
+ $X2=0 $Y2=0
cc_1171 N_A_2586_249#_c_1573_n N_VGND_c_2545_n 0.0156992f $X=14.985 $Y=0.685
+ $X2=0 $Y2=0
cc_1172 N_A_2586_249#_c_1574_n N_VGND_c_2545_n 0.00370233f $X=14.185 $Y=0.685
+ $X2=0 $Y2=0
cc_1173 N_A_2586_249#_c_1576_n N_VGND_c_2545_n 0.115743f $X=16.93 $Y=0.34 $X2=0
+ $Y2=0
cc_1174 N_A_2586_249#_c_1577_n N_VGND_c_2545_n 0.0220501f $X=15.315 $Y=0.34
+ $X2=0 $Y2=0
cc_1175 N_A_2586_249#_c_1582_n N_VGND_c_2546_n 0.0147561f $X=18.18 $Y=0.575
+ $X2=0 $Y2=0
cc_1176 N_A_2586_249#_M1047_g N_VGND_c_2548_n 7.88961e-19 $X=13.075 $Y=0.805
+ $X2=0 $Y2=0
cc_1177 N_A_2586_249#_c_1573_n N_VGND_c_2548_n 0.0203144f $X=14.985 $Y=0.685
+ $X2=0 $Y2=0
cc_1178 N_A_2586_249#_c_1574_n N_VGND_c_2548_n 0.00462134f $X=14.185 $Y=0.685
+ $X2=0 $Y2=0
cc_1179 N_A_2586_249#_c_1576_n N_VGND_c_2548_n 0.065378f $X=16.93 $Y=0.34 $X2=0
+ $Y2=0
cc_1180 N_A_2586_249#_c_1577_n N_VGND_c_2548_n 0.0112289f $X=15.315 $Y=0.34
+ $X2=0 $Y2=0
cc_1181 N_A_2586_249#_c_1579_n N_VGND_c_2548_n 0.0176204f $X=17.895 $Y=0.865
+ $X2=0 $Y2=0
cc_1182 N_A_2586_249#_c_1582_n N_VGND_c_2548_n 0.0119945f $X=18.18 $Y=0.575
+ $X2=0 $Y2=0
cc_1183 N_A_2586_249#_c_1584_n N_VGND_c_2548_n 0.00498951f $X=18.12 $Y=0.865
+ $X2=0 $Y2=0
cc_1184 N_A_2586_249#_M1047_g N_A_2544_119#_c_2791_n 2.08092e-19 $X=13.075
+ $Y=0.805 $X2=0 $Y2=0
cc_1185 N_A_2586_249#_M1047_g N_A_2544_119#_c_2792_n 0.0138587f $X=13.075
+ $Y=0.805 $X2=0 $Y2=0
cc_1186 N_A_2586_249#_c_1570_n N_A_2544_119#_c_2792_n 0.0675896f $X=14.015
+ $Y=1.41 $X2=0 $Y2=0
cc_1187 N_A_2586_249#_c_1571_n N_A_2544_119#_c_2792_n 0.00403997f $X=13.095
+ $Y=1.41 $X2=0 $Y2=0
cc_1188 N_A_2586_249#_c_1572_n N_A_2544_119#_c_2792_n 0.014296f $X=14.1 $Y=1.32
+ $X2=0 $Y2=0
cc_1189 N_A_2586_249#_c_1570_n N_A_2544_119#_c_2793_n 0.00119838f $X=14.015
+ $Y=1.41 $X2=0 $Y2=0
cc_1190 N_A_2586_249#_c_1571_n N_A_2544_119#_c_2793_n 3.8029e-19 $X=13.095
+ $Y=1.41 $X2=0 $Y2=0
cc_1191 N_A_2586_249#_c_1572_n N_A_2544_119#_c_2794_n 0.0154587f $X=14.1 $Y=1.32
+ $X2=0 $Y2=0
cc_1192 N_A_2586_249#_c_1574_n N_A_2544_119#_c_2794_n 0.0141315f $X=14.185
+ $Y=0.685 $X2=0 $Y2=0
cc_1193 N_A_2586_249#_c_1578_n A_3407_97# 0.00336847f $X=17.015 $Y=0.78
+ $X2=-0.19 $Y2=-0.245
cc_1194 N_A_2586_249#_c_1579_n A_3407_97# 0.00165852f $X=17.895 $Y=0.865
+ $X2=-0.19 $Y2=-0.245
cc_1195 N_RESET_B_M1045_g N_VPWR_c_2101_n 0.00441827f $X=4.375 $Y=2.65 $X2=0
+ $Y2=0
cc_1196 N_RESET_B_M1041_g N_VPWR_c_2103_n 0.00951574f $X=15.65 $Y=2.45 $X2=0
+ $Y2=0
cc_1197 N_RESET_B_M1045_g N_VPWR_c_2093_n 0.00389802f $X=4.375 $Y=2.65 $X2=0
+ $Y2=0
cc_1198 N_RESET_B_M1041_g N_VPWR_c_2093_n 0.00531456f $X=15.65 $Y=2.45 $X2=0
+ $Y2=0
cc_1199 N_RESET_B_M1045_g N_A_332_136#_c_2251_n 0.0139228f $X=4.375 $Y=2.65
+ $X2=0 $Y2=0
cc_1200 RESET_B N_A_332_136#_c_2251_n 0.0203984f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_1201 N_RESET_B_c_1736_n N_A_332_136#_c_2251_n 0.00398551f $X=4.375 $Y=1.715
+ $X2=0 $Y2=0
cc_1202 N_RESET_B_M1045_g N_A_332_136#_c_2252_n 0.0266202f $X=4.375 $Y=2.65
+ $X2=0 $Y2=0
cc_1203 N_RESET_B_M1023_g N_A_332_136#_c_2242_n 6.12381e-19 $X=3.995 $Y=0.81
+ $X2=0 $Y2=0
cc_1204 N_RESET_B_c_1721_n N_A_332_136#_c_2242_n 0.00383523f $X=4.495 $Y=1.55
+ $X2=0 $Y2=0
cc_1205 RESET_B N_A_332_136#_c_2242_n 0.015854f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_1206 N_RESET_B_c_1736_n N_A_332_136#_c_2242_n 0.0122411f $X=4.375 $Y=1.715
+ $X2=0 $Y2=0
cc_1207 N_RESET_B_M1023_g N_A_332_136#_c_2244_n 2.78067e-19 $X=3.995 $Y=0.81
+ $X2=0 $Y2=0
cc_1208 N_RESET_B_c_1721_n N_A_332_136#_c_2244_n 0.00655441f $X=4.495 $Y=1.55
+ $X2=0 $Y2=0
cc_1209 N_RESET_B_c_1721_n N_A_332_136#_c_2245_n 0.00169412f $X=4.495 $Y=1.55
+ $X2=0 $Y2=0
cc_1210 N_RESET_B_M1045_g N_A_332_136#_c_2256_n 0.00388924f $X=4.375 $Y=2.65
+ $X2=0 $Y2=0
cc_1211 N_RESET_B_c_1736_n N_A_332_136#_c_2256_n 0.00360305f $X=4.375 $Y=1.715
+ $X2=0 $Y2=0
cc_1212 N_RESET_B_M1041_g N_KAPWR_c_2380_n 0.00176698f $X=15.65 $Y=2.45 $X2=0
+ $Y2=0
cc_1213 N_RESET_B_M1045_g N_KAPWR_c_2381_n 0.00699735f $X=4.375 $Y=2.65 $X2=0
+ $Y2=0
cc_1214 N_RESET_B_M1043_g N_KAPWR_c_2381_n 0.00303235f $X=6.615 $Y=2.33 $X2=0
+ $Y2=0
cc_1215 N_RESET_B_M1041_g N_KAPWR_c_2381_n 0.00924297f $X=15.65 $Y=2.45 $X2=0
+ $Y2=0
cc_1216 N_RESET_B_M1023_g N_VGND_c_2526_n 0.00593262f $X=3.995 $Y=0.81 $X2=0
+ $Y2=0
cc_1217 N_RESET_B_c_1723_n N_VGND_c_2526_n 0.00783761f $X=4.57 $Y=0.18 $X2=0
+ $Y2=0
cc_1218 N_RESET_B_M1042_g N_VGND_c_2527_n 0.0168202f $X=7 $Y=0.805 $X2=0 $Y2=0
cc_1219 N_RESET_B_c_1726_n N_VGND_c_2527_n 0.0177874f $X=13.47 $Y=0.18 $X2=0
+ $Y2=0
cc_1220 N_RESET_B_c_1731_n N_VGND_c_2527_n 0.00460513f $X=7 $Y=0.18 $X2=0 $Y2=0
cc_1221 N_RESET_B_c_1726_n N_VGND_c_2528_n 0.0247016f $X=13.47 $Y=0.18 $X2=0
+ $Y2=0
cc_1222 N_RESET_B_c_1726_n N_VGND_c_2529_n 0.0258253f $X=13.47 $Y=0.18 $X2=0
+ $Y2=0
cc_1223 N_RESET_B_c_1726_n N_VGND_c_2530_n 0.0237543f $X=13.47 $Y=0.18 $X2=0
+ $Y2=0
cc_1224 N_RESET_B_M1007_g N_VGND_c_2530_n 0.0125947f $X=13.545 $Y=0.805 $X2=0
+ $Y2=0
cc_1225 N_RESET_B_M1023_g N_VGND_c_2537_n 0.00412501f $X=3.995 $Y=0.81 $X2=0
+ $Y2=0
cc_1226 N_RESET_B_c_1723_n N_VGND_c_2537_n 0.0645079f $X=4.57 $Y=0.18 $X2=0
+ $Y2=0
cc_1227 N_RESET_B_c_1726_n N_VGND_c_2539_n 0.0197523f $X=13.47 $Y=0.18 $X2=0
+ $Y2=0
cc_1228 N_RESET_B_c_1726_n N_VGND_c_2541_n 0.0803837f $X=13.47 $Y=0.18 $X2=0
+ $Y2=0
cc_1229 N_RESET_B_c_1726_n N_VGND_c_2544_n 0.0439306f $X=13.47 $Y=0.18 $X2=0
+ $Y2=0
cc_1230 N_RESET_B_c_1726_n N_VGND_c_2545_n 0.0590637f $X=13.47 $Y=0.18 $X2=0
+ $Y2=0
cc_1231 N_RESET_B_M1023_g N_VGND_c_2548_n 0.00476395f $X=3.995 $Y=0.81 $X2=0
+ $Y2=0
cc_1232 N_RESET_B_c_1722_n N_VGND_c_2548_n 0.064943f $X=6.925 $Y=0.18 $X2=0
+ $Y2=0
cc_1233 N_RESET_B_c_1723_n N_VGND_c_2548_n 0.0116041f $X=4.57 $Y=0.18 $X2=0
+ $Y2=0
cc_1234 N_RESET_B_c_1726_n N_VGND_c_2548_n 0.180227f $X=13.47 $Y=0.18 $X2=0
+ $Y2=0
cc_1235 N_RESET_B_c_1728_n N_VGND_c_2548_n 0.0636382f $X=15.625 $Y=0.18 $X2=0
+ $Y2=0
cc_1236 N_RESET_B_c_1731_n N_VGND_c_2548_n 0.00749832f $X=7 $Y=0.18 $X2=0 $Y2=0
cc_1237 N_RESET_B_c_1733_n N_VGND_c_2548_n 0.00903773f $X=13.545 $Y=0.18 $X2=0
+ $Y2=0
cc_1238 N_RESET_B_M1023_g N_noxref_31_c_2723_n 0.0152948f $X=3.995 $Y=0.81 $X2=0
+ $Y2=0
cc_1239 N_RESET_B_c_1721_n N_noxref_31_c_2723_n 0.00189393f $X=4.495 $Y=1.55
+ $X2=0 $Y2=0
cc_1240 RESET_B N_noxref_31_c_2723_n 0.0260446f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_1241 N_RESET_B_c_1736_n N_noxref_31_c_2723_n 0.00442248f $X=4.375 $Y=1.715
+ $X2=0 $Y2=0
cc_1242 N_RESET_B_M1023_g N_noxref_31_c_2725_n 0.0156029f $X=3.995 $Y=0.81 $X2=0
+ $Y2=0
cc_1243 N_RESET_B_c_1721_n N_noxref_31_c_2725_n 0.00687666f $X=4.495 $Y=1.55
+ $X2=0 $Y2=0
cc_1244 N_RESET_B_c_1721_n N_A_929_152#_c_2755_n 0.0135097f $X=4.495 $Y=1.55
+ $X2=0 $Y2=0
cc_1245 N_RESET_B_c_1722_n N_A_929_152#_c_2756_n 0.0363931f $X=6.925 $Y=0.18
+ $X2=0 $Y2=0
cc_1246 N_RESET_B_M1042_g N_A_929_152#_c_2756_n 0.00332376f $X=7 $Y=0.805 $X2=0
+ $Y2=0
cc_1247 N_RESET_B_c_1721_n N_A_929_152#_c_2757_n 0.00799075f $X=4.495 $Y=1.55
+ $X2=0 $Y2=0
cc_1248 N_RESET_B_c_1722_n N_A_929_152#_c_2757_n 0.00707995f $X=6.925 $Y=0.18
+ $X2=0 $Y2=0
cc_1249 N_RESET_B_M1042_g N_A_929_152#_c_2758_n 0.00175158f $X=7 $Y=0.805 $X2=0
+ $Y2=0
cc_1250 N_RESET_B_c_1726_n N_A_2544_119#_c_2791_n 0.00455256f $X=13.47 $Y=0.18
+ $X2=0 $Y2=0
cc_1251 N_RESET_B_M1007_g N_A_2544_119#_c_2792_n 0.0158464f $X=13.545 $Y=0.805
+ $X2=0 $Y2=0
cc_1252 N_RESET_B_M1007_g N_A_2544_119#_c_2794_n 7.37117e-19 $X=13.545 $Y=0.805
+ $X2=0 $Y2=0
cc_1253 N_RESET_B_c_1728_n N_A_2544_119#_c_2794_n 0.00268246f $X=15.625 $Y=0.18
+ $X2=0 $Y2=0
cc_1254 N_CLK_M1048_g N_SLEEP_B_c_1931_n 0.0483985f $X=16.6 $Y=0.695 $X2=-0.19
+ $Y2=-0.245
cc_1255 N_CLK_M1024_g N_SLEEP_B_M1027_g 0.0252484f $X=16.775 $Y=2.27 $X2=0 $Y2=0
cc_1256 CLK N_SLEEP_B_M1027_g 0.00267493f $X=16.955 $Y=1.58 $X2=0 $Y2=0
cc_1257 N_CLK_c_1889_n N_SLEEP_B_M1027_g 0.0162534f $X=16.755 $Y=1.625 $X2=0
+ $Y2=0
cc_1258 N_CLK_M1048_g N_SLEEP_B_c_1935_n 0.00760632f $X=16.6 $Y=0.695 $X2=0
+ $Y2=0
cc_1259 CLK N_SLEEP_B_c_1935_n 0.00130246f $X=16.955 $Y=1.58 $X2=0 $Y2=0
cc_1260 N_CLK_c_1889_n N_SLEEP_B_c_1935_n 0.00141089f $X=16.755 $Y=1.625 $X2=0
+ $Y2=0
cc_1261 N_CLK_M1024_g N_VPWR_c_2103_n 0.00240442f $X=16.775 $Y=2.27 $X2=0 $Y2=0
cc_1262 N_CLK_M1024_g N_VPWR_c_2093_n 6.78815e-19 $X=16.775 $Y=2.27 $X2=0 $Y2=0
cc_1263 N_CLK_M1024_g N_KAPWR_c_2380_n 2.69918e-19 $X=16.775 $Y=2.27 $X2=0 $Y2=0
cc_1264 N_CLK_M1024_g N_KAPWR_c_2381_n 0.00392702f $X=16.775 $Y=2.27 $X2=0 $Y2=0
cc_1265 N_CLK_M1024_g N_KAPWR_c_2382_n 2.18323e-19 $X=16.775 $Y=2.27 $X2=0 $Y2=0
cc_1266 N_CLK_M1048_g N_VGND_c_2545_n 7.35405e-19 $X=16.6 $Y=0.695 $X2=0 $Y2=0
cc_1267 SLEEP_B N_A_3751_367#_c_2024_n 0.00203388f $X=18.395 $Y=1.21 $X2=0 $Y2=0
cc_1268 N_SLEEP_B_c_1942_n N_A_3751_367#_c_2024_n 0.0118808f $X=18.4 $Y=1.285
+ $X2=0 $Y2=0
cc_1269 N_SLEEP_B_M1014_g N_A_3751_367#_c_2025_n 0.0010233f $X=18.755 $Y=0.575
+ $X2=0 $Y2=0
cc_1270 N_SLEEP_B_M1025_g N_A_3751_367#_c_2032_n 0.00220169f $X=17.945 $Y=2.45
+ $X2=0 $Y2=0
cc_1271 N_SLEEP_B_c_1944_n N_A_3751_367#_c_2027_n 0.00117047f $X=17.945 $Y=1.815
+ $X2=0 $Y2=0
cc_1272 SLEEP_B N_A_3751_367#_c_2027_n 0.0229225f $X=18.395 $Y=1.21 $X2=0 $Y2=0
cc_1273 N_SLEEP_B_c_1942_n N_A_3751_367#_c_2027_n 0.00114849f $X=18.4 $Y=1.285
+ $X2=0 $Y2=0
cc_1274 N_SLEEP_B_M1027_g N_VPWR_c_2103_n 4.54171e-19 $X=17.235 $Y=2.27 $X2=0
+ $Y2=0
cc_1275 N_SLEEP_B_M1025_g N_VPWR_c_2103_n 0.00951574f $X=17.945 $Y=2.45 $X2=0
+ $Y2=0
cc_1276 N_SLEEP_B_M1025_g N_VPWR_c_2093_n 0.00531456f $X=17.945 $Y=2.45 $X2=0
+ $Y2=0
cc_1277 N_SLEEP_B_M1027_g N_KAPWR_c_2381_n 0.00167138f $X=17.235 $Y=2.27 $X2=0
+ $Y2=0
cc_1278 N_SLEEP_B_M1025_g N_KAPWR_c_2381_n 0.0145849f $X=17.945 $Y=2.45 $X2=0
+ $Y2=0
cc_1279 N_SLEEP_B_M1027_g N_KAPWR_c_2382_n 0.00532945f $X=17.235 $Y=2.27 $X2=0
+ $Y2=0
cc_1280 N_SLEEP_B_M1025_g N_KAPWR_c_2382_n 0.0123909f $X=17.945 $Y=2.45 $X2=0
+ $Y2=0
cc_1281 N_SLEEP_B_c_1933_n N_VGND_c_2531_n 0.0063279f $X=17.32 $Y=1.015 $X2=0
+ $Y2=0
cc_1282 N_SLEEP_B_M1012_g N_VGND_c_2531_n 0.0032554f $X=18.395 $Y=0.575 $X2=0
+ $Y2=0
cc_1283 N_SLEEP_B_M1012_g N_VGND_c_2532_n 0.00184114f $X=18.395 $Y=0.575 $X2=0
+ $Y2=0
cc_1284 N_SLEEP_B_M1014_g N_VGND_c_2532_n 0.0117013f $X=18.755 $Y=0.575 $X2=0
+ $Y2=0
cc_1285 N_SLEEP_B_c_1931_n N_VGND_c_2545_n 7.52779e-19 $X=16.96 $Y=1.015 $X2=0
+ $Y2=0
cc_1286 N_SLEEP_B_c_1933_n N_VGND_c_2545_n 0.00497279f $X=17.32 $Y=1.015 $X2=0
+ $Y2=0
cc_1287 N_SLEEP_B_M1012_g N_VGND_c_2546_n 0.00438034f $X=18.395 $Y=0.575 $X2=0
+ $Y2=0
cc_1288 N_SLEEP_B_M1014_g N_VGND_c_2546_n 0.00386543f $X=18.755 $Y=0.575 $X2=0
+ $Y2=0
cc_1289 N_SLEEP_B_c_1933_n N_VGND_c_2548_n 0.00509887f $X=17.32 $Y=1.015 $X2=0
+ $Y2=0
cc_1290 N_SLEEP_B_M1012_g N_VGND_c_2548_n 0.00838734f $X=18.395 $Y=0.575 $X2=0
+ $Y2=0
cc_1291 N_SLEEP_B_M1014_g N_VGND_c_2548_n 0.00759904f $X=18.755 $Y=0.575 $X2=0
+ $Y2=0
cc_1292 N_A_3751_367#_M1016_g N_VPWR_c_2098_n 0.0208453f $X=19.945 $Y=2.465
+ $X2=0 $Y2=0
cc_1293 N_A_3751_367#_c_2028_n N_VPWR_c_2098_n 6.78817e-19 $X=19.46 $Y=1.06
+ $X2=0 $Y2=0
cc_1294 N_A_3751_367#_c_2029_n N_VPWR_c_2098_n 0.0267814f $X=19.855 $Y=1.48
+ $X2=0 $Y2=0
cc_1295 N_A_3751_367#_c_2030_n N_VPWR_c_2098_n 0.00312162f $X=19.945 $Y=1.48
+ $X2=0 $Y2=0
cc_1296 N_A_3751_367#_M1016_g N_VPWR_c_2107_n 0.0054895f $X=19.945 $Y=2.465
+ $X2=0 $Y2=0
cc_1297 N_A_3751_367#_M1016_g N_VPWR_c_2093_n 0.0075719f $X=19.945 $Y=2.465
+ $X2=0 $Y2=0
cc_1298 N_A_3751_367#_M1016_g N_KAPWR_c_2381_n 0.0106059f $X=19.945 $Y=2.465
+ $X2=0 $Y2=0
cc_1299 N_A_3751_367#_M1016_g N_Q_c_2504_n 0.0121474f $X=19.945 $Y=2.465 $X2=0
+ $Y2=0
cc_1300 N_A_3751_367#_M1016_g Q 0.00439596f $X=19.945 $Y=2.465 $X2=0 $Y2=0
cc_1301 N_A_3751_367#_c_2029_n Q 0.00187828f $X=19.855 $Y=1.48 $X2=0 $Y2=0
cc_1302 N_A_3751_367#_c_2030_n Q 0.00649369f $X=19.945 $Y=1.48 $X2=0 $Y2=0
cc_1303 N_A_3751_367#_M1049_g N_Q_c_2503_n 0.0204893f $X=20.155 $Y=0.705 $X2=0
+ $Y2=0
cc_1304 N_A_3751_367#_c_2026_n N_Q_c_2503_n 0.00546917f $X=19.6 $Y=1.315 $X2=0
+ $Y2=0
cc_1305 N_A_3751_367#_c_2029_n N_Q_c_2503_n 0.0246274f $X=19.855 $Y=1.48 $X2=0
+ $Y2=0
cc_1306 N_A_3751_367#_c_2030_n N_Q_c_2503_n 0.0135894f $X=19.945 $Y=1.48 $X2=0
+ $Y2=0
cc_1307 N_A_3751_367#_c_2023_n N_VGND_c_2532_n 0.0125468f $X=19.235 $Y=1.06
+ $X2=0 $Y2=0
cc_1308 N_A_3751_367#_c_2024_n N_VGND_c_2532_n 0.00905894f $X=18.905 $Y=1.06
+ $X2=0 $Y2=0
cc_1309 N_A_3751_367#_c_2025_n N_VGND_c_2532_n 0.018744f $X=19.4 $Y=0.575 $X2=0
+ $Y2=0
cc_1310 N_A_3751_367#_c_2025_n N_VGND_c_2533_n 0.0203268f $X=19.4 $Y=0.575 $X2=0
+ $Y2=0
cc_1311 N_A_3751_367#_M1049_g N_VGND_c_2534_n 0.00770538f $X=20.155 $Y=0.705
+ $X2=0 $Y2=0
cc_1312 N_A_3751_367#_c_2025_n N_VGND_c_2534_n 0.0503232f $X=19.4 $Y=0.575 $X2=0
+ $Y2=0
cc_1313 N_A_3751_367#_c_2028_n N_VGND_c_2534_n 0.0141582f $X=19.46 $Y=1.06 $X2=0
+ $Y2=0
cc_1314 N_A_3751_367#_c_2029_n N_VGND_c_2534_n 0.0138307f $X=19.855 $Y=1.48
+ $X2=0 $Y2=0
cc_1315 N_A_3751_367#_c_2030_n N_VGND_c_2534_n 0.00451949f $X=19.945 $Y=1.48
+ $X2=0 $Y2=0
cc_1316 N_A_3751_367#_M1049_g N_VGND_c_2547_n 0.00502664f $X=20.155 $Y=0.705
+ $X2=0 $Y2=0
cc_1317 N_A_3751_367#_M1049_g N_VGND_c_2548_n 0.0109703f $X=20.155 $Y=0.705
+ $X2=0 $Y2=0
cc_1318 N_A_3751_367#_c_2025_n N_VGND_c_2548_n 0.0164802f $X=19.4 $Y=0.575 $X2=0
+ $Y2=0
cc_1319 N_VPWR_M1034_d N_A_332_136#_c_2267_n 0.00421102f $X=0.64 $Y=2.33 $X2=0
+ $Y2=0
cc_1320 N_VPWR_c_2094_n N_A_332_136#_c_2267_n 0.0101446f $X=0.785 $Y=2.665 $X2=0
+ $Y2=0
cc_1321 N_VPWR_c_2095_n N_A_332_136#_c_2251_n 0.0232094f $X=3.41 $Y=2.715 $X2=0
+ $Y2=0
cc_1322 N_VPWR_c_2101_n N_A_332_136#_c_2252_n 0.0151738f $X=6.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1323 N_VPWR_c_2093_n N_A_332_136#_c_2252_n 0.00320222f $X=20.4 $Y=3.33 $X2=0
+ $Y2=0
cc_1324 N_VPWR_c_2095_n N_A_332_136#_c_2254_n 0.0100786f $X=3.41 $Y=2.715 $X2=0
+ $Y2=0
cc_1325 N_VPWR_c_2099_n N_A_332_136#_c_2255_n 0.0151738f $X=3.245 $Y=3.33 $X2=0
+ $Y2=0
cc_1326 N_VPWR_c_2093_n N_A_332_136#_c_2255_n 0.00320222f $X=20.4 $Y=3.33 $X2=0
+ $Y2=0
cc_1327 N_VPWR_c_2103_n N_KAPWR_c_2379_n 0.0176805f $X=19.495 $Y=3.33 $X2=0
+ $Y2=0
cc_1328 N_VPWR_c_2093_n N_KAPWR_c_2379_n 0.00386549f $X=20.4 $Y=3.33 $X2=0 $Y2=0
cc_1329 N_VPWR_c_2103_n N_KAPWR_c_2380_n 0.0157848f $X=19.495 $Y=3.33 $X2=0
+ $Y2=0
cc_1330 N_VPWR_c_2093_n N_KAPWR_c_2380_n 0.00347494f $X=20.4 $Y=3.33 $X2=0 $Y2=0
cc_1331 N_VPWR_M1034_d N_KAPWR_c_2381_n 0.010686f $X=0.64 $Y=2.33 $X2=0 $Y2=0
cc_1332 N_VPWR_M1009_d N_KAPWR_c_2381_n 0.0157298f $X=3.27 $Y=2.33 $X2=0 $Y2=0
cc_1333 N_VPWR_M1020_d N_KAPWR_c_2381_n 0.00225196f $X=6.03 $Y=2.12 $X2=0 $Y2=0
cc_1334 N_VPWR_M1001_d N_KAPWR_c_2381_n 0.00132014f $X=7.795 $Y=1.865 $X2=0
+ $Y2=0
cc_1335 N_VPWR_M1051_d N_KAPWR_c_2381_n 0.00199666f $X=19.19 $Y=1.835 $X2=0
+ $Y2=0
cc_1336 N_VPWR_c_2094_n N_KAPWR_c_2381_n 0.0316311f $X=0.785 $Y=2.665 $X2=0
+ $Y2=0
cc_1337 N_VPWR_c_2095_n N_KAPWR_c_2381_n 0.0340722f $X=3.41 $Y=2.715 $X2=0 $Y2=0
cc_1338 N_VPWR_c_2096_n N_KAPWR_c_2381_n 0.0244927f $X=6.285 $Y=2.855 $X2=0
+ $Y2=0
cc_1339 N_VPWR_c_2097_n N_KAPWR_c_2381_n 0.0316566f $X=8.015 $Y=2.77 $X2=0 $Y2=0
cc_1340 N_VPWR_c_2098_n N_KAPWR_c_2381_n 0.0448539f $X=19.66 $Y=1.98 $X2=0 $Y2=0
cc_1341 N_VPWR_c_2099_n N_KAPWR_c_2381_n 0.0106424f $X=3.245 $Y=3.33 $X2=0 $Y2=0
cc_1342 N_VPWR_c_2101_n N_KAPWR_c_2381_n 0.00930822f $X=6.12 $Y=3.33 $X2=0 $Y2=0
cc_1343 N_VPWR_c_2103_n N_KAPWR_c_2381_n 0.0278584f $X=19.495 $Y=3.33 $X2=0
+ $Y2=0
cc_1344 N_VPWR_c_2105_n N_KAPWR_c_2381_n 0.0014101f $X=0.62 $Y=3.33 $X2=0 $Y2=0
cc_1345 N_VPWR_c_2106_n N_KAPWR_c_2381_n 0.00493877f $X=7.85 $Y=3.33 $X2=0 $Y2=0
cc_1346 N_VPWR_c_2107_n N_KAPWR_c_2381_n 0.00240987f $X=20.4 $Y=3.33 $X2=0 $Y2=0
cc_1347 N_VPWR_c_2093_n N_KAPWR_c_2381_n 2.16755f $X=20.4 $Y=3.33 $X2=0 $Y2=0
cc_1348 N_VPWR_c_2103_n N_KAPWR_c_2382_n 0.0413895f $X=19.495 $Y=3.33 $X2=0
+ $Y2=0
cc_1349 N_VPWR_c_2093_n N_KAPWR_c_2382_n 0.00720145f $X=20.4 $Y=3.33 $X2=0 $Y2=0
cc_1350 N_VPWR_c_2093_n N_Q_M1016_d 0.00119401f $X=20.4 $Y=3.33 $X2=0 $Y2=0
cc_1351 N_VPWR_c_2098_n N_Q_c_2504_n 0.0382483f $X=19.66 $Y=1.98 $X2=0 $Y2=0
cc_1352 N_VPWR_c_2107_n N_Q_c_2504_n 0.0210192f $X=20.4 $Y=3.33 $X2=0 $Y2=0
cc_1353 N_VPWR_c_2093_n N_Q_c_2504_n 0.00303861f $X=20.4 $Y=3.33 $X2=0 $Y2=0
cc_1354 N_VPWR_c_2098_n Q 0.0142958f $X=19.66 $Y=1.98 $X2=0 $Y2=0
cc_1355 A_313_466# N_A_332_136#_c_2266_n 0.0029684f $X=1.565 $Y=2.33 $X2=2.305
+ $Y2=2.425
cc_1356 A_313_466# N_KAPWR_c_2381_n 0.00318255f $X=1.565 $Y=2.33 $X2=2.635
+ $Y2=2.185
cc_1357 N_A_332_136#_M1039_d N_KAPWR_c_2381_n 0.00529062f $X=1.955 $Y=2.33 $X2=0
+ $Y2=0
cc_1358 N_A_332_136#_c_2266_n N_KAPWR_c_2381_n 0.0420077f $X=2.305 $Y=2.425
+ $X2=0 $Y2=0
cc_1359 N_A_332_136#_c_2267_n N_KAPWR_c_2381_n 0.00946083f $X=1.395 $Y=2.425
+ $X2=0 $Y2=0
cc_1360 N_A_332_136#_c_2251_n N_KAPWR_c_2381_n 0.0550803f $X=4.425 $Y=2.185
+ $X2=0 $Y2=0
cc_1361 N_A_332_136#_c_2252_n N_KAPWR_c_2381_n 0.0444408f $X=4.59 $Y=2.475 $X2=0
+ $Y2=0
cc_1362 N_A_332_136#_c_2255_n N_KAPWR_c_2381_n 0.044676f $X=2.47 $Y=2.475 $X2=0
+ $Y2=0
cc_1363 N_A_332_136#_c_2244_n N_noxref_31_c_2723_n 0.0115635f $X=4.715 $Y=1.335
+ $X2=0 $Y2=0
cc_1364 N_A_332_136#_c_2245_n N_noxref_31_c_2723_n 0.00122295f $X=5.12 $Y=1.25
+ $X2=0 $Y2=0
cc_1365 N_A_332_136#_c_2245_n N_noxref_31_c_2725_n 0.00373889f $X=5.12 $Y=1.25
+ $X2=0 $Y2=0
cc_1366 N_A_332_136#_c_2245_n N_A_929_152#_M1033_s 0.00518279f $X=5.12 $Y=1.25
+ $X2=-0.19 $Y2=-0.245
cc_1367 N_A_332_136#_c_2243_n N_A_929_152#_c_2755_n 0.012283f $X=5.035 $Y=1.335
+ $X2=0 $Y2=0
cc_1368 N_A_332_136#_c_2244_n N_A_929_152#_c_2755_n 0.00915231f $X=4.715
+ $Y=1.335 $X2=0 $Y2=0
cc_1369 N_A_332_136#_c_2245_n N_A_929_152#_c_2755_n 0.0236018f $X=5.12 $Y=1.25
+ $X2=0 $Y2=0
cc_1370 N_A_332_136#_c_2247_n N_A_929_152#_c_2755_n 0.0147378f $X=5.205 $Y=0.68
+ $X2=0 $Y2=0
cc_1371 N_A_332_136#_c_2246_n N_A_929_152#_c_2756_n 0.0628184f $X=5.725 $Y=0.68
+ $X2=0 $Y2=0
cc_1372 N_A_332_136#_c_2247_n N_A_929_152#_c_2756_n 0.0134299f $X=5.205 $Y=0.68
+ $X2=0 $Y2=0
cc_1373 N_A_332_136#_c_2246_n N_A_929_152#_c_2758_n 0.0131778f $X=5.725 $Y=0.68
+ $X2=0 $Y2=0
cc_1374 N_A_332_136#_c_2248_n N_A_929_152#_c_2758_n 0.00507506f $X=5.89 $Y=1.035
+ $X2=0 $Y2=0
cc_1375 A_552_466# N_KAPWR_c_2381_n 0.00579478f $X=2.76 $Y=2.33 $X2=17.04
+ $Y2=2.82
cc_1376 A_2836_390# N_KAPWR_c_2381_n 0.00316235f $X=14.18 $Y=1.95 $X2=11.43
+ $Y2=1.24
cc_1377 N_KAPWR_c_2381_n A_3063_390# 0.00276706f $X=17.04 $Y=2.82 $X2=-0.19
+ $Y2=1.655
cc_1378 N_KAPWR_c_2381_n N_Q_c_2504_n 0.029525f $X=17.04 $Y=2.82 $X2=0 $Y2=0
cc_1379 N_KAPWR_c_2381_n Q 0.00845277f $X=17.04 $Y=2.82 $X2=0 $Y2=0
cc_1380 N_Q_c_2503_n N_VGND_c_2534_n 0.0329135f $X=20.37 $Y=0.43 $X2=0 $Y2=0
cc_1381 N_Q_c_2503_n N_VGND_c_2547_n 0.0220321f $X=20.37 $Y=0.43 $X2=0 $Y2=0
cc_1382 N_Q_c_2503_n N_VGND_c_2548_n 0.0125808f $X=20.37 $Y=0.43 $X2=0 $Y2=0
cc_1383 N_VGND_c_2525_n N_noxref_29_c_2697_n 0.040374f $X=0.7 $Y=0.76 $X2=0
+ $Y2=0
cc_1384 N_VGND_c_2526_n N_noxref_29_c_2698_n 0.0127057f $X=3.78 $Y=0.81 $X2=0
+ $Y2=0
cc_1385 N_VGND_c_2535_n N_noxref_29_c_2698_n 0.136071f $X=3.615 $Y=0 $X2=0 $Y2=0
cc_1386 N_VGND_c_2548_n N_noxref_29_c_2698_n 0.0787034f $X=20.4 $Y=0 $X2=0 $Y2=0
cc_1387 N_VGND_c_2525_n N_noxref_29_c_2699_n 0.0131781f $X=0.7 $Y=0.76 $X2=0
+ $Y2=0
cc_1388 N_VGND_c_2535_n N_noxref_29_c_2699_n 0.0179217f $X=3.615 $Y=0 $X2=0
+ $Y2=0
cc_1389 N_VGND_c_2548_n N_noxref_29_c_2699_n 0.00971942f $X=20.4 $Y=0 $X2=0
+ $Y2=0
cc_1390 N_VGND_c_2526_n N_noxref_29_c_2700_n 0.0423098f $X=3.78 $Y=0.81 $X2=0
+ $Y2=0
cc_1391 N_VGND_c_2526_n N_noxref_31_c_2723_n 0.0209461f $X=3.78 $Y=0.81 $X2=0
+ $Y2=0
cc_1392 N_VGND_c_2526_n N_noxref_31_c_2725_n 0.0179429f $X=3.78 $Y=0.81 $X2=0
+ $Y2=0
cc_1393 N_VGND_c_2537_n N_noxref_31_c_2725_n 0.00742154f $X=7.05 $Y=0 $X2=0
+ $Y2=0
cc_1394 N_VGND_c_2548_n N_noxref_31_c_2725_n 0.0103348f $X=20.4 $Y=0 $X2=0 $Y2=0
cc_1395 N_VGND_c_2527_n N_A_929_152#_c_2756_n 0.00679944f $X=7.215 $Y=0.745
+ $X2=0 $Y2=0
cc_1396 N_VGND_c_2537_n N_A_929_152#_c_2756_n 0.112015f $X=7.05 $Y=0 $X2=0 $Y2=0
cc_1397 N_VGND_c_2548_n N_A_929_152#_c_2756_n 0.0581495f $X=20.4 $Y=0 $X2=0
+ $Y2=0
cc_1398 N_VGND_c_2537_n N_A_929_152#_c_2757_n 0.0170431f $X=7.05 $Y=0 $X2=0
+ $Y2=0
cc_1399 N_VGND_c_2548_n N_A_929_152#_c_2757_n 0.00857552f $X=20.4 $Y=0 $X2=0
+ $Y2=0
cc_1400 N_VGND_c_2527_n N_A_929_152#_c_2758_n 0.0138627f $X=7.215 $Y=0.745 $X2=0
+ $Y2=0
cc_1401 N_VGND_c_2530_n N_A_2544_119#_c_2791_n 0.00915068f $X=13.29 $Y=0.725
+ $X2=0 $Y2=0
cc_1402 N_VGND_c_2544_n N_A_2544_119#_c_2791_n 0.00558311f $X=13.125 $Y=0 $X2=0
+ $Y2=0
cc_1403 N_VGND_c_2548_n N_A_2544_119#_c_2791_n 0.00679464f $X=20.4 $Y=0 $X2=0
+ $Y2=0
cc_1404 N_VGND_M1047_d N_A_2544_119#_c_2792_n 0.00218982f $X=13.15 $Y=0.595
+ $X2=0 $Y2=0
cc_1405 N_VGND_c_2530_n N_A_2544_119#_c_2792_n 0.0185459f $X=13.29 $Y=0.725
+ $X2=0 $Y2=0
cc_1406 N_VGND_c_2530_n N_A_2544_119#_c_2794_n 0.00125617f $X=13.29 $Y=0.725
+ $X2=0 $Y2=0
cc_1407 N_VGND_c_2545_n N_A_2544_119#_c_2794_n 0.00382082f $X=17.475 $Y=0 $X2=0
+ $Y2=0
cc_1408 N_VGND_c_2548_n N_A_2544_119#_c_2794_n 0.00462135f $X=20.4 $Y=0 $X2=0
+ $Y2=0
cc_1409 N_noxref_29_c_2698_n N_noxref_31_c_2726_n 0.0125216f $X=3.155 $Y=0.34
+ $X2=0 $Y2=0
cc_1410 N_noxref_29_c_2700_n N_noxref_31_c_2723_n 0.020085f $X=3.24 $Y=0.85
+ $X2=0 $Y2=0
cc_1411 N_noxref_31_c_2725_n N_A_929_152#_c_2755_n 0.0320088f $X=4.21 $Y=0.81
+ $X2=0 $Y2=0
