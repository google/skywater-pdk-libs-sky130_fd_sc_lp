* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 a_670_125# a_270_465# a_778_447# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND GATE_N a_270_465# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR a_47_47# a_598_447# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 VGND a_47_47# a_598_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_820_99# a_670_125# a_1040_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR GATE_N a_270_465# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VPWR a_820_99# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_670_125# a_387_385# a_756_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_1040_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_778_447# a_820_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_820_99# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VPWR a_670_125# a_820_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND a_820_99# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_598_447# a_387_385# a_670_125# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_387_385# a_270_465# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_598_125# a_270_465# a_670_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_756_125# a_820_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_47_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_387_385# a_270_465# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_47_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
