* File: sky130_fd_sc_lp__clkinv_16.pxi.spice
* Created: Wed Sep  2 09:40:19 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINV_16%A N_A_M1000_g N_A_M1001_g N_A_M1002_g
+ N_A_M1003_g N_A_M1006_g N_A_M1004_g N_A_M1007_g N_A_M1005_g N_A_M1008_g
+ N_A_M1009_g N_A_M1010_g N_A_M1013_g N_A_M1011_g N_A_M1014_g N_A_M1012_g
+ N_A_M1016_g N_A_M1015_g N_A_M1018_g N_A_M1017_g N_A_M1019_g N_A_M1022_g
+ N_A_M1020_g N_A_M1028_g N_A_M1021_g N_A_M1029_g N_A_M1023_g N_A_M1031_g
+ N_A_M1024_g N_A_M1032_g N_A_M1025_g N_A_M1035_g N_A_M1026_g N_A_M1037_g
+ N_A_M1027_g N_A_M1039_g N_A_M1030_g N_A_M1033_g N_A_M1034_g N_A_M1036_g
+ N_A_M1038_g A N_A_c_206_n N_A_c_207_n N_A_c_208_n N_A_c_209_n N_A_c_210_n
+ N_A_c_211_n N_A_c_212_n N_A_c_213_n N_A_c_214_n N_A_c_215_n N_A_c_216_n
+ PM_SKY130_FD_SC_LP__CLKINV_16%A
x_PM_SKY130_FD_SC_LP__CLKINV_16%VPWR N_VPWR_M1000_s N_VPWR_M1001_s
+ N_VPWR_M1003_s N_VPWR_M1005_s N_VPWR_M1013_s N_VPWR_M1016_s N_VPWR_M1019_s
+ N_VPWR_M1021_s N_VPWR_M1024_s N_VPWR_M1026_s N_VPWR_M1030_s N_VPWR_M1034_s
+ N_VPWR_M1038_s N_VPWR_c_541_n N_VPWR_c_542_n N_VPWR_c_543_n N_VPWR_c_544_n
+ N_VPWR_c_545_n N_VPWR_c_546_n N_VPWR_c_547_n N_VPWR_c_548_n N_VPWR_c_549_n
+ N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_554_n
+ N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n
+ N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n
+ N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n
+ N_VPWR_c_570_n N_VPWR_c_571_n VPWR N_VPWR_c_572_n N_VPWR_c_573_n
+ N_VPWR_c_574_n N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n
+ N_VPWR_c_579_n N_VPWR_c_540_n PM_SKY130_FD_SC_LP__CLKINV_16%VPWR
x_PM_SKY130_FD_SC_LP__CLKINV_16%Y N_Y_M1006_s N_Y_M1008_s N_Y_M1011_s
+ N_Y_M1015_s N_Y_M1022_s N_Y_M1029_s N_Y_M1032_s N_Y_M1037_s N_Y_M1000_d
+ N_Y_M1002_d N_Y_M1004_d N_Y_M1009_d N_Y_M1014_d N_Y_M1018_d N_Y_M1020_d
+ N_Y_M1023_d N_Y_M1025_d N_Y_M1027_d N_Y_M1033_d N_Y_M1036_d N_Y_c_768_n
+ N_Y_c_796_n Y N_Y_c_777_n N_Y_c_778_n N_Y_c_769_n N_Y_c_770_n N_Y_c_771_n
+ N_Y_c_940_n N_Y_c_772_n N_Y_c_773_n N_Y_c_774_n N_Y_c_775_n N_Y_c_786_n
+ N_Y_c_787_n N_Y_c_873_n PM_SKY130_FD_SC_LP__CLKINV_16%Y
x_PM_SKY130_FD_SC_LP__CLKINV_16%VGND N_VGND_M1006_d N_VGND_M1007_d
+ N_VGND_M1010_d N_VGND_M1012_d N_VGND_M1017_d N_VGND_M1028_d N_VGND_M1031_d
+ N_VGND_M1035_d N_VGND_M1039_d N_VGND_c_1005_n N_VGND_c_1006_n N_VGND_c_1007_n
+ N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n N_VGND_c_1011_n
+ N_VGND_c_1012_n N_VGND_c_1013_n N_VGND_c_1014_n N_VGND_c_1015_n
+ N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n
+ N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n N_VGND_c_1023_n
+ N_VGND_c_1024_n N_VGND_c_1025_n N_VGND_c_1026_n VGND N_VGND_c_1027_n
+ N_VGND_c_1028_n N_VGND_c_1029_n N_VGND_c_1030_n N_VGND_c_1031_n
+ N_VGND_c_1032_n N_VGND_c_1033_n PM_SKY130_FD_SC_LP__CLKINV_16%VGND
cc_1 VNB N_A_M1000_g 0.00233375f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_2 VNB N_A_M1001_g 0.00147483f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=2.465
cc_3 VNB N_A_M1002_g 0.00147483f $X=-0.19 $Y=-0.245 $X2=1.525 $Y2=2.465
cc_4 VNB N_A_M1003_g 0.0014732f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.465
cc_5 VNB N_A_M1006_g 0.0519398f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=0.56
cc_6 VNB N_A_M1004_g 0.00146538f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=2.465
cc_7 VNB N_A_M1007_g 0.037035f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.56
cc_8 VNB N_A_M1005_g 0.00146373f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=2.465
cc_9 VNB N_A_M1008_g 0.0370346f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=0.56
cc_10 VNB N_A_M1009_g 0.00146369f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=2.465
cc_11 VNB N_A_M1010_g 0.037035f $X=-0.19 $Y=-0.245 $X2=3.675 $Y2=0.56
cc_12 VNB N_A_M1013_g 0.00146373f $X=-0.19 $Y=-0.245 $X2=3.675 $Y2=2.465
cc_13 VNB N_A_M1011_g 0.0370346f $X=-0.19 $Y=-0.245 $X2=4.105 $Y2=0.56
cc_14 VNB N_A_M1014_g 0.00146369f $X=-0.19 $Y=-0.245 $X2=4.105 $Y2=2.465
cc_15 VNB N_A_M1012_g 0.037035f $X=-0.19 $Y=-0.245 $X2=4.535 $Y2=0.56
cc_16 VNB N_A_M1016_g 0.00146373f $X=-0.19 $Y=-0.245 $X2=4.535 $Y2=2.465
cc_17 VNB N_A_M1015_g 0.0370346f $X=-0.19 $Y=-0.245 $X2=4.965 $Y2=0.56
cc_18 VNB N_A_M1018_g 0.00146369f $X=-0.19 $Y=-0.245 $X2=4.965 $Y2=2.465
cc_19 VNB N_A_M1017_g 0.037035f $X=-0.19 $Y=-0.245 $X2=5.395 $Y2=0.56
cc_20 VNB N_A_M1019_g 0.00146373f $X=-0.19 $Y=-0.245 $X2=5.395 $Y2=2.465
cc_21 VNB N_A_M1022_g 0.0370346f $X=-0.19 $Y=-0.245 $X2=5.825 $Y2=0.56
cc_22 VNB N_A_M1020_g 0.00146369f $X=-0.19 $Y=-0.245 $X2=5.825 $Y2=2.465
cc_23 VNB N_A_M1028_g 0.037035f $X=-0.19 $Y=-0.245 $X2=6.255 $Y2=0.56
cc_24 VNB N_A_M1021_g 0.00146373f $X=-0.19 $Y=-0.245 $X2=6.255 $Y2=2.465
cc_25 VNB N_A_M1029_g 0.0370346f $X=-0.19 $Y=-0.245 $X2=6.685 $Y2=0.56
cc_26 VNB N_A_M1023_g 0.00146369f $X=-0.19 $Y=-0.245 $X2=6.685 $Y2=2.465
cc_27 VNB N_A_M1031_g 0.037035f $X=-0.19 $Y=-0.245 $X2=7.115 $Y2=0.56
cc_28 VNB N_A_M1024_g 0.00146373f $X=-0.19 $Y=-0.245 $X2=7.115 $Y2=2.465
cc_29 VNB N_A_M1032_g 0.0370346f $X=-0.19 $Y=-0.245 $X2=7.545 $Y2=0.56
cc_30 VNB N_A_M1025_g 0.00146369f $X=-0.19 $Y=-0.245 $X2=7.545 $Y2=2.465
cc_31 VNB N_A_M1035_g 0.037035f $X=-0.19 $Y=-0.245 $X2=7.975 $Y2=0.56
cc_32 VNB N_A_M1026_g 0.00146373f $X=-0.19 $Y=-0.245 $X2=7.975 $Y2=2.465
cc_33 VNB N_A_M1037_g 0.0370346f $X=-0.19 $Y=-0.245 $X2=8.405 $Y2=0.56
cc_34 VNB N_A_M1027_g 0.00146369f $X=-0.19 $Y=-0.245 $X2=8.405 $Y2=2.465
cc_35 VNB N_A_M1039_g 0.0519399f $X=-0.19 $Y=-0.245 $X2=8.835 $Y2=0.56
cc_36 VNB N_A_M1030_g 0.00146537f $X=-0.19 $Y=-0.245 $X2=8.835 $Y2=2.465
cc_37 VNB N_A_M1033_g 0.00147314f $X=-0.19 $Y=-0.245 $X2=9.265 $Y2=2.465
cc_38 VNB N_A_M1034_g 0.00147483f $X=-0.19 $Y=-0.245 $X2=9.695 $Y2=2.465
cc_39 VNB N_A_M1036_g 0.00147483f $X=-0.19 $Y=-0.245 $X2=10.125 $Y2=2.465
cc_40 VNB N_A_M1038_g 0.00233375f $X=-0.19 $Y=-0.245 $X2=10.555 $Y2=2.465
cc_41 VNB N_A_c_206_n 0.597321f $X=-0.19 $Y=-0.245 $X2=10.555 $Y2=1.46
cc_42 VNB N_A_c_207_n 0.0693329f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.295
cc_43 VNB N_A_c_208_n 0.00550596f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.295
cc_44 VNB N_A_c_209_n 0.00550596f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=1.295
cc_45 VNB N_A_c_210_n 0.00550596f $X=-0.19 $Y=-0.245 $X2=4.755 $Y2=1.295
cc_46 VNB N_A_c_211_n 0.00550596f $X=-0.19 $Y=-0.245 $X2=5.61 $Y2=1.295
cc_47 VNB N_A_c_212_n 0.00550596f $X=-0.19 $Y=-0.245 $X2=6.475 $Y2=1.295
cc_48 VNB N_A_c_213_n 0.00550596f $X=-0.19 $Y=-0.245 $X2=7.335 $Y2=1.295
cc_49 VNB N_A_c_214_n 0.00550596f $X=-0.19 $Y=-0.245 $X2=8.195 $Y2=1.295
cc_50 VNB N_A_c_215_n 0.0659587f $X=-0.19 $Y=-0.245 $X2=9.3 $Y2=1.295
cc_51 VNB N_A_c_216_n 0.0131001f $X=-0.19 $Y=-0.245 $X2=10.38 $Y2=1.295
cc_52 VNB N_VPWR_c_540_n 0.462217f $X=-0.19 $Y=-0.245 $X2=7.115 $Y2=1.46
cc_53 VNB N_Y_c_768_n 0.011055f $X=-0.19 $Y=-0.245 $X2=4.535 $Y2=2.465
cc_54 VNB N_Y_c_769_n 0.0116226f $X=-0.19 $Y=-0.245 $X2=5.825 $Y2=2.465
cc_55 VNB N_Y_c_770_n 0.011055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Y_c_771_n 0.011055f $X=-0.19 $Y=-0.245 $X2=7.115 $Y2=0.56
cc_57 VNB N_Y_c_772_n 0.011055f $X=-0.19 $Y=-0.245 $X2=7.975 $Y2=0.56
cc_58 VNB N_Y_c_773_n 0.011055f $X=-0.19 $Y=-0.245 $X2=8.405 $Y2=1.625
cc_59 VNB N_Y_c_774_n 0.011055f $X=-0.19 $Y=-0.245 $X2=8.835 $Y2=2.465
cc_60 VNB N_Y_c_775_n 0.0116221f $X=-0.19 $Y=-0.245 $X2=10.125 $Y2=1.625
cc_61 VNB N_VGND_c_1005_n 0.0245466f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=2.465
cc_62 VNB N_VGND_c_1006_n 0.00701118f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=0.56
cc_63 VNB N_VGND_c_1007_n 0.00701118f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=2.465
cc_64 VNB N_VGND_c_1008_n 0.00701118f $X=-0.19 $Y=-0.245 $X2=3.675 $Y2=0.56
cc_65 VNB N_VGND_c_1009_n 0.0170098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1010_n 0.00701118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1011_n 0.00701118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1012_n 0.00701118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1013_n 0.00701118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1014_n 0.0244578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1015_n 0.0170098f $X=-0.19 $Y=-0.245 $X2=4.965 $Y2=0.56
cc_72 VNB N_VGND_c_1016_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1017_n 0.0170098f $X=-0.19 $Y=-0.245 $X2=4.965 $Y2=2.465
cc_74 VNB N_VGND_c_1018_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=4.965 $Y2=2.465
cc_75 VNB N_VGND_c_1019_n 0.0170098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1020_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=5.395 $Y2=1.295
cc_77 VNB N_VGND_c_1021_n 0.0170098f $X=-0.19 $Y=-0.245 $X2=5.395 $Y2=0.56
cc_78 VNB N_VGND_c_1022_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1023_n 0.0170098f $X=-0.19 $Y=-0.245 $X2=5.395 $Y2=2.465
cc_80 VNB N_VGND_c_1024_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=5.395 $Y2=2.465
cc_81 VNB N_VGND_c_1025_n 0.0170098f $X=-0.19 $Y=-0.245 $X2=5.825 $Y2=1.295
cc_82 VNB N_VGND_c_1026_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=5.825 $Y2=0.56
cc_83 VNB N_VGND_c_1027_n 0.0669011f $X=-0.19 $Y=-0.245 $X2=5.825 $Y2=1.625
cc_84 VNB N_VGND_c_1028_n 0.0170098f $X=-0.19 $Y=-0.245 $X2=6.685 $Y2=2.465
cc_85 VNB N_VGND_c_1029_n 0.0611731f $X=-0.19 $Y=-0.245 $X2=7.975 $Y2=0.56
cc_86 VNB N_VGND_c_1030_n 0.690211f $X=-0.19 $Y=-0.245 $X2=7.975 $Y2=0.56
cc_87 VNB N_VGND_c_1031_n 0.00519339f $X=-0.19 $Y=-0.245 $X2=7.975 $Y2=2.465
cc_88 VNB N_VGND_c_1032_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=8.405 $Y2=1.295
cc_89 VNB N_VGND_c_1033_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VPB N_A_M1000_g 0.0277951f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_91 VPB N_A_M1001_g 0.0198162f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=2.465
cc_92 VPB N_A_M1002_g 0.0198162f $X=-0.19 $Y=1.655 $X2=1.525 $Y2=2.465
cc_93 VPB N_A_M1003_g 0.0198061f $X=-0.19 $Y=1.655 $X2=1.955 $Y2=2.465
cc_94 VPB N_A_M1004_g 0.0197576f $X=-0.19 $Y=1.655 $X2=2.385 $Y2=2.465
cc_95 VPB N_A_M1005_g 0.0197473f $X=-0.19 $Y=1.655 $X2=2.815 $Y2=2.465
cc_96 VPB N_A_M1009_g 0.0197471f $X=-0.19 $Y=1.655 $X2=3.245 $Y2=2.465
cc_97 VPB N_A_M1013_g 0.0197473f $X=-0.19 $Y=1.655 $X2=3.675 $Y2=2.465
cc_98 VPB N_A_M1014_g 0.0197471f $X=-0.19 $Y=1.655 $X2=4.105 $Y2=2.465
cc_99 VPB N_A_M1016_g 0.0197473f $X=-0.19 $Y=1.655 $X2=4.535 $Y2=2.465
cc_100 VPB N_A_M1018_g 0.0197471f $X=-0.19 $Y=1.655 $X2=4.965 $Y2=2.465
cc_101 VPB N_A_M1019_g 0.0197473f $X=-0.19 $Y=1.655 $X2=5.395 $Y2=2.465
cc_102 VPB N_A_M1020_g 0.0197471f $X=-0.19 $Y=1.655 $X2=5.825 $Y2=2.465
cc_103 VPB N_A_M1021_g 0.0197473f $X=-0.19 $Y=1.655 $X2=6.255 $Y2=2.465
cc_104 VPB N_A_M1023_g 0.0197471f $X=-0.19 $Y=1.655 $X2=6.685 $Y2=2.465
cc_105 VPB N_A_M1024_g 0.0197473f $X=-0.19 $Y=1.655 $X2=7.115 $Y2=2.465
cc_106 VPB N_A_M1025_g 0.0197471f $X=-0.19 $Y=1.655 $X2=7.545 $Y2=2.465
cc_107 VPB N_A_M1026_g 0.0197473f $X=-0.19 $Y=1.655 $X2=7.975 $Y2=2.465
cc_108 VPB N_A_M1027_g 0.0197471f $X=-0.19 $Y=1.655 $X2=8.405 $Y2=2.465
cc_109 VPB N_A_M1030_g 0.0197575f $X=-0.19 $Y=1.655 $X2=8.835 $Y2=2.465
cc_110 VPB N_A_M1033_g 0.0198057f $X=-0.19 $Y=1.655 $X2=9.265 $Y2=2.465
cc_111 VPB N_A_M1034_g 0.0198162f $X=-0.19 $Y=1.655 $X2=9.695 $Y2=2.465
cc_112 VPB N_A_M1036_g 0.0198162f $X=-0.19 $Y=1.655 $X2=10.125 $Y2=2.465
cc_113 VPB N_A_M1038_g 0.0277951f $X=-0.19 $Y=1.655 $X2=10.555 $Y2=2.465
cc_114 VPB N_VPWR_c_541_n 0.0132644f $X=-0.19 $Y=1.655 $X2=3.675 $Y2=0.56
cc_115 VPB N_VPWR_c_542_n 0.0167406f $X=-0.19 $Y=1.655 $X2=3.675 $Y2=2.465
cc_116 VPB N_VPWR_c_543_n 0.00521585f $X=-0.19 $Y=1.655 $X2=4.105 $Y2=0.56
cc_117 VPB N_VPWR_c_544_n 0.00521585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_545_n 0.00521585f $X=-0.19 $Y=1.655 $X2=4.535 $Y2=2.465
cc_119 VPB N_VPWR_c_546_n 0.00521585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_547_n 0.00521585f $X=-0.19 $Y=1.655 $X2=5.395 $Y2=0.56
cc_121 VPB N_VPWR_c_548_n 0.0166954f $X=-0.19 $Y=1.655 $X2=5.395 $Y2=2.465
cc_122 VPB N_VPWR_c_549_n 0.00521585f $X=-0.19 $Y=1.655 $X2=5.825 $Y2=0.56
cc_123 VPB N_VPWR_c_550_n 0.00521585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_551_n 0.00521585f $X=-0.19 $Y=1.655 $X2=6.255 $Y2=2.465
cc_125 VPB N_VPWR_c_552_n 0.00521585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_553_n 0.00521585f $X=-0.19 $Y=1.655 $X2=7.115 $Y2=0.56
cc_127 VPB N_VPWR_c_554_n 0.0167406f $X=-0.19 $Y=1.655 $X2=7.115 $Y2=2.465
cc_128 VPB N_VPWR_c_555_n 0.00521585f $X=-0.19 $Y=1.655 $X2=7.545 $Y2=0.56
cc_129 VPB N_VPWR_c_556_n 0.0117052f $X=-0.19 $Y=1.655 $X2=7.545 $Y2=2.465
cc_130 VPB N_VPWR_c_557_n 0.013033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_558_n 0.0123263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_559_n 0.00497514f $X=-0.19 $Y=1.655 $X2=7.975 $Y2=1.625
cc_133 VPB N_VPWR_c_560_n 0.0167406f $X=-0.19 $Y=1.655 $X2=7.975 $Y2=2.465
cc_134 VPB N_VPWR_c_561_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_562_n 0.0167406f $X=-0.19 $Y=1.655 $X2=8.405 $Y2=0.56
cc_136 VPB N_VPWR_c_563_n 0.00497514f $X=-0.19 $Y=1.655 $X2=8.405 $Y2=0.56
cc_137 VPB N_VPWR_c_564_n 0.0167406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_565_n 0.00497514f $X=-0.19 $Y=1.655 $X2=8.405 $Y2=1.625
cc_139 VPB N_VPWR_c_566_n 0.0167406f $X=-0.19 $Y=1.655 $X2=8.405 $Y2=2.465
cc_140 VPB N_VPWR_c_567_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_568_n 0.0167406f $X=-0.19 $Y=1.655 $X2=8.835 $Y2=0.56
cc_142 VPB N_VPWR_c_569_n 0.00497514f $X=-0.19 $Y=1.655 $X2=8.835 $Y2=0.56
cc_143 VPB N_VPWR_c_570_n 0.0167406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_571_n 0.00497514f $X=-0.19 $Y=1.655 $X2=8.835 $Y2=1.625
cc_145 VPB N_VPWR_c_572_n 0.0167406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_573_n 0.0167406f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.46
cc_147 VPB N_VPWR_c_574_n 0.0166954f $X=-0.19 $Y=1.655 $X2=3.035 $Y2=1.46
cc_148 VPB N_VPWR_c_575_n 0.00497514f $X=-0.19 $Y=1.655 $X2=4.105 $Y2=1.46
cc_149 VPB N_VPWR_c_576_n 0.00497514f $X=-0.19 $Y=1.655 $X2=4.755 $Y2=1.46
cc_150 VPB N_VPWR_c_577_n 0.00497514f $X=-0.19 $Y=1.655 $X2=5.395 $Y2=1.46
cc_151 VPB N_VPWR_c_578_n 0.00497514f $X=-0.19 $Y=1.655 $X2=5.61 $Y2=1.46
cc_152 VPB N_VPWR_c_579_n 0.00497514f $X=-0.19 $Y=1.655 $X2=6.475 $Y2=1.46
cc_153 VPB N_VPWR_c_540_n 0.0552847f $X=-0.19 $Y=1.655 $X2=7.115 $Y2=1.46
cc_154 VPB N_Y_c_768_n 0.00318723f $X=-0.19 $Y=1.655 $X2=4.535 $Y2=2.465
cc_155 VPB N_Y_c_777_n 0.00120588f $X=-0.19 $Y=1.655 $X2=4.965 $Y2=2.465
cc_156 VPB N_Y_c_778_n 0.00120588f $X=-0.19 $Y=1.655 $X2=5.395 $Y2=2.465
cc_157 VPB N_Y_c_769_n 0.00342968f $X=-0.19 $Y=1.655 $X2=5.825 $Y2=2.465
cc_158 VPB N_Y_c_770_n 0.00318723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_Y_c_771_n 0.00318723f $X=-0.19 $Y=1.655 $X2=7.115 $Y2=0.56
cc_160 VPB N_Y_c_772_n 0.00318723f $X=-0.19 $Y=1.655 $X2=7.975 $Y2=0.56
cc_161 VPB N_Y_c_773_n 0.00318723f $X=-0.19 $Y=1.655 $X2=8.405 $Y2=1.625
cc_162 VPB N_Y_c_774_n 0.00318723f $X=-0.19 $Y=1.655 $X2=8.835 $Y2=2.465
cc_163 VPB N_Y_c_775_n 0.00342949f $X=-0.19 $Y=1.655 $X2=10.125 $Y2=1.625
cc_164 VPB N_Y_c_786_n 0.00120588f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.46
cc_165 VPB N_Y_c_787_n 0.00120588f $X=-0.19 $Y=1.655 $X2=2.22 $Y2=1.46
cc_166 N_A_M1000_g N_VPWR_c_541_n 0.00520924f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A_M1000_g N_VPWR_c_542_n 0.00585385f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A_M1001_g N_VPWR_c_542_n 0.00585385f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_M1001_g N_VPWR_c_543_n 0.00237003f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_M1002_g N_VPWR_c_543_n 0.00237871f $X=1.525 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A_c_206_n N_VPWR_c_543_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_172 N_A_c_207_n N_VPWR_c_543_n 0.0124345f $X=0.86 $Y=1.295 $X2=0 $Y2=0
cc_173 N_A_c_216_n N_VPWR_c_543_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_174 N_A_M1003_g N_VPWR_c_544_n 0.00237003f $X=1.955 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A_M1004_g N_VPWR_c_544_n 0.00237871f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_c_206_n N_VPWR_c_544_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_177 N_A_c_207_n N_VPWR_c_544_n 0.0124345f $X=0.86 $Y=1.295 $X2=0 $Y2=0
cc_178 N_A_c_216_n N_VPWR_c_544_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_179 N_A_M1005_g N_VPWR_c_545_n 0.00237003f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_M1009_g N_VPWR_c_545_n 0.00237871f $X=3.245 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A_c_206_n N_VPWR_c_545_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_182 N_A_c_208_n N_VPWR_c_545_n 0.0124345f $X=3.035 $Y=1.295 $X2=0 $Y2=0
cc_183 N_A_c_216_n N_VPWR_c_545_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_184 N_A_M1013_g N_VPWR_c_546_n 0.00237003f $X=3.675 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_M1014_g N_VPWR_c_546_n 0.00237871f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_c_206_n N_VPWR_c_546_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_187 N_A_c_209_n N_VPWR_c_546_n 0.0124345f $X=3.89 $Y=1.295 $X2=0 $Y2=0
cc_188 N_A_c_216_n N_VPWR_c_546_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_189 N_A_M1016_g N_VPWR_c_547_n 0.00237003f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A_M1018_g N_VPWR_c_547_n 0.00237003f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_c_206_n N_VPWR_c_547_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_192 N_A_c_210_n N_VPWR_c_547_n 0.0124345f $X=4.755 $Y=1.295 $X2=0 $Y2=0
cc_193 N_A_c_216_n N_VPWR_c_547_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_194 N_A_M1018_g N_VPWR_c_548_n 0.00585385f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A_M1019_g N_VPWR_c_548_n 0.00585385f $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A_M1019_g N_VPWR_c_549_n 0.00237003f $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A_M1020_g N_VPWR_c_549_n 0.00237871f $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A_c_206_n N_VPWR_c_549_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_199 N_A_c_211_n N_VPWR_c_549_n 0.0124345f $X=5.61 $Y=1.295 $X2=0 $Y2=0
cc_200 N_A_c_216_n N_VPWR_c_549_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_201 N_A_M1021_g N_VPWR_c_550_n 0.00237003f $X=6.255 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A_M1023_g N_VPWR_c_550_n 0.00237871f $X=6.685 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A_c_206_n N_VPWR_c_550_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_204 N_A_c_212_n N_VPWR_c_550_n 0.0124345f $X=6.475 $Y=1.295 $X2=0 $Y2=0
cc_205 N_A_c_216_n N_VPWR_c_550_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_206 N_A_M1024_g N_VPWR_c_551_n 0.00237003f $X=7.115 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_M1025_g N_VPWR_c_551_n 0.00237871f $X=7.545 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A_c_206_n N_VPWR_c_551_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_209 N_A_c_213_n N_VPWR_c_551_n 0.0124345f $X=7.335 $Y=1.295 $X2=0 $Y2=0
cc_210 N_A_c_216_n N_VPWR_c_551_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_211 N_A_M1026_g N_VPWR_c_552_n 0.00237003f $X=7.975 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A_M1027_g N_VPWR_c_552_n 0.00237871f $X=8.405 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A_c_206_n N_VPWR_c_552_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_214 N_A_c_214_n N_VPWR_c_552_n 0.0124345f $X=8.195 $Y=1.295 $X2=0 $Y2=0
cc_215 N_A_c_216_n N_VPWR_c_552_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_216 N_A_M1030_g N_VPWR_c_553_n 0.00237003f $X=8.835 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_M1033_g N_VPWR_c_553_n 0.00237871f $X=9.265 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A_c_206_n N_VPWR_c_553_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_219 N_A_c_215_n N_VPWR_c_553_n 0.0124345f $X=9.3 $Y=1.295 $X2=0 $Y2=0
cc_220 N_A_c_216_n N_VPWR_c_553_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_221 N_A_M1033_g N_VPWR_c_554_n 0.00585385f $X=9.265 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A_M1034_g N_VPWR_c_554_n 0.00585385f $X=9.695 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A_M1034_g N_VPWR_c_555_n 0.00237003f $X=9.695 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_M1036_g N_VPWR_c_555_n 0.00237003f $X=10.125 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A_c_206_n N_VPWR_c_555_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_226 N_A_c_215_n N_VPWR_c_555_n 0.0124345f $X=9.3 $Y=1.295 $X2=0 $Y2=0
cc_227 N_A_c_216_n N_VPWR_c_555_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_228 N_A_M1038_g N_VPWR_c_557_n 0.00520659f $X=10.555 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A_M1004_g N_VPWR_c_560_n 0.00585385f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A_M1005_g N_VPWR_c_560_n 0.00585385f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_M1009_g N_VPWR_c_562_n 0.00585385f $X=3.245 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A_M1013_g N_VPWR_c_562_n 0.00585385f $X=3.675 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A_M1014_g N_VPWR_c_564_n 0.00585385f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A_M1016_g N_VPWR_c_564_n 0.00585385f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A_M1023_g N_VPWR_c_566_n 0.00585385f $X=6.685 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A_M1024_g N_VPWR_c_566_n 0.00585385f $X=7.115 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A_M1025_g N_VPWR_c_568_n 0.00585385f $X=7.545 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A_M1026_g N_VPWR_c_568_n 0.00585385f $X=7.975 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A_M1027_g N_VPWR_c_570_n 0.00585385f $X=8.405 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_M1030_g N_VPWR_c_570_n 0.00585385f $X=8.835 $Y=2.465 $X2=0 $Y2=0
cc_241 N_A_M1002_g N_VPWR_c_572_n 0.00585385f $X=1.525 $Y=2.465 $X2=0 $Y2=0
cc_242 N_A_M1003_g N_VPWR_c_572_n 0.00585385f $X=1.955 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A_M1020_g N_VPWR_c_573_n 0.00585385f $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A_M1021_g N_VPWR_c_573_n 0.00585385f $X=6.255 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A_M1036_g N_VPWR_c_574_n 0.00585385f $X=10.125 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A_M1038_g N_VPWR_c_574_n 0.00585385f $X=10.555 $Y=2.465 $X2=0 $Y2=0
cc_247 N_A_M1000_g N_VPWR_c_540_n 0.011797f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A_M1001_g N_VPWR_c_540_n 0.0106452f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A_M1002_g N_VPWR_c_540_n 0.0106452f $X=1.525 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A_M1003_g N_VPWR_c_540_n 0.0106452f $X=1.955 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A_M1004_g N_VPWR_c_540_n 0.0106452f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_252 N_A_M1005_g N_VPWR_c_540_n 0.0106452f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_253 N_A_M1009_g N_VPWR_c_540_n 0.0106452f $X=3.245 $Y=2.465 $X2=0 $Y2=0
cc_254 N_A_M1013_g N_VPWR_c_540_n 0.0106452f $X=3.675 $Y=2.465 $X2=0 $Y2=0
cc_255 N_A_M1014_g N_VPWR_c_540_n 0.0106452f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_256 N_A_M1016_g N_VPWR_c_540_n 0.0106452f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A_M1018_g N_VPWR_c_540_n 0.0106452f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A_M1019_g N_VPWR_c_540_n 0.0106452f $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A_M1020_g N_VPWR_c_540_n 0.0106452f $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A_M1021_g N_VPWR_c_540_n 0.0106452f $X=6.255 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A_M1023_g N_VPWR_c_540_n 0.0106452f $X=6.685 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A_M1024_g N_VPWR_c_540_n 0.0106452f $X=7.115 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A_M1025_g N_VPWR_c_540_n 0.0106452f $X=7.545 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A_M1026_g N_VPWR_c_540_n 0.0106452f $X=7.975 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A_M1027_g N_VPWR_c_540_n 0.0106452f $X=8.405 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A_M1030_g N_VPWR_c_540_n 0.0106452f $X=8.835 $Y=2.465 $X2=0 $Y2=0
cc_267 N_A_M1033_g N_VPWR_c_540_n 0.0106452f $X=9.265 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A_M1034_g N_VPWR_c_540_n 0.0106452f $X=9.695 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A_M1036_g N_VPWR_c_540_n 0.0106452f $X=10.125 $Y=2.465 $X2=0 $Y2=0
cc_270 N_A_M1038_g N_VPWR_c_540_n 0.0116596f $X=10.555 $Y=2.465 $X2=0 $Y2=0
cc_271 N_A_M1015_g N_Y_c_768_n 0.00656691f $X=4.965 $Y=0.56 $X2=0 $Y2=0
cc_272 N_A_M1018_g N_Y_c_768_n 0.00303055f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A_M1017_g N_Y_c_768_n 0.00663665f $X=5.395 $Y=0.56 $X2=0 $Y2=0
cc_274 N_A_M1019_g N_Y_c_768_n 0.00370846f $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A_c_206_n N_Y_c_768_n 0.0205099f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_276 N_A_c_210_n N_Y_c_768_n 0.0328715f $X=4.755 $Y=1.295 $X2=0 $Y2=0
cc_277 N_A_c_211_n N_Y_c_768_n 0.0328715f $X=5.61 $Y=1.295 $X2=0 $Y2=0
cc_278 N_A_c_216_n N_Y_c_768_n 0.0321248f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_279 N_A_M1018_g N_Y_c_796_n 6.4719e-19 $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_280 N_A_M1000_g N_Y_c_777_n 6.94171e-19 $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_281 N_A_M1001_g N_Y_c_777_n 6.9407e-19 $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_282 N_A_c_206_n N_Y_c_777_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_283 N_A_c_207_n N_Y_c_777_n 0.0122997f $X=0.86 $Y=1.295 $X2=0 $Y2=0
cc_284 N_A_c_216_n N_Y_c_777_n 9.17266e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_285 N_A_M1002_g N_Y_c_778_n 6.94171e-19 $X=1.525 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A_M1003_g N_Y_c_778_n 6.9407e-19 $X=1.955 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A_c_206_n N_Y_c_778_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_288 N_A_c_207_n N_Y_c_778_n 0.0122997f $X=0.86 $Y=1.295 $X2=0 $Y2=0
cc_289 N_A_c_216_n N_Y_c_778_n 9.17266e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_290 N_A_M1006_g N_Y_c_769_n 0.0115656f $X=2.385 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A_M1004_g N_Y_c_769_n 0.00636465f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A_M1007_g N_Y_c_769_n 0.00663665f $X=2.815 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A_M1005_g N_Y_c_769_n 0.00370909f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A_c_206_n N_Y_c_769_n 0.0205099f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_295 N_A_c_207_n N_Y_c_769_n 0.0343615f $X=0.86 $Y=1.295 $X2=0 $Y2=0
cc_296 N_A_c_208_n N_Y_c_769_n 0.0328715f $X=3.035 $Y=1.295 $X2=0 $Y2=0
cc_297 N_A_c_216_n N_Y_c_769_n 0.0321248f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_298 N_A_M1008_g N_Y_c_770_n 0.00656691f $X=3.245 $Y=0.56 $X2=0 $Y2=0
cc_299 N_A_M1009_g N_Y_c_770_n 0.00367895f $X=3.245 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A_M1010_g N_Y_c_770_n 0.00663665f $X=3.675 $Y=0.56 $X2=0 $Y2=0
cc_301 N_A_M1013_g N_Y_c_770_n 0.00370909f $X=3.675 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A_c_206_n N_Y_c_770_n 0.0205099f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_303 N_A_c_208_n N_Y_c_770_n 0.0328715f $X=3.035 $Y=1.295 $X2=0 $Y2=0
cc_304 N_A_c_209_n N_Y_c_770_n 0.0328715f $X=3.89 $Y=1.295 $X2=0 $Y2=0
cc_305 N_A_c_216_n N_Y_c_770_n 0.0321248f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_306 N_A_M1011_g N_Y_c_771_n 0.00656691f $X=4.105 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A_M1014_g N_Y_c_771_n 0.00367895f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_308 N_A_M1012_g N_Y_c_771_n 0.00663665f $X=4.535 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A_M1016_g N_Y_c_771_n 0.00370909f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_310 N_A_c_206_n N_Y_c_771_n 0.0205099f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_311 N_A_c_209_n N_Y_c_771_n 0.0328715f $X=3.89 $Y=1.295 $X2=0 $Y2=0
cc_312 N_A_c_210_n N_Y_c_771_n 0.0328715f $X=4.755 $Y=1.295 $X2=0 $Y2=0
cc_313 N_A_c_216_n N_Y_c_771_n 0.0321248f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_314 N_A_M1022_g N_Y_c_772_n 0.00656691f $X=5.825 $Y=0.56 $X2=0 $Y2=0
cc_315 N_A_M1020_g N_Y_c_772_n 0.00367895f $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_316 N_A_M1028_g N_Y_c_772_n 0.00663665f $X=6.255 $Y=0.56 $X2=0 $Y2=0
cc_317 N_A_M1021_g N_Y_c_772_n 0.00370909f $X=6.255 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A_c_206_n N_Y_c_772_n 0.0205099f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_319 N_A_c_211_n N_Y_c_772_n 0.0328715f $X=5.61 $Y=1.295 $X2=0 $Y2=0
cc_320 N_A_c_212_n N_Y_c_772_n 0.0328715f $X=6.475 $Y=1.295 $X2=0 $Y2=0
cc_321 N_A_c_216_n N_Y_c_772_n 0.0321248f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_322 N_A_M1029_g N_Y_c_773_n 0.00656691f $X=6.685 $Y=0.56 $X2=0 $Y2=0
cc_323 N_A_M1023_g N_Y_c_773_n 0.00367895f $X=6.685 $Y=2.465 $X2=0 $Y2=0
cc_324 N_A_M1031_g N_Y_c_773_n 0.00663665f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_325 N_A_M1024_g N_Y_c_773_n 0.00370909f $X=7.115 $Y=2.465 $X2=0 $Y2=0
cc_326 N_A_c_206_n N_Y_c_773_n 0.0205099f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_327 N_A_c_212_n N_Y_c_773_n 0.0328715f $X=6.475 $Y=1.295 $X2=0 $Y2=0
cc_328 N_A_c_213_n N_Y_c_773_n 0.0328715f $X=7.335 $Y=1.295 $X2=0 $Y2=0
cc_329 N_A_c_216_n N_Y_c_773_n 0.0321248f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_330 N_A_M1032_g N_Y_c_774_n 0.00656691f $X=7.545 $Y=0.56 $X2=0 $Y2=0
cc_331 N_A_M1025_g N_Y_c_774_n 0.00367895f $X=7.545 $Y=2.465 $X2=0 $Y2=0
cc_332 N_A_M1035_g N_Y_c_774_n 0.00663665f $X=7.975 $Y=0.56 $X2=0 $Y2=0
cc_333 N_A_M1026_g N_Y_c_774_n 0.00370909f $X=7.975 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A_c_206_n N_Y_c_774_n 0.0205099f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_335 N_A_c_213_n N_Y_c_774_n 0.0328715f $X=7.335 $Y=1.295 $X2=0 $Y2=0
cc_336 N_A_c_214_n N_Y_c_774_n 0.0328715f $X=8.195 $Y=1.295 $X2=0 $Y2=0
cc_337 N_A_c_216_n N_Y_c_774_n 0.0321248f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_338 N_A_M1037_g N_Y_c_775_n 0.00656691f $X=8.405 $Y=0.56 $X2=0 $Y2=0
cc_339 N_A_M1027_g N_Y_c_775_n 0.00367895f $X=8.405 $Y=2.465 $X2=0 $Y2=0
cc_340 N_A_M1039_g N_Y_c_775_n 0.0116468f $X=8.835 $Y=0.56 $X2=0 $Y2=0
cc_341 N_A_M1030_g N_Y_c_775_n 0.00640091f $X=8.835 $Y=2.465 $X2=0 $Y2=0
cc_342 N_A_c_206_n N_Y_c_775_n 0.0205099f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_343 N_A_c_214_n N_Y_c_775_n 0.0328715f $X=8.195 $Y=1.295 $X2=0 $Y2=0
cc_344 N_A_c_215_n N_Y_c_775_n 0.0343615f $X=9.3 $Y=1.295 $X2=0 $Y2=0
cc_345 N_A_c_216_n N_Y_c_775_n 0.0321248f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_346 N_A_M1033_g N_Y_c_786_n 6.94171e-19 $X=9.265 $Y=2.465 $X2=0 $Y2=0
cc_347 N_A_M1034_g N_Y_c_786_n 6.9407e-19 $X=9.695 $Y=2.465 $X2=0 $Y2=0
cc_348 N_A_c_206_n N_Y_c_786_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_349 N_A_c_215_n N_Y_c_786_n 0.0122997f $X=9.3 $Y=1.295 $X2=0 $Y2=0
cc_350 N_A_c_216_n N_Y_c_786_n 9.17266e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_351 N_A_M1036_g N_Y_c_787_n 6.94851e-19 $X=10.125 $Y=2.465 $X2=0 $Y2=0
cc_352 N_A_M1038_g N_Y_c_787_n 6.94851e-19 $X=10.555 $Y=2.465 $X2=0 $Y2=0
cc_353 N_A_c_206_n N_Y_c_787_n 7.70873e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_354 N_A_c_215_n N_Y_c_787_n 0.0124345f $X=9.3 $Y=1.295 $X2=0 $Y2=0
cc_355 N_A_c_216_n N_Y_c_787_n 9.35394e-19 $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_356 N_A_M1000_g N_Y_c_873_n 0.00197372f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_357 N_A_M1001_g N_Y_c_873_n 0.0078518f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_358 N_A_M1002_g N_Y_c_873_n 0.0078518f $X=1.525 $Y=2.465 $X2=0 $Y2=0
cc_359 N_A_M1003_g N_Y_c_873_n 0.0078518f $X=1.955 $Y=2.465 $X2=0 $Y2=0
cc_360 N_A_M1004_g N_Y_c_873_n 0.00875712f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_361 N_A_M1005_g N_Y_c_873_n 0.00875712f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_362 N_A_M1009_g N_Y_c_873_n 0.00875712f $X=3.245 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A_M1013_g N_Y_c_873_n 0.00875712f $X=3.675 $Y=2.465 $X2=0 $Y2=0
cc_364 N_A_M1014_g N_Y_c_873_n 0.00875712f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_365 N_A_M1016_g N_Y_c_873_n 0.00875712f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_366 N_A_M1018_g N_Y_c_873_n 0.00875712f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_367 N_A_M1019_g N_Y_c_873_n 0.00875712f $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_368 N_A_M1020_g N_Y_c_873_n 0.00875712f $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_369 N_A_M1021_g N_Y_c_873_n 0.00875712f $X=6.255 $Y=2.465 $X2=0 $Y2=0
cc_370 N_A_M1023_g N_Y_c_873_n 0.00875712f $X=6.685 $Y=2.465 $X2=0 $Y2=0
cc_371 N_A_M1024_g N_Y_c_873_n 0.00875712f $X=7.115 $Y=2.465 $X2=0 $Y2=0
cc_372 N_A_M1025_g N_Y_c_873_n 0.00875712f $X=7.545 $Y=2.465 $X2=0 $Y2=0
cc_373 N_A_M1026_g N_Y_c_873_n 0.00875712f $X=7.975 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A_M1027_g N_Y_c_873_n 0.00875712f $X=8.405 $Y=2.465 $X2=0 $Y2=0
cc_375 N_A_M1030_g N_Y_c_873_n 0.00875712f $X=8.835 $Y=2.465 $X2=0 $Y2=0
cc_376 N_A_M1033_g N_Y_c_873_n 0.0078518f $X=9.265 $Y=2.465 $X2=0 $Y2=0
cc_377 N_A_M1034_g N_Y_c_873_n 0.0078518f $X=9.695 $Y=2.465 $X2=0 $Y2=0
cc_378 N_A_M1036_g N_Y_c_873_n 0.0078518f $X=10.125 $Y=2.465 $X2=0 $Y2=0
cc_379 N_A_M1038_g N_Y_c_873_n 0.00197372f $X=10.555 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A_c_207_n N_Y_c_873_n 0.0182758f $X=0.86 $Y=1.295 $X2=0 $Y2=0
cc_381 N_A_c_208_n N_Y_c_873_n 0.0011189f $X=3.035 $Y=1.295 $X2=0 $Y2=0
cc_382 N_A_c_209_n N_Y_c_873_n 0.0011189f $X=3.89 $Y=1.295 $X2=0 $Y2=0
cc_383 N_A_c_210_n N_Y_c_873_n 0.0011189f $X=4.755 $Y=1.295 $X2=0 $Y2=0
cc_384 N_A_c_211_n N_Y_c_873_n 0.0011189f $X=5.61 $Y=1.295 $X2=0 $Y2=0
cc_385 N_A_c_212_n N_Y_c_873_n 0.0011189f $X=6.475 $Y=1.295 $X2=0 $Y2=0
cc_386 N_A_c_213_n N_Y_c_873_n 0.0011189f $X=7.335 $Y=1.295 $X2=0 $Y2=0
cc_387 N_A_c_214_n N_Y_c_873_n 0.0011189f $X=8.195 $Y=1.295 $X2=0 $Y2=0
cc_388 N_A_c_215_n N_Y_c_873_n 0.0180332f $X=9.3 $Y=1.295 $X2=0 $Y2=0
cc_389 N_A_c_216_n N_Y_c_873_n 0.436174f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_390 N_A_M1006_g N_VGND_c_1005_n 0.00411636f $X=2.385 $Y=0.56 $X2=0 $Y2=0
cc_391 N_A_c_206_n N_VGND_c_1005_n 0.00129197f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_392 N_A_c_207_n N_VGND_c_1005_n 0.00921969f $X=0.86 $Y=1.295 $X2=0 $Y2=0
cc_393 N_A_c_216_n N_VGND_c_1005_n 0.00208709f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_394 N_A_M1007_g N_VGND_c_1006_n 0.00187708f $X=2.815 $Y=0.56 $X2=0 $Y2=0
cc_395 N_A_M1008_g N_VGND_c_1006_n 0.00189723f $X=3.245 $Y=0.56 $X2=0 $Y2=0
cc_396 N_A_c_206_n N_VGND_c_1006_n 5.50763e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_397 N_A_c_208_n N_VGND_c_1006_n 0.00837841f $X=3.035 $Y=1.295 $X2=0 $Y2=0
cc_398 N_A_c_216_n N_VGND_c_1006_n 0.00204815f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_399 N_A_M1010_g N_VGND_c_1007_n 0.00187708f $X=3.675 $Y=0.56 $X2=0 $Y2=0
cc_400 N_A_M1011_g N_VGND_c_1007_n 0.00189723f $X=4.105 $Y=0.56 $X2=0 $Y2=0
cc_401 N_A_c_206_n N_VGND_c_1007_n 5.50763e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_402 N_A_c_209_n N_VGND_c_1007_n 0.00837841f $X=3.89 $Y=1.295 $X2=0 $Y2=0
cc_403 N_A_c_216_n N_VGND_c_1007_n 0.00204815f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_404 N_A_M1012_g N_VGND_c_1008_n 0.00187708f $X=4.535 $Y=0.56 $X2=0 $Y2=0
cc_405 N_A_M1015_g N_VGND_c_1008_n 0.00189723f $X=4.965 $Y=0.56 $X2=0 $Y2=0
cc_406 N_A_c_206_n N_VGND_c_1008_n 5.50763e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_407 N_A_c_210_n N_VGND_c_1008_n 0.00837841f $X=4.755 $Y=1.295 $X2=0 $Y2=0
cc_408 N_A_c_216_n N_VGND_c_1008_n 0.00204815f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_409 N_A_M1015_g N_VGND_c_1009_n 0.00478016f $X=4.965 $Y=0.56 $X2=0 $Y2=0
cc_410 N_A_M1017_g N_VGND_c_1009_n 0.00478016f $X=5.395 $Y=0.56 $X2=0 $Y2=0
cc_411 N_A_M1017_g N_VGND_c_1010_n 0.00187708f $X=5.395 $Y=0.56 $X2=0 $Y2=0
cc_412 N_A_M1022_g N_VGND_c_1010_n 0.00189723f $X=5.825 $Y=0.56 $X2=0 $Y2=0
cc_413 N_A_c_206_n N_VGND_c_1010_n 5.50763e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_414 N_A_c_211_n N_VGND_c_1010_n 0.00837841f $X=5.61 $Y=1.295 $X2=0 $Y2=0
cc_415 N_A_c_216_n N_VGND_c_1010_n 0.00204815f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_416 N_A_M1028_g N_VGND_c_1011_n 0.00187708f $X=6.255 $Y=0.56 $X2=0 $Y2=0
cc_417 N_A_M1029_g N_VGND_c_1011_n 0.00189723f $X=6.685 $Y=0.56 $X2=0 $Y2=0
cc_418 N_A_c_206_n N_VGND_c_1011_n 5.50763e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_419 N_A_c_212_n N_VGND_c_1011_n 0.00837841f $X=6.475 $Y=1.295 $X2=0 $Y2=0
cc_420 N_A_c_216_n N_VGND_c_1011_n 0.00204815f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_421 N_A_M1031_g N_VGND_c_1012_n 0.00187708f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_422 N_A_M1032_g N_VGND_c_1012_n 0.00189723f $X=7.545 $Y=0.56 $X2=0 $Y2=0
cc_423 N_A_c_206_n N_VGND_c_1012_n 5.50763e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_424 N_A_c_213_n N_VGND_c_1012_n 0.00837841f $X=7.335 $Y=1.295 $X2=0 $Y2=0
cc_425 N_A_c_216_n N_VGND_c_1012_n 0.00204815f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_426 N_A_M1035_g N_VGND_c_1013_n 0.00187708f $X=7.975 $Y=0.56 $X2=0 $Y2=0
cc_427 N_A_M1037_g N_VGND_c_1013_n 0.00189723f $X=8.405 $Y=0.56 $X2=0 $Y2=0
cc_428 N_A_c_206_n N_VGND_c_1013_n 5.50763e-19 $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_429 N_A_c_214_n N_VGND_c_1013_n 0.00837841f $X=8.195 $Y=1.295 $X2=0 $Y2=0
cc_430 N_A_c_216_n N_VGND_c_1013_n 0.00204815f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_431 N_A_M1039_g N_VGND_c_1014_n 0.00408131f $X=8.835 $Y=0.56 $X2=0 $Y2=0
cc_432 N_A_c_206_n N_VGND_c_1014_n 0.00128203f $X=10.555 $Y=1.46 $X2=0 $Y2=0
cc_433 N_A_c_215_n N_VGND_c_1014_n 0.00910469f $X=9.3 $Y=1.295 $X2=0 $Y2=0
cc_434 N_A_c_216_n N_VGND_c_1014_n 0.00204815f $X=10.38 $Y=1.295 $X2=0 $Y2=0
cc_435 N_A_M1006_g N_VGND_c_1015_n 0.00478016f $X=2.385 $Y=0.56 $X2=0 $Y2=0
cc_436 N_A_M1007_g N_VGND_c_1015_n 0.00478016f $X=2.815 $Y=0.56 $X2=0 $Y2=0
cc_437 N_A_M1008_g N_VGND_c_1017_n 0.00478016f $X=3.245 $Y=0.56 $X2=0 $Y2=0
cc_438 N_A_M1010_g N_VGND_c_1017_n 0.00478016f $X=3.675 $Y=0.56 $X2=0 $Y2=0
cc_439 N_A_M1011_g N_VGND_c_1019_n 0.00478016f $X=4.105 $Y=0.56 $X2=0 $Y2=0
cc_440 N_A_M1012_g N_VGND_c_1019_n 0.00478016f $X=4.535 $Y=0.56 $X2=0 $Y2=0
cc_441 N_A_M1029_g N_VGND_c_1021_n 0.00478016f $X=6.685 $Y=0.56 $X2=0 $Y2=0
cc_442 N_A_M1031_g N_VGND_c_1021_n 0.00478016f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_443 N_A_M1032_g N_VGND_c_1023_n 0.00478016f $X=7.545 $Y=0.56 $X2=0 $Y2=0
cc_444 N_A_M1035_g N_VGND_c_1023_n 0.00478016f $X=7.975 $Y=0.56 $X2=0 $Y2=0
cc_445 N_A_M1037_g N_VGND_c_1025_n 0.00478016f $X=8.405 $Y=0.56 $X2=0 $Y2=0
cc_446 N_A_M1039_g N_VGND_c_1025_n 0.00478016f $X=8.835 $Y=0.56 $X2=0 $Y2=0
cc_447 N_A_M1022_g N_VGND_c_1028_n 0.00478016f $X=5.825 $Y=0.56 $X2=0 $Y2=0
cc_448 N_A_M1028_g N_VGND_c_1028_n 0.00478016f $X=6.255 $Y=0.56 $X2=0 $Y2=0
cc_449 N_A_M1006_g N_VGND_c_1030_n 0.0095996f $X=2.385 $Y=0.56 $X2=0 $Y2=0
cc_450 N_A_M1007_g N_VGND_c_1030_n 0.00935526f $X=2.815 $Y=0.56 $X2=0 $Y2=0
cc_451 N_A_M1008_g N_VGND_c_1030_n 0.00934966f $X=3.245 $Y=0.56 $X2=0 $Y2=0
cc_452 N_A_M1010_g N_VGND_c_1030_n 0.00935526f $X=3.675 $Y=0.56 $X2=0 $Y2=0
cc_453 N_A_M1011_g N_VGND_c_1030_n 0.00934966f $X=4.105 $Y=0.56 $X2=0 $Y2=0
cc_454 N_A_M1012_g N_VGND_c_1030_n 0.00935526f $X=4.535 $Y=0.56 $X2=0 $Y2=0
cc_455 N_A_M1015_g N_VGND_c_1030_n 0.00934966f $X=4.965 $Y=0.56 $X2=0 $Y2=0
cc_456 N_A_M1017_g N_VGND_c_1030_n 0.00935526f $X=5.395 $Y=0.56 $X2=0 $Y2=0
cc_457 N_A_M1022_g N_VGND_c_1030_n 0.00934966f $X=5.825 $Y=0.56 $X2=0 $Y2=0
cc_458 N_A_M1028_g N_VGND_c_1030_n 0.00935526f $X=6.255 $Y=0.56 $X2=0 $Y2=0
cc_459 N_A_M1029_g N_VGND_c_1030_n 0.00934966f $X=6.685 $Y=0.56 $X2=0 $Y2=0
cc_460 N_A_M1031_g N_VGND_c_1030_n 0.00935526f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_461 N_A_M1032_g N_VGND_c_1030_n 0.00934966f $X=7.545 $Y=0.56 $X2=0 $Y2=0
cc_462 N_A_M1035_g N_VGND_c_1030_n 0.00935526f $X=7.975 $Y=0.56 $X2=0 $Y2=0
cc_463 N_A_M1037_g N_VGND_c_1030_n 0.00934966f $X=8.405 $Y=0.56 $X2=0 $Y2=0
cc_464 N_A_M1039_g N_VGND_c_1030_n 0.0096052f $X=8.835 $Y=0.56 $X2=0 $Y2=0
cc_465 N_VPWR_c_540_n N_Y_M1000_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_466 N_VPWR_c_540_n N_Y_M1002_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_467 N_VPWR_c_540_n N_Y_M1004_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_468 N_VPWR_c_540_n N_Y_M1009_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_469 N_VPWR_c_540_n N_Y_M1014_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_470 N_VPWR_c_540_n N_Y_M1018_d 0.00293778f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_471 N_VPWR_c_540_n N_Y_M1020_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_472 N_VPWR_c_540_n N_Y_M1023_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_473 N_VPWR_c_540_n N_Y_M1025_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_474 N_VPWR_c_540_n N_Y_M1027_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_475 N_VPWR_c_540_n N_Y_M1033_d 0.00311159f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_476 N_VPWR_c_540_n N_Y_M1036_d 0.00293778f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_c_547_n N_Y_c_796_n 0.00820394f $X=4.75 $Y=2.04 $X2=0 $Y2=0
cc_478 N_VPWR_c_549_n N_Y_c_796_n 0.00820394f $X=5.61 $Y=2.04 $X2=0 $Y2=0
cc_479 N_VPWR_c_542_n N_Y_c_777_n 0.0131021f $X=1.18 $Y=3.33 $X2=0 $Y2=0
cc_480 N_VPWR_c_543_n N_Y_c_777_n 0.0082193f $X=1.31 $Y=2.04 $X2=0 $Y2=0
cc_481 N_VPWR_c_540_n N_Y_c_777_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_482 N_VPWR_c_543_n N_Y_c_778_n 0.0079844f $X=1.31 $Y=2.04 $X2=0 $Y2=0
cc_483 N_VPWR_c_544_n N_Y_c_778_n 0.0082193f $X=2.17 $Y=2.04 $X2=0 $Y2=0
cc_484 N_VPWR_c_572_n N_Y_c_778_n 0.0131021f $X=2.04 $Y=3.33 $X2=0 $Y2=0
cc_485 N_VPWR_c_540_n N_Y_c_778_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_486 N_VPWR_c_544_n N_Y_c_769_n 0.0079844f $X=2.17 $Y=2.04 $X2=0 $Y2=0
cc_487 N_VPWR_c_545_n N_Y_c_769_n 0.0082193f $X=3.03 $Y=2.04 $X2=0 $Y2=0
cc_488 N_VPWR_c_560_n N_Y_c_769_n 0.0131021f $X=2.9 $Y=3.33 $X2=0 $Y2=0
cc_489 N_VPWR_c_540_n N_Y_c_769_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_490 N_VPWR_c_545_n N_Y_c_770_n 0.0079844f $X=3.03 $Y=2.04 $X2=0 $Y2=0
cc_491 N_VPWR_c_546_n N_Y_c_770_n 0.0082193f $X=3.89 $Y=2.04 $X2=0 $Y2=0
cc_492 N_VPWR_c_562_n N_Y_c_770_n 0.0131021f $X=3.76 $Y=3.33 $X2=0 $Y2=0
cc_493 N_VPWR_c_540_n N_Y_c_770_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_494 N_VPWR_c_546_n N_Y_c_771_n 0.0079844f $X=3.89 $Y=2.04 $X2=0 $Y2=0
cc_495 N_VPWR_c_547_n N_Y_c_771_n 0.0082193f $X=4.75 $Y=2.04 $X2=0 $Y2=0
cc_496 N_VPWR_c_564_n N_Y_c_771_n 0.0131021f $X=4.62 $Y=3.33 $X2=0 $Y2=0
cc_497 N_VPWR_c_540_n N_Y_c_771_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_498 N_VPWR_c_548_n N_Y_c_940_n 0.0132609f $X=5.48 $Y=3.33 $X2=0 $Y2=0
cc_499 N_VPWR_c_540_n N_Y_c_940_n 0.00993371f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_500 N_VPWR_c_549_n N_Y_c_772_n 0.0079844f $X=5.61 $Y=2.04 $X2=0 $Y2=0
cc_501 N_VPWR_c_550_n N_Y_c_772_n 0.0082193f $X=6.47 $Y=2.04 $X2=0 $Y2=0
cc_502 N_VPWR_c_573_n N_Y_c_772_n 0.0131021f $X=6.34 $Y=3.33 $X2=0 $Y2=0
cc_503 N_VPWR_c_540_n N_Y_c_772_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_504 N_VPWR_c_550_n N_Y_c_773_n 0.0079844f $X=6.47 $Y=2.04 $X2=0 $Y2=0
cc_505 N_VPWR_c_551_n N_Y_c_773_n 0.0082193f $X=7.33 $Y=2.04 $X2=0 $Y2=0
cc_506 N_VPWR_c_566_n N_Y_c_773_n 0.0131021f $X=7.2 $Y=3.33 $X2=0 $Y2=0
cc_507 N_VPWR_c_540_n N_Y_c_773_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_508 N_VPWR_c_551_n N_Y_c_774_n 0.0079844f $X=7.33 $Y=2.04 $X2=0 $Y2=0
cc_509 N_VPWR_c_552_n N_Y_c_774_n 0.0082193f $X=8.19 $Y=2.04 $X2=0 $Y2=0
cc_510 N_VPWR_c_568_n N_Y_c_774_n 0.0131021f $X=8.06 $Y=3.33 $X2=0 $Y2=0
cc_511 N_VPWR_c_540_n N_Y_c_774_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_512 N_VPWR_c_552_n N_Y_c_775_n 0.0079844f $X=8.19 $Y=2.04 $X2=0 $Y2=0
cc_513 N_VPWR_c_553_n N_Y_c_775_n 0.0082193f $X=9.05 $Y=2.04 $X2=0 $Y2=0
cc_514 N_VPWR_c_570_n N_Y_c_775_n 0.0131021f $X=8.92 $Y=3.33 $X2=0 $Y2=0
cc_515 N_VPWR_c_540_n N_Y_c_775_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_516 N_VPWR_c_553_n N_Y_c_786_n 0.0079844f $X=9.05 $Y=2.04 $X2=0 $Y2=0
cc_517 N_VPWR_c_554_n N_Y_c_786_n 0.0131021f $X=9.78 $Y=3.33 $X2=0 $Y2=0
cc_518 N_VPWR_c_555_n N_Y_c_786_n 0.0082193f $X=9.91 $Y=2.04 $X2=0 $Y2=0
cc_519 N_VPWR_c_540_n N_Y_c_786_n 0.0097412f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_520 N_VPWR_c_555_n N_Y_c_787_n 0.00822181f $X=9.91 $Y=2.04 $X2=0 $Y2=0
cc_521 N_VPWR_c_574_n N_Y_c_787_n 0.0132609f $X=10.64 $Y=3.33 $X2=0 $Y2=0
cc_522 N_VPWR_c_540_n N_Y_c_787_n 0.00993371f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_523 N_VPWR_M1001_s N_Y_c_873_n 7.61922e-19 $X=1.17 $Y=1.835 $X2=0 $Y2=0
cc_524 N_VPWR_M1003_s N_Y_c_873_n 7.69148e-19 $X=2.03 $Y=1.835 $X2=0 $Y2=0
cc_525 N_VPWR_M1005_s N_Y_c_873_n 8.17926e-19 $X=2.89 $Y=1.835 $X2=0 $Y2=0
cc_526 N_VPWR_M1013_s N_Y_c_873_n 8.17926e-19 $X=3.75 $Y=1.835 $X2=0 $Y2=0
cc_527 N_VPWR_M1016_s N_Y_c_873_n 8.17926e-19 $X=4.61 $Y=1.835 $X2=0 $Y2=0
cc_528 N_VPWR_M1019_s N_Y_c_873_n 8.17926e-19 $X=5.47 $Y=1.835 $X2=0 $Y2=0
cc_529 N_VPWR_M1021_s N_Y_c_873_n 8.17926e-19 $X=6.33 $Y=1.835 $X2=0 $Y2=0
cc_530 N_VPWR_M1024_s N_Y_c_873_n 8.17926e-19 $X=7.19 $Y=1.835 $X2=0 $Y2=0
cc_531 N_VPWR_M1026_s N_Y_c_873_n 8.17926e-19 $X=8.05 $Y=1.835 $X2=0 $Y2=0
cc_532 N_VPWR_M1030_s N_Y_c_873_n 8.10699e-19 $X=8.91 $Y=1.835 $X2=0 $Y2=0
cc_533 N_VPWR_M1034_s N_Y_c_873_n 7.61922e-19 $X=9.77 $Y=1.835 $X2=0 $Y2=0
cc_534 N_VPWR_c_541_n N_Y_c_873_n 0.00691811f $X=0.45 $Y=2.04 $X2=0 $Y2=0
cc_535 N_VPWR_c_543_n N_Y_c_873_n 0.0296667f $X=1.31 $Y=2.04 $X2=0 $Y2=0
cc_536 N_VPWR_c_544_n N_Y_c_873_n 0.0296667f $X=2.17 $Y=2.04 $X2=0 $Y2=0
cc_537 N_VPWR_c_545_n N_Y_c_873_n 0.0296667f $X=3.03 $Y=2.04 $X2=0 $Y2=0
cc_538 N_VPWR_c_546_n N_Y_c_873_n 0.0296667f $X=3.89 $Y=2.04 $X2=0 $Y2=0
cc_539 N_VPWR_c_547_n N_Y_c_873_n 0.0296101f $X=4.75 $Y=2.04 $X2=0 $Y2=0
cc_540 N_VPWR_c_549_n N_Y_c_873_n 0.0296667f $X=5.61 $Y=2.04 $X2=0 $Y2=0
cc_541 N_VPWR_c_550_n N_Y_c_873_n 0.0296667f $X=6.47 $Y=2.04 $X2=0 $Y2=0
cc_542 N_VPWR_c_551_n N_Y_c_873_n 0.0296667f $X=7.33 $Y=2.04 $X2=0 $Y2=0
cc_543 N_VPWR_c_552_n N_Y_c_873_n 0.0296667f $X=8.19 $Y=2.04 $X2=0 $Y2=0
cc_544 N_VPWR_c_553_n N_Y_c_873_n 0.0296667f $X=9.05 $Y=2.04 $X2=0 $Y2=0
cc_545 N_VPWR_c_555_n N_Y_c_873_n 0.0296101f $X=9.91 $Y=2.04 $X2=0 $Y2=0
cc_546 N_VPWR_c_557_n N_Y_c_873_n 0.00689488f $X=10.77 $Y=2.04 $X2=0 $Y2=0
cc_547 N_Y_c_768_n N_VGND_c_1009_n 0.00778443f $X=5.18 $Y=0.56 $X2=0 $Y2=0
cc_548 N_Y_c_769_n N_VGND_c_1015_n 0.00778443f $X=2.6 $Y=0.56 $X2=0 $Y2=0
cc_549 N_Y_c_770_n N_VGND_c_1017_n 0.00778443f $X=3.46 $Y=0.56 $X2=0 $Y2=0
cc_550 N_Y_c_771_n N_VGND_c_1019_n 0.00778443f $X=4.32 $Y=0.56 $X2=0 $Y2=0
cc_551 N_Y_c_773_n N_VGND_c_1021_n 0.00778443f $X=6.9 $Y=0.56 $X2=0 $Y2=0
cc_552 N_Y_c_774_n N_VGND_c_1023_n 0.00778443f $X=7.76 $Y=0.56 $X2=0 $Y2=0
cc_553 N_Y_c_775_n N_VGND_c_1025_n 0.00778443f $X=8.62 $Y=0.56 $X2=0 $Y2=0
cc_554 N_Y_c_772_n N_VGND_c_1028_n 0.00778443f $X=6.04 $Y=0.56 $X2=0 $Y2=0
cc_555 N_Y_c_768_n N_VGND_c_1030_n 0.00908624f $X=5.18 $Y=0.56 $X2=0 $Y2=0
cc_556 N_Y_c_769_n N_VGND_c_1030_n 0.00908624f $X=2.6 $Y=0.56 $X2=0 $Y2=0
cc_557 N_Y_c_770_n N_VGND_c_1030_n 0.00908624f $X=3.46 $Y=0.56 $X2=0 $Y2=0
cc_558 N_Y_c_771_n N_VGND_c_1030_n 0.00908624f $X=4.32 $Y=0.56 $X2=0 $Y2=0
cc_559 N_Y_c_772_n N_VGND_c_1030_n 0.00908624f $X=6.04 $Y=0.56 $X2=0 $Y2=0
cc_560 N_Y_c_773_n N_VGND_c_1030_n 0.00908624f $X=6.9 $Y=0.56 $X2=0 $Y2=0
cc_561 N_Y_c_774_n N_VGND_c_1030_n 0.00908624f $X=7.76 $Y=0.56 $X2=0 $Y2=0
cc_562 N_Y_c_775_n N_VGND_c_1030_n 0.00908624f $X=8.62 $Y=0.56 $X2=0 $Y2=0
