* File: sky130_fd_sc_lp__o221ai_1.spice
* Created: Wed Sep  2 10:19:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221ai_1.pex.spice"
.subckt sky130_fd_sc_lp__o221ai_1  VNB VPB C1 B1 B2 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1002 N_A_114_47#_M1002_d N_C1_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_A_114_47#_M1008_d N_B1_M1008_g N_A_221_49#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1638 AS=0.2226 PD=1.23 PS=2.21 NRD=7.848 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1001 N_A_221_49#_M1001_d N_B2_M1001_g N_A_114_47#_M1008_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1638 PD=1.12 PS=1.23 NRD=0 NRS=7.848 M=1 R=5.6
+ SA=75000.7 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_221_49#_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=4.284 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1003 N_A_221_49#_M1003_d N_A1_M1003_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1344 PD=2.21 PS=1.16 NRD=0 NRS=1.428 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_C1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.3339 PD=1.88 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1007 A_304_367# N_B1_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3906 PD=1.47 PS=1.88 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1009 N_Y_M1009_d N_B2_M1009_g A_304_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.3591
+ AS=0.1323 PD=1.83 PS=1.47 NRD=21.0987 NRS=7.8012 M=1 R=8.4 SA=75001.3
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1004 A_520_367# N_A2_M1004_g N_Y_M1009_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.3591 PD=1.47 PS=1.83 NRD=7.8012 NRS=24.231 M=1 R=8.4 SA=75002 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g A_520_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o221ai_1.pxi.spice"
*
.ends
*
*
