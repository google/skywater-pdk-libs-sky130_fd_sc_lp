* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxbp_lp2 D GATE VGND VNB VPB VPWR Q Q_N
X0 a_978_393# a_934_29# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VPWR a_784_55# a_934_29# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VGND GATE a_278_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_461_55# a_278_409# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_886_55# a_934_29# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1860_92# a_1662_57# Q_N VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_27_57# a_717_393# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 Q a_934_29# a_1432_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR GATE a_278_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VPWR a_934_29# a_1662_57# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_1162_55# a_784_55# a_934_29# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1432_57# a_934_29# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_717_393# a_278_409# a_784_55# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 VGND a_934_29# a_1590_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_706_55# a_461_55# a_784_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_278_57# GATE a_278_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 Q a_934_29# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 VGND a_1662_57# a_1860_92# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_548_55# a_278_409# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_784_55# a_278_409# a_886_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_461_55# a_278_409# a_548_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VGND a_784_55# a_1162_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_114_57# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_27_57# D a_114_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VGND a_27_57# a_706_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_784_55# a_461_55# a_978_393# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X26 a_27_57# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 VPWR a_1662_57# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X28 a_1590_57# a_934_29# a_1662_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
