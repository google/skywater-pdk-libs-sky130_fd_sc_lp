* NGSPICE file created from sky130_fd_sc_lp__or2_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or2_lp A B VGND VNB VPB VPWR X
M1000 a_196_114# B a_154_468# VPB phighvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1001 a_196_114# A a_118_114# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.008e+11p ps=1.32e+06u
M1002 a_282_114# B a_196_114# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1003 X a_196_114# a_484_114# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1004 a_118_114# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.297e+11p ps=3.25e+06u
M1005 a_484_114# a_196_114# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_154_468# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.82e+06u
M1007 X a_196_114# a_435_490# VPB phighvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1008 VGND B a_282_114# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_435_490# a_196_114# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

