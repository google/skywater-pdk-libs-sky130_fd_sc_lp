* File: sky130_fd_sc_lp__a2111o_2.spice
* Created: Wed Sep  2 09:16:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111o_2.pex.spice"
.subckt sky130_fd_sc_lp__a2111o_2  VNB VPB D1 C1 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1003 N_X_M1003_d N_A_86_275#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1006 N_X_M1003_d N_A_86_275#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3759 PD=1.12 PS=1.735 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_86_275#_M1004_d N_D1_M1004_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3759 PD=1.12 PS=1.735 NRD=0 NRS=0 M=1 R=5.6 SA=75001.7
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_C1_M1009_g N_A_86_275#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1575 AS=0.1176 PD=1.215 PS=1.12 NRD=7.14 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1000 N_A_86_275#_M1000_d N_B1_M1000_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1407 AS=0.1575 PD=1.175 PS=1.215 NRD=0 NRS=6.42 M=1 R=5.6 SA=75002.6
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1013 A_715_49# N_A1_M1013_g N_A_86_275#_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1407 PD=1.23 PS=1.175 NRD=19.992 NRS=7.848 M=1 R=5.6 SA=75003.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g A_715_49# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6 SA=75003.6 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1005 N_X_M1005_d N_A_86_275#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_X_M1005_d N_A_86_275#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1008 A_427_367# N_D1_M1008_g N_A_86_275#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1011 A_499_367# N_C1_M1011_g A_427_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1001 N_A_607_367#_M1001_d N_B1_M1001_g A_499_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=9.3772 NRS=21.8867 M=1 R=8.4
+ SA=75001.1 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_607_367#_M1001_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=8.5892 NRS=7.8012 M=1 R=8.4
+ SA=75001.6 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1012 N_A_607_367#_M1012_d N_A2_M1012_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=8.5892 M=1 R=8.4
+ SA=75002.2 SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__a2111o_2.pxi.spice"
*
.ends
*
*
