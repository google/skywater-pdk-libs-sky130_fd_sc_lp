* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__ha_1 A B VGND VNB VPB VPWR COUT SUM
X0 a_401_428# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR B a_223_320# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_80_30# a_223_320# a_307_62# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_307_62# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_223_320# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR a_223_320# a_80_30# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_223_320# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND A a_307_62# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 SUM a_80_30# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_223_320# B a_675_146# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_80_30# B a_401_428# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 SUM a_80_30# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_675_146# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_223_320# COUT VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
