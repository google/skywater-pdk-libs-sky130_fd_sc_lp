* File: sky130_fd_sc_lp__o311a_4.pxi.spice
* Created: Wed Sep  2 10:23:09 2020
* 
x_PM_SKY130_FD_SC_LP__O311A_4%A_81_23# N_A_81_23#_M1012_d N_A_81_23#_M1007_s
+ N_A_81_23#_M1010_d N_A_81_23#_M1004_s N_A_81_23#_M1000_g N_A_81_23#_M1003_g
+ N_A_81_23#_M1006_g N_A_81_23#_M1014_g N_A_81_23#_M1008_g N_A_81_23#_M1018_g
+ N_A_81_23#_M1021_g N_A_81_23#_M1024_g N_A_81_23#_c_204_p N_A_81_23#_c_134_n
+ N_A_81_23#_c_187_p N_A_81_23#_c_135_n N_A_81_23#_c_155_p N_A_81_23#_c_142_n
+ N_A_81_23#_c_136_n N_A_81_23#_c_194_p N_A_81_23#_c_144_n N_A_81_23#_c_145_n
+ N_A_81_23#_c_230_p N_A_81_23#_c_146_n N_A_81_23#_c_137_n
+ PM_SKY130_FD_SC_LP__O311A_4%A_81_23#
x_PM_SKY130_FD_SC_LP__O311A_4%C1 N_C1_M1007_g N_C1_c_260_n N_C1_M1012_g
+ N_C1_M1027_g N_C1_c_262_n N_C1_M1022_g C1 N_C1_c_264_n
+ PM_SKY130_FD_SC_LP__O311A_4%C1
x_PM_SKY130_FD_SC_LP__O311A_4%B1 N_B1_M1010_g N_B1_c_306_n N_B1_M1001_g
+ N_B1_M1025_g N_B1_c_308_n N_B1_M1009_g B1 N_B1_c_310_n
+ PM_SKY130_FD_SC_LP__O311A_4%B1
x_PM_SKY130_FD_SC_LP__O311A_4%A3 N_A3_M1004_g N_A3_c_349_n N_A3_M1015_g
+ N_A3_M1019_g N_A3_c_351_n N_A3_M1017_g N_A3_c_352_n N_A3_c_353_n A3 A3 A3 A3
+ PM_SKY130_FD_SC_LP__O311A_4%A3
x_PM_SKY130_FD_SC_LP__O311A_4%A2 N_A2_M1002_g N_A2_M1011_g N_A2_M1016_g
+ N_A2_M1026_g A2 A2 A2 N_A2_c_402_n PM_SKY130_FD_SC_LP__O311A_4%A2
x_PM_SKY130_FD_SC_LP__O311A_4%A1 N_A1_M1013_g N_A1_M1005_g N_A1_M1023_g
+ N_A1_M1020_g A1 A1 N_A1_c_458_n PM_SKY130_FD_SC_LP__O311A_4%A1
x_PM_SKY130_FD_SC_LP__O311A_4%VPWR N_VPWR_M1003_d N_VPWR_M1014_d N_VPWR_M1024_d
+ N_VPWR_M1027_d N_VPWR_M1025_s N_VPWR_M1005_s N_VPWR_c_494_n N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n
+ N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n VPWR
+ N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_493_n
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n
+ PM_SKY130_FD_SC_LP__O311A_4%VPWR
x_PM_SKY130_FD_SC_LP__O311A_4%X N_X_M1000_d N_X_M1008_d N_X_M1003_s N_X_M1018_s
+ N_X_c_602_n N_X_c_607_n N_X_c_608_n N_X_c_653_p N_X_c_603_n N_X_c_640_n
+ N_X_c_609_n N_X_c_652_p N_X_c_644_n N_X_c_604_n N_X_c_610_n X X N_X_c_605_n X
+ PM_SKY130_FD_SC_LP__O311A_4%X
x_PM_SKY130_FD_SC_LP__O311A_4%A_910_345# N_A_910_345#_M1004_d
+ N_A_910_345#_M1019_d N_A_910_345#_M1011_d N_A_910_345#_c_658_n
+ N_A_910_345#_c_659_n N_A_910_345#_c_660_n N_A_910_345#_c_661_n
+ N_A_910_345#_c_662_n N_A_910_345#_c_682_n N_A_910_345#_c_663_n
+ PM_SKY130_FD_SC_LP__O311A_4%A_910_345#
x_PM_SKY130_FD_SC_LP__O311A_4%A_1196_367# N_A_1196_367#_M1011_s
+ N_A_1196_367#_M1026_s N_A_1196_367#_M1020_d N_A_1196_367#_c_701_n
+ N_A_1196_367#_c_702_n N_A_1196_367#_c_706_n N_A_1196_367#_c_720_n
+ N_A_1196_367#_c_710_n N_A_1196_367#_c_703_n N_A_1196_367#_c_704_n
+ N_A_1196_367#_c_711_n PM_SKY130_FD_SC_LP__O311A_4%A_1196_367#
x_PM_SKY130_FD_SC_LP__O311A_4%VGND N_VGND_M1000_s N_VGND_M1006_s N_VGND_M1021_s
+ N_VGND_M1015_d N_VGND_M1002_d N_VGND_M1013_s N_VGND_c_733_n N_VGND_c_734_n
+ N_VGND_c_735_n N_VGND_c_736_n N_VGND_c_737_n N_VGND_c_738_n N_VGND_c_739_n
+ N_VGND_c_740_n VGND N_VGND_c_741_n N_VGND_c_742_n N_VGND_c_743_n
+ N_VGND_c_744_n N_VGND_c_745_n N_VGND_c_746_n N_VGND_c_747_n N_VGND_c_748_n
+ N_VGND_c_749_n N_VGND_c_750_n PM_SKY130_FD_SC_LP__O311A_4%VGND
x_PM_SKY130_FD_SC_LP__O311A_4%A_476_47# N_A_476_47#_M1012_s N_A_476_47#_M1022_s
+ N_A_476_47#_M1009_s N_A_476_47#_c_845_n N_A_476_47#_c_855_n
+ N_A_476_47#_c_856_n N_A_476_47#_c_866_n N_A_476_47#_c_846_n
+ PM_SKY130_FD_SC_LP__O311A_4%A_476_47#
x_PM_SKY130_FD_SC_LP__O311A_4%A_731_47# N_A_731_47#_M1001_d N_A_731_47#_M1015_s
+ N_A_731_47#_M1017_s N_A_731_47#_M1016_s N_A_731_47#_M1023_d
+ N_A_731_47#_c_876_n N_A_731_47#_c_877_n N_A_731_47#_c_892_n
+ N_A_731_47#_c_928_n N_A_731_47#_c_878_n N_A_731_47#_c_906_n
+ N_A_731_47#_c_879_n N_A_731_47#_c_880_n N_A_731_47#_c_884_n
+ N_A_731_47#_c_881_n N_A_731_47#_c_882_n N_A_731_47#_c_883_n
+ PM_SKY130_FD_SC_LP__O311A_4%A_731_47#
cc_1 VNB N_A_81_23#_M1000_g 0.0258992f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.665
cc_2 VNB N_A_81_23#_M1006_g 0.0213077f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.665
cc_3 VNB N_A_81_23#_M1008_g 0.0213292f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.665
cc_4 VNB N_A_81_23#_M1021_g 0.0277381f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=0.665
cc_5 VNB N_A_81_23#_c_134_n 0.00506167f $X=-0.19 $Y=-0.245 $X2=2.557 $Y2=1.405
cc_6 VNB N_A_81_23#_c_135_n 0.00309477f $X=-0.19 $Y=-0.245 $X2=2.795 $Y2=0.89
cc_7 VNB N_A_81_23#_c_136_n 0.00532838f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.79
cc_8 VNB N_A_81_23#_c_137_n 0.0965064f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=1.49
cc_9 VNB N_C1_M1007_g 0.00549113f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.835
cc_10 VNB N_C1_c_260_n 0.0200087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C1_M1027_g 0.00709761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C1_c_262_n 0.0164274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB C1 0.00437061f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.665
cc_14 VNB N_C1_c_264_n 0.0473265f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.325
cc_15 VNB N_B1_M1010_g 0.00436542f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.835
cc_16 VNB N_B1_c_306_n 0.0169694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_M1025_g 0.00635747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_308_n 0.0228862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB B1 0.00228955f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.665
cc_20 VNB N_B1_c_310_n 0.054779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A3_M1004_g 0.00233375f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.835
cc_22 VNB N_A3_c_349_n 0.0271196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A3_M1019_g 0.00176052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A3_c_351_n 0.0214434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A3_c_352_n 0.0417029f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.665
cc_26 VNB N_A3_c_353_n 0.0533735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A3 0.0179547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_M1002_g 0.0229513f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.835
cc_29 VNB N_A2_M1016_g 0.0229523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB A2 0.00734919f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_31 VNB N_A2_c_402_n 0.0328533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_M1013_g 0.0229349f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.835
cc_33 VNB N_A1_M1023_g 0.0306331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB A1 0.0171091f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_35 VNB N_A1_c_458_n 0.0369905f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_36 VNB N_VPWR_c_493_n 0.342803f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.49
cc_37 VNB N_X_c_602_n 9.73185e-19 $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.325
cc_38 VNB N_X_c_603_n 0.00670746f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.325
cc_39 VNB N_X_c_604_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=2.465
cc_40 VNB N_X_c_605_n 0.00918763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB X 0.0218909f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=1.49
cc_42 VNB N_VGND_c_733_n 0.010601f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_43 VNB N_VGND_c_734_n 0.0281524f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.325
cc_44 VNB N_VGND_c_735_n 4.82391e-19 $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.655
cc_45 VNB N_VGND_c_736_n 0.016264f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.325
cc_46 VNB N_VGND_c_737_n 3.08929e-19 $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.655
cc_47 VNB N_VGND_c_738_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.325
cc_48 VNB N_VGND_c_739_n 0.014949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_740_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=1.655
cc_50 VNB N_VGND_c_741_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_742_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=2.79 $Y2=1.98
cc_52 VNB N_VGND_c_743_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=2.935 $Y2=0.89
cc_53 VNB N_VGND_c_744_n 0.0177625f $X=-0.19 $Y=-0.245 $X2=3.725 $Y2=1.98
cc_54 VNB N_VGND_c_745_n 0.40227f $X=-0.19 $Y=-0.245 $X2=3.707 $Y2=2.91
cc_55 VNB N_VGND_c_746_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=5.122 $Y2=2.57
cc_56 VNB N_VGND_c_747_n 0.0676848f $X=-0.19 $Y=-0.245 $X2=3.707 $Y2=1.79
cc_57 VNB N_VGND_c_748_n 0.0162594f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.49
cc_58 VNB N_VGND_c_749_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.49
cc_59 VNB N_VGND_c_750_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.49
cc_60 VNB N_A_476_47#_c_845_n 0.00371693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_476_47#_c_846_n 0.00447166f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.665
cc_62 VNB N_A_731_47#_c_876_n 0.00735052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_731_47#_c_877_n 0.00611325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_731_47#_c_878_n 0.00901485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_731_47#_c_879_n 0.0190171f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=2.465
cc_66 VNB N_A_731_47#_c_880_n 0.0315826f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=0.665
cc_67 VNB N_A_731_47#_c_881_n 6.49321e-19 $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=2.465
cc_68 VNB N_A_731_47#_c_882_n 0.00387368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_731_47#_c_883_n 0.00178419f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.49
cc_70 VPB N_A_81_23#_M1003_g 0.0229319f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.465
cc_71 VPB N_A_81_23#_M1014_g 0.0188632f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.465
cc_72 VPB N_A_81_23#_M1018_g 0.0188558f $X=-0.19 $Y=1.655 $X2=1.715 $Y2=2.465
cc_73 VPB N_A_81_23#_M1024_g 0.0187985f $X=-0.19 $Y=1.655 $X2=2.145 $Y2=2.465
cc_74 VPB N_A_81_23#_c_142_n 0.00721189f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=1.79
cc_75 VPB N_A_81_23#_c_136_n 0.00452497f $X=-0.19 $Y=1.655 $X2=2.925 $Y2=1.79
cc_76 VPB N_A_81_23#_c_144_n 0.0187798f $X=-0.19 $Y=1.655 $X2=5.01 $Y2=1.79
cc_77 VPB N_A_81_23#_c_145_n 0.00203797f $X=-0.19 $Y=1.655 $X2=5.122 $Y2=1.875
cc_78 VPB N_A_81_23#_c_146_n 0.002093f $X=-0.19 $Y=1.655 $X2=3.707 $Y2=1.79
cc_79 VPB N_A_81_23#_c_137_n 0.0165201f $X=-0.19 $Y=1.655 $X2=2.145 $Y2=1.49
cc_80 VPB N_C1_M1007_g 0.0180918f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=1.835
cc_81 VPB N_C1_M1027_g 0.0196727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_B1_M1010_g 0.0196802f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=1.835
cc_83 VPB N_B1_M1025_g 0.0239519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A3_M1004_g 0.026762f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=1.835
cc_85 VPB N_A3_M1019_g 0.0237698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A2_M1011_g 0.0228913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A2_M1026_g 0.0182425f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.665
cc_88 VPB A2 0.0130168f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.465
cc_89 VPB N_A2_c_402_n 0.00492723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A1_M1005_g 0.0183636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A1_M1020_g 0.0240279f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.665
cc_92 VPB A1 0.0138655f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.465
cc_93 VPB N_A1_c_458_n 0.00492723f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.465
cc_94 VPB N_VPWR_c_494_n 0.0414999f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.325
cc_95 VPB N_VPWR_c_495_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.465
cc_96 VPB N_VPWR_c_496_n 3.16049e-19 $X=-0.19 $Y=1.655 $X2=1.715 $Y2=1.655
cc_97 VPB N_VPWR_c_497_n 0.0148832f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=1.325
cc_98 VPB N_VPWR_c_498_n 0.00431378f $X=-0.19 $Y=1.655 $X2=2.145 $Y2=1.655
cc_99 VPB N_VPWR_c_499_n 0.0126203f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.49
cc_100 VPB N_VPWR_c_500_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=2.557 $Y2=1.015
cc_101 VPB N_VPWR_c_501_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.81 $Y2=1.98
cc_102 VPB N_VPWR_c_502_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.79 $Y2=1.98
cc_103 VPB N_VPWR_c_503_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.81 $Y2=2.91
cc_104 VPB N_VPWR_c_504_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.79 $Y2=2.91
cc_105 VPB N_VPWR_c_505_n 0.0172587f $X=-0.19 $Y=1.655 $X2=2.935 $Y2=0.89
cc_106 VPB N_VPWR_c_506_n 0.0147711f $X=-0.19 $Y=1.655 $X2=3.82 $Y2=1.79
cc_107 VPB N_VPWR_c_507_n 0.0685841f $X=-0.19 $Y=1.655 $X2=2.557 $Y2=1.64
cc_108 VPB N_VPWR_c_508_n 0.0177625f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=1.49
cc_109 VPB N_VPWR_c_493_n 0.0806139f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=1.49
cc_110 VPB N_VPWR_c_510_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=1.49
cc_111 VPB N_VPWR_c_511_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_512_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_513_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_X_c_607_n 0.0088321f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.665
cc_115 VPB N_X_c_608_n 0.0197681f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_X_c_609_n 0.00507419f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=1.325
cc_117 VPB N_X_c_610_n 0.00144314f $X=-0.19 $Y=1.655 $X2=2.145 $Y2=2.465
cc_118 VPB X 0.00582661f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=1.49
cc_119 VPB N_A_910_345#_c_658_n 0.0080373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_910_345#_c_659_n 0.00205771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_910_345#_c_660_n 0.00404106f $X=-0.19 $Y=1.655 $X2=0.855
+ $Y2=1.655
cc_122 VPB N_A_910_345#_c_661_n 0.0150943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_910_345#_c_662_n 0.0132763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_910_345#_c_663_n 0.00241061f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=0.665
cc_125 VPB N_A_1196_367#_c_701_n 0.00203846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_1196_367#_c_702_n 0.00663726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_1196_367#_c_703_n 0.0075508f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.665
cc_128 VPB N_A_1196_367#_c_704_n 0.0369431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 N_A_81_23#_M1024_g N_C1_M1007_g 0.0163861f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A_81_23#_c_136_n N_C1_M1007_g 0.0186809f $X=2.925 $Y=1.79 $X2=0 $Y2=0
cc_131 N_A_81_23#_c_134_n N_C1_c_260_n 0.00736922f $X=2.557 $Y=1.405 $X2=0 $Y2=0
cc_132 N_A_81_23#_c_135_n N_C1_c_260_n 0.0107825f $X=2.795 $Y=0.89 $X2=0 $Y2=0
cc_133 N_A_81_23#_c_142_n N_C1_M1027_g 0.0159635f $X=3.595 $Y=1.79 $X2=0 $Y2=0
cc_134 N_A_81_23#_c_136_n N_C1_M1027_g 0.005042f $X=2.925 $Y=1.79 $X2=0 $Y2=0
cc_135 N_A_81_23#_c_134_n N_C1_c_262_n 6.79588e-19 $X=2.557 $Y=1.405 $X2=0 $Y2=0
cc_136 N_A_81_23#_c_155_p N_C1_c_262_n 0.00319283f $X=2.935 $Y=0.88 $X2=0 $Y2=0
cc_137 N_A_81_23#_c_134_n C1 0.016057f $X=2.557 $Y=1.405 $X2=0 $Y2=0
cc_138 N_A_81_23#_c_155_p C1 0.00758217f $X=2.935 $Y=0.88 $X2=0 $Y2=0
cc_139 N_A_81_23#_c_142_n C1 0.021285f $X=3.595 $Y=1.79 $X2=0 $Y2=0
cc_140 N_A_81_23#_c_136_n C1 0.00951341f $X=2.925 $Y=1.79 $X2=0 $Y2=0
cc_141 N_A_81_23#_c_134_n N_C1_c_264_n 0.0140114f $X=2.557 $Y=1.405 $X2=0 $Y2=0
cc_142 N_A_81_23#_c_155_p N_C1_c_264_n 0.00399944f $X=2.935 $Y=0.88 $X2=0 $Y2=0
cc_143 N_A_81_23#_c_142_n N_C1_c_264_n 9.96329e-19 $X=3.595 $Y=1.79 $X2=0 $Y2=0
cc_144 N_A_81_23#_c_136_n N_C1_c_264_n 0.00999574f $X=2.925 $Y=1.79 $X2=0 $Y2=0
cc_145 N_A_81_23#_c_137_n N_C1_c_264_n 0.017623f $X=2.145 $Y=1.49 $X2=0 $Y2=0
cc_146 N_A_81_23#_c_142_n N_B1_M1010_g 0.0149464f $X=3.595 $Y=1.79 $X2=0 $Y2=0
cc_147 N_A_81_23#_c_144_n N_B1_M1025_g 0.0186522f $X=5.01 $Y=1.79 $X2=0 $Y2=0
cc_148 N_A_81_23#_c_142_n B1 0.0109013f $X=3.595 $Y=1.79 $X2=0 $Y2=0
cc_149 N_A_81_23#_c_146_n B1 0.0153391f $X=3.707 $Y=1.79 $X2=0 $Y2=0
cc_150 N_A_81_23#_c_144_n N_B1_c_310_n 0.00195096f $X=5.01 $Y=1.79 $X2=0 $Y2=0
cc_151 N_A_81_23#_c_146_n N_B1_c_310_n 0.00277011f $X=3.707 $Y=1.79 $X2=0 $Y2=0
cc_152 N_A_81_23#_c_144_n N_A3_M1004_g 0.0146156f $X=5.01 $Y=1.79 $X2=0 $Y2=0
cc_153 N_A_81_23#_c_145_n N_A3_c_352_n 0.00257648f $X=5.122 $Y=1.875 $X2=0 $Y2=0
cc_154 N_A_81_23#_c_144_n A3 0.0746894f $X=5.01 $Y=1.79 $X2=0 $Y2=0
cc_155 N_A_81_23#_c_145_n A3 0.0173628f $X=5.122 $Y=1.875 $X2=0 $Y2=0
cc_156 N_A_81_23#_c_136_n N_VPWR_M1024_d 0.00183167f $X=2.925 $Y=1.79 $X2=0
+ $Y2=0
cc_157 N_A_81_23#_c_142_n N_VPWR_M1027_d 0.00256188f $X=3.595 $Y=1.79 $X2=0
+ $Y2=0
cc_158 N_A_81_23#_c_144_n N_VPWR_M1025_s 0.00239457f $X=5.01 $Y=1.79 $X2=0 $Y2=0
cc_159 N_A_81_23#_M1003_g N_VPWR_c_494_n 0.0153838f $X=0.855 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_81_23#_M1014_g N_VPWR_c_494_n 7.27171e-19 $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_81_23#_M1003_g N_VPWR_c_495_n 7.24342e-19 $X=0.855 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_81_23#_M1014_g N_VPWR_c_495_n 0.0141881f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_81_23#_M1018_g N_VPWR_c_495_n 0.0141881f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_81_23#_M1024_g N_VPWR_c_495_n 7.24342e-19 $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_81_23#_M1018_g N_VPWR_c_496_n 7.41316e-19 $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_81_23#_M1024_g N_VPWR_c_496_n 0.0151578f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_81_23#_c_136_n N_VPWR_c_496_n 0.0187866f $X=2.925 $Y=1.79 $X2=0 $Y2=0
cc_168 N_A_81_23#_c_187_p N_VPWR_c_497_n 0.0138717f $X=2.79 $Y=1.98 $X2=0 $Y2=0
cc_169 N_A_81_23#_c_142_n N_VPWR_c_498_n 0.0196074f $X=3.595 $Y=1.79 $X2=0 $Y2=0
cc_170 N_A_81_23#_c_144_n N_VPWR_c_499_n 0.0220026f $X=5.01 $Y=1.79 $X2=0 $Y2=0
cc_171 N_A_81_23#_M1003_g N_VPWR_c_501_n 0.00486043f $X=0.855 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_81_23#_M1014_g N_VPWR_c_501_n 0.00486043f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_81_23#_M1018_g N_VPWR_c_503_n 0.00486043f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_174 N_A_81_23#_M1024_g N_VPWR_c_503_n 0.00486043f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A_81_23#_c_194_p N_VPWR_c_506_n 0.0136943f $X=3.725 $Y=1.98 $X2=0 $Y2=0
cc_176 N_A_81_23#_M1007_s N_VPWR_c_493_n 0.00397496f $X=2.65 $Y=1.835 $X2=0
+ $Y2=0
cc_177 N_A_81_23#_M1010_d N_VPWR_c_493_n 0.0041489f $X=3.585 $Y=1.835 $X2=0
+ $Y2=0
cc_178 N_A_81_23#_M1003_g N_VPWR_c_493_n 0.00824727f $X=0.855 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A_81_23#_M1014_g N_VPWR_c_493_n 0.00824727f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_81_23#_M1018_g N_VPWR_c_493_n 0.00824727f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_81_23#_M1024_g N_VPWR_c_493_n 0.00824727f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_81_23#_c_187_p N_VPWR_c_493_n 0.00886411f $X=2.79 $Y=1.98 $X2=0 $Y2=0
cc_183 N_A_81_23#_c_194_p N_VPWR_c_493_n 0.00866972f $X=3.725 $Y=1.98 $X2=0
+ $Y2=0
cc_184 N_A_81_23#_M1000_g N_X_c_602_n 0.0169287f $X=0.48 $Y=0.665 $X2=0 $Y2=0
cc_185 N_A_81_23#_c_204_p N_X_c_602_n 0.00491911f $X=2.195 $Y=1.495 $X2=0 $Y2=0
cc_186 N_A_81_23#_M1003_g N_X_c_607_n 0.0151995f $X=0.855 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A_81_23#_c_204_p N_X_c_607_n 0.0313614f $X=2.195 $Y=1.495 $X2=0 $Y2=0
cc_188 N_A_81_23#_c_137_n N_X_c_607_n 0.0108194f $X=2.145 $Y=1.49 $X2=0 $Y2=0
cc_189 N_A_81_23#_M1006_g N_X_c_603_n 0.0140083f $X=0.91 $Y=0.665 $X2=0 $Y2=0
cc_190 N_A_81_23#_M1008_g N_X_c_603_n 0.0137655f $X=1.34 $Y=0.665 $X2=0 $Y2=0
cc_191 N_A_81_23#_M1021_g N_X_c_603_n 0.00246848f $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_192 N_A_81_23#_c_204_p N_X_c_603_n 0.0655553f $X=2.195 $Y=1.495 $X2=0 $Y2=0
cc_193 N_A_81_23#_c_134_n N_X_c_603_n 0.0046745f $X=2.557 $Y=1.405 $X2=0 $Y2=0
cc_194 N_A_81_23#_c_137_n N_X_c_603_n 0.00550536f $X=2.145 $Y=1.49 $X2=0 $Y2=0
cc_195 N_A_81_23#_M1014_g N_X_c_609_n 0.0131755f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A_81_23#_M1018_g N_X_c_609_n 0.0130133f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A_81_23#_M1024_g N_X_c_609_n 6.54275e-19 $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A_81_23#_c_204_p N_X_c_609_n 0.0623153f $X=2.195 $Y=1.495 $X2=0 $Y2=0
cc_199 N_A_81_23#_c_136_n N_X_c_609_n 0.00877753f $X=2.925 $Y=1.79 $X2=0 $Y2=0
cc_200 N_A_81_23#_c_137_n N_X_c_609_n 0.00520544f $X=2.145 $Y=1.49 $X2=0 $Y2=0
cc_201 N_A_81_23#_c_204_p N_X_c_604_n 0.015388f $X=2.195 $Y=1.495 $X2=0 $Y2=0
cc_202 N_A_81_23#_c_137_n N_X_c_604_n 0.00256759f $X=2.145 $Y=1.49 $X2=0 $Y2=0
cc_203 N_A_81_23#_c_204_p N_X_c_610_n 0.0153881f $X=2.195 $Y=1.495 $X2=0 $Y2=0
cc_204 N_A_81_23#_c_137_n N_X_c_610_n 0.00277027f $X=2.145 $Y=1.49 $X2=0 $Y2=0
cc_205 N_A_81_23#_M1000_g X 0.0167765f $X=0.48 $Y=0.665 $X2=0 $Y2=0
cc_206 N_A_81_23#_M1003_g X 0.00275692f $X=0.855 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_81_23#_c_204_p X 0.0147324f $X=2.195 $Y=1.495 $X2=0 $Y2=0
cc_208 N_A_81_23#_c_144_n N_A_910_345#_M1004_d 0.00291209f $X=5.01 $Y=1.79
+ $X2=-0.19 $Y2=-0.245
cc_209 N_A_81_23#_c_144_n N_A_910_345#_c_658_n 0.0220026f $X=5.01 $Y=1.79 $X2=0
+ $Y2=0
cc_210 N_A_81_23#_M1004_s N_A_910_345#_c_659_n 0.00176461f $X=4.965 $Y=1.725
+ $X2=0 $Y2=0
cc_211 N_A_81_23#_c_230_p N_A_910_345#_c_659_n 0.0126348f $X=5.105 $Y=2.57 $X2=0
+ $Y2=0
cc_212 N_A_81_23#_c_145_n N_A_910_345#_c_661_n 0.00165793f $X=5.122 $Y=1.875
+ $X2=0 $Y2=0
cc_213 N_A_81_23#_M1000_g N_VGND_c_734_n 0.0116205f $X=0.48 $Y=0.665 $X2=0 $Y2=0
cc_214 N_A_81_23#_M1006_g N_VGND_c_734_n 6.10117e-19 $X=0.91 $Y=0.665 $X2=0
+ $Y2=0
cc_215 N_A_81_23#_M1000_g N_VGND_c_735_n 6.12946e-19 $X=0.48 $Y=0.665 $X2=0
+ $Y2=0
cc_216 N_A_81_23#_M1006_g N_VGND_c_735_n 0.0110192f $X=0.91 $Y=0.665 $X2=0 $Y2=0
cc_217 N_A_81_23#_M1008_g N_VGND_c_735_n 0.011105f $X=1.34 $Y=0.665 $X2=0 $Y2=0
cc_218 N_A_81_23#_M1021_g N_VGND_c_735_n 6.28047e-19 $X=1.77 $Y=0.665 $X2=0
+ $Y2=0
cc_219 N_A_81_23#_M1021_g N_VGND_c_736_n 0.00698774f $X=1.77 $Y=0.665 $X2=0
+ $Y2=0
cc_220 N_A_81_23#_c_204_p N_VGND_c_736_n 0.0153018f $X=2.195 $Y=1.495 $X2=0
+ $Y2=0
cc_221 N_A_81_23#_c_134_n N_VGND_c_736_n 0.00758963f $X=2.557 $Y=1.405 $X2=0
+ $Y2=0
cc_222 N_A_81_23#_c_135_n N_VGND_c_736_n 0.0219126f $X=2.795 $Y=0.89 $X2=0 $Y2=0
cc_223 N_A_81_23#_c_137_n N_VGND_c_736_n 0.00756387f $X=2.145 $Y=1.49 $X2=0
+ $Y2=0
cc_224 N_A_81_23#_M1008_g N_VGND_c_739_n 0.00477554f $X=1.34 $Y=0.665 $X2=0
+ $Y2=0
cc_225 N_A_81_23#_M1021_g N_VGND_c_739_n 0.00575161f $X=1.77 $Y=0.665 $X2=0
+ $Y2=0
cc_226 N_A_81_23#_M1000_g N_VGND_c_741_n 0.00477554f $X=0.48 $Y=0.665 $X2=0
+ $Y2=0
cc_227 N_A_81_23#_M1006_g N_VGND_c_741_n 0.00477554f $X=0.91 $Y=0.665 $X2=0
+ $Y2=0
cc_228 N_A_81_23#_M1012_d N_VGND_c_745_n 0.00225186f $X=2.795 $Y=0.235 $X2=0
+ $Y2=0
cc_229 N_A_81_23#_M1000_g N_VGND_c_745_n 0.00825815f $X=0.48 $Y=0.665 $X2=0
+ $Y2=0
cc_230 N_A_81_23#_M1006_g N_VGND_c_745_n 0.00825815f $X=0.91 $Y=0.665 $X2=0
+ $Y2=0
cc_231 N_A_81_23#_M1008_g N_VGND_c_745_n 0.00825815f $X=1.34 $Y=0.665 $X2=0
+ $Y2=0
cc_232 N_A_81_23#_M1021_g N_VGND_c_745_n 0.0118487f $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_233 N_A_81_23#_c_135_n N_VGND_c_745_n 0.00172834f $X=2.795 $Y=0.89 $X2=0
+ $Y2=0
cc_234 N_A_81_23#_c_134_n N_A_476_47#_M1012_s 2.77582e-19 $X=2.557 $Y=1.405
+ $X2=-0.19 $Y2=-0.245
cc_235 N_A_81_23#_c_135_n N_A_476_47#_M1012_s 0.00343667f $X=2.795 $Y=0.89
+ $X2=-0.19 $Y2=-0.245
cc_236 N_A_81_23#_M1012_d N_A_476_47#_c_845_n 0.00330375f $X=2.795 $Y=0.235
+ $X2=0 $Y2=0
cc_237 N_A_81_23#_c_135_n N_A_476_47#_c_845_n 0.0320809f $X=2.795 $Y=0.89 $X2=0
+ $Y2=0
cc_238 N_A_81_23#_c_155_p N_A_476_47#_c_845_n 0.0144025f $X=2.935 $Y=0.88 $X2=0
+ $Y2=0
cc_239 N_A_81_23#_c_146_n N_A_731_47#_c_884_n 0.00115675f $X=3.707 $Y=1.79 $X2=0
+ $Y2=0
cc_240 N_C1_c_262_n N_B1_c_306_n 0.015406f $X=3.15 $Y=1.185 $X2=0 $Y2=0
cc_241 C1 B1 0.0260314f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_242 N_C1_c_264_n B1 3.77007e-19 $X=3.06 $Y=1.36 $X2=0 $Y2=0
cc_243 N_C1_M1027_g N_B1_c_310_n 0.0202902f $X=3.005 $Y=2.465 $X2=0 $Y2=0
cc_244 C1 N_B1_c_310_n 0.00201123f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_245 N_C1_c_264_n N_B1_c_310_n 0.0217737f $X=3.06 $Y=1.36 $X2=0 $Y2=0
cc_246 N_C1_M1007_g N_VPWR_c_496_n 0.0152497f $X=2.575 $Y=2.465 $X2=0 $Y2=0
cc_247 N_C1_M1027_g N_VPWR_c_496_n 7.57541e-19 $X=3.005 $Y=2.465 $X2=0 $Y2=0
cc_248 N_C1_M1007_g N_VPWR_c_497_n 0.00486043f $X=2.575 $Y=2.465 $X2=0 $Y2=0
cc_249 N_C1_M1027_g N_VPWR_c_497_n 0.00585385f $X=3.005 $Y=2.465 $X2=0 $Y2=0
cc_250 N_C1_M1027_g N_VPWR_c_498_n 0.00194641f $X=3.005 $Y=2.465 $X2=0 $Y2=0
cc_251 N_C1_M1007_g N_VPWR_c_493_n 0.00824727f $X=2.575 $Y=2.465 $X2=0 $Y2=0
cc_252 N_C1_M1027_g N_VPWR_c_493_n 0.0107317f $X=3.005 $Y=2.465 $X2=0 $Y2=0
cc_253 N_C1_c_260_n N_VGND_c_736_n 0.0077455f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_254 N_C1_c_260_n N_VGND_c_745_n 0.00665089f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_255 N_C1_c_262_n N_VGND_c_745_n 0.00537654f $X=3.15 $Y=1.185 $X2=0 $Y2=0
cc_256 N_C1_c_260_n N_VGND_c_747_n 0.00357877f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_257 N_C1_c_262_n N_VGND_c_747_n 0.00357877f $X=3.15 $Y=1.185 $X2=0 $Y2=0
cc_258 N_C1_c_260_n N_A_476_47#_c_845_n 0.0121141f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_259 N_C1_c_262_n N_A_476_47#_c_845_n 0.0139071f $X=3.15 $Y=1.185 $X2=0 $Y2=0
cc_260 C1 N_A_476_47#_c_845_n 0.00398364f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_261 B1 A3 0.0242902f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_262 N_B1_c_310_n A3 0.0189192f $X=4.01 $Y=1.385 $X2=0 $Y2=0
cc_263 N_B1_M1010_g N_VPWR_c_498_n 0.0019647f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_264 N_B1_M1010_g N_VPWR_c_499_n 7.55536e-19 $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_265 N_B1_M1025_g N_VPWR_c_499_n 0.0166795f $X=3.94 $Y=2.465 $X2=0 $Y2=0
cc_266 N_B1_M1010_g N_VPWR_c_506_n 0.00585385f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_267 N_B1_M1025_g N_VPWR_c_506_n 0.00486043f $X=3.94 $Y=2.465 $X2=0 $Y2=0
cc_268 N_B1_M1010_g N_VPWR_c_493_n 0.010718f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_269 N_B1_M1025_g N_VPWR_c_493_n 0.00824727f $X=3.94 $Y=2.465 $X2=0 $Y2=0
cc_270 N_B1_M1025_g N_A_910_345#_c_658_n 0.00142977f $X=3.94 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_B1_c_306_n N_VGND_c_745_n 0.00537654f $X=3.58 $Y=1.195 $X2=0 $Y2=0
cc_272 N_B1_c_308_n N_VGND_c_745_n 0.0068216f $X=4.01 $Y=1.195 $X2=0 $Y2=0
cc_273 N_B1_c_306_n N_VGND_c_747_n 0.00357877f $X=3.58 $Y=1.195 $X2=0 $Y2=0
cc_274 N_B1_c_308_n N_VGND_c_747_n 0.00357877f $X=4.01 $Y=1.195 $X2=0 $Y2=0
cc_275 B1 N_A_476_47#_c_855_n 0.00141301f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_276 N_B1_c_306_n N_A_476_47#_c_856_n 0.0117305f $X=3.58 $Y=1.195 $X2=0 $Y2=0
cc_277 N_B1_c_308_n N_A_476_47#_c_856_n 0.0100985f $X=4.01 $Y=1.195 $X2=0 $Y2=0
cc_278 N_B1_c_308_n N_A_731_47#_c_876_n 0.0110228f $X=4.01 $Y=1.195 $X2=0 $Y2=0
cc_279 N_B1_c_308_n N_A_731_47#_c_877_n 0.00276351f $X=4.01 $Y=1.195 $X2=0 $Y2=0
cc_280 N_B1_c_306_n N_A_731_47#_c_884_n 0.00579274f $X=3.58 $Y=1.195 $X2=0 $Y2=0
cc_281 N_B1_c_308_n N_A_731_47#_c_884_n 0.00725026f $X=4.01 $Y=1.195 $X2=0 $Y2=0
cc_282 B1 N_A_731_47#_c_884_n 0.00982986f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_283 N_B1_c_310_n N_A_731_47#_c_884_n 0.00261823f $X=4.01 $Y=1.385 $X2=0 $Y2=0
cc_284 N_A3_c_351_n N_A2_M1002_g 0.01591f $X=5.89 $Y=1.185 $X2=0 $Y2=0
cc_285 A3 N_A2_M1002_g 6.73103e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_286 N_A3_M1019_g A2 0.00586916f $X=5.32 $Y=2.355 $X2=0 $Y2=0
cc_287 N_A3_c_353_n A2 0.00804767f $X=5.815 $Y=1.35 $X2=0 $Y2=0
cc_288 A3 A2 0.00744928f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_289 N_A3_c_353_n N_A2_c_402_n 0.01591f $X=5.815 $Y=1.35 $X2=0 $Y2=0
cc_290 N_A3_M1004_g N_VPWR_c_499_n 0.00255381f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_291 N_A3_M1004_g N_VPWR_c_507_n 0.00291444f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_292 N_A3_M1019_g N_VPWR_c_507_n 0.0029147f $X=5.32 $Y=2.355 $X2=0 $Y2=0
cc_293 N_A3_M1004_g N_VPWR_c_493_n 0.00428623f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_294 N_A3_M1019_g N_VPWR_c_493_n 0.00428625f $X=5.32 $Y=2.355 $X2=0 $Y2=0
cc_295 N_A3_M1004_g N_A_910_345#_c_658_n 0.0103497f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_296 N_A3_M1019_g N_A_910_345#_c_658_n 6.37286e-19 $X=5.32 $Y=2.355 $X2=0
+ $Y2=0
cc_297 N_A3_M1004_g N_A_910_345#_c_659_n 0.0101655f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_298 N_A3_M1019_g N_A_910_345#_c_659_n 0.0139445f $X=5.32 $Y=2.355 $X2=0 $Y2=0
cc_299 N_A3_M1004_g N_A_910_345#_c_660_n 0.00233316f $X=4.89 $Y=2.355 $X2=0
+ $Y2=0
cc_300 N_A3_M1019_g N_A_910_345#_c_661_n 0.00429211f $X=5.32 $Y=2.355 $X2=0
+ $Y2=0
cc_301 N_A3_c_353_n N_A_910_345#_c_661_n 0.00629614f $X=5.815 $Y=1.35 $X2=0
+ $Y2=0
cc_302 A3 N_A_910_345#_c_661_n 0.0210636f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_303 N_A3_c_351_n N_VGND_c_737_n 6.23782e-19 $X=5.89 $Y=1.185 $X2=0 $Y2=0
cc_304 N_A3_c_351_n N_VGND_c_742_n 0.00486043f $X=5.89 $Y=1.185 $X2=0 $Y2=0
cc_305 N_A3_c_349_n N_VGND_c_745_n 0.00949812f $X=4.96 $Y=1.185 $X2=0 $Y2=0
cc_306 N_A3_c_351_n N_VGND_c_745_n 0.00822376f $X=5.89 $Y=1.185 $X2=0 $Y2=0
cc_307 N_A3_c_349_n N_VGND_c_747_n 0.00486043f $X=4.96 $Y=1.185 $X2=0 $Y2=0
cc_308 N_A3_c_349_n N_VGND_c_748_n 0.015448f $X=4.96 $Y=1.185 $X2=0 $Y2=0
cc_309 N_A3_c_351_n N_VGND_c_748_n 0.0137202f $X=5.89 $Y=1.185 $X2=0 $Y2=0
cc_310 A3 N_A_731_47#_c_876_n 0.0456404f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_311 N_A3_c_349_n N_A_731_47#_c_892_n 0.0142704f $X=4.96 $Y=1.185 $X2=0 $Y2=0
cc_312 N_A3_c_351_n N_A_731_47#_c_892_n 0.0161285f $X=5.89 $Y=1.185 $X2=0 $Y2=0
cc_313 N_A3_c_352_n N_A_731_47#_c_892_n 0.0155017f $X=5.395 $Y=1.35 $X2=0 $Y2=0
cc_314 A3 N_A_731_47#_c_892_n 0.0575065f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_315 A3 N_A_731_47#_c_884_n 3.82325e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_316 N_A3_c_352_n N_A_731_47#_c_881_n 6.63067e-19 $X=5.395 $Y=1.35 $X2=0 $Y2=0
cc_317 A3 N_A_731_47#_c_881_n 0.0218414f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_318 N_A3_c_351_n N_A_731_47#_c_882_n 0.00396556f $X=5.89 $Y=1.185 $X2=0 $Y2=0
cc_319 A3 N_A_731_47#_c_882_n 0.00220918f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_320 N_A2_M1016_g N_A1_M1013_g 0.0192777f $X=6.75 $Y=0.655 $X2=0 $Y2=0
cc_321 N_A2_M1026_g N_A1_M1005_g 0.0192777f $X=6.75 $Y=2.465 $X2=0 $Y2=0
cc_322 A2 N_A1_M1005_g 0.00187199f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_323 A2 A1 0.0285236f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_324 A2 N_A1_c_458_n 0.00694149f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_325 N_A2_c_402_n N_A1_c_458_n 0.0192777f $X=6.75 $Y=1.51 $X2=0 $Y2=0
cc_326 N_A2_M1026_g N_VPWR_c_500_n 0.00131998f $X=6.75 $Y=2.465 $X2=0 $Y2=0
cc_327 N_A2_M1011_g N_VPWR_c_507_n 0.00357842f $X=6.32 $Y=2.465 $X2=0 $Y2=0
cc_328 N_A2_M1026_g N_VPWR_c_507_n 0.00547432f $X=6.75 $Y=2.465 $X2=0 $Y2=0
cc_329 N_A2_M1011_g N_VPWR_c_493_n 0.00675085f $X=6.32 $Y=2.465 $X2=0 $Y2=0
cc_330 N_A2_M1026_g N_VPWR_c_493_n 0.00990114f $X=6.75 $Y=2.465 $X2=0 $Y2=0
cc_331 N_A2_M1011_g N_A_910_345#_c_661_n 0.00808884f $X=6.32 $Y=2.465 $X2=0
+ $Y2=0
cc_332 A2 N_A_910_345#_c_661_n 0.00471539f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_333 N_A2_M1011_g N_A_910_345#_c_662_n 0.0131423f $X=6.32 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A2_M1026_g N_A_910_345#_c_662_n 0.00192258f $X=6.75 $Y=2.465 $X2=0
+ $Y2=0
cc_335 N_A2_M1011_g N_A_910_345#_c_682_n 0.0141764f $X=6.32 $Y=2.465 $X2=0 $Y2=0
cc_336 N_A2_M1026_g N_A_910_345#_c_682_n 0.00830481f $X=6.75 $Y=2.465 $X2=0
+ $Y2=0
cc_337 A2 N_A_1196_367#_c_701_n 0.0220966f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_338 N_A2_M1011_g N_A_1196_367#_c_706_n 0.0122595f $X=6.32 $Y=2.465 $X2=0
+ $Y2=0
cc_339 N_A2_M1026_g N_A_1196_367#_c_706_n 0.0122595f $X=6.75 $Y=2.465 $X2=0
+ $Y2=0
cc_340 A2 N_A_1196_367#_c_706_n 0.0428505f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_341 N_A2_c_402_n N_A_1196_367#_c_706_n 5.64665e-19 $X=6.75 $Y=1.51 $X2=0
+ $Y2=0
cc_342 A2 N_A_1196_367#_c_710_n 0.00255894f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_343 A2 N_A_1196_367#_c_711_n 0.0154122f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_344 N_A2_M1002_g N_VGND_c_737_n 0.0117053f $X=6.32 $Y=0.655 $X2=0 $Y2=0
cc_345 N_A2_M1016_g N_VGND_c_737_n 0.0117077f $X=6.75 $Y=0.655 $X2=0 $Y2=0
cc_346 N_A2_M1016_g N_VGND_c_738_n 6.36641e-19 $X=6.75 $Y=0.655 $X2=0 $Y2=0
cc_347 N_A2_M1002_g N_VGND_c_742_n 0.00486043f $X=6.32 $Y=0.655 $X2=0 $Y2=0
cc_348 N_A2_M1016_g N_VGND_c_743_n 0.00486043f $X=6.75 $Y=0.655 $X2=0 $Y2=0
cc_349 N_A2_M1002_g N_VGND_c_745_n 0.0082726f $X=6.32 $Y=0.655 $X2=0 $Y2=0
cc_350 N_A2_M1016_g N_VGND_c_745_n 0.0082726f $X=6.75 $Y=0.655 $X2=0 $Y2=0
cc_351 N_A2_M1002_g N_VGND_c_748_n 5.92296e-19 $X=6.32 $Y=0.655 $X2=0 $Y2=0
cc_352 A2 N_A_731_47#_c_892_n 0.00507253f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_353 N_A2_M1002_g N_A_731_47#_c_878_n 0.0130736f $X=6.32 $Y=0.655 $X2=0 $Y2=0
cc_354 N_A2_M1016_g N_A_731_47#_c_878_n 0.0142467f $X=6.75 $Y=0.655 $X2=0 $Y2=0
cc_355 A2 N_A_731_47#_c_878_n 0.0496265f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_356 N_A2_c_402_n N_A_731_47#_c_878_n 0.00246472f $X=6.75 $Y=1.51 $X2=0 $Y2=0
cc_357 N_A2_M1016_g N_A_731_47#_c_906_n 6.32385e-19 $X=6.75 $Y=0.655 $X2=0 $Y2=0
cc_358 A2 N_A_731_47#_c_879_n 0.00424945f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_359 N_A2_M1002_g N_A_731_47#_c_882_n 0.00103683f $X=6.32 $Y=0.655 $X2=0 $Y2=0
cc_360 A2 N_A_731_47#_c_882_n 0.0174998f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_361 A2 N_A_731_47#_c_883_n 0.0168258f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_362 N_A1_M1005_g N_VPWR_c_500_n 0.0156897f $X=7.18 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A1_M1020_g N_VPWR_c_500_n 0.0163814f $X=7.61 $Y=2.465 $X2=0 $Y2=0
cc_364 N_A1_M1005_g N_VPWR_c_507_n 0.00486043f $X=7.18 $Y=2.465 $X2=0 $Y2=0
cc_365 N_A1_M1020_g N_VPWR_c_508_n 0.00486043f $X=7.61 $Y=2.465 $X2=0 $Y2=0
cc_366 N_A1_M1005_g N_VPWR_c_493_n 0.0082726f $X=7.18 $Y=2.465 $X2=0 $Y2=0
cc_367 N_A1_M1020_g N_VPWR_c_493_n 0.00924348f $X=7.61 $Y=2.465 $X2=0 $Y2=0
cc_368 N_A1_M1005_g N_A_1196_367#_c_710_n 0.0144012f $X=7.18 $Y=2.465 $X2=0
+ $Y2=0
cc_369 N_A1_M1020_g N_A_1196_367#_c_710_n 0.0122595f $X=7.61 $Y=2.465 $X2=0
+ $Y2=0
cc_370 A1 N_A_1196_367#_c_710_n 0.0290298f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A1_c_458_n N_A_1196_367#_c_710_n 5.64665e-19 $X=7.61 $Y=1.51 $X2=0
+ $Y2=0
cc_372 A1 N_A_1196_367#_c_703_n 0.0220966f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_373 N_A1_M1013_g N_VGND_c_737_n 6.36641e-19 $X=7.18 $Y=0.655 $X2=0 $Y2=0
cc_374 N_A1_M1013_g N_VGND_c_738_n 0.0117077f $X=7.18 $Y=0.655 $X2=0 $Y2=0
cc_375 N_A1_M1023_g N_VGND_c_738_n 0.0135126f $X=7.61 $Y=0.655 $X2=0 $Y2=0
cc_376 N_A1_M1013_g N_VGND_c_743_n 0.00486043f $X=7.18 $Y=0.655 $X2=0 $Y2=0
cc_377 N_A1_M1023_g N_VGND_c_744_n 0.00486043f $X=7.61 $Y=0.655 $X2=0 $Y2=0
cc_378 N_A1_M1013_g N_VGND_c_745_n 0.0082726f $X=7.18 $Y=0.655 $X2=0 $Y2=0
cc_379 N_A1_M1023_g N_VGND_c_745_n 0.00924348f $X=7.61 $Y=0.655 $X2=0 $Y2=0
cc_380 N_A1_M1013_g N_A_731_47#_c_906_n 6.32385e-19 $X=7.18 $Y=0.655 $X2=0 $Y2=0
cc_381 N_A1_M1013_g N_A_731_47#_c_879_n 0.016435f $X=7.18 $Y=0.655 $X2=0 $Y2=0
cc_382 N_A1_M1023_g N_A_731_47#_c_879_n 0.0157274f $X=7.61 $Y=0.655 $X2=0 $Y2=0
cc_383 A1 N_A_731_47#_c_879_n 0.0560965f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_384 N_A1_c_458_n N_A_731_47#_c_879_n 0.00246472f $X=7.61 $Y=1.51 $X2=0 $Y2=0
cc_385 N_A1_M1023_g N_A_731_47#_c_880_n 0.00259704f $X=7.61 $Y=0.655 $X2=0 $Y2=0
cc_386 N_VPWR_c_493_n N_X_M1003_s 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_387 N_VPWR_c_493_n N_X_M1018_s 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_388 N_VPWR_M1003_d N_X_c_607_n 0.00262981f $X=0.515 $Y=1.835 $X2=0 $Y2=0
cc_389 N_VPWR_c_494_n N_X_c_607_n 0.0220025f $X=0.64 $Y=2.18 $X2=0 $Y2=0
cc_390 N_VPWR_c_501_n N_X_c_640_n 0.0124525f $X=1.335 $Y=3.33 $X2=0 $Y2=0
cc_391 N_VPWR_c_493_n N_X_c_640_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_392 N_VPWR_M1014_d N_X_c_609_n 0.00180746f $X=1.36 $Y=1.835 $X2=0 $Y2=0
cc_393 N_VPWR_c_495_n N_X_c_609_n 0.0163515f $X=1.5 $Y=2.19 $X2=0 $Y2=0
cc_394 N_VPWR_c_503_n N_X_c_644_n 0.0124525f $X=2.195 $Y=3.33 $X2=0 $Y2=0
cc_395 N_VPWR_c_493_n N_X_c_644_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_396 N_VPWR_c_493_n N_A_910_345#_M1011_d 0.00223559f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_499_n N_A_910_345#_c_658_n 0.0661835f $X=4.155 $Y=2.13 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_507_n N_A_910_345#_c_659_n 0.0355404f $X=7.23 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_493_n N_A_910_345#_c_659_n 0.0199839f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_499_n N_A_910_345#_c_660_n 0.0139f $X=4.155 $Y=2.13 $X2=0 $Y2=0
cc_401 N_VPWR_c_507_n N_A_910_345#_c_660_n 0.0235688f $X=7.23 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_493_n N_A_910_345#_c_660_n 0.0127152f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_507_n N_A_910_345#_c_662_n 0.0611478f $X=7.23 $Y=3.33 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_493_n N_A_910_345#_c_662_n 0.0378113f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_507_n N_A_910_345#_c_663_n 0.0197139f $X=7.23 $Y=3.33 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_493_n N_A_910_345#_c_663_n 0.0106914f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_493_n N_A_1196_367#_M1011_s 0.0021598f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_408 N_VPWR_c_493_n N_A_1196_367#_M1026_s 0.00536646f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_493_n N_A_1196_367#_M1020_d 0.00371702f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_507_n N_A_1196_367#_c_720_n 0.0124525f $X=7.23 $Y=3.33 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_493_n N_A_1196_367#_c_720_n 0.00730901f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_412 N_VPWR_M1005_s N_A_1196_367#_c_710_n 0.00333177f $X=7.255 $Y=1.835 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_500_n N_A_1196_367#_c_710_n 0.0170777f $X=7.395 $Y=2.39 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_508_n N_A_1196_367#_c_704_n 0.0178111f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_493_n N_A_1196_367#_c_704_n 0.0100304f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_416 N_X_c_605_n N_VGND_M1000_s 0.00244292f $X=0.222 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_417 N_X_c_603_n N_VGND_M1006_s 0.00176461f $X=1.46 $Y=1.15 $X2=0 $Y2=0
cc_418 N_X_c_602_n N_VGND_c_734_n 0.0017933f $X=0.6 $Y=1.145 $X2=0 $Y2=0
cc_419 N_X_c_605_n N_VGND_c_734_n 0.0224079f $X=0.222 $Y=1.235 $X2=0 $Y2=0
cc_420 N_X_c_603_n N_VGND_c_735_n 0.0170777f $X=1.46 $Y=1.15 $X2=0 $Y2=0
cc_421 N_X_c_603_n N_VGND_c_736_n 0.00166417f $X=1.46 $Y=1.15 $X2=0 $Y2=0
cc_422 N_X_c_652_p N_VGND_c_739_n 0.0138717f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_423 N_X_c_653_p N_VGND_c_741_n 0.0124525f $X=0.695 $Y=0.42 $X2=0 $Y2=0
cc_424 N_X_M1000_d N_VGND_c_745_n 0.00536646f $X=0.555 $Y=0.245 $X2=0 $Y2=0
cc_425 N_X_M1008_d N_VGND_c_745_n 0.00397496f $X=1.415 $Y=0.245 $X2=0 $Y2=0
cc_426 N_X_c_653_p N_VGND_c_745_n 0.00730901f $X=0.695 $Y=0.42 $X2=0 $Y2=0
cc_427 N_X_c_652_p N_VGND_c_745_n 0.00886411f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_428 N_A_910_345#_c_662_n N_A_1196_367#_M1011_s 0.00495471f $X=6.37 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_429 N_A_910_345#_c_661_n N_A_1196_367#_c_701_n 0.0110282f $X=5.535 $Y=1.87
+ $X2=0 $Y2=0
cc_430 N_A_910_345#_c_661_n N_A_1196_367#_c_702_n 0.0380785f $X=5.535 $Y=1.87
+ $X2=0 $Y2=0
cc_431 N_A_910_345#_c_662_n N_A_1196_367#_c_702_n 0.0189128f $X=6.37 $Y=2.99
+ $X2=0 $Y2=0
cc_432 N_A_910_345#_M1011_d N_A_1196_367#_c_706_n 0.00333177f $X=6.395 $Y=1.835
+ $X2=0 $Y2=0
cc_433 N_A_910_345#_c_682_n N_A_1196_367#_c_706_n 0.0170777f $X=6.535 $Y=2.39
+ $X2=0 $Y2=0
cc_434 N_A_1196_367#_c_710_n N_A_731_47#_c_879_n 0.00342491f $X=7.73 $Y=2.015
+ $X2=0 $Y2=0
cc_435 N_VGND_c_745_n N_A_476_47#_M1012_s 0.00215176f $X=7.92 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_436 N_VGND_c_745_n N_A_476_47#_M1022_s 0.00223565f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_745_n N_A_476_47#_M1009_s 0.00215161f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_438 N_VGND_c_736_n N_A_476_47#_c_845_n 0.0273835f $X=1.985 $Y=0.39 $X2=0
+ $Y2=0
cc_439 N_VGND_c_745_n N_A_476_47#_c_845_n 0.033994f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_747_n N_A_476_47#_c_845_n 0.0544569f $X=5.01 $Y=0.307 $X2=0
+ $Y2=0
cc_441 N_VGND_c_745_n N_A_476_47#_c_856_n 0.0237806f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_442 N_VGND_c_747_n N_A_476_47#_c_856_n 0.0362529f $X=5.01 $Y=0.307 $X2=0
+ $Y2=0
cc_443 N_VGND_c_745_n N_A_476_47#_c_866_n 0.00738676f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_444 N_VGND_c_747_n N_A_476_47#_c_866_n 0.0125234f $X=5.01 $Y=0.307 $X2=0
+ $Y2=0
cc_445 N_VGND_c_745_n N_A_476_47#_c_846_n 0.00991423f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_747_n N_A_476_47#_c_846_n 0.017241f $X=5.01 $Y=0.307 $X2=0 $Y2=0
cc_447 N_VGND_c_745_n N_A_731_47#_M1001_d 0.00225186f $X=7.92 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_448 N_VGND_c_745_n N_A_731_47#_M1015_s 0.00371702f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_449 N_VGND_c_745_n N_A_731_47#_M1017_s 0.00536646f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_450 N_VGND_c_745_n N_A_731_47#_M1016_s 0.00536646f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_745_n N_A_731_47#_M1023_d 0.00371702f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_745_n N_A_731_47#_c_876_n 0.00739898f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_453 N_VGND_c_745_n N_A_731_47#_c_877_n 0.0100304f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_454 N_VGND_c_747_n N_A_731_47#_c_877_n 0.0178111f $X=5.01 $Y=0.307 $X2=0
+ $Y2=0
cc_455 N_VGND_M1015_d N_A_731_47#_c_892_n 0.0175406f $X=5.035 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_VGND_c_748_n N_A_731_47#_c_892_n 0.0576541f $X=5.84 $Y=0.307 $X2=0
+ $Y2=0
cc_457 N_VGND_c_742_n N_A_731_47#_c_928_n 0.0124525f $X=6.37 $Y=0 $X2=0 $Y2=0
cc_458 N_VGND_c_745_n N_A_731_47#_c_928_n 0.00730901f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_459 N_VGND_c_737_n N_A_731_47#_c_878_n 0.0216087f $X=6.535 $Y=0.38 $X2=0
+ $Y2=0
cc_460 N_VGND_c_743_n N_A_731_47#_c_906_n 0.0124525f $X=7.23 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_745_n N_A_731_47#_c_906_n 0.00730901f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_462 N_VGND_c_738_n N_A_731_47#_c_879_n 0.0216087f $X=7.395 $Y=0.38 $X2=0
+ $Y2=0
cc_463 N_VGND_c_744_n N_A_731_47#_c_880_n 0.0178111f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_464 N_VGND_c_745_n N_A_731_47#_c_880_n 0.0100304f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_465 N_A_476_47#_c_856_n N_A_731_47#_M1001_d 0.00337224f $X=4.13 $Y=0.345
+ $X2=-0.19 $Y2=-0.245
cc_466 N_A_476_47#_M1009_s N_A_731_47#_c_876_n 0.00527241f $X=4.085 $Y=0.235
+ $X2=0 $Y2=0
cc_467 N_A_476_47#_c_856_n N_A_731_47#_c_876_n 0.00350393f $X=4.13 $Y=0.345
+ $X2=0 $Y2=0
cc_468 N_A_476_47#_c_846_n N_A_731_47#_c_876_n 0.0191744f $X=4.26 $Y=0.345 $X2=0
+ $Y2=0
cc_469 N_A_476_47#_c_846_n N_A_731_47#_c_877_n 0.0319372f $X=4.26 $Y=0.345 $X2=0
+ $Y2=0
cc_470 N_A_476_47#_c_856_n N_A_731_47#_c_884_n 0.0148612f $X=4.13 $Y=0.345 $X2=0
+ $Y2=0
