# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__and3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.470000 0.805000 2.120000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425000 1.345000 3.695000 1.750000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 1.345000 3.255000 1.750000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.075000 2.455000 1.245000 ;
        RECT 0.985000 1.245000 1.155000 1.815000 ;
        RECT 0.985000 1.815000 2.445000 2.145000 ;
        RECT 1.365000 0.255000 1.595000 1.075000 ;
        RECT 2.265000 0.255000 2.455000 1.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.205000  0.700000 0.455000 2.315000 ;
      RECT 0.205000  2.315000 2.455000 2.430000 ;
      RECT 0.205000  2.430000 4.035000 2.485000 ;
      RECT 0.905000  2.655000 1.235000 3.245000 ;
      RECT 0.975000  0.085000 1.195000 0.905000 ;
      RECT 1.335000  1.425000 2.795000 1.595000 ;
      RECT 1.765000  0.085000 2.095000 0.895000 ;
      RECT 1.765000  2.655000 2.095000 3.245000 ;
      RECT 2.265000  2.485000 4.035000 2.610000 ;
      RECT 2.625000  0.995000 4.690000 1.165000 ;
      RECT 2.625000  1.165000 2.795000 1.425000 ;
      RECT 2.625000  1.595000 2.795000 1.930000 ;
      RECT 2.625000  1.930000 3.400000 2.260000 ;
      RECT 2.625000  2.780000 2.955000 3.245000 ;
      RECT 2.695000  0.085000 3.025000 0.825000 ;
      RECT 3.330000  0.255000 4.690000 0.995000 ;
      RECT 3.560000  2.780000 3.890000 3.245000 ;
      RECT 3.865000  1.335000 4.340000 1.645000 ;
      RECT 3.865000  1.645000 4.035000 2.430000 ;
      RECT 4.205000  1.815000 4.690000 3.075000 ;
      RECT 4.520000  1.165000 4.690000 1.815000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__and3b_4
END LIBRARY
