* File: sky130_fd_sc_lp__decapkapwr_8.pex.spice
* Created: Wed Sep  2 09:42:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_8%VGND 1 12 15 17 18 22 26 30 31 41 42 45
+ 48
r31 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r32 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r33 42 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r34 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r35 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=0 $X2=3.095
+ $Y2=0
r36 39 41 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.26 $Y=0 $X2=3.6
+ $Y2=0
r37 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r38 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r40 34 37 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r41 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r43 32 34 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r44 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=0 $X2=3.095
+ $Y2=0
r45 31 37 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.93 $Y=0 $X2=2.64
+ $Y2=0
r46 26 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r47 26 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r48 22 24 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.095 $Y=0.36
+ $X2=3.095 $Y2=1.04
r49 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0
r50 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0.36
r51 18 30 22.4154 $w=1.774e-06 $l=1.03959e-06 $layer=POLY_cond $X=1.395 $Y=1.77
+ $X2=1.88 $Y2=2.595
r52 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.395
+ $Y=1.77 $X2=1.395 $Y2=1.77
r53 15 17 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.98 $Y=1.77
+ $X2=1.395 $Y2=1.77
r54 12 14 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.815 $Y=0.38
+ $X2=0.815 $Y2=1.06
r55 10 15 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=0.815 $Y=1.605
+ $X2=0.98 $Y2=1.77
r56 10 14 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.815 $Y=1.605
+ $X2=0.815 $Y2=1.06
r57 9 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r58 9 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.38
r59 1 24 121.333 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=3.095 $Y2=1.04
r60 1 22 121.333 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=3.095 $Y2=0.36
r61 1 14 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=0.815 $Y2=1.06
r62 1 12 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=0.815 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_8%KAPWR 1 7 9 11 13 16 22 24 25 28 36 41
r34 35 36 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.11 $Y=2.81
+ $X2=3.11 $Y2=2.81
r35 32 41 0.669526 $w=2.7e-07 $l=1.225e-06 $layer=MET1_cond $X=0.66 $Y=2.81
+ $X2=1.885 $Y2=2.81
r36 31 32 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.66 $Y=2.81
+ $X2=0.66 $Y2=2.81
r37 25 36 0.650397 $w=2.7e-07 $l=1.19e-06 $layer=MET1_cond $X=1.92 $Y=2.81
+ $X2=3.11 $Y2=2.81
r38 25 41 0.0191293 $w=2.7e-07 $l=3.5e-08 $layer=MET1_cond $X=1.92 $Y=2.81
+ $X2=1.885 $Y2=2.81
r39 22 35 3.05012 $w=4.2e-07 $l=2e-07 $layer=LI1_cond $X=3.075 $Y=2.675
+ $X2=3.075 $Y2=2.875
r40 22 24 10.5641 $w=4.18e-07 $l=3.85e-07 $layer=LI1_cond $X=3.075 $Y=2.675
+ $X2=3.075 $Y2=2.29
r41 21 24 16.8751 $w=4.18e-07 $l=6.15e-07 $layer=LI1_cond $X=3.075 $Y=1.675
+ $X2=3.075 $Y2=2.29
r42 16 28 20.7068 $w=1.804e-06 $l=7.75e-07 $layer=POLY_cond $X=1.96 $Y=1.51
+ $X2=1.96 $Y2=0.735
r43 16 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=1.51 $X2=2.8 $Y2=1.51
r44 15 19 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=2.12 $Y=1.507
+ $X2=2.8 $Y2=1.507
r45 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.12
+ $Y=1.51 $X2=2.12 $Y2=1.51
r46 13 21 6.92947 $w=3.35e-07 $l=2.81745e-07 $layer=LI1_cond $X=2.865 $Y=1.507
+ $X2=3.075 $Y2=1.675
r47 13 19 2.23608 $w=3.33e-07 $l=6.5e-08 $layer=LI1_cond $X=2.865 $Y=1.507
+ $X2=2.8 $Y2=1.507
r48 12 31 4.13568 $w=2.7e-07 $l=2.35266e-07 $layer=LI1_cond $X=0.905 $Y=2.81
+ $X2=0.7 $Y2=2.875
r49 11 35 4.19392 $w=2.7e-07 $l=2.40312e-07 $layer=LI1_cond $X=2.865 $Y=2.81
+ $X2=3.075 $Y2=2.875
r50 11 12 83.6588 $w=2.68e-07 $l=1.96e-06 $layer=LI1_cond $X=2.865 $Y=2.81
+ $X2=0.905 $Y2=2.81
r51 7 31 3.06347 $w=4.1e-07 $l=2e-07 $layer=LI1_cond $X=0.7 $Y=2.675 $X2=0.7
+ $Y2=2.875
r52 7 9 11.3839 $w=4.08e-07 $l=4.05e-07 $layer=LI1_cond $X=0.7 $Y=2.675 $X2=0.7
+ $Y2=2.27
r53 1 35 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=2.095 $X2=3.03 $Y2=2.97
r54 1 31 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=2.095 $X2=0.74 $Y2=2.95
r55 1 24 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=2.095 $X2=3.03 $Y2=2.29
r56 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=2.095 $X2=0.74 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_8%VPWR 1 8 14
r14 5 14 0.00397135 $w=3.84e-06 $l=1.22e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.92 $Y2=3.208
r15 5 8 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r16 4 8 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=3.6
+ $Y2=3.33
r17 4 5 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r18 1 14 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=3.207
+ $X2=1.92 $Y2=3.208
.ends

