* File: sky130_fd_sc_lp__or4bb_4.pex.spice
* Created: Wed Sep  2 10:33:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4BB_4%C_N 1 3 6 8 9 10 11
c28 1 0 3.72547e-20 $X=0.735 $Y=1.215
r29 10 11 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r30 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.38 $X2=0.27 $Y2=1.38
r31 8 15 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=0.66 $Y=1.38 $X2=0.27
+ $Y2=1.38
r32 8 9 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.66 $Y=1.38 $X2=0.735
+ $Y2=1.38
r33 4 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.735 $Y=1.545
+ $X2=0.735 $Y2=1.38
r34 4 6 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.735 $Y=1.545 $X2=0.735
+ $Y2=2.045
r35 1 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.735 $Y=1.215
+ $X2=0.735 $Y2=1.38
r36 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.735 $Y=1.215
+ $X2=0.735 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_4%A 3 6 8 9 13 15
c37 8 0 3.72547e-20 $X=1.2 $Y=1.295
r38 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.38
+ $X2=1.185 $Y2=1.545
r39 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.38
+ $X2=1.185 $Y2=1.215
r40 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.187 $Y=1.295
+ $X2=1.187 $Y2=1.665
r41 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.185
+ $Y=1.38 $X2=1.185 $Y2=1.38
r42 6 16 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=1.275 $Y=2.465
+ $X2=1.275 $Y2=1.545
r43 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.275 $Y=0.685
+ $X2=1.275 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_4%B 3 7 9 12 13
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.51
+ $X2=1.725 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.51 $X2=1.725 $Y2=1.51
r40 9 13 4.89394 $w=3.63e-07 $l=1.55e-07 $layer=LI1_cond $X=1.707 $Y=1.665
+ $X2=1.707 $Y2=1.51
r41 7 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.765 $Y=0.685
+ $X2=1.765 $Y2=1.345
r42 1 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.675
+ $X2=1.725 $Y2=1.51
r43 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.725 $Y=1.675
+ $X2=1.725 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_4%A_79_137# 1 2 9 13 16 17 18 21 22 27
r75 30 31 4.31095 $w=2.83e-07 $l=1e-07 $layer=LI1_cond $X=0.52 $Y=2.065 $X2=0.62
+ $Y2=2.065
r76 25 27 3.71756 $w=3.08e-07 $l=1e-07 $layer=LI1_cond $X=0.52 $Y=0.885 $X2=0.62
+ $Y2=0.885
r77 22 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.51
+ $X2=2.265 $Y2=1.675
r78 22 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.51
+ $X2=2.265 $Y2=1.345
r79 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.265
+ $Y=1.51 $X2=2.265 $Y2=1.51
r80 19 21 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=2.225 $Y=1.925
+ $X2=2.225 $Y2=1.51
r81 18 31 5.59441 $w=2.83e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.705 $Y=2.01
+ $X2=0.62 $Y2=2.065
r82 17 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.1 $Y=2.01
+ $X2=2.225 $Y2=1.925
r83 17 18 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.1 $Y=2.01
+ $X2=0.705 $Y2=2.01
r84 16 31 3.71884 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.62 $Y=1.92
+ $X2=0.62 $Y2=2.065
r85 15 27 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.62 $Y=1.04
+ $X2=0.62 $Y2=0.885
r86 15 16 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.62 $Y=1.04
+ $X2=0.62 $Y2=1.92
r87 13 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.285 $Y=0.685
+ $X2=2.285 $Y2=1.345
r88 9 34 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.175 $Y=2.465
+ $X2=2.175 $Y2=1.675
r89 2 30 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=1.835 $X2=0.52 $Y2=2.045
r90 1 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.395
+ $Y=0.685 $X2=0.52 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_4%A_528_27# 1 2 7 9 12 16 17 19 20 21 22 29
c89 22 0 1.68898e-19 $X=5.607 $Y=1.92
r90 26 29 3.69577 $w=2.88e-07 $l=9.3e-08 $layer=LI1_cond $X=5.607 $Y=2.065
+ $X2=5.7 $Y2=2.065
r91 24 25 5.99107 $w=3.36e-07 $l=1.65e-07 $layer=LI1_cond $X=5.687 $Y=0.475
+ $X2=5.687 $Y2=0.64
r92 22 26 3.08157 $w=1.95e-07 $l=1.45e-07 $layer=LI1_cond $X=5.607 $Y=1.92
+ $X2=5.607 $Y2=2.065
r93 21 25 5.2167 $w=3.36e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.607 $Y=0.725
+ $X2=5.687 $Y2=0.64
r94 21 22 67.9674 $w=1.93e-07 $l=1.195e-06 $layer=LI1_cond $X=5.607 $Y=0.725
+ $X2=5.607 $Y2=1.92
r95 19 25 4.73076 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=5.51 $Y=0.64
+ $X2=5.687 $Y2=0.64
r96 19 20 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=5.51 $Y=0.64
+ $X2=3.13 $Y2=0.64
r97 17 31 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.965 $Y=1.38
+ $X2=2.715 $Y2=1.38
r98 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.38 $X2=2.965 $Y2=1.38
r99 14 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3 $Y=0.725
+ $X2=3.13 $Y2=0.64
r100 14 16 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=3 $Y=0.725 $X2=3
+ $Y2=1.38
r101 10 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.545
+ $X2=2.715 $Y2=1.38
r102 10 12 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=2.715 $Y=1.545
+ $X2=2.715 $Y2=2.465
r103 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.215
+ $X2=2.715 $Y2=1.38
r104 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.715 $Y=1.215
+ $X2=2.715 $Y2=0.685
r105 2 29 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.56
+ $Y=1.835 $X2=5.7 $Y2=2.045
r106 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.265 $X2=5.7 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_4%A_270_53# 1 2 3 12 16 20 24 28 32 36 40 44
+ 46 47 50 53 56 60 61 62 63 66 69 84
c152 40 0 1.68898e-19 $X=4.96 $Y=2.465
r153 81 82 20.8558 $w=3.12e-07 $l=1.35e-07 $layer=POLY_cond $X=4.395 $Y=1.49
+ $X2=4.53 $Y2=1.49
r154 80 81 45.5737 $w=3.12e-07 $l=2.95e-07 $layer=POLY_cond $X=4.1 $Y=1.49
+ $X2=4.395 $Y2=1.49
r155 79 80 39.3942 $w=3.12e-07 $l=2.55e-07 $layer=POLY_cond $X=3.845 $Y=1.49
+ $X2=4.1 $Y2=1.49
r156 78 79 27.0353 $w=3.12e-07 $l=1.75e-07 $layer=POLY_cond $X=3.67 $Y=1.49
+ $X2=3.845 $Y2=1.49
r157 75 78 20.8558 $w=3.12e-07 $l=1.35e-07 $layer=POLY_cond $X=3.535 $Y=1.49
+ $X2=3.67 $Y2=1.49
r158 75 76 18.5385 $w=3.12e-07 $l=1.2e-07 $layer=POLY_cond $X=3.535 $Y=1.49
+ $X2=3.415 $Y2=1.49
r159 74 75 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.535
+ $Y=1.49 $X2=3.535 $Y2=1.49
r160 67 84 41.7115 $w=3.12e-07 $l=2.7e-07 $layer=POLY_cond $X=4.555 $Y=1.49
+ $X2=4.825 $Y2=1.49
r161 67 82 3.86218 $w=3.12e-07 $l=2.5e-08 $layer=POLY_cond $X=4.555 $Y=1.49
+ $X2=4.53 $Y2=1.49
r162 66 67 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.555
+ $Y=1.49 $X2=4.555 $Y2=1.49
r163 64 74 3.3405 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=3.54 $Y=1.45 $X2=3.42
+ $Y2=1.45
r164 64 66 46.7892 $w=2.48e-07 $l=1.015e-06 $layer=LI1_cond $X=3.54 $Y=1.45
+ $X2=4.555 $Y2=1.45
r165 62 74 3.47969 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=3.42 $Y=1.575
+ $X2=3.42 $Y2=1.45
r166 62 63 8.64332 $w=2.38e-07 $l=1.8e-07 $layer=LI1_cond $X=3.42 $Y=1.575
+ $X2=3.42 $Y2=1.755
r167 60 63 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.3 $Y=1.84
+ $X2=3.42 $Y2=1.755
r168 60 61 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.3 $Y=1.84
+ $X2=3.095 $Y2=1.84
r169 56 58 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=2.93 $Y=1.98
+ $X2=2.93 $Y2=2.91
r170 54 61 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=1.84
+ $X2=3.095 $Y2=1.84
r171 54 70 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.93 $Y=1.84
+ $X2=2.615 $Y2=1.84
r172 54 56 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=2.93 $Y=1.925
+ $X2=2.93 $Y2=1.98
r173 53 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=1.755
+ $X2=2.615 $Y2=1.84
r174 52 69 3.67481 $w=2.52e-07 $l=1.19499e-07 $layer=LI1_cond $X=2.615 $Y=1.165
+ $X2=2.532 $Y2=1.08
r175 52 53 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.615 $Y=1.165
+ $X2=2.615 $Y2=1.755
r176 48 69 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=2.532 $Y=0.995
+ $X2=2.532 $Y2=1.08
r177 48 50 19.7807 $w=3.33e-07 $l=5.75e-07 $layer=LI1_cond $X=2.532 $Y=0.995
+ $X2=2.532 $Y2=0.42
r178 46 69 2.79892 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.365 $Y=1.08
+ $X2=2.532 $Y2=1.08
r179 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.365 $Y=1.08
+ $X2=1.695 $Y2=1.08
r180 42 47 23.4276 $w=8.2e-08 $l=2.03101e-07 $layer=LI1_cond $X=1.53 $Y=0.995
+ $X2=1.695 $Y2=1.08
r181 42 44 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=0.42
r182 38 84 20.8558 $w=3.12e-07 $l=2.22486e-07 $layer=POLY_cond $X=4.96 $Y=1.655
+ $X2=4.825 $Y2=1.49
r183 38 40 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.96 $Y=1.655
+ $X2=4.96 $Y2=2.465
r184 34 84 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.825 $Y=1.325
+ $X2=4.825 $Y2=1.49
r185 34 36 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.825 $Y=1.325
+ $X2=4.825 $Y2=0.685
r186 30 82 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.53 $Y=1.655
+ $X2=4.53 $Y2=1.49
r187 30 32 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.53 $Y=1.655
+ $X2=4.53 $Y2=2.465
r188 26 81 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.325
+ $X2=4.395 $Y2=1.49
r189 26 28 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.395 $Y=1.325
+ $X2=4.395 $Y2=0.685
r190 22 80 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.1 $Y=1.655
+ $X2=4.1 $Y2=1.49
r191 22 24 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.1 $Y=1.655 $X2=4.1
+ $Y2=2.465
r192 18 79 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.325
+ $X2=3.845 $Y2=1.49
r193 18 20 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.845 $Y=1.325
+ $X2=3.845 $Y2=0.685
r194 14 78 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.655
+ $X2=3.67 $Y2=1.49
r195 14 16 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.67 $Y=1.655
+ $X2=3.67 $Y2=2.465
r196 10 76 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=1.325
+ $X2=3.415 $Y2=1.49
r197 10 12 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.415 $Y=1.325
+ $X2=3.415 $Y2=0.685
r198 3 58 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.835 $X2=2.93 $Y2=2.91
r199 3 56 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.835 $X2=2.93 $Y2=1.98
r200 2 50 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.265 $X2=2.5 $Y2=0.42
r201 1 44 91 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_NDIFF $count=2 $X=1.35
+ $Y=0.265 $X2=1.525 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_4%D_N 3 7 9 10 14 15
r25 14 17 75.2115 $w=7.25e-07 $l=5.05e-07 $layer=POLY_cond $X=5.772 $Y=1.12
+ $X2=5.772 $Y2=1.625
r26 14 16 51.0986 $w=7.25e-07 $l=1.65e-07 $layer=POLY_cond $X=5.772 $Y=1.12
+ $X2=5.772 $Y2=0.955
r27 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.97
+ $Y=1.12 $X2=5.97 $Y2=1.12
r28 9 10 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=6.015 $Y=1.295
+ $X2=6.015 $Y2=1.665
r29 9 15 7.20277 $w=2.78e-07 $l=1.75e-07 $layer=LI1_cond $X=6.015 $Y=1.295
+ $X2=6.015 $Y2=1.12
r30 7 17 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=5.485 $Y=2.045
+ $X2=5.485 $Y2=1.625
r31 3 16 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.485 $Y=0.475
+ $X2=5.485 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_4%VPWR 1 2 3 4 15 19 25 29 33 38 39 40 41 42
+ 44 58 59 62 65
r68 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r69 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 59 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r71 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r72 56 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.34 $Y=3.33
+ $X2=5.175 $Y2=3.33
r73 56 58 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.34 $Y=3.33 $X2=6
+ $Y2=3.33
r74 55 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r75 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 49 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.06 $Y2=3.33
r77 49 51 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=3.12 $Y2=3.33
r78 47 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r79 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 44 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.06 $Y2=3.33
r81 44 46 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.72 $Y2=3.33
r82 42 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r83 42 63 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=1.2 $Y2=3.33
r84 42 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 40 54 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.15 $Y=3.33 $X2=4.08
+ $Y2=3.33
r86 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=4.315 $Y2=3.33
r87 38 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.29 $Y=3.33
+ $X2=3.12 $Y2=3.33
r88 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=3.33
+ $X2=3.455 $Y2=3.33
r89 37 54 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.62 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=3.33
+ $X2=3.455 $Y2=3.33
r91 33 36 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.175 $Y=2.17
+ $X2=5.175 $Y2=2.555
r92 31 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.175 $Y=3.245
+ $X2=5.175 $Y2=3.33
r93 31 36 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.175 $Y=3.245
+ $X2=5.175 $Y2=2.555
r94 30 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.48 $Y=3.33
+ $X2=4.315 $Y2=3.33
r95 29 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=5.175 $Y2=3.33
r96 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=4.48 $Y2=3.33
r97 25 28 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=4.315 $Y=2.17
+ $X2=4.315 $Y2=2.95
r98 23 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=3.245
+ $X2=4.315 $Y2=3.33
r99 23 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.315 $Y=3.245
+ $X2=4.315 $Y2=2.95
r100 19 22 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.455 $Y=2.18
+ $X2=3.455 $Y2=2.95
r101 17 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=3.245
+ $X2=3.455 $Y2=3.33
r102 17 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.455 $Y=3.245
+ $X2=3.455 $Y2=2.95
r103 13 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=3.245
+ $X2=1.06 $Y2=3.33
r104 13 15 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=1.06 $Y=3.245
+ $X2=1.06 $Y2=2.395
r105 4 36 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=5.035
+ $Y=1.835 $X2=5.175 $Y2=2.555
r106 4 33 600 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=5.035
+ $Y=1.835 $X2=5.175 $Y2=2.17
r107 3 28 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=1.835 $X2=4.315 $Y2=2.95
r108 3 25 400 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=1.835 $X2=4.315 $Y2=2.17
r109 2 22 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=1.835 $X2=3.455 $Y2=2.95
r110 2 19 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=1.835 $X2=3.455 $Y2=2.18
r111 1 15 300 $w=1.7e-07 $l=6.73498e-07 $layer=licon1_PDIFF $count=2 $X=0.81
+ $Y=1.835 $X2=1.06 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_4%X 1 2 3 4 13 21 25 26 29 34 35 39 44
r52 39 44 2.7521 $w=3.33e-07 $l=8e-08 $layer=LI1_cond $X=5.057 $Y=1.745
+ $X2=5.057 $Y2=1.665
r53 35 39 1.10909 $w=1.68e-07 $l=1.7e-08 $layer=LI1_cond $X=5.04 $Y=1.83
+ $X2=5.057 $Y2=1.83
r54 35 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.04 $Y=1.83
+ $X2=4.745 $Y2=1.83
r55 35 44 0.103204 $w=3.33e-07 $l=3e-09 $layer=LI1_cond $X=5.057 $Y=1.662
+ $X2=5.057 $Y2=1.665
r56 34 35 12.6253 $w=3.33e-07 $l=3.67e-07 $layer=LI1_cond $X=5.057 $Y=1.295
+ $X2=5.057 $Y2=1.662
r57 33 34 5.16019 $w=3.33e-07 $l=1.5e-07 $layer=LI1_cond $X=5.057 $Y=1.145
+ $X2=5.057 $Y2=1.295
r58 29 31 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=4.745 $Y=1.98
+ $X2=4.745 $Y2=2.91
r59 27 45 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.745 $Y=1.915
+ $X2=4.745 $Y2=1.83
r60 27 29 3.79426 $w=1.88e-07 $l=6.5e-08 $layer=LI1_cond $X=4.745 $Y=1.915
+ $X2=4.745 $Y2=1.98
r61 25 45 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.65 $Y=1.83
+ $X2=4.745 $Y2=1.83
r62 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.65 $Y=1.83
+ $X2=3.98 $Y2=1.83
r63 21 23 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.885 $Y=1.98
+ $X2=3.885 $Y2=2.91
r64 19 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.885 $Y=1.915
+ $X2=3.98 $Y2=1.83
r65 19 21 3.79426 $w=1.88e-07 $l=6.5e-08 $layer=LI1_cond $X=3.885 $Y=1.915
+ $X2=3.885 $Y2=1.98
r66 15 18 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=3.63 $Y=1.02
+ $X2=4.61 $Y2=1.02
r67 13 33 7.00535 $w=2.5e-07 $l=2.20826e-07 $layer=LI1_cond $X=4.89 $Y=1.02
+ $X2=5.057 $Y2=1.145
r68 13 18 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=4.89 $Y=1.02
+ $X2=4.61 $Y2=1.02
r69 4 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.605
+ $Y=1.835 $X2=4.745 $Y2=2.91
r70 4 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.605
+ $Y=1.835 $X2=4.745 $Y2=1.98
r71 3 23 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.835 $X2=3.885 $Y2=2.91
r72 3 21 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.835 $X2=3.885 $Y2=1.98
r73 2 18 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=4.47
+ $Y=0.265 $X2=4.61 $Y2=0.98
r74 1 15 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=3.49
+ $Y=0.265 $X2=3.63 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_4%VGND 1 2 3 4 5 18 24 26 29 30 32 33 34 43 47
+ 54 55 59 66 73
r79 73 76 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=5.155
+ $Y2=0.28
r80 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r81 67 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r82 66 69 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.12 $Y=0 $X2=4.12
+ $Y2=0.28
r83 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r84 59 62 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.045
+ $Y2=0.28
r85 55 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r86 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r87 52 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.155
+ $Y2=0
r88 52 54 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.32 $Y=0 $X2=6
+ $Y2=0
r89 51 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r90 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r91 48 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.21 $Y=0 $X2=3.045
+ $Y2=0
r92 48 50 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.21 $Y=0 $X2=3.6
+ $Y2=0
r93 47 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=0 $X2=4.12
+ $Y2=0
r94 47 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=0 $X2=3.6
+ $Y2=0
r95 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r96 43 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=3.045
+ $Y2=0
r97 43 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r98 42 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r99 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r100 38 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r101 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r102 34 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r103 34 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r104 34 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r105 32 41 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=1.68 $Y2=0
r106 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.03
+ $Y2=0
r107 31 45 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.195 $Y=0
+ $X2=2.64 $Y2=0
r108 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.03
+ $Y2=0
r109 29 37 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.72 $Y2=0
r110 29 30 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.035
+ $Y2=0
r111 28 41 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.195 $Y=0
+ $X2=1.68 $Y2=0
r112 28 30 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.035
+ $Y2=0
r113 27 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.12
+ $Y2=0
r114 26 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.99 $Y=0 $X2=5.155
+ $Y2=0
r115 26 27 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.99 $Y=0
+ $X2=4.285 $Y2=0
r116 22 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0
r117 22 24 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0.39
r118 18 20 16.7464 $w=3.18e-07 $l=4.65e-07 $layer=LI1_cond $X=1.035 $Y=0.41
+ $X2=1.035 $Y2=0.875
r119 16 30 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.085
+ $X2=1.035 $Y2=0
r120 16 18 11.7045 $w=3.18e-07 $l=3.25e-07 $layer=LI1_cond $X=1.035 $Y=0.085
+ $X2=1.035 $Y2=0.41
r121 5 76 182 $w=1.7e-07 $l=2.62393e-07 $layer=licon1_NDIFF $count=1 $X=4.9
+ $Y=0.265 $X2=5.155 $Y2=0.28
r122 4 69 182 $w=1.7e-07 $l=2.07364e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.265 $X2=4.12 $Y2=0.28
r123 3 62 182 $w=1.7e-07 $l=2.62393e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.265 $X2=3.045 $Y2=0.28
r124 2 24 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.265 $X2=2.03 $Y2=0.39
r125 1 20 182 $w=1.7e-07 $l=2.54165e-07 $layer=licon1_NDIFF $count=1 $X=0.81
+ $Y=0.685 $X2=0.96 $Y2=0.875
r126 1 18 182 $w=1.7e-07 $l=3.79967e-07 $layer=licon1_NDIFF $count=1 $X=0.81
+ $Y=0.685 $X2=1.06 $Y2=0.41
.ends

