* File: sky130_fd_sc_lp__einvp_0.spice
* Created: Wed Sep  2 09:52:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvp_0.pex.spice"
.subckt sky130_fd_sc_lp__einvp_0  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_TE_M1003_g N_A_32_70#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1004 A_201_70# N_TE_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_Z_M1005_d N_A_M1005_g A_201_70# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_TE_M1000_g N_A_32_70#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0855057 AS=0.1113 PD=0.80434 PS=1.37 NRD=39.8531 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 A_220_484# N_A_32_70#_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.130294 PD=0.88 PS=1.22566 NRD=19.9955 NRS=3.8415 M=1 R=4.26667
+ SA=75000.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g A_220_484# VPB PHIGHVT L=0.15 W=0.64 AD=0.1824
+ AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75000.9
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.2895 P=8.33
*
.include "sky130_fd_sc_lp__einvp_0.pxi.spice"
*
.ends
*
*
