* File: sky130_fd_sc_lp__clkinv_8.pex.spice
* Created: Fri Aug 28 10:18:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKINV_8%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55
+ 59 63 67 71 75 79 81 82 83 84 85 86 87 88 89 90 119
r167 117 119 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.1 $Y=1.375
+ $X2=5.275 $Y2=1.375
r168 115 117 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=4.845 $Y=1.375
+ $X2=5.1 $Y2=1.375
r169 114 115 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.415 $Y=1.375
+ $X2=4.845 $Y2=1.375
r170 113 114 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.985 $Y=1.375
+ $X2=4.415 $Y2=1.375
r171 112 113 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.555 $Y=1.375
+ $X2=3.985 $Y2=1.375
r172 111 112 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.125 $Y=1.375
+ $X2=3.555 $Y2=1.375
r173 110 111 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.695 $Y=1.375
+ $X2=3.125 $Y2=1.375
r174 109 110 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.265 $Y=1.375
+ $X2=2.695 $Y2=1.375
r175 108 109 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.835 $Y=1.375
+ $X2=2.265 $Y2=1.375
r176 107 108 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.405 $Y=1.375
+ $X2=1.835 $Y2=1.375
r177 106 107 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.975 $Y=1.375
+ $X2=1.405 $Y2=1.375
r178 104 106 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=0.68 $Y=1.375
+ $X2=0.975 $Y2=1.375
r179 101 104 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.545 $Y=1.375
+ $X2=0.68 $Y2=1.375
r180 90 117 20.7543 $w=1.7e-07 $l=1.19e-06 $layer=licon1_POLY $count=7 $X=5.1
+ $Y=1.375 $X2=5.1 $Y2=1.375
r181 89 90 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.375
+ $X2=5.04 $Y2=1.375
r182 88 89 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.375
+ $X2=4.56 $Y2=1.375
r183 87 88 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.375
+ $X2=4.08 $Y2=1.375
r184 86 87 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.375
+ $X2=3.6 $Y2=1.375
r185 85 86 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.375
+ $X2=3.12 $Y2=1.375
r186 84 85 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.375
+ $X2=2.64 $Y2=1.375
r187 83 84 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.375
+ $X2=2.16 $Y2=1.375
r188 82 83 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.375
+ $X2=1.68 $Y2=1.375
r189 81 82 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=0.68 $Y=1.375
+ $X2=1.2 $Y2=1.375
r190 81 104 20.7543 $w=1.7e-07 $l=1.19e-06 $layer=licon1_POLY $count=7 $X=0.68
+ $Y=1.375 $X2=0.68 $Y2=1.375
r191 77 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.275 $Y=1.54
+ $X2=5.275 $Y2=1.375
r192 77 79 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=5.275 $Y=1.54
+ $X2=5.275 $Y2=2.465
r193 73 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.845 $Y=1.54
+ $X2=4.845 $Y2=1.375
r194 73 75 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=4.845 $Y=1.54
+ $X2=4.845 $Y2=2.465
r195 69 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.54
+ $X2=4.415 $Y2=1.375
r196 69 71 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=4.415 $Y=1.54
+ $X2=4.415 $Y2=2.465
r197 65 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.21
+ $X2=4.415 $Y2=1.375
r198 65 67 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=4.415 $Y=1.21
+ $X2=4.415 $Y2=0.56
r199 61 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.54
+ $X2=3.985 $Y2=1.375
r200 61 63 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.985 $Y=1.54
+ $X2=3.985 $Y2=2.465
r201 57 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.21
+ $X2=3.985 $Y2=1.375
r202 57 59 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.985 $Y=1.21
+ $X2=3.985 $Y2=0.56
r203 53 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.555 $Y=1.54
+ $X2=3.555 $Y2=1.375
r204 53 55 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.555 $Y=1.54
+ $X2=3.555 $Y2=2.465
r205 49 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.555 $Y=1.21
+ $X2=3.555 $Y2=1.375
r206 49 51 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.555 $Y=1.21
+ $X2=3.555 $Y2=0.56
r207 45 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.54
+ $X2=3.125 $Y2=1.375
r208 45 47 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.125 $Y=1.54
+ $X2=3.125 $Y2=2.465
r209 41 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.21
+ $X2=3.125 $Y2=1.375
r210 41 43 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.125 $Y=1.21
+ $X2=3.125 $Y2=0.56
r211 37 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.54
+ $X2=2.695 $Y2=1.375
r212 37 39 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.695 $Y=1.54
+ $X2=2.695 $Y2=2.465
r213 33 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.21
+ $X2=2.695 $Y2=1.375
r214 33 35 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.695 $Y=1.21
+ $X2=2.695 $Y2=0.56
r215 29 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.54
+ $X2=2.265 $Y2=1.375
r216 29 31 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.265 $Y=1.54
+ $X2=2.265 $Y2=2.465
r217 25 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.21
+ $X2=2.265 $Y2=1.375
r218 25 27 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.265 $Y=1.21
+ $X2=2.265 $Y2=0.56
r219 21 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.54
+ $X2=1.835 $Y2=1.375
r220 21 23 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.835 $Y=1.54
+ $X2=1.835 $Y2=2.465
r221 17 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.21
+ $X2=1.835 $Y2=1.375
r222 17 19 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.835 $Y=1.21
+ $X2=1.835 $Y2=0.56
r223 13 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.54
+ $X2=1.405 $Y2=1.375
r224 13 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.405 $Y=1.54
+ $X2=1.405 $Y2=2.465
r225 9 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.21
+ $X2=1.405 $Y2=1.375
r226 9 11 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.405 $Y=1.21
+ $X2=1.405 $Y2=0.56
r227 5 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.54
+ $X2=0.975 $Y2=1.375
r228 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.975 $Y=1.54
+ $X2=0.975 $Y2=2.465
r229 1 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.54
+ $X2=0.545 $Y2=1.375
r230 1 3 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.545 $Y=1.54
+ $X2=0.545 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_8%VPWR 1 2 3 4 5 6 7 22 24 30 36 42 48 52 56
+ 60 62 67 68 70 71 72 73 74 76 91 100 103 107
r92 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r95 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r96 95 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 95 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r98 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r99 92 103 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=4.63 $Y2=3.33
r100 92 94 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=5.04 $Y2=3.33
r101 91 106 4.00962 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=5.36 $Y=3.33 $X2=5.56
+ $Y2=3.33
r102 91 94 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.36 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 90 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r104 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 84 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r108 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 81 100 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.19 $Y2=3.33
r110 81 83 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.68 $Y2=3.33
r111 80 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 80 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r114 77 97 3.99713 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.23 $Y2=3.33
r115 77 79 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 76 100 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=1.19 $Y2=3.33
r117 76 79 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 74 90 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r119 74 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 72 89 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r121 72 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.64 $Y=3.33
+ $X2=3.77 $Y2=3.33
r122 70 86 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.78 $Y=3.33
+ $X2=2.64 $Y2=3.33
r123 70 71 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.78 $Y=3.33
+ $X2=2.91 $Y2=3.33
r124 69 89 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r125 69 71 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.04 $Y=3.33
+ $X2=2.91 $Y2=3.33
r126 67 83 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 67 68 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=2.05 $Y2=3.33
r128 66 86 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.18 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 66 68 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.18 $Y=3.33
+ $X2=2.05 $Y2=3.33
r130 62 65 31.4097 $w=2.53e-07 $l=6.95e-07 $layer=LI1_cond $X=5.487 $Y=2.22
+ $X2=5.487 $Y2=2.915
r131 60 106 3.1676 $w=2.55e-07 $l=1.15888e-07 $layer=LI1_cond $X=5.487 $Y=3.245
+ $X2=5.56 $Y2=3.33
r132 60 65 14.914 $w=2.53e-07 $l=3.3e-07 $layer=LI1_cond $X=5.487 $Y=3.245
+ $X2=5.487 $Y2=2.915
r133 56 59 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=4.63 $Y=2.22
+ $X2=4.63 $Y2=2.915
r134 54 103 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=3.245
+ $X2=4.63 $Y2=3.33
r135 54 59 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=4.63 $Y=3.245
+ $X2=4.63 $Y2=2.915
r136 53 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.9 $Y=3.33 $X2=3.77
+ $Y2=3.33
r137 52 103 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.5 $Y=3.33
+ $X2=4.63 $Y2=3.33
r138 52 53 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.5 $Y=3.33 $X2=3.9
+ $Y2=3.33
r139 48 51 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=3.77 $Y=2.22
+ $X2=3.77 $Y2=2.915
r140 46 73 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=3.245
+ $X2=3.77 $Y2=3.33
r141 46 51 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=3.77 $Y=3.245
+ $X2=3.77 $Y2=2.915
r142 42 45 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=2.91 $Y=2.22
+ $X2=2.91 $Y2=2.915
r143 40 71 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=3.245
+ $X2=2.91 $Y2=3.33
r144 40 45 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=2.91 $Y=3.245
+ $X2=2.91 $Y2=2.915
r145 36 39 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=2.05 $Y=2.22
+ $X2=2.05 $Y2=2.915
r146 34 68 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=3.245
+ $X2=2.05 $Y2=3.33
r147 34 39 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=2.05 $Y=3.245
+ $X2=2.05 $Y2=2.915
r148 30 33 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=1.19 $Y=2.22
+ $X2=1.19 $Y2=2.915
r149 28 100 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=3.33
r150 28 33 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=2.915
r151 24 27 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=0.33 $Y=2.22
+ $X2=0.33 $Y2=2.915
r152 22 97 3.21509 $w=2.6e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.23 $Y2=3.33
r153 22 27 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.33 $Y2=2.915
r154 7 65 400 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.835 $X2=5.49 $Y2=2.915
r155 7 62 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.835 $X2=5.49 $Y2=2.22
r156 6 59 400 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=4.49
+ $Y=1.835 $X2=4.63 $Y2=2.915
r157 6 56 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=4.49
+ $Y=1.835 $X2=4.63 $Y2=2.22
r158 5 51 400 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=3.63
+ $Y=1.835 $X2=3.77 $Y2=2.915
r159 5 48 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=3.63
+ $Y=1.835 $X2=3.77 $Y2=2.22
r160 4 45 400 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.835 $X2=2.91 $Y2=2.915
r161 4 42 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.835 $X2=2.91 $Y2=2.22
r162 3 39 400 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=2.915
r163 3 36 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=2.22
r164 2 33 400 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.915
r165 2 30 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.22
r166 1 27 400 $w=1.7e-07 $l=1.14079e-06 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.915
r167 1 24 400 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_8%Y 1 2 3 4 5 6 7 8 9 10 32 33 34 35 36 39 43
+ 47 51 55 57 61 65 69 71 75 79 83 85 89 93 97 101 105 107 108 109 110 111 112
+ 113 115 116 117 119 120 124
r161 120 124 15.2875 $w=1.83e-07 $l=2.55e-07 $layer=LI1_cond $X=5.527 $Y=1.295
+ $X2=5.527 $Y2=1.04
r162 119 124 3.55727 $w=1.85e-07 $l=1e-07 $layer=LI1_cond $X=5.527 $Y=0.94
+ $X2=5.527 $Y2=1.04
r163 118 120 24.8796 $w=1.83e-07 $l=4.15e-07 $layer=LI1_cond $X=5.527 $Y=1.71
+ $X2=5.527 $Y2=1.295
r164 114 119 35.7429 $w=3.68e-07 $l=1.105e-06 $layer=LI1_cond $X=4.33 $Y=0.94
+ $X2=5.435 $Y2=0.94
r165 114 115 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=4.33 $Y=0.94 $X2=4.2
+ $Y2=0.94
r166 106 117 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=5.19 $Y=1.797
+ $X2=5.06 $Y2=1.797
r167 105 118 6.82334 $w=1.75e-07 $l=1.28328e-07 $layer=LI1_cond $X=5.435
+ $Y=1.797 $X2=5.527 $Y2=1.71
r168 105 106 15.5273 $w=1.73e-07 $l=2.45e-07 $layer=LI1_cond $X=5.435 $Y=1.797
+ $X2=5.19 $Y2=1.797
r169 101 103 39.0058 $w=2.58e-07 $l=8.8e-07 $layer=LI1_cond $X=5.06 $Y=2
+ $X2=5.06 $Y2=2.88
r170 99 117 0.0359085 $w=2.6e-07 $l=8.8e-08 $layer=LI1_cond $X=5.06 $Y=1.885
+ $X2=5.06 $Y2=1.797
r171 99 101 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=5.06 $Y=1.885
+ $X2=5.06 $Y2=2
r172 98 116 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=4.33 $Y=1.797
+ $X2=4.202 $Y2=1.797
r173 97 117 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=4.93 $Y=1.797
+ $X2=5.06 $Y2=1.797
r174 97 98 38.026 $w=1.73e-07 $l=6e-07 $layer=LI1_cond $X=4.93 $Y=1.797 $X2=4.33
+ $Y2=1.797
r175 93 95 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=4.202 $Y=2
+ $X2=4.202 $Y2=2.88
r176 91 116 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=4.202 $Y=1.885
+ $X2=4.202 $Y2=1.797
r177 91 93 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=4.202 $Y=1.885
+ $X2=4.202 $Y2=2
r178 87 115 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=4.2 $Y=0.84 $X2=4.2
+ $Y2=0.94
r179 87 89 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=4.2 $Y=0.84 $X2=4.2
+ $Y2=0.56
r180 86 113 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=3.47 $Y=1.797
+ $X2=3.342 $Y2=1.797
r181 85 116 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=4.075 $Y=1.797
+ $X2=4.202 $Y2=1.797
r182 85 86 38.3429 $w=1.73e-07 $l=6.05e-07 $layer=LI1_cond $X=4.075 $Y=1.797
+ $X2=3.47 $Y2=1.797
r183 84 112 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=3.47 $Y=0.94 $X2=3.34
+ $Y2=0.94
r184 83 115 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=4.07 $Y=0.94 $X2=4.2
+ $Y2=0.94
r185 83 84 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=4.07 $Y=0.94 $X2=3.47
+ $Y2=0.94
r186 79 81 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=3.342 $Y=2
+ $X2=3.342 $Y2=2.88
r187 77 113 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=3.342 $Y=1.885
+ $X2=3.342 $Y2=1.797
r188 77 79 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=3.342 $Y=1.885
+ $X2=3.342 $Y2=2
r189 73 112 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=3.34 $Y=0.84
+ $X2=3.34 $Y2=0.94
r190 73 75 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=3.34 $Y=0.84
+ $X2=3.34 $Y2=0.56
r191 72 111 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=2.61 $Y=1.797
+ $X2=2.482 $Y2=1.797
r192 71 113 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=3.215 $Y=1.797
+ $X2=3.342 $Y2=1.797
r193 71 72 38.3429 $w=1.73e-07 $l=6.05e-07 $layer=LI1_cond $X=3.215 $Y=1.797
+ $X2=2.61 $Y2=1.797
r194 70 110 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=2.61 $Y=0.94 $X2=2.48
+ $Y2=0.94
r195 69 112 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=3.21 $Y=0.94 $X2=3.34
+ $Y2=0.94
r196 69 70 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=3.21 $Y=0.94 $X2=2.61
+ $Y2=0.94
r197 65 67 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=2.482 $Y=2
+ $X2=2.482 $Y2=2.88
r198 63 111 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=2.482 $Y=1.885
+ $X2=2.482 $Y2=1.797
r199 63 65 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=2.482 $Y=1.885
+ $X2=2.482 $Y2=2
r200 59 110 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=2.48 $Y=0.84
+ $X2=2.48 $Y2=0.94
r201 59 61 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=2.48 $Y=0.84
+ $X2=2.48 $Y2=0.56
r202 58 109 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=1.75 $Y=1.797
+ $X2=1.622 $Y2=1.797
r203 57 111 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=2.355 $Y=1.797
+ $X2=2.482 $Y2=1.797
r204 57 58 38.3429 $w=1.73e-07 $l=6.05e-07 $layer=LI1_cond $X=2.355 $Y=1.797
+ $X2=1.75 $Y2=1.797
r205 56 108 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.75 $Y=0.94 $X2=1.62
+ $Y2=0.94
r206 55 110 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=2.35 $Y=0.94 $X2=2.48
+ $Y2=0.94
r207 55 56 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=2.35 $Y=0.94 $X2=1.75
+ $Y2=0.94
r208 51 53 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=1.622 $Y=2
+ $X2=1.622 $Y2=2.88
r209 49 109 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=1.622 $Y=1.885
+ $X2=1.622 $Y2=1.797
r210 49 51 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=1.622 $Y=1.885
+ $X2=1.622 $Y2=2
r211 45 108 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=1.62 $Y=0.84
+ $X2=1.62 $Y2=0.94
r212 45 47 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=1.62 $Y=0.84
+ $X2=1.62 $Y2=0.56
r213 44 107 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=0.89 $Y=1.797
+ $X2=0.762 $Y2=1.797
r214 43 109 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=1.495 $Y=1.797
+ $X2=1.622 $Y2=1.797
r215 43 44 38.3429 $w=1.73e-07 $l=6.05e-07 $layer=LI1_cond $X=1.495 $Y=1.797
+ $X2=0.89 $Y2=1.797
r216 39 41 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=0.762 $Y=2
+ $X2=0.762 $Y2=2.88
r217 37 107 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=0.762 $Y=1.885
+ $X2=0.762 $Y2=1.797
r218 37 39 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=0.762 $Y=1.885
+ $X2=0.762 $Y2=2
r219 35 107 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=0.635 $Y=1.797
+ $X2=0.762 $Y2=1.797
r220 35 36 18.3792 $w=1.73e-07 $l=2.9e-07 $layer=LI1_cond $X=0.635 $Y=1.797
+ $X2=0.345 $Y2=1.797
r221 33 108 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.49 $Y=0.94 $X2=1.62
+ $Y2=0.94
r222 33 34 63.4955 $w=1.98e-07 $l=1.145e-06 $layer=LI1_cond $X=1.49 $Y=0.94
+ $X2=0.345 $Y2=0.94
r223 32 36 6.81835 $w=1.75e-07 $l=1.22327e-07 $layer=LI1_cond $X=0.26 $Y=1.71
+ $X2=0.345 $Y2=1.797
r224 31 34 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.26 $Y=1.04
+ $X2=0.345 $Y2=0.94
r225 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.26 $Y=1.04
+ $X2=0.26 $Y2=1.71
r226 10 103 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.835 $X2=5.06 $Y2=2.88
r227 10 101 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.835 $X2=5.06 $Y2=2
r228 9 95 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=4.06
+ $Y=1.835 $X2=4.2 $Y2=2.88
r229 9 93 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=4.06
+ $Y=1.835 $X2=4.2 $Y2=2
r230 8 81 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.835 $X2=3.34 $Y2=2.88
r231 8 79 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.835 $X2=3.34 $Y2=2
r232 7 67 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=1.835 $X2=2.48 $Y2=2.88
r233 7 65 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=1.835 $X2=2.48 $Y2=2
r234 6 53 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=2.88
r235 6 51 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=2
r236 5 41 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2.88
r237 5 39 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2
r238 4 89 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.35 $X2=4.2 $Y2=0.56
r239 3 75 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.35 $X2=3.34 $Y2=0.56
r240 2 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.34
+ $Y=0.35 $X2=2.48 $Y2=0.56
r241 1 47 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.35 $X2=1.62 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_8%VGND 1 2 3 4 5 18 22 26 30 32 36 39 40 42
+ 43 44 45 46 48 65 66 69 72
r61 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r62 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r63 66 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r64 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r65 63 72 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.647
+ $Y2=0
r66 63 65 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=5.52
+ $Y2=0
r67 62 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r68 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r69 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r70 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r71 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r72 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r73 53 69 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.172
+ $Y2=0
r74 53 55 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.68
+ $Y2=0
r75 51 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r76 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r77 48 69 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.172
+ $Y2=0
r78 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=0.72
+ $Y2=0
r79 46 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r80 46 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r81 44 61 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.6
+ $Y2=0
r82 44 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.77
+ $Y2=0
r83 42 58 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.64
+ $Y2=0
r84 42 43 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.91
+ $Y2=0
r85 41 61 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.6
+ $Y2=0
r86 41 43 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.91
+ $Y2=0
r87 39 55 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r88 39 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=2.05
+ $Y2=0
r89 38 58 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.64
+ $Y2=0
r90 38 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.05
+ $Y2=0
r91 34 72 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.647 $Y=0.085
+ $X2=4.647 $Y2=0
r92 34 36 16.4077 $w=2.93e-07 $l=4.2e-07 $layer=LI1_cond $X=4.647 $Y=0.085
+ $X2=4.647 $Y2=0.505
r93 33 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.9 $Y=0 $X2=3.77
+ $Y2=0
r94 32 72 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=4.647
+ $Y2=0
r95 32 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=3.9 $Y2=0
r96 28 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=0.085
+ $X2=3.77 $Y2=0
r97 28 30 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=3.77 $Y=0.085
+ $X2=3.77 $Y2=0.505
r98 24 43 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.91 $Y2=0
r99 24 26 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.91 $Y2=0.505
r100 20 40 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=0.085
+ $X2=2.05 $Y2=0
r101 20 22 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=2.05 $Y=0.085
+ $X2=2.05 $Y2=0.505
r102 16 69 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.172 $Y=0.085
+ $X2=1.172 $Y2=0
r103 16 18 16.4077 $w=2.93e-07 $l=4.2e-07 $layer=LI1_cond $X=1.172 $Y=0.085
+ $X2=1.172 $Y2=0.505
r104 5 36 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.49
+ $Y=0.35 $X2=4.63 $Y2=0.505
r105 4 30 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.35 $X2=3.77 $Y2=0.505
r106 3 26 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.77
+ $Y=0.35 $X2=2.91 $Y2=0.505
r107 2 22 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.35 $X2=2.05 $Y2=0.505
r108 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.35 $X2=1.19 $Y2=0.505
.ends

