# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 1.550000 2.735000 1.760000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.115000 0.255000 13.375000 1.065000 ;
        RECT 13.115000 1.755000 13.375000 3.075000 ;
        RECT 13.200000 1.065000 13.375000 1.755000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.795000 1.950000 6.125000 2.305000 ;
        RECT 5.795000 2.305000 6.925000 2.475000 ;
        RECT 6.755000 2.475000 6.925000 2.525000 ;
        RECT 6.755000 2.525000 9.405000 2.695000 ;
        RECT 9.075000 2.250000 9.405000 2.525000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.210000 3.285000 2.130000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 1.200000 2.735000 1.380000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 11.630000 1.415000 12.005000 2.490000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.920000 0.085000 ;
        RECT  0.565000  0.085000  0.895000 0.690000 ;
        RECT  3.405000  0.085000  3.735000 0.665000 ;
        RECT  6.145000  0.085000  6.475000 0.615000 ;
        RECT  8.470000  0.085000  8.800000 0.955000 ;
        RECT 10.880000  0.085000 11.210000 0.475000 ;
        RECT 12.615000  0.085000 12.945000 0.475000 ;
        RECT 13.545000  0.085000 13.815000 1.095000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.920000 3.415000 ;
        RECT  1.205000 2.320000  1.475000 3.245000 ;
        RECT  2.970000 2.640000  3.300000 3.245000 ;
        RECT  4.855000 2.515000  5.185000 3.245000 ;
        RECT  6.245000 2.645000  6.575000 3.245000 ;
        RECT  8.410000 2.865000  9.140000 3.245000 ;
        RECT  9.925000 2.705000 10.175000 3.245000 ;
        RECT 10.805000 2.665000 11.120000 3.245000 ;
        RECT 12.545000 2.015000 12.945000 3.245000 ;
        RECT 13.545000 1.815000 13.815000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.135000 0.415000  0.395000 0.860000 ;
      RECT  0.135000 0.860000  1.510000 1.030000 ;
      RECT  0.135000 1.030000  0.405000 1.930000 ;
      RECT  0.135000 1.930000  2.560000 2.130000 ;
      RECT  0.135000 2.130000  1.035000 3.000000 ;
      RECT  1.085000 0.265000  3.225000 0.435000 ;
      RECT  1.085000 0.435000  1.415000 0.625000 ;
      RECT  1.990000 0.605000  2.320000 0.835000 ;
      RECT  1.990000 0.835000  4.215000 1.005000 ;
      RECT  1.995000 2.300000  3.885000 2.470000 ;
      RECT  1.995000 2.470000  2.325000 3.000000 ;
      RECT  2.895000 0.435000  3.225000 0.665000 ;
      RECT  3.455000 1.005000  3.680000 2.300000 ;
      RECT  3.510000 2.470000  3.885000 2.970000 ;
      RECT  3.850000 1.175000  4.215000 1.995000 ;
      RECT  3.955000 0.640000  4.215000 0.835000 ;
      RECT  4.055000 2.175000  5.625000 2.345000 ;
      RECT  4.055000 2.345000  4.385000 2.695000 ;
      RECT  4.385000 0.640000  4.800000 0.785000 ;
      RECT  4.385000 0.785000  6.475000 0.995000 ;
      RECT  4.385000 0.995000  4.555000 2.175000 ;
      RECT  4.725000 1.600000  6.835000 1.770000 ;
      RECT  4.725000 1.770000  5.010000 1.995000 ;
      RECT  4.735000 1.165000  5.200000 1.430000 ;
      RECT  5.355000 2.345000  5.625000 2.695000 ;
      RECT  6.145000 0.995000  6.475000 1.430000 ;
      RECT  6.645000 0.325000  6.835000 1.600000 ;
      RECT  6.655000 1.770000  6.835000 1.945000 ;
      RECT  6.655000 1.945000  7.100000 2.135000 ;
      RECT  7.005000 0.325000  8.235000 0.925000 ;
      RECT  7.005000 0.925000  7.175000 1.605000 ;
      RECT  7.005000 1.605000  7.555000 1.775000 ;
      RECT  7.270000 1.775000  7.555000 2.355000 ;
      RECT  7.345000 1.095000  7.895000 1.425000 ;
      RECT  7.725000 1.425000  7.895000 2.095000 ;
      RECT  7.725000 2.095000  8.075000 2.355000 ;
      RECT  8.065000 0.925000  8.235000 1.205000 ;
      RECT  8.065000 1.205000 10.000000 1.375000 ;
      RECT  8.065000 1.555000  8.245000 1.560000 ;
      RECT  8.065000 1.560000 10.105000 1.730000 ;
      RECT  8.065000 1.730000  8.325000 1.885000 ;
      RECT  8.535000 1.910000  9.755000 2.080000 ;
      RECT  8.535000 2.080000  8.865000 2.275000 ;
      RECT  9.310000 2.865000  9.755000 3.075000 ;
      RECT  9.380000 0.255000 10.110000 0.475000 ;
      RECT  9.380000 0.475000  9.660000 0.970000 ;
      RECT  9.585000 2.080000  9.755000 2.865000 ;
      RECT  9.830000 0.645000 12.070000 0.815000 ;
      RECT  9.830000 0.815000 10.000000 1.205000 ;
      RECT  9.935000 1.730000 10.105000 2.325000 ;
      RECT  9.935000 2.325000 11.460000 2.495000 ;
      RECT 10.210000 0.985000 10.700000 1.165000 ;
      RECT 10.210000 1.165000 10.635000 1.425000 ;
      RECT 10.375000 1.425000 10.635000 2.155000 ;
      RECT 10.805000 1.345000 11.460000 2.325000 ;
      RECT 11.290000 0.985000 11.720000 1.245000 ;
      RECT 11.290000 1.245000 11.460000 1.345000 ;
      RECT 11.290000 2.495000 11.460000 2.660000 ;
      RECT 11.290000 2.660000 11.720000 2.940000 ;
      RECT 11.900000 0.815000 12.070000 0.995000 ;
      RECT 11.900000 0.995000 12.540000 1.245000 ;
      RECT 12.115000 0.275000 12.445000 0.465000 ;
      RECT 12.175000 1.675000 12.890000 1.845000 ;
      RECT 12.175000 1.845000 12.375000 2.495000 ;
      RECT 12.210000 1.245000 12.540000 1.505000 ;
      RECT 12.275000 0.465000 12.445000 0.645000 ;
      RECT 12.275000 0.645000 12.945000 0.815000 ;
      RECT 12.720000 0.815000 12.945000 1.245000 ;
      RECT 12.720000 1.245000 13.030000 1.575000 ;
      RECT 12.720000 1.575000 12.890000 1.675000 ;
    LAYER mcon ;
      RECT  3.995000 1.210000  4.165000 1.380000 ;
      RECT  4.955000 1.210000  5.125000 1.380000 ;
      RECT  7.355000 1.210000  7.525000 1.380000 ;
      RECT 10.235000 1.210000 10.405000 1.380000 ;
    LAYER met1 ;
      RECT  3.935000 1.180000  4.225000 1.225000 ;
      RECT  3.935000 1.225000 10.465000 1.365000 ;
      RECT  3.935000 1.365000  4.225000 1.410000 ;
      RECT  4.895000 1.180000  5.185000 1.225000 ;
      RECT  4.895000 1.365000  5.185000 1.410000 ;
      RECT  7.295000 1.180000  7.585000 1.225000 ;
      RECT  7.295000 1.365000  7.585000 1.410000 ;
      RECT 10.175000 1.180000 10.465000 1.225000 ;
      RECT 10.175000 1.365000 10.465000 1.410000 ;
  END
END sky130_fd_sc_lp__sdfrtp_2
