* File: sky130_fd_sc_lp__clkinv_1.spice
* Created: Wed Sep  2 09:40:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkinv_1.pex.spice"
.subckt sky130_fd_sc_lp__clkinv_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX3_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__clkinv_1.pxi.spice"
*
.ends
*
*
