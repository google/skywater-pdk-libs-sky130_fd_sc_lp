* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o22a_m A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 VPWR a_88_187# X VPB phighvt w=420000u l=150000u
+  ad=5.124e+11p pd=4.12e+06u as=1.197e+11p ps=1.41e+06u
M1001 a_88_187# B2 a_339_535# VPB phighvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=8.82e+10p ps=1.26e+06u
M1002 VGND a_88_187# X VNB nshort w=420000u l=150000u
+  ad=3.213e+11p pd=3.21e+06u as=1.197e+11p ps=1.41e+06u
M1003 VGND A2 a_237_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.024e+11p ps=3.12e+06u
M1004 a_339_535# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A1 a_519_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_519_535# A2 a_88_187# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_237_81# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_88_187# B1 a_237_81# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1009 a_237_81# B2 a_88_187# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
