* File: sky130_fd_sc_lp__and3_0.spice
* Created: Fri Aug 28 10:05:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and3_0.pex.spice"
.subckt sky130_fd_sc_lp__and3_0  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 A_157_65# N_A_M1005_g N_A_68_65#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1239 PD=0.63 PS=1.43 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1003 A_229_65# N_B_M1003_g A_157_65# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_C_M1001_g A_229_65# VNB NSHORT L=0.15 W=0.42 AD=0.17325
+ AS=0.0441 PD=1.245 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.9 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_68_65#_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.17325 PD=1.37 PS=1.245 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_68_65#_M1007_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_68_65#_M1002_d N_B_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_A_68_65#_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.14066 AS=0.0588 PD=0.998491 PS=0.7 NRD=53.9386 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_68_65#_M1004_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.176 AS=0.21434 PD=1.83 PS=1.52151 NRD=0 NRS=17.6906 M=1 R=4.26667
+ SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__and3_0.pxi.spice"
*
.ends
*
*
