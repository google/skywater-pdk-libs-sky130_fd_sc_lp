# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__buf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.890000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.365000 1.385000 2.735000 1.585000 ;
        RECT 1.905000 1.205000 2.255000 1.385000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  4.704000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.225000 1.920000 9.535000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.195000  0.085000  0.490000 1.075000 ;
      RECT 0.195000  1.815000  0.490000 3.245000 ;
      RECT 0.660000  0.425000  0.920000 1.045000 ;
      RECT 0.660000  1.045000  1.735000 1.215000 ;
      RECT 0.660000  1.755000  3.095000 1.925000 ;
      RECT 0.660000  1.925000  0.920000 3.075000 ;
      RECT 1.090000  0.085000  1.360000 0.875000 ;
      RECT 1.090000  2.095000  1.350000 3.245000 ;
      RECT 1.520000  1.925000  1.780000 3.075000 ;
      RECT 1.530000  0.425000  1.745000 0.865000 ;
      RECT 1.530000  0.865000  2.640000 1.035000 ;
      RECT 1.530000  1.035000  1.735000 1.045000 ;
      RECT 1.915000  0.085000  2.245000 0.695000 ;
      RECT 1.950000  2.095000  2.210000 3.245000 ;
      RECT 2.380000  1.925000  2.640000 3.075000 ;
      RECT 2.415000  0.425000  2.640000 0.865000 ;
      RECT 2.425000  1.035000  2.640000 1.045000 ;
      RECT 2.425000  1.045000  3.095000 1.215000 ;
      RECT 2.810000  0.085000  3.095000 0.875000 ;
      RECT 2.810000  2.095000  3.095000 3.245000 ;
      RECT 2.905000  1.215000  3.095000 1.755000 ;
      RECT 3.265000  0.255000  3.500000 3.075000 ;
      RECT 3.670000  0.085000  3.930000 1.075000 ;
      RECT 3.670000  1.325000  3.930000 1.750000 ;
      RECT 3.670000  1.920000  3.930000 3.245000 ;
      RECT 4.100000  0.255000  4.360000 3.075000 ;
      RECT 4.530000  0.085000  4.790000 1.075000 ;
      RECT 4.530000  1.325000  4.790000 1.750000 ;
      RECT 4.530000  1.920000  4.790000 3.245000 ;
      RECT 4.960000  0.255000  5.220000 3.075000 ;
      RECT 5.390000  0.085000  5.650000 1.075000 ;
      RECT 5.390000  1.325000  5.650000 1.750000 ;
      RECT 5.390000  1.920000  5.650000 3.245000 ;
      RECT 5.820000  0.255000  6.080000 3.075000 ;
      RECT 6.250000  0.085000  6.510000 1.075000 ;
      RECT 6.250000  1.325000  6.510000 1.750000 ;
      RECT 6.250000  1.920000  6.510000 3.245000 ;
      RECT 6.680000  0.255000  6.940000 3.075000 ;
      RECT 7.110000  0.085000  7.370000 1.075000 ;
      RECT 7.110000  1.325000  7.370000 1.750000 ;
      RECT 7.110000  1.920000  7.370000 3.245000 ;
      RECT 7.540000  0.255000  7.800000 3.075000 ;
      RECT 7.970000  0.085000  8.230000 1.075000 ;
      RECT 7.970000  1.325000  8.230000 1.750000 ;
      RECT 7.970000  1.920000  8.230000 3.245000 ;
      RECT 8.400000  0.255000  8.660000 3.075000 ;
      RECT 8.830000  0.085000  9.090000 1.075000 ;
      RECT 8.830000  1.325000  9.090000 1.750000 ;
      RECT 8.830000  1.920000  9.090000 3.245000 ;
      RECT 9.260000  0.255000  9.520000 3.075000 ;
      RECT 9.690000  0.085000  9.985000 1.075000 ;
      RECT 9.690000  1.920000  9.985000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 2.915000  1.580000 3.085000 1.750000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.285000  1.950000 3.455000 2.120000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.715000  1.580000 3.885000 1.750000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.145000  1.950000 4.315000 2.120000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.575000  1.580000 4.745000 1.750000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.005000  1.950000 5.175000 2.120000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  1.580000 5.605000 1.750000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.865000  1.950000 6.035000 2.120000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.295000  1.580000 6.465000 1.750000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.725000  1.950000 6.895000 2.120000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.155000  1.580000 7.325000 1.750000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.585000  1.950000 7.755000 2.120000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.015000  1.580000 8.185000 1.750000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.445000  1.950000 8.615000 2.120000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 8.875000  1.580000 9.045000 1.750000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.305000  1.950000 9.475000 2.120000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
    LAYER met1 ;
      RECT 2.855000 1.550000 9.105000 1.780000 ;
  END
END sky130_fd_sc_lp__buf_16
END LIBRARY
