* File: sky130_fd_sc_lp__inputiso0p_lp.spice
* Created: Wed Sep  2 09:55:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__inputiso0p_lp.pex.spice"
.subckt sky130_fd_sc_lp__inputiso0p_lp  VNB VPB SLEEP A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* SLEEP	SLEEP
* VPB	VPB
* VNB	VNB
MM1012 A_112_93# N_SLEEP_M1012_g N_A_27_93#_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1155 PD=0.63 PS=1.39 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_SLEEP_M1006_g A_112_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.1323 AS=0.0441 PD=1.05 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1007 A_340_93# N_A_27_93#_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1323 PD=0.63 PS=1.05 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_342_489#_M1001_d N_A_M1001_g A_340_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_602_93# N_A_342_489#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_342_489#_M1004_g A_602_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_112_489# N_SLEEP_M1005_g N_A_27_93#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1155 PD=0.63 PS=1.39 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_SLEEP_M1002_g A_112_489# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1011 A_270_489# N_A_27_93#_M1011_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_342_489#_M1013_d N_A_27_93#_M1013_g A_270_489# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.063 AS=0.0441 PD=0.72 PS=0.63 NRD=9.3772 NRS=23.443 M=1 R=2.8
+ SA=75001.3 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 A_432_489# N_A_M1000_g N_A_342_489#_M1013_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.063 PD=0.63 PS=0.72 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g A_432_489# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09135 AS=0.0441 PD=0.8 PS=0.63 NRD=30.4759 NRS=23.443 M=1 R=2.8
+ SA=75002.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_602_367# N_A_342_489#_M1008_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.27405 PD=1.47 PS=2.4 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_X_M1009_d N_A_342_489#_M1009_g A_602_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.86097 P=12.16
c_32 VNB 0 1.49298e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__inputiso0p_lp.pxi.spice"
*
.ends
*
*
