* File: sky130_fd_sc_lp__o2111ai_lp.spice
* Created: Fri Aug 28 11:01:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111ai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o2111ai_lp  VNB VPB D1 C1 B1 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1002 A_167_57# N_D1_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1003 A_245_57# N_C1_M1003_g A_167_57# VNB NSHORT L=0.15 W=0.42 AD=0.0756
+ AS=0.0504 PD=0.78 PS=0.66 NRD=35.712 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_347_57#_M1007_d N_B1_M1007_g A_245_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0756 PD=0.84 PS=0.78 NRD=25.704 NRS=35.712 M=1 R=2.8 SA=75001.1
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_347_57#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0882 PD=0.81 PS=0.84 NRD=8.568 NRS=14.28 M=1 R=2.8 SA=75001.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_347_57#_M1005_d N_A1_M1005_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0819 PD=1.41 PS=0.81 NRD=0 NRS=22.848 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_D1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1004 N_VPWR_M1004_d N_C1_M1004_g N_Y_M1008_d VPB PHIGHVT L=0.25 W=1 AD=0.15
+ AS=0.14 PD=1.3 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_VPWR_M1004_d VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.15 PD=1.28 PS=1.3 NRD=0 NRS=3.9203 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1000 A_483_409# N_A2_M1000_g N_Y_M1006_d VPB PHIGHVT L=0.25 W=1 AD=0.125
+ AS=0.14 PD=1.25 PS=1.28 NRD=13.7703 NRS=0 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_483_409# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.125 PD=2.57 PS=1.25 NRD=0 NRS=13.7703 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o2111ai_lp.pxi.spice"
*
.ends
*
*
