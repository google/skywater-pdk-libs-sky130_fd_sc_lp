* NGSPICE file created from sky130_fd_sc_lp__dlygate4s50_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlygate4s50_1 A VGND VNB VPB VPWR X
M1000 X a_405_136# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=4.179e+11p ps=3.98e+06u
M1001 X a_405_136# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=5.292e+11p ps=4.82e+06u
M1002 VPWR A a_27_52# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 VGND A a_27_52# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 VGND a_288_52# a_405_136# VNB nshort w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 a_288_52# a_27_52# VGND VNB nshort w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 a_288_52# a_27_52# VPWR VPB phighvt w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 VPWR a_288_52# a_405_136# VPB phighvt w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

