* File: sky130_fd_sc_lp__o21a_0.pxi.spice
* Created: Fri Aug 28 11:03:33 2020
* 
x_PM_SKY130_FD_SC_LP__O21A_0%A_80_23# N_A_80_23#_M1002_s N_A_80_23#_M1006_d
+ N_A_80_23#_M1004_g N_A_80_23#_c_65_n N_A_80_23#_M1003_g N_A_80_23#_c_67_n
+ N_A_80_23#_c_68_n N_A_80_23#_c_69_n N_A_80_23#_c_70_n N_A_80_23#_c_76_n
+ N_A_80_23#_c_77_n N_A_80_23#_c_71_n N_A_80_23#_c_78_n N_A_80_23#_c_72_n
+ N_A_80_23#_c_73_n PM_SKY130_FD_SC_LP__O21A_0%A_80_23#
x_PM_SKY130_FD_SC_LP__O21A_0%B1 N_B1_M1006_g N_B1_c_136_n N_B1_M1002_g
+ N_B1_c_137_n N_B1_c_138_n N_B1_c_139_n N_B1_c_140_n B1 B1 N_B1_c_142_n
+ PM_SKY130_FD_SC_LP__O21A_0%B1
x_PM_SKY130_FD_SC_LP__O21A_0%A2 N_A2_c_189_n N_A2_M1005_g N_A2_M1007_g
+ N_A2_c_195_n A2 A2 A2 A2 A2 N_A2_c_192_n PM_SKY130_FD_SC_LP__O21A_0%A2
x_PM_SKY130_FD_SC_LP__O21A_0%A1 N_A1_M1000_g N_A1_M1001_g N_A1_c_241_n A1 A1 A1
+ N_A1_c_239_n PM_SKY130_FD_SC_LP__O21A_0%A1
x_PM_SKY130_FD_SC_LP__O21A_0%X N_X_M1004_s N_X_M1003_s N_X_c_266_n X X X X X X
+ PM_SKY130_FD_SC_LP__O21A_0%X
x_PM_SKY130_FD_SC_LP__O21A_0%VPWR N_VPWR_M1003_d N_VPWR_M1000_d N_VPWR_c_284_n
+ N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n VPWR N_VPWR_c_288_n
+ N_VPWR_c_289_n N_VPWR_c_283_n N_VPWR_c_291_n PM_SKY130_FD_SC_LP__O21A_0%VPWR
x_PM_SKY130_FD_SC_LP__O21A_0%VGND N_VGND_M1004_d N_VGND_M1007_d N_VGND_c_319_n
+ N_VGND_c_320_n N_VGND_c_321_n N_VGND_c_322_n VGND N_VGND_c_323_n
+ N_VGND_c_324_n N_VGND_c_325_n N_VGND_c_326_n PM_SKY130_FD_SC_LP__O21A_0%VGND
x_PM_SKY130_FD_SC_LP__O21A_0%A_300_58# N_A_300_58#_M1002_d N_A_300_58#_M1001_d
+ N_A_300_58#_c_356_n N_A_300_58#_c_357_n N_A_300_58#_c_358_n
+ N_A_300_58#_c_359_n PM_SKY130_FD_SC_LP__O21A_0%A_300_58#
cc_1 VNB N_A_80_23#_c_65_n 0.0259287f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.268
cc_2 VNB N_A_80_23#_M1003_g 0.012105f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.735
cc_3 VNB N_A_80_23#_c_67_n 0.0226118f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.445
cc_4 VNB N_A_80_23#_c_68_n 0.00201975f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.955
cc_5 VNB N_A_80_23#_c_69_n 0.00341193f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.045
cc_6 VNB N_A_80_23#_c_70_n 0.0149454f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.865
cc_7 VNB N_A_80_23#_c_71_n 0.00126444f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.5
cc_8 VNB N_A_80_23#_c_72_n 0.0199798f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.94
cc_9 VNB N_A_80_23#_c_73_n 0.0232126f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=0.775
cc_10 VNB N_B1_c_136_n 0.0197126f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.775
cc_11 VNB N_B1_c_137_n 0.00991137f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.268
cc_12 VNB N_B1_c_138_n 0.0215953f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.445
cc_13 VNB N_B1_c_139_n 0.00161501f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.735
cc_14 VNB N_B1_c_140_n 0.0243116f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.445
cc_15 VNB B1 0.00591959f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.045
cc_16 VNB N_B1_c_142_n 0.0162688f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.775
cc_17 VNB N_A2_c_189_n 0.0190996f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.415
cc_18 VNB N_A2_M1007_g 0.037458f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_19 VNB A2 0.00197008f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.445
cc_20 VNB N_A2_c_192_n 0.022237f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.775
cc_21 VNB N_A1_M1001_g 0.0669572f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.775
cc_22 VNB A1 0.0257391f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.445
cc_23 VNB N_A1_c_239_n 0.0126581f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.775
cc_24 VNB N_X_c_266_n 0.0131963f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_25 VNB X 0.0529411f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.445
cc_26 VNB N_VPWR_c_283_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.865
cc_27 VNB N_VGND_c_319_n 0.0100501f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_28 VNB N_VGND_c_320_n 0.00694515f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.735
cc_29 VNB N_VGND_c_321_n 0.0303431f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.445
cc_30 VNB N_VGND_c_322_n 0.00519339f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.955
cc_31 VNB N_VGND_c_323_n 0.0174373f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.865
cc_32 VNB N_VGND_c_324_n 0.021255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_325_n 0.183128f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.865
cc_34 VNB N_VGND_c_326_n 0.00545644f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=0.94
cc_35 VNB N_A_300_58#_c_356_n 0.00205974f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_36 VNB N_A_300_58#_c_357_n 0.021357f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.268
cc_37 VNB N_A_300_58#_c_358_n 0.00427031f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.445
cc_38 VNB N_A_300_58#_c_359_n 0.0207446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A_80_23#_M1003_g 0.0588771f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.735
cc_40 VPB N_A_80_23#_c_69_n 0.00734901f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.045
cc_41 VPB N_A_80_23#_c_76_n 0.0175838f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=2.13
cc_42 VPB N_A_80_23#_c_77_n 0.003178f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=2.13
cc_43 VPB N_A_80_23#_c_78_n 0.00328409f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=2.56
cc_44 VPB N_B1_M1006_g 0.0443381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_B1_c_139_n 0.0141528f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.735
cc_46 VPB B1 0.00329813f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.045
cc_47 VPB N_A2_c_189_n 0.00206317f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.415
cc_48 VPB N_A2_M1005_g 0.0383557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A2_c_195_n 0.0236254f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.268
cc_50 VPB A2 0.00391864f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.445
cc_51 VPB N_A1_M1000_g 0.0232723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A1_c_241_n 0.0748048f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.445
cc_53 VPB A1 0.0277195f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.445
cc_54 VPB N_A1_c_239_n 0.00488866f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=0.775
cc_55 VPB X 0.038769f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.445
cc_56 VPB X 0.0434734f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.94
cc_57 VPB N_VPWR_c_284_n 0.00926957f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.455
cc_58 VPB N_VPWR_c_285_n 0.032187f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.735
cc_59 VPB N_VPWR_c_286_n 0.0210228f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.445
cc_60 VPB N_VPWR_c_287_n 0.00516416f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.955
cc_61 VPB N_VPWR_c_288_n 0.0271332f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=0.5
cc_62 VPB N_VPWR_c_289_n 0.0190089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_283_n 0.0771187f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.865
cc_64 VPB N_VPWR_c_291_n 0.00541171f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=0.94
cc_65 N_A_80_23#_M1003_g N_B1_M1006_g 0.0265235f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_66 N_A_80_23#_c_69_n N_B1_M1006_g 0.00489886f $X=0.63 $Y=2.045 $X2=0 $Y2=0
cc_67 N_A_80_23#_c_76_n N_B1_M1006_g 0.0143858f $X=1.175 $Y=2.13 $X2=0 $Y2=0
cc_68 N_A_80_23#_c_78_n N_B1_M1006_g 0.0126839f $X=1.34 $Y=2.56 $X2=0 $Y2=0
cc_69 N_A_80_23#_c_70_n N_B1_c_136_n 5.75042e-19 $X=1.105 $Y=0.865 $X2=0 $Y2=0
cc_70 N_A_80_23#_c_71_n N_B1_c_136_n 0.00183047f $X=1.21 $Y=0.5 $X2=0 $Y2=0
cc_71 N_A_80_23#_c_72_n N_B1_c_136_n 5.47469e-19 $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_72 N_A_80_23#_c_65_n N_B1_c_137_n 0.00443633f $X=0.577 $Y=1.268 $X2=0 $Y2=0
cc_73 N_A_80_23#_M1003_g N_B1_c_138_n 0.0151861f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_74 N_A_80_23#_c_67_n N_B1_c_138_n 0.00830261f $X=0.577 $Y=1.445 $X2=0 $Y2=0
cc_75 N_A_80_23#_c_69_n N_B1_c_138_n 0.00222351f $X=0.63 $Y=2.045 $X2=0 $Y2=0
cc_76 N_A_80_23#_c_76_n N_B1_c_139_n 0.00128205f $X=1.175 $Y=2.13 $X2=0 $Y2=0
cc_77 N_A_80_23#_c_69_n N_B1_c_140_n 9.65908e-19 $X=0.63 $Y=2.045 $X2=0 $Y2=0
cc_78 N_A_80_23#_c_70_n N_B1_c_140_n 0.0115169f $X=1.105 $Y=0.865 $X2=0 $Y2=0
cc_79 N_A_80_23#_c_72_n N_B1_c_140_n 0.00443633f $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_80 N_A_80_23#_c_65_n B1 0.00119008f $X=0.577 $Y=1.268 $X2=0 $Y2=0
cc_81 N_A_80_23#_M1003_g B1 4.23935e-19 $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_82 N_A_80_23#_c_69_n B1 0.0390508f $X=0.63 $Y=2.045 $X2=0 $Y2=0
cc_83 N_A_80_23#_c_70_n B1 0.0292524f $X=1.105 $Y=0.865 $X2=0 $Y2=0
cc_84 N_A_80_23#_c_76_n B1 0.0228338f $X=1.175 $Y=2.13 $X2=0 $Y2=0
cc_85 N_A_80_23#_c_65_n N_B1_c_142_n 0.00830261f $X=0.577 $Y=1.268 $X2=0 $Y2=0
cc_86 N_A_80_23#_c_69_n N_B1_c_142_n 0.00117583f $X=0.63 $Y=2.045 $X2=0 $Y2=0
cc_87 N_A_80_23#_c_70_n N_B1_c_142_n 0.00129995f $X=1.105 $Y=0.865 $X2=0 $Y2=0
cc_88 N_A_80_23#_c_76_n N_A2_M1005_g 0.00133491f $X=1.175 $Y=2.13 $X2=0 $Y2=0
cc_89 N_A_80_23#_c_78_n N_A2_M1005_g 0.003844f $X=1.34 $Y=2.56 $X2=0 $Y2=0
cc_90 N_A_80_23#_c_76_n A2 0.0140495f $X=1.175 $Y=2.13 $X2=0 $Y2=0
cc_91 N_A_80_23#_c_78_n A2 0.0563579f $X=1.34 $Y=2.56 $X2=0 $Y2=0
cc_92 N_A_80_23#_M1003_g X 0.0108589f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_93 N_A_80_23#_c_68_n X 0.0146669f $X=0.63 $Y=0.955 $X2=0 $Y2=0
cc_94 N_A_80_23#_c_69_n X 0.0849547f $X=0.63 $Y=2.045 $X2=0 $Y2=0
cc_95 N_A_80_23#_c_77_n X 0.014744f $X=0.755 $Y=2.13 $X2=0 $Y2=0
cc_96 N_A_80_23#_c_73_n X 0.0236175f $X=0.577 $Y=0.775 $X2=0 $Y2=0
cc_97 N_A_80_23#_M1003_g X 9.24391e-19 $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_98 N_A_80_23#_c_77_n X 0.00526223f $X=0.755 $Y=2.13 $X2=0 $Y2=0
cc_99 N_A_80_23#_M1003_g N_VPWR_c_284_n 0.00296605f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_100 N_A_80_23#_c_76_n N_VPWR_c_284_n 0.0201589f $X=1.175 $Y=2.13 $X2=0 $Y2=0
cc_101 N_A_80_23#_c_77_n N_VPWR_c_284_n 0.00166412f $X=0.755 $Y=2.13 $X2=0 $Y2=0
cc_102 N_A_80_23#_c_78_n N_VPWR_c_284_n 0.0259861f $X=1.34 $Y=2.56 $X2=0 $Y2=0
cc_103 N_A_80_23#_c_78_n N_VPWR_c_285_n 0.00299946f $X=1.34 $Y=2.56 $X2=0 $Y2=0
cc_104 N_A_80_23#_M1003_g N_VPWR_c_286_n 0.00545548f $X=0.64 $Y=2.735 $X2=0
+ $Y2=0
cc_105 N_A_80_23#_c_78_n N_VPWR_c_288_n 0.017694f $X=1.34 $Y=2.56 $X2=0 $Y2=0
cc_106 N_A_80_23#_M1003_g N_VPWR_c_283_n 0.0112526f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_107 N_A_80_23#_c_78_n N_VPWR_c_283_n 0.00953185f $X=1.34 $Y=2.56 $X2=0 $Y2=0
cc_108 N_A_80_23#_c_68_n N_VGND_c_319_n 0.013994f $X=0.63 $Y=0.955 $X2=0 $Y2=0
cc_109 N_A_80_23#_c_70_n N_VGND_c_319_n 0.00802642f $X=1.105 $Y=0.865 $X2=0
+ $Y2=0
cc_110 N_A_80_23#_c_71_n N_VGND_c_319_n 0.0161745f $X=1.21 $Y=0.5 $X2=0 $Y2=0
cc_111 N_A_80_23#_c_72_n N_VGND_c_319_n 0.00132584f $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_112 N_A_80_23#_c_73_n N_VGND_c_319_n 0.0047323f $X=0.577 $Y=0.775 $X2=0 $Y2=0
cc_113 N_A_80_23#_c_71_n N_VGND_c_321_n 0.00983021f $X=1.21 $Y=0.5 $X2=0 $Y2=0
cc_114 N_A_80_23#_c_73_n N_VGND_c_323_n 0.00575161f $X=0.577 $Y=0.775 $X2=0
+ $Y2=0
cc_115 N_A_80_23#_c_68_n N_VGND_c_325_n 0.00291585f $X=0.63 $Y=0.955 $X2=0 $Y2=0
cc_116 N_A_80_23#_c_70_n N_VGND_c_325_n 0.00956759f $X=1.105 $Y=0.865 $X2=0
+ $Y2=0
cc_117 N_A_80_23#_c_71_n N_VGND_c_325_n 0.00884167f $X=1.21 $Y=0.5 $X2=0 $Y2=0
cc_118 N_A_80_23#_c_73_n N_VGND_c_325_n 0.0114421f $X=0.577 $Y=0.775 $X2=0 $Y2=0
cc_119 N_A_80_23#_c_70_n N_A_300_58#_c_356_n 0.00509314f $X=1.105 $Y=0.865 $X2=0
+ $Y2=0
cc_120 N_A_80_23#_c_71_n N_A_300_58#_c_356_n 0.0050507f $X=1.21 $Y=0.5 $X2=0
+ $Y2=0
cc_121 N_A_80_23#_c_70_n N_A_300_58#_c_358_n 0.0106968f $X=1.105 $Y=0.865 $X2=0
+ $Y2=0
cc_122 N_B1_c_138_n N_A2_c_189_n 0.0123095f $X=1.16 $Y=1.63 $X2=0 $Y2=0
cc_123 N_B1_c_136_n N_A2_M1007_g 0.0175973f $X=1.425 $Y=0.82 $X2=0 $Y2=0
cc_124 N_B1_c_137_n N_A2_M1007_g 0.00647097f $X=1.16 $Y=1.125 $X2=0 $Y2=0
cc_125 B1 N_A2_M1007_g 0.00106358f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B1_M1006_g N_A2_c_195_n 0.0263633f $X=1.125 $Y=2.735 $X2=0 $Y2=0
cc_127 N_B1_c_139_n N_A2_c_195_n 0.0123095f $X=1.16 $Y=1.795 $X2=0 $Y2=0
cc_128 N_B1_M1006_g A2 0.00181451f $X=1.125 $Y=2.735 $X2=0 $Y2=0
cc_129 B1 A2 0.038788f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_130 N_B1_c_142_n A2 7.51419e-19 $X=1.16 $Y=1.29 $X2=0 $Y2=0
cc_131 B1 N_A2_c_192_n 0.0038936f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_c_142_n N_A2_c_192_n 0.0123095f $X=1.16 $Y=1.29 $X2=0 $Y2=0
cc_133 N_B1_M1006_g N_VPWR_c_284_n 0.00282811f $X=1.125 $Y=2.735 $X2=0 $Y2=0
cc_134 N_B1_M1006_g N_VPWR_c_288_n 0.00511358f $X=1.125 $Y=2.735 $X2=0 $Y2=0
cc_135 N_B1_M1006_g N_VPWR_c_283_n 0.00973667f $X=1.125 $Y=2.735 $X2=0 $Y2=0
cc_136 N_B1_c_136_n N_VGND_c_319_n 0.00383707f $X=1.425 $Y=0.82 $X2=0 $Y2=0
cc_137 N_B1_c_136_n N_VGND_c_321_n 0.00531318f $X=1.425 $Y=0.82 $X2=0 $Y2=0
cc_138 N_B1_c_136_n N_VGND_c_325_n 0.0112385f $X=1.425 $Y=0.82 $X2=0 $Y2=0
cc_139 N_B1_c_136_n N_A_300_58#_c_356_n 0.00105525f $X=1.425 $Y=0.82 $X2=0 $Y2=0
cc_140 N_B1_c_137_n N_A_300_58#_c_358_n 9.9541e-19 $X=1.16 $Y=1.125 $X2=0 $Y2=0
cc_141 N_B1_c_140_n N_A_300_58#_c_358_n 0.00167046f $X=1.425 $Y=0.895 $X2=0
+ $Y2=0
cc_142 N_A2_M1007_g N_A1_M1001_g 0.0445528f $X=1.855 $Y=0.5 $X2=0 $Y2=0
cc_143 A2 N_A1_M1001_g 3.08094e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A2_M1005_g N_A1_c_241_n 0.0688243f $X=1.61 $Y=2.735 $X2=0 $Y2=0
cc_145 N_A2_c_195_n N_A1_c_241_n 0.0111341f $X=1.732 $Y=1.88 $X2=0 $Y2=0
cc_146 A2 N_A1_c_241_n 0.00759132f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A2_M1005_g A1 8.14066e-19 $X=1.61 $Y=2.735 $X2=0 $Y2=0
cc_148 N_A2_M1007_g A1 0.0056876f $X=1.855 $Y=0.5 $X2=0 $Y2=0
cc_149 A2 A1 0.085567f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_150 N_A2_c_189_n N_A1_c_239_n 0.00854244f $X=1.732 $Y=1.683 $X2=0 $Y2=0
cc_151 A2 N_A1_c_239_n 2.68989e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A2_M1005_g N_VPWR_c_285_n 0.00165403f $X=1.61 $Y=2.735 $X2=0 $Y2=0
cc_153 A2 N_VPWR_c_285_n 0.0213345f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A2_M1005_g N_VPWR_c_288_n 0.00429963f $X=1.61 $Y=2.735 $X2=0 $Y2=0
cc_155 A2 N_VPWR_c_288_n 0.00884202f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A2_M1005_g N_VPWR_c_283_n 0.00727785f $X=1.61 $Y=2.735 $X2=0 $Y2=0
cc_157 A2 N_VPWR_c_283_n 0.00848288f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_158 A2 A_337_483# 0.00116033f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_159 N_A2_M1007_g N_VGND_c_320_n 0.00329318f $X=1.855 $Y=0.5 $X2=0 $Y2=0
cc_160 N_A2_M1007_g N_VGND_c_321_n 0.00531318f $X=1.855 $Y=0.5 $X2=0 $Y2=0
cc_161 N_A2_M1007_g N_VGND_c_325_n 0.00568855f $X=1.855 $Y=0.5 $X2=0 $Y2=0
cc_162 N_A2_M1007_g N_A_300_58#_c_356_n 0.00183624f $X=1.855 $Y=0.5 $X2=0 $Y2=0
cc_163 N_A2_M1007_g N_A_300_58#_c_357_n 0.0144163f $X=1.855 $Y=0.5 $X2=0 $Y2=0
cc_164 A2 N_A_300_58#_c_357_n 0.00572326f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_165 A2 N_A_300_58#_c_358_n 0.0158148f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_166 N_A2_c_192_n N_A_300_58#_c_358_n 0.00401332f $X=1.73 $Y=1.375 $X2=0 $Y2=0
cc_167 N_A1_M1000_g N_VPWR_c_285_n 0.0138831f $X=1.97 $Y=2.735 $X2=0 $Y2=0
cc_168 N_A1_c_241_n N_VPWR_c_285_n 0.00777454f $X=2.335 $Y=2.12 $X2=0 $Y2=0
cc_169 A1 N_VPWR_c_285_n 0.0291329f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A1_M1000_g N_VPWR_c_288_n 0.00452967f $X=1.97 $Y=2.735 $X2=0 $Y2=0
cc_171 N_A1_M1000_g N_VPWR_c_283_n 0.00803025f $X=1.97 $Y=2.735 $X2=0 $Y2=0
cc_172 N_A1_M1001_g N_VGND_c_320_n 0.00329318f $X=2.285 $Y=0.5 $X2=0 $Y2=0
cc_173 N_A1_M1001_g N_VGND_c_324_n 0.00531318f $X=2.285 $Y=0.5 $X2=0 $Y2=0
cc_174 N_A1_M1001_g N_VGND_c_325_n 0.00634412f $X=2.285 $Y=0.5 $X2=0 $Y2=0
cc_175 N_A1_M1001_g N_A_300_58#_c_357_n 0.0132615f $X=2.285 $Y=0.5 $X2=0 $Y2=0
cc_176 A1 N_A_300_58#_c_357_n 0.0462163f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A1_c_239_n N_A_300_58#_c_357_n 6.14691e-19 $X=2.335 $Y=1.72 $X2=0 $Y2=0
cc_178 N_A1_M1001_g N_A_300_58#_c_359_n 0.00403984f $X=2.285 $Y=0.5 $X2=0 $Y2=0
cc_179 X N_VPWR_c_284_n 0.0313844f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_180 X N_VPWR_c_286_n 0.0342663f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_181 X N_VPWR_c_283_n 0.0185835f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_182 N_X_c_266_n N_VGND_c_323_n 0.0178269f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_183 N_X_M1004_s N_VGND_c_325_n 0.00212959f $X=0.135 $Y=0.245 $X2=0 $Y2=0
cc_184 N_X_c_266_n N_VGND_c_325_n 0.0120043f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_185 N_VGND_c_321_n N_A_300_58#_c_356_n 0.0096594f $X=1.935 $Y=0 $X2=0 $Y2=0
cc_186 N_VGND_c_325_n N_A_300_58#_c_356_n 0.0092367f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_187 N_VGND_c_320_n N_A_300_58#_c_357_n 0.0170782f $X=2.07 $Y=0.5 $X2=0 $Y2=0
cc_188 N_VGND_c_325_n N_A_300_58#_c_357_n 0.0105521f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_189 N_VGND_c_324_n N_A_300_58#_c_359_n 0.012454f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_190 N_VGND_c_325_n N_A_300_58#_c_359_n 0.0107265f $X=2.64 $Y=0 $X2=0 $Y2=0
