* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfstp_lp CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_750_108# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_2006_125# a_986_409# a_2206_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_1425_99# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VPWR SET_B a_2006_125# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 VPWR a_1199_419# a_1928_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VGND a_27_409# a_368_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_352_406# a_750_108# a_1199_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_2767_57# a_2006_125# a_2854_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_2767_57# a_2006_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_2584_57# a_2006_125# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_245_406# a_27_409# a_352_406# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 VPWR a_1199_419# a_1425_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_2854_57# a_2006_125# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1928_419# a_750_108# a_2006_125# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VGND a_2767_57# a_3012_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_352_406# a_986_409# a_1199_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_1001_108# a_750_108# a_986_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1736_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1371_419# a_1425_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X19 a_2124_66# a_2172_40# a_2202_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_27_409# SCE a_144_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_27_409# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_3012_57# a_2767_57# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_144_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_1383_125# a_1425_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_1199_419# a_1928_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR a_750_108# a_986_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 a_1425_99# a_1199_419# a_1736_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_2172_40# a_2006_125# a_2584_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_837_108# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_1199_419# a_986_409# a_1383_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VPWR SCD a_245_406# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X32 a_1928_125# a_986_409# a_2006_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 VPWR a_2767_57# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X34 a_2006_125# a_750_108# a_2124_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_352_406# D a_458_406# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X36 a_1199_419# a_750_108# a_1371_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X37 a_368_47# D a_352_406# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_352_406# SCE a_532_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_458_406# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X40 a_750_108# CLK a_837_108# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_2172_40# a_2006_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X42 a_2206_419# a_2172_40# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X43 a_532_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 VGND a_750_108# a_1001_108# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 a_2202_66# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
