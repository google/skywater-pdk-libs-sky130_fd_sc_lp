* File: sky130_fd_sc_lp__a21bo_0.spice
* Created: Fri Aug 28 09:49:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21bo_0.pex.spice"
.subckt sky130_fd_sc_lp__a21bo_0  VNB VPB B1_N A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_72_212#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_216_526#_M1008_d N_B1_N_M1008_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_72_212#_M1004_d N_A_216_526#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 A_533_52# N_A1_M1009_g N_A_72_212#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0588 PD=0.8 PS=0.7 NRD=38.568 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g A_533_52# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0798 PD=1.37 PS=0.8 NRD=0 NRS=38.568 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_72_212#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.130294 AS=0.1696 PD=1.22566 PS=1.81 NRD=7.683 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1005 N_A_216_526#_M1005_d N_B1_N_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0855057 PD=1.37 PS=0.80434 NRD=0 NRS=34.0022 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_467_458#_M1001_d N_A_216_526#_M1001_g N_A_72_212#_M1001_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_467_458#_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1003 N_A_467_458#_M1003_d N_A2_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a21bo_0.pxi.spice"
*
.ends
*
*
