* File: sky130_fd_sc_lp__a2bb2o_lp.pex.spice
* Created: Wed Sep  2 09:24:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%B2 3 7 11 12 13 15 22
r35 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.335 $X2=0.585 $Y2=1.335
r36 15 23 2.41001 $w=6.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.505
+ $X2=0.585 $Y2=1.505
r37 13 23 6.15891 $w=6.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.505
+ $X2=0.585 $Y2=1.505
r38 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.585 $Y=1.675
+ $X2=0.585 $Y2=1.335
r39 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.675
+ $X2=0.585 $Y2=1.84
r40 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.17
+ $X2=0.585 $Y2=1.335
r41 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.675 $Y=0.495
+ $X2=0.675 $Y2=1.17
r42 3 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.625 $Y=2.54 $X2=0.625
+ $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%B1 3 6 9 11 12 13 17
r45 17 19 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.167 $Y=1.335
+ $X2=1.167 $Y2=1.17
r46 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=1.295
+ $X2=1.18 $Y2=1.665
r47 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.18
+ $Y=1.335 $X2=1.18 $Y2=1.335
r48 9 11 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.155 $Y=2.54 $X2=1.155
+ $Y2=1.84
r49 6 11 31.6765 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=1.167 $Y=1.663
+ $X2=1.167 $Y2=1.84
r50 5 17 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=1.167 $Y=1.347
+ $X2=1.167 $Y2=1.335
r51 5 6 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=1.167 $Y=1.347
+ $X2=1.167 $Y2=1.663
r52 3 19 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.065 $Y=0.495
+ $X2=1.065 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%A_284_31# 1 2 7 9 10 11 13 16 18 20 23 24
+ 27 28 31 32 33 35 36 38 43 47
c112 28 0 4.19057e-20 $X=1.765 $Y=1.335
c113 27 0 1.45652e-19 $X=1.765 $Y=1.335
r114 43 45 6.46358 $w=6.04e-07 $l=3.2e-07 $layer=LI1_cond $X=4.43 $Y=2.58
+ $X2=4.43 $Y2=2.9
r115 42 43 7.87748 $w=6.04e-07 $l=3.9e-07 $layer=LI1_cond $X=4.43 $Y=2.19
+ $X2=4.43 $Y2=2.58
r116 38 40 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.21 $Y=0.58
+ $X2=4.21 $Y2=0.81
r117 35 42 10.3858 $w=6.04e-07 $l=3.22102e-07 $layer=LI1_cond $X=4.18 $Y=2.025
+ $X2=4.43 $Y2=2.19
r118 35 40 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=4.18 $Y=2.025
+ $X2=4.18 $Y2=0.81
r119 32 43 8.35964 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=4.095 $Y=2.58
+ $X2=4.43 $Y2=2.58
r120 32 33 140.92 $w=1.68e-07 $l=2.16e-06 $layer=LI1_cond $X=4.095 $Y=2.58
+ $X2=1.935 $Y2=2.58
r121 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.85 $Y=2.495
+ $X2=1.935 $Y2=2.58
r122 31 36 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.85 $Y=2.495
+ $X2=1.85 $Y2=1.84
r123 28 47 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.757 $Y=1.335
+ $X2=1.757 $Y2=1.17
r124 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.765
+ $Y=1.335 $X2=1.765 $Y2=1.335
r125 25 36 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=1.767 $Y=1.673
+ $X2=1.767 $Y2=1.84
r126 25 27 11.6276 $w=3.33e-07 $l=3.38e-07 $layer=LI1_cond $X=1.767 $Y=1.673
+ $X2=1.767 $Y2=1.335
r127 21 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.855 $Y=0.93
+ $X2=1.855 $Y2=0.855
r128 21 47 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.855 $Y=0.93
+ $X2=1.855 $Y2=1.17
r129 18 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.855 $Y=0.78
+ $X2=1.855 $Y2=0.855
r130 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.855 $Y=0.78
+ $X2=1.855 $Y2=0.495
r131 16 23 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.71 $Y=2.54 $X2=1.71
+ $Y2=1.84
r132 13 23 33.2433 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=1.757 $Y=1.668
+ $X2=1.757 $Y2=1.84
r133 12 28 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=1.757 $Y=1.342
+ $X2=1.757 $Y2=1.335
r134 12 13 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=1.757 $Y=1.342
+ $X2=1.757 $Y2=1.668
r135 10 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.78 $Y=0.855
+ $X2=1.855 $Y2=0.855
r136 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.78 $Y=0.855
+ $X2=1.57 $Y2=0.855
r137 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.495 $Y=0.78
+ $X2=1.57 $Y2=0.855
r138 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.495 $Y=0.78
+ $X2=1.495 $Y2=0.495
r139 2 45 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=2.045 $X2=4.6 $Y2=2.9
r140 2 42 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=2.045 $X2=4.6 $Y2=2.19
r141 1 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.07
+ $Y=0.37 $X2=4.21 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%A_63_57# 1 2 3 10 11 14 18 22 27 31 33 34
+ 37 39 40 43 48 49
c95 39 0 4.19057e-20 $X=2.307 $Y=1.182
r96 43 49 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.28 $Y=2.185
+ $X2=2.28 $Y2=1.66
r97 40 49 6.01482 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=2.307 $Y=1.468
+ $X2=2.307 $Y2=1.66
r98 39 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.335
+ $Y=1.155 $X2=2.335 $Y2=1.155
r99 39 40 8.56101 $w=3.83e-07 $l=2.86e-07 $layer=LI1_cond $X=2.307 $Y=1.182
+ $X2=2.307 $Y2=1.468
r100 35 39 12.4629 $w=2.32e-07 $l=3.14748e-07 $layer=LI1_cond $X=2.07 $Y=0.82
+ $X2=2.307 $Y2=1.001
r101 35 37 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.07 $Y=0.82
+ $X2=2.07 $Y2=0.495
r102 33 35 9.57122 $w=2.32e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.905 $Y=0.905
+ $X2=2.07 $Y2=0.82
r103 33 34 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=1.905 $Y=0.905
+ $X2=0.625 $Y2=0.905
r104 29 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.46 $Y=0.82
+ $X2=0.625 $Y2=0.905
r105 29 31 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.46 $Y=0.82
+ $X2=0.46 $Y2=0.495
r106 24 48 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.335 $Y=1.14
+ $X2=2.335 $Y2=1.155
r107 20 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.205 $Y=0.99
+ $X2=3.205 $Y2=1.065
r108 20 22 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.205 $Y=0.99
+ $X2=3.205 $Y2=0.58
r109 16 27 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=3.155 $Y=1.065
+ $X2=3.205 $Y2=1.065
r110 16 25 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=3.155 $Y=1.065
+ $X2=2.845 $Y2=1.065
r111 16 18 349.077 $w=2.5e-07 $l=1.405e-06 $layer=POLY_cond $X=3.155 $Y=1.14
+ $X2=3.155 $Y2=2.545
r112 12 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.845 $Y=0.99
+ $X2=2.845 $Y2=1.065
r113 12 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.845 $Y=0.99
+ $X2=2.845 $Y2=0.58
r114 11 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.5 $Y=1.065
+ $X2=2.335 $Y2=1.14
r115 10 25 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.77 $Y=1.065
+ $X2=2.845 $Y2=1.065
r116 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.77 $Y=1.065
+ $X2=2.5 $Y2=1.065
r117 3 43 600 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=2.04 $X2=2.28 $Y2=2.185
r118 2 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.285 $X2=2.07 $Y2=0.495
r119 1 31 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.315
+ $Y=0.285 $X2=0.46 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%A1_N 3 7 11 15 17 18 19 20 25
r43 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.725
+ $Y=1.345 $X2=3.725 $Y2=1.345
r44 19 20 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.687 $Y=1.665
+ $X2=3.687 $Y2=2.035
r45 19 26 9.10572 $w=4.03e-07 $l=3.2e-07 $layer=LI1_cond $X=3.687 $Y=1.665
+ $X2=3.687 $Y2=1.345
r46 18 26 1.42277 $w=4.03e-07 $l=5e-08 $layer=LI1_cond $X=3.687 $Y=1.295
+ $X2=3.687 $Y2=1.345
r47 16 25 40.6942 $w=4.1e-07 $l=3e-07 $layer=POLY_cond $X=3.765 $Y=1.645
+ $X2=3.765 $Y2=1.345
r48 16 17 36.2176 $w=4.1e-07 $l=2.05e-07 $layer=POLY_cond $X=3.765 $Y=1.645
+ $X2=3.765 $Y2=1.85
r49 15 25 2.03471 $w=4.1e-07 $l=1.5e-08 $layer=POLY_cond $X=3.765 $Y=1.33
+ $X2=3.765 $Y2=1.345
r50 7 17 172.675 $w=2.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.845 $Y=2.545
+ $X2=3.845 $Y2=1.85
r51 1 15 24.4548 $w=4.1e-07 $l=1.5e-07 $layer=POLY_cond $X=3.815 $Y=1.18
+ $X2=3.815 $Y2=1.33
r52 1 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.995 $Y=1.18 $X2=3.995
+ $Y2=0.58
r53 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.635 $Y=1.18 $X2=3.635
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%A2_N 1 3 7 11 13 15
r31 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.695
+ $Y=1.275 $X2=4.695 $Y2=1.275
r32 15 23 6.15891 $w=6.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.04 $Y=1.445
+ $X2=4.695 $Y2=1.445
r33 13 23 2.41001 $w=6.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.56 $Y=1.445
+ $X2=4.695 $Y2=1.445
r34 9 22 29.9477 $w=2.9e-07 $l=3.22102e-07 $layer=POLY_cond $X=4.785 $Y=1.11
+ $X2=4.535 $Y2=1.275
r35 9 11 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.785 $Y=1.11
+ $X2=4.785 $Y2=0.58
r36 5 22 29.9477 $w=2.9e-07 $l=2.13014e-07 $layer=POLY_cond $X=4.425 $Y=1.11
+ $X2=4.535 $Y2=1.275
r37 5 7 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.425 $Y=1.11
+ $X2=4.425 $Y2=0.58
r38 1 22 57.8488 $w=5.81e-07 $l=5.96678e-07 $layer=POLY_cond $X=4.335 $Y=1.78
+ $X2=4.535 $Y2=1.275
r39 1 3 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=4.335 $Y=1.78
+ $X2=4.335 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%A_43_408# 1 2 7 9 11 13 15
r33 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=2.19 $X2=1.42
+ $Y2=2.105
r34 13 15 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.42 $Y=2.19
+ $X2=1.42 $Y2=2.895
r35 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=2.105
+ $X2=0.36 $Y2=2.105
r36 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=2.105
+ $X2=1.42 $Y2=2.105
r37 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.255 $Y=2.105
+ $X2=0.525 $Y2=2.105
r38 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.36 $Y=2.19 $X2=0.36
+ $Y2=2.105
r39 7 9 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.36 $Y=2.19 $X2=0.36
+ $Y2=2.895
r40 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.28
+ $Y=2.04 $X2=1.42 $Y2=2.185
r41 2 15 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.28
+ $Y=2.04 $X2=1.42 $Y2=2.895
r42 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=2.04 $X2=0.36 $Y2=2.185
r43 1 9 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=2.04 $X2=0.36 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%VPWR 1 2 9 13 16 17 18 24 33 34 37
r45 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r46 34 38 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r48 31 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.5 $Y2=3.33
r49 31 33 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=5.04 $Y2=3.33
r50 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r51 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 26 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.5 $Y2=3.33
r55 24 29 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 18 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 18 27 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 16 21 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.89 $Y2=3.33
r62 15 26 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.89 $Y2=3.33
r64 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=3.33
r65 11 13 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.5 $Y=3.245
+ $X2=3.5 $Y2=2.92
r66 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245 $X2=0.89
+ $Y2=3.33
r67 7 9 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.89 $Y=3.245 $X2=0.89
+ $Y2=2.535
r68 2 13 600 $w=1.7e-07 $l=9.78839e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=2.045 $X2=3.5 $Y2=2.92
r69 1 9 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=0.75
+ $Y=2.04 $X2=0.89 $Y2=2.535
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%X 1 2 8 10 13
r30 15 17 4.38218 $w=3.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.765 $Y=2.122
+ $X2=2.89 $Y2=2.122
r31 13 17 8.06322 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=3.12 $Y=2.122
+ $X2=2.89 $Y2=2.122
r32 10 12 10.5346 $w=3.83e-07 $l=2.3e-07 $layer=LI1_cond $X=2.657 $Y=0.58
+ $X2=2.657 $Y2=0.81
r33 8 15 4.93978 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=2.765 $Y=1.92
+ $X2=2.765 $Y2=2.122
r34 8 12 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=2.765 $Y=1.92
+ $X2=2.765 $Y2=0.81
r35 2 17 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=2.045 $X2=2.89 $Y2=2.19
r36 1 10 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.37 $X2=2.63 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_LP%VGND 1 2 3 12 16 18 20 23 24 25 27 39 47
+ 51
r60 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r61 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r62 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r63 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r64 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r65 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r66 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r67 39 50 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5.057
+ $Y2=0
r68 39 44 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.56
+ $Y2=0
r69 38 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r70 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r71 35 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r72 34 37 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r73 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 32 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r75 32 34 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.68
+ $Y2=0
r76 30 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r77 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r78 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r79 27 29 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.72
+ $Y2=0
r80 25 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r81 25 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r82 23 37 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.12
+ $Y2=0
r83 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r84 22 41 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.6
+ $Y2=0
r85 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r86 18 50 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5 $Y=0.085
+ $X2=5.057 $Y2=0
r87 18 20 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.58
r88 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r89 14 16 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.58
r90 10 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r91 10 12 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.45
r92 3 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5 $Y2=0.58
r93 2 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.37 $X2=3.42 $Y2=0.58
r94 1 12 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.285 $X2=1.28 $Y2=0.45
.ends

