* File: sky130_fd_sc_lp__a311o_lp.pex.spice
* Created: Wed Sep  2 09:25:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311O_LP%A_85_21# 1 2 3 12 16 18 22 26 28 29 32 36
+ 38 42 46 51 52 53 55 56 57
c115 57 0 1.35038e-19 $X=3.995 $Y=0.935
c116 18 0 4.93603e-20 $X=0.63 $Y=2.57
r117 55 56 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.957 $Y=2.215
+ $X2=3.957 $Y2=2.05
r118 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.62
+ $Y=1.015 $X2=0.62 $Y2=1.015
r119 48 57 3.70735 $w=2.5e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.1 $Y=1.02
+ $X2=3.995 $Y2=0.935
r120 48 56 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=4.1 $Y=1.02
+ $X2=4.1 $Y2=2.05
r121 44 57 3.70735 $w=2.5e-07 $l=9.66954e-08 $layer=LI1_cond $X=3.97 $Y=0.85
+ $X2=3.995 $Y2=0.935
r122 44 46 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=3.97 $Y=0.85
+ $X2=3.97 $Y2=0.47
r123 40 55 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=3.957 $Y=2.277
+ $X2=3.957 $Y2=2.215
r124 40 42 16.3771 $w=4.53e-07 $l=6.23e-07 $layer=LI1_cond $X=3.957 $Y=2.277
+ $X2=3.957 $Y2=2.9
r125 39 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.555 $Y=0.935
+ $X2=2.39 $Y2=0.935
r126 38 57 2.76166 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=0.935
+ $X2=3.995 $Y2=0.935
r127 38 39 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.805 $Y=0.935
+ $X2=2.555 $Y2=0.935
r128 34 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=0.85
+ $X2=2.39 $Y2=0.935
r129 34 36 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.39 $Y=0.85
+ $X2=2.39 $Y2=0.47
r130 33 51 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=0.935
+ $X2=0.62 $Y2=0.935
r131 32 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=0.935
+ $X2=2.39 $Y2=0.935
r132 32 33 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.225 $Y=0.935
+ $X2=0.785 $Y2=0.935
r133 28 29 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.58 $Y=1.52
+ $X2=0.58 $Y2=1.76
r134 27 52 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=0.605 $Y=1.34
+ $X2=0.605 $Y2=1.015
r135 27 28 40.28 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.605 $Y=1.34
+ $X2=0.605 $Y2=1.52
r136 26 52 8.81592 $w=3.6e-07 $l=5.5e-08 $layer=POLY_cond $X=0.605 $Y=0.96
+ $X2=0.605 $Y2=1.015
r137 16 29 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.63 $Y=1.885
+ $X2=0.63 $Y2=1.76
r138 16 18 170.191 $w=2.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.63 $Y=1.885
+ $X2=0.63 $Y2=2.57
r139 10 26 25.8164 $w=3.6e-07 $l=1.5e-07 $layer=POLY_cond $X=0.68 $Y=0.81
+ $X2=0.68 $Y2=0.96
r140 10 22 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.86 $Y=0.81
+ $X2=0.86 $Y2=0.445
r141 10 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.5 $Y=0.81 $X2=0.5
+ $Y2=0.445
r142 3 55 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=2.07 $X2=3.895 $Y2=2.215
r143 3 42 400 $w=1.7e-07 $l=8.97274e-07 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=2.07 $X2=3.895 $Y2=2.9
r144 2 46 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.83
+ $Y=0.235 $X2=3.97 $Y2=0.47
r145 1 36 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.235 $X2=2.39 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_LP%A3 1 3 7 9 11 12 15 17 20 21
c53 7 0 1.12422e-19 $X=1.395 $Y=0.73
r54 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=1.365 $X2=1.16 $Y2=1.365
r55 17 21 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.16 $Y=1.665 $X2=1.16
+ $Y2=1.365
r56 13 15 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.25 $Y=0.805
+ $X2=1.395 $Y2=0.805
r57 12 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.16 $Y=1.705
+ $X2=1.16 $Y2=1.365
r58 11 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.2
+ $X2=1.16 $Y2=1.365
r59 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=0.73
+ $X2=1.395 $Y2=0.805
r60 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.395 $Y=0.73 $X2=1.395
+ $Y2=0.445
r61 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.25 $Y=0.88 $X2=1.25
+ $Y2=0.805
r62 5 11 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.25 $Y=0.88 $X2=1.25
+ $Y2=1.2
r63 1 12 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.87
+ $X2=1.16 $Y2=1.705
r64 1 3 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.16 $Y=1.87 $X2=1.16
+ $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_LP%A2 3 7 11 12 13 16 17
r45 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.7
+ $Y=1.365 $X2=1.7 $Y2=1.365
r46 13 17 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.7 $Y=1.665 $X2=1.7
+ $Y2=1.365
r47 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.7 $Y=1.705 $X2=1.7
+ $Y2=1.365
r48 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.705
+ $X2=1.7 $Y2=1.87
r49 10 16 45.2978 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.2 $X2=1.7
+ $Y2=1.365
r50 7 10 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.785 $Y=0.445
+ $X2=1.785 $Y2=1.2
r51 3 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.69 $Y=2.57 $X2=1.69
+ $Y2=1.87
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_LP%A1 3 7 10 12 13 14 15 16 20 22
c54 13 0 1.15418e-20 $X=2.177 $Y=0.88
r55 20 22 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=2.277 $Y=1.365
+ $X2=2.277 $Y2=1.2
r56 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.27
+ $Y=1.365 $X2=2.27 $Y2=1.365
r57 16 21 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.535
+ $X2=2.27 $Y2=1.535
r58 15 21 1.96371 $w=6.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.16 $Y=1.535
+ $X2=2.27 $Y2=1.535
r59 13 22 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.18 $Y=0.88
+ $X2=2.18 $Y2=1.2
r60 12 13 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=2.177 $Y=0.73
+ $X2=2.177 $Y2=0.88
r61 10 14 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.325 $Y=2.57
+ $X2=2.325 $Y2=1.87
r62 7 14 33.2433 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=2.277 $Y=1.698
+ $X2=2.277 $Y2=1.87
r63 6 20 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=2.277 $Y=1.372
+ $X2=2.277 $Y2=1.365
r64 6 7 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=2.277 $Y=1.372
+ $X2=2.277 $Y2=1.698
r65 3 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.175 $Y=0.445
+ $X2=2.175 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_LP%B1 1 3 8 10 12 16 18 19 20 21 27 28 29
r58 27 30 65.7961 $w=5.35e-07 $l=5.05e-07 $layer=POLY_cond $X=2.997 $Y=1.405
+ $X2=2.997 $Y2=1.91
r59 27 29 47.5561 $w=5.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.997 $Y=1.405
+ $X2=2.997 $Y2=1.24
r60 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.1
+ $Y=1.405 $X2=3.1 $Y2=1.405
r61 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=2.405 $X2=3.1
+ $Y2=2.775
r62 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=2.035 $X2=3.1
+ $Y2=2.405
r63 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=1.665 $X2=3.1
+ $Y2=2.035
r64 18 28 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=3.1 $Y=1.665 $X2=3.1
+ $Y2=1.405
r65 15 16 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.805 $Y=0.805
+ $X2=2.965 $Y2=0.805
r66 13 15 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.605 $Y=0.805
+ $X2=2.805 $Y2=0.805
r67 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.965 $Y=0.73
+ $X2=2.965 $Y2=0.805
r68 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.965 $Y=0.73
+ $X2=2.965 $Y2=0.445
r69 8 30 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.855 $Y=2.57
+ $X2=2.855 $Y2=1.91
r70 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.805 $Y=0.88
+ $X2=2.805 $Y2=0.805
r71 4 29 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.805 $Y=0.88
+ $X2=2.805 $Y2=1.24
r72 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.605 $Y=0.73
+ $X2=2.605 $Y2=0.805
r73 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.605 $Y=0.73 $X2=2.605
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_LP%C1 1 3 8 10 12 16 19 20 21 22 25 26
c48 25 0 1.35038e-19 $X=3.67 $Y=1.365
r49 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.67
+ $Y=1.365 $X2=3.67 $Y2=1.365
r50 22 26 9.87808 $w=3.48e-07 $l=3e-07 $layer=LI1_cond $X=3.66 $Y=1.665 $X2=3.66
+ $Y2=1.365
r51 20 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.67 $Y=1.705
+ $X2=3.67 $Y2=1.365
r52 20 21 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.705
+ $X2=3.67 $Y2=1.87
r53 19 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.2
+ $X2=3.67 $Y2=1.365
r54 15 16 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.58 $Y=0.805
+ $X2=3.755 $Y2=0.805
r55 13 15 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=3.395 $Y=0.805
+ $X2=3.58 $Y2=0.805
r56 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.755 $Y=0.73
+ $X2=3.755 $Y2=0.805
r57 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.755 $Y=0.73
+ $X2=3.755 $Y2=0.445
r58 8 21 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.63 $Y=2.57 $X2=3.63
+ $Y2=1.87
r59 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.58 $Y=0.88 $X2=3.58
+ $Y2=0.805
r60 4 19 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.58 $Y=0.88 $X2=3.58
+ $Y2=1.2
r61 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.395 $Y=0.73
+ $X2=3.395 $Y2=0.805
r62 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.395 $Y=0.73 $X2=3.395
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_LP%X 1 2 7 11 14 15 16 17
c29 17 0 1.12422e-19 $X=0.72 $Y=0.555
r30 21 23 0.284554 $w=4.03e-07 $l=1e-08 $layer=LI1_cond $X=0.275 $Y=0.467
+ $X2=0.285 $Y2=0.467
r31 16 21 2.48344 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.19 $Y=0.467
+ $X2=0.275 $Y2=0.467
r32 16 17 11.9513 $w=4.03e-07 $l=4.2e-07 $layer=LI1_cond $X=0.3 $Y=0.467
+ $X2=0.72 $Y2=0.467
r33 16 23 0.426831 $w=4.03e-07 $l=1.5e-08 $layer=LI1_cond $X=0.3 $Y=0.467
+ $X2=0.285 $Y2=0.467
r34 14 15 8.76046 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=0.317 $Y=2.215
+ $X2=0.317 $Y2=2.05
r35 9 14 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=0.317 $Y=2.262
+ $X2=0.317 $Y2=2.215
r36 9 11 17.3002 $w=4.23e-07 $l=6.38e-07 $layer=LI1_cond $X=0.317 $Y=2.262
+ $X2=0.317 $Y2=2.9
r37 7 16 5.93104 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.19 $Y=0.67 $X2=0.19
+ $Y2=0.467
r38 7 15 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.19 $Y=0.67
+ $X2=0.19 $Y2=2.05
r39 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=2.07 $X2=0.365 $Y2=2.215
r40 2 11 400 $w=1.7e-07 $l=8.99583e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=2.07 $X2=0.365 $Y2=2.9
r41 1 23 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.235 $X2=0.285 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_LP%VPWR 1 2 9 15 18 19 21 22 23 36 37
r48 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r49 33 36 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 27 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 23 37 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 23 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 23 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 21 30 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.79 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=3.33
+ $X2=1.955 $Y2=3.33
r58 20 33 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.12 $Y=3.33 $X2=2.16
+ $Y2=3.33
r59 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=3.33
+ $X2=1.955 $Y2=3.33
r60 18 26 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=0.73 $Y=3.33 $X2=0.72
+ $Y2=3.33
r61 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=3.33
+ $X2=0.895 $Y2=3.33
r62 17 30 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.895 $Y2=3.33
r64 13 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=3.245
+ $X2=1.955 $Y2=3.33
r65 13 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.955 $Y=3.245
+ $X2=1.955 $Y2=2.565
r66 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.895 $Y=2.215
+ $X2=0.895 $Y2=2.925
r67 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=3.245
+ $X2=0.895 $Y2=3.33
r68 7 12 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.895 $Y=3.245
+ $X2=0.895 $Y2=2.925
r69 2 15 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=1.815
+ $Y=2.07 $X2=1.955 $Y2=2.565
r70 1 12 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=2.07 $X2=0.895 $Y2=2.925
r71 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=2.07 $X2=0.895 $Y2=2.215
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_LP%A_257_414# 1 2 7 9 11 13 15
c36 7 0 4.93603e-20 $X=1.425 $Y=2.22
r37 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=2.22 $X2=2.59
+ $Y2=2.135
r38 13 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.59 $Y=2.22
+ $X2=2.59 $Y2=2.9
r39 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.59 $Y=2.135
+ $X2=1.425 $Y2=2.135
r40 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=2.135
+ $X2=2.59 $Y2=2.135
r41 11 12 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.425 $Y=2.135
+ $X2=1.59 $Y2=2.135
r42 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.425 $Y=2.22 $X2=1.425
+ $Y2=2.135
r43 7 9 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.425 $Y=2.22
+ $X2=1.425 $Y2=2.9
r44 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=2.07 $X2=2.59 $Y2=2.215
r45 2 15 400 $w=1.7e-07 $l=8.97274e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=2.07 $X2=2.59 $Y2=2.9
r46 1 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.285
+ $Y=2.07 $X2=1.425 $Y2=2.215
r47 1 9 400 $w=1.7e-07 $l=8.97274e-07 $layer=licon1_PDIFF $count=1 $X=1.285
+ $Y=2.07 $X2=1.425 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_LP%VGND 1 2 9 13 15 17 22 32 33 36 39
c62 22 0 1.15418e-20 $X=3.015 $Y=0
r63 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r64 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r65 33 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r66 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r67 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=0 $X2=3.18
+ $Y2=0
r68 30 32 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.345 $Y=0 $X2=4.08
+ $Y2=0
r69 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r70 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r71 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r72 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r73 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.18
+ $Y2=0
r75 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.68
+ $Y2=0
r76 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.18
+ $Y2=0
r77 22 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.015 $Y=0 $X2=2.64
+ $Y2=0
r78 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r79 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r80 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.18
+ $Y2=0
r81 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.72
+ $Y2=0
r82 15 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r83 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r84 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=0.085
+ $X2=3.18 $Y2=0
r85 11 13 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.18 $Y=0.085
+ $X2=3.18 $Y2=0.44
r86 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085 $X2=1.18
+ $Y2=0
r87 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.44
r88 2 13 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.04
+ $Y=0.235 $X2=3.18 $Y2=0.44
r89 1 9 182 $w=1.7e-07 $l=3.32039e-07 $layer=licon1_NDIFF $count=1 $X=0.935
+ $Y=0.235 $X2=1.18 $Y2=0.44
.ends

