* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2111o_lp A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_114_47# D1 a_27_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND D1 a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_436_47# a_27_409# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_27_409# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 VGND A2 a_868_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_27_409# C1 a_278_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_409# B1 a_710_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_27_409# D1 a_134_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_134_409# C1 a_232_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_739_409# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_278_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_232_409# B1 a_739_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_868_57# A1 a_27_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR A1 a_739_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VGND a_27_409# a_436_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_710_57# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
