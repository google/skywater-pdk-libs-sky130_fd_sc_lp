* NGSPICE file created from sky130_fd_sc_lp__nor4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
M1000 VGND A Y VNB nshort w=840000u l=150000u
+  ad=1.071e+12p pd=8.31e+06u as=5.082e+11p ps=4.57e+06u
M1001 VGND a_375_269# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR D_N a_27_508# VPB phighvt w=420000u l=150000u
+  ad=4.977e+11p pd=4.67e+06u as=1.113e+11p ps=1.37e+06u
M1003 a_375_269# C_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1004 a_333_367# a_27_508# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=3.339e+11p ps=3.05e+06u
M1005 a_513_367# B a_405_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.914e+11p pd=3.3e+06u as=4.914e+11p ps=3.3e+06u
M1006 VGND D_N a_27_508# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 Y B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A a_513_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_508# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_375_269# C_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 a_405_367# a_375_269# a_333_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

