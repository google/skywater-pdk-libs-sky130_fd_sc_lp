# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__clkbuflp_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.775000 0.695000 1.565000 ;
        RECT 0.125000 1.565000 0.370000 1.805000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.010000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.805000 1.920000 11.555000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.480000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.480000 0.085000 ;
      RECT  0.000000  3.245000 12.480000 3.415000 ;
      RECT  0.095000  2.065000  0.425000 3.245000 ;
      RECT  0.125000  0.085000  0.425000 0.605000 ;
      RECT  0.595000  2.015000  1.055000 3.075000 ;
      RECT  0.885000  0.265000  1.230000 1.205000 ;
      RECT  0.885000  1.205000  3.910000 1.535000 ;
      RECT  0.885000  1.535000  1.055000 2.015000 ;
      RECT  1.225000  2.065000  1.485000 3.245000 ;
      RECT  1.675000  0.085000  2.005000 0.605000 ;
      RECT  1.685000  1.535000  2.015000 3.075000 ;
      RECT  2.215000  2.085000  2.545000 3.245000 ;
      RECT  2.450000  0.265000  2.795000 1.180000 ;
      RECT  2.450000  1.180000  3.910000 1.205000 ;
      RECT  2.745000  1.535000  3.075000 3.075000 ;
      RECT  3.255000  0.085000  3.585000 0.605000 ;
      RECT  3.275000  2.085000  3.605000 3.245000 ;
      RECT  3.805000  1.705000  4.395000 1.875000 ;
      RECT  3.805000  1.875000  4.135000 3.075000 ;
      RECT  4.065000  0.265000  4.395000 1.035000 ;
      RECT  4.080000  1.035000  4.395000 1.705000 ;
      RECT  4.335000  2.085000  4.665000 3.245000 ;
      RECT  4.585000  1.180000  5.390000 1.510000 ;
      RECT  4.855000  0.085000  5.185000 0.605000 ;
      RECT  4.865000  1.920000  5.195000 3.075000 ;
      RECT  5.395000  2.085000  5.725000 3.245000 ;
      RECT  5.645000  0.265000  5.975000 1.170000 ;
      RECT  5.645000  1.170000  6.255000 1.790000 ;
      RECT  5.925000  1.790000  6.255000 3.075000 ;
      RECT  6.435000  0.085000  6.765000 0.605000 ;
      RECT  6.455000  2.085000  6.785000 3.245000 ;
      RECT  6.470000  1.180000  6.800000 1.510000 ;
      RECT  6.985000  1.170000  7.555000 1.790000 ;
      RECT  6.985000  1.790000  7.315000 3.075000 ;
      RECT  7.225000  0.265000  7.555000 1.170000 ;
      RECT  7.515000  2.085000  7.845000 3.245000 ;
      RECT  7.750000  1.180000  8.555000 1.510000 ;
      RECT  8.015000  0.085000  8.345000 0.605000 ;
      RECT  8.045000  1.920000  8.375000 3.075000 ;
      RECT  8.575000  2.085000  8.905000 3.245000 ;
      RECT  8.805000  0.265000  9.135000 1.170000 ;
      RECT  8.805000  1.170000  9.435000 1.790000 ;
      RECT  9.105000  1.790000  9.435000 3.075000 ;
      RECT  9.595000  0.085000  9.925000 0.605000 ;
      RECT  9.635000  2.085000  9.965000 3.245000 ;
      RECT  9.650000  1.180000  9.980000 1.510000 ;
      RECT 10.165000  1.170000 10.715000 1.790000 ;
      RECT 10.165000  1.790000 10.495000 3.075000 ;
      RECT 10.385000  0.265000 10.715000 1.170000 ;
      RECT 10.695000  2.085000 11.025000 3.245000 ;
      RECT 10.910000  1.180000 11.920000 1.510000 ;
      RECT 11.175000  0.085000 11.505000 0.605000 ;
      RECT 11.225000  1.920000 11.555000 3.075000 ;
      RECT 11.755000  2.085000 12.085000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.210000  3.205000 1.380000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  1.210000  3.685000 1.380000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.885000  1.950000  4.055000 2.120000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.210000  5.125000 1.380000 ;
      RECT  4.955000  1.950000  5.125000 2.120000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.005000  1.950000  6.175000 2.120000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.550000  1.210000  6.720000 1.380000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.070000  1.950000  7.240000 2.120000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.210000  8.005000 1.380000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.130000  1.950000  8.300000 2.120000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.210000  8.485000 1.380000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.190000  1.950000  9.360000 2.120000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.210000  9.925000 1.380000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  1.950000 10.405000 2.120000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  1.210000 11.365000 1.380000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.305000  1.950000 11.475000 2.120000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  1.210000 11.845000 1.380000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
    LAYER met1 ;
      RECT 2.975000 1.180000 11.905000 1.410000 ;
  END
END sky130_fd_sc_lp__clkbuflp_16
END LIBRARY
