* File: sky130_fd_sc_lp__nor4_4.pxi.spice
* Created: Fri Aug 28 10:57:42 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4_4%A N_A_M1002_g N_A_c_117_n N_A_M1004_g N_A_M1006_g
+ N_A_c_119_n N_A_M1011_g N_A_M1014_g N_A_c_121_n N_A_M1012_g N_A_M1019_g
+ N_A_c_123_n N_A_M1023_g A A A A N_A_c_124_n N_A_c_125_n N_A_c_126_n
+ PM_SKY130_FD_SC_LP__NOR4_4%A
x_PM_SKY130_FD_SC_LP__NOR4_4%B N_B_c_200_n N_B_M1009_g N_B_c_201_n N_B_M1020_g
+ N_B_c_194_n N_B_M1005_g N_B_c_202_n N_B_M1022_g N_B_c_195_n N_B_M1015_g
+ N_B_c_203_n N_B_M1031_g N_B_c_196_n N_B_M1026_g N_B_c_197_n N_B_M1028_g B B
+ N_B_c_198_n N_B_c_199_n PM_SKY130_FD_SC_LP__NOR4_4%B
x_PM_SKY130_FD_SC_LP__NOR4_4%C N_C_c_277_n N_C_M1007_g N_C_M1003_g N_C_c_279_n
+ N_C_M1018_g N_C_M1010_g N_C_c_281_n N_C_M1024_g N_C_M1017_g N_C_c_283_n
+ N_C_M1030_g N_C_M1025_g C C C N_C_c_286_n PM_SKY130_FD_SC_LP__NOR4_4%C
x_PM_SKY130_FD_SC_LP__NOR4_4%D N_D_M1013_g N_D_M1000_g N_D_M1016_g N_D_M1001_g
+ N_D_M1027_g N_D_M1008_g N_D_M1029_g N_D_M1021_g N_D_c_418_p D D N_D_c_374_n
+ N_D_c_375_n D N_D_c_376_n PM_SKY130_FD_SC_LP__NOR4_4%D
x_PM_SKY130_FD_SC_LP__NOR4_4%A_72_367# N_A_72_367#_M1002_d N_A_72_367#_M1006_d
+ N_A_72_367#_M1019_d N_A_72_367#_M1020_d N_A_72_367#_M1031_d
+ N_A_72_367#_c_454_n N_A_72_367#_c_455_n N_A_72_367#_c_460_n
+ N_A_72_367#_c_486_p N_A_72_367#_c_464_n N_A_72_367#_c_468_n
+ N_A_72_367#_c_489_p N_A_72_367#_c_471_n N_A_72_367#_c_473_n
+ N_A_72_367#_c_478_n N_A_72_367#_c_456_n N_A_72_367#_c_457_n
+ N_A_72_367#_c_469_n N_A_72_367#_c_480_n PM_SKY130_FD_SC_LP__NOR4_4%A_72_367#
x_PM_SKY130_FD_SC_LP__NOR4_4%VPWR N_VPWR_M1002_s N_VPWR_M1014_s N_VPWR_c_518_n
+ N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n VPWR
+ N_VPWR_c_523_n N_VPWR_c_517_n N_VPWR_c_525_n PM_SKY130_FD_SC_LP__NOR4_4%VPWR
x_PM_SKY130_FD_SC_LP__NOR4_4%A_499_367# N_A_499_367#_M1009_s
+ N_A_499_367#_M1022_s N_A_499_367#_M1003_d N_A_499_367#_M1017_d
+ N_A_499_367#_c_645_n N_A_499_367#_c_622_n N_A_499_367#_c_617_n
+ N_A_499_367#_c_648_n N_A_499_367#_c_618_n N_A_499_367#_c_659_p
+ N_A_499_367#_c_619_n N_A_499_367#_c_662_p N_A_499_367#_c_632_n
+ N_A_499_367#_c_620_n PM_SKY130_FD_SC_LP__NOR4_4%A_499_367#
x_PM_SKY130_FD_SC_LP__NOR4_4%A_864_367# N_A_864_367#_M1003_s
+ N_A_864_367#_M1010_s N_A_864_367#_M1025_s N_A_864_367#_M1001_s
+ N_A_864_367#_M1021_s N_A_864_367#_c_665_n N_A_864_367#_c_666_n
+ N_A_864_367#_c_672_n N_A_864_367#_c_674_n N_A_864_367#_c_678_n
+ N_A_864_367#_c_680_n N_A_864_367#_c_689_n N_A_864_367#_c_691_n
+ N_A_864_367#_c_695_n N_A_864_367#_c_667_n N_A_864_367#_c_668_n
+ N_A_864_367#_c_683_n N_A_864_367#_c_685_n N_A_864_367#_c_701_n
+ PM_SKY130_FD_SC_LP__NOR4_4%A_864_367#
x_PM_SKY130_FD_SC_LP__NOR4_4%Y N_Y_M1004_d N_Y_M1012_d N_Y_M1005_s N_Y_M1026_s
+ N_Y_M1007_d N_Y_M1024_d N_Y_M1013_s N_Y_M1027_s N_Y_M1000_d N_Y_M1008_d
+ N_Y_c_848_p N_Y_c_745_n N_Y_c_746_n N_Y_c_854_p N_Y_c_763_n N_Y_c_851_p
+ N_Y_c_771_n N_Y_c_849_p N_Y_c_775_n N_Y_c_850_p N_Y_c_784_n N_Y_c_844_p
+ N_Y_c_788_n N_Y_c_852_p N_Y_c_825_n N_Y_c_747_n N_Y_c_751_n N_Y_c_752_n
+ N_Y_c_853_p N_Y_c_828_n N_Y_c_748_n N_Y_c_753_n N_Y_c_749_n N_Y_c_778_n
+ N_Y_c_780_n N_Y_c_790_n N_Y_c_792_n N_Y_c_813_n N_Y_c_754_n Y
+ PM_SKY130_FD_SC_LP__NOR4_4%Y
x_PM_SKY130_FD_SC_LP__NOR4_4%VGND N_VGND_M1004_s N_VGND_M1011_s N_VGND_M1023_s
+ N_VGND_M1015_d N_VGND_M1028_d N_VGND_M1018_s N_VGND_M1030_s N_VGND_M1016_d
+ N_VGND_M1029_d N_VGND_c_872_n N_VGND_c_873_n N_VGND_c_874_n N_VGND_c_875_n
+ N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n N_VGND_c_879_n N_VGND_c_880_n
+ N_VGND_c_881_n N_VGND_c_882_n N_VGND_c_883_n N_VGND_c_884_n N_VGND_c_885_n
+ N_VGND_c_886_n N_VGND_c_887_n N_VGND_c_888_n N_VGND_c_889_n VGND
+ N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n N_VGND_c_894_n
+ N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n N_VGND_c_898_n
+ PM_SKY130_FD_SC_LP__NOR4_4%VGND
cc_1 VNB N_A_M1002_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.465
cc_2 VNB N_A_c_117_n 0.0214749f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.185
cc_3 VNB N_A_M1006_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=2.465
cc_4 VNB N_A_c_119_n 0.015136f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.185
cc_5 VNB N_A_M1014_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=2.465
cc_6 VNB N_A_c_121_n 0.015136f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.185
cc_7 VNB N_A_M1019_g 0.00123444f $X=-0.19 $Y=-0.245 $X2=1.99 $Y2=2.465
cc_8 VNB N_A_c_123_n 0.021212f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.185
cc_9 VNB N_A_c_124_n 0.0765425f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.405
cc_10 VNB N_A_c_125_n 0.0152569f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.46
cc_11 VNB N_A_c_126_n 0.0957194f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.405
cc_12 VNB N_B_c_194_n 0.0212715f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=0.655
cc_13 VNB N_B_c_195_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.655
cc_14 VNB N_B_c_196_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.185
cc_15 VNB N_B_c_197_n 0.016201f $X=-0.19 $Y=-0.245 $X2=1.99 $Y2=1.625
cc_16 VNB N_B_c_198_n 0.148412f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_17 VNB N_B_c_199_n 0.00528532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C_c_277_n 0.016201f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.625
cc_19 VNB N_C_M1003_g 0.0092958f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=0.655
cc_20 VNB N_C_c_279_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.625
cc_21 VNB N_C_M1010_g 0.00691852f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.655
cc_22 VNB N_C_c_281_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=1.625
cc_23 VNB N_C_M1017_g 0.00691852f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=0.655
cc_24 VNB N_C_c_283_n 0.016201f $X=-0.19 $Y=-0.245 $X2=1.99 $Y2=1.625
cc_25 VNB N_C_M1025_g 0.00712556f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.655
cc_26 VNB C 0.0130403f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_27 VNB N_C_c_286_n 0.0763278f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.46
cc_28 VNB N_D_M1013_g 0.0203018f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.465
cc_29 VNB N_D_M1000_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=0.655
cc_30 VNB N_D_M1016_g 0.0200323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_D_M1001_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=1.625
cc_32 VNB N_D_M1027_g 0.0204894f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.185
cc_33 VNB N_D_M1008_g 0.00249019f $X=-0.19 $Y=-0.245 $X2=1.99 $Y2=2.465
cc_34 VNB N_D_M1029_g 0.0235981f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.655
cc_35 VNB N_D_M1021_g 0.00268533f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_36 VNB N_D_c_374_n 0.0786635f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.405
cc_37 VNB N_D_c_375_n 0.00574211f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.46
cc_38 VNB N_D_c_376_n 0.0021425f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.547
cc_39 VNB N_VPWR_c_517_n 0.342803f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_40 VNB N_Y_c_745_n 0.00303808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_746_n 0.00290472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_747_n 0.00306427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_748_n 0.0106203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_749_n 0.00240588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB Y 0.0237196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_872_n 0.0399184f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_47 VNB N_VGND_c_873_n 3.13331e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_874_n 3.09829e-19 $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_49 VNB N_VGND_c_875_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.405
cc_50 VNB N_VGND_c_876_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.405
cc_51 VNB N_VGND_c_877_n 0.012974f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.405
cc_52 VNB N_VGND_c_878_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.99 $Y2=1.405
cc_53 VNB N_VGND_c_879_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_880_n 0.0108441f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.547
cc_55 VNB N_VGND_c_881_n 0.0261041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_882_n 0.0145539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_883_n 0.0058666f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.547
cc_58 VNB N_VGND_c_884_n 0.0145469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_885_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.547
cc_60 VNB N_VGND_c_886_n 0.012974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_887_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_888_n 0.012974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_889_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_890_n 0.0130811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_891_n 0.012974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_892_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_893_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_894_n 0.0148602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_895_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_896_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_897_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_898_n 0.399827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VPB N_A_M1002_g 0.0254689f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.465
cc_74 VPB N_A_M1006_g 0.0188311f $X=-0.19 $Y=1.655 $X2=1.13 $Y2=2.465
cc_75 VPB N_A_M1014_g 0.0188311f $X=-0.19 $Y=1.655 $X2=1.56 $Y2=2.465
cc_76 VPB N_A_M1019_g 0.019032f $X=-0.19 $Y=1.655 $X2=1.99 $Y2=2.465
cc_77 VPB N_A_c_125_n 0.0243168f $X=-0.19 $Y=1.655 $X2=1.97 $Y2=1.46
cc_78 VPB N_B_c_200_n 0.0164031f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.625
cc_79 VPB N_B_c_201_n 0.0152515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_B_c_202_n 0.0152515f $X=-0.19 $Y=1.655 $X2=1.13 $Y2=2.465
cc_81 VPB N_B_c_203_n 0.0195571f $X=-0.19 $Y=1.655 $X2=1.56 $Y2=2.465
cc_82 VPB N_B_c_198_n 0.0240097f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_83 VPB N_C_M1003_g 0.0248182f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=0.655
cc_84 VPB N_C_M1010_g 0.018695f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=0.655
cc_85 VPB N_C_M1017_g 0.018695f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=0.655
cc_86 VPB N_C_M1025_g 0.0201271f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.655
cc_87 VPB N_D_M1000_g 0.0201244f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=0.655
cc_88 VPB N_D_M1001_g 0.0186114f $X=-0.19 $Y=1.655 $X2=1.56 $Y2=1.625
cc_89 VPB N_D_M1008_g 0.0185925f $X=-0.19 $Y=1.655 $X2=1.99 $Y2=2.465
cc_90 VPB N_D_M1021_g 0.023518f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_91 VPB N_A_72_367#_c_454_n 0.00743726f $X=-0.19 $Y=1.655 $X2=1.56 $Y2=2.465
cc_92 VPB N_A_72_367#_c_455_n 0.0369481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_72_367#_c_456_n 0.0018321f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.405
cc_94 VPB N_A_72_367#_c_457_n 0.00777165f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_95 VPB N_VPWR_c_518_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.13 $Y2=2.465
cc_96 VPB N_VPWR_c_519_n 0.012974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_520_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.56 $Y2=1.625
cc_98 VPB N_VPWR_c_521_n 0.0225828f $X=-0.19 $Y=1.655 $X2=1.56 $Y2=2.465
cc_99 VPB N_VPWR_c_522_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_523_n 0.144209f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_101 VPB N_VPWR_c_517_n 0.0641831f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_102 VPB N_VPWR_c_525_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_499_367#_c_617_n 0.00109676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_499_367#_c_618_n 0.0170883f $X=-0.19 $Y=1.655 $X2=1.99 $Y2=2.465
cc_105 VPB N_A_499_367#_c_619_n 0.00591333f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_106 VPB N_A_499_367#_c_620_n 0.00146483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_864_367#_c_665_n 0.00189498f $X=-0.19 $Y=1.655 $X2=1.56 $Y2=2.465
cc_108 VPB N_A_864_367#_c_666_n 0.00786202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_864_367#_c_667_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_110 VPB N_A_864_367#_c_668_n 0.0332384f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.405
cc_111 VPB N_Y_c_751_n 0.0030392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_Y_c_752_n 0.0030854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_Y_c_753_n 0.0107706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_Y_c_754_n 0.00143206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB Y 0.00198241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 N_A_M1019_g N_B_c_198_n 0.0197728f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_c_125_n N_B_c_198_n 0.00355017f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_118 N_A_c_126_n N_B_c_198_n 0.0296078f $X=2.06 $Y=1.405 $X2=0 $Y2=0
cc_119 N_A_c_125_n N_B_c_199_n 0.0134142f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_120 N_A_c_126_n N_B_c_199_n 0.00126268f $X=2.06 $Y=1.405 $X2=0 $Y2=0
cc_121 N_A_c_124_n N_A_72_367#_c_454_n 0.00148159f $X=0.625 $Y=1.405 $X2=0 $Y2=0
cc_122 N_A_c_125_n N_A_72_367#_c_454_n 0.0224133f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_123 N_A_M1002_g N_A_72_367#_c_460_n 0.0122595f $X=0.7 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_M1006_g N_A_72_367#_c_460_n 0.0122595f $X=1.13 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_c_125_n N_A_72_367#_c_460_n 0.0436322f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_126 N_A_c_126_n N_A_72_367#_c_460_n 5.1019e-19 $X=2.06 $Y=1.405 $X2=0 $Y2=0
cc_127 N_A_M1014_g N_A_72_367#_c_464_n 0.0122129f $X=1.56 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_M1019_g N_A_72_367#_c_464_n 0.0122595f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A_c_125_n N_A_72_367#_c_464_n 0.0436322f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_130 N_A_c_126_n N_A_72_367#_c_464_n 5.1019e-19 $X=2.06 $Y=1.405 $X2=0 $Y2=0
cc_131 N_A_c_125_n N_A_72_367#_c_468_n 0.00166155f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_132 N_A_c_125_n N_A_72_367#_c_469_n 0.0156438f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_133 N_A_c_126_n N_A_72_367#_c_469_n 5.77956e-19 $X=2.06 $Y=1.405 $X2=0 $Y2=0
cc_134 N_A_M1002_g N_VPWR_c_518_n 0.0163935f $X=0.7 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_M1006_g N_VPWR_c_518_n 0.0142502f $X=1.13 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_M1014_g N_VPWR_c_518_n 6.85495e-19 $X=1.56 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_M1006_g N_VPWR_c_519_n 0.00486043f $X=1.13 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A_M1014_g N_VPWR_c_519_n 0.00486043f $X=1.56 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_M1006_g N_VPWR_c_520_n 6.85495e-19 $X=1.13 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A_M1014_g N_VPWR_c_520_n 0.0147919f $X=1.56 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_M1019_g N_VPWR_c_520_n 0.015973f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_M1002_g N_VPWR_c_521_n 0.00486043f $X=0.7 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_M1019_g N_VPWR_c_523_n 0.00486043f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_M1002_g N_VPWR_c_517_n 0.00933443f $X=0.7 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1006_g N_VPWR_c_517_n 0.00824727f $X=1.13 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_M1014_g N_VPWR_c_517_n 0.00824727f $X=1.56 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_M1019_g N_VPWR_c_517_n 0.0082726f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_c_125_n N_A_499_367#_c_617_n 0.00225308f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_149 N_A_c_119_n N_Y_c_745_n 0.0131987f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_150 N_A_c_121_n N_Y_c_745_n 0.0131251f $X=1.63 $Y=1.185 $X2=0 $Y2=0
cc_151 N_A_c_125_n N_Y_c_745_n 0.0499599f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_152 N_A_c_126_n N_Y_c_745_n 0.00309344f $X=2.06 $Y=1.405 $X2=0 $Y2=0
cc_153 N_A_c_117_n N_Y_c_746_n 0.00281332f $X=0.77 $Y=1.185 $X2=0 $Y2=0
cc_154 N_A_c_125_n N_Y_c_746_n 0.0183905f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_155 N_A_c_126_n N_Y_c_746_n 0.00321567f $X=2.06 $Y=1.405 $X2=0 $Y2=0
cc_156 N_A_c_123_n N_Y_c_763_n 0.0150307f $X=2.06 $Y=1.185 $X2=0 $Y2=0
cc_157 N_A_c_125_n N_Y_c_763_n 0.00789415f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_158 N_A_c_123_n N_Y_c_749_n 0.00313693f $X=2.06 $Y=1.185 $X2=0 $Y2=0
cc_159 N_A_c_125_n N_Y_c_749_n 0.0153962f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_160 N_A_c_126_n N_Y_c_749_n 0.00321567f $X=2.06 $Y=1.405 $X2=0 $Y2=0
cc_161 N_A_c_117_n N_VGND_c_872_n 0.00712293f $X=0.77 $Y=1.185 $X2=0 $Y2=0
cc_162 N_A_c_124_n N_VGND_c_872_n 0.00886009f $X=0.625 $Y=1.405 $X2=0 $Y2=0
cc_163 N_A_c_125_n N_VGND_c_872_n 0.0193926f $X=1.97 $Y=1.46 $X2=0 $Y2=0
cc_164 N_A_c_117_n N_VGND_c_873_n 6.24197e-19 $X=0.77 $Y=1.185 $X2=0 $Y2=0
cc_165 N_A_c_119_n N_VGND_c_873_n 0.0102349f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A_c_121_n N_VGND_c_873_n 0.0101747f $X=1.63 $Y=1.185 $X2=0 $Y2=0
cc_167 N_A_c_123_n N_VGND_c_873_n 6.13597e-19 $X=2.06 $Y=1.185 $X2=0 $Y2=0
cc_168 N_A_c_117_n N_VGND_c_884_n 0.00583607f $X=0.77 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A_c_119_n N_VGND_c_884_n 0.00486043f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_170 N_A_c_121_n N_VGND_c_893_n 0.00486043f $X=1.63 $Y=1.185 $X2=0 $Y2=0
cc_171 N_A_c_123_n N_VGND_c_893_n 0.00486043f $X=2.06 $Y=1.185 $X2=0 $Y2=0
cc_172 N_A_c_121_n N_VGND_c_894_n 5.92296e-19 $X=1.63 $Y=1.185 $X2=0 $Y2=0
cc_173 N_A_c_123_n N_VGND_c_894_n 0.0129947f $X=2.06 $Y=1.185 $X2=0 $Y2=0
cc_174 N_A_c_117_n N_VGND_c_898_n 0.0115976f $X=0.77 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A_c_119_n N_VGND_c_898_n 0.00824727f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_176 N_A_c_121_n N_VGND_c_898_n 0.00824727f $X=1.63 $Y=1.185 $X2=0 $Y2=0
cc_177 N_A_c_123_n N_VGND_c_898_n 0.00819843f $X=2.06 $Y=1.185 $X2=0 $Y2=0
cc_178 N_B_c_197_n N_C_c_277_n 0.0314022f $X=4.23 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_179 N_B_c_198_n C 3.4996e-19 $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_180 N_B_c_199_n C 0.0172618f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_181 N_B_c_198_n N_C_c_286_n 0.0267093f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_182 N_B_c_199_n N_C_c_286_n 0.00135597f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_183 N_B_c_200_n N_A_72_367#_c_471_n 0.0123048f $X=2.42 $Y=1.725 $X2=0 $Y2=0
cc_184 N_B_c_201_n N_A_72_367#_c_471_n 0.0105303f $X=2.85 $Y=1.725 $X2=0 $Y2=0
cc_185 N_B_c_200_n N_A_72_367#_c_473_n 6.29579e-19 $X=2.42 $Y=1.725 $X2=0 $Y2=0
cc_186 N_B_c_201_n N_A_72_367#_c_473_n 0.0101309f $X=2.85 $Y=1.725 $X2=0 $Y2=0
cc_187 N_B_c_202_n N_A_72_367#_c_473_n 0.0101309f $X=3.28 $Y=1.725 $X2=0 $Y2=0
cc_188 N_B_c_203_n N_A_72_367#_c_473_n 6.29579e-19 $X=3.71 $Y=1.725 $X2=0 $Y2=0
cc_189 N_B_c_198_n N_A_72_367#_c_473_n 5.48305e-19 $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_190 N_B_c_202_n N_A_72_367#_c_478_n 0.0105769f $X=3.28 $Y=1.725 $X2=0 $Y2=0
cc_191 N_B_c_203_n N_A_72_367#_c_478_n 0.0123048f $X=3.71 $Y=1.725 $X2=0 $Y2=0
cc_192 N_B_c_201_n N_A_72_367#_c_480_n 6.00691e-19 $X=2.85 $Y=1.725 $X2=0 $Y2=0
cc_193 N_B_c_202_n N_A_72_367#_c_480_n 6.00691e-19 $X=3.28 $Y=1.725 $X2=0 $Y2=0
cc_194 N_B_c_200_n N_VPWR_c_520_n 0.0011194f $X=2.42 $Y=1.725 $X2=0 $Y2=0
cc_195 N_B_c_200_n N_VPWR_c_523_n 0.00359964f $X=2.42 $Y=1.725 $X2=0 $Y2=0
cc_196 N_B_c_201_n N_VPWR_c_523_n 0.0035993f $X=2.85 $Y=1.725 $X2=0 $Y2=0
cc_197 N_B_c_202_n N_VPWR_c_523_n 0.0035993f $X=3.28 $Y=1.725 $X2=0 $Y2=0
cc_198 N_B_c_203_n N_VPWR_c_523_n 0.00359964f $X=3.71 $Y=1.725 $X2=0 $Y2=0
cc_199 N_B_c_200_n N_VPWR_c_517_n 0.00537821f $X=2.42 $Y=1.725 $X2=0 $Y2=0
cc_200 N_B_c_201_n N_VPWR_c_517_n 0.00535284f $X=2.85 $Y=1.725 $X2=0 $Y2=0
cc_201 N_B_c_202_n N_VPWR_c_517_n 0.00535284f $X=3.28 $Y=1.725 $X2=0 $Y2=0
cc_202 N_B_c_203_n N_VPWR_c_517_n 0.00665257f $X=3.71 $Y=1.725 $X2=0 $Y2=0
cc_203 N_B_c_201_n N_A_499_367#_c_622_n 0.0107712f $X=2.85 $Y=1.725 $X2=0 $Y2=0
cc_204 N_B_c_202_n N_A_499_367#_c_622_n 0.0109695f $X=3.28 $Y=1.725 $X2=0 $Y2=0
cc_205 N_B_c_198_n N_A_499_367#_c_622_n 0.0120729f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_206 N_B_c_199_n N_A_499_367#_c_622_n 0.0477199f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_207 N_B_c_200_n N_A_499_367#_c_617_n 0.00311996f $X=2.42 $Y=1.725 $X2=0 $Y2=0
cc_208 N_B_c_198_n N_A_499_367#_c_617_n 0.00628811f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_209 N_B_c_199_n N_A_499_367#_c_617_n 0.0171434f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_210 N_B_c_203_n N_A_499_367#_c_618_n 0.0135323f $X=3.71 $Y=1.725 $X2=0 $Y2=0
cc_211 N_B_c_198_n N_A_499_367#_c_618_n 0.0188264f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_212 N_B_c_199_n N_A_499_367#_c_618_n 0.0563797f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_213 N_B_c_198_n N_A_499_367#_c_632_n 0.00603335f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_214 N_B_c_199_n N_A_499_367#_c_632_n 0.0171434f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_215 N_B_c_194_n N_Y_c_763_n 0.0153277f $X=2.94 $Y=1.185 $X2=0 $Y2=0
cc_216 N_B_c_198_n N_Y_c_763_n 0.0138217f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_217 N_B_c_199_n N_Y_c_763_n 0.048476f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_218 N_B_c_195_n N_Y_c_771_n 0.013164f $X=3.37 $Y=1.185 $X2=0 $Y2=0
cc_219 N_B_c_196_n N_Y_c_771_n 0.013164f $X=3.8 $Y=1.185 $X2=0 $Y2=0
cc_220 N_B_c_198_n N_Y_c_771_n 0.00269787f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_221 N_B_c_199_n N_Y_c_771_n 0.0412767f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_222 N_B_c_197_n N_Y_c_775_n 0.0131174f $X=4.23 $Y=1.185 $X2=0 $Y2=0
cc_223 N_B_c_198_n N_Y_c_775_n 0.00154121f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_224 N_B_c_199_n N_Y_c_775_n 0.0154758f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_225 N_B_c_198_n N_Y_c_778_n 0.00279027f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_226 N_B_c_199_n N_Y_c_778_n 0.0147846f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_227 N_B_c_198_n N_Y_c_780_n 0.00248163f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_228 N_B_c_199_n N_Y_c_780_n 0.0145966f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_229 N_B_c_194_n N_VGND_c_874_n 5.8251e-19 $X=2.94 $Y=1.185 $X2=0 $Y2=0
cc_230 N_B_c_195_n N_VGND_c_874_n 0.0101643f $X=3.37 $Y=1.185 $X2=0 $Y2=0
cc_231 N_B_c_196_n N_VGND_c_874_n 0.0101622f $X=3.8 $Y=1.185 $X2=0 $Y2=0
cc_232 N_B_c_197_n N_VGND_c_874_n 5.80819e-19 $X=4.23 $Y=1.185 $X2=0 $Y2=0
cc_233 N_B_c_196_n N_VGND_c_875_n 5.80819e-19 $X=3.8 $Y=1.185 $X2=0 $Y2=0
cc_234 N_B_c_197_n N_VGND_c_875_n 0.0100971f $X=4.23 $Y=1.185 $X2=0 $Y2=0
cc_235 N_B_c_196_n N_VGND_c_886_n 0.00486043f $X=3.8 $Y=1.185 $X2=0 $Y2=0
cc_236 N_B_c_197_n N_VGND_c_886_n 0.00486043f $X=4.23 $Y=1.185 $X2=0 $Y2=0
cc_237 N_B_c_194_n N_VGND_c_890_n 0.00505556f $X=2.94 $Y=1.185 $X2=0 $Y2=0
cc_238 N_B_c_195_n N_VGND_c_890_n 0.00486043f $X=3.37 $Y=1.185 $X2=0 $Y2=0
cc_239 N_B_c_194_n N_VGND_c_894_n 0.0127123f $X=2.94 $Y=1.185 $X2=0 $Y2=0
cc_240 N_B_c_195_n N_VGND_c_894_n 5.9197e-19 $X=3.37 $Y=1.185 $X2=0 $Y2=0
cc_241 N_B_c_194_n N_VGND_c_898_n 0.00850734f $X=2.94 $Y=1.185 $X2=0 $Y2=0
cc_242 N_B_c_195_n N_VGND_c_898_n 0.00824727f $X=3.37 $Y=1.185 $X2=0 $Y2=0
cc_243 N_B_c_196_n N_VGND_c_898_n 0.00824727f $X=3.8 $Y=1.185 $X2=0 $Y2=0
cc_244 N_B_c_197_n N_VGND_c_898_n 0.00824727f $X=4.23 $Y=1.185 $X2=0 $Y2=0
cc_245 N_C_c_283_n N_D_M1013_g 0.0245111f $X=5.95 $Y=1.185 $X2=0 $Y2=0
cc_246 C N_D_M1013_g 0.00133638f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_247 N_C_M1025_g N_D_M1000_g 0.0245111f $X=5.95 $Y=2.465 $X2=0 $Y2=0
cc_248 C N_D_c_374_n 2.72706e-19 $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_249 N_C_c_286_n N_D_c_374_n 0.0245111f $X=5.95 $Y=1.35 $X2=0 $Y2=0
cc_250 C N_D_c_375_n 0.0229335f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_251 N_C_c_286_n N_D_c_375_n 3.55129e-19 $X=5.95 $Y=1.35 $X2=0 $Y2=0
cc_252 N_C_M1003_g N_A_72_367#_c_457_n 0.00129321f $X=4.66 $Y=2.465 $X2=0 $Y2=0
cc_253 N_C_M1003_g N_VPWR_c_523_n 0.00357842f $X=4.66 $Y=2.465 $X2=0 $Y2=0
cc_254 N_C_M1010_g N_VPWR_c_523_n 0.00357842f $X=5.09 $Y=2.465 $X2=0 $Y2=0
cc_255 N_C_M1017_g N_VPWR_c_523_n 0.00357842f $X=5.52 $Y=2.465 $X2=0 $Y2=0
cc_256 N_C_M1025_g N_VPWR_c_523_n 0.00357842f $X=5.95 $Y=2.465 $X2=0 $Y2=0
cc_257 N_C_M1003_g N_VPWR_c_517_n 0.00665087f $X=4.66 $Y=2.465 $X2=0 $Y2=0
cc_258 N_C_M1010_g N_VPWR_c_517_n 0.00535118f $X=5.09 $Y=2.465 $X2=0 $Y2=0
cc_259 N_C_M1017_g N_VPWR_c_517_n 0.00535118f $X=5.52 $Y=2.465 $X2=0 $Y2=0
cc_260 N_C_M1025_g N_VPWR_c_517_n 0.00537652f $X=5.95 $Y=2.465 $X2=0 $Y2=0
cc_261 N_C_M1003_g N_A_499_367#_c_618_n 0.0172219f $X=4.66 $Y=2.465 $X2=0 $Y2=0
cc_262 C N_A_499_367#_c_618_n 0.00780537f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_263 N_C_M1010_g N_A_499_367#_c_619_n 0.0137774f $X=5.09 $Y=2.465 $X2=0 $Y2=0
cc_264 N_C_M1017_g N_A_499_367#_c_619_n 0.0134566f $X=5.52 $Y=2.465 $X2=0 $Y2=0
cc_265 N_C_M1025_g N_A_499_367#_c_619_n 0.00215072f $X=5.95 $Y=2.465 $X2=0 $Y2=0
cc_266 C N_A_499_367#_c_619_n 0.0665248f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_267 N_C_c_286_n N_A_499_367#_c_619_n 0.00141664f $X=5.95 $Y=1.35 $X2=0 $Y2=0
cc_268 C N_A_499_367#_c_620_n 0.0167876f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_269 N_C_c_286_n N_A_499_367#_c_620_n 7.50045e-19 $X=5.95 $Y=1.35 $X2=0 $Y2=0
cc_270 N_C_M1003_g N_A_864_367#_c_665_n 5.81207e-19 $X=4.66 $Y=2.465 $X2=0 $Y2=0
cc_271 N_C_M1003_g N_A_864_367#_c_666_n 0.0102648f $X=4.66 $Y=2.465 $X2=0 $Y2=0
cc_272 N_C_M1010_g N_A_864_367#_c_666_n 6.27227e-19 $X=5.09 $Y=2.465 $X2=0 $Y2=0
cc_273 N_C_M1003_g N_A_864_367#_c_672_n 0.0105205f $X=4.66 $Y=2.465 $X2=0 $Y2=0
cc_274 N_C_M1010_g N_A_864_367#_c_672_n 0.0105205f $X=5.09 $Y=2.465 $X2=0 $Y2=0
cc_275 N_C_M1003_g N_A_864_367#_c_674_n 6.27227e-19 $X=4.66 $Y=2.465 $X2=0 $Y2=0
cc_276 N_C_M1010_g N_A_864_367#_c_674_n 0.0102236f $X=5.09 $Y=2.465 $X2=0 $Y2=0
cc_277 N_C_M1017_g N_A_864_367#_c_674_n 0.0102236f $X=5.52 $Y=2.465 $X2=0 $Y2=0
cc_278 N_C_M1025_g N_A_864_367#_c_674_n 6.27227e-19 $X=5.95 $Y=2.465 $X2=0 $Y2=0
cc_279 N_C_M1017_g N_A_864_367#_c_678_n 0.0105205f $X=5.52 $Y=2.465 $X2=0 $Y2=0
cc_280 N_C_M1025_g N_A_864_367#_c_678_n 0.0105205f $X=5.95 $Y=2.465 $X2=0 $Y2=0
cc_281 N_C_M1017_g N_A_864_367#_c_680_n 6.37774e-19 $X=5.52 $Y=2.465 $X2=0 $Y2=0
cc_282 N_C_M1025_g N_A_864_367#_c_680_n 0.0106544f $X=5.95 $Y=2.465 $X2=0 $Y2=0
cc_283 C N_A_864_367#_c_680_n 0.00195743f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_284 N_C_M1010_g N_A_864_367#_c_683_n 5.81207e-19 $X=5.09 $Y=2.465 $X2=0 $Y2=0
cc_285 N_C_M1017_g N_A_864_367#_c_683_n 5.81207e-19 $X=5.52 $Y=2.465 $X2=0 $Y2=0
cc_286 N_C_M1025_g N_A_864_367#_c_685_n 5.81207e-19 $X=5.95 $Y=2.465 $X2=0 $Y2=0
cc_287 N_C_c_277_n N_Y_c_775_n 0.0144748f $X=4.66 $Y=1.185 $X2=0 $Y2=0
cc_288 C N_Y_c_775_n 0.00596406f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_289 N_C_c_279_n N_Y_c_784_n 0.013164f $X=5.09 $Y=1.185 $X2=0 $Y2=0
cc_290 N_C_c_281_n N_Y_c_784_n 0.013164f $X=5.52 $Y=1.185 $X2=0 $Y2=0
cc_291 C N_Y_c_784_n 0.0412767f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_292 N_C_c_286_n N_Y_c_784_n 0.00230884f $X=5.95 $Y=1.35 $X2=0 $Y2=0
cc_293 N_C_c_283_n N_Y_c_788_n 0.0131174f $X=5.95 $Y=1.185 $X2=0 $Y2=0
cc_294 C N_Y_c_788_n 0.0149846f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_295 C N_Y_c_790_n 0.0145966f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_296 N_C_c_286_n N_Y_c_790_n 0.00240082f $X=5.95 $Y=1.35 $X2=0 $Y2=0
cc_297 C N_Y_c_792_n 0.0145966f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_298 N_C_c_286_n N_Y_c_792_n 0.00240082f $X=5.95 $Y=1.35 $X2=0 $Y2=0
cc_299 N_C_c_277_n N_VGND_c_875_n 0.0100971f $X=4.66 $Y=1.185 $X2=0 $Y2=0
cc_300 N_C_c_279_n N_VGND_c_875_n 5.80819e-19 $X=5.09 $Y=1.185 $X2=0 $Y2=0
cc_301 N_C_c_277_n N_VGND_c_876_n 5.80819e-19 $X=4.66 $Y=1.185 $X2=0 $Y2=0
cc_302 N_C_c_279_n N_VGND_c_876_n 0.0101622f $X=5.09 $Y=1.185 $X2=0 $Y2=0
cc_303 N_C_c_281_n N_VGND_c_876_n 0.0101622f $X=5.52 $Y=1.185 $X2=0 $Y2=0
cc_304 N_C_c_283_n N_VGND_c_876_n 5.80819e-19 $X=5.95 $Y=1.185 $X2=0 $Y2=0
cc_305 N_C_c_281_n N_VGND_c_877_n 0.00486043f $X=5.52 $Y=1.185 $X2=0 $Y2=0
cc_306 N_C_c_283_n N_VGND_c_877_n 0.00486043f $X=5.95 $Y=1.185 $X2=0 $Y2=0
cc_307 N_C_c_281_n N_VGND_c_878_n 5.80819e-19 $X=5.52 $Y=1.185 $X2=0 $Y2=0
cc_308 N_C_c_283_n N_VGND_c_878_n 0.0100971f $X=5.95 $Y=1.185 $X2=0 $Y2=0
cc_309 N_C_c_277_n N_VGND_c_888_n 0.00486043f $X=4.66 $Y=1.185 $X2=0 $Y2=0
cc_310 N_C_c_279_n N_VGND_c_888_n 0.00486043f $X=5.09 $Y=1.185 $X2=0 $Y2=0
cc_311 N_C_c_277_n N_VGND_c_898_n 0.00824727f $X=4.66 $Y=1.185 $X2=0 $Y2=0
cc_312 N_C_c_279_n N_VGND_c_898_n 0.00824727f $X=5.09 $Y=1.185 $X2=0 $Y2=0
cc_313 N_C_c_281_n N_VGND_c_898_n 0.00824727f $X=5.52 $Y=1.185 $X2=0 $Y2=0
cc_314 N_C_c_283_n N_VGND_c_898_n 0.00824727f $X=5.95 $Y=1.185 $X2=0 $Y2=0
cc_315 N_D_M1000_g N_VPWR_c_523_n 0.00357842f $X=6.38 $Y=2.465 $X2=0 $Y2=0
cc_316 N_D_M1001_g N_VPWR_c_523_n 0.00357842f $X=6.81 $Y=2.465 $X2=0 $Y2=0
cc_317 N_D_M1008_g N_VPWR_c_523_n 0.00357842f $X=7.24 $Y=2.465 $X2=0 $Y2=0
cc_318 N_D_M1021_g N_VPWR_c_523_n 0.00357842f $X=7.67 $Y=2.465 $X2=0 $Y2=0
cc_319 N_D_M1000_g N_VPWR_c_517_n 0.00537652f $X=6.38 $Y=2.465 $X2=0 $Y2=0
cc_320 N_D_M1001_g N_VPWR_c_517_n 0.00535118f $X=6.81 $Y=2.465 $X2=0 $Y2=0
cc_321 N_D_M1008_g N_VPWR_c_517_n 0.00535118f $X=7.24 $Y=2.465 $X2=0 $Y2=0
cc_322 N_D_M1021_g N_VPWR_c_517_n 0.00629769f $X=7.67 $Y=2.465 $X2=0 $Y2=0
cc_323 N_D_M1000_g N_A_864_367#_c_680_n 0.0105046f $X=6.38 $Y=2.465 $X2=0 $Y2=0
cc_324 N_D_M1001_g N_A_864_367#_c_680_n 6.27227e-19 $X=6.81 $Y=2.465 $X2=0 $Y2=0
cc_325 N_D_c_375_n N_A_864_367#_c_680_n 7.33789e-19 $X=6.988 $Y=1.367 $X2=0
+ $Y2=0
cc_326 N_D_M1000_g N_A_864_367#_c_689_n 0.0105205f $X=6.38 $Y=2.465 $X2=0 $Y2=0
cc_327 N_D_M1001_g N_A_864_367#_c_689_n 0.0105205f $X=6.81 $Y=2.465 $X2=0 $Y2=0
cc_328 N_D_M1000_g N_A_864_367#_c_691_n 6.27227e-19 $X=6.38 $Y=2.465 $X2=0 $Y2=0
cc_329 N_D_M1001_g N_A_864_367#_c_691_n 0.0102236f $X=6.81 $Y=2.465 $X2=0 $Y2=0
cc_330 N_D_M1008_g N_A_864_367#_c_691_n 0.0102236f $X=7.24 $Y=2.465 $X2=0 $Y2=0
cc_331 N_D_M1021_g N_A_864_367#_c_691_n 6.27227e-19 $X=7.67 $Y=2.465 $X2=0 $Y2=0
cc_332 N_D_M1008_g N_A_864_367#_c_695_n 0.0105205f $X=7.24 $Y=2.465 $X2=0 $Y2=0
cc_333 N_D_M1021_g N_A_864_367#_c_695_n 0.0105205f $X=7.67 $Y=2.465 $X2=0 $Y2=0
cc_334 N_D_M1021_g N_A_864_367#_c_667_n 5.81207e-19 $X=7.67 $Y=2.465 $X2=0 $Y2=0
cc_335 N_D_M1008_g N_A_864_367#_c_668_n 6.27227e-19 $X=7.24 $Y=2.465 $X2=0 $Y2=0
cc_336 N_D_M1021_g N_A_864_367#_c_668_n 0.0102648f $X=7.67 $Y=2.465 $X2=0 $Y2=0
cc_337 N_D_M1000_g N_A_864_367#_c_685_n 5.81207e-19 $X=6.38 $Y=2.465 $X2=0 $Y2=0
cc_338 N_D_M1001_g N_A_864_367#_c_701_n 5.81207e-19 $X=6.81 $Y=2.465 $X2=0 $Y2=0
cc_339 N_D_M1008_g N_A_864_367#_c_701_n 5.81207e-19 $X=7.24 $Y=2.465 $X2=0 $Y2=0
cc_340 N_D_M1013_g N_Y_c_788_n 0.0123951f $X=6.38 $Y=0.655 $X2=0 $Y2=0
cc_341 N_D_c_375_n N_Y_c_788_n 0.0125324f $X=6.988 $Y=1.367 $X2=0 $Y2=0
cc_342 N_D_M1016_g N_Y_c_747_n 0.0124417f $X=6.81 $Y=0.655 $X2=0 $Y2=0
cc_343 N_D_M1027_g N_Y_c_747_n 0.0160392f $X=7.24 $Y=0.655 $X2=0 $Y2=0
cc_344 N_D_M1029_g N_Y_c_747_n 2.39666e-19 $X=7.67 $Y=0.655 $X2=0 $Y2=0
cc_345 N_D_c_418_p N_Y_c_747_n 0.0251555f $X=7.49 $Y=1.44 $X2=0 $Y2=0
cc_346 N_D_c_374_n N_Y_c_747_n 0.00317504f $X=7.67 $Y=1.44 $X2=0 $Y2=0
cc_347 N_D_c_375_n N_Y_c_747_n 0.0292687f $X=6.988 $Y=1.367 $X2=0 $Y2=0
cc_348 N_D_M1001_g N_Y_c_751_n 0.0138775f $X=6.81 $Y=2.465 $X2=0 $Y2=0
cc_349 N_D_M1008_g N_Y_c_751_n 0.0141975f $X=7.24 $Y=2.465 $X2=0 $Y2=0
cc_350 N_D_c_374_n N_Y_c_751_n 0.00246815f $X=7.67 $Y=1.44 $X2=0 $Y2=0
cc_351 N_D_c_375_n N_Y_c_751_n 0.0483976f $X=6.988 $Y=1.367 $X2=0 $Y2=0
cc_352 N_D_M1000_g N_Y_c_752_n 0.00251344f $X=6.38 $Y=2.465 $X2=0 $Y2=0
cc_353 N_D_c_374_n N_Y_c_752_n 0.00256759f $X=7.67 $Y=1.44 $X2=0 $Y2=0
cc_354 N_D_c_375_n N_Y_c_752_n 0.0159733f $X=6.988 $Y=1.367 $X2=0 $Y2=0
cc_355 N_D_M1029_g N_Y_c_748_n 0.0155321f $X=7.67 $Y=0.655 $X2=0 $Y2=0
cc_356 N_D_c_418_p N_Y_c_748_n 0.00731891f $X=7.49 $Y=1.44 $X2=0 $Y2=0
cc_357 N_D_M1021_g N_Y_c_753_n 0.0167171f $X=7.67 $Y=2.465 $X2=0 $Y2=0
cc_358 N_D_c_418_p N_Y_c_753_n 0.00728094f $X=7.49 $Y=1.44 $X2=0 $Y2=0
cc_359 N_D_c_374_n N_Y_c_813_n 6.68767e-19 $X=7.67 $Y=1.44 $X2=0 $Y2=0
cc_360 N_D_c_375_n N_Y_c_813_n 0.0153383f $X=6.988 $Y=1.367 $X2=0 $Y2=0
cc_361 N_D_c_418_p N_Y_c_754_n 0.0153308f $X=7.49 $Y=1.44 $X2=0 $Y2=0
cc_362 N_D_c_374_n N_Y_c_754_n 0.00256759f $X=7.67 $Y=1.44 $X2=0 $Y2=0
cc_363 N_D_M1029_g Y 0.0196656f $X=7.67 $Y=0.655 $X2=0 $Y2=0
cc_364 N_D_c_418_p Y 0.0137867f $X=7.49 $Y=1.44 $X2=0 $Y2=0
cc_365 N_D_M1013_g N_VGND_c_878_n 0.0100971f $X=6.38 $Y=0.655 $X2=0 $Y2=0
cc_366 N_D_M1016_g N_VGND_c_878_n 5.80819e-19 $X=6.81 $Y=0.655 $X2=0 $Y2=0
cc_367 N_D_M1013_g N_VGND_c_879_n 5.80819e-19 $X=6.38 $Y=0.655 $X2=0 $Y2=0
cc_368 N_D_M1016_g N_VGND_c_879_n 0.0101622f $X=6.81 $Y=0.655 $X2=0 $Y2=0
cc_369 N_D_M1027_g N_VGND_c_879_n 0.0100888f $X=7.24 $Y=0.655 $X2=0 $Y2=0
cc_370 N_D_M1029_g N_VGND_c_879_n 5.75816e-19 $X=7.67 $Y=0.655 $X2=0 $Y2=0
cc_371 N_D_M1027_g N_VGND_c_881_n 6.14008e-19 $X=7.24 $Y=0.655 $X2=0 $Y2=0
cc_372 N_D_M1029_g N_VGND_c_881_n 0.0112405f $X=7.67 $Y=0.655 $X2=0 $Y2=0
cc_373 N_D_M1013_g N_VGND_c_891_n 0.00486043f $X=6.38 $Y=0.655 $X2=0 $Y2=0
cc_374 N_D_M1016_g N_VGND_c_891_n 0.00486043f $X=6.81 $Y=0.655 $X2=0 $Y2=0
cc_375 N_D_M1027_g N_VGND_c_892_n 0.00486043f $X=7.24 $Y=0.655 $X2=0 $Y2=0
cc_376 N_D_M1029_g N_VGND_c_892_n 0.00486043f $X=7.67 $Y=0.655 $X2=0 $Y2=0
cc_377 N_D_M1013_g N_VGND_c_898_n 0.00824727f $X=6.38 $Y=0.655 $X2=0 $Y2=0
cc_378 N_D_M1016_g N_VGND_c_898_n 0.00824727f $X=6.81 $Y=0.655 $X2=0 $Y2=0
cc_379 N_D_M1027_g N_VGND_c_898_n 0.00824727f $X=7.24 $Y=0.655 $X2=0 $Y2=0
cc_380 N_D_M1029_g N_VGND_c_898_n 0.00824727f $X=7.67 $Y=0.655 $X2=0 $Y2=0
cc_381 N_A_72_367#_c_460_n N_VPWR_M1002_s 0.00334576f $X=1.25 $Y=2.005 $X2=-0.19
+ $Y2=1.655
cc_382 N_A_72_367#_c_464_n N_VPWR_M1014_s 0.00334576f $X=2.11 $Y=2.005 $X2=0
+ $Y2=0
cc_383 N_A_72_367#_c_460_n N_VPWR_c_518_n 0.0170777f $X=1.25 $Y=2.005 $X2=0
+ $Y2=0
cc_384 N_A_72_367#_c_486_p N_VPWR_c_519_n 0.0117038f $X=1.345 $Y=2.9 $X2=0 $Y2=0
cc_385 N_A_72_367#_c_464_n N_VPWR_c_520_n 0.0170777f $X=2.11 $Y=2.005 $X2=0
+ $Y2=0
cc_386 N_A_72_367#_c_455_n N_VPWR_c_521_n 0.0167395f $X=0.485 $Y=2.9 $X2=0 $Y2=0
cc_387 N_A_72_367#_c_489_p N_VPWR_c_523_n 0.0132784f $X=2.227 $Y=2.895 $X2=0
+ $Y2=0
cc_388 N_A_72_367#_c_471_n N_VPWR_c_523_n 0.0295311f $X=2.9 $Y=2.98 $X2=0 $Y2=0
cc_389 N_A_72_367#_c_478_n N_VPWR_c_523_n 0.0295311f $X=3.785 $Y=2.98 $X2=0
+ $Y2=0
cc_390 N_A_72_367#_c_456_n N_VPWR_c_523_n 0.018348f $X=3.937 $Y=2.895 $X2=0
+ $Y2=0
cc_391 N_A_72_367#_c_480_n N_VPWR_c_523_n 0.0179231f $X=3.065 $Y=2.9 $X2=0 $Y2=0
cc_392 N_A_72_367#_M1002_d N_VPWR_c_517_n 0.00371907f $X=0.36 $Y=1.835 $X2=0
+ $Y2=0
cc_393 N_A_72_367#_M1006_d N_VPWR_c_517_n 0.00536823f $X=1.205 $Y=1.835 $X2=0
+ $Y2=0
cc_394 N_A_72_367#_M1019_d N_VPWR_c_517_n 0.00376843f $X=2.065 $Y=1.835 $X2=0
+ $Y2=0
cc_395 N_A_72_367#_M1020_d N_VPWR_c_517_n 0.00223819f $X=2.925 $Y=1.835 $X2=0
+ $Y2=0
cc_396 N_A_72_367#_M1031_d N_VPWR_c_517_n 0.00215406f $X=3.785 $Y=1.835 $X2=0
+ $Y2=0
cc_397 N_A_72_367#_c_455_n N_VPWR_c_517_n 0.00998284f $X=0.485 $Y=2.9 $X2=0
+ $Y2=0
cc_398 N_A_72_367#_c_486_p N_VPWR_c_517_n 0.00727431f $X=1.345 $Y=2.9 $X2=0
+ $Y2=0
cc_399 N_A_72_367#_c_489_p N_VPWR_c_517_n 0.0090542f $X=2.227 $Y=2.895 $X2=0
+ $Y2=0
cc_400 N_A_72_367#_c_471_n N_VPWR_c_517_n 0.0194467f $X=2.9 $Y=2.98 $X2=0 $Y2=0
cc_401 N_A_72_367#_c_478_n N_VPWR_c_517_n 0.0194467f $X=3.785 $Y=2.98 $X2=0
+ $Y2=0
cc_402 N_A_72_367#_c_456_n N_VPWR_c_517_n 0.0117627f $X=3.937 $Y=2.895 $X2=0
+ $Y2=0
cc_403 N_A_72_367#_c_480_n N_VPWR_c_517_n 0.0123929f $X=3.065 $Y=2.9 $X2=0 $Y2=0
cc_404 N_A_72_367#_c_471_n N_A_499_367#_M1009_s 0.00335807f $X=2.9 $Y=2.98
+ $X2=-0.19 $Y2=1.655
cc_405 N_A_72_367#_c_478_n N_A_499_367#_M1022_s 0.00335807f $X=3.785 $Y=2.98
+ $X2=0 $Y2=0
cc_406 N_A_72_367#_c_471_n N_A_499_367#_c_645_n 0.012662f $X=2.9 $Y=2.98 $X2=0
+ $Y2=0
cc_407 N_A_72_367#_M1020_d N_A_499_367#_c_622_n 0.00180746f $X=2.925 $Y=1.835
+ $X2=0 $Y2=0
cc_408 N_A_72_367#_c_473_n N_A_499_367#_c_622_n 0.0163514f $X=3.065 $Y=2.22
+ $X2=0 $Y2=0
cc_409 N_A_72_367#_c_478_n N_A_499_367#_c_648_n 0.012662f $X=3.785 $Y=2.98 $X2=0
+ $Y2=0
cc_410 N_A_72_367#_M1031_d N_A_499_367#_c_618_n 0.00244825f $X=3.785 $Y=1.835
+ $X2=0 $Y2=0
cc_411 N_A_72_367#_c_457_n N_A_499_367#_c_618_n 0.0193774f $X=3.925 $Y=2.22
+ $X2=0 $Y2=0
cc_412 N_A_72_367#_c_456_n N_A_864_367#_c_665_n 0.0138501f $X=3.937 $Y=2.895
+ $X2=0 $Y2=0
cc_413 N_A_72_367#_c_456_n N_A_864_367#_c_666_n 7.79003e-19 $X=3.937 $Y=2.895
+ $X2=0 $Y2=0
cc_414 N_A_72_367#_c_457_n N_A_864_367#_c_666_n 0.0642607f $X=3.925 $Y=2.22
+ $X2=0 $Y2=0
cc_415 N_VPWR_c_517_n N_A_499_367#_M1009_s 0.00225465f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_416 N_VPWR_c_517_n N_A_499_367#_M1022_s 0.00225465f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_517_n N_A_499_367#_M1003_d 0.00225186f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_517_n N_A_499_367#_M1017_d 0.00225186f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_517_n N_A_864_367#_M1003_s 0.00215158f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_420 N_VPWR_c_517_n N_A_864_367#_M1010_s 0.00223559f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_517_n N_A_864_367#_M1025_s 0.00223559f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_517_n N_A_864_367#_M1001_s 0.00223559f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_517_n N_A_864_367#_M1021_s 0.00215158f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_523_n N_A_864_367#_c_665_n 0.0211538f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_517_n N_A_864_367#_c_665_n 0.0126374f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_523_n N_A_864_367#_c_672_n 0.0298674f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_517_n N_A_864_367#_c_672_n 0.0187823f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_523_n N_A_864_367#_c_678_n 0.0298674f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_517_n N_A_864_367#_c_678_n 0.0187823f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_523_n N_A_864_367#_c_689_n 0.0298674f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_517_n N_A_864_367#_c_689_n 0.0187823f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_523_n N_A_864_367#_c_695_n 0.0298674f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_517_n N_A_864_367#_c_695_n 0.0187823f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_523_n N_A_864_367#_c_667_n 0.0211538f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_517_n N_A_864_367#_c_667_n 0.0126374f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_523_n N_A_864_367#_c_683_n 0.0189946f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_517_n N_A_864_367#_c_683_n 0.0124451f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_523_n N_A_864_367#_c_685_n 0.0189946f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_517_n N_A_864_367#_c_685_n 0.0124451f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_523_n N_A_864_367#_c_701_n 0.0189946f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_517_n N_A_864_367#_c_701_n 0.0124451f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_517_n N_Y_M1000_d 0.00225186f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_443 N_VPWR_c_517_n N_Y_M1008_d 0.00225186f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_444 N_A_499_367#_c_618_n N_A_864_367#_M1003_s 0.00244825f $X=4.78 $Y=1.79
+ $X2=-0.19 $Y2=1.655
cc_445 N_A_499_367#_c_619_n N_A_864_367#_M1010_s 0.00180746f $X=5.64 $Y=1.79
+ $X2=0 $Y2=0
cc_446 N_A_499_367#_c_618_n N_A_864_367#_c_666_n 0.021083f $X=4.78 $Y=1.79 $X2=0
+ $Y2=0
cc_447 N_A_499_367#_M1003_d N_A_864_367#_c_672_n 0.00332344f $X=4.735 $Y=1.835
+ $X2=0 $Y2=0
cc_448 N_A_499_367#_c_659_p N_A_864_367#_c_672_n 0.0126348f $X=4.875 $Y=1.98
+ $X2=0 $Y2=0
cc_449 N_A_499_367#_c_619_n N_A_864_367#_c_674_n 0.0163515f $X=5.64 $Y=1.79
+ $X2=0 $Y2=0
cc_450 N_A_499_367#_M1017_d N_A_864_367#_c_678_n 0.00332344f $X=5.595 $Y=1.835
+ $X2=0 $Y2=0
cc_451 N_A_499_367#_c_662_p N_A_864_367#_c_678_n 0.0126348f $X=5.735 $Y=1.98
+ $X2=0 $Y2=0
cc_452 N_A_499_367#_c_618_n N_Y_c_775_n 0.00699269f $X=4.78 $Y=1.79 $X2=0 $Y2=0
cc_453 N_A_499_367#_c_619_n N_Y_c_752_n 0.00445637f $X=5.64 $Y=1.79 $X2=0 $Y2=0
cc_454 N_A_864_367#_c_689_n N_Y_M1000_d 0.00332344f $X=6.86 $Y=2.99 $X2=0 $Y2=0
cc_455 N_A_864_367#_c_695_n N_Y_M1008_d 0.00332344f $X=7.72 $Y=2.99 $X2=0 $Y2=0
cc_456 N_A_864_367#_c_689_n N_Y_c_825_n 0.0126348f $X=6.86 $Y=2.99 $X2=0 $Y2=0
cc_457 N_A_864_367#_M1001_s N_Y_c_751_n 0.00181066f $X=6.885 $Y=1.835 $X2=0
+ $Y2=0
cc_458 N_A_864_367#_c_691_n N_Y_c_751_n 0.0164152f $X=7.025 $Y=2.14 $X2=0 $Y2=0
cc_459 N_A_864_367#_c_695_n N_Y_c_828_n 0.0126348f $X=7.72 $Y=2.99 $X2=0 $Y2=0
cc_460 N_A_864_367#_M1021_s N_Y_c_753_n 0.00252559f $X=7.745 $Y=1.835 $X2=0
+ $Y2=0
cc_461 N_A_864_367#_c_668_n N_Y_c_753_n 0.0229629f $X=7.885 $Y=2.14 $X2=0 $Y2=0
cc_462 N_Y_c_745_n N_VGND_M1011_s 0.00176461f $X=1.75 $Y=1.09 $X2=0 $Y2=0
cc_463 N_Y_c_763_n N_VGND_M1023_s 0.0195227f $X=3.055 $Y=0.955 $X2=0 $Y2=0
cc_464 N_Y_c_771_n N_VGND_M1015_d 0.00329816f $X=3.92 $Y=0.955 $X2=0 $Y2=0
cc_465 N_Y_c_775_n N_VGND_M1028_d 0.00508883f $X=4.78 $Y=0.955 $X2=0 $Y2=0
cc_466 N_Y_c_784_n N_VGND_M1018_s 0.00329816f $X=5.64 $Y=0.955 $X2=0 $Y2=0
cc_467 N_Y_c_788_n N_VGND_M1030_s 0.00798397f $X=6.5 $Y=0.955 $X2=0 $Y2=0
cc_468 N_Y_c_747_n N_VGND_M1016_d 0.003325f $X=7.315 $Y=0.955 $X2=0 $Y2=0
cc_469 N_Y_c_748_n N_VGND_M1029_d 0.00261087f $X=7.825 $Y=1.095 $X2=0 $Y2=0
cc_470 N_Y_c_746_n N_VGND_c_872_n 0.00455995f $X=1.08 $Y=1.09 $X2=0 $Y2=0
cc_471 N_Y_c_745_n N_VGND_c_873_n 0.0170777f $X=1.75 $Y=1.09 $X2=0 $Y2=0
cc_472 N_Y_c_771_n N_VGND_c_874_n 0.0170777f $X=3.92 $Y=0.955 $X2=0 $Y2=0
cc_473 N_Y_c_775_n N_VGND_c_875_n 0.0170777f $X=4.78 $Y=0.955 $X2=0 $Y2=0
cc_474 N_Y_c_784_n N_VGND_c_876_n 0.0170777f $X=5.64 $Y=0.955 $X2=0 $Y2=0
cc_475 N_Y_c_844_p N_VGND_c_877_n 0.0117038f $X=5.735 $Y=0.43 $X2=0 $Y2=0
cc_476 N_Y_c_788_n N_VGND_c_878_n 0.0170777f $X=6.5 $Y=0.955 $X2=0 $Y2=0
cc_477 N_Y_c_747_n N_VGND_c_879_n 0.0170777f $X=7.315 $Y=0.955 $X2=0 $Y2=0
cc_478 N_Y_c_748_n N_VGND_c_881_n 0.0239691f $X=7.825 $Y=1.095 $X2=0 $Y2=0
cc_479 N_Y_c_848_p N_VGND_c_884_n 0.0133395f $X=0.985 $Y=0.42 $X2=0 $Y2=0
cc_480 N_Y_c_849_p N_VGND_c_886_n 0.0117038f $X=4.015 $Y=0.43 $X2=0 $Y2=0
cc_481 N_Y_c_850_p N_VGND_c_888_n 0.0117038f $X=4.875 $Y=0.43 $X2=0 $Y2=0
cc_482 N_Y_c_851_p N_VGND_c_890_n 0.0118713f $X=3.155 $Y=0.43 $X2=0 $Y2=0
cc_483 N_Y_c_852_p N_VGND_c_891_n 0.0117038f $X=6.595 $Y=0.43 $X2=0 $Y2=0
cc_484 N_Y_c_853_p N_VGND_c_892_n 0.0124525f $X=7.455 $Y=0.42 $X2=0 $Y2=0
cc_485 N_Y_c_854_p N_VGND_c_893_n 0.0124525f $X=1.845 $Y=0.42 $X2=0 $Y2=0
cc_486 N_Y_c_763_n N_VGND_c_894_n 0.0532249f $X=3.055 $Y=0.955 $X2=0 $Y2=0
cc_487 N_Y_M1004_d N_VGND_c_898_n 0.00449678f $X=0.845 $Y=0.235 $X2=0 $Y2=0
cc_488 N_Y_M1012_d N_VGND_c_898_n 0.00536646f $X=1.705 $Y=0.235 $X2=0 $Y2=0
cc_489 N_Y_M1005_s N_VGND_c_898_n 0.00519434f $X=3.015 $Y=0.235 $X2=0 $Y2=0
cc_490 N_Y_M1026_s N_VGND_c_898_n 0.00536823f $X=3.875 $Y=0.235 $X2=0 $Y2=0
cc_491 N_Y_M1007_d N_VGND_c_898_n 0.00536823f $X=4.735 $Y=0.235 $X2=0 $Y2=0
cc_492 N_Y_M1024_d N_VGND_c_898_n 0.00536823f $X=5.595 $Y=0.235 $X2=0 $Y2=0
cc_493 N_Y_M1013_s N_VGND_c_898_n 0.00536823f $X=6.455 $Y=0.235 $X2=0 $Y2=0
cc_494 N_Y_M1027_s N_VGND_c_898_n 0.00536646f $X=7.315 $Y=0.235 $X2=0 $Y2=0
cc_495 N_Y_c_848_p N_VGND_c_898_n 0.00828095f $X=0.985 $Y=0.42 $X2=0 $Y2=0
cc_496 N_Y_c_854_p N_VGND_c_898_n 0.00730901f $X=1.845 $Y=0.42 $X2=0 $Y2=0
cc_497 N_Y_c_851_p N_VGND_c_898_n 0.00746778f $X=3.155 $Y=0.43 $X2=0 $Y2=0
cc_498 N_Y_c_849_p N_VGND_c_898_n 0.00727431f $X=4.015 $Y=0.43 $X2=0 $Y2=0
cc_499 N_Y_c_850_p N_VGND_c_898_n 0.00727431f $X=4.875 $Y=0.43 $X2=0 $Y2=0
cc_500 N_Y_c_844_p N_VGND_c_898_n 0.00727431f $X=5.735 $Y=0.43 $X2=0 $Y2=0
cc_501 N_Y_c_852_p N_VGND_c_898_n 0.00727431f $X=6.595 $Y=0.43 $X2=0 $Y2=0
cc_502 N_Y_c_853_p N_VGND_c_898_n 0.00730901f $X=7.455 $Y=0.42 $X2=0 $Y2=0
