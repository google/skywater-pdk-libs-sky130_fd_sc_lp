* File: sky130_fd_sc_lp__clkinvlp_2.pex.spice
* Created: Wed Sep  2 09:41:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKINVLP_2%A 3 5 7 8 10 13 15 17 28
r38 27 28 30.5162 $w=6.16e-07 $l=3.9e-07 $layer=POLY_cond $X=0.85 $Y=1.33
+ $X2=1.24 $Y2=1.33
r39 26 27 1.56494 $w=6.16e-07 $l=2e-08 $layer=POLY_cond $X=0.83 $Y=1.33 $X2=0.85
+ $Y2=1.33
r40 24 26 10.9545 $w=6.16e-07 $l=1.4e-07 $layer=POLY_cond $X=0.69 $Y=1.33
+ $X2=0.83 $Y2=1.33
r41 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.16 $X2=0.69 $Y2=1.16
r42 17 25 0.4571 $w=7.83e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=1.387 $X2=0.69
+ $Y2=1.387
r43 15 25 6.8565 $w=7.83e-07 $l=4.5e-07 $layer=LI1_cond $X=0.24 $Y=1.387
+ $X2=0.69 $Y2=1.387
r44 11 28 9.38961 $w=6.16e-07 $l=3.90416e-07 $layer=POLY_cond $X=1.36 $Y=1.665
+ $X2=1.24 $Y2=1.33
r45 11 13 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=1.36 $Y=1.665
+ $X2=1.36 $Y2=2.48
r46 8 28 36.7582 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.24 $Y=0.995
+ $X2=1.24 $Y2=1.33
r47 8 10 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.24 $Y=0.995
+ $X2=1.24 $Y2=0.61
r48 5 27 36.7582 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.85 $Y=0.995
+ $X2=0.85 $Y2=1.33
r49 5 7 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.85 $Y=0.995
+ $X2=0.85 $Y2=0.61
r50 1 26 23.9406 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.83 $Y=1.665
+ $X2=0.83 $Y2=1.33
r51 1 3 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=0.83 $Y=1.665 $X2=0.83
+ $Y2=2.48
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_2%VPWR 1 2 9 13 15 20 21 22 28 34
r21 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r22 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r23 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r24 28 33 4.42822 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.49 $Y=3.33
+ $X2=1.705 $Y2=3.33
r25 28 30 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.49 $Y=3.33 $X2=1.2
+ $Y2=3.33
r26 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 22 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r28 22 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 20 25 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.24
+ $Y2=3.33
r30 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.4 $Y=3.33
+ $X2=0.565 $Y2=3.33
r31 19 30 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=0.73 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=3.33
+ $X2=0.565 $Y2=3.33
r33 15 18 27.2745 $w=2.98e-07 $l=7.1e-07 $layer=LI1_cond $X=1.64 $Y=2.125
+ $X2=1.64 $Y2=2.835
r34 13 33 3.08945 $w=3e-07 $l=1.12916e-07 $layer=LI1_cond $X=1.64 $Y=3.245
+ $X2=1.705 $Y2=3.33
r35 13 18 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=1.64 $Y=3.245
+ $X2=1.64 $Y2=2.835
r36 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.565 $Y=2.125
+ $X2=0.565 $Y2=2.835
r37 7 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.565 $Y=3.245
+ $X2=0.565 $Y2=3.33
r38 7 12 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.565 $Y=3.245
+ $X2=0.565 $Y2=2.835
r39 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.98 $X2=1.625 $Y2=2.835
r40 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.98 $X2=1.625 $Y2=2.125
r41 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.44
+ $Y=1.98 $X2=0.565 $Y2=2.835
r42 1 9 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.44
+ $Y=1.98 $X2=0.565 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_2%Y 1 2 11 13 14 15 16 17 18 43
r27 43 44 3.07301 $w=3.88e-07 $l=7.5e-08 $layer=LI1_cond $X=1.125 $Y=2.035
+ $X2=1.125 $Y2=1.96
r28 34 47 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=1.125 $Y=2.155
+ $X2=1.125 $Y2=2.125
r29 18 40 1.77299 $w=3.88e-07 $l=6e-08 $layer=LI1_cond $X=1.125 $Y=2.775
+ $X2=1.125 $Y2=2.835
r30 17 18 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.125 $Y=2.405
+ $X2=1.125 $Y2=2.775
r31 17 34 7.38745 $w=3.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.125 $Y=2.405
+ $X2=1.125 $Y2=2.155
r32 16 47 2.51173 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=2.04
+ $X2=1.125 $Y2=2.125
r33 16 43 0.147749 $w=3.88e-07 $l=5e-09 $layer=LI1_cond $X=1.125 $Y=2.04
+ $X2=1.125 $Y2=2.035
r34 16 44 0.202183 $w=2.83e-07 $l=5e-09 $layer=LI1_cond $X=1.177 $Y=1.955
+ $X2=1.177 $Y2=1.96
r35 15 16 11.7266 $w=2.83e-07 $l=2.9e-07 $layer=LI1_cond $X=1.177 $Y=1.665
+ $X2=1.177 $Y2=1.955
r36 14 15 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.177 $Y=1.295
+ $X2=1.177 $Y2=1.665
r37 13 14 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.177 $Y=0.925
+ $X2=1.177 $Y2=1.295
r38 8 13 5.86331 $w=2.83e-07 $l=1.45e-07 $layer=LI1_cond $X=1.177 $Y=0.78
+ $X2=1.177 $Y2=0.925
r39 7 11 7.15075 $w=4.63e-07 $l=2.78e-07 $layer=LI1_cond $X=1.177 $Y=0.547
+ $X2=1.455 $Y2=0.547
r40 7 8 3.61438 $w=2.85e-07 $l=2.33e-07 $layer=LI1_cond $X=1.177 $Y=0.547
+ $X2=1.177 $Y2=0.78
r41 2 47 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.955
+ $Y=1.98 $X2=1.095 $Y2=2.125
r42 2 40 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.955
+ $Y=1.98 $X2=1.095 $Y2=2.835
r43 1 11 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.315
+ $Y=0.335 $X2=1.455 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_2%VGND 1 6 8 10 17 18 21
r16 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r17 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r18 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.8 $Y=0 $X2=0.635
+ $Y2=0
r19 15 17 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.8 $Y=0 $X2=1.68
+ $Y2=0
r20 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r21 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r22 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.635
+ $Y2=0
r23 10 12 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.24
+ $Y2=0
r24 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r25 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r26 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.635 $Y=0.085
+ $X2=0.635 $Y2=0
r27 4 6 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.635 $Y=0.085
+ $X2=0.635 $Y2=0.61
r28 1 6 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.49
+ $Y=0.335 $X2=0.635 $Y2=0.61
.ends

