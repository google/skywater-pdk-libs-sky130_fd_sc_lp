* File: sky130_fd_sc_lp__and4bb_2.pxi.spice
* Created: Fri Aug 28 10:09:20 2020
* 
x_PM_SKY130_FD_SC_LP__AND4BB_2%A_N N_A_N_M1013_g N_A_N_c_100_n N_A_N_M1009_g A_N
+ N_A_N_c_101_n PM_SKY130_FD_SC_LP__AND4BB_2%A_N
x_PM_SKY130_FD_SC_LP__AND4BB_2%A_185_23# N_A_185_23#_M1015_s N_A_185_23#_M1008_d
+ N_A_185_23#_M1002_d N_A_185_23#_M1006_g N_A_185_23#_M1003_g
+ N_A_185_23#_c_125_n N_A_185_23#_M1010_g N_A_185_23#_c_127_n
+ N_A_185_23#_M1012_g N_A_185_23#_c_129_n N_A_185_23#_c_130_n
+ N_A_185_23#_c_217_p N_A_185_23#_c_136_n N_A_185_23#_c_188_p
+ N_A_185_23#_c_131_n N_A_185_23#_c_132_n N_A_185_23#_c_137_n
+ N_A_185_23#_c_133_n PM_SKY130_FD_SC_LP__AND4BB_2%A_185_23#
x_PM_SKY130_FD_SC_LP__AND4BB_2%A_27_133# N_A_27_133#_M1013_s N_A_27_133#_M1009_s
+ N_A_27_133#_M1015_g N_A_27_133#_M1008_g N_A_27_133#_c_234_n
+ N_A_27_133#_c_235_n N_A_27_133#_c_236_n N_A_27_133#_c_244_n
+ N_A_27_133#_c_237_n N_A_27_133#_c_238_n N_A_27_133#_c_239_n
+ N_A_27_133#_c_276_n N_A_27_133#_c_278_n N_A_27_133#_c_246_n
+ N_A_27_133#_c_247_n N_A_27_133#_c_240_n N_A_27_133#_c_290_n
+ PM_SKY130_FD_SC_LP__AND4BB_2%A_27_133#
x_PM_SKY130_FD_SC_LP__AND4BB_2%A_558_99# N_A_558_99#_M1005_d N_A_558_99#_M1007_d
+ N_A_558_99#_M1011_g N_A_558_99#_M1004_g N_A_558_99#_c_335_n
+ N_A_558_99#_c_336_n N_A_558_99#_c_344_n N_A_558_99#_c_357_n
+ N_A_558_99#_c_337_n N_A_558_99#_c_338_n N_A_558_99#_c_339_n
+ N_A_558_99#_c_340_n N_A_558_99#_c_347_n N_A_558_99#_c_341_n
+ PM_SKY130_FD_SC_LP__AND4BB_2%A_558_99#
x_PM_SKY130_FD_SC_LP__AND4BB_2%C N_C_M1001_g N_C_M1002_g C N_C_c_413_n
+ PM_SKY130_FD_SC_LP__AND4BB_2%C
x_PM_SKY130_FD_SC_LP__AND4BB_2%D N_D_M1014_g N_D_M1000_g D D N_D_c_445_n
+ N_D_c_446_n PM_SKY130_FD_SC_LP__AND4BB_2%D
x_PM_SKY130_FD_SC_LP__AND4BB_2%B_N N_B_N_M1005_g N_B_N_M1007_g N_B_N_c_484_n
+ N_B_N_c_485_n N_B_N_c_490_n B_N B_N N_B_N_c_487_n
+ PM_SKY130_FD_SC_LP__AND4BB_2%B_N
x_PM_SKY130_FD_SC_LP__AND4BB_2%VPWR N_VPWR_M1009_d N_VPWR_M1012_s N_VPWR_M1004_d
+ N_VPWR_M1000_d N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n
+ N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n VPWR N_VPWR_c_535_n
+ N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_527_n N_VPWR_c_539_n N_VPWR_c_540_n
+ N_VPWR_c_541_n PM_SKY130_FD_SC_LP__AND4BB_2%VPWR
x_PM_SKY130_FD_SC_LP__AND4BB_2%X N_X_M1006_d N_X_M1003_d N_X_c_603_n X X
+ N_X_c_601_n PM_SKY130_FD_SC_LP__AND4BB_2%X
x_PM_SKY130_FD_SC_LP__AND4BB_2%VGND N_VGND_M1013_d N_VGND_M1010_s N_VGND_M1014_d
+ N_VGND_c_627_n N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_664_n N_VGND_c_665_n
+ VGND N_VGND_c_630_n N_VGND_c_631_n N_VGND_c_632_n N_VGND_c_633_n
+ N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n N_VGND_c_637_n
+ PM_SKY130_FD_SC_LP__AND4BB_2%VGND
cc_1 VNB N_A_N_M1013_g 0.0332265f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.875
cc_2 VNB N_A_N_c_100_n 0.035645f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.675
cc_3 VNB N_A_N_c_101_n 0.0104537f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_4 VNB N_A_185_23#_M1006_g 0.0242581f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_5 VNB N_A_185_23#_M1003_g 0.0113815f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_6 VNB N_A_185_23#_c_125_n 0.00920232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_185_23#_M1010_g 0.0246632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_185_23#_c_127_n 0.0342354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_185_23#_M1012_g 0.00218363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_185_23#_c_129_n 0.0104645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_185_23#_c_130_n 0.00436379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_185_23#_c_131_n 0.0174869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_185_23#_c_132_n 0.00838102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_185_23#_c_133_n 0.00242388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_133#_M1015_g 0.0306571f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_A_27_133#_c_234_n 0.033573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_133#_c_235_n 0.0101733f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_18 VNB N_A_27_133#_c_236_n 0.0142618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_133#_c_237_n 0.00458406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_133#_c_238_n 0.00966895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_133#_c_239_n 0.00807664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_133#_c_240_n 0.00241892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_558_99#_c_335_n 0.0184164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_558_99#_c_336_n 0.0212341f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_25 VNB N_A_558_99#_c_337_n 0.0211552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_558_99#_c_338_n 0.0136064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_558_99#_c_339_n 4.82926e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_558_99#_c_340_n 0.0308863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_558_99#_c_341_n 0.00309688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_M1001_g 0.0397608f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.875
cc_31 VNB N_D_M1000_g 0.00876642f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.045
cc_32 VNB D 0.00840728f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_33 VNB N_D_c_445_n 0.0286909f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_34 VNB N_D_c_446_n 0.0166793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_N_M1005_g 0.0140215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_N_c_484_n 0.0109596f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_37 VNB N_B_N_c_485_n 0.0217301f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_38 VNB B_N 0.0208805f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_39 VNB N_B_N_c_487_n 0.0471932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_527_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_601_n 0.00392608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_627_n 0.017202f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_43 VNB N_VGND_c_628_n 0.0177247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_629_n 0.0180547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_630_n 0.0178607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_631_n 0.014949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_632_n 0.0498445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_633_n 0.0279842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_634_n 0.308945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_635_n 0.00740538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_636_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_637_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_A_N_c_100_n 0.00886429f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.675
cc_54 VPB N_A_N_M1009_g 0.0283179f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_55 VPB N_A_N_c_101_n 0.0092752f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_56 VPB N_A_185_23#_M1003_g 0.0216409f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_57 VPB N_A_185_23#_M1012_g 0.0228346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_185_23#_c_136_n 0.00698388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_185_23#_c_137_n 0.0107233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_185_23#_c_133_n 0.00237682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_27_133#_M1008_g 0.0369406f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_62 VPB N_A_27_133#_c_234_n 0.0187169f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_27_133#_c_235_n 6.56333e-19 $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_64 VPB N_A_27_133#_c_244_n 0.0354134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_27_133#_c_239_n 0.00332194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_27_133#_c_246_n 0.0120868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_27_133#_c_247_n 0.00193356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_27_133#_c_240_n 0.002077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_558_99#_M1004_g 0.0232769f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_70 VPB N_A_558_99#_c_336_n 7.75211e-19 $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_71 VPB N_A_558_99#_c_344_n 0.014556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_558_99#_c_338_n 0.0108705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_558_99#_c_339_n 7.51985e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_558_99#_c_347_n 0.0287175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_558_99#_c_341_n 0.00486653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_C_M1001_g 0.0317501f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.875
cc_77 VPB C 0.00580827f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_78 VPB N_C_c_413_n 0.0418098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_D_M1000_g 0.033649f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_80 VPB N_B_N_M1007_g 0.0287238f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_81 VPB N_B_N_c_485_n 0.00409126f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_82 VPB N_B_N_c_490_n 0.0112212f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.51
cc_83 VPB N_VPWR_c_528_n 0.0173181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_529_n 0.009635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_530_n 0.0287891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_531_n 0.032669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_532_n 0.00271811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_533_n 0.024312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_534_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_535_n 0.0147344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_536_n 0.0204301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_537_n 0.0217138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_527_n 0.121998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_539_n 0.0290503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_540_n 0.0413818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_541_n 0.00535984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_X_c_601_n 0.00163178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 N_A_N_M1013_g N_A_185_23#_M1006_g 0.00922272f $X=0.475 $Y=0.875 $X2=0
+ $Y2=0
cc_99 N_A_N_c_100_n N_A_185_23#_M1003_g 0.0234423f $X=0.54 $Y=1.675 $X2=0 $Y2=0
cc_100 N_A_N_c_100_n N_A_185_23#_c_129_n 0.00922272f $X=0.54 $Y=1.675 $X2=0
+ $Y2=0
cc_101 N_A_N_c_100_n N_A_27_133#_c_244_n 0.00139419f $X=0.54 $Y=1.675 $X2=0
+ $Y2=0
cc_102 N_A_N_M1009_g N_A_27_133#_c_244_n 0.0236845f $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_103 N_A_N_c_101_n N_A_27_133#_c_244_n 0.0297735f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_104 N_A_N_M1013_g N_A_27_133#_c_237_n 0.015703f $X=0.475 $Y=0.875 $X2=0 $Y2=0
cc_105 N_A_N_c_100_n N_A_27_133#_c_237_n 0.00287757f $X=0.54 $Y=1.675 $X2=0
+ $Y2=0
cc_106 N_A_N_c_101_n N_A_27_133#_c_237_n 0.0134159f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_107 N_A_N_c_100_n N_A_27_133#_c_238_n 0.00341464f $X=0.54 $Y=1.675 $X2=0
+ $Y2=0
cc_108 N_A_N_c_101_n N_A_27_133#_c_238_n 0.0211855f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A_N_M1013_g N_A_27_133#_c_239_n 0.00469497f $X=0.475 $Y=0.875 $X2=0
+ $Y2=0
cc_110 N_A_N_c_100_n N_A_27_133#_c_239_n 0.00576256f $X=0.54 $Y=1.675 $X2=0
+ $Y2=0
cc_111 N_A_N_c_101_n N_A_27_133#_c_239_n 0.0239842f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_112 N_A_N_M1009_g N_X_c_603_n 2.11244e-19 $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_113 N_A_N_M1013_g N_VGND_c_627_n 0.0124161f $X=0.475 $Y=0.875 $X2=0 $Y2=0
cc_114 N_A_N_M1013_g N_VGND_c_630_n 0.0032821f $X=0.475 $Y=0.875 $X2=0 $Y2=0
cc_115 N_A_N_M1013_g N_VGND_c_634_n 0.00385154f $X=0.475 $Y=0.875 $X2=0 $Y2=0
cc_116 N_A_185_23#_c_127_n N_A_27_133#_M1015_g 7.91673e-19 $X=1.495 $Y=1.615
+ $X2=0 $Y2=0
cc_117 N_A_185_23#_c_130_n N_A_27_133#_M1015_g 6.06825e-19 $X=1.585 $Y=1.45
+ $X2=0 $Y2=0
cc_118 N_A_185_23#_c_132_n N_A_27_133#_M1015_g 0.0194887f $X=2.475 $Y=0.922
+ $X2=0 $Y2=0
cc_119 N_A_185_23#_c_133_n N_A_27_133#_M1015_g 0.00619132f $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_120 N_A_185_23#_c_137_n N_A_27_133#_M1008_g 0.0239691f $X=2.602 $Y=2.02 $X2=0
+ $Y2=0
cc_121 N_A_185_23#_c_133_n N_A_27_133#_M1008_g 0.00964685f $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_122 N_A_185_23#_c_127_n N_A_27_133#_c_234_n 0.0176205f $X=1.495 $Y=1.615
+ $X2=0 $Y2=0
cc_123 N_A_185_23#_M1012_g N_A_27_133#_c_234_n 0.00183704f $X=1.495 $Y=2.465
+ $X2=0 $Y2=0
cc_124 N_A_185_23#_c_130_n N_A_27_133#_c_234_n 0.00106019f $X=1.585 $Y=1.45
+ $X2=0 $Y2=0
cc_125 N_A_185_23#_c_131_n N_A_27_133#_c_234_n 0.0018796f $X=2.125 $Y=0.922
+ $X2=0 $Y2=0
cc_126 N_A_185_23#_c_132_n N_A_27_133#_c_234_n 0.00749475f $X=2.475 $Y=0.922
+ $X2=0 $Y2=0
cc_127 N_A_185_23#_c_133_n N_A_27_133#_c_234_n 0.00720551f $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_128 N_A_185_23#_c_133_n N_A_27_133#_c_235_n 0.0060528f $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_129 N_A_185_23#_M1006_g N_A_27_133#_c_237_n 0.00167043f $X=1 $Y=0.665 $X2=0
+ $Y2=0
cc_130 N_A_185_23#_M1006_g N_A_27_133#_c_239_n 0.00204964f $X=1 $Y=0.665 $X2=0
+ $Y2=0
cc_131 N_A_185_23#_M1003_g N_A_27_133#_c_239_n 0.00382384f $X=1.065 $Y=2.465
+ $X2=0 $Y2=0
cc_132 N_A_185_23#_M1003_g N_A_27_133#_c_276_n 0.015497f $X=1.065 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_185_23#_M1012_g N_A_27_133#_c_276_n 0.0164441f $X=1.495 $Y=2.465
+ $X2=0 $Y2=0
cc_134 N_A_185_23#_c_137_n N_A_27_133#_c_278_n 0.00432482f $X=2.602 $Y=2.02
+ $X2=0 $Y2=0
cc_135 N_A_185_23#_c_131_n N_A_27_133#_c_246_n 0.00534668f $X=2.125 $Y=0.922
+ $X2=0 $Y2=0
cc_136 N_A_185_23#_c_133_n N_A_27_133#_c_246_n 0.0143487f $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_137 N_A_185_23#_c_127_n N_A_27_133#_c_247_n 0.00105269f $X=1.495 $Y=1.615
+ $X2=0 $Y2=0
cc_138 N_A_185_23#_M1012_g N_A_27_133#_c_247_n 0.00354552f $X=1.495 $Y=2.465
+ $X2=0 $Y2=0
cc_139 N_A_185_23#_c_130_n N_A_27_133#_c_247_n 0.011363f $X=1.585 $Y=1.45 $X2=0
+ $Y2=0
cc_140 N_A_185_23#_c_131_n N_A_27_133#_c_247_n 0.00118668f $X=2.125 $Y=0.922
+ $X2=0 $Y2=0
cc_141 N_A_185_23#_c_127_n N_A_27_133#_c_240_n 9.91333e-19 $X=1.495 $Y=1.615
+ $X2=0 $Y2=0
cc_142 N_A_185_23#_M1012_g N_A_27_133#_c_240_n 0.00246085f $X=1.495 $Y=2.465
+ $X2=0 $Y2=0
cc_143 N_A_185_23#_c_130_n N_A_27_133#_c_240_n 0.0165449f $X=1.585 $Y=1.45 $X2=0
+ $Y2=0
cc_144 N_A_185_23#_c_131_n N_A_27_133#_c_240_n 0.0211194f $X=2.125 $Y=0.922
+ $X2=0 $Y2=0
cc_145 N_A_185_23#_c_133_n N_A_27_133#_c_240_n 0.0324174f $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_146 N_A_185_23#_M1003_g N_A_27_133#_c_290_n 0.00799335f $X=1.065 $Y=2.465
+ $X2=0 $Y2=0
cc_147 N_A_185_23#_c_136_n N_A_558_99#_M1004_g 0.0128089f $X=3.485 $Y=2.02 $X2=0
+ $Y2=0
cc_148 N_A_185_23#_c_137_n N_A_558_99#_M1004_g 3.38716e-19 $X=2.602 $Y=2.02
+ $X2=0 $Y2=0
cc_149 N_A_185_23#_c_133_n N_A_558_99#_M1004_g 6.00027e-19 $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_150 N_A_185_23#_c_132_n N_A_558_99#_c_335_n 0.00317461f $X=2.475 $Y=0.922
+ $X2=0 $Y2=0
cc_151 N_A_185_23#_c_133_n N_A_558_99#_c_336_n 2.2098e-19 $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_152 N_A_185_23#_c_136_n N_A_558_99#_c_344_n 0.00438503f $X=3.485 $Y=2.02
+ $X2=0 $Y2=0
cc_153 N_A_185_23#_c_137_n N_A_558_99#_c_344_n 7.04201e-19 $X=2.602 $Y=2.02
+ $X2=0 $Y2=0
cc_154 N_A_185_23#_c_133_n N_A_558_99#_c_344_n 4.80068e-19 $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_155 N_A_185_23#_c_133_n N_A_558_99#_c_357_n 0.0189834f $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_156 N_A_185_23#_c_133_n N_A_558_99#_c_337_n 0.00162974f $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_157 N_A_185_23#_c_136_n N_A_558_99#_c_338_n 0.0471208f $X=3.485 $Y=2.02 $X2=0
+ $Y2=0
cc_158 N_A_185_23#_c_136_n N_A_558_99#_c_339_n 0.0233f $X=3.485 $Y=2.02 $X2=0
+ $Y2=0
cc_159 N_A_185_23#_c_137_n N_A_558_99#_c_339_n 0.00205458f $X=2.602 $Y=2.02
+ $X2=0 $Y2=0
cc_160 N_A_185_23#_c_133_n N_A_558_99#_c_339_n 0.0106953f $X=2.602 $Y=1.935
+ $X2=0 $Y2=0
cc_161 N_A_185_23#_c_136_n N_A_558_99#_c_347_n 0.00528519f $X=3.485 $Y=2.02
+ $X2=0 $Y2=0
cc_162 N_A_185_23#_c_188_p N_A_558_99#_c_347_n 3.94582e-19 $X=3.62 $Y=2.285
+ $X2=0 $Y2=0
cc_163 N_A_185_23#_c_136_n N_C_M1001_g 0.0123167f $X=3.485 $Y=2.02 $X2=0 $Y2=0
cc_164 N_A_185_23#_c_136_n C 0.00379006f $X=3.485 $Y=2.02 $X2=0 $Y2=0
cc_165 N_A_185_23#_c_188_p C 0.0142911f $X=3.62 $Y=2.285 $X2=0 $Y2=0
cc_166 N_A_185_23#_c_136_n N_C_c_413_n 2.15682e-19 $X=3.485 $Y=2.02 $X2=0 $Y2=0
cc_167 N_A_185_23#_c_188_p N_C_c_413_n 0.00202174f $X=3.62 $Y=2.285 $X2=0 $Y2=0
cc_168 N_A_185_23#_c_136_n N_D_M1000_g 0.00267298f $X=3.485 $Y=2.02 $X2=0 $Y2=0
cc_169 N_A_185_23#_c_136_n N_VPWR_M1004_d 0.00217806f $X=3.485 $Y=2.02 $X2=0
+ $Y2=0
cc_170 N_A_185_23#_M1003_g N_VPWR_c_528_n 0.0129267f $X=1.065 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_185_23#_M1012_g N_VPWR_c_528_n 0.00151645f $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_185_23#_M1012_g N_VPWR_c_529_n 0.00484924f $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_185_23#_c_188_p N_VPWR_c_531_n 0.0247708f $X=3.62 $Y=2.285 $X2=0
+ $Y2=0
cc_174 N_A_185_23#_c_136_n N_VPWR_c_532_n 0.017091f $X=3.485 $Y=2.02 $X2=0 $Y2=0
cc_175 N_A_185_23#_M1003_g N_VPWR_c_535_n 0.00486043f $X=1.065 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_185_23#_M1012_g N_VPWR_c_535_n 0.00487821f $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_185_23#_M1003_g N_VPWR_c_527_n 0.00448287f $X=1.065 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_185_23#_M1012_g N_VPWR_c_527_n 0.00448292f $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A_185_23#_M1003_g N_VPWR_c_540_n 0.0015287f $X=1.065 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_185_23#_M1012_g N_VPWR_c_540_n 0.0135993f $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_185_23#_M1003_g N_X_c_603_n 0.00457203f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A_185_23#_c_125_n N_X_c_603_n 8.28374e-19 $X=1.355 $Y=1.36 $X2=0 $Y2=0
cc_183 N_A_185_23#_M1012_g N_X_c_603_n 0.00443291f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_185_23#_M1006_g N_X_c_601_n 0.00223038f $X=1 $Y=0.665 $X2=0 $Y2=0
cc_185 N_A_185_23#_M1003_g N_X_c_601_n 0.0103328f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_185_23#_c_125_n N_X_c_601_n 0.00867609f $X=1.355 $Y=1.36 $X2=0 $Y2=0
cc_187 N_A_185_23#_M1010_g N_X_c_601_n 0.0020178f $X=1.43 $Y=0.665 $X2=0 $Y2=0
cc_188 N_A_185_23#_c_127_n N_X_c_601_n 0.00450245f $X=1.495 $Y=1.615 $X2=0 $Y2=0
cc_189 N_A_185_23#_c_129_n N_X_c_601_n 0.00219459f $X=1.032 $Y=1.36 $X2=0 $Y2=0
cc_190 N_A_185_23#_c_130_n N_X_c_601_n 0.032687f $X=1.585 $Y=1.45 $X2=0 $Y2=0
cc_191 N_A_185_23#_c_217_p N_X_c_601_n 0.0111029f $X=1.75 $Y=1.085 $X2=0 $Y2=0
cc_192 N_A_185_23#_c_217_p N_VGND_M1010_s 0.00238736f $X=1.75 $Y=1.085 $X2=0
+ $Y2=0
cc_193 N_A_185_23#_c_131_n N_VGND_M1010_s 2.95928e-19 $X=2.125 $Y=0.922 $X2=0
+ $Y2=0
cc_194 N_A_185_23#_M1006_g N_VGND_c_627_n 0.0052368f $X=1 $Y=0.665 $X2=0 $Y2=0
cc_195 N_A_185_23#_M1006_g N_VGND_c_628_n 6.08243e-19 $X=1 $Y=0.665 $X2=0 $Y2=0
cc_196 N_A_185_23#_M1010_g N_VGND_c_628_n 0.011099f $X=1.43 $Y=0.665 $X2=0 $Y2=0
cc_197 N_A_185_23#_c_127_n N_VGND_c_628_n 9.253e-19 $X=1.495 $Y=1.615 $X2=0
+ $Y2=0
cc_198 N_A_185_23#_c_217_p N_VGND_c_628_n 0.0188108f $X=1.75 $Y=1.085 $X2=0
+ $Y2=0
cc_199 N_A_185_23#_c_131_n N_VGND_c_628_n 0.00490349f $X=2.125 $Y=0.922 $X2=0
+ $Y2=0
cc_200 N_A_185_23#_c_132_n N_VGND_c_628_n 0.00856491f $X=2.475 $Y=0.922 $X2=0
+ $Y2=0
cc_201 N_A_185_23#_M1006_g N_VGND_c_631_n 0.00575161f $X=1 $Y=0.665 $X2=0 $Y2=0
cc_202 N_A_185_23#_M1010_g N_VGND_c_631_n 0.00477554f $X=1.43 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_185_23#_c_132_n N_VGND_c_632_n 0.00697628f $X=2.475 $Y=0.922 $X2=0
+ $Y2=0
cc_204 N_A_185_23#_M1006_g N_VGND_c_634_n 0.0118487f $X=1 $Y=0.665 $X2=0 $Y2=0
cc_205 N_A_185_23#_M1010_g N_VGND_c_634_n 0.00825815f $X=1.43 $Y=0.665 $X2=0
+ $Y2=0
cc_206 N_A_185_23#_c_132_n N_VGND_c_634_n 0.0125029f $X=2.475 $Y=0.922 $X2=0
+ $Y2=0
cc_207 N_A_27_133#_M1008_g N_A_558_99#_M1004_g 0.0175743f $X=2.505 $Y=2.285
+ $X2=0 $Y2=0
cc_208 N_A_27_133#_M1015_g N_A_558_99#_c_335_n 0.0277438f $X=2.505 $Y=0.835
+ $X2=0 $Y2=0
cc_209 N_A_27_133#_M1008_g N_A_558_99#_c_336_n 0.0277438f $X=2.505 $Y=2.285
+ $X2=0 $Y2=0
cc_210 N_A_27_133#_M1015_g N_A_558_99#_c_357_n 0.00125794f $X=2.505 $Y=0.835
+ $X2=0 $Y2=0
cc_211 N_A_27_133#_c_235_n N_A_558_99#_c_337_n 0.0277438f $X=2.505 $Y=1.51 $X2=0
+ $Y2=0
cc_212 N_A_27_133#_c_235_n N_A_558_99#_c_339_n 6.29756e-19 $X=2.505 $Y=1.51
+ $X2=0 $Y2=0
cc_213 N_A_27_133#_c_244_n N_VPWR_M1009_d 0.0011474f $X=0.73 $Y=2.152 $X2=-0.19
+ $Y2=-0.245
cc_214 N_A_27_133#_c_239_n N_VPWR_M1009_d 0.0021297f $X=0.815 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A_27_133#_c_276_n N_VPWR_M1009_d 0.00155461f $X=1.615 $Y=2.47 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A_27_133#_c_290_n N_VPWR_M1009_d 0.0162358f $X=0.815 $Y=2.237 $X2=-0.19
+ $Y2=-0.245
cc_217 N_A_27_133#_c_276_n N_VPWR_M1012_s 0.00378709f $X=1.615 $Y=2.47 $X2=0
+ $Y2=0
cc_218 N_A_27_133#_c_278_n N_VPWR_M1012_s 0.0078292f $X=1.7 $Y=2.385 $X2=0 $Y2=0
cc_219 N_A_27_133#_c_246_n N_VPWR_M1012_s 0.00216525f $X=1.96 $Y=1.88 $X2=0
+ $Y2=0
cc_220 N_A_27_133#_c_247_n N_VPWR_M1012_s 0.00113247f $X=1.785 $Y=1.88 $X2=0
+ $Y2=0
cc_221 N_A_27_133#_c_244_n N_VPWR_c_528_n 0.00242386f $X=0.73 $Y=2.152 $X2=0
+ $Y2=0
cc_222 N_A_27_133#_c_276_n N_VPWR_c_528_n 0.00431593f $X=1.615 $Y=2.47 $X2=0
+ $Y2=0
cc_223 N_A_27_133#_c_290_n N_VPWR_c_528_n 0.0147871f $X=0.815 $Y=2.237 $X2=0
+ $Y2=0
cc_224 N_A_27_133#_M1008_g N_VPWR_c_529_n 0.00813662f $X=2.505 $Y=2.285 $X2=0
+ $Y2=0
cc_225 N_A_27_133#_c_234_n N_VPWR_c_529_n 0.00108803f $X=2.43 $Y=1.51 $X2=0
+ $Y2=0
cc_226 N_A_27_133#_c_276_n N_VPWR_c_529_n 0.0143446f $X=1.615 $Y=2.47 $X2=0
+ $Y2=0
cc_227 N_A_27_133#_c_278_n N_VPWR_c_529_n 0.018746f $X=1.7 $Y=2.385 $X2=0 $Y2=0
cc_228 N_A_27_133#_c_246_n N_VPWR_c_529_n 0.0236431f $X=1.96 $Y=1.88 $X2=0 $Y2=0
cc_229 N_A_27_133#_M1008_g N_VPWR_c_530_n 5.16824e-19 $X=2.505 $Y=2.285 $X2=0
+ $Y2=0
cc_230 N_A_27_133#_M1008_g N_VPWR_c_532_n 2.72131e-19 $X=2.505 $Y=2.285 $X2=0
+ $Y2=0
cc_231 N_A_27_133#_M1008_g N_VPWR_c_533_n 0.00320058f $X=2.505 $Y=2.285 $X2=0
+ $Y2=0
cc_232 N_A_27_133#_M1008_g N_VPWR_c_527_n 0.00415093f $X=2.505 $Y=2.285 $X2=0
+ $Y2=0
cc_233 N_A_27_133#_c_276_n N_VPWR_c_527_n 0.0189497f $X=1.615 $Y=2.47 $X2=0
+ $Y2=0
cc_234 N_A_27_133#_c_290_n N_VPWR_c_527_n 6.78937e-19 $X=0.815 $Y=2.237 $X2=0
+ $Y2=0
cc_235 N_A_27_133#_c_276_n N_VPWR_c_540_n 0.0155592f $X=1.615 $Y=2.47 $X2=0
+ $Y2=0
cc_236 N_A_27_133#_c_276_n N_X_M1003_d 0.00491884f $X=1.615 $Y=2.47 $X2=0 $Y2=0
cc_237 N_A_27_133#_c_276_n N_X_c_603_n 0.0184057f $X=1.615 $Y=2.47 $X2=0 $Y2=0
cc_238 N_A_27_133#_c_290_n N_X_c_603_n 0.0222221f $X=0.815 $Y=2.237 $X2=0 $Y2=0
cc_239 N_A_27_133#_c_237_n N_X_c_601_n 0.0131561f $X=0.73 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_27_133#_c_239_n N_X_c_601_n 0.0472211f $X=0.815 $Y=1.92 $X2=0 $Y2=0
cc_241 N_A_27_133#_c_247_n N_X_c_601_n 0.00471491f $X=1.785 $Y=1.88 $X2=0 $Y2=0
cc_242 N_A_27_133#_c_240_n N_X_c_601_n 0.00530776f $X=2.125 $Y=1.51 $X2=0 $Y2=0
cc_243 N_A_27_133#_c_290_n N_X_c_601_n 0.00115595f $X=0.815 $Y=2.237 $X2=0 $Y2=0
cc_244 N_A_27_133#_c_237_n N_VGND_M1013_d 0.00290041f $X=0.73 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_245 N_A_27_133#_c_237_n N_VGND_c_627_n 0.024199f $X=0.73 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A_27_133#_M1015_g N_VGND_c_628_n 0.00376765f $X=2.505 $Y=0.835 $X2=0
+ $Y2=0
cc_247 N_A_27_133#_c_236_n N_VGND_c_630_n 0.00412822f $X=0.26 $Y=0.875 $X2=0
+ $Y2=0
cc_248 N_A_27_133#_M1015_g N_VGND_c_632_n 0.00335368f $X=2.505 $Y=0.835 $X2=0
+ $Y2=0
cc_249 N_A_27_133#_M1015_g N_VGND_c_634_n 0.00469432f $X=2.505 $Y=0.835 $X2=0
+ $Y2=0
cc_250 N_A_27_133#_c_236_n N_VGND_c_634_n 0.00732126f $X=0.26 $Y=0.875 $X2=0
+ $Y2=0
cc_251 N_A_558_99#_M1004_g N_C_M1001_g 0.017809f $X=2.935 $Y=2.285 $X2=0 $Y2=0
cc_252 N_A_558_99#_c_335_n N_C_M1001_g 0.022465f $X=2.955 $Y=1.165 $X2=0 $Y2=0
cc_253 N_A_558_99#_c_357_n N_C_M1001_g 0.00168012f $X=2.955 $Y=1.33 $X2=0 $Y2=0
cc_254 N_A_558_99#_c_337_n N_C_M1001_g 0.0425666f $X=2.955 $Y=1.33 $X2=0 $Y2=0
cc_255 N_A_558_99#_c_338_n N_C_M1001_g 0.0129624f $X=4.355 $Y=1.675 $X2=0 $Y2=0
cc_256 N_A_558_99#_c_338_n N_D_M1000_g 0.0148479f $X=4.355 $Y=1.675 $X2=0 $Y2=0
cc_257 N_A_558_99#_c_340_n N_D_M1000_g 5.02215e-19 $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_258 N_A_558_99#_c_347_n N_D_M1000_g 0.00132177f $X=4.52 $Y=2.285 $X2=0 $Y2=0
cc_259 N_A_558_99#_c_357_n D 0.00876031f $X=2.955 $Y=1.33 $X2=0 $Y2=0
cc_260 N_A_558_99#_c_337_n D 8.93757e-19 $X=2.955 $Y=1.33 $X2=0 $Y2=0
cc_261 N_A_558_99#_c_338_n D 0.0576745f $X=4.355 $Y=1.675 $X2=0 $Y2=0
cc_262 N_A_558_99#_c_340_n D 0.0196092f $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_263 N_A_558_99#_c_338_n N_D_c_445_n 0.00483619f $X=4.355 $Y=1.675 $X2=0 $Y2=0
cc_264 N_A_558_99#_c_340_n N_D_c_445_n 7.25864e-19 $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_265 N_A_558_99#_c_340_n N_D_c_446_n 5.85067e-19 $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_266 N_A_558_99#_c_340_n N_B_N_M1005_g 0.00751726f $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_267 N_A_558_99#_c_347_n N_B_N_M1007_g 0.0132951f $X=4.52 $Y=2.285 $X2=0 $Y2=0
cc_268 N_A_558_99#_c_338_n N_B_N_c_484_n 6.34754e-19 $X=4.355 $Y=1.675 $X2=0
+ $Y2=0
cc_269 N_A_558_99#_c_340_n N_B_N_c_484_n 0.00558255f $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_270 N_A_558_99#_c_338_n N_B_N_c_485_n 0.00717957f $X=4.355 $Y=1.675 $X2=0
+ $Y2=0
cc_271 N_A_558_99#_c_340_n N_B_N_c_485_n 0.0103046f $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_272 N_A_558_99#_c_341_n N_B_N_c_485_n 0.00346199f $X=4.52 $Y=1.675 $X2=0
+ $Y2=0
cc_273 N_A_558_99#_c_338_n N_B_N_c_490_n 0.00673912f $X=4.355 $Y=1.675 $X2=0
+ $Y2=0
cc_274 N_A_558_99#_c_347_n N_B_N_c_490_n 0.00515908f $X=4.52 $Y=2.285 $X2=0
+ $Y2=0
cc_275 N_A_558_99#_c_341_n N_B_N_c_490_n 9.96256e-19 $X=4.52 $Y=1.675 $X2=0
+ $Y2=0
cc_276 N_A_558_99#_M1005_d B_N 0.00335558f $X=4.38 $Y=0.625 $X2=0 $Y2=0
cc_277 N_A_558_99#_c_340_n B_N 0.0192952f $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_278 N_A_558_99#_c_340_n N_B_N_c_487_n 3.15414e-19 $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_279 N_A_558_99#_M1004_g N_VPWR_c_530_n 0.00333885f $X=2.935 $Y=2.285 $X2=0
+ $Y2=0
cc_280 N_A_558_99#_c_338_n N_VPWR_c_531_n 0.0115477f $X=4.355 $Y=1.675 $X2=0
+ $Y2=0
cc_281 N_A_558_99#_M1004_g N_VPWR_c_532_n 0.00370625f $X=2.935 $Y=2.285 $X2=0
+ $Y2=0
cc_282 N_A_558_99#_M1004_g N_VPWR_c_533_n 0.00266097f $X=2.935 $Y=2.285 $X2=0
+ $Y2=0
cc_283 N_A_558_99#_M1004_g N_VPWR_c_527_n 0.00348678f $X=2.935 $Y=2.285 $X2=0
+ $Y2=0
cc_284 N_A_558_99#_c_335_n N_VGND_c_629_n 0.00155542f $X=2.955 $Y=1.165 $X2=0
+ $Y2=0
cc_285 N_A_558_99#_c_335_n N_VGND_c_664_n 9.04178e-19 $X=2.955 $Y=1.165 $X2=0
+ $Y2=0
cc_286 N_A_558_99#_c_340_n N_VGND_c_665_n 0.0132351f $X=4.52 $Y=0.92 $X2=0 $Y2=0
cc_287 N_A_558_99#_c_335_n N_VGND_c_632_n 0.00415323f $X=2.955 $Y=1.165 $X2=0
+ $Y2=0
cc_288 N_A_558_99#_c_335_n N_VGND_c_634_n 0.00469432f $X=2.955 $Y=1.165 $X2=0
+ $Y2=0
cc_289 N_A_558_99#_c_340_n N_VGND_c_634_n 0.00210288f $X=4.52 $Y=0.92 $X2=0
+ $Y2=0
cc_290 N_C_M1001_g N_D_M1000_g 0.0295066f $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_291 N_C_M1001_g D 0.00890406f $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_292 N_C_M1001_g N_D_c_446_n 0.0643349f $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_293 N_C_M1001_g N_VPWR_c_530_n 0.0043984f $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_294 C N_VPWR_c_530_n 0.0240707f $X=3.515 $Y=2.69 $X2=0 $Y2=0
cc_295 N_C_c_413_n N_VPWR_c_530_n 0.00810943f $X=3.42 $Y=2.855 $X2=0 $Y2=0
cc_296 N_C_M1001_g N_VPWR_c_531_n 0.00255181f $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_297 C N_VPWR_c_531_n 0.0275035f $X=3.515 $Y=2.69 $X2=0 $Y2=0
cc_298 N_C_c_413_n N_VPWR_c_531_n 0.00166495f $X=3.42 $Y=2.855 $X2=0 $Y2=0
cc_299 N_C_M1001_g N_VPWR_c_532_n 3.5651e-19 $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_300 N_C_c_413_n N_VPWR_c_532_n 0.00234537f $X=3.42 $Y=2.855 $X2=0 $Y2=0
cc_301 C N_VPWR_c_536_n 0.0193391f $X=3.515 $Y=2.69 $X2=0 $Y2=0
cc_302 N_C_c_413_n N_VPWR_c_536_n 0.00832175f $X=3.42 $Y=2.855 $X2=0 $Y2=0
cc_303 C N_VPWR_c_527_n 0.0146107f $X=3.515 $Y=2.69 $X2=0 $Y2=0
cc_304 N_C_c_413_n N_VPWR_c_527_n 0.0108081f $X=3.42 $Y=2.855 $X2=0 $Y2=0
cc_305 N_C_M1001_g N_VGND_c_629_n 0.0108953f $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_306 N_C_M1001_g N_VGND_c_664_n 0.00668728f $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_307 N_C_M1001_g N_VGND_c_632_n 0.00289833f $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_308 N_C_M1001_g N_VGND_c_634_n 0.00331732f $X=3.405 $Y=0.835 $X2=0 $Y2=0
cc_309 N_D_c_446_n N_B_N_M1005_g 0.0130192f $X=3.855 $Y=1.155 $X2=0 $Y2=0
cc_310 D N_B_N_c_484_n 9.19193e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_311 N_D_c_445_n N_B_N_c_484_n 0.00904343f $X=3.855 $Y=1.32 $X2=0 $Y2=0
cc_312 N_D_M1000_g N_B_N_c_485_n 0.00939986f $X=3.87 $Y=2.285 $X2=0 $Y2=0
cc_313 D N_B_N_c_485_n 7.84305e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_314 N_D_c_445_n N_B_N_c_485_n 0.00933596f $X=3.855 $Y=1.32 $X2=0 $Y2=0
cc_315 N_D_M1000_g N_B_N_c_490_n 0.0213509f $X=3.87 $Y=2.285 $X2=0 $Y2=0
cc_316 D B_N 0.0012153f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_317 N_D_c_446_n B_N 0.00129289f $X=3.855 $Y=1.155 $X2=0 $Y2=0
cc_318 N_D_c_446_n N_B_N_c_487_n 7.35477e-19 $X=3.855 $Y=1.155 $X2=0 $Y2=0
cc_319 N_D_M1000_g N_VPWR_c_531_n 0.0103104f $X=3.87 $Y=2.285 $X2=0 $Y2=0
cc_320 N_D_M1000_g N_VPWR_c_536_n 0.00234092f $X=3.87 $Y=2.285 $X2=0 $Y2=0
cc_321 N_D_M1000_g N_VPWR_c_527_n 0.00307168f $X=3.87 $Y=2.285 $X2=0 $Y2=0
cc_322 N_D_c_446_n N_VGND_c_629_n 0.0112137f $X=3.855 $Y=1.155 $X2=0 $Y2=0
cc_323 D N_VGND_c_664_n 0.0226929f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_324 N_D_c_446_n N_VGND_c_664_n 0.00444032f $X=3.855 $Y=1.155 $X2=0 $Y2=0
cc_325 D N_VGND_c_665_n 0.0250001f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_326 N_D_c_445_n N_VGND_c_665_n 0.00445684f $X=3.855 $Y=1.32 $X2=0 $Y2=0
cc_327 N_D_c_446_n N_VGND_c_665_n 0.00335672f $X=3.855 $Y=1.155 $X2=0 $Y2=0
cc_328 N_D_c_446_n N_VGND_c_633_n 0.0017908f $X=3.855 $Y=1.155 $X2=0 $Y2=0
cc_329 N_D_c_446_n N_VGND_c_634_n 0.0020655f $X=3.855 $Y=1.155 $X2=0 $Y2=0
cc_330 N_B_N_M1007_g N_VPWR_c_531_n 0.00350877f $X=4.305 $Y=2.285 $X2=0 $Y2=0
cc_331 N_B_N_M1007_g N_VPWR_c_537_n 0.00320058f $X=4.305 $Y=2.285 $X2=0 $Y2=0
cc_332 N_B_N_M1007_g N_VPWR_c_527_n 0.00415093f $X=4.305 $Y=2.285 $X2=0 $Y2=0
cc_333 B_N N_VGND_M1014_d 0.00283965f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_334 N_B_N_M1005_g N_VGND_c_629_n 9.80689e-19 $X=4.305 $Y=0.835 $X2=0 $Y2=0
cc_335 B_N N_VGND_c_629_n 0.0342374f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_336 N_B_N_c_487_n N_VGND_c_629_n 0.00276853f $X=4.305 $Y=0.35 $X2=0 $Y2=0
cc_337 N_B_N_M1005_g N_VGND_c_665_n 0.00181674f $X=4.305 $Y=0.835 $X2=0 $Y2=0
cc_338 B_N N_VGND_c_665_n 0.0152284f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_339 B_N N_VGND_c_633_n 0.0467974f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_340 N_B_N_c_487_n N_VGND_c_633_n 0.00647615f $X=4.305 $Y=0.35 $X2=0 $Y2=0
cc_341 B_N N_VGND_c_634_n 0.0253178f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_342 N_B_N_c_487_n N_VGND_c_634_n 0.00988008f $X=4.305 $Y=0.35 $X2=0 $Y2=0
cc_343 N_VPWR_c_527_n N_X_M1003_d 0.00383613f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_344 N_X_c_601_n N_VGND_c_631_n 0.0138717f $X=1.215 $Y=0.42 $X2=0 $Y2=0
cc_345 N_X_M1006_d N_VGND_c_634_n 0.00397496f $X=1.075 $Y=0.245 $X2=0 $Y2=0
cc_346 N_X_c_601_n N_VGND_c_634_n 0.00886411f $X=1.215 $Y=0.42 $X2=0 $Y2=0
cc_347 N_VGND_c_664_n A_696_125# 0.00106497f $X=3.775 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
