* NGSPICE file created from sky130_fd_sc_lp__a221oi_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a221oi_m A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_296_535# VPB phighvt w=420000u l=150000u
+  ad=1.974e+11p pd=1.78e+06u as=2.352e+11p ps=2.8e+06u
M1001 a_226_55# B2 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.289e+11p ps=2.77e+06u
M1002 Y B1 a_226_55# VNB nshort w=420000u l=150000u
+  ad=2.751e+11p pd=2.99e+06u as=0p ps=0u
M1003 a_210_535# B1 a_296_535# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1004 a_406_55# A1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 a_296_535# B2 a_210_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_406_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_210_535# C1 Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 a_296_535# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

