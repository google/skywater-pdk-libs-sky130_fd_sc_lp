* File: sky130_fd_sc_lp__decapkapwr_8.pxi.spice
* Created: Wed Sep  2 09:42:47 2020
* 
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_8%VGND N_VGND_M1000_s N_VGND_c_26_n
+ N_VGND_c_27_n N_VGND_c_28_n N_VGND_c_29_n N_VGND_c_30_n VGND N_VGND_M1001_g
+ N_VGND_c_31_n N_VGND_c_32_n N_VGND_c_33_n N_VGND_c_34_n N_VGND_c_35_n
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_8%VGND
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_8%KAPWR N_KAPWR_M1001_s N_KAPWR_c_59_n
+ N_KAPWR_c_60_n N_KAPWR_c_69_n N_KAPWR_c_57_n N_KAPWR_c_58_n N_KAPWR_c_63_n
+ N_KAPWR_c_64_n KAPWR N_KAPWR_M1000_g N_KAPWR_c_65_n KAPWR
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_8%KAPWR
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_8%VPWR VPWR N_VPWR_c_93_n VPWR
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_8%VPWR
cc_1 VNB N_VGND_c_26_n 0.0651019f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=0.38
cc_2 VNB N_VGND_c_27_n 0.00211035f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.77
cc_3 VNB N_VGND_c_28_n 4.60769e-19 $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.77
cc_4 VNB N_VGND_c_29_n 0.0193278f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.77
cc_5 VNB N_VGND_c_30_n 0.0365902f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=0.36
cc_6 VNB N_VGND_c_31_n 0.0598957f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=0
cc_7 VNB N_VGND_c_32_n 0.0206f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=0
cc_8 VNB N_VGND_c_33_n 0.2505f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=0
cc_9 VNB N_VGND_c_34_n 0.0279619f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_10 VNB N_VGND_c_35_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=0
cc_11 VNB N_KAPWR_c_57_n 0.0287929f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.06
cc_12 VNB N_KAPWR_c_58_n 0.209886f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.77
cc_13 VNB VPWR 0.163682f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.235
cc_14 VPB N_VGND_c_27_n 0.0140672f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.77
cc_15 VPB N_VGND_c_28_n 0.00877216f $X=-0.19 $Y=1.655 $X2=1.395 $Y2=1.77
cc_16 VPB N_VGND_c_29_n 0.222588f $X=-0.19 $Y=1.655 $X2=1.395 $Y2=1.77
cc_17 VPB N_KAPWR_c_59_n 0.0111229f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_18 VPB N_KAPWR_c_60_n 0.0291277f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=0.085
cc_19 VPB N_KAPWR_c_57_n 0.00109678f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=1.06
cc_20 VPB N_KAPWR_c_58_n 0.0210044f $X=-0.19 $Y=1.655 $X2=1.395 $Y2=1.77
cc_21 VPB N_KAPWR_c_63_n 0.0109168f $X=-0.19 $Y=1.655 $X2=3.095 $Y2=0.36
cc_22 VPB N_KAPWR_c_64_n 0.0514848f $X=-0.19 $Y=1.655 $X2=3.095 $Y2=1.04
cc_23 VPB N_KAPWR_c_65_n 0.0648142f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=0
cc_24 VPB VPWR 0.051391f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.235
cc_25 VPB N_VPWR_c_93_n 0.104947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 N_VGND_c_29_n N_KAPWR_c_59_n 0.00701606f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_27 N_VGND_c_27_n N_KAPWR_c_60_n 0.0205458f $X=0.98 $Y=1.77 $X2=0 $Y2=0
cc_28 N_VGND_c_29_n N_KAPWR_c_60_n 0.0287446f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_29 N_VGND_c_29_n N_KAPWR_c_69_n 0.117197f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_30 N_VGND_c_28_n N_KAPWR_c_57_n 0.00290374f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_31 N_VGND_c_29_n N_KAPWR_c_57_n 0.00707553f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_32 N_VGND_c_30_n N_KAPWR_c_57_n 0.0230356f $X=3.095 $Y=0.36 $X2=0 $Y2=0
cc_33 N_VGND_c_26_n N_KAPWR_c_58_n 0.0654854f $X=0.815 $Y=0.38 $X2=0 $Y2=0
cc_34 N_VGND_c_28_n N_KAPWR_c_58_n 0.00447085f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_35 N_VGND_c_29_n N_KAPWR_c_58_n 0.127128f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_36 N_VGND_c_30_n N_KAPWR_c_58_n 0.0510144f $X=3.095 $Y=0.36 $X2=0 $Y2=0
cc_37 N_VGND_c_31_n N_KAPWR_c_58_n 0.0760645f $X=2.93 $Y=0 $X2=0 $Y2=0
cc_38 N_VGND_c_33_n N_KAPWR_c_58_n 0.120027f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_39 N_VGND_c_29_n N_KAPWR_c_63_n 0.00748742f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_40 N_VGND_c_29_n N_KAPWR_c_64_n 0.0451651f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_41 N_VGND_c_29_n N_KAPWR_c_65_n 0.0972887f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_42 N_VGND_c_29_n VPWR 0.046619f $X=1.395 $Y=1.77 $X2=-0.19 $Y2=-0.245
cc_43 N_VGND_c_29_n N_VPWR_c_93_n 0.0524183f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_44 N_KAPWR_M1001_s VPWR 0.00234386f $X=0.615 $Y=2.095 $X2=-0.19 $Y2=-0.245
cc_45 N_KAPWR_c_59_n VPWR 0.00381888f $X=0.7 $Y=2.675 $X2=-0.19 $Y2=-0.245
cc_46 N_KAPWR_c_69_n VPWR 0.0106097f $X=2.865 $Y=2.81 $X2=-0.19 $Y2=-0.245
cc_47 N_KAPWR_c_63_n VPWR 0.00389737f $X=3.075 $Y=2.675 $X2=-0.19 $Y2=-0.245
cc_48 N_KAPWR_c_65_n VPWR 0.395208f $X=3.11 $Y=2.81 $X2=-0.19 $Y2=-0.245
cc_49 N_KAPWR_c_59_n N_VPWR_c_93_n 0.0269429f $X=0.7 $Y=2.675 $X2=0 $Y2=0
cc_50 N_KAPWR_c_69_n N_VPWR_c_93_n 0.0690021f $X=2.865 $Y=2.81 $X2=0 $Y2=0
cc_51 N_KAPWR_c_63_n N_VPWR_c_93_n 0.0275782f $X=3.075 $Y=2.675 $X2=0 $Y2=0
cc_52 N_KAPWR_c_65_n N_VPWR_c_93_n 0.0103135f $X=3.11 $Y=2.81 $X2=0 $Y2=0
