* File: sky130_fd_sc_lp__mux4_4.pxi.spice
* Created: Wed Sep  2 10:02:07 2020
* 
x_PM_SKY130_FD_SC_LP__MUX4_4%A_84_277# N_A_84_277#_M1007_s N_A_84_277#_M1016_s
+ N_A_84_277#_M1031_g N_A_84_277#_c_177_n N_A_84_277#_c_178_n
+ N_A_84_277#_M1006_g N_A_84_277#_c_180_n N_A_84_277#_c_181_n
+ N_A_84_277#_c_187_n N_A_84_277#_c_182_n N_A_84_277#_c_183_n
+ N_A_84_277#_c_184_n N_A_84_277#_c_185_n PM_SKY130_FD_SC_LP__MUX4_4%A_84_277#
x_PM_SKY130_FD_SC_LP__MUX4_4%S1 N_S1_M1008_g N_S1_c_233_n N_S1_c_234_n
+ N_S1_c_238_n N_S1_M1009_g N_S1_c_239_n N_S1_c_240_n N_S1_M1016_g N_S1_M1007_g
+ S1 S1 S1 N_S1_c_237_n PM_SKY130_FD_SC_LP__MUX4_4%S1
x_PM_SKY130_FD_SC_LP__MUX4_4%A_114_119# N_A_114_119#_M1008_d
+ N_A_114_119#_M1031_d N_A_114_119#_M1005_g N_A_114_119#_c_301_n
+ N_A_114_119#_M1014_g N_A_114_119#_M1011_g N_A_114_119#_c_302_n
+ N_A_114_119#_M1015_g N_A_114_119#_M1018_g N_A_114_119#_c_303_n
+ N_A_114_119#_M1024_g N_A_114_119#_M1022_g N_A_114_119#_c_304_n
+ N_A_114_119#_M1027_g N_A_114_119#_c_305_n N_A_114_119#_c_306_n
+ N_A_114_119#_c_307_n N_A_114_119#_c_308_n N_A_114_119#_c_359_p
+ N_A_114_119#_c_325_n N_A_114_119#_c_309_n N_A_114_119#_c_310_n
+ N_A_114_119#_c_395_p N_A_114_119#_c_311_n
+ PM_SKY130_FD_SC_LP__MUX4_4%A_114_119#
x_PM_SKY130_FD_SC_LP__MUX4_4%A1 N_A1_M1001_g N_A1_M1004_g A1 A1 N_A1_c_439_n
+ PM_SKY130_FD_SC_LP__MUX4_4%A1
x_PM_SKY130_FD_SC_LP__MUX4_4%A_1041_333# N_A_1041_333#_M1021_d
+ N_A_1041_333#_M1026_d N_A_1041_333#_M1000_g N_A_1041_333#_M1002_g
+ N_A_1041_333#_M1013_g N_A_1041_333#_M1023_g N_A_1041_333#_c_482_n
+ N_A_1041_333#_c_483_n N_A_1041_333#_c_484_n N_A_1041_333#_c_485_n
+ N_A_1041_333#_c_497_n N_A_1041_333#_c_486_n N_A_1041_333#_c_487_n
+ N_A_1041_333#_c_488_n N_A_1041_333#_c_499_n N_A_1041_333#_c_538_p
+ N_A_1041_333#_c_500_n N_A_1041_333#_c_501_n N_A_1041_333#_c_489_n
+ N_A_1041_333#_c_490_n N_A_1041_333#_c_491_n N_A_1041_333#_c_492_n
+ PM_SKY130_FD_SC_LP__MUX4_4%A_1041_333#
x_PM_SKY130_FD_SC_LP__MUX4_4%A0 N_A0_c_626_n N_A0_M1030_g N_A0_c_627_n
+ N_A0_c_628_n N_A0_M1019_g A0 N_A0_c_630_n N_A0_c_631_n
+ PM_SKY130_FD_SC_LP__MUX4_4%A0
x_PM_SKY130_FD_SC_LP__MUX4_4%A3 N_A3_M1025_g N_A3_M1012_g A3 N_A3_c_670_n
+ PM_SKY130_FD_SC_LP__MUX4_4%A3
x_PM_SKY130_FD_SC_LP__MUX4_4%A2 N_A2_M1028_g N_A2_M1003_g A2 A2 A2 A2
+ N_A2_c_706_n N_A2_c_707_n PM_SKY130_FD_SC_LP__MUX4_4%A2
x_PM_SKY130_FD_SC_LP__MUX4_4%S0 N_S0_M1029_g N_S0_c_751_n N_S0_c_752_n
+ N_S0_M1020_g N_S0_c_762_n N_S0_c_763_n N_S0_M1017_g N_S0_c_754_n N_S0_M1010_g
+ N_S0_c_765_n N_S0_c_755_n N_S0_M1026_g N_S0_M1021_g N_S0_c_757_n N_S0_c_767_n
+ N_S0_c_758_n S0 S0 S0 S0 N_S0_c_760_n PM_SKY130_FD_SC_LP__MUX4_4%S0
x_PM_SKY130_FD_SC_LP__MUX4_4%A_27_119# N_A_27_119#_M1008_s N_A_27_119#_M1017_d
+ N_A_27_119#_M1031_s N_A_27_119#_M1013_d N_A_27_119#_c_860_n
+ N_A_27_119#_c_870_n N_A_27_119#_c_909_n N_A_27_119#_c_861_n
+ N_A_27_119#_c_862_n N_A_27_119#_c_916_n N_A_27_119#_c_863_n
+ N_A_27_119#_c_871_n N_A_27_119#_c_864_n N_A_27_119#_c_865_n
+ N_A_27_119#_c_866_n N_A_27_119#_c_867_n N_A_27_119#_c_868_n
+ PM_SKY130_FD_SC_LP__MUX4_4%A_27_119#
x_PM_SKY130_FD_SC_LP__MUX4_4%A_200_119# N_A_200_119#_M1006_d
+ N_A_200_119#_M1029_d N_A_200_119#_M1009_d N_A_200_119#_M1000_d
+ N_A_200_119#_c_1027_n N_A_200_119#_c_1025_n N_A_200_119#_c_1029_n
+ N_A_200_119#_c_1056_n N_A_200_119#_c_1030_n N_A_200_119#_c_1058_n
+ N_A_200_119#_c_1026_n N_A_200_119#_c_1069_n N_A_200_119#_c_1070_n
+ N_A_200_119#_c_1076_n N_A_200_119#_c_1071_n N_A_200_119#_c_1032_n
+ PM_SKY130_FD_SC_LP__MUX4_4%A_200_119#
x_PM_SKY130_FD_SC_LP__MUX4_4%VPWR N_VPWR_M1016_d N_VPWR_M1011_d N_VPWR_M1022_d
+ N_VPWR_M1019_d N_VPWR_M1003_d N_VPWR_c_1128_n N_VPWR_c_1129_n N_VPWR_c_1130_n
+ N_VPWR_c_1131_n N_VPWR_c_1132_n N_VPWR_c_1133_n N_VPWR_c_1134_n
+ N_VPWR_c_1135_n N_VPWR_c_1136_n N_VPWR_c_1137_n N_VPWR_c_1138_n VPWR
+ N_VPWR_c_1139_n N_VPWR_c_1140_n N_VPWR_c_1141_n N_VPWR_c_1127_n
+ N_VPWR_c_1143_n N_VPWR_c_1144_n PM_SKY130_FD_SC_LP__MUX4_4%VPWR
x_PM_SKY130_FD_SC_LP__MUX4_4%X N_X_M1014_d N_X_M1024_d N_X_M1005_s N_X_M1018_s
+ N_X_c_1231_n N_X_c_1240_n N_X_c_1241_n N_X_c_1245_n N_X_c_1263_n X X
+ N_X_c_1233_n X PM_SKY130_FD_SC_LP__MUX4_4%X
x_PM_SKY130_FD_SC_LP__MUX4_4%VGND N_VGND_M1007_d N_VGND_M1015_s N_VGND_M1027_s
+ N_VGND_M1030_d N_VGND_M1028_d N_VGND_c_1291_n N_VGND_c_1292_n N_VGND_c_1293_n
+ N_VGND_c_1294_n N_VGND_c_1295_n N_VGND_c_1296_n N_VGND_c_1297_n
+ N_VGND_c_1298_n N_VGND_c_1299_n N_VGND_c_1300_n N_VGND_c_1301_n VGND
+ N_VGND_c_1302_n N_VGND_c_1303_n N_VGND_c_1304_n N_VGND_c_1305_n
+ N_VGND_c_1306_n N_VGND_c_1307_n PM_SKY130_FD_SC_LP__MUX4_4%VGND
cc_1 VNB N_A_84_277#_M1031_g 0.00694864f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.33
cc_2 VNB N_A_84_277#_c_177_n 0.020756f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.46
cc_3 VNB N_A_84_277#_c_178_n 0.00889375f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.46
cc_4 VNB N_A_84_277#_M1006_g 0.0320005f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.805
cc_5 VNB N_A_84_277#_c_180_n 0.0187927f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.46
cc_6 VNB N_A_84_277#_c_181_n 0.00577252f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.46
cc_7 VNB N_A_84_277#_c_182_n 0.00848481f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.315
cc_8 VNB N_A_84_277#_c_183_n 0.0401213f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.315
cc_9 VNB N_A_84_277#_c_184_n 0.00360773f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.15
cc_10 VNB N_A_84_277#_c_185_n 0.00789037f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.805
cc_11 VNB N_S1_M1008_g 0.0363355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_S1_c_233_n 0.114665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_S1_c_234_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_S1_M1007_g 0.0354764f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.46
cc_15 VNB S1 4.74806e-19 $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.82
cc_16 VNB N_S1_c_237_n 0.0288418f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.315
cc_17 VNB N_A_114_119#_c_301_n 0.0176359f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.46
cc_18 VNB N_A_114_119#_c_302_n 0.0161943f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.46
cc_19 VNB N_A_114_119#_c_303_n 0.016172f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.15
cc_20 VNB N_A_114_119#_c_304_n 0.0194272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_114_119#_c_305_n 0.011932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_114_119#_c_306_n 0.024261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_114_119#_c_307_n 0.0039519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_114_119#_c_308_n 0.00140392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_114_119#_c_309_n 0.00190841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_114_119#_c_310_n 0.0020659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_114_119#_c_311_n 0.0767775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_M1001_g 0.0203487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A1_M1004_g 0.00375278f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.535
cc_30 VNB A1 0.00259188f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.33
cc_31 VNB N_A1_c_439_n 0.0434495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1041_333#_M1002_g 0.0335322f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.385
cc_33 VNB N_A_1041_333#_c_482_n 0.00572514f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.15
cc_34 VNB N_A_1041_333#_c_483_n 0.0144119f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.315
cc_35 VNB N_A_1041_333#_c_484_n 0.0295651f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.15
cc_36 VNB N_A_1041_333#_c_485_n 0.00688416f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.82
cc_37 VNB N_A_1041_333#_c_486_n 0.0272953f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.805
cc_38 VNB N_A_1041_333#_c_487_n 0.0295282f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.315
cc_39 VNB N_A_1041_333#_c_488_n 0.00431647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1041_333#_c_489_n 0.0376813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1041_333#_c_490_n 0.00117897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1041_333#_c_491_n 0.0186837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1041_333#_c_492_n 0.0202836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A0_c_626_n 0.0180176f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=0.655
cc_45 VNB N_A0_c_627_n 0.024763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A0_c_628_n 0.00804771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB A0 0.00130524f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.46
cc_48 VNB N_A0_c_630_n 0.00922834f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.805
cc_49 VNB N_A0_c_631_n 0.017978f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.46
cc_50 VNB N_A3_M1025_g 0.0463279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB A3 9.74971e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.33
cc_52 VNB N_A3_c_670_n 0.00973515f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.46
cc_53 VNB N_A2_M1028_g 0.0399096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A2_c_706_n 0.0249034f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.46
cc_55 VNB N_A2_c_707_n 0.00374129f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.82
cc_56 VNB N_S0_M1029_g 0.0355228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_S0_c_751_n 0.138765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_S0_c_752_n 0.0125859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_S0_M1017_g 0.0385379f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.805
cc_60 VNB N_S0_c_754_n 0.156353f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.46
cc_61 VNB N_S0_c_755_n 0.0234592f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.315
cc_62 VNB N_S0_M1021_g 0.0338004f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.805
cc_63 VNB N_S0_c_757_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_S0_c_758_n 0.00725219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB S0 0.00987272f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.46
cc_66 VNB N_S0_c_760_n 0.0333201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_27_119#_c_860_n 0.00230212f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.805
cc_68 VNB N_A_27_119#_c_861_n 0.00478163f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.46
cc_69 VNB N_A_27_119#_c_862_n 0.00646844f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.46
cc_70 VNB N_A_27_119#_c_863_n 0.00201292f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.97
cc_71 VNB N_A_27_119#_c_864_n 0.0269475f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.82
cc_72 VNB N_A_27_119#_c_865_n 0.0122483f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.805
cc_73 VNB N_A_27_119#_c_866_n 0.0365234f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.805
cc_74 VNB N_A_27_119#_c_867_n 0.00202061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_27_119#_c_868_n 0.00357604f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.46
cc_76 VNB N_A_200_119#_c_1025_n 0.00884369f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=0.805
cc_77 VNB N_A_200_119#_c_1026_n 0.00628681f $X=-0.19 $Y=-0.245 $X2=1.66
+ $Y2=1.315
cc_78 VNB N_VPWR_c_1127_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB X 0.00303781f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.15
cc_80 VNB N_VGND_c_1291_n 0.00429877f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.46
cc_81 VNB N_VGND_c_1292_n 0.00385266f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.105
cc_82 VNB N_VGND_c_1293_n 0.00441053f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.315
cc_83 VNB N_VGND_c_1294_n 0.0202243f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.82
cc_84 VNB N_VGND_c_1295_n 0.0151289f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.805
cc_85 VNB N_VGND_c_1296_n 0.0190273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1297_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.46
cc_87 VNB N_VGND_c_1298_n 0.0190273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1299_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1300_n 0.0497514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1301_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1302_n 0.0666225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1303_n 0.0446284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1304_n 0.0381228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1305_n 0.459108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1306_n 0.00362723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1307_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VPB N_A_84_277#_M1031_g 0.0356888f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.33
cc_98 VPB N_A_84_277#_c_187_n 0.00388057f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.105
cc_99 VPB N_A_84_277#_c_182_n 0.00356164f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.315
cc_100 VPB N_A_84_277#_c_183_n 0.0255524f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.315
cc_101 VPB N_S1_c_238_n 0.0190925f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.535
cc_102 VPB N_S1_c_239_n 0.0759956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_S1_c_240_n 0.0143744f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.46
cc_104 VPB N_S1_M1016_g 0.042298f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.805
cc_105 VPB S1 0.00290737f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.82
cc_106 VPB N_S1_c_237_n 0.0103336f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.315
cc_107 VPB N_A_114_119#_M1005_g 0.0209612f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.33
cc_108 VPB N_A_114_119#_M1011_g 0.0177998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_114_119#_M1018_g 0.0177858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_114_119#_M1022_g 0.0203677f $X=-0.19 $Y=1.655 $X2=1.66 $Y2=1.82
cc_111 VPB N_A_114_119#_c_305_n 0.00994035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_114_119#_c_311_n 0.0114889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A1_M1004_g 0.0445876f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.535
cc_114 VPB A1 0.00209787f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.33
cc_115 VPB N_A1_c_439_n 0.014869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_1041_333#_M1000_g 0.029607f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.33
cc_117 VPB N_A_1041_333#_M1013_g 0.0273045f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.46
cc_118 VPB N_A_1041_333#_c_482_n 0.0249169f $X=-0.19 $Y=1.655 $X2=1.81 $Y2=1.15
cc_119 VPB N_A_1041_333#_c_485_n 0.00535874f $X=-0.19 $Y=1.655 $X2=1.66 $Y2=1.82
cc_120 VPB N_A_1041_333#_c_497_n 0.00293684f $X=-0.19 $Y=1.655 $X2=1.94
+ $Y2=0.805
cc_121 VPB N_A_1041_333#_c_488_n 0.00225584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_1041_333#_c_499_n 0.00429647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_1041_333#_c_500_n 0.00305622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_1041_333#_c_501_n 0.0242653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_1041_333#_c_489_n 0.0161157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_1041_333#_c_492_n 0.0339554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A0_M1019_g 0.0249593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB A0 0.00243862f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.46
cc_129 VPB N_A0_c_630_n 0.0238822f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.805
cc_130 VPB N_A3_M1012_g 0.0213038f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.535
cc_131 VPB A3 0.00264979f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.33
cc_132 VPB N_A3_c_670_n 0.0203965f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.46
cc_133 VPB N_A2_M1003_g 0.023951f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.535
cc_134 VPB N_A2_c_706_n 0.021132f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.46
cc_135 VPB N_A2_c_707_n 0.0099597f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.82
cc_136 VPB N_S0_M1020_g 0.0304842f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.33
cc_137 VPB N_S0_c_762_n 0.160008f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.46
cc_138 VPB N_S0_c_763_n 0.012806f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.46
cc_139 VPB N_S0_M1010_g 0.0358263f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.105
cc_140 VPB N_S0_c_765_n 0.0665969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_S0_M1026_g 0.0453462f $X=-0.19 $Y=1.655 $X2=1.66 $Y2=1.82
cc_142 VPB N_S0_c_767_n 0.00749069f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.315
cc_143 VPB N_S0_c_758_n 0.0207957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB S0 9.47981e-19 $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.46
cc_145 VPB N_A_27_119#_c_860_n 0.00791059f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.805
cc_146 VPB N_A_27_119#_c_870_n 0.0224469f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.805
cc_147 VPB N_A_27_119#_c_871_n 0.0034628f $X=-0.19 $Y=1.655 $X2=1.66 $Y2=1.15
cc_148 VPB N_A_27_119#_c_866_n 0.0209065f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=0.805
cc_149 VPB N_A_200_119#_c_1027_n 0.00297297f $X=-0.19 $Y=1.655 $X2=0.925
+ $Y2=1.385
cc_150 VPB N_A_200_119#_c_1025_n 0.00811073f $X=-0.19 $Y=1.655 $X2=0.925
+ $Y2=0.805
cc_151 VPB N_A_200_119#_c_1029_n 0.0288089f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.46
cc_152 VPB N_A_200_119#_c_1030_n 0.00197915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_200_119#_c_1026_n 0.00204419f $X=-0.19 $Y=1.655 $X2=1.66
+ $Y2=1.315
cc_154 VPB N_A_200_119#_c_1032_n 9.7648e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_1128_n 0.013716f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.46
cc_156 VPB N_VPWR_c_1129_n 0.00434709f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.105
cc_157 VPB N_VPWR_c_1130_n 0.0176046f $X=-0.19 $Y=1.655 $X2=1.66 $Y2=1.315
cc_158 VPB N_VPWR_c_1131_n 0.0133906f $X=-0.19 $Y=1.655 $X2=1.66 $Y2=1.82
cc_159 VPB N_VPWR_c_1132_n 0.00854505f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=0.805
cc_160 VPB N_VPWR_c_1133_n 0.0735785f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1134_n 0.00632207f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=1.46
cc_162 VPB N_VPWR_c_1135_n 0.016802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1136_n 0.00632207f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1137_n 0.0542918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1138_n 0.00277066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1139_n 0.0279397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1140_n 0.0444619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1141_n 0.0287137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1127_n 0.138924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1143_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1144_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_X_c_1231_n 0.00563683f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.385
cc_173 VPB X 0.00275081f $X=-0.19 $Y=1.655 $X2=1.66 $Y2=1.15
cc_174 VPB N_X_c_1233_n 0.00214215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 N_A_84_277#_c_178_n N_S1_M1008_g 0.0111069f $X=0.57 $Y=1.46 $X2=0 $Y2=0
cc_176 N_A_84_277#_M1006_g N_S1_M1008_g 0.0135639f $X=0.925 $Y=0.805 $X2=0 $Y2=0
cc_177 N_A_84_277#_M1006_g N_S1_c_233_n 0.00881852f $X=0.925 $Y=0.805 $X2=0
+ $Y2=0
cc_178 N_A_84_277#_M1031_g N_S1_c_238_n 0.0110475f $X=0.495 $Y=2.33 $X2=0 $Y2=0
cc_179 N_A_84_277#_c_181_n N_S1_c_238_n 0.00799915f $X=0.925 $Y=1.46 $X2=0 $Y2=0
cc_180 N_A_84_277#_c_187_n N_S1_M1016_g 0.00254128f $X=1.73 $Y=2.105 $X2=0 $Y2=0
cc_181 N_A_84_277#_c_182_n N_S1_M1016_g 0.00340825f $X=1.51 $Y=1.315 $X2=0 $Y2=0
cc_182 N_A_84_277#_c_183_n N_S1_M1016_g 0.00814743f $X=1.51 $Y=1.315 $X2=0 $Y2=0
cc_183 N_A_84_277#_c_183_n N_S1_M1007_g 7.81725e-19 $X=1.51 $Y=1.315 $X2=0 $Y2=0
cc_184 N_A_84_277#_c_184_n N_S1_M1007_g 0.00585945f $X=1.66 $Y=1.15 $X2=0 $Y2=0
cc_185 N_A_84_277#_c_185_n N_S1_M1007_g 0.00130816f $X=1.94 $Y=0.805 $X2=0 $Y2=0
cc_186 N_A_84_277#_c_182_n S1 0.054458f $X=1.51 $Y=1.315 $X2=0 $Y2=0
cc_187 N_A_84_277#_c_183_n S1 7.00019e-19 $X=1.51 $Y=1.315 $X2=0 $Y2=0
cc_188 N_A_84_277#_c_182_n N_S1_c_237_n 0.00281599f $X=1.51 $Y=1.315 $X2=0 $Y2=0
cc_189 N_A_84_277#_c_183_n N_S1_c_237_n 0.0117264f $X=1.51 $Y=1.315 $X2=0 $Y2=0
cc_190 N_A_84_277#_c_185_n N_S1_c_237_n 0.00115542f $X=1.94 $Y=0.805 $X2=0 $Y2=0
cc_191 N_A_84_277#_M1031_g N_A_114_119#_c_305_n 0.00931102f $X=0.495 $Y=2.33
+ $X2=0 $Y2=0
cc_192 N_A_84_277#_c_177_n N_A_114_119#_c_305_n 0.0147082f $X=0.85 $Y=1.46 $X2=0
+ $Y2=0
cc_193 N_A_84_277#_M1006_g N_A_114_119#_c_305_n 0.00989317f $X=0.925 $Y=0.805
+ $X2=0 $Y2=0
cc_194 N_A_84_277#_M1006_g N_A_114_119#_c_306_n 0.00389216f $X=0.925 $Y=0.805
+ $X2=0 $Y2=0
cc_195 N_A_84_277#_c_183_n N_A_114_119#_c_306_n 0.00489041f $X=1.51 $Y=1.315
+ $X2=0 $Y2=0
cc_196 N_A_84_277#_c_185_n N_A_114_119#_c_306_n 0.0172575f $X=1.94 $Y=0.805
+ $X2=0 $Y2=0
cc_197 N_A_84_277#_c_185_n N_A_114_119#_c_308_n 0.0136852f $X=1.94 $Y=0.805
+ $X2=0 $Y2=0
cc_198 N_A_84_277#_c_184_n N_A_114_119#_c_325_n 0.00170694f $X=1.66 $Y=1.15
+ $X2=0 $Y2=0
cc_199 N_A_84_277#_c_185_n N_A_114_119#_c_325_n 0.0104097f $X=1.94 $Y=0.805
+ $X2=0 $Y2=0
cc_200 N_A_84_277#_M1006_g N_A_27_119#_c_864_n 0.00988487f $X=0.925 $Y=0.805
+ $X2=0 $Y2=0
cc_201 N_A_84_277#_c_182_n N_A_27_119#_c_864_n 0.010236f $X=1.51 $Y=1.315 $X2=0
+ $Y2=0
cc_202 N_A_84_277#_c_183_n N_A_27_119#_c_864_n 0.0018075f $X=1.51 $Y=1.315 $X2=0
+ $Y2=0
cc_203 N_A_84_277#_c_185_n N_A_27_119#_c_864_n 0.00928745f $X=1.94 $Y=0.805
+ $X2=0 $Y2=0
cc_204 N_A_84_277#_c_178_n N_A_27_119#_c_866_n 0.0159017f $X=0.57 $Y=1.46 $X2=0
+ $Y2=0
cc_205 N_A_84_277#_M1006_g N_A_200_119#_c_1025_n 0.00570008f $X=0.925 $Y=0.805
+ $X2=0 $Y2=0
cc_206 N_A_84_277#_c_180_n N_A_200_119#_c_1025_n 0.0163389f $X=1.345 $Y=1.46
+ $X2=0 $Y2=0
cc_207 N_A_84_277#_c_187_n N_A_200_119#_c_1025_n 0.0189198f $X=1.73 $Y=2.105
+ $X2=0 $Y2=0
cc_208 N_A_84_277#_c_182_n N_A_200_119#_c_1025_n 0.0497699f $X=1.51 $Y=1.315
+ $X2=0 $Y2=0
cc_209 N_A_84_277#_c_183_n N_A_200_119#_c_1025_n 0.00897112f $X=1.51 $Y=1.315
+ $X2=0 $Y2=0
cc_210 N_A_84_277#_c_184_n N_A_200_119#_c_1025_n 0.00663173f $X=1.66 $Y=1.15
+ $X2=0 $Y2=0
cc_211 N_A_84_277#_c_185_n N_A_200_119#_c_1025_n 0.0122994f $X=1.94 $Y=0.805
+ $X2=0 $Y2=0
cc_212 N_A_84_277#_c_187_n N_A_200_119#_c_1029_n 0.0260475f $X=1.73 $Y=2.105
+ $X2=0 $Y2=0
cc_213 N_A_84_277#_c_182_n N_A_200_119#_c_1029_n 0.00454075f $X=1.51 $Y=1.315
+ $X2=0 $Y2=0
cc_214 N_A_84_277#_c_183_n N_A_200_119#_c_1029_n 0.00332828f $X=1.51 $Y=1.315
+ $X2=0 $Y2=0
cc_215 N_A_84_277#_M1031_g N_VPWR_c_1133_n 0.0038748f $X=0.495 $Y=2.33 $X2=0
+ $Y2=0
cc_216 N_A_84_277#_M1031_g N_VPWR_c_1127_n 0.00454494f $X=0.495 $Y=2.33 $X2=0
+ $Y2=0
cc_217 N_S1_M1016_g N_A_114_119#_M1005_g 0.0373197f $X=2.16 $Y=1.995 $X2=0 $Y2=0
cc_218 S1 N_A_114_119#_M1005_g 0.00376812f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_219 N_S1_c_233_n N_A_114_119#_c_301_n 0.0164326f $X=2.1 $Y=0.18 $X2=0 $Y2=0
cc_220 N_S1_M1008_g N_A_114_119#_c_305_n 0.00272799f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_221 N_S1_c_238_n N_A_114_119#_c_305_n 0.00112621f $X=0.925 $Y=2.76 $X2=0
+ $Y2=0
cc_222 N_S1_c_233_n N_A_114_119#_c_306_n 0.0255354f $X=2.1 $Y=0.18 $X2=0 $Y2=0
cc_223 N_S1_M1007_g N_A_114_119#_c_306_n 0.0113462f $X=2.175 $Y=0.865 $X2=0
+ $Y2=0
cc_224 N_S1_M1008_g N_A_114_119#_c_307_n 0.008099f $X=0.495 $Y=0.805 $X2=0 $Y2=0
cc_225 N_S1_c_233_n N_A_114_119#_c_307_n 0.00329158f $X=2.1 $Y=0.18 $X2=0 $Y2=0
cc_226 N_S1_M1007_g N_A_114_119#_c_308_n 0.0115179f $X=2.175 $Y=0.865 $X2=0
+ $Y2=0
cc_227 N_S1_M1007_g N_A_114_119#_c_325_n 0.00617678f $X=2.175 $Y=0.865 $X2=0
+ $Y2=0
cc_228 S1 N_A_114_119#_c_325_n 0.00306186f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_229 N_S1_c_237_n N_A_114_119#_c_325_n 0.00193244f $X=2.16 $Y=1.35 $X2=0 $Y2=0
cc_230 N_S1_M1007_g N_A_114_119#_c_309_n 0.00324945f $X=2.175 $Y=0.865 $X2=0
+ $Y2=0
cc_231 S1 N_A_114_119#_c_309_n 0.00318627f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_232 N_S1_c_237_n N_A_114_119#_c_309_n 5.52573e-19 $X=2.16 $Y=1.35 $X2=0 $Y2=0
cc_233 S1 N_A_114_119#_c_310_n 0.00770634f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_234 N_S1_c_237_n N_A_114_119#_c_310_n 0.0014175f $X=2.16 $Y=1.35 $X2=0 $Y2=0
cc_235 S1 N_A_114_119#_c_311_n 7.88151e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_236 N_S1_c_237_n N_A_114_119#_c_311_n 0.0138371f $X=2.16 $Y=1.35 $X2=0 $Y2=0
cc_237 N_S1_M1008_g N_A_27_119#_c_864_n 0.00905163f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_238 N_S1_M1007_g N_A_27_119#_c_864_n 0.00443064f $X=2.175 $Y=0.865 $X2=0
+ $Y2=0
cc_239 S1 N_A_27_119#_c_864_n 0.00399281f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_240 N_S1_c_237_n N_A_27_119#_c_864_n 9.79667e-19 $X=2.16 $Y=1.35 $X2=0 $Y2=0
cc_241 N_S1_M1008_g N_A_27_119#_c_865_n 0.00116153f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_242 N_S1_M1008_g N_A_27_119#_c_866_n 0.00717262f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_243 N_S1_c_238_n N_A_200_119#_c_1027_n 6.41154e-19 $X=0.925 $Y=2.76 $X2=0
+ $Y2=0
cc_244 N_S1_c_239_n N_A_200_119#_c_1027_n 0.00443957f $X=2.085 $Y=2.835 $X2=0
+ $Y2=0
cc_245 N_S1_c_238_n N_A_200_119#_c_1025_n 0.0030815f $X=0.925 $Y=2.76 $X2=0
+ $Y2=0
cc_246 N_S1_c_239_n N_A_200_119#_c_1029_n 0.0243162f $X=2.085 $Y=2.835 $X2=0
+ $Y2=0
cc_247 N_S1_M1016_g N_A_200_119#_c_1029_n 0.014667f $X=2.16 $Y=1.995 $X2=0 $Y2=0
cc_248 S1 N_A_200_119#_c_1029_n 0.00890299f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_249 N_S1_M1016_g N_VPWR_c_1128_n 0.00538712f $X=2.16 $Y=1.995 $X2=0 $Y2=0
cc_250 N_S1_c_240_n N_VPWR_c_1133_n 0.0351973f $X=1 $Y=2.835 $X2=0 $Y2=0
cc_251 N_S1_c_240_n N_VPWR_c_1127_n 0.0392491f $X=1 $Y=2.835 $X2=0 $Y2=0
cc_252 S1 N_X_c_1231_n 0.00100849f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_253 N_S1_c_233_n N_VGND_c_1291_n 0.00299233f $X=2.1 $Y=0.18 $X2=0 $Y2=0
cc_254 N_S1_M1007_g N_VGND_c_1291_n 7.0505e-19 $X=2.175 $Y=0.865 $X2=0 $Y2=0
cc_255 N_S1_c_234_n N_VGND_c_1302_n 0.0421819f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_256 N_S1_c_233_n N_VGND_c_1305_n 0.0336876f $X=2.1 $Y=0.18 $X2=0 $Y2=0
cc_257 N_S1_c_234_n N_VGND_c_1305_n 0.00589026f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_258 N_A_114_119#_c_304_n N_A1_M1001_g 0.0137144f $X=4.145 $Y=1.185 $X2=0
+ $Y2=0
cc_259 N_A_114_119#_M1022_g A1 0.00115418f $X=3.995 $Y=2.305 $X2=0 $Y2=0
cc_260 N_A_114_119#_c_311_n A1 8.03683e-19 $X=3.995 $Y=1.35 $X2=0 $Y2=0
cc_261 N_A_114_119#_c_311_n N_A1_c_439_n 0.0163462f $X=3.995 $Y=1.35 $X2=0 $Y2=0
cc_262 N_A_114_119#_M1008_d N_A_27_119#_c_864_n 0.003271f $X=0.57 $Y=0.595 $X2=0
+ $Y2=0
cc_263 N_A_114_119#_c_301_n N_A_27_119#_c_864_n 0.0077552f $X=2.855 $Y=1.185
+ $X2=0 $Y2=0
cc_264 N_A_114_119#_c_302_n N_A_27_119#_c_864_n 0.0030285f $X=3.285 $Y=1.185
+ $X2=0 $Y2=0
cc_265 N_A_114_119#_c_303_n N_A_27_119#_c_864_n 0.0030285f $X=3.715 $Y=1.185
+ $X2=0 $Y2=0
cc_266 N_A_114_119#_c_304_n N_A_27_119#_c_864_n 0.00489944f $X=4.145 $Y=1.185
+ $X2=0 $Y2=0
cc_267 N_A_114_119#_c_305_n N_A_27_119#_c_864_n 0.0220735f $X=0.71 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_114_119#_c_306_n N_A_27_119#_c_864_n 0.0328529f $X=2.205 $Y=0.375
+ $X2=0 $Y2=0
cc_269 N_A_114_119#_c_308_n N_A_27_119#_c_864_n 0.0163939f $X=2.29 $Y=0.835
+ $X2=0 $Y2=0
cc_270 N_A_114_119#_c_359_p N_A_27_119#_c_864_n 0.0148929f $X=2.615 $Y=0.92
+ $X2=0 $Y2=0
cc_271 N_A_114_119#_c_305_n N_A_27_119#_c_865_n 0.00213704f $X=0.71 $Y=0.74
+ $X2=0 $Y2=0
cc_272 N_A_114_119#_c_307_n N_A_27_119#_c_865_n 0.00106697f $X=0.795 $Y=0.375
+ $X2=0 $Y2=0
cc_273 N_A_114_119#_c_305_n N_A_27_119#_c_866_n 0.0677075f $X=0.71 $Y=0.74 $X2=0
+ $Y2=0
cc_274 N_A_114_119#_c_305_n N_A_200_119#_c_1027_n 5.47165e-19 $X=0.71 $Y=0.74
+ $X2=0 $Y2=0
cc_275 N_A_114_119#_c_305_n N_A_200_119#_c_1025_n 0.0590108f $X=0.71 $Y=0.74
+ $X2=0 $Y2=0
cc_276 N_A_114_119#_c_306_n N_A_200_119#_c_1025_n 0.0118084f $X=2.205 $Y=0.375
+ $X2=0 $Y2=0
cc_277 N_A_114_119#_M1005_g N_A_200_119#_c_1029_n 0.0166576f $X=2.705 $Y=2.305
+ $X2=0 $Y2=0
cc_278 N_A_114_119#_M1011_g N_A_200_119#_c_1029_n 0.0126945f $X=3.135 $Y=2.305
+ $X2=0 $Y2=0
cc_279 N_A_114_119#_M1018_g N_A_200_119#_c_1029_n 0.0126479f $X=3.565 $Y=2.305
+ $X2=0 $Y2=0
cc_280 N_A_114_119#_M1022_g N_A_200_119#_c_1029_n 0.0138794f $X=3.995 $Y=2.305
+ $X2=0 $Y2=0
cc_281 N_A_114_119#_M1018_g N_A_200_119#_c_1056_n 0.00100351f $X=3.565 $Y=2.305
+ $X2=0 $Y2=0
cc_282 N_A_114_119#_M1022_g N_A_200_119#_c_1056_n 0.00698234f $X=3.995 $Y=2.305
+ $X2=0 $Y2=0
cc_283 N_A_114_119#_M1018_g N_A_200_119#_c_1058_n 7.78212e-19 $X=3.565 $Y=2.305
+ $X2=0 $Y2=0
cc_284 N_A_114_119#_M1022_g N_A_200_119#_c_1058_n 0.00784118f $X=3.995 $Y=2.305
+ $X2=0 $Y2=0
cc_285 N_A_114_119#_c_311_n N_A_200_119#_c_1058_n 0.00163843f $X=3.995 $Y=1.35
+ $X2=0 $Y2=0
cc_286 N_A_114_119#_M1005_g N_VPWR_c_1128_n 0.00939796f $X=2.705 $Y=2.305 $X2=0
+ $Y2=0
cc_287 N_A_114_119#_M1011_g N_VPWR_c_1128_n 0.0010009f $X=3.135 $Y=2.305 $X2=0
+ $Y2=0
cc_288 N_A_114_119#_M1005_g N_VPWR_c_1129_n 0.0010009f $X=2.705 $Y=2.305 $X2=0
+ $Y2=0
cc_289 N_A_114_119#_M1011_g N_VPWR_c_1129_n 0.00833447f $X=3.135 $Y=2.305 $X2=0
+ $Y2=0
cc_290 N_A_114_119#_M1018_g N_VPWR_c_1129_n 0.00861369f $X=3.565 $Y=2.305 $X2=0
+ $Y2=0
cc_291 N_A_114_119#_M1022_g N_VPWR_c_1129_n 0.00165793f $X=3.995 $Y=2.305 $X2=0
+ $Y2=0
cc_292 N_A_114_119#_M1022_g N_VPWR_c_1130_n 0.0175462f $X=3.995 $Y=2.305 $X2=0
+ $Y2=0
cc_293 N_A_114_119#_c_305_n N_VPWR_c_1133_n 0.00354692f $X=0.71 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_114_119#_M1005_g N_VPWR_c_1135_n 0.00465077f $X=2.705 $Y=2.305 $X2=0
+ $Y2=0
cc_295 N_A_114_119#_M1011_g N_VPWR_c_1135_n 0.00465077f $X=3.135 $Y=2.305 $X2=0
+ $Y2=0
cc_296 N_A_114_119#_M1018_g N_VPWR_c_1139_n 0.00465077f $X=3.565 $Y=2.305 $X2=0
+ $Y2=0
cc_297 N_A_114_119#_M1022_g N_VPWR_c_1139_n 0.00559701f $X=3.995 $Y=2.305 $X2=0
+ $Y2=0
cc_298 N_A_114_119#_M1005_g N_VPWR_c_1127_n 0.00451796f $X=2.705 $Y=2.305 $X2=0
+ $Y2=0
cc_299 N_A_114_119#_M1011_g N_VPWR_c_1127_n 0.00451796f $X=3.135 $Y=2.305 $X2=0
+ $Y2=0
cc_300 N_A_114_119#_M1018_g N_VPWR_c_1127_n 0.00451796f $X=3.565 $Y=2.305 $X2=0
+ $Y2=0
cc_301 N_A_114_119#_M1022_g N_VPWR_c_1127_n 0.00537853f $X=3.995 $Y=2.305 $X2=0
+ $Y2=0
cc_302 N_A_114_119#_c_305_n N_VPWR_c_1127_n 0.00555956f $X=0.71 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_A_114_119#_M1005_g N_X_c_1231_n 4.44852e-19 $X=2.705 $Y=2.305 $X2=0
+ $Y2=0
cc_304 N_A_114_119#_M1011_g N_X_c_1231_n 0.0146578f $X=3.135 $Y=2.305 $X2=0
+ $Y2=0
cc_305 N_A_114_119#_M1018_g N_X_c_1231_n 0.0146729f $X=3.565 $Y=2.305 $X2=0
+ $Y2=0
cc_306 N_A_114_119#_c_395_p N_X_c_1231_n 0.05209f $X=3.475 $Y=1.35 $X2=0 $Y2=0
cc_307 N_A_114_119#_c_311_n N_X_c_1231_n 0.00572418f $X=3.995 $Y=1.35 $X2=0
+ $Y2=0
cc_308 N_A_114_119#_c_308_n N_X_c_1240_n 0.00409765f $X=2.29 $Y=0.835 $X2=0
+ $Y2=0
cc_309 N_A_114_119#_c_302_n N_X_c_1241_n 0.00922533f $X=3.285 $Y=1.185 $X2=0
+ $Y2=0
cc_310 N_A_114_119#_c_303_n N_X_c_1241_n 0.0107007f $X=3.715 $Y=1.185 $X2=0
+ $Y2=0
cc_311 N_A_114_119#_c_395_p N_X_c_1241_n 0.0208115f $X=3.475 $Y=1.35 $X2=0 $Y2=0
cc_312 N_A_114_119#_c_311_n N_X_c_1241_n 0.00275994f $X=3.995 $Y=1.35 $X2=0
+ $Y2=0
cc_313 N_A_114_119#_c_395_p N_X_c_1245_n 0.0113592f $X=3.475 $Y=1.35 $X2=0 $Y2=0
cc_314 N_A_114_119#_c_311_n N_X_c_1245_n 0.00287453f $X=3.995 $Y=1.35 $X2=0
+ $Y2=0
cc_315 N_A_114_119#_M1018_g X 0.00279028f $X=3.565 $Y=2.305 $X2=0 $Y2=0
cc_316 N_A_114_119#_c_303_n X 0.00346214f $X=3.715 $Y=1.185 $X2=0 $Y2=0
cc_317 N_A_114_119#_M1022_g X 0.00431048f $X=3.995 $Y=2.305 $X2=0 $Y2=0
cc_318 N_A_114_119#_c_304_n X 0.00273439f $X=4.145 $Y=1.185 $X2=0 $Y2=0
cc_319 N_A_114_119#_c_395_p X 0.010603f $X=3.475 $Y=1.35 $X2=0 $Y2=0
cc_320 N_A_114_119#_c_311_n X 0.0285917f $X=3.995 $Y=1.35 $X2=0 $Y2=0
cc_321 N_A_114_119#_M1022_g N_X_c_1233_n 0.00930382f $X=3.995 $Y=2.305 $X2=0
+ $Y2=0
cc_322 N_A_114_119#_c_311_n N_X_c_1233_n 0.00337022f $X=3.995 $Y=1.35 $X2=0
+ $Y2=0
cc_323 N_A_114_119#_c_308_n N_VGND_M1007_d 0.00281436f $X=2.29 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_324 N_A_114_119#_c_359_p N_VGND_M1007_d 0.0151679f $X=2.615 $Y=0.92 $X2=-0.19
+ $Y2=-0.245
cc_325 N_A_114_119#_c_325_n N_VGND_M1007_d 0.00247357f $X=2.375 $Y=0.92
+ $X2=-0.19 $Y2=-0.245
cc_326 N_A_114_119#_c_309_n N_VGND_M1007_d 9.40899e-19 $X=2.7 $Y=1.265 $X2=-0.19
+ $Y2=-0.245
cc_327 N_A_114_119#_c_301_n N_VGND_c_1291_n 0.00199501f $X=2.855 $Y=1.185 $X2=0
+ $Y2=0
cc_328 N_A_114_119#_c_306_n N_VGND_c_1291_n 0.0136568f $X=2.205 $Y=0.375 $X2=0
+ $Y2=0
cc_329 N_A_114_119#_c_308_n N_VGND_c_1291_n 0.00570278f $X=2.29 $Y=0.835 $X2=0
+ $Y2=0
cc_330 N_A_114_119#_c_359_p N_VGND_c_1291_n 0.00661924f $X=2.615 $Y=0.92 $X2=0
+ $Y2=0
cc_331 N_A_114_119#_c_311_n N_VGND_c_1291_n 3.07899e-19 $X=3.995 $Y=1.35 $X2=0
+ $Y2=0
cc_332 N_A_114_119#_c_302_n N_VGND_c_1292_n 0.0016604f $X=3.285 $Y=1.185 $X2=0
+ $Y2=0
cc_333 N_A_114_119#_c_303_n N_VGND_c_1292_n 0.0016604f $X=3.715 $Y=1.185 $X2=0
+ $Y2=0
cc_334 N_A_114_119#_c_304_n N_VGND_c_1293_n 0.00351171f $X=4.145 $Y=1.185 $X2=0
+ $Y2=0
cc_335 N_A_114_119#_c_301_n N_VGND_c_1296_n 0.00585385f $X=2.855 $Y=1.185 $X2=0
+ $Y2=0
cc_336 N_A_114_119#_c_302_n N_VGND_c_1296_n 0.00585385f $X=3.285 $Y=1.185 $X2=0
+ $Y2=0
cc_337 N_A_114_119#_c_303_n N_VGND_c_1298_n 0.00585385f $X=3.715 $Y=1.185 $X2=0
+ $Y2=0
cc_338 N_A_114_119#_c_304_n N_VGND_c_1298_n 0.00585385f $X=4.145 $Y=1.185 $X2=0
+ $Y2=0
cc_339 N_A_114_119#_c_306_n N_VGND_c_1302_n 0.0840212f $X=2.205 $Y=0.375 $X2=0
+ $Y2=0
cc_340 N_A_114_119#_c_307_n N_VGND_c_1302_n 0.0111417f $X=0.795 $Y=0.375 $X2=0
+ $Y2=0
cc_341 N_A_114_119#_c_301_n N_VGND_c_1305_n 0.00594448f $X=2.855 $Y=1.185 $X2=0
+ $Y2=0
cc_342 N_A_114_119#_c_302_n N_VGND_c_1305_n 0.00516778f $X=3.285 $Y=1.185 $X2=0
+ $Y2=0
cc_343 N_A_114_119#_c_303_n N_VGND_c_1305_n 0.00516778f $X=3.715 $Y=1.185 $X2=0
+ $Y2=0
cc_344 N_A_114_119#_c_304_n N_VGND_c_1305_n 0.00677528f $X=4.145 $Y=1.185 $X2=0
+ $Y2=0
cc_345 N_A_114_119#_c_306_n N_VGND_c_1305_n 0.0159237f $X=2.205 $Y=0.375 $X2=0
+ $Y2=0
cc_346 N_A_114_119#_c_307_n N_VGND_c_1305_n 0.00215088f $X=0.795 $Y=0.375 $X2=0
+ $Y2=0
cc_347 N_A1_M1001_g N_A_1041_333#_M1002_g 0.00271217f $X=4.685 $Y=0.805 $X2=0
+ $Y2=0
cc_348 N_A1_c_439_n N_A_1041_333#_M1002_g 0.00381455f $X=4.685 $Y=1.36 $X2=0
+ $Y2=0
cc_349 N_A1_M1004_g N_A_1041_333#_c_492_n 0.0811006f $X=4.92 $Y=2.475 $X2=0
+ $Y2=0
cc_350 N_A1_M1001_g N_S0_M1029_g 0.041468f $X=4.685 $Y=0.805 $X2=0 $Y2=0
cc_351 N_A1_c_439_n N_S0_M1029_g 0.00138617f $X=4.685 $Y=1.36 $X2=0 $Y2=0
cc_352 N_A1_M1004_g N_A_27_119#_c_860_n 4.28076e-19 $X=4.92 $Y=2.475 $X2=0 $Y2=0
cc_353 N_A1_c_439_n N_A_27_119#_c_860_n 8.08842e-19 $X=4.685 $Y=1.36 $X2=0 $Y2=0
cc_354 N_A1_M1001_g N_A_27_119#_c_864_n 0.00763193f $X=4.685 $Y=0.805 $X2=0
+ $Y2=0
cc_355 A1 N_A_27_119#_c_864_n 0.00622349f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_356 N_A1_c_439_n N_A_27_119#_c_864_n 2.32902e-19 $X=4.685 $Y=1.36 $X2=0 $Y2=0
cc_357 N_A1_M1004_g N_A_200_119#_c_1056_n 0.0038421f $X=4.92 $Y=2.475 $X2=0
+ $Y2=0
cc_358 N_A1_M1004_g N_A_200_119#_c_1030_n 0.0100992f $X=4.92 $Y=2.475 $X2=0
+ $Y2=0
cc_359 A1 N_A_200_119#_c_1030_n 0.0124086f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_360 N_A1_c_439_n N_A_200_119#_c_1030_n 0.00676092f $X=4.685 $Y=1.36 $X2=0
+ $Y2=0
cc_361 N_A1_M1001_g N_A_200_119#_c_1026_n 0.0071553f $X=4.685 $Y=0.805 $X2=0
+ $Y2=0
cc_362 N_A1_M1004_g N_A_200_119#_c_1026_n 0.0169383f $X=4.92 $Y=2.475 $X2=0
+ $Y2=0
cc_363 A1 N_A_200_119#_c_1026_n 0.0325329f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_364 N_A1_c_439_n N_A_200_119#_c_1026_n 0.00650597f $X=4.685 $Y=1.36 $X2=0
+ $Y2=0
cc_365 N_A1_M1004_g N_A_200_119#_c_1069_n 0.0106307f $X=4.92 $Y=2.475 $X2=0
+ $Y2=0
cc_366 N_A1_M1004_g N_A_200_119#_c_1070_n 0.0094102f $X=4.92 $Y=2.475 $X2=0
+ $Y2=0
cc_367 N_A1_M1001_g N_A_200_119#_c_1071_n 0.0041444f $X=4.685 $Y=0.805 $X2=0
+ $Y2=0
cc_368 N_A1_M1004_g N_A_200_119#_c_1032_n 0.00208048f $X=4.92 $Y=2.475 $X2=0
+ $Y2=0
cc_369 A1 N_VPWR_M1022_d 0.0046236f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_370 N_A1_M1004_g N_VPWR_c_1130_n 0.0149132f $X=4.92 $Y=2.475 $X2=0 $Y2=0
cc_371 N_A1_M1004_g N_VPWR_c_1140_n 0.00398025f $X=4.92 $Y=2.475 $X2=0 $Y2=0
cc_372 N_A1_M1004_g N_VPWR_c_1127_n 0.00495025f $X=4.92 $Y=2.475 $X2=0 $Y2=0
cc_373 A1 X 0.0217878f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_374 N_A1_c_439_n X 0.00204325f $X=4.685 $Y=1.36 $X2=0 $Y2=0
cc_375 N_A1_M1004_g N_X_c_1233_n 0.00180697f $X=4.92 $Y=2.475 $X2=0 $Y2=0
cc_376 A1 N_X_c_1233_n 0.00565454f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_377 N_A1_M1001_g N_VGND_c_1293_n 0.00573413f $X=4.685 $Y=0.805 $X2=0 $Y2=0
cc_378 N_A1_c_439_n N_VGND_c_1293_n 0.00132312f $X=4.685 $Y=1.36 $X2=0 $Y2=0
cc_379 N_A1_M1001_g N_VGND_c_1303_n 0.00431487f $X=4.685 $Y=0.805 $X2=0 $Y2=0
cc_380 N_A1_M1001_g N_VGND_c_1305_n 0.00290123f $X=4.685 $Y=0.805 $X2=0 $Y2=0
cc_381 N_A_1041_333#_M1002_g N_A0_c_626_n 0.0513125f $X=5.475 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_382 N_A_1041_333#_c_484_n N_A0_c_627_n 0.00537366f $X=7.485 $Y=1.315 $X2=0
+ $Y2=0
cc_383 N_A_1041_333#_c_485_n N_A0_c_627_n 0.00472145f $X=6.045 $Y=1.315 $X2=0
+ $Y2=0
cc_384 N_A_1041_333#_c_485_n N_A0_c_628_n 0.00282394f $X=6.045 $Y=1.315 $X2=0
+ $Y2=0
cc_385 N_A_1041_333#_c_492_n N_A0_c_628_n 0.0063381f $X=5.475 $Y=1.65 $X2=0
+ $Y2=0
cc_386 N_A_1041_333#_c_484_n A0 0.0245868f $X=7.485 $Y=1.315 $X2=0 $Y2=0
cc_387 N_A_1041_333#_c_485_n A0 0.0183596f $X=6.045 $Y=1.315 $X2=0 $Y2=0
cc_388 N_A_1041_333#_c_484_n N_A0_c_630_n 0.00400978f $X=7.485 $Y=1.315 $X2=0
+ $Y2=0
cc_389 N_A_1041_333#_M1002_g N_A0_c_631_n 0.00265335f $X=5.475 $Y=0.805 $X2=0
+ $Y2=0
cc_390 N_A_1041_333#_c_484_n N_A0_c_631_n 0.00999292f $X=7.485 $Y=1.315 $X2=0
+ $Y2=0
cc_391 N_A_1041_333#_c_485_n N_A0_c_631_n 0.00670874f $X=6.045 $Y=1.315 $X2=0
+ $Y2=0
cc_392 N_A_1041_333#_c_492_n N_A0_c_631_n 0.013216f $X=5.475 $Y=1.65 $X2=0 $Y2=0
cc_393 N_A_1041_333#_c_484_n N_A3_M1025_g 0.0153019f $X=7.485 $Y=1.315 $X2=0
+ $Y2=0
cc_394 N_A_1041_333#_c_497_n N_A3_M1025_g 8.0893e-19 $X=7.57 $Y=1.63 $X2=0 $Y2=0
cc_395 N_A_1041_333#_c_490_n N_A3_M1025_g 4.01131e-19 $X=7.57 $Y=1.29 $X2=0
+ $Y2=0
cc_396 N_A_1041_333#_c_491_n N_A3_M1025_g 0.00878367f $X=7.57 $Y=1.29 $X2=0
+ $Y2=0
cc_397 N_A_1041_333#_M1013_g N_A3_M1012_g 0.0381602f $X=7.3 $Y=2.415 $X2=0 $Y2=0
cc_398 N_A_1041_333#_c_482_n A3 0.00382826f $X=7.57 $Y=1.645 $X2=0 $Y2=0
cc_399 N_A_1041_333#_c_484_n A3 0.0200175f $X=7.485 $Y=1.315 $X2=0 $Y2=0
cc_400 N_A_1041_333#_c_497_n A3 0.00784895f $X=7.57 $Y=1.63 $X2=0 $Y2=0
cc_401 N_A_1041_333#_c_486_n A3 4.96653e-19 $X=7.57 $Y=1.63 $X2=0 $Y2=0
cc_402 N_A_1041_333#_c_482_n N_A3_c_670_n 0.0381602f $X=7.57 $Y=1.645 $X2=0
+ $Y2=0
cc_403 N_A_1041_333#_c_484_n N_A3_c_670_n 0.00459442f $X=7.485 $Y=1.315 $X2=0
+ $Y2=0
cc_404 N_A_1041_333#_c_486_n N_A3_c_670_n 0.00185187f $X=7.57 $Y=1.63 $X2=0
+ $Y2=0
cc_405 N_A_1041_333#_c_483_n N_A2_M1028_g 0.0253094f $X=7.57 $Y=1.125 $X2=0
+ $Y2=0
cc_406 N_A_1041_333#_c_497_n N_A2_M1028_g 4.68321e-19 $X=7.57 $Y=1.63 $X2=0
+ $Y2=0
cc_407 N_A_1041_333#_c_487_n N_A2_M1028_g 0.0150425f $X=8.445 $Y=1.21 $X2=0
+ $Y2=0
cc_408 N_A_1041_333#_c_488_n N_A2_M1028_g 0.00362448f $X=8.53 $Y=1.975 $X2=0
+ $Y2=0
cc_409 N_A_1041_333#_c_490_n N_A2_M1028_g 5.73382e-19 $X=7.57 $Y=1.29 $X2=0
+ $Y2=0
cc_410 N_A_1041_333#_c_491_n N_A2_M1028_g 0.0163002f $X=7.57 $Y=1.29 $X2=0 $Y2=0
cc_411 N_A_1041_333#_c_488_n N_A2_M1003_g 0.00278221f $X=8.53 $Y=1.975 $X2=0
+ $Y2=0
cc_412 N_A_1041_333#_c_538_p N_A2_M1003_g 0.00410043f $X=8.615 $Y=2.06 $X2=0
+ $Y2=0
cc_413 N_A_1041_333#_M1013_g N_A2_c_706_n 2.37237e-19 $X=7.3 $Y=2.415 $X2=0
+ $Y2=0
cc_414 N_A_1041_333#_c_497_n N_A2_c_706_n 2.69288e-19 $X=7.57 $Y=1.63 $X2=0
+ $Y2=0
cc_415 N_A_1041_333#_c_486_n N_A2_c_706_n 0.0233057f $X=7.57 $Y=1.63 $X2=0 $Y2=0
cc_416 N_A_1041_333#_c_487_n N_A2_c_706_n 0.00834032f $X=8.445 $Y=1.21 $X2=0
+ $Y2=0
cc_417 N_A_1041_333#_c_488_n N_A2_c_706_n 0.00764168f $X=8.53 $Y=1.975 $X2=0
+ $Y2=0
cc_418 N_A_1041_333#_M1013_g N_A2_c_707_n 0.00740468f $X=7.3 $Y=2.415 $X2=0
+ $Y2=0
cc_419 N_A_1041_333#_c_497_n N_A2_c_707_n 0.0228972f $X=7.57 $Y=1.63 $X2=0 $Y2=0
cc_420 N_A_1041_333#_c_486_n N_A2_c_707_n 0.00235692f $X=7.57 $Y=1.63 $X2=0
+ $Y2=0
cc_421 N_A_1041_333#_c_487_n N_A2_c_707_n 0.031368f $X=8.445 $Y=1.21 $X2=0 $Y2=0
cc_422 N_A_1041_333#_c_488_n N_A2_c_707_n 0.0347682f $X=8.53 $Y=1.975 $X2=0
+ $Y2=0
cc_423 N_A_1041_333#_c_538_p N_A2_c_707_n 0.011807f $X=8.615 $Y=2.06 $X2=0 $Y2=0
cc_424 N_A_1041_333#_M1002_g N_S0_M1029_g 0.0129015f $X=5.475 $Y=0.805 $X2=0
+ $Y2=0
cc_425 N_A_1041_333#_M1002_g N_S0_c_751_n 0.0101977f $X=5.475 $Y=0.805 $X2=0
+ $Y2=0
cc_426 N_A_1041_333#_M1000_g N_S0_M1020_g 0.0239664f $X=5.28 $Y=2.475 $X2=0
+ $Y2=0
cc_427 N_A_1041_333#_c_485_n N_S0_M1020_g 6.32967e-19 $X=6.045 $Y=1.315 $X2=0
+ $Y2=0
cc_428 N_A_1041_333#_c_492_n N_S0_M1020_g 0.0100075f $X=5.475 $Y=1.65 $X2=0
+ $Y2=0
cc_429 N_A_1041_333#_M1013_g N_S0_c_762_n 0.0104164f $X=7.3 $Y=2.415 $X2=0 $Y2=0
cc_430 N_A_1041_333#_c_483_n N_S0_M1017_g 0.0157105f $X=7.57 $Y=1.125 $X2=0
+ $Y2=0
cc_431 N_A_1041_333#_c_484_n N_S0_M1017_g 0.00467401f $X=7.485 $Y=1.315 $X2=0
+ $Y2=0
cc_432 N_A_1041_333#_c_491_n N_S0_M1017_g 0.0012997f $X=7.57 $Y=1.29 $X2=0 $Y2=0
cc_433 N_A_1041_333#_c_483_n N_S0_c_754_n 0.0100282f $X=7.57 $Y=1.125 $X2=0
+ $Y2=0
cc_434 N_A_1041_333#_M1013_g N_S0_M1010_g 0.0119972f $X=7.3 $Y=2.415 $X2=0 $Y2=0
cc_435 N_A_1041_333#_c_489_n N_S0_c_755_n 0.0082777f $X=9.33 $Y=0.87 $X2=0 $Y2=0
cc_436 N_A_1041_333#_c_499_n N_S0_M1026_g 0.0176207f $X=8.92 $Y=2.06 $X2=0 $Y2=0
cc_437 N_A_1041_333#_c_500_n N_S0_M1026_g 2.30416e-19 $X=9.025 $Y=2.24 $X2=0
+ $Y2=0
cc_438 N_A_1041_333#_c_489_n N_S0_M1026_g 0.00373674f $X=9.33 $Y=0.87 $X2=0
+ $Y2=0
cc_439 N_A_1041_333#_c_489_n N_S0_M1021_g 0.00611172f $X=9.33 $Y=0.87 $X2=0
+ $Y2=0
cc_440 N_A_1041_333#_c_499_n N_S0_c_758_n 6.78821e-19 $X=8.92 $Y=2.06 $X2=0
+ $Y2=0
cc_441 N_A_1041_333#_c_501_n N_S0_c_758_n 0.007459f $X=9.33 $Y=1.975 $X2=0 $Y2=0
cc_442 N_A_1041_333#_c_489_n N_S0_c_758_n 0.00767632f $X=9.33 $Y=0.87 $X2=0
+ $Y2=0
cc_443 N_A_1041_333#_c_487_n S0 0.0132343f $X=8.445 $Y=1.21 $X2=0 $Y2=0
cc_444 N_A_1041_333#_c_488_n S0 0.0344337f $X=8.53 $Y=1.975 $X2=0 $Y2=0
cc_445 N_A_1041_333#_c_499_n S0 0.0140128f $X=8.92 $Y=2.06 $X2=0 $Y2=0
cc_446 N_A_1041_333#_c_489_n S0 0.0628153f $X=9.33 $Y=0.87 $X2=0 $Y2=0
cc_447 N_A_1041_333#_c_487_n N_S0_c_760_n 0.0021959f $X=8.445 $Y=1.21 $X2=0
+ $Y2=0
cc_448 N_A_1041_333#_c_488_n N_S0_c_760_n 0.0063559f $X=8.53 $Y=1.975 $X2=0
+ $Y2=0
cc_449 N_A_1041_333#_c_489_n N_S0_c_760_n 0.00767632f $X=9.33 $Y=0.87 $X2=0
+ $Y2=0
cc_450 N_A_1041_333#_M1000_g N_A_27_119#_c_860_n 0.00774874f $X=5.28 $Y=2.475
+ $X2=0 $Y2=0
cc_451 N_A_1041_333#_M1002_g N_A_27_119#_c_860_n 0.00518227f $X=5.475 $Y=0.805
+ $X2=0 $Y2=0
cc_452 N_A_1041_333#_c_485_n N_A_27_119#_c_860_n 0.0297862f $X=6.045 $Y=1.315
+ $X2=0 $Y2=0
cc_453 N_A_1041_333#_c_492_n N_A_27_119#_c_860_n 0.0148858f $X=5.475 $Y=1.65
+ $X2=0 $Y2=0
cc_454 N_A_1041_333#_M1013_g N_A_27_119#_c_870_n 0.0163692f $X=7.3 $Y=2.415
+ $X2=0 $Y2=0
cc_455 N_A_1041_333#_c_482_n N_A_27_119#_c_870_n 0.00106332f $X=7.57 $Y=1.645
+ $X2=0 $Y2=0
cc_456 N_A_1041_333#_c_485_n N_A_27_119#_c_870_n 0.0238578f $X=6.045 $Y=1.315
+ $X2=0 $Y2=0
cc_457 N_A_1041_333#_c_492_n N_A_27_119#_c_870_n 0.00727793f $X=5.475 $Y=1.65
+ $X2=0 $Y2=0
cc_458 N_A_1041_333#_M1000_g N_A_27_119#_c_909_n 0.00607006f $X=5.28 $Y=2.475
+ $X2=0 $Y2=0
cc_459 N_A_1041_333#_c_484_n N_A_27_119#_c_861_n 0.0292587f $X=7.485 $Y=1.315
+ $X2=0 $Y2=0
cc_460 N_A_1041_333#_c_485_n N_A_27_119#_c_861_n 0.0186442f $X=6.045 $Y=1.315
+ $X2=0 $Y2=0
cc_461 N_A_1041_333#_c_492_n N_A_27_119#_c_861_n 4.55688e-19 $X=5.475 $Y=1.65
+ $X2=0 $Y2=0
cc_462 N_A_1041_333#_M1002_g N_A_27_119#_c_862_n 0.0197881f $X=5.475 $Y=0.805
+ $X2=0 $Y2=0
cc_463 N_A_1041_333#_c_485_n N_A_27_119#_c_862_n 0.0133532f $X=6.045 $Y=1.315
+ $X2=0 $Y2=0
cc_464 N_A_1041_333#_c_492_n N_A_27_119#_c_862_n 0.00294395f $X=5.475 $Y=1.65
+ $X2=0 $Y2=0
cc_465 N_A_1041_333#_c_484_n N_A_27_119#_c_916_n 0.0189446f $X=7.485 $Y=1.315
+ $X2=0 $Y2=0
cc_466 N_A_1041_333#_c_484_n N_A_27_119#_c_863_n 0.0124637f $X=7.485 $Y=1.315
+ $X2=0 $Y2=0
cc_467 N_A_1041_333#_M1013_g N_A_27_119#_c_871_n 6.61294e-19 $X=7.3 $Y=2.415
+ $X2=0 $Y2=0
cc_468 N_A_1041_333#_c_482_n N_A_27_119#_c_871_n 0.00414283f $X=7.57 $Y=1.645
+ $X2=0 $Y2=0
cc_469 N_A_1041_333#_c_497_n N_A_27_119#_c_871_n 0.00788212f $X=7.57 $Y=1.63
+ $X2=0 $Y2=0
cc_470 N_A_1041_333#_M1002_g N_A_27_119#_c_864_n 0.00478503f $X=5.475 $Y=0.805
+ $X2=0 $Y2=0
cc_471 N_A_1041_333#_c_484_n N_A_27_119#_c_864_n 0.00226957f $X=7.485 $Y=1.315
+ $X2=0 $Y2=0
cc_472 N_A_1041_333#_c_483_n N_A_27_119#_c_867_n 0.00334831f $X=7.57 $Y=1.125
+ $X2=0 $Y2=0
cc_473 N_A_1041_333#_c_484_n N_A_27_119#_c_867_n 8.45747e-19 $X=7.485 $Y=1.315
+ $X2=0 $Y2=0
cc_474 N_A_1041_333#_c_490_n N_A_27_119#_c_867_n 0.00226363f $X=7.57 $Y=1.29
+ $X2=0 $Y2=0
cc_475 N_A_1041_333#_c_483_n N_A_27_119#_c_868_n 0.00988304f $X=7.57 $Y=1.125
+ $X2=0 $Y2=0
cc_476 N_A_1041_333#_c_484_n N_A_27_119#_c_868_n 0.00907616f $X=7.485 $Y=1.315
+ $X2=0 $Y2=0
cc_477 N_A_1041_333#_c_490_n N_A_27_119#_c_868_n 0.00239769f $X=7.57 $Y=1.29
+ $X2=0 $Y2=0
cc_478 N_A_1041_333#_c_491_n N_A_27_119#_c_868_n 0.00163631f $X=7.57 $Y=1.29
+ $X2=0 $Y2=0
cc_479 N_A_1041_333#_M1002_g N_A_200_119#_c_1026_n 0.00192944f $X=5.475 $Y=0.805
+ $X2=0 $Y2=0
cc_480 N_A_1041_333#_c_492_n N_A_200_119#_c_1026_n 0.00190736f $X=5.475 $Y=1.65
+ $X2=0 $Y2=0
cc_481 N_A_1041_333#_M1000_g N_A_200_119#_c_1069_n 0.00424204f $X=5.28 $Y=2.475
+ $X2=0 $Y2=0
cc_482 N_A_1041_333#_M1000_g N_A_200_119#_c_1076_n 0.013721f $X=5.28 $Y=2.475
+ $X2=0 $Y2=0
cc_483 N_A_1041_333#_c_492_n N_A_200_119#_c_1076_n 3.4112e-19 $X=5.475 $Y=1.65
+ $X2=0 $Y2=0
cc_484 N_A_1041_333#_M1000_g N_A_200_119#_c_1032_n 0.0010653f $X=5.28 $Y=2.475
+ $X2=0 $Y2=0
cc_485 N_A_1041_333#_c_499_n N_VPWR_M1003_d 8.27517e-19 $X=8.92 $Y=2.06 $X2=0
+ $Y2=0
cc_486 N_A_1041_333#_c_538_p N_VPWR_M1003_d 0.00143441f $X=8.615 $Y=2.06 $X2=0
+ $Y2=0
cc_487 N_A_1041_333#_c_499_n N_VPWR_c_1132_n 0.00351911f $X=8.92 $Y=2.06 $X2=0
+ $Y2=0
cc_488 N_A_1041_333#_c_538_p N_VPWR_c_1132_n 0.00641018f $X=8.615 $Y=2.06 $X2=0
+ $Y2=0
cc_489 N_A_1041_333#_c_500_n N_VPWR_c_1132_n 5.83564e-19 $X=9.025 $Y=2.24 $X2=0
+ $Y2=0
cc_490 N_A_1041_333#_M1000_g N_VPWR_c_1140_n 0.00352758f $X=5.28 $Y=2.475 $X2=0
+ $Y2=0
cc_491 N_A_1041_333#_c_500_n N_VPWR_c_1141_n 0.00464591f $X=9.025 $Y=2.24 $X2=0
+ $Y2=0
cc_492 N_A_1041_333#_M1000_g N_VPWR_c_1127_n 0.00495025f $X=5.28 $Y=2.475 $X2=0
+ $Y2=0
cc_493 N_A_1041_333#_M1013_g N_VPWR_c_1127_n 9.39239e-19 $X=7.3 $Y=2.415 $X2=0
+ $Y2=0
cc_494 N_A_1041_333#_c_500_n N_VPWR_c_1127_n 0.00651069f $X=9.025 $Y=2.24 $X2=0
+ $Y2=0
cc_495 N_A_1041_333#_c_483_n N_VGND_c_1295_n 0.00114854f $X=7.57 $Y=1.125 $X2=0
+ $Y2=0
cc_496 N_A_1041_333#_c_487_n N_VGND_c_1295_n 0.016976f $X=8.445 $Y=1.21 $X2=0
+ $Y2=0
cc_497 N_A_1041_333#_M1002_g N_VGND_c_1305_n 4.63031e-19 $X=5.475 $Y=0.805 $X2=0
+ $Y2=0
cc_498 N_A_1041_333#_c_483_n N_VGND_c_1305_n 3.69739e-19 $X=7.57 $Y=1.125 $X2=0
+ $Y2=0
cc_499 N_A_1041_333#_c_489_n N_VGND_c_1305_n 0.0137519f $X=9.33 $Y=0.87 $X2=0
+ $Y2=0
cc_500 N_A0_c_627_n N_A3_M1025_g 0.0152456f $X=6.145 $Y=1.2 $X2=0 $Y2=0
cc_501 N_A0_M1019_g N_A3_M1012_g 0.0155107f $X=6.22 $Y=2.415 $X2=0 $Y2=0
cc_502 A0 A3 0.0229602f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_503 N_A0_c_630_n A3 3.07797e-19 $X=6.31 $Y=1.745 $X2=0 $Y2=0
cc_504 A0 N_A3_c_670_n 0.00219587f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_505 N_A0_c_630_n N_A3_c_670_n 0.0205108f $X=6.31 $Y=1.745 $X2=0 $Y2=0
cc_506 N_A0_c_626_n N_S0_c_751_n 0.0100906f $X=5.835 $Y=1.125 $X2=0 $Y2=0
cc_507 N_A0_M1019_g N_S0_M1020_g 0.0290784f $X=6.22 $Y=2.415 $X2=0 $Y2=0
cc_508 N_A0_M1019_g N_S0_c_762_n 0.0103107f $X=6.22 $Y=2.415 $X2=0 $Y2=0
cc_509 N_A0_M1019_g N_A_27_119#_c_870_n 0.0180864f $X=6.22 $Y=2.415 $X2=0 $Y2=0
cc_510 A0 N_A_27_119#_c_870_n 0.0245868f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_511 N_A0_c_630_n N_A_27_119#_c_870_n 0.00400978f $X=6.31 $Y=1.745 $X2=0 $Y2=0
cc_512 N_A0_c_626_n N_A_27_119#_c_861_n 0.01119f $X=5.835 $Y=1.125 $X2=0 $Y2=0
cc_513 N_A0_c_627_n N_A_27_119#_c_861_n 0.00946491f $X=6.145 $Y=1.2 $X2=0 $Y2=0
cc_514 N_A0_c_626_n N_A_27_119#_c_862_n 0.00499735f $X=5.835 $Y=1.125 $X2=0
+ $Y2=0
cc_515 N_A0_c_626_n N_A_27_119#_c_863_n 0.00366313f $X=5.835 $Y=1.125 $X2=0
+ $Y2=0
cc_516 N_A0_c_626_n N_A_27_119#_c_864_n 0.00564173f $X=5.835 $Y=1.125 $X2=0
+ $Y2=0
cc_517 N_A0_M1019_g N_VPWR_c_1131_n 0.0101766f $X=6.22 $Y=2.415 $X2=0 $Y2=0
cc_518 N_A0_M1019_g N_VPWR_c_1127_n 7.88961e-19 $X=6.22 $Y=2.415 $X2=0 $Y2=0
cc_519 N_A0_c_626_n N_VGND_c_1294_n 0.00684327f $X=5.835 $Y=1.125 $X2=0 $Y2=0
cc_520 N_A0_c_626_n N_VGND_c_1305_n 4.63031e-19 $X=5.835 $Y=1.125 $X2=0 $Y2=0
cc_521 N_A3_M1025_g N_S0_c_751_n 0.00992583f $X=6.76 $Y=0.805 $X2=0 $Y2=0
cc_522 N_A3_M1012_g N_S0_c_762_n 0.0104164f $X=6.94 $Y=2.415 $X2=0 $Y2=0
cc_523 N_A3_M1025_g N_S0_M1017_g 0.0438952f $X=6.76 $Y=0.805 $X2=0 $Y2=0
cc_524 N_A3_M1012_g N_A_27_119#_c_870_n 0.0154483f $X=6.94 $Y=2.415 $X2=0 $Y2=0
cc_525 A3 N_A_27_119#_c_870_n 0.0197155f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_526 N_A3_c_670_n N_A_27_119#_c_870_n 0.00578533f $X=6.85 $Y=1.745 $X2=0 $Y2=0
cc_527 N_A3_M1025_g N_A_27_119#_c_916_n 0.0118868f $X=6.76 $Y=0.805 $X2=0 $Y2=0
cc_528 N_A3_M1025_g N_A_27_119#_c_863_n 0.0035227f $X=6.76 $Y=0.805 $X2=0 $Y2=0
cc_529 N_A3_M1025_g N_A_27_119#_c_864_n 0.00570797f $X=6.76 $Y=0.805 $X2=0 $Y2=0
cc_530 N_A3_M1012_g N_VPWR_c_1131_n 0.00888388f $X=6.94 $Y=2.415 $X2=0 $Y2=0
cc_531 N_A3_M1012_g N_VPWR_c_1127_n 9.39239e-19 $X=6.94 $Y=2.415 $X2=0 $Y2=0
cc_532 N_A3_M1025_g N_VGND_c_1294_n 0.00547728f $X=6.76 $Y=0.805 $X2=0 $Y2=0
cc_533 N_A3_M1025_g N_VGND_c_1305_n 4.63031e-19 $X=6.76 $Y=0.805 $X2=0 $Y2=0
cc_534 N_A2_M1028_g N_S0_c_754_n 0.0103107f $X=8.02 $Y=0.805 $X2=0 $Y2=0
cc_535 N_A2_M1003_g N_S0_M1010_g 0.0236847f $X=8.38 $Y=2.415 $X2=0 $Y2=0
cc_536 N_A2_c_707_n N_S0_M1010_g 0.0306909f $X=8.18 $Y=1.65 $X2=0 $Y2=0
cc_537 N_A2_M1003_g N_S0_c_765_n 0.0104164f $X=8.38 $Y=2.415 $X2=0 $Y2=0
cc_538 N_A2_c_707_n N_S0_c_765_n 0.00502333f $X=8.18 $Y=1.65 $X2=0 $Y2=0
cc_539 N_A2_c_706_n N_S0_c_755_n 0.0216494f $X=8.18 $Y=1.65 $X2=0 $Y2=0
cc_540 N_A2_M1003_g N_S0_c_758_n 0.0216494f $X=8.38 $Y=2.415 $X2=0 $Y2=0
cc_541 N_A2_c_706_n S0 2.76309e-19 $X=8.18 $Y=1.65 $X2=0 $Y2=0
cc_542 N_A2_M1028_g N_S0_c_760_n 0.00412836f $X=8.02 $Y=0.805 $X2=0 $Y2=0
cc_543 N_A2_c_707_n N_A_27_119#_c_871_n 0.0438543f $X=8.18 $Y=1.65 $X2=0 $Y2=0
cc_544 N_A2_M1028_g N_A_27_119#_c_867_n 0.00104645f $X=8.02 $Y=0.805 $X2=0 $Y2=0
cc_545 N_A2_M1028_g N_A_27_119#_c_868_n 0.00167977f $X=8.02 $Y=0.805 $X2=0 $Y2=0
cc_546 N_A2_M1003_g N_VPWR_c_1132_n 0.0011622f $X=8.38 $Y=2.415 $X2=0 $Y2=0
cc_547 N_A2_c_707_n N_VPWR_c_1132_n 0.00836902f $X=8.18 $Y=1.65 $X2=0 $Y2=0
cc_548 N_A2_c_707_n N_VPWR_c_1137_n 0.0125423f $X=8.18 $Y=1.65 $X2=0 $Y2=0
cc_549 N_A2_M1003_g N_VPWR_c_1127_n 9.39239e-19 $X=8.38 $Y=2.415 $X2=0 $Y2=0
cc_550 N_A2_c_707_n N_VPWR_c_1127_n 0.0127744f $X=8.18 $Y=1.65 $X2=0 $Y2=0
cc_551 N_A2_c_707_n A_1589_431# 0.00458965f $X=8.18 $Y=1.65 $X2=-0.19 $Y2=-0.245
cc_552 N_A2_M1028_g N_VGND_c_1295_n 0.0099495f $X=8.02 $Y=0.805 $X2=0 $Y2=0
cc_553 N_A2_M1028_g N_VGND_c_1305_n 7.88961e-19 $X=8.02 $Y=0.805 $X2=0 $Y2=0
cc_554 N_S0_M1020_g N_A_27_119#_c_860_n 0.00126386f $X=5.71 $Y=2.475 $X2=0 $Y2=0
cc_555 N_S0_M1020_g N_A_27_119#_c_870_n 0.0146283f $X=5.71 $Y=2.475 $X2=0 $Y2=0
cc_556 N_S0_c_751_n N_A_27_119#_c_861_n 0.00603594f $X=7.045 $Y=0.18 $X2=0 $Y2=0
cc_557 N_S0_M1029_g N_A_27_119#_c_862_n 5.16498e-19 $X=5.045 $Y=0.805 $X2=0
+ $Y2=0
cc_558 N_S0_c_751_n N_A_27_119#_c_862_n 0.00278424f $X=7.045 $Y=0.18 $X2=0 $Y2=0
cc_559 N_S0_c_751_n N_A_27_119#_c_916_n 0.0020557f $X=7.045 $Y=0.18 $X2=0 $Y2=0
cc_560 N_S0_M1017_g N_A_27_119#_c_916_n 0.00951763f $X=7.12 $Y=0.805 $X2=0 $Y2=0
cc_561 N_S0_c_751_n N_A_27_119#_c_863_n 0.0027666f $X=7.045 $Y=0.18 $X2=0 $Y2=0
cc_562 N_S0_c_762_n N_A_27_119#_c_871_n 0.00422132f $X=7.795 $Y=3.15 $X2=0 $Y2=0
cc_563 N_S0_M1010_g N_A_27_119#_c_871_n 0.00520417f $X=7.87 $Y=2.475 $X2=0 $Y2=0
cc_564 N_S0_M1029_g N_A_27_119#_c_864_n 0.0045807f $X=5.045 $Y=0.805 $X2=0 $Y2=0
cc_565 N_S0_c_751_n N_A_27_119#_c_864_n 0.01252f $X=7.045 $Y=0.18 $X2=0 $Y2=0
cc_566 N_S0_M1017_g N_A_27_119#_c_864_n 0.00423616f $X=7.12 $Y=0.805 $X2=0 $Y2=0
cc_567 N_S0_M1017_g N_A_27_119#_c_867_n 7.01026e-19 $X=7.12 $Y=0.805 $X2=0 $Y2=0
cc_568 N_S0_c_754_n N_A_27_119#_c_867_n 0.00257847f $X=9.02 $Y=0.18 $X2=0 $Y2=0
cc_569 N_S0_M1017_g N_A_27_119#_c_868_n 0.00313613f $X=7.12 $Y=0.805 $X2=0 $Y2=0
cc_570 N_S0_c_754_n N_A_27_119#_c_868_n 0.00398847f $X=9.02 $Y=0.18 $X2=0 $Y2=0
cc_571 N_S0_M1029_g N_A_200_119#_c_1026_n 0.00720592f $X=5.045 $Y=0.805 $X2=0
+ $Y2=0
cc_572 N_S0_M1029_g N_A_200_119#_c_1071_n 0.010973f $X=5.045 $Y=0.805 $X2=0
+ $Y2=0
cc_573 N_S0_c_751_n N_A_200_119#_c_1071_n 0.00249633f $X=7.045 $Y=0.18 $X2=0
+ $Y2=0
cc_574 N_S0_M1020_g N_VPWR_c_1131_n 0.00692722f $X=5.71 $Y=2.475 $X2=0 $Y2=0
cc_575 N_S0_c_762_n N_VPWR_c_1131_n 0.0254387f $X=7.795 $Y=3.15 $X2=0 $Y2=0
cc_576 N_S0_M1010_g N_VPWR_c_1132_n 0.00498297f $X=7.87 $Y=2.475 $X2=0 $Y2=0
cc_577 N_S0_c_765_n N_VPWR_c_1132_n 0.0173925f $X=8.735 $Y=3.15 $X2=0 $Y2=0
cc_578 N_S0_M1026_g N_VPWR_c_1132_n 0.01166f $X=8.81 $Y=2.415 $X2=0 $Y2=0
cc_579 N_S0_c_762_n N_VPWR_c_1137_n 0.0601747f $X=7.795 $Y=3.15 $X2=0 $Y2=0
cc_580 N_S0_c_763_n N_VPWR_c_1140_n 0.0232701f $X=5.785 $Y=3.15 $X2=0 $Y2=0
cc_581 N_S0_c_765_n N_VPWR_c_1141_n 0.00718072f $X=8.735 $Y=3.15 $X2=0 $Y2=0
cc_582 N_S0_c_762_n N_VPWR_c_1127_n 0.0771075f $X=7.795 $Y=3.15 $X2=0 $Y2=0
cc_583 N_S0_c_763_n N_VPWR_c_1127_n 0.0116041f $X=5.785 $Y=3.15 $X2=0 $Y2=0
cc_584 N_S0_c_765_n N_VPWR_c_1127_n 0.0300227f $X=8.735 $Y=3.15 $X2=0 $Y2=0
cc_585 N_S0_c_767_n N_VPWR_c_1127_n 0.00540001f $X=7.87 $Y=3.15 $X2=0 $Y2=0
cc_586 S0 N_VGND_M1028_d 0.0138089f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_587 N_S0_c_752_n N_VGND_c_1293_n 0.00797946f $X=5.12 $Y=0.18 $X2=0 $Y2=0
cc_588 N_S0_c_751_n N_VGND_c_1294_n 0.0254714f $X=7.045 $Y=0.18 $X2=0 $Y2=0
cc_589 N_S0_c_754_n N_VGND_c_1295_n 0.0255272f $X=9.02 $Y=0.18 $X2=0 $Y2=0
cc_590 N_S0_M1021_g N_VGND_c_1295_n 0.00383582f $X=9.095 $Y=0.805 $X2=0 $Y2=0
cc_591 S0 N_VGND_c_1295_n 0.0159357f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_592 N_S0_c_751_n N_VGND_c_1300_n 0.0528188f $X=7.045 $Y=0.18 $X2=0 $Y2=0
cc_593 N_S0_c_752_n N_VGND_c_1303_n 0.0319333f $X=5.12 $Y=0.18 $X2=0 $Y2=0
cc_594 N_S0_c_754_n N_VGND_c_1304_n 0.0256944f $X=9.02 $Y=0.18 $X2=0 $Y2=0
cc_595 S0 N_VGND_c_1304_n 0.00563096f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_596 N_S0_c_751_n N_VGND_c_1305_n 0.032005f $X=7.045 $Y=0.18 $X2=0 $Y2=0
cc_597 N_S0_c_752_n N_VGND_c_1305_n 0.00585472f $X=5.12 $Y=0.18 $X2=0 $Y2=0
cc_598 N_S0_c_754_n N_VGND_c_1305_n 0.0694898f $X=9.02 $Y=0.18 $X2=0 $Y2=0
cc_599 N_S0_c_757_n N_VGND_c_1305_n 0.00360983f $X=7.12 $Y=0.18 $X2=0 $Y2=0
cc_600 S0 N_VGND_c_1305_n 0.00567022f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_601 N_A_27_119#_c_864_n N_A_200_119#_M1006_d 0.00370184f $X=7.295 $Y=0.555
+ $X2=-0.19 $Y2=-0.245
cc_602 N_A_27_119#_c_864_n N_A_200_119#_M1029_d 0.00181506f $X=7.295 $Y=0.555
+ $X2=0 $Y2=0
cc_603 N_A_27_119#_c_870_n N_A_200_119#_M1000_d 0.00165893f $X=7.41 $Y=2.175
+ $X2=0 $Y2=0
cc_604 N_A_27_119#_c_864_n N_A_200_119#_c_1025_n 0.00659353f $X=7.295 $Y=0.555
+ $X2=0 $Y2=0
cc_605 N_A_27_119#_c_860_n N_A_200_119#_c_1026_n 0.0485383f $X=5.34 $Y=2.09
+ $X2=0 $Y2=0
cc_606 N_A_27_119#_c_862_n N_A_200_119#_c_1026_n 0.0191698f $X=5.695 $Y=0.965
+ $X2=0 $Y2=0
cc_607 N_A_27_119#_c_909_n N_A_200_119#_c_1069_n 0.00710653f $X=5.425 $Y=2.175
+ $X2=0 $Y2=0
cc_608 N_A_27_119#_c_870_n N_A_200_119#_c_1076_n 0.0111713f $X=7.41 $Y=2.175
+ $X2=0 $Y2=0
cc_609 N_A_27_119#_c_909_n N_A_200_119#_c_1076_n 0.00860732f $X=5.425 $Y=2.175
+ $X2=0 $Y2=0
cc_610 N_A_27_119#_c_862_n N_A_200_119#_c_1071_n 0.00711279f $X=5.695 $Y=0.965
+ $X2=0 $Y2=0
cc_611 N_A_27_119#_c_864_n N_A_200_119#_c_1071_n 0.0163182f $X=7.295 $Y=0.555
+ $X2=0 $Y2=0
cc_612 N_A_27_119#_c_860_n N_A_200_119#_c_1032_n 0.00730991f $X=5.34 $Y=2.09
+ $X2=0 $Y2=0
cc_613 N_A_27_119#_c_909_n N_A_200_119#_c_1032_n 0.00638402f $X=5.425 $Y=2.175
+ $X2=0 $Y2=0
cc_614 N_A_27_119#_c_870_n N_VPWR_M1019_d 0.0128502f $X=7.41 $Y=2.175 $X2=0
+ $Y2=0
cc_615 N_A_27_119#_c_870_n N_VPWR_c_1131_n 0.0177446f $X=7.41 $Y=2.175 $X2=0
+ $Y2=0
cc_616 N_A_27_119#_c_866_n N_VPWR_c_1133_n 0.00392426f $X=0.24 $Y=0.555 $X2=0
+ $Y2=0
cc_617 N_A_27_119#_c_871_n N_VPWR_c_1137_n 0.00476636f $X=7.515 $Y=2.255 $X2=0
+ $Y2=0
cc_618 N_A_27_119#_c_871_n N_VPWR_c_1127_n 0.00578995f $X=7.515 $Y=2.255 $X2=0
+ $Y2=0
cc_619 N_A_27_119#_c_866_n N_VPWR_c_1127_n 0.00615101f $X=0.24 $Y=0.555 $X2=0
+ $Y2=0
cc_620 N_A_27_119#_c_864_n N_X_M1014_d 0.00195104f $X=7.295 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_621 N_A_27_119#_c_864_n N_X_M1024_d 0.00112111f $X=7.295 $Y=0.555 $X2=0 $Y2=0
cc_622 N_A_27_119#_c_864_n N_X_c_1240_n 0.0188308f $X=7.295 $Y=0.555 $X2=0 $Y2=0
cc_623 N_A_27_119#_c_864_n N_X_c_1241_n 0.0216587f $X=7.295 $Y=0.555 $X2=0 $Y2=0
cc_624 N_A_27_119#_c_864_n N_X_c_1263_n 0.0185492f $X=7.295 $Y=0.555 $X2=0 $Y2=0
cc_625 N_A_27_119#_c_864_n X 0.00368039f $X=7.295 $Y=0.555 $X2=0 $Y2=0
cc_626 N_A_27_119#_c_870_n A_1157_431# 0.00938627f $X=7.41 $Y=2.175 $X2=-0.19
+ $Y2=-0.245
cc_627 N_A_27_119#_c_870_n A_1403_419# 0.00366293f $X=7.41 $Y=2.175 $X2=-0.19
+ $Y2=-0.245
cc_628 N_A_27_119#_c_864_n N_VGND_M1007_d 0.00264513f $X=7.295 $Y=0.555
+ $X2=-0.19 $Y2=-0.245
cc_629 N_A_27_119#_c_864_n N_VGND_M1015_s 0.00279618f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_630 N_A_27_119#_c_864_n N_VGND_M1027_s 0.0034847f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_631 N_A_27_119#_c_861_n N_VGND_M1030_d 0.00737346f $X=6.475 $Y=0.965 $X2=0
+ $Y2=0
cc_632 N_A_27_119#_c_863_n N_VGND_M1030_d 0.00530059f $X=6.56 $Y=0.82 $X2=0
+ $Y2=0
cc_633 N_A_27_119#_c_864_n N_VGND_M1030_d 0.00370396f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_634 N_A_27_119#_c_864_n N_VGND_c_1291_n 0.00715658f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_635 N_A_27_119#_c_864_n N_VGND_c_1292_n 0.00804044f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_636 N_A_27_119#_c_864_n N_VGND_c_1293_n 0.0218917f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_637 N_A_27_119#_c_861_n N_VGND_c_1294_n 0.0235419f $X=6.475 $Y=0.965 $X2=0
+ $Y2=0
cc_638 N_A_27_119#_c_864_n N_VGND_c_1294_n 0.0243335f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_639 N_A_27_119#_c_867_n N_VGND_c_1295_n 0.0054979f $X=7.44 $Y=0.555 $X2=0
+ $Y2=0
cc_640 N_A_27_119#_c_868_n N_VGND_c_1295_n 0.00792839f $X=7.44 $Y=0.555 $X2=0
+ $Y2=0
cc_641 N_A_27_119#_c_864_n N_VGND_c_1296_n 0.00228771f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_642 N_A_27_119#_c_864_n N_VGND_c_1298_n 0.00228771f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_643 N_A_27_119#_c_916_n N_VGND_c_1300_n 0.00597284f $X=7.23 $Y=0.82 $X2=0
+ $Y2=0
cc_644 N_A_27_119#_c_863_n N_VGND_c_1300_n 0.00202153f $X=6.56 $Y=0.82 $X2=0
+ $Y2=0
cc_645 N_A_27_119#_c_864_n N_VGND_c_1300_n 0.0034697f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_646 N_A_27_119#_c_867_n N_VGND_c_1300_n 0.00105355f $X=7.44 $Y=0.555 $X2=0
+ $Y2=0
cc_647 N_A_27_119#_c_868_n N_VGND_c_1300_n 0.00886512f $X=7.44 $Y=0.555 $X2=0
+ $Y2=0
cc_648 N_A_27_119#_c_864_n N_VGND_c_1302_n 0.00274162f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_649 N_A_27_119#_c_865_n N_VGND_c_1302_n 0.00110095f $X=0.385 $Y=0.555 $X2=0
+ $Y2=0
cc_650 N_A_27_119#_c_866_n N_VGND_c_1302_n 0.00658194f $X=0.24 $Y=0.555 $X2=0
+ $Y2=0
cc_651 N_A_27_119#_c_864_n N_VGND_c_1303_n 0.00669128f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_652 N_A_27_119#_c_864_n N_VGND_c_1305_n 0.547138f $X=7.295 $Y=0.555 $X2=0
+ $Y2=0
cc_653 N_A_27_119#_c_865_n N_VGND_c_1305_n 0.0273116f $X=0.385 $Y=0.555 $X2=0
+ $Y2=0
cc_654 N_A_27_119#_c_866_n N_VGND_c_1305_n 9.51068e-19 $X=0.24 $Y=0.555 $X2=0
+ $Y2=0
cc_655 N_A_27_119#_c_867_n N_VGND_c_1305_n 0.0268291f $X=7.44 $Y=0.555 $X2=0
+ $Y2=0
cc_656 N_A_27_119#_c_868_n N_VGND_c_1305_n 0.00170736f $X=7.44 $Y=0.555 $X2=0
+ $Y2=0
cc_657 N_A_27_119#_c_864_n A_952_119# 0.00556504f $X=7.295 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_658 N_A_27_119#_c_862_n A_1110_119# 6.23616e-19 $X=5.695 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_659 N_A_27_119#_c_864_n A_1110_119# 0.0018284f $X=7.295 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_660 N_A_27_119#_c_916_n A_1367_119# 0.00266715f $X=7.23 $Y=0.82 $X2=-0.19
+ $Y2=-0.245
cc_661 N_A_27_119#_c_864_n A_1367_119# 0.00156881f $X=7.295 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_662 N_A_200_119#_c_1029_n N_VPWR_M1016_d 0.0114899f $X=4.045 $Y=2.455
+ $X2=-0.19 $Y2=-0.245
cc_663 N_A_200_119#_c_1029_n N_VPWR_M1011_d 0.00440501f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_664 N_A_200_119#_c_1029_n N_VPWR_M1022_d 0.00372468f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_665 N_A_200_119#_c_1056_n N_VPWR_M1022_d 0.00331509f $X=4.13 $Y=2.37 $X2=0
+ $Y2=0
cc_666 N_A_200_119#_c_1030_n N_VPWR_M1022_d 0.0277268f $X=4.905 $Y=2.08 $X2=0
+ $Y2=0
cc_667 N_A_200_119#_c_1058_n N_VPWR_M1022_d 0.00139724f $X=4.215 $Y=2.08 $X2=0
+ $Y2=0
cc_668 N_A_200_119#_c_1029_n N_VPWR_c_1128_n 0.0199326f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_669 N_A_200_119#_c_1029_n N_VPWR_c_1129_n 0.0154997f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_670 N_A_200_119#_c_1029_n N_VPWR_c_1130_n 0.0138718f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_671 N_A_200_119#_c_1056_n N_VPWR_c_1130_n 0.00179625f $X=4.13 $Y=2.37 $X2=0
+ $Y2=0
cc_672 N_A_200_119#_c_1030_n N_VPWR_c_1130_n 0.0255687f $X=4.905 $Y=2.08 $X2=0
+ $Y2=0
cc_673 N_A_200_119#_c_1069_n N_VPWR_c_1130_n 0.00669417f $X=4.99 $Y=2.44 $X2=0
+ $Y2=0
cc_674 N_A_200_119#_c_1070_n N_VPWR_c_1130_n 0.0260542f $X=5.075 $Y=2.605 $X2=0
+ $Y2=0
cc_675 N_A_200_119#_c_1027_n N_VPWR_c_1133_n 0.00400008f $X=1.14 $Y=2.37 $X2=0
+ $Y2=0
cc_676 N_A_200_119#_c_1070_n N_VPWR_c_1140_n 0.00313099f $X=5.075 $Y=2.605 $X2=0
+ $Y2=0
cc_677 N_A_200_119#_c_1076_n N_VPWR_c_1140_n 0.00985599f $X=5.495 $Y=2.605 $X2=0
+ $Y2=0
cc_678 N_A_200_119#_c_1027_n N_VPWR_c_1127_n 0.00624159f $X=1.14 $Y=2.37 $X2=0
+ $Y2=0
cc_679 N_A_200_119#_c_1029_n N_VPWR_c_1127_n 0.0842472f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_680 N_A_200_119#_c_1070_n N_VPWR_c_1127_n 0.00534071f $X=5.075 $Y=2.605 $X2=0
+ $Y2=0
cc_681 N_A_200_119#_c_1076_n N_VPWR_c_1127_n 0.0161257f $X=5.495 $Y=2.605 $X2=0
+ $Y2=0
cc_682 N_A_200_119#_c_1029_n N_X_M1005_s 0.00580401f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_683 N_A_200_119#_c_1029_n N_X_M1018_s 0.00580046f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_684 N_A_200_119#_c_1029_n N_X_c_1231_n 0.0250254f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_685 N_A_200_119#_c_1029_n N_X_c_1233_n 0.0105453f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_686 N_A_200_119#_c_1058_n N_X_c_1233_n 0.00517053f $X=4.215 $Y=2.08 $X2=0
+ $Y2=0
cc_687 N_A_200_119#_c_1069_n A_999_431# 0.00281033f $X=4.99 $Y=2.44 $X2=-0.19
+ $Y2=-0.245
cc_688 N_A_200_119#_c_1070_n A_999_431# 3.81944e-19 $X=5.075 $Y=2.605 $X2=-0.19
+ $Y2=-0.245
cc_689 N_A_200_119#_c_1076_n A_999_431# 0.00414458f $X=5.495 $Y=2.605 $X2=-0.19
+ $Y2=-0.245
cc_690 N_A_200_119#_c_1071_n N_VGND_c_1293_n 0.0101896f $X=5.26 $Y=0.79 $X2=0
+ $Y2=0
cc_691 N_A_200_119#_c_1071_n N_VGND_c_1303_n 0.00634659f $X=5.26 $Y=0.79 $X2=0
+ $Y2=0
cc_692 N_A_200_119#_c_1026_n A_952_119# 7.05114e-19 $X=4.99 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_693 N_A_200_119#_c_1071_n A_952_119# 0.00432011f $X=5.26 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_694 N_VPWR_M1011_d N_X_c_1231_n 0.00267082f $X=3.21 $Y=1.675 $X2=0 $Y2=0
cc_695 N_VPWR_M1022_d N_X_c_1233_n 0.00279815f $X=4.07 $Y=1.675 $X2=0 $Y2=0
cc_696 N_X_c_1241_n N_VGND_M1015_s 0.00387652f $X=3.825 $Y=0.945 $X2=0 $Y2=0
cc_697 N_X_c_1240_n N_VGND_c_1291_n 0.00165123f $X=3.07 $Y=0.525 $X2=0 $Y2=0
cc_698 N_X_c_1240_n N_VGND_c_1292_n 0.00165384f $X=3.07 $Y=0.525 $X2=0 $Y2=0
cc_699 N_X_c_1241_n N_VGND_c_1292_n 0.00589743f $X=3.825 $Y=0.945 $X2=0 $Y2=0
cc_700 N_X_c_1263_n N_VGND_c_1292_n 0.00165384f $X=3.93 $Y=0.525 $X2=0 $Y2=0
cc_701 N_X_c_1263_n N_VGND_c_1293_n 0.00385895f $X=3.93 $Y=0.525 $X2=0 $Y2=0
cc_702 N_X_c_1240_n N_VGND_c_1296_n 0.00784537f $X=3.07 $Y=0.525 $X2=0 $Y2=0
cc_703 N_X_c_1263_n N_VGND_c_1298_n 0.00785174f $X=3.93 $Y=0.525 $X2=0 $Y2=0
cc_704 N_X_M1014_d N_VGND_c_1305_n 0.00165127f $X=2.93 $Y=0.235 $X2=0 $Y2=0
cc_705 N_X_M1024_d N_VGND_c_1305_n 0.00165127f $X=3.79 $Y=0.235 $X2=0 $Y2=0
cc_706 N_X_c_1240_n N_VGND_c_1305_n 0.00250034f $X=3.07 $Y=0.525 $X2=0 $Y2=0
cc_707 N_X_c_1263_n N_VGND_c_1305_n 0.00250354f $X=3.93 $Y=0.525 $X2=0 $Y2=0
