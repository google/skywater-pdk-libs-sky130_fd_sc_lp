* File: sky130_fd_sc_lp__a211o_1.spice
* Created: Wed Sep  2 09:17:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a211o_1.pex.spice"
.subckt sky130_fd_sc_lp__a211o_1  VNB VPB A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_80_237#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.3066 AS=0.2226 PD=1.57 PS=2.21 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1002 A_294_47# N_A2_M1002_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.3066 PD=1.08 PS=1.57 NRD=9.276 NRS=0 M=1 R=5.6 SA=75001.1 SB=75001.7
+ A=0.126 P=1.98 MULT=1
MM1001 N_A_80_237#_M1001_d N_A1_M1001_g A_294_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1764 AS=0.1008 PD=1.26 PS=1.08 NRD=9.996 NRS=9.276 M=1 R=5.6 SA=75001.5
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_B1_M1006_g N_A_80_237#_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1764 PD=1.2 PS=1.26 NRD=5.712 NRS=9.996 M=1 R=5.6 SA=75002
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1007 N_A_80_237#_M1007_d N_C1_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1512 PD=2.21 PS=1.2 NRD=0 NRS=5.712 M=1 R=5.6 SA=75002.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A_80_237#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_217_367#_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.3339 PD=1.62 PS=3.05 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1004 N_A_217_367#_M1004_d N_A1_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.2268 PD=1.62 PS=1.62 NRD=7.0329 NRS=6.2449 M=1 R=8.4
+ SA=75000.7 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 A_504_367# N_B1_M1005_g N_A_217_367#_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1701 AS=0.2268 PD=1.53 PS=1.62 NRD=12.4898 NRS=5.4569 M=1 R=8.4
+ SA=75001.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_A_80_237#_M1000_d N_C1_M1000_g A_504_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1701 PD=3.05 PS=1.53 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75001.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a211o_1.pxi.spice"
*
.ends
*
*
