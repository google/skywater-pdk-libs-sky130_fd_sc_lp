* File: sky130_fd_sc_lp__a31oi_4.pex.spice
* Created: Wed Sep  2 09:27:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31OI_4%A3 3 7 11 15 19 23 27 31 33 34 35 36 37 38
+ 64
c82 38 0 8.15747e-20 $X=2.64 $Y=1.665
r83 63 64 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.835 $Y2=1.51
r84 61 63 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.745 $Y=1.51
+ $X2=1.765 $Y2=1.51
r85 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.745
+ $Y=1.51 $X2=1.745 $Y2=1.51
r86 58 61 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.405 $Y=1.51
+ $X2=1.745 $Y2=1.51
r87 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.405
+ $Y=1.51 $X2=1.405 $Y2=1.51
r88 56 58 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.405 $Y2=1.51
r89 55 56 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=0.975 $Y=1.51
+ $X2=1.335 $Y2=1.51
r90 54 55 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=0.975 $Y2=1.51
r91 52 54 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.725 $Y=1.51
+ $X2=0.905 $Y2=1.51
r92 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=1.51 $X2=0.725 $Y2=1.51
r93 50 52 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.545 $Y=1.51
+ $X2=0.725 $Y2=1.51
r94 49 50 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.475 $Y=1.51
+ $X2=0.545 $Y2=1.51
r95 46 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.385 $Y=1.51
+ $X2=0.475 $Y2=1.51
r96 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.51 $X2=0.385 $Y2=1.51
r97 37 38 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=2.64 $Y2=1.592
r98 37 62 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=1.745 $Y2=1.592
r99 36 62 2.23608 $w=3.33e-07 $l=6.5e-08 $layer=LI1_cond $X=1.68 $Y=1.592
+ $X2=1.745 $Y2=1.592
r100 36 59 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=1.68 $Y=1.592
+ $X2=1.405 $Y2=1.592
r101 35 59 7.05226 $w=3.33e-07 $l=2.05e-07 $layer=LI1_cond $X=1.2 $Y=1.592
+ $X2=1.405 $Y2=1.592
r102 35 53 16.3406 $w=3.33e-07 $l=4.75e-07 $layer=LI1_cond $X=1.2 $Y=1.592
+ $X2=0.725 $Y2=1.592
r103 34 53 0.172006 $w=3.33e-07 $l=5e-09 $layer=LI1_cond $X=0.72 $Y=1.592
+ $X2=0.725 $Y2=1.592
r104 34 47 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=1.592
+ $X2=0.385 $Y2=1.592
r105 33 47 4.98819 $w=3.33e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.592
+ $X2=0.385 $Y2=1.592
r106 29 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.675
+ $X2=1.835 $Y2=1.51
r107 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.835 $Y=1.675
+ $X2=1.835 $Y2=2.465
r108 25 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=1.51
r109 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=0.765
r110 21 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.675
+ $X2=1.405 $Y2=1.51
r111 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.405 $Y=1.675
+ $X2=1.405 $Y2=2.465
r112 17 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.345
+ $X2=1.335 $Y2=1.51
r113 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.335 $Y=1.345
+ $X2=1.335 $Y2=0.765
r114 13 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.675
+ $X2=0.975 $Y2=1.51
r115 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.975 $Y=1.675
+ $X2=0.975 $Y2=2.465
r116 9 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=1.51
r117 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=0.765
r118 5 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.675
+ $X2=0.545 $Y2=1.51
r119 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.545 $Y=1.675
+ $X2=0.545 $Y2=2.465
r120 1 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=1.51
r121 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_4%A2 3 7 11 15 19 23 25 26 29 33 35 36 37 54
c90 33 0 6.59418e-20 $X=4.095 $Y=2.465
c91 26 0 8.70781e-20 $X=3.21 $Y=1.51
c92 19 0 8.15747e-20 $X=3.125 $Y=2.465
r93 52 54 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=3.775 $Y=1.51
+ $X2=4.095 $Y2=1.51
r94 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.775
+ $Y=1.51 $X2=3.775 $Y2=1.51
r95 50 52 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=3.645 $Y=1.51
+ $X2=3.775 $Y2=1.51
r96 48 49 1.51572 $w=3.18e-07 $l=1e-08 $layer=POLY_cond $X=3.125 $Y=1.51
+ $X2=3.135 $Y2=1.51
r97 46 48 4.54717 $w=3.18e-07 $l=3e-08 $layer=POLY_cond $X=3.095 $Y=1.51
+ $X2=3.125 $Y2=1.51
r98 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=1.51 $X2=3.095 $Y2=1.51
r99 44 46 60.6289 $w=3.18e-07 $l=4e-07 $layer=POLY_cond $X=2.695 $Y=1.51
+ $X2=3.095 $Y2=1.51
r100 43 44 10.6101 $w=3.18e-07 $l=7e-08 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.695 $Y2=1.51
r101 42 43 54.566 $w=3.18e-07 $l=3.6e-07 $layer=POLY_cond $X=2.265 $Y=1.51
+ $X2=2.625 $Y2=1.51
r102 41 42 10.6101 $w=3.18e-07 $l=7e-08 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.265 $Y2=1.51
r103 37 53 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=4.08 $Y=1.592
+ $X2=3.775 $Y2=1.592
r104 36 53 6.02022 $w=3.33e-07 $l=1.75e-07 $layer=LI1_cond $X=3.6 $Y=1.592
+ $X2=3.775 $Y2=1.592
r105 35 36 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.592
+ $X2=3.6 $Y2=1.592
r106 35 47 0.860032 $w=3.33e-07 $l=2.5e-08 $layer=LI1_cond $X=3.12 $Y=1.592
+ $X2=3.095 $Y2=1.592
r107 31 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.095 $Y=1.675
+ $X2=4.095 $Y2=1.51
r108 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.095 $Y=1.675
+ $X2=4.095 $Y2=2.465
r109 27 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.345
+ $X2=3.645 $Y2=1.51
r110 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.645 $Y=1.345
+ $X2=3.645 $Y2=0.765
r111 26 49 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.21 $Y=1.51
+ $X2=3.135 $Y2=1.51
r112 25 50 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.57 $Y=1.51
+ $X2=3.645 $Y2=1.51
r113 25 26 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.57 $Y=1.51
+ $X2=3.21 $Y2=1.51
r114 21 49 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.135 $Y=1.345
+ $X2=3.135 $Y2=1.51
r115 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.135 $Y=1.345
+ $X2=3.135 $Y2=0.765
r116 17 48 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.675
+ $X2=3.125 $Y2=1.51
r117 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.125 $Y=1.675
+ $X2=3.125 $Y2=2.465
r118 13 44 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.675
+ $X2=2.695 $Y2=1.51
r119 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.695 $Y=1.675
+ $X2=2.695 $Y2=2.465
r120 9 43 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=1.51
r121 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=0.765
r122 5 42 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.675
+ $X2=2.265 $Y2=1.51
r123 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.265 $Y=1.675
+ $X2=2.265 $Y2=2.465
r124 1 41 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=1.51
r125 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_4%A1 3 7 11 15 19 23 27 31 33 34 35 36 53
c88 53 0 1.39361e-19 $X=5.815 $Y=1.485
c89 23 0 5.49369e-20 $X=5.535 $Y=0.745
c90 15 0 2.06194e-19 $X=5.105 $Y=0.745
c91 7 0 5.39005e-20 $X=4.675 $Y=0.745
r92 53 54 20.1955 $w=3.58e-07 $l=1.5e-07 $layer=POLY_cond $X=5.815 $Y=1.485
+ $X2=5.965 $Y2=1.485
r93 51 53 2.01955 $w=3.58e-07 $l=1.5e-08 $layer=POLY_cond $X=5.8 $Y=1.485
+ $X2=5.815 $Y2=1.485
r94 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.8 $Y=1.51
+ $X2=5.8 $Y2=1.51
r95 49 51 35.6788 $w=3.58e-07 $l=2.65e-07 $layer=POLY_cond $X=5.535 $Y=1.485
+ $X2=5.8 $Y2=1.485
r96 48 49 20.1955 $w=3.58e-07 $l=1.5e-07 $layer=POLY_cond $X=5.385 $Y=1.485
+ $X2=5.535 $Y2=1.485
r97 46 48 35.6788 $w=3.58e-07 $l=2.65e-07 $layer=POLY_cond $X=5.12 $Y=1.485
+ $X2=5.385 $Y2=1.485
r98 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.51 $X2=5.12 $Y2=1.51
r99 44 46 2.01955 $w=3.58e-07 $l=1.5e-08 $layer=POLY_cond $X=5.105 $Y=1.485
+ $X2=5.12 $Y2=1.485
r100 43 44 20.1955 $w=3.58e-07 $l=1.5e-07 $layer=POLY_cond $X=4.955 $Y=1.485
+ $X2=5.105 $Y2=1.485
r101 42 43 37.6983 $w=3.58e-07 $l=2.8e-07 $layer=POLY_cond $X=4.675 $Y=1.485
+ $X2=4.955 $Y2=1.485
r102 35 36 15.5823 $w=3.53e-07 $l=4.8e-07 $layer=LI1_cond $X=6 $Y=1.602 $X2=6.48
+ $Y2=1.602
r103 35 52 6.49264 $w=3.53e-07 $l=2e-07 $layer=LI1_cond $X=6 $Y=1.602 $X2=5.8
+ $Y2=1.602
r104 34 52 9.08969 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=5.52 $Y=1.602
+ $X2=5.8 $Y2=1.602
r105 34 47 12.9853 $w=3.53e-07 $l=4e-07 $layer=LI1_cond $X=5.52 $Y=1.602
+ $X2=5.12 $Y2=1.602
r106 33 47 2.59705 $w=3.53e-07 $l=8e-08 $layer=LI1_cond $X=5.04 $Y=1.602
+ $X2=5.12 $Y2=1.602
r107 29 54 23.1716 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.965 $Y=1.295
+ $X2=5.965 $Y2=1.485
r108 29 31 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.965 $Y=1.295
+ $X2=5.965 $Y2=0.745
r109 25 53 23.1716 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.815 $Y2=1.485
r110 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.815 $Y2=2.465
r111 21 49 23.1716 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.535 $Y=1.295
+ $X2=5.535 $Y2=1.485
r112 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.535 $Y=1.295
+ $X2=5.535 $Y2=0.745
r113 17 48 23.1716 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=1.485
r114 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=2.465
r115 13 44 23.1716 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.105 $Y=1.295
+ $X2=5.105 $Y2=1.485
r116 13 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.105 $Y=1.295
+ $X2=5.105 $Y2=0.745
r117 9 43 23.1716 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=4.955 $Y2=1.485
r118 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=4.955 $Y2=2.465
r119 5 42 23.1716 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.675 $Y=1.295
+ $X2=4.675 $Y2=1.485
r120 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.675 $Y=1.295
+ $X2=4.675 $Y2=0.745
r121 1 42 20.1955 $w=3.58e-07 $l=2.54165e-07 $layer=POLY_cond $X=4.525 $Y=1.675
+ $X2=4.675 $Y2=1.485
r122 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.525 $Y=1.675
+ $X2=4.525 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_4%B1 3 7 11 15 19 23 27 31 33 34 35 51
c75 51 0 2.32723e-19 $X=7.615 $Y=1.515
r76 51 52 10.1934 $w=3.31e-07 $l=7e-08 $layer=POLY_cond $X=7.615 $Y=1.515
+ $X2=7.685 $Y2=1.515
r77 49 51 2.91239 $w=3.31e-07 $l=2e-08 $layer=POLY_cond $X=7.595 $Y=1.515
+ $X2=7.615 $Y2=1.515
r78 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.595
+ $Y=1.51 $X2=7.595 $Y2=1.51
r79 47 49 49.5106 $w=3.31e-07 $l=3.4e-07 $layer=POLY_cond $X=7.255 $Y=1.515
+ $X2=7.595 $Y2=1.515
r80 46 47 10.1934 $w=3.31e-07 $l=7e-08 $layer=POLY_cond $X=7.185 $Y=1.515
+ $X2=7.255 $Y2=1.515
r81 44 46 39.3172 $w=3.31e-07 $l=2.7e-07 $layer=POLY_cond $X=6.915 $Y=1.515
+ $X2=7.185 $Y2=1.515
r82 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.915
+ $Y=1.51 $X2=6.915 $Y2=1.51
r83 42 44 13.1057 $w=3.31e-07 $l=9e-08 $layer=POLY_cond $X=6.825 $Y=1.515
+ $X2=6.915 $Y2=1.515
r84 41 42 10.1934 $w=3.31e-07 $l=7e-08 $layer=POLY_cond $X=6.755 $Y=1.515
+ $X2=6.825 $Y2=1.515
r85 40 41 52.423 $w=3.31e-07 $l=3.6e-07 $layer=POLY_cond $X=6.395 $Y=1.515
+ $X2=6.755 $Y2=1.515
r86 39 40 10.1934 $w=3.31e-07 $l=7e-08 $layer=POLY_cond $X=6.325 $Y=1.515
+ $X2=6.395 $Y2=1.515
r87 35 50 10.5505 $w=3.53e-07 $l=3.25e-07 $layer=LI1_cond $X=7.92 $Y=1.602
+ $X2=7.595 $Y2=1.602
r88 34 50 5.03179 $w=3.53e-07 $l=1.55e-07 $layer=LI1_cond $X=7.44 $Y=1.602
+ $X2=7.595 $Y2=1.602
r89 33 34 15.5823 $w=3.53e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.602
+ $X2=7.44 $Y2=1.602
r90 33 45 1.46084 $w=3.53e-07 $l=4.5e-08 $layer=LI1_cond $X=6.96 $Y=1.602
+ $X2=6.915 $Y2=1.602
r91 29 52 21.295 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.685 $Y=1.345
+ $X2=7.685 $Y2=1.515
r92 29 31 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.685 $Y=1.345
+ $X2=7.685 $Y2=0.745
r93 25 51 21.295 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.615 $Y=1.685
+ $X2=7.615 $Y2=1.515
r94 25 27 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.615 $Y=1.685
+ $X2=7.615 $Y2=2.465
r95 21 47 21.295 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.255 $Y=1.345
+ $X2=7.255 $Y2=1.515
r96 21 23 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.255 $Y=1.345
+ $X2=7.255 $Y2=0.745
r97 17 46 21.295 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.185 $Y=1.685
+ $X2=7.185 $Y2=1.515
r98 17 19 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.185 $Y=1.685
+ $X2=7.185 $Y2=2.465
r99 13 42 21.295 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.825 $Y=1.345
+ $X2=6.825 $Y2=1.515
r100 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.825 $Y=1.345
+ $X2=6.825 $Y2=0.745
r101 9 41 21.295 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.755 $Y=1.685
+ $X2=6.755 $Y2=1.515
r102 9 11 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.755 $Y=1.685
+ $X2=6.755 $Y2=2.465
r103 5 40 21.295 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.395 $Y=1.345
+ $X2=6.395 $Y2=1.515
r104 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.395 $Y=1.345 $X2=6.395
+ $Y2=0.745
r105 1 39 21.295 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.325 $Y=1.685
+ $X2=6.325 $Y2=1.515
r106 1 3 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.325 $Y=1.685
+ $X2=6.325 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_4%A_41_367# 1 2 3 4 5 6 7 8 9 28 30 32 36 38
+ 42 44 48 50 53 54 56 60 62 64 65 68 70 72 74 79 81 83 88 90 93
c100 81 0 8.70781e-20 $X=2.05 $Y=2.095
c101 74 0 8.37457e-20 $X=7.83 $Y=2.115
c102 56 0 1.39361e-19 $X=5.075 $Y=2.375
r103 72 95 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=2.905
+ $X2=7.87 $Y2=2.99
r104 72 74 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=7.87 $Y=2.905
+ $X2=7.87 $Y2=2.115
r105 71 93 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.065 $Y=2.99
+ $X2=6.97 $Y2=2.99
r106 70 95 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.745 $Y=2.99
+ $X2=7.87 $Y2=2.99
r107 70 71 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.745 $Y=2.99
+ $X2=7.065 $Y2=2.99
r108 66 93 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=2.905
+ $X2=6.97 $Y2=2.99
r109 66 68 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=6.97 $Y=2.905
+ $X2=6.97 $Y2=2.455
r110 64 93 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.875 $Y=2.99
+ $X2=6.97 $Y2=2.99
r111 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.875 $Y=2.99
+ $X2=6.205 $Y2=2.99
r112 63 65 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=6.07 $Y=2.905
+ $X2=6.205 $Y2=2.99
r113 62 92 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=2.46
+ $X2=6.07 $Y2=2.375
r114 62 63 18.994 $w=2.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.07 $Y=2.46
+ $X2=6.07 $Y2=2.905
r115 61 90 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.265 $Y=2.375
+ $X2=5.17 $Y2=2.375
r116 60 92 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.935 $Y=2.375
+ $X2=6.07 $Y2=2.375
r117 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.935 $Y=2.375
+ $X2=5.265 $Y2=2.375
r118 56 90 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.075 $Y=2.375
+ $X2=5.17 $Y2=2.375
r119 56 88 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.075 $Y=2.375
+ $X2=4.405 $Y2=2.375
r120 54 88 6.82456 $w=1.78e-07 $l=1.1e-07 $layer=LI1_cond $X=4.295 $Y=2.38
+ $X2=4.405 $Y2=2.38
r121 54 84 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=4.295 $Y=2.38
+ $X2=4.1 $Y2=2.38
r122 53 84 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.1 $Y=2.29 $X2=4.1
+ $Y2=2.38
r123 52 53 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.1 $Y=2.1 $X2=4.1
+ $Y2=2.29
r124 51 83 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.005 $Y=2.015
+ $X2=2.91 $Y2=2.015
r125 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=2.015
+ $X2=4.1 $Y2=2.1
r126 50 51 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.015 $Y=2.015
+ $X2=3.005 $Y2=2.015
r127 46 83 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=2.1
+ $X2=2.91 $Y2=2.015
r128 46 48 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=2.91 $Y=2.1
+ $X2=2.91 $Y2=2.91
r129 45 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.145 $Y=2.015
+ $X2=2.05 $Y2=2.015
r130 44 83 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.815 $Y=2.015
+ $X2=2.91 $Y2=2.015
r131 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.815 $Y=2.015
+ $X2=2.145 $Y2=2.015
r132 40 81 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=2.1
+ $X2=2.05 $Y2=2.015
r133 40 42 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=2.05 $Y=2.1
+ $X2=2.05 $Y2=2.91
r134 39 79 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.285 $Y=2.015
+ $X2=1.19 $Y2=2.015
r135 38 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.955 $Y=2.015
+ $X2=2.05 $Y2=2.015
r136 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.955 $Y=2.015
+ $X2=1.285 $Y2=2.015
r137 34 79 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=2.1
+ $X2=1.19 $Y2=2.015
r138 34 36 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=1.19 $Y=2.1
+ $X2=1.19 $Y2=2.91
r139 33 77 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.425 $Y=2.015
+ $X2=0.295 $Y2=2.015
r140 32 79 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.095 $Y=2.015
+ $X2=1.19 $Y2=2.015
r141 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.095 $Y=2.015
+ $X2=0.425 $Y2=2.015
r142 28 77 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.295 $Y=2.1
+ $X2=0.295 $Y2=2.015
r143 28 30 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=0.295 $Y=2.1
+ $X2=0.295 $Y2=2.91
r144 9 95 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.69
+ $Y=1.835 $X2=7.83 $Y2=2.91
r145 9 74 400 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=7.69
+ $Y=1.835 $X2=7.83 $Y2=2.115
r146 8 68 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=6.83
+ $Y=1.835 $X2=6.97 $Y2=2.455
r147 7 92 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=5.89
+ $Y=1.835 $X2=6.03 $Y2=2.455
r148 6 90 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=5.03
+ $Y=1.835 $X2=5.17 $Y2=2.455
r149 5 54 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=4.17
+ $Y=1.835 $X2=4.31 $Y2=2.455
r150 4 83 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.835 $X2=2.91 $Y2=2.095
r151 4 48 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.835 $X2=2.91 $Y2=2.91
r152 3 81 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=2.095
r153 3 42 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=2.91
r154 2 79 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.095
r155 2 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.91
r156 1 77 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.095
r157 1 30 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 40 41 43 44
+ 45 47 52 61 69 78 79 82 85 92 95
r124 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r125 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r126 90 92 5.90573 $w=7.85e-07 $l=3.8e-07 $layer=LI1_cond $X=3.595 $Y=2.95
+ $X2=3.595 $Y2=3.33
r127 88 90 9.24713 $w=7.85e-07 $l=5.95e-07 $layer=LI1_cond $X=3.595 $Y=2.355
+ $X2=3.595 $Y2=2.95
r128 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 76 79 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r132 76 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r133 75 78 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.92
+ $Y2=3.33
r134 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r135 73 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.6 $Y2=3.33
r136 73 75 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=6 $Y2=3.33
r137 72 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r138 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r139 69 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.6 $Y2=3.33
r140 69 71 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.04 $Y2=3.33
r141 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r142 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 65 92 10.0822 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=3.595 $Y2=3.33
r144 65 67 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=4.56 $Y2=3.33
r145 64 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r146 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r147 61 92 10.0822 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.595 $Y2=3.33
r148 61 63 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.12 $Y2=3.33
r149 60 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r150 60 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r151 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r152 57 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.62 $Y2=3.33
r153 57 59 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=2.16 $Y2=3.33
r154 56 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r155 56 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r156 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r157 53 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.76 $Y2=3.33
r158 53 55 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.2 $Y2=3.33
r159 52 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=3.33
+ $X2=1.62 $Y2=3.33
r160 52 55 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.455 $Y=3.33
+ $X2=1.2 $Y2=3.33
r161 50 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r162 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r163 47 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.76 $Y2=3.33
r164 47 49 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.24 $Y2=3.33
r165 45 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r166 45 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r167 43 67 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.56 $Y2=3.33
r168 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.74 $Y2=3.33
r169 42 71 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=5.04 $Y2=3.33
r170 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=4.74 $Y2=3.33
r171 40 59 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.16 $Y2=3.33
r172 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.48 $Y2=3.33
r173 39 63 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=3.12 $Y2=3.33
r174 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.48 $Y2=3.33
r175 35 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.6 $Y=3.245 $X2=5.6
+ $Y2=3.33
r176 35 37 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.6 $Y=3.245
+ $X2=5.6 $Y2=2.75
r177 31 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.74 $Y=3.245
+ $X2=4.74 $Y2=3.33
r178 31 33 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.74 $Y=3.245
+ $X2=4.74 $Y2=2.75
r179 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=3.245
+ $X2=2.48 $Y2=3.33
r180 27 29 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=2.48 $Y=3.245
+ $X2=2.48 $Y2=2.395
r181 23 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=3.245
+ $X2=1.62 $Y2=3.33
r182 23 25 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=1.62 $Y=3.245
+ $X2=1.62 $Y2=2.395
r183 19 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=3.33
r184 19 21 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=2.395
r185 6 37 600 $w=1.7e-07 $l=9.8251e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.75
r186 5 33 600 $w=1.7e-07 $l=9.8251e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.835 $X2=4.74 $Y2=2.75
r187 4 90 300 $w=1.7e-07 $l=1.41472e-06 $layer=licon1_PDIFF $count=2 $X=3.2
+ $Y=1.835 $X2=3.88 $Y2=2.95
r188 4 88 300 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=2 $X=3.2
+ $Y=1.835 $X2=3.34 $Y2=2.355
r189 3 29 300 $w=1.7e-07 $l=6.26099e-07 $layer=licon1_PDIFF $count=2 $X=2.34
+ $Y=1.835 $X2=2.48 $Y2=2.395
r190 2 25 300 $w=1.7e-07 $l=6.26099e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=2.395
r191 1 21 300 $w=1.7e-07 $l=6.26099e-07 $layer=licon1_PDIFF $count=2 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_4%Y 1 2 3 4 5 6 7 22 24 26 30 32 36 40 42 48
+ 51 56 58 59 61 62 64 65 72 75
c128 75 0 6.59418e-20 $X=4.56 $Y=1.295
c129 56 0 1.48977e-19 $X=6.175 $Y=1.152
c130 26 0 5.44556e-20 $X=6.075 $Y=1.152
c131 22 0 5.49369e-20 $X=5.155 $Y=1.047
r132 72 75 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=4.53 $Y=1.255
+ $X2=4.53 $Y2=1.295
r133 64 65 7.83892 $w=5.18e-07 $l=2.85e-07 $layer=LI1_cond $X=4.53 $Y=1.665
+ $X2=4.53 $Y2=1.95
r134 62 72 3.73677 $w=3.5e-07 $l=2.08e-07 $layer=LI1_cond $X=4.53 $Y=1.047
+ $X2=4.53 $Y2=1.255
r135 62 64 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=4.53 $Y=1.317
+ $X2=4.53 $Y2=1.665
r136 62 75 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=4.53 $Y=1.317
+ $X2=4.53 $Y2=1.295
r137 46 48 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=7.94 $Y=1.075
+ $X2=7.94 $Y2=0.47
r138 43 59 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=7.135 $Y=1.165
+ $X2=7.04 $Y2=1.165
r139 42 46 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=7.815 $Y=1.165
+ $X2=7.94 $Y2=1.075
r140 42 43 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=1.165
+ $X2=7.135 $Y2=1.165
r141 38 59 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=7.04 $Y=1.075 $X2=7.04
+ $Y2=1.165
r142 38 40 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=7.04 $Y=1.075
+ $X2=7.04 $Y2=0.45
r143 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.705 $Y=2.035
+ $X2=6.54 $Y2=2.035
r144 36 61 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.235 $Y=2.035
+ $X2=7.4 $Y2=2.035
r145 36 37 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.235 $Y=2.035
+ $X2=6.705 $Y2=2.035
r146 33 56 5.33237 $w=1.92e-07 $l=1.06301e-07 $layer=LI1_cond $X=6.275 $Y=1.165
+ $X2=6.175 $Y2=1.152
r147 32 59 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.945 $Y=1.165
+ $X2=7.04 $Y2=1.165
r148 32 33 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=6.945 $Y=1.165
+ $X2=6.275 $Y2=1.165
r149 28 56 1.20529 $w=2e-07 $l=1.02e-07 $layer=LI1_cond $X=6.175 $Y=1.05
+ $X2=6.175 $Y2=1.152
r150 28 30 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=6.175 $Y=1.05
+ $X2=6.175 $Y2=0.45
r151 27 54 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=5.485 $Y=1.152
+ $X2=5.32 $Y2=1.152
r152 26 56 5.33237 $w=1.92e-07 $l=1e-07 $layer=LI1_cond $X=6.075 $Y=1.152
+ $X2=6.175 $Y2=1.152
r153 26 27 31.9202 $w=2.03e-07 $l=5.9e-07 $layer=LI1_cond $X=6.075 $Y=1.152
+ $X2=5.485 $Y2=1.152
r154 25 65 5.34211 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.705 $Y=2.035
+ $X2=4.53 $Y2=2.035
r155 24 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=2.035
+ $X2=6.54 $Y2=2.035
r156 24 25 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=6.375 $Y=2.035
+ $X2=4.705 $Y2=2.035
r157 23 62 3.14392 $w=4.15e-07 $l=1.75e-07 $layer=LI1_cond $X=4.705 $Y=1.047
+ $X2=4.53 $Y2=1.047
r158 22 54 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=5.32 $Y=1.047
+ $X2=5.32 $Y2=1.152
r159 22 51 12.8166 $w=3.28e-07 $l=3.67e-07 $layer=LI1_cond $X=5.32 $Y=1.047
+ $X2=5.32 $Y2=0.68
r160 22 23 12.4964 $w=4.13e-07 $l=4.5e-07 $layer=LI1_cond $X=5.155 $Y=1.047
+ $X2=4.705 $Y2=1.047
r161 7 61 300 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=2 $X=7.26
+ $Y=1.835 $X2=7.4 $Y2=2.115
r162 6 58 300 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=2 $X=6.4
+ $Y=1.835 $X2=6.54 $Y2=2.115
r163 5 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.76
+ $Y=0.325 $X2=7.9 $Y2=0.47
r164 4 40 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.9
+ $Y=0.325 $X2=7.04 $Y2=0.45
r165 3 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.04
+ $Y=0.325 $X2=6.18 $Y2=0.45
r166 2 51 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=5.18
+ $Y=0.325 $X2=5.32 $Y2=0.68
r167 1 62 182 $w=1.7e-07 $l=7.39865e-07 $layer=licon1_NDIFF $count=1 $X=4.335
+ $Y=0.325 $X2=4.46 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_4%A_27_69# 1 2 3 4 5 18 20 21 24 26 30 32 36
+ 38 42 44 45 46
r79 40 42 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.94 $Y=1.085
+ $X2=3.94 $Y2=0.69
r80 39 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=1.17
+ $X2=2.92 $Y2=1.17
r81 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.775 $Y=1.17
+ $X2=3.94 $Y2=1.085
r82 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.775 $Y=1.17
+ $X2=3.085 $Y2=1.17
r83 34 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=1.085
+ $X2=2.92 $Y2=1.17
r84 34 36 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.92 $Y=1.085
+ $X2=2.92 $Y2=0.69
r85 33 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.075 $Y=1.17
+ $X2=1.98 $Y2=1.17
r86 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=1.17
+ $X2=2.92 $Y2=1.17
r87 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.755 $Y=1.17
+ $X2=2.075 $Y2=1.17
r88 28 45 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=1.085
+ $X2=1.98 $Y2=1.17
r89 28 30 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=1.98 $Y=1.085
+ $X2=1.98 $Y2=0.49
r90 27 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.215 $Y=1.17
+ $X2=1.12 $Y2=1.17
r91 26 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.885 $Y=1.17
+ $X2=1.98 $Y2=1.17
r92 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.885 $Y=1.17
+ $X2=1.215 $Y2=1.17
r93 22 44 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.085
+ $X2=1.12 $Y2=1.17
r94 22 24 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=1.12 $Y=1.085
+ $X2=1.12 $Y2=0.49
r95 20 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.025 $Y=1.17
+ $X2=1.12 $Y2=1.17
r96 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.025 $Y=1.17
+ $X2=0.345 $Y2=1.17
r97 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=1.085
+ $X2=0.345 $Y2=1.17
r98 16 18 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=0.22 $Y=1.085
+ $X2=0.22 $Y2=0.49
r99 5 42 91 $w=1.7e-07 $l=4.41503e-07 $layer=licon1_NDIFF $count=2 $X=3.72
+ $Y=0.345 $X2=3.94 $Y2=0.69
r100 4 36 91 $w=1.7e-07 $l=4.41503e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.345 $X2=2.92 $Y2=0.69
r101 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.345 $X2=1.98 $Y2=0.49
r102 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.345 $X2=1.12 $Y2=0.49
r103 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.345 $X2=0.26 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_4%VGND 1 2 3 4 15 19 21 25 29 31 33 38 43 50
+ 51 54 57 60 63
r103 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r104 60 61 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r105 57 58 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r106 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r107 51 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r108 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r109 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.635 $Y=0 $X2=7.47
+ $Y2=0
r110 48 50 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.635 $Y=0
+ $X2=7.92 $Y2=0
r111 47 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r112 47 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r113 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r114 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.61
+ $Y2=0
r115 44 46 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.775 $Y=0
+ $X2=6.96 $Y2=0
r116 43 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=0 $X2=7.47
+ $Y2=0
r117 43 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.305 $Y=0 $X2=6.96
+ $Y2=0
r118 42 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r119 42 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r120 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r121 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r122 39 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r123 38 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.55
+ $Y2=0
r124 38 41 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.2
+ $Y2=0
r125 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r126 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r127 33 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r128 33 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.24 $Y2=0
r129 31 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6.48
+ $Y2=0
r130 31 58 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=1.68
+ $Y2=0
r131 27 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=0.085
+ $X2=7.47 $Y2=0
r132 27 29 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.47 $Y=0.085
+ $X2=7.47 $Y2=0.45
r133 23 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0
r134 23 25 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0.45
r135 22 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=0 $X2=1.55
+ $Y2=0
r136 21 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.61
+ $Y2=0
r137 21 22 308.588 $w=1.68e-07 $l=4.73e-06 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=1.715 $Y2=0
r138 17 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0
r139 17 19 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0.47
r140 13 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r141 13 15 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.47
r142 4 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.33
+ $Y=0.325 $X2=7.47 $Y2=0.45
r143 3 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.47
+ $Y=0.325 $X2=6.61 $Y2=0.45
r144 2 19 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.345 $X2=1.55 $Y2=0.47
r145 1 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.345 $X2=0.69 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_4%A_454_69# 1 2 3 4 15 17 18 21 23 25 29 31 32
c61 32 0 1.51739e-19 $X=4.855 $Y=0.34
c62 25 0 5.39005e-20 $X=5.655 $Y=0.34
r63 32 35 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=0.34
+ $X2=4.855 $Y2=0.505
r64 27 29 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=5.755 $Y=0.425
+ $X2=5.755 $Y2=0.715
r65 26 32 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.985 $Y=0.34
+ $X2=4.855 $Y2=0.34
r66 25 27 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.655 $Y=0.34
+ $X2=5.755 $Y2=0.425
r67 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.655 $Y=0.34
+ $X2=4.985 $Y2=0.34
r68 24 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0.34
+ $X2=3.43 $Y2=0.34
r69 23 32 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.725 $Y=0.34
+ $X2=4.855 $Y2=0.34
r70 23 24 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=4.725 $Y=0.34
+ $X2=3.595 $Y2=0.34
r71 19 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=0.425
+ $X2=3.43 $Y2=0.34
r72 19 21 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.43 $Y=0.425
+ $X2=3.43 $Y2=0.47
r73 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=0.34
+ $X2=3.43 $Y2=0.34
r74 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.265 $Y=0.34
+ $X2=2.575 $Y2=0.34
r75 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.41 $Y=0.425
+ $X2=2.575 $Y2=0.34
r76 13 15 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.41 $Y=0.425
+ $X2=2.41 $Y2=0.47
r77 4 29 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.325 $X2=5.75 $Y2=0.715
r78 3 35 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.75 $Y=0.325
+ $X2=4.89 $Y2=0.505
r79 2 21 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=3.21
+ $Y=0.345 $X2=3.43 $Y2=0.47
r80 1 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.345 $X2=2.41 $Y2=0.47
.ends

