* File: sky130_fd_sc_lp__a21oi_4.pex.spice
* Created: Wed Sep  2 09:20:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21OI_4%A2 3 7 11 15 19 23 27 31 34 35 38 40 41 42
+ 43 61 66
c110 34 0 1.17145e-19 $X=3.51 $Y=1.51
c111 31 0 9.49247e-20 $X=3.53 $Y=2.465
r112 60 66 7.58926 $w=4.08e-07 $l=2.7e-07 $layer=LI1_cond $X=1.29 $Y=1.58
+ $X2=1.56 $Y2=1.58
r113 59 61 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.29 $Y=1.46 $X2=1.34
+ $Y2=1.46
r114 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.29
+ $Y=1.46 $X2=1.29 $Y2=1.46
r115 57 59 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=0.91 $Y=1.46
+ $X2=1.29 $Y2=1.46
r116 55 57 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=0.61 $Y=1.46 $X2=0.91
+ $Y2=1.46
r117 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.46 $X2=0.61 $Y2=1.46
r118 53 55 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=0.48 $Y=1.46
+ $X2=0.61 $Y2=1.46
r119 51 56 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=0.27 $Y=1.58
+ $X2=0.61 $Y2=1.58
r120 50 53 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.48 $Y2=1.46
r121 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.46 $X2=0.27 $Y2=1.46
r122 43 66 3.373 $w=4.08e-07 $l=1.2e-07 $layer=LI1_cond $X=1.68 $Y=1.58 $X2=1.56
+ $Y2=1.58
r123 42 60 2.52975 $w=4.08e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.58 $X2=1.29
+ $Y2=1.58
r124 41 42 13.492 $w=4.08e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.58 $X2=1.2
+ $Y2=1.58
r125 41 56 3.09192 $w=4.08e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.58
+ $X2=0.61 $Y2=1.58
r126 40 51 0.843251 $w=4.08e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=1.58
+ $X2=0.27 $Y2=1.58
r127 38 43 63.0764 $w=3.03e-07 $l=1.635e-06 $layer=LI1_cond $X=3.4 $Y=1.7
+ $X2=1.765 $Y2=1.7
r128 35 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=1.51
+ $X2=3.51 $Y2=1.675
r129 35 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=1.51
+ $X2=3.51 $Y2=1.345
r130 34 38 7.96233 $w=2.73e-07 $l=1.9e-07 $layer=LI1_cond $X=3.537 $Y=1.51
+ $X2=3.537 $Y2=1.7
r131 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.51
+ $Y=1.51 $X2=3.51 $Y2=1.51
r132 31 65 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.53 $Y=2.465
+ $X2=3.53 $Y2=1.675
r133 27 64 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.49 $Y=0.655
+ $X2=3.49 $Y2=1.345
r134 21 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.625
+ $X2=1.34 $Y2=1.46
r135 21 23 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.34 $Y=1.625
+ $X2=1.34 $Y2=2.465
r136 17 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.295
+ $X2=1.34 $Y2=1.46
r137 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.34 $Y=1.295
+ $X2=1.34 $Y2=0.655
r138 13 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.625
+ $X2=0.91 $Y2=1.46
r139 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.91 $Y=1.625
+ $X2=0.91 $Y2=2.465
r140 9 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.295
+ $X2=0.91 $Y2=1.46
r141 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.91 $Y=1.295
+ $X2=0.91 $Y2=0.655
r142 5 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.625
+ $X2=0.48 $Y2=1.46
r143 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.48 $Y=1.625
+ $X2=0.48 $Y2=2.465
r144 1 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.295
+ $X2=0.48 $Y2=1.46
r145 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.48 $Y=1.295 $X2=0.48
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 45
c77 27 0 1.17145e-19 $X=3.06 $Y=2.465
r78 43 45 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=2.82 $Y=1.35
+ $X2=3.06 $Y2=1.35
r79 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.35 $X2=2.82 $Y2=1.35
r80 41 43 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.63 $Y=1.35
+ $X2=2.82 $Y2=1.35
r81 40 41 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.2 $Y=1.35 $X2=2.63
+ $Y2=1.35
r82 38 40 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.14 $Y=1.35 $X2=2.2
+ $Y2=1.35
r83 35 38 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=1.77 $Y=1.35
+ $X2=2.14 $Y2=1.35
r84 31 44 14.712 $w=2.33e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.317 $X2=2.82
+ $Y2=1.317
r85 30 44 8.82722 $w=2.33e-07 $l=1.8e-07 $layer=LI1_cond $X=2.64 $Y=1.317
+ $X2=2.82 $Y2=1.317
r86 29 30 24.5201 $w=2.33e-07 $l=5e-07 $layer=LI1_cond $X=2.14 $Y=1.317 $X2=2.64
+ $Y2=1.317
r87 29 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.35 $X2=2.14 $Y2=1.35
r88 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.515
+ $X2=3.06 $Y2=1.35
r89 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.06 $Y=1.515
+ $X2=3.06 $Y2=2.465
r90 22 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.185
+ $X2=3.06 $Y2=1.35
r91 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.06 $Y=1.185
+ $X2=3.06 $Y2=0.655
r92 18 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.63 $Y=1.515
+ $X2=2.63 $Y2=1.35
r93 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.63 $Y=1.515
+ $X2=2.63 $Y2=2.465
r94 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.63 $Y=1.185
+ $X2=2.63 $Y2=1.35
r95 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.63 $Y=1.185
+ $X2=2.63 $Y2=0.655
r96 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.515
+ $X2=2.2 $Y2=1.35
r97 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.2 $Y=1.515 $X2=2.2
+ $Y2=2.465
r98 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.185 $X2=2.2
+ $Y2=1.35
r99 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.2 $Y=1.185 $X2=2.2
+ $Y2=0.655
r100 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.515
+ $X2=1.77 $Y2=1.35
r101 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.77 $Y=1.515
+ $X2=1.77 $Y2=2.465
r102 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.185
+ $X2=1.77 $Y2=1.35
r103 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.77 $Y=1.185
+ $X2=1.77 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_4%B1 3 7 11 15 19 23 27 31 33 34 35 50 51
c75 50 0 9.49247e-20 $X=5.07 $Y=1.51
r76 49 51 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.07 $Y=1.51 $X2=5.25
+ $Y2=1.51
r77 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.07
+ $Y=1.51 $X2=5.07 $Y2=1.51
r78 47 49 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=4.82 $Y=1.51
+ $X2=5.07 $Y2=1.51
r79 45 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.73 $Y=1.51 $X2=4.82
+ $Y2=1.51
r80 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.73
+ $Y=1.51 $X2=4.73 $Y2=1.51
r81 42 45 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.39 $Y=1.51
+ $X2=4.73 $Y2=1.51
r82 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.39
+ $Y=1.51 $X2=4.39 $Y2=1.51
r83 39 42 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.96 $Y=1.51
+ $X2=4.39 $Y2=1.51
r84 35 50 1.03204 $w=3.33e-07 $l=3e-08 $layer=LI1_cond $X=5.04 $Y=1.592 $X2=5.07
+ $Y2=1.592
r85 35 46 10.6644 $w=3.33e-07 $l=3.1e-07 $layer=LI1_cond $X=5.04 $Y=1.592
+ $X2=4.73 $Y2=1.592
r86 34 46 5.84822 $w=3.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.56 $Y=1.592
+ $X2=4.73 $Y2=1.592
r87 34 43 5.84822 $w=3.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.56 $Y=1.592
+ $X2=4.39 $Y2=1.592
r88 33 43 10.6644 $w=3.33e-07 $l=3.1e-07 $layer=LI1_cond $X=4.08 $Y=1.592
+ $X2=4.39 $Y2=1.592
r89 29 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.25 $Y=1.675
+ $X2=5.25 $Y2=1.51
r90 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.25 $Y=1.675
+ $X2=5.25 $Y2=2.465
r91 25 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.25 $Y=1.345
+ $X2=5.25 $Y2=1.51
r92 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.25 $Y=1.345
+ $X2=5.25 $Y2=0.655
r93 21 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.82 $Y=1.675
+ $X2=4.82 $Y2=1.51
r94 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.82 $Y=1.675
+ $X2=4.82 $Y2=2.465
r95 17 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.82 $Y=1.345
+ $X2=4.82 $Y2=1.51
r96 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.82 $Y=1.345
+ $X2=4.82 $Y2=0.655
r97 13 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.39 $Y=1.675
+ $X2=4.39 $Y2=1.51
r98 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.39 $Y=1.675
+ $X2=4.39 $Y2=2.465
r99 9 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.39 $Y=1.345
+ $X2=4.39 $Y2=1.51
r100 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.39 $Y=1.345
+ $X2=4.39 $Y2=0.655
r101 5 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.96 $Y=1.675
+ $X2=3.96 $Y2=1.51
r102 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.96 $Y=1.675
+ $X2=3.96 $Y2=2.465
r103 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.96 $Y=1.345
+ $X2=3.96 $Y2=1.51
r104 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.96 $Y=1.345
+ $X2=3.96 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_4%A_28_367# 1 2 3 4 5 6 7 22 24 26 30 32 36 38
+ 42 44 46 47 48 52 54 58 63 65 67 72
r71 56 58 16.4365 $w=3.03e-07 $l=4.35e-07 $layer=LI1_cond $X=5.477 $Y=2.905
+ $X2=5.477 $Y2=2.47
r72 55 72 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=4.74 $Y=2.99
+ $X2=4.602 $Y2=2.99
r73 54 56 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=5.325 $Y=2.99
+ $X2=5.477 $Y2=2.905
r74 54 55 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.325 $Y=2.99
+ $X2=4.74 $Y2=2.99
r75 50 72 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.602 $Y=2.905
+ $X2=4.602 $Y2=2.99
r76 50 52 18.2296 $w=2.73e-07 $l=4.35e-07 $layer=LI1_cond $X=4.602 $Y=2.905
+ $X2=4.602 $Y2=2.47
r77 49 71 4.53113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=3.885 $Y=2.99
+ $X2=3.747 $Y2=2.99
r78 48 72 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.465 $Y=2.99
+ $X2=4.602 $Y2=2.99
r79 48 49 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.465 $Y=2.99
+ $X2=3.885 $Y2=2.99
r80 47 71 2.79091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=3.747 $Y=2.905
+ $X2=3.747 $Y2=2.99
r81 46 69 2.80348 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=3.747 $Y=2.125
+ $X2=3.747 $Y2=2.04
r82 46 47 32.6875 $w=2.73e-07 $l=7.8e-07 $layer=LI1_cond $X=3.747 $Y=2.125
+ $X2=3.747 $Y2=2.905
r83 45 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.94 $Y=2.04
+ $X2=2.845 $Y2=2.04
r84 44 69 4.51856 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=3.61 $Y=2.04
+ $X2=3.747 $Y2=2.04
r85 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.61 $Y=2.04
+ $X2=2.94 $Y2=2.04
r86 40 67 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=2.125
+ $X2=2.845 $Y2=2.04
r87 40 42 45.823 $w=1.88e-07 $l=7.85e-07 $layer=LI1_cond $X=2.845 $Y=2.125
+ $X2=2.845 $Y2=2.91
r88 39 65 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.08 $Y=2.04 $X2=1.99
+ $Y2=2.04
r89 38 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.75 $Y=2.04
+ $X2=2.845 $Y2=2.04
r90 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.75 $Y=2.04
+ $X2=2.08 $Y2=2.04
r91 34 65 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=2.125
+ $X2=1.99 $Y2=2.04
r92 34 36 48.3687 $w=1.78e-07 $l=7.85e-07 $layer=LI1_cond $X=1.99 $Y=2.125
+ $X2=1.99 $Y2=2.91
r93 33 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.22 $Y=2.04
+ $X2=1.125 $Y2=2.04
r94 32 65 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.9 $Y=2.04 $X2=1.99
+ $Y2=2.04
r95 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.9 $Y=2.04 $X2=1.22
+ $Y2=2.04
r96 28 63 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=2.125
+ $X2=1.125 $Y2=2.04
r97 28 30 45.823 $w=1.88e-07 $l=7.85e-07 $layer=LI1_cond $X=1.125 $Y=2.125
+ $X2=1.125 $Y2=2.91
r98 27 61 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.36 $Y=2.04 $X2=0.23
+ $Y2=2.04
r99 26 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.03 $Y=2.04
+ $X2=1.125 $Y2=2.04
r100 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.03 $Y=2.04
+ $X2=0.36 $Y2=2.04
r101 22 61 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=2.125
+ $X2=0.23 $Y2=2.04
r102 22 24 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=0.23 $Y=2.125
+ $X2=0.23 $Y2=2.91
r103 7 58 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=5.325
+ $Y=1.835 $X2=5.465 $Y2=2.47
r104 6 52 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=4.465
+ $Y=1.835 $X2=4.605 $Y2=2.47
r105 5 71 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.605
+ $Y=1.835 $X2=3.745 $Y2=2.91
r106 5 69 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=3.605
+ $Y=1.835 $X2=3.745 $Y2=2.12
r107 4 67 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.835 $X2=2.845 $Y2=2.12
r108 4 42 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.835 $X2=2.845 $Y2=2.91
r109 3 65 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.835 $X2=1.985 $Y2=2.12
r110 3 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.835 $X2=1.985 $Y2=2.91
r111 2 63 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.12
r112 2 30 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.91
r113 1 61 400 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.12
r114 1 24 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_4%VPWR 1 2 3 4 15 19 23 25 29 32 33 34 35 36
+ 38 55 56 59 62
r86 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r87 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r88 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r89 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 53 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r91 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r92 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r93 50 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.44 $Y=3.33
+ $X2=3.275 $Y2=3.33
r94 50 52 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.44 $Y=3.33 $X2=3.6
+ $Y2=3.33
r95 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r96 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r97 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r99 43 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=3.33
+ $X2=0.695 $Y2=3.33
r100 43 45 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.86 $Y=3.33
+ $X2=1.2 $Y2=3.33
r101 41 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r103 38 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.695 $Y2=3.33
r104 38 40 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 36 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 36 49 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r107 34 48 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.25 $Y=3.33 $X2=2.16
+ $Y2=3.33
r108 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=2.415 $Y2=3.33
r109 32 45 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.555 $Y2=3.33
r111 31 48 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r112 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=1.555 $Y2=3.33
r113 27 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=3.245
+ $X2=3.275 $Y2=3.33
r114 27 29 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=3.275 $Y=3.245
+ $X2=3.275 $Y2=2.41
r115 26 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=3.33
+ $X2=2.415 $Y2=3.33
r116 25 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=3.33
+ $X2=3.275 $Y2=3.33
r117 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.11 $Y=3.33
+ $X2=2.58 $Y2=3.33
r118 21 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=3.245
+ $X2=2.415 $Y2=3.33
r119 21 23 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=2.415 $Y=3.245
+ $X2=2.415 $Y2=2.41
r120 17 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=3.245
+ $X2=1.555 $Y2=3.33
r121 17 19 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=1.555 $Y=3.245
+ $X2=1.555 $Y2=2.41
r122 13 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=3.33
r123 13 15 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=2.41
r124 4 29 300 $w=1.7e-07 $l=6.4119e-07 $layer=licon1_PDIFF $count=2 $X=3.135
+ $Y=1.835 $X2=3.275 $Y2=2.41
r125 3 23 300 $w=1.7e-07 $l=6.4119e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=1.835 $X2=2.415 $Y2=2.41
r126 2 19 300 $w=1.7e-07 $l=6.4119e-07 $layer=licon1_PDIFF $count=2 $X=1.415
+ $Y=1.835 $X2=1.555 $Y2=2.41
r127 1 15 300 $w=1.7e-07 $l=6.4119e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.835 $X2=0.695 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_4%Y 1 2 3 4 5 6 23 25 27 33 35 37 40 42 44 45
+ 46 47 48 49 50 57
c73 33 0 1.4697e-19 $X=5.035 $Y=0.42
r74 50 75 15.4072 $w=1.94e-07 $l=2.45e-07 $layer=LI1_cond $X=4.16 $Y=0.925
+ $X2=4.16 $Y2=1.17
r75 50 57 0.227314 $w=2.1e-07 $l=1e-07 $layer=LI1_cond $X=4.16 $Y=0.925 $X2=4.06
+ $Y2=0.925
r76 50 57 1.74286 $w=2.08e-07 $l=3.3e-08 $layer=LI1_cond $X=4.027 $Y=0.925
+ $X2=4.06 $Y2=0.925
r77 49 50 22.5515 $w=2.08e-07 $l=4.27e-07 $layer=LI1_cond $X=3.6 $Y=0.925
+ $X2=4.027 $Y2=0.925
r78 48 49 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=0.925
+ $X2=3.6 $Y2=0.925
r79 48 66 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=3.12 $Y=0.925
+ $X2=2.845 $Y2=0.925
r80 47 66 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=2.64 $Y=0.925
+ $X2=2.845 $Y2=0.925
r81 46 47 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=2.64 $Y2=0.925
r82 46 59 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=1.985 $Y2=0.925
r83 39 40 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.5 $Y=1.255
+ $X2=5.5 $Y2=1.93
r84 38 44 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=5.155 $Y=2.015
+ $X2=5.032 $Y2=2.015
r85 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=2.015
+ $X2=5.5 $Y2=1.93
r86 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.415 $Y=2.015
+ $X2=5.155 $Y2=2.015
r87 36 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.13 $Y=1.17
+ $X2=5.035 $Y2=1.17
r88 35 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=1.17
+ $X2=5.5 $Y2=1.255
r89 35 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.415 $Y=1.17
+ $X2=5.13 $Y2=1.17
r90 31 45 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.035 $Y=1.085
+ $X2=5.035 $Y2=1.17
r91 31 33 38.8182 $w=1.88e-07 $l=6.65e-07 $layer=LI1_cond $X=5.035 $Y=1.085
+ $X2=5.035 $Y2=0.42
r92 28 42 4.1433 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.295 $Y=2.015
+ $X2=4.175 $Y2=2.015
r93 27 44 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=4.91 $Y=2.015
+ $X2=5.032 $Y2=2.015
r94 27 28 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.91 $Y=2.015
+ $X2=4.295 $Y2=2.015
r95 26 75 1.50975 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.26 $Y=1.17 $X2=4.16
+ $Y2=1.17
r96 25 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.94 $Y=1.17
+ $X2=5.035 $Y2=1.17
r97 25 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.94 $Y=1.17
+ $X2=4.26 $Y2=1.17
r98 21 50 6.405 $w=2e-07 $l=1.05e-07 $layer=LI1_cond $X=4.16 $Y=0.82 $X2=4.16
+ $Y2=0.925
r99 21 23 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=4.16 $Y=0.82 $X2=4.16
+ $Y2=0.42
r100 6 44 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=4.895
+ $Y=1.835 $X2=5.035 $Y2=2.095
r101 5 42 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=1.835 $X2=4.175 $Y2=2.095
r102 4 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.895
+ $Y=0.235 $X2=5.035 $Y2=0.42
r103 3 50 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=4.035
+ $Y=0.235 $X2=4.175 $Y2=0.93
r104 3 23 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.035
+ $Y=0.235 $X2=4.175 $Y2=0.42
r105 2 66 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=2.705
+ $Y=0.235 $X2=2.845 $Y2=0.925
r106 1 59 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.235 $X2=1.985 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_4%VGND 1 2 3 4 5 16 18 22 26 30 32 34 36 38 43
+ 48 53 62 65 68 72
r82 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r83 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r84 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r85 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r86 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r87 57 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r88 57 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r89 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r90 54 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.77 $Y=0 $X2=4.605
+ $Y2=0
r91 54 56 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.77 $Y=0 $X2=5.04
+ $Y2=0
r92 53 71 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.53
+ $Y2=0
r93 53 56 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.04
+ $Y2=0
r94 52 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r95 52 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r96 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r97 49 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=3.725
+ $Y2=0
r98 49 51 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.08
+ $Y2=0
r99 48 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.605
+ $Y2=0
r100 48 51 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.08
+ $Y2=0
r101 47 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r102 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r103 44 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.125
+ $Y2=0
r104 44 46 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.68
+ $Y2=0
r105 43 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=0 $X2=3.725
+ $Y2=0
r106 43 46 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=3.56 $Y=0 $X2=1.68
+ $Y2=0
r107 42 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r108 42 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r109 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r110 39 59 4.39509 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r111 39 41 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.72
+ $Y2=0
r112 38 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.125
+ $Y2=0
r113 38 41 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r114 36 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r115 36 47 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.68
+ $Y2=0
r116 32 71 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=5.465 $Y=0.085
+ $X2=5.53 $Y2=0
r117 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.465 $Y=0.085
+ $X2=5.465 $Y2=0.38
r118 28 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.605 $Y=0.085
+ $X2=4.605 $Y2=0
r119 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.605 $Y=0.085
+ $X2=4.605 $Y2=0.38
r120 24 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0
r121 24 26 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0.525
r122 20 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0
r123 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0.38
r124 16 59 3.04275 $w=2.9e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.195 $Y2=0
r125 16 18 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.245 $Y2=0.38
r126 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.325
+ $Y=0.235 $X2=5.465 $Y2=0.38
r127 4 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.465
+ $Y=0.235 $X2=4.605 $Y2=0.38
r128 3 26 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=3.565
+ $Y=0.235 $X2=3.725 $Y2=0.525
r129 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.235 $X2=1.125 $Y2=0.38
r130 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_4%A_111_47# 1 2 3 4 15 17 18 19 27
r32 25 27 25.7429 $w=3.83e-07 $l=8.6e-07 $layer=LI1_cond $X=2.415 $Y=0.447
+ $X2=3.275 $Y2=0.447
r33 23 30 2.60241 $w=3.85e-07 $l=9.5e-08 $layer=LI1_cond $X=1.65 $Y=0.447
+ $X2=1.555 $Y2=0.447
r34 23 25 22.8992 $w=3.83e-07 $l=7.65e-07 $layer=LI1_cond $X=1.65 $Y=0.447
+ $X2=2.415 $Y2=0.447
r35 20 22 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=1.555 $Y=1.035
+ $X2=1.555 $Y2=0.93
r36 19 30 5.287 $w=1.9e-07 $l=1.93e-07 $layer=LI1_cond $X=1.555 $Y=0.64
+ $X2=1.555 $Y2=0.447
r37 19 22 16.9282 $w=1.88e-07 $l=2.9e-07 $layer=LI1_cond $X=1.555 $Y=0.64
+ $X2=1.555 $Y2=0.93
r38 17 20 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.46 $Y=1.12
+ $X2=1.555 $Y2=1.035
r39 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.46 $Y=1.12
+ $X2=0.79 $Y2=1.12
r40 13 18 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.675 $Y=1.035
+ $X2=0.79 $Y2=1.12
r41 13 15 30.8153 $w=2.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.675 $Y=1.035
+ $X2=0.675 $Y2=0.42
r42 4 27 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=3.135
+ $Y=0.235 $X2=3.275 $Y2=0.475
r43 3 25 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.235 $X2=2.415 $Y2=0.475
r44 2 30 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.235 $X2=1.555 $Y2=0.42
r45 2 22 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.235 $X2=1.555 $Y2=0.93
r46 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.235 $X2=0.695 $Y2=0.42
.ends

