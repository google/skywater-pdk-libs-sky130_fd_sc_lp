* File: sky130_fd_sc_lp__a2111oi_4.pex.spice
* Created: Fri Aug 28 09:46:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111OI_4%D1 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 31 45
r87 43 45 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.675 $Y=1.35
+ $X2=1.765 $Y2=1.35
r88 41 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.335 $Y=1.35
+ $X2=1.675 $Y2=1.35
r89 40 41 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.905 $Y=1.35
+ $X2=1.335 $Y2=1.35
r90 38 40 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.655 $Y=1.35
+ $X2=0.905 $Y2=1.35
r91 35 38 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.475 $Y=1.35
+ $X2=0.655 $Y2=1.35
r92 31 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.675
+ $Y=1.35 $X2=1.675 $Y2=1.35
r93 30 31 24.3294 $w=2.23e-07 $l=4.75e-07 $layer=LI1_cond $X=1.2 $Y=1.322
+ $X2=1.675 $Y2=1.322
r94 29 30 27.9147 $w=2.23e-07 $l=5.45e-07 $layer=LI1_cond $X=0.655 $Y=1.322
+ $X2=1.2 $Y2=1.322
r95 29 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.655
+ $Y=1.35 $X2=0.655 $Y2=1.35
r96 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.515
+ $X2=1.765 $Y2=1.35
r97 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.765 $Y=1.515
+ $X2=1.765 $Y2=2.465
r98 22 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=1.35
r99 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=0.655
r100 18 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.515
+ $X2=1.335 $Y2=1.35
r101 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.335 $Y=1.515
+ $X2=1.335 $Y2=2.465
r102 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.185
+ $X2=1.335 $Y2=1.35
r103 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.335 $Y=1.185
+ $X2=1.335 $Y2=0.655
r104 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.515
+ $X2=0.905 $Y2=1.35
r105 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.905 $Y=1.515
+ $X2=0.905 $Y2=2.465
r106 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=1.35
r107 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=0.655
r108 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=1.35
r109 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=2.465
r110 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=1.35
r111 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%C1 3 7 11 15 19 23 27 31 33 34 35 36 56
r100 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.575
+ $Y=1.51 $X2=3.575 $Y2=1.51
r101 54 56 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.485 $Y=1.51
+ $X2=3.575 $Y2=1.51
r102 53 57 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=3.235 $Y=1.592
+ $X2=3.575 $Y2=1.592
r103 52 54 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.235 $Y=1.51
+ $X2=3.485 $Y2=1.51
r104 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.235
+ $Y=1.51 $X2=3.235 $Y2=1.51
r105 50 52 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.055 $Y=1.51
+ $X2=3.235 $Y2=1.51
r106 48 50 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.895 $Y=1.51
+ $X2=3.055 $Y2=1.51
r107 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.895
+ $Y=1.51 $X2=2.895 $Y2=1.51
r108 46 48 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.895 $Y2=1.51
r109 44 46 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.555 $Y=1.51
+ $X2=2.625 $Y2=1.51
r110 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.555
+ $Y=1.51 $X2=2.555 $Y2=1.51
r111 41 44 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.555 $Y2=1.51
r112 36 57 0.860032 $w=3.33e-07 $l=2.5e-08 $layer=LI1_cond $X=3.6 $Y=1.592
+ $X2=3.575 $Y2=1.592
r113 35 53 3.95615 $w=3.33e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.592
+ $X2=3.235 $Y2=1.592
r114 35 49 7.74029 $w=3.33e-07 $l=2.25e-07 $layer=LI1_cond $X=3.12 $Y=1.592
+ $X2=2.895 $Y2=1.592
r115 34 49 8.77233 $w=3.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.64 $Y=1.592
+ $X2=2.895 $Y2=1.592
r116 34 45 2.92411 $w=3.33e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.592
+ $X2=2.555 $Y2=1.592
r117 33 45 13.5885 $w=3.33e-07 $l=3.95e-07 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=2.555 $Y2=1.592
r118 29 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.675
+ $X2=3.485 $Y2=1.51
r119 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.485 $Y=1.675
+ $X2=3.485 $Y2=2.465
r120 25 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.345
+ $X2=3.485 $Y2=1.51
r121 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.485 $Y=1.345
+ $X2=3.485 $Y2=0.655
r122 21 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.675
+ $X2=3.055 $Y2=1.51
r123 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.055 $Y=1.675
+ $X2=3.055 $Y2=2.465
r124 17 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.345
+ $X2=3.055 $Y2=1.51
r125 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.055 $Y=1.345
+ $X2=3.055 $Y2=0.655
r126 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.675
+ $X2=2.625 $Y2=1.51
r127 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.625 $Y=1.675
+ $X2=2.625 $Y2=2.465
r128 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=1.51
r129 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=0.655
r130 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.675
+ $X2=2.195 $Y2=1.51
r131 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.195 $Y=1.675
+ $X2=2.195 $Y2=2.465
r132 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=1.51
r133 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%B1 3 7 11 15 19 23 27 31 33 34 35 36 58
r97 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.475
+ $Y=1.51 $X2=5.475 $Y2=1.51
r98 56 58 24.5605 $w=3.14e-07 $l=1.6e-07 $layer=POLY_cond $X=5.315 $Y=1.51
+ $X2=5.475 $Y2=1.51
r99 55 56 3.07006 $w=3.14e-07 $l=2e-08 $layer=POLY_cond $X=5.295 $Y=1.51
+ $X2=5.315 $Y2=1.51
r100 54 59 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=5.135 $Y=1.592
+ $X2=5.475 $Y2=1.592
r101 53 55 24.5605 $w=3.14e-07 $l=1.6e-07 $layer=POLY_cond $X=5.135 $Y=1.51
+ $X2=5.295 $Y2=1.51
r102 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.135
+ $Y=1.51 $X2=5.135 $Y2=1.51
r103 51 53 38.3758 $w=3.14e-07 $l=2.5e-07 $layer=POLY_cond $X=4.885 $Y=1.51
+ $X2=5.135 $Y2=1.51
r104 50 51 3.07006 $w=3.14e-07 $l=2e-08 $layer=POLY_cond $X=4.865 $Y=1.51
+ $X2=4.885 $Y2=1.51
r105 48 50 10.7452 $w=3.14e-07 $l=7e-08 $layer=POLY_cond $X=4.795 $Y=1.51
+ $X2=4.865 $Y2=1.51
r106 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.795
+ $Y=1.51 $X2=4.795 $Y2=1.51
r107 46 48 52.1911 $w=3.14e-07 $l=3.4e-07 $layer=POLY_cond $X=4.455 $Y=1.51
+ $X2=4.795 $Y2=1.51
r108 45 46 3.07006 $w=3.14e-07 $l=2e-08 $layer=POLY_cond $X=4.435 $Y=1.51
+ $X2=4.455 $Y2=1.51
r109 43 45 49.121 $w=3.14e-07 $l=3.2e-07 $layer=POLY_cond $X=4.115 $Y=1.51
+ $X2=4.435 $Y2=1.51
r110 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.51 $X2=4.115 $Y2=1.51
r111 41 43 13.8153 $w=3.14e-07 $l=9e-08 $layer=POLY_cond $X=4.025 $Y=1.51
+ $X2=4.115 $Y2=1.51
r112 36 59 1.54806 $w=3.33e-07 $l=4.5e-08 $layer=LI1_cond $X=5.52 $Y=1.592
+ $X2=5.475 $Y2=1.592
r113 35 54 3.26812 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=5.04 $Y=1.592
+ $X2=5.135 $Y2=1.592
r114 35 49 8.42831 $w=3.33e-07 $l=2.45e-07 $layer=LI1_cond $X=5.04 $Y=1.592
+ $X2=4.795 $Y2=1.592
r115 34 49 8.0843 $w=3.33e-07 $l=2.35e-07 $layer=LI1_cond $X=4.56 $Y=1.592
+ $X2=4.795 $Y2=1.592
r116 34 44 15.3086 $w=3.33e-07 $l=4.45e-07 $layer=LI1_cond $X=4.56 $Y=1.592
+ $X2=4.115 $Y2=1.592
r117 33 44 1.20404 $w=3.33e-07 $l=3.5e-08 $layer=LI1_cond $X=4.08 $Y=1.592
+ $X2=4.115 $Y2=1.592
r118 29 58 38.3758 $w=3.14e-07 $l=3.22102e-07 $layer=POLY_cond $X=5.725 $Y=1.675
+ $X2=5.475 $Y2=1.51
r119 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.725 $Y=1.675
+ $X2=5.725 $Y2=2.465
r120 25 56 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.315 $Y=1.345
+ $X2=5.315 $Y2=1.51
r121 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.315 $Y=1.345
+ $X2=5.315 $Y2=0.655
r122 21 55 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.295 $Y=1.675
+ $X2=5.295 $Y2=1.51
r123 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.295 $Y=1.675
+ $X2=5.295 $Y2=2.465
r124 17 51 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.885 $Y=1.345
+ $X2=4.885 $Y2=1.51
r125 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.885 $Y=1.345
+ $X2=4.885 $Y2=0.655
r126 13 50 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.865 $Y=1.675
+ $X2=4.865 $Y2=1.51
r127 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.865 $Y=1.675
+ $X2=4.865 $Y2=2.465
r128 9 46 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=1.345
+ $X2=4.455 $Y2=1.51
r129 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.455 $Y=1.345
+ $X2=4.455 $Y2=0.655
r130 5 45 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.435 $Y=1.675
+ $X2=4.435 $Y2=1.51
r131 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.435 $Y=1.675
+ $X2=4.435 $Y2=2.465
r132 1 41 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.345
+ $X2=4.025 $Y2=1.51
r133 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.025 $Y=1.345
+ $X2=4.025 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%A1 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 50 51
r90 49 51 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=7.535 $Y=1.35
+ $X2=7.655 $Y2=1.35
r91 49 50 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=7.535
+ $Y=1.35 $X2=7.535 $Y2=1.35
r92 47 49 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.465 $Y=1.35
+ $X2=7.535 $Y2=1.35
r93 46 47 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=7.225 $Y=1.35
+ $X2=7.465 $Y2=1.35
r94 45 46 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.015 $Y=1.35
+ $X2=7.225 $Y2=1.35
r95 44 45 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=6.795 $Y=1.35
+ $X2=7.015 $Y2=1.35
r96 43 44 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=6.585 $Y=1.35
+ $X2=6.795 $Y2=1.35
r97 42 43 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=6.365 $Y=1.35
+ $X2=6.585 $Y2=1.35
r98 40 42 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=6.175 $Y=1.35
+ $X2=6.365 $Y2=1.35
r99 40 41 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.175
+ $Y=1.35 $X2=6.175 $Y2=1.35
r100 37 40 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=6.155 $Y=1.35
+ $X2=6.175 $Y2=1.35
r101 32 50 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=7.44 $Y=1.322
+ $X2=7.535 $Y2=1.322
r102 31 32 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.322
+ $X2=7.44 $Y2=1.322
r103 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.322
+ $X2=6.96 $Y2=1.322
r104 30 41 15.622 $w=2.23e-07 $l=3.05e-07 $layer=LI1_cond $X=6.48 $Y=1.322
+ $X2=6.175 $Y2=1.322
r105 29 41 8.96345 $w=2.23e-07 $l=1.75e-07 $layer=LI1_cond $X=6 $Y=1.322
+ $X2=6.175 $Y2=1.322
r106 26 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.185
+ $X2=7.655 $Y2=1.35
r107 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.655 $Y=1.185
+ $X2=7.655 $Y2=0.655
r108 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.465 $Y=1.515
+ $X2=7.465 $Y2=1.35
r109 22 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.465 $Y=1.515
+ $X2=7.465 $Y2=2.465
r110 19 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.225 $Y=1.185
+ $X2=7.225 $Y2=1.35
r111 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.225 $Y=1.185
+ $X2=7.225 $Y2=0.655
r112 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.015 $Y=1.515
+ $X2=7.015 $Y2=1.35
r113 15 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.015 $Y=1.515
+ $X2=7.015 $Y2=2.465
r114 12 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.185
+ $X2=6.795 $Y2=1.35
r115 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.795 $Y=1.185
+ $X2=6.795 $Y2=0.655
r116 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.585 $Y=1.515
+ $X2=6.585 $Y2=1.35
r117 8 10 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.585 $Y=1.515
+ $X2=6.585 $Y2=2.465
r118 5 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.185
+ $X2=6.365 $Y2=1.35
r119 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.365 $Y=1.185
+ $X2=6.365 $Y2=0.655
r120 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.155 $Y=1.515
+ $X2=6.155 $Y2=1.35
r121 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.155 $Y=1.515
+ $X2=6.155 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%A2 3 7 11 15 19 23 27 31 38 39 41 43 63
r82 57 58 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.395 $Y=1.46
+ $X2=9.47 $Y2=1.46
r83 56 57 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=9.04 $Y=1.46
+ $X2=9.395 $Y2=1.46
r84 55 56 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.965 $Y=1.46
+ $X2=9.04 $Y2=1.46
r85 52 63 4.69757 $w=3.83e-07 $l=3.5e-08 $layer=LI1_cond $X=8.45 $Y=1.567
+ $X2=8.485 $Y2=1.567
r86 51 53 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=8.45 $Y=1.46
+ $X2=8.61 $Y2=1.46
r87 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.45
+ $Y=1.46 $X2=8.45 $Y2=1.46
r88 49 51 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=8.445 $Y=1.46
+ $X2=8.45 $Y2=1.46
r89 48 49 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=8.18 $Y=1.46
+ $X2=8.445 $Y2=1.46
r90 46 48 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.015 $Y=1.46
+ $X2=8.18 $Y2=1.46
r91 43 58 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.545 $Y=1.46
+ $X2=9.47 $Y2=1.46
r92 41 52 1.49668 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=8.4 $Y=1.567 $X2=8.45
+ $Y2=1.567
r93 39 43 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=9.81 $Y=1.46
+ $X2=9.545 $Y2=1.46
r94 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.81
+ $Y=1.46 $X2=9.81 $Y2=1.46
r95 36 55 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=8.79 $Y=1.46
+ $X2=8.965 $Y2=1.46
r96 36 53 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=8.79 $Y=1.46 $X2=8.61
+ $Y2=1.46
r97 35 38 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.79 $Y=1.46
+ $X2=9.81 $Y2=1.46
r98 35 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.79 $Y=1.46
+ $X2=8.485 $Y2=1.46
r99 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.79
+ $Y=1.46 $X2=8.79 $Y2=1.46
r100 29 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.47 $Y=1.295
+ $X2=9.47 $Y2=1.46
r101 29 31 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=9.47 $Y=1.295
+ $X2=9.47 $Y2=0.655
r102 25 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.395 $Y=1.625
+ $X2=9.395 $Y2=1.46
r103 25 27 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=9.395 $Y=1.625
+ $X2=9.395 $Y2=2.465
r104 21 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.04 $Y=1.295
+ $X2=9.04 $Y2=1.46
r105 21 23 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=9.04 $Y=1.295
+ $X2=9.04 $Y2=0.655
r106 17 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.965 $Y=1.625
+ $X2=8.965 $Y2=1.46
r107 17 19 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.965 $Y=1.625
+ $X2=8.965 $Y2=2.465
r108 13 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.61 $Y=1.295
+ $X2=8.61 $Y2=1.46
r109 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=8.61 $Y=1.295
+ $X2=8.61 $Y2=0.655
r110 9 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.625
+ $X2=8.445 $Y2=1.46
r111 9 11 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.445 $Y=1.625
+ $X2=8.445 $Y2=2.465
r112 5 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.18 $Y=1.295
+ $X2=8.18 $Y2=1.46
r113 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=8.18 $Y=1.295 $X2=8.18
+ $Y2=0.655
r114 1 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.015 $Y=1.625
+ $X2=8.015 $Y2=1.46
r115 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.015 $Y=1.625
+ $X2=8.015 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%A_27_367# 1 2 3 4 5 16 18 20 24 28 32 36
+ 40 42 46 50 51 52
r80 44 46 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.7 $Y=2.905 $X2=3.7
+ $Y2=2.385
r81 43 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=2.99
+ $X2=2.84 $Y2=2.99
r82 42 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.535 $Y=2.99
+ $X2=3.7 $Y2=2.905
r83 42 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.535 $Y=2.99
+ $X2=3.005 $Y2=2.99
r84 38 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=2.905
+ $X2=2.84 $Y2=2.99
r85 38 40 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=2.84 $Y=2.905
+ $X2=2.84 $Y2=2.385
r86 37 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=2.99
+ $X2=1.98 $Y2=2.99
r87 36 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=2.99
+ $X2=2.84 $Y2=2.99
r88 36 37 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.675 $Y=2.99
+ $X2=2.145 $Y2=2.99
r89 32 35 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=1.98 $Y=2.015
+ $X2=1.98 $Y2=2.9
r90 30 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.905
+ $X2=1.98 $Y2=2.99
r91 30 35 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.98 $Y=2.905
+ $X2=1.98 $Y2=2.9
r92 29 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=2.99
+ $X2=1.12 $Y2=2.99
r93 28 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=2.99
+ $X2=1.98 $Y2=2.99
r94 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.815 $Y=2.99
+ $X2=1.285 $Y2=2.99
r95 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.12 $Y=2.13
+ $X2=1.12 $Y2=2.9
r96 22 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.905
+ $X2=1.12 $Y2=2.99
r97 22 27 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.12 $Y=2.905
+ $X2=1.12 $Y2=2.9
r98 21 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=2.99
+ $X2=0.26 $Y2=2.99
r99 20 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=2.99
+ $X2=1.12 $Y2=2.99
r100 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.955 $Y=2.99
+ $X2=0.425 $Y2=2.99
r101 16 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.905
+ $X2=0.26 $Y2=2.99
r102 16 18 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=0.26 $Y=2.905
+ $X2=0.26 $Y2=2.13
r103 5 46 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.385
r104 4 40 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.385
r105 3 35 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.9
r106 3 32 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.015
r107 2 27 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.9
r108 2 24 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.13
r109 1 49 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r110 1 18 400 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%Y 1 2 3 4 5 6 7 8 9 10 32 33 34 35 36 39
+ 43 45 47 51 55 57 61 63 67 69 73 75 77 81 83 85 86 87 88 92 93 94 96 100 101
+ 107 113 115
c153 73 0 6.54577e-20 $X=4.24 $Y=0.42
c154 67 0 6.86963e-20 $X=3.27 $Y=0.42
r155 115 116 10.75 $w=2.44e-07 $l=2.15e-07 $layer=LI1_cond $X=5.07 $Y=0.955
+ $X2=5.07 $Y2=1.17
r156 105 113 2.684 $w=2.5e-07 $l=5.5e-08 $layer=LI1_cond $X=5.07 $Y=0.87
+ $X2=5.07 $Y2=0.925
r157 101 115 0.75 $w=2.44e-07 $l=1.5e-08 $layer=LI1_cond $X=5.07 $Y=0.94
+ $X2=5.07 $Y2=0.955
r158 101 113 0.75 $w=2.44e-07 $l=1.5e-08 $layer=LI1_cond $X=5.07 $Y=0.94
+ $X2=5.07 $Y2=0.925
r159 101 105 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=5.07 $Y=0.855
+ $X2=5.07 $Y2=0.87
r160 100 101 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=5.07 $Y=0.555
+ $X2=5.07 $Y2=0.855
r161 100 107 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=5.07 $Y=0.555
+ $X2=5.07 $Y2=0.42
r162 88 90 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=2.405 $Y=0.955
+ $X2=2.405 $Y2=1.17
r163 88 89 4.75232 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=0.955
+ $X2=2.405 $Y2=0.87
r164 84 94 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=6.705 $Y=0.955
+ $X2=6.582 $Y2=0.955
r165 83 96 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=7.457 $Y=0.955
+ $X2=7.457 $Y2=0.76
r166 83 84 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.31 $Y=0.955
+ $X2=6.705 $Y2=0.955
r167 79 94 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=6.582 $Y=0.87
+ $X2=6.582 $Y2=0.955
r168 79 81 5.17423 $w=2.43e-07 $l=1.1e-07 $layer=LI1_cond $X=6.582 $Y=0.87
+ $X2=6.582 $Y2=0.76
r169 78 115 2.85362 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.195 $Y=0.955
+ $X2=5.07 $Y2=0.955
r170 77 94 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=6.46 $Y=0.955
+ $X2=6.582 $Y2=0.955
r171 77 78 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=6.46 $Y=0.955
+ $X2=5.195 $Y2=0.955
r172 76 93 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.335 $Y=1.17
+ $X2=4.215 $Y2=1.17
r173 75 116 2.85362 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.945 $Y=1.17
+ $X2=5.07 $Y2=1.17
r174 75 76 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.945 $Y=1.17
+ $X2=4.335 $Y2=1.17
r175 71 93 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=1.085
+ $X2=4.215 $Y2=1.17
r176 71 73 31.9323 $w=2.38e-07 $l=6.65e-07 $layer=LI1_cond $X=4.215 $Y=1.085
+ $X2=4.215 $Y2=0.42
r177 70 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.425 $Y=1.17
+ $X2=3.3 $Y2=1.17
r178 69 93 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.095 $Y=1.17
+ $X2=4.215 $Y2=1.17
r179 69 70 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.095 $Y=1.17
+ $X2=3.425 $Y2=1.17
r180 65 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=1.085
+ $X2=3.3 $Y2=1.17
r181 65 67 30.655 $w=2.48e-07 $l=6.65e-07 $layer=LI1_cond $X=3.3 $Y=1.085
+ $X2=3.3 $Y2=0.42
r182 64 90 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.505 $Y=1.17
+ $X2=2.405 $Y2=1.17
r183 63 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.175 $Y=1.17
+ $X2=3.3 $Y2=1.17
r184 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.175 $Y=1.17
+ $X2=2.505 $Y2=1.17
r185 61 89 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=2.41 $Y=0.42
+ $X2=2.41 $Y2=0.87
r186 58 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.645 $Y=0.955
+ $X2=1.55 $Y2=0.955
r187 57 88 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.305 $Y=0.955
+ $X2=2.405 $Y2=0.955
r188 57 58 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.305 $Y=0.955
+ $X2=1.645 $Y2=0.955
r189 53 55 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=1.55 $Y=1.875
+ $X2=1.55 $Y2=1.98
r190 49 87 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.87
+ $X2=1.55 $Y2=0.955
r191 49 51 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=1.55 $Y=0.87
+ $X2=1.55 $Y2=0.42
r192 48 86 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.785 $Y=1.79
+ $X2=0.69 $Y2=1.79
r193 47 53 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.455 $Y=1.79
+ $X2=1.55 $Y2=1.875
r194 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.455 $Y=1.79
+ $X2=0.785 $Y2=1.79
r195 46 85 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.785 $Y=0.955
+ $X2=0.69 $Y2=0.955
r196 45 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.455 $Y=0.955
+ $X2=1.55 $Y2=0.955
r197 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.455 $Y=0.955
+ $X2=0.785 $Y2=0.955
r198 41 86 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.875
+ $X2=0.69 $Y2=1.79
r199 41 43 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=0.69 $Y=1.875
+ $X2=0.69 $Y2=1.98
r200 37 85 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.87
+ $X2=0.69 $Y2=0.955
r201 37 39 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=0.87
+ $X2=0.69 $Y2=0.42
r202 35 86 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.595 $Y=1.79
+ $X2=0.69 $Y2=1.79
r203 35 36 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.595 $Y=1.79
+ $X2=0.32 $Y2=1.79
r204 33 85 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.595 $Y=0.955
+ $X2=0.69 $Y2=0.955
r205 33 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.595 $Y=0.955
+ $X2=0.32 $Y2=0.955
r206 32 36 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.23 $Y=1.705
+ $X2=0.32 $Y2=1.79
r207 31 34 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.23 $Y=1.04
+ $X2=0.32 $Y2=0.955
r208 31 32 40.9747 $w=1.78e-07 $l=6.65e-07 $layer=LI1_cond $X=0.23 $Y=1.04
+ $X2=0.23 $Y2=1.705
r209 10 55 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=1.98
r210 9 43 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=1.98
r211 8 96 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=7.3
+ $Y=0.235 $X2=7.44 $Y2=0.76
r212 7 81 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=6.44
+ $Y=0.235 $X2=6.58 $Y2=0.76
r213 6 107 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.96
+ $Y=0.235 $X2=5.1 $Y2=0.42
r214 5 73 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.1
+ $Y=0.235 $X2=4.24 $Y2=0.42
r215 4 67 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.42
r216 3 61 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.42
r217 2 51 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.42
r218 1 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%A_454_367# 1 2 3 4 15 19 23 28 30 32 34
r47 24 32 6.30264 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=4.785 $Y=2.025
+ $X2=4.67 $Y2=2.025
r48 23 34 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.345 $Y=2.025
+ $X2=5.51 $Y2=2.025
r49 23 24 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=5.345 $Y=2.025
+ $X2=4.785 $Y2=2.025
r50 20 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.365 $Y=2.015
+ $X2=3.27 $Y2=2.015
r51 19 32 6.30264 $w=1.8e-07 $l=1.19896e-07 $layer=LI1_cond $X=4.555 $Y=2.015
+ $X2=4.67 $Y2=2.025
r52 19 20 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=4.555 $Y=2.015
+ $X2=3.365 $Y2=2.015
r53 16 28 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.505 $Y=2.015
+ $X2=2.41 $Y2=2.015
r54 15 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.175 $Y=2.015
+ $X2=3.27 $Y2=2.015
r55 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.175 $Y=2.015
+ $X2=2.505 $Y2=2.015
r56 4 34 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=5.37
+ $Y=1.835 $X2=5.51 $Y2=2.095
r57 3 32 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=4.51
+ $Y=1.835 $X2=4.65 $Y2=2.095
r58 2 30 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.095
r59 1 28 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%A_819_367# 1 2 3 4 5 6 7 24 26 27 30 32 35
+ 37 38 39 42 46 49 52 54 56 58 60 64 68 71
r99 76 77 1.86463 $w=2.29e-07 $l=3.5e-08 $layer=LI1_cond $X=8.705 $Y=1.98
+ $X2=8.705 $Y2=2.015
r100 74 76 9.58952 $w=2.29e-07 $l=1.8e-07 $layer=LI1_cond $X=8.705 $Y=1.8
+ $X2=8.705 $Y2=1.98
r101 64 66 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=9.645 $Y=1.98
+ $X2=9.645 $Y2=2.91
r102 62 64 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=9.645 $Y=1.885
+ $X2=9.645 $Y2=1.98
r103 61 74 2.48377 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.845 $Y=1.8
+ $X2=8.705 $Y2=1.8
r104 60 62 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.515 $Y=1.8
+ $X2=9.645 $Y2=1.885
r105 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.515 $Y=1.8
+ $X2=8.845 $Y2=1.8
r106 56 77 4.14435 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.705 $Y=2.1
+ $X2=8.705 $Y2=2.015
r107 56 58 14.6113 $w=2.78e-07 $l=3.55e-07 $layer=LI1_cond $X=8.705 $Y=2.1
+ $X2=8.705 $Y2=2.455
r108 55 73 3.05049 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.895 $Y=2.015
+ $X2=7.73 $Y2=2.015
r109 54 77 2.48377 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.565 $Y=2.015
+ $X2=8.705 $Y2=2.015
r110 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.565 $Y=2.015
+ $X2=7.895 $Y2=2.015
r111 50 73 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.73 $Y=2.1 $X2=7.73
+ $Y2=2.015
r112 50 52 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=7.73 $Y=2.1
+ $X2=7.73 $Y2=2.475
r113 49 73 3.46198 $w=2.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=7.67 $Y=1.93
+ $X2=7.73 $Y2=2.015
r114 48 49 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=7.67 $Y=1.775
+ $X2=7.67 $Y2=1.93
r115 47 71 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.895 $Y=1.69
+ $X2=6.8 $Y2=1.69
r116 46 48 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.565 $Y=1.69
+ $X2=7.67 $Y2=1.775
r117 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.565 $Y=1.69
+ $X2=6.895 $Y2=1.69
r118 42 44 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.8 $Y=1.98 $X2=6.8
+ $Y2=2.91
r119 40 71 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.8 $Y=1.775
+ $X2=6.8 $Y2=1.69
r120 40 42 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=6.8 $Y=1.775
+ $X2=6.8 $Y2=1.98
r121 38 71 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.705 $Y=1.69
+ $X2=6.8 $Y2=1.69
r122 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.705 $Y=1.69
+ $X2=6.035 $Y2=1.69
r123 35 70 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=2.905
+ $X2=5.94 $Y2=2.99
r124 35 37 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=5.94 $Y=2.905
+ $X2=5.94 $Y2=1.98
r125 34 39 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.94 $Y=1.775
+ $X2=6.035 $Y2=1.69
r126 34 37 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=5.94 $Y=1.775
+ $X2=5.94 $Y2=1.98
r127 33 68 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=5.175 $Y=2.99
+ $X2=5.065 $Y2=2.99
r128 32 70 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.845 $Y=2.99
+ $X2=5.94 $Y2=2.99
r129 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.845 $Y=2.99
+ $X2=5.175 $Y2=2.99
r130 28 68 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=2.905
+ $X2=5.065 $Y2=2.99
r131 28 30 22.7869 $w=2.18e-07 $l=4.35e-07 $layer=LI1_cond $X=5.065 $Y=2.905
+ $X2=5.065 $Y2=2.47
r132 26 68 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.955 $Y=2.99
+ $X2=5.065 $Y2=2.99
r133 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.955 $Y=2.99
+ $X2=4.385 $Y2=2.99
r134 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.22 $Y=2.905
+ $X2=4.385 $Y2=2.99
r135 22 24 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=4.22 $Y=2.905
+ $X2=4.22 $Y2=2.385
r136 7 66 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.47
+ $Y=1.835 $X2=9.61 $Y2=2.91
r137 7 64 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.47
+ $Y=1.835 $X2=9.61 $Y2=1.98
r138 6 76 600 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_PDIFF $count=1 $X=8.52
+ $Y=1.835 $X2=8.75 $Y2=1.98
r139 6 58 300 $w=1.7e-07 $l=7.0647e-07 $layer=licon1_PDIFF $count=2 $X=8.52
+ $Y=1.835 $X2=8.705 $Y2=2.455
r140 5 73 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=1.835 $X2=7.68 $Y2=1.98
r141 5 52 300 $w=1.7e-07 $l=7.28835e-07 $layer=licon1_PDIFF $count=2 $X=7.54
+ $Y=1.835 $X2=7.73 $Y2=2.475
r142 4 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.66
+ $Y=1.835 $X2=6.8 $Y2=2.91
r143 4 42 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.66
+ $Y=1.835 $X2=6.8 $Y2=1.98
r144 3 70 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.8
+ $Y=1.835 $X2=5.94 $Y2=2.91
r145 3 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.8
+ $Y=1.835 $X2=5.94 $Y2=1.98
r146 2 30 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=4.94
+ $Y=1.835 $X2=5.08 $Y2=2.47
r147 1 24 300 $w=1.7e-07 $l=6.09303e-07 $layer=licon1_PDIFF $count=2 $X=4.095
+ $Y=1.835 $X2=4.22 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%VPWR 1 2 3 4 15 21 27 31 36 37 39 40 42 43
+ 45 46 47 66 67
r128 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r129 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r130 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r131 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r132 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r133 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r135 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r136 54 55 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r137 50 54 375.786 $w=1.68e-07 $l=5.76e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=6
+ $Y2=3.33
r138 50 51 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 47 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r140 47 51 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=0.24 $Y2=3.33
r141 45 63 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=9.015 $Y=3.33
+ $X2=8.88 $Y2=3.33
r142 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.015 $Y=3.33
+ $X2=9.18 $Y2=3.33
r143 44 66 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.345 $Y=3.33
+ $X2=9.84 $Y2=3.33
r144 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.345 $Y=3.33
+ $X2=9.18 $Y2=3.33
r145 42 60 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.065 $Y=3.33
+ $X2=7.92 $Y2=3.33
r146 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.065 $Y=3.33
+ $X2=8.23 $Y2=3.33
r147 41 63 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.395 $Y=3.33
+ $X2=8.88 $Y2=3.33
r148 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.395 $Y=3.33
+ $X2=8.23 $Y2=3.33
r149 39 57 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.065 $Y=3.33
+ $X2=6.96 $Y2=3.33
r150 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.065 $Y=3.33
+ $X2=7.23 $Y2=3.33
r151 38 60 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=7.395 $Y=3.33
+ $X2=7.92 $Y2=3.33
r152 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.395 $Y=3.33
+ $X2=7.23 $Y2=3.33
r153 36 54 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.205 $Y=3.33
+ $X2=6 $Y2=3.33
r154 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.205 $Y=3.33
+ $X2=6.37 $Y2=3.33
r155 35 57 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.535 $Y=3.33
+ $X2=6.96 $Y2=3.33
r156 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=3.33
+ $X2=6.37 $Y2=3.33
r157 31 34 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=9.18 $Y=2.14
+ $X2=9.18 $Y2=2.95
r158 29 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.18 $Y=3.245
+ $X2=9.18 $Y2=3.33
r159 29 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.18 $Y=3.245
+ $X2=9.18 $Y2=2.95
r160 25 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.23 $Y=3.245
+ $X2=8.23 $Y2=3.33
r161 25 27 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=8.23 $Y=3.245
+ $X2=8.23 $Y2=2.38
r162 21 24 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=7.23 $Y=2.03
+ $X2=7.23 $Y2=2.95
r163 19 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.23 $Y=3.245
+ $X2=7.23 $Y2=3.33
r164 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.23 $Y=3.245
+ $X2=7.23 $Y2=2.95
r165 15 18 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=6.37 $Y=2.03
+ $X2=6.37 $Y2=2.95
r166 13 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=3.245
+ $X2=6.37 $Y2=3.33
r167 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.37 $Y=3.245
+ $X2=6.37 $Y2=2.95
r168 4 34 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.04
+ $Y=1.835 $X2=9.18 $Y2=2.95
r169 4 31 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=9.04
+ $Y=1.835 $X2=9.18 $Y2=2.14
r170 3 27 300 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=2 $X=8.09
+ $Y=1.835 $X2=8.23 $Y2=2.38
r171 2 24 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.09
+ $Y=1.835 $X2=7.23 $Y2=2.95
r172 2 21 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=7.09
+ $Y=1.835 $X2=7.23 $Y2=2.03
r173 1 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.23
+ $Y=1.835 $X2=6.37 $Y2=2.95
r174 1 15 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=6.23
+ $Y=1.835 $X2=6.37 $Y2=2.03
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 44
+ 48 50 54 58 62 66 69 70 71 72 74 75 76 78 90 95 108 109 115 118 121 124 127
r155 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r156 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r157 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r158 119 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.56 $Y2=0
r159 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r160 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r161 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r162 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r163 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.84 $Y2=0
r164 106 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=8.4 $Y2=0
r165 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r166 103 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.56 $Y=0
+ $X2=8.395 $Y2=0
r167 103 105 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.56 $Y=0 $X2=8.88
+ $Y2=0
r168 102 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r169 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r170 99 102 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=7.92
+ $Y2=0
r171 99 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r172 98 101 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=0 $X2=7.92
+ $Y2=0
r173 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r174 96 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.695 $Y=0
+ $X2=5.53 $Y2=0
r175 96 98 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.695 $Y=0 $X2=6
+ $Y2=0
r176 95 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.23 $Y=0
+ $X2=8.395 $Y2=0
r177 95 101 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.23 $Y=0 $X2=7.92
+ $Y2=0
r178 91 121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.775 $Y=0
+ $X2=4.64 $Y2=0
r179 91 93 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.775 $Y=0
+ $X2=5.04 $Y2=0
r180 90 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=0
+ $X2=5.53 $Y2=0
r181 90 93 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.365 $Y=0
+ $X2=5.04 $Y2=0
r182 89 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r183 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r184 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r185 86 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r186 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r187 83 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.12 $Y2=0
r188 83 85 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.68 $Y2=0
r189 82 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r190 82 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r191 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r192 79 112 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r193 79 81 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r194 78 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0
+ $X2=1.12 $Y2=0
r195 78 81 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=0
+ $X2=0.72 $Y2=0
r196 76 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r197 76 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r198 76 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r199 74 105 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.09 $Y=0 $X2=8.88
+ $Y2=0
r200 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.09 $Y=0 $X2=9.255
+ $Y2=0
r201 73 108 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.42 $Y=0 $X2=9.84
+ $Y2=0
r202 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.42 $Y=0 $X2=9.255
+ $Y2=0
r203 71 88 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.64
+ $Y2=0
r204 71 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.84
+ $Y2=0
r205 69 85 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=0
+ $X2=1.68 $Y2=0
r206 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.98
+ $Y2=0
r207 68 88 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.145 $Y=0
+ $X2=2.64 $Y2=0
r208 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=1.98
+ $Y2=0
r209 64 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.255 $Y=0.085
+ $X2=9.255 $Y2=0
r210 64 66 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.255 $Y=0.085
+ $X2=9.255 $Y2=0.38
r211 60 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.395 $Y=0.085
+ $X2=8.395 $Y2=0
r212 60 62 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.395 $Y=0.085
+ $X2=8.395 $Y2=0.38
r213 56 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=0.085
+ $X2=5.53 $Y2=0
r214 56 58 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.53 $Y=0.085
+ $X2=5.53 $Y2=0.565
r215 52 121 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0
r216 52 54 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0.38
r217 51 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=0
+ $X2=3.76 $Y2=0
r218 50 121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.505 $Y=0
+ $X2=4.64 $Y2=0
r219 50 51 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.505 $Y=0
+ $X2=3.925 $Y2=0
r220 46 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.76 $Y2=0
r221 46 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.76 $Y2=0.38
r222 45 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=0 $X2=2.84
+ $Y2=0
r223 44 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=3.76 $Y2=0
r224 44 45 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.595 $Y=0 $X2=3.005
+ $Y2=0
r225 40 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r226 40 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.38
r227 36 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r228 36 38 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.575
r229 32 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r230 32 34 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.575
r231 28 112 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r232 28 30 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.575
r233 9 66 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.115
+ $Y=0.235 $X2=9.255 $Y2=0.38
r234 8 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.255
+ $Y=0.235 $X2=8.395 $Y2=0.38
r235 7 58 182 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_NDIFF $count=1 $X=5.39
+ $Y=0.235 $X2=5.53 $Y2=0.565
r236 6 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.53
+ $Y=0.235 $X2=4.67 $Y2=0.38
r237 5 48 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.235 $X2=3.76 $Y2=0.38
r238 4 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.38
r239 3 38 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.575
r240 2 34 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.575
r241 1 30 182 $w=1.7e-07 $l=3.97618e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_4%A_1201_47# 1 2 3 4 5 16 20 22 24 25 26 27
+ 30 32 36 38 43 46
r63 38 41 6.91466 $w=3.23e-07 $l=1.95e-07 $layer=LI1_cond $X=6.127 $Y=0.34
+ $X2=6.127 $Y2=0.535
r64 34 36 27.2597 $w=2.58e-07 $l=6.15e-07 $layer=LI1_cond $X=9.72 $Y=1.035
+ $X2=9.72 $Y2=0.42
r65 33 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.92 $Y=1.12
+ $X2=8.825 $Y2=1.12
r66 32 34 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.59 $Y=1.12
+ $X2=9.72 $Y2=1.035
r67 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.59 $Y=1.12
+ $X2=8.92 $Y2=1.12
r68 28 46 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.825 $Y=1.035
+ $X2=8.825 $Y2=1.12
r69 28 30 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=8.825 $Y=1.035
+ $X2=8.825 $Y2=0.42
r70 26 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.73 $Y=1.12
+ $X2=8.825 $Y2=1.12
r71 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.73 $Y=1.12
+ $X2=8.06 $Y2=1.12
r72 25 27 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.965 $Y=1.035
+ $X2=8.06 $Y2=1.12
r73 24 45 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.965 $Y=0.425
+ $X2=7.965 $Y2=0.34
r74 24 25 35.6077 $w=1.88e-07 $l=6.1e-07 $layer=LI1_cond $X=7.965 $Y=0.425
+ $X2=7.965 $Y2=1.035
r75 23 43 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=7.14 $Y=0.34
+ $X2=7.007 $Y2=0.34
r76 22 45 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.87 $Y=0.34
+ $X2=7.965 $Y2=0.34
r77 22 23 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.87 $Y=0.34
+ $X2=7.14 $Y2=0.34
r78 18 43 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.007 $Y=0.425
+ $X2=7.007 $Y2=0.34
r79 18 20 4.78373 $w=2.63e-07 $l=1.1e-07 $layer=LI1_cond $X=7.007 $Y=0.425
+ $X2=7.007 $Y2=0.535
r80 17 38 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=6.29 $Y=0.34
+ $X2=6.127 $Y2=0.34
r81 16 43 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=6.875 $Y=0.34
+ $X2=7.007 $Y2=0.34
r82 16 17 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=6.875 $Y=0.34
+ $X2=6.29 $Y2=0.34
r83 5 36 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.545
+ $Y=0.235 $X2=9.685 $Y2=0.42
r84 4 30 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.685
+ $Y=0.235 $X2=8.825 $Y2=0.42
r85 3 45 91 $w=1.7e-07 $l=3.0895e-07 $layer=licon1_NDIFF $count=2 $X=7.73
+ $Y=0.235 $X2=7.96 $Y2=0.42
r86 2 20 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=6.87
+ $Y=0.235 $X2=7.01 $Y2=0.535
r87 1 41 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=6.005
+ $Y=0.235 $X2=6.13 $Y2=0.535
.ends

