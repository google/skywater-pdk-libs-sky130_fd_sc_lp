* File: sky130_fd_sc_lp__inputiso1p_lp.pex.spice
* Created: Fri Aug 28 10:37:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INPUTISO1P_LP%A 1 3 4 6 8 10 11 12
r35 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.06
+ $Y=1.48 $X2=1.06 $Y2=1.48
r36 12 17 4.10364 $w=5.5e-07 $l=1.85e-07 $layer=LI1_cond $X=0.89 $Y=1.665
+ $X2=0.89 $Y2=1.48
r37 11 17 4.10364 $w=5.5e-07 $l=2.56271e-07 $layer=LI1_cond $X=0.72 $Y=1.295
+ $X2=0.89 $Y2=1.48
r38 8 16 88.9511 $w=2.9e-07 $l=6.40937e-07 $layer=POLY_cond $X=1.17 $Y=0.96
+ $X2=0.9 $Y2=1.48
r39 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.17 $Y=0.96 $X2=1.17
+ $Y2=0.675
r40 4 16 44.0725 $w=5.81e-07 $l=3.22102e-07 $layer=POLY_cond $X=1.15 $Y=1.645
+ $X2=0.9 $Y2=1.48
r41 4 6 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.15 $Y=1.645
+ $X2=1.15 $Y2=2.655
r42 1 16 88.9511 $w=2.9e-07 $l=5.63205e-07 $layer=POLY_cond $X=0.81 $Y=0.96
+ $X2=0.9 $Y2=1.48
r43 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.81 $Y=0.96 $X2=0.81
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO1P_LP%SLEEP 3 7 11 13 20 21
c40 20 0 7.06387e-20 $X=1.94 $Y=1.48
r41 19 21 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.94 $Y=1.48 $X2=1.96
+ $Y2=1.48
r42 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.94
+ $Y=1.48 $X2=1.94 $Y2=1.48
r43 17 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.6 $Y=1.48 $X2=1.94
+ $Y2=1.48
r44 15 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.51 $Y=1.48 $X2=1.6
+ $Y2=1.48
r45 13 20 3.3026 $w=6.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.77 $Y=1.665
+ $X2=1.77 $Y2=1.48
r46 9 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.315
+ $X2=1.96 $Y2=1.48
r47 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.96 $Y=1.315 $X2=1.96
+ $Y2=0.675
r48 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.6 $Y=1.315 $X2=1.6
+ $Y2=1.48
r49 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.6 $Y=1.315 $X2=1.6
+ $Y2=0.675
r50 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.51 $Y=1.645
+ $X2=1.51 $Y2=1.48
r51 1 3 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.51 $Y=1.645
+ $X2=1.51 $Y2=2.655
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO1P_LP%A_161_489# 1 2 7 9 12 14 16 19 23 25
+ 26 29 31 32 33 34 37
r64 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.515
+ $Y=1.17 $X2=2.515 $Y2=1.17
r65 33 36 2.63384 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.517 $Y=1.18
+ $X2=2.517 $Y2=1.095
r66 33 34 26.661 $w=3.33e-07 $l=7.75e-07 $layer=LI1_cond $X=2.517 $Y=1.18
+ $X2=2.517 $Y2=1.955
r67 31 36 5.17472 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.35 $Y=1.095
+ $X2=2.517 $Y2=1.095
r68 31 32 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.35 $Y=1.095
+ $X2=1.49 $Y2=1.095
r69 27 32 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.385 $Y=1.01
+ $X2=1.49 $Y2=1.095
r70 27 29 15.316 $w=2.08e-07 $l=2.9e-07 $layer=LI1_cond $X=1.385 $Y=1.01
+ $X2=1.385 $Y2=0.72
r71 25 34 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=2.35 $Y=2.04
+ $X2=2.517 $Y2=1.955
r72 25 26 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.35 $Y=2.04
+ $X2=1.1 $Y2=2.04
r73 21 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.935 $Y=2.125
+ $X2=1.1 $Y2=2.04
r74 21 23 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.935 $Y=2.125
+ $X2=0.935 $Y2=2.655
r75 17 37 97.1997 $w=2.55e-07 $l=5.88154e-07 $layer=POLY_cond $X=2.75 $Y=1.675
+ $X2=2.57 $Y2=1.17
r76 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.75 $Y=1.675
+ $X2=2.75 $Y2=2.465
r77 14 37 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=2.75 $Y=1.005
+ $X2=2.57 $Y2=1.17
r78 14 16 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.75 $Y=1.005
+ $X2=2.75 $Y2=0.675
r79 10 37 97.1997 $w=2.55e-07 $l=5.88154e-07 $layer=POLY_cond $X=2.39 $Y=1.675
+ $X2=2.57 $Y2=1.17
r80 10 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.39 $Y=1.675
+ $X2=2.39 $Y2=2.465
r81 7 37 32.933 $w=2.55e-07 $l=1.8e-07 $layer=POLY_cond $X=2.39 $Y=1.17 $X2=2.57
+ $Y2=1.17
r82 7 9 106.04 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.39 $Y=1.17 $X2=2.39
+ $Y2=0.675
r83 2 23 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=0.805
+ $Y=2.445 $X2=0.935 $Y2=2.655
r84 1 29 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.245
+ $Y=0.465 $X2=1.385 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO1P_LP%VPWR 1 6 10 12 22 23 26
r27 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 23 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r30 20 26 14.6804 $w=1.7e-07 $l=4.03e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=1.962 $Y2=3.33
r31 20 22 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 18 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 15 19 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r34 14 18 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 12 26 14.6804 $w=1.7e-07 $l=4.02e-07 $layer=LI1_cond $X=1.56 $Y=3.33
+ $X2=1.962 $Y2=3.33
r37 12 18 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.56 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 10 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 10 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 6 9 4.08598 $w=8.03e-07 $l=2.75e-07 $layer=LI1_cond $X=1.962 $Y=2.38
+ $X2=1.962 $Y2=2.655
r41 4 26 3.14386 $w=8.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.962 $Y=3.245
+ $X2=1.962 $Y2=3.33
r42 4 9 8.76629 $w=8.03e-07 $l=5.9e-07 $layer=LI1_cond $X=1.962 $Y=3.245
+ $X2=1.962 $Y2=2.655
r43 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=2.445 $X2=1.725 $Y2=2.655
r44 1 6 300 $w=1.7e-07 $l=6.21651e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=2.445 $X2=2.175 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO1P_LP%X 1 2 7 8 9 10 11 18 21 24 27 30 35
r10 33 35 7.54576 $w=4.18e-07 $l=2.75e-07 $layer=LI1_cond $X=3.065 $Y=2.125
+ $X2=3.065 $Y2=2.4
r11 18 21 5.48782 $w=4.18e-07 $l=2e-07 $layer=LI1_cond $X=3.065 $Y=0.72
+ $X2=3.065 $Y2=0.92
r12 11 38 13.5824 $w=4.18e-07 $l=4.95e-07 $layer=LI1_cond $X=3.065 $Y=2.405
+ $X2=3.065 $Y2=2.9
r13 11 35 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=2.405
+ $X2=3.065 $Y2=2.4
r14 10 33 2.46952 $w=4.18e-07 $l=9e-08 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=3.065 $Y2=2.125
r15 10 30 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=3.065 $Y2=2.03
r16 9 30 10.0153 $w=4.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.065 $Y=1.665
+ $X2=3.065 $Y2=2.03
r17 9 27 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=1.665
+ $X2=3.065 $Y2=1.66
r18 8 27 10.0153 $w=4.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.065 $Y=1.295
+ $X2=3.065 $Y2=1.66
r19 8 24 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=1.295
+ $X2=3.065 $Y2=1.29
r20 7 24 10.0153 $w=4.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.065 $Y=0.925
+ $X2=3.065 $Y2=1.29
r21 7 21 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=0.925
+ $X2=3.065 $Y2=0.92
r22 2 38 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.835 $X2=2.965 $Y2=2.9
r23 2 33 400 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.835 $X2=2.965 $Y2=2.125
r24 1 18 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.465 $X2=2.965 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO1P_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r35 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r36 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r37 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.175
+ $Y2=0
r40 27 29 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=3.12
+ $Y2=0
r41 23 33 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.61
+ $Y2=0
r42 23 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.76 $Y=0 $X2=1.68
+ $Y2=0
r43 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.175
+ $Y2=0
r44 22 25 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.68
+ $Y2=0
r45 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r46 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 17 33 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.61
+ $Y2=0
r48 17 19 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.24
+ $Y2=0
r49 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r50 15 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r51 15 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0
r53 11 13 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0.675
r54 7 33 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=0.085 $X2=0.61
+ $Y2=0
r55 7 9 22.6647 $w=2.98e-07 $l=5.9e-07 $layer=LI1_cond $X=0.61 $Y=0.085 $X2=0.61
+ $Y2=0.675
r56 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.035
+ $Y=0.465 $X2=2.175 $Y2=0.675
r57 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.47
+ $Y=0.465 $X2=0.595 $Y2=0.675
.ends

