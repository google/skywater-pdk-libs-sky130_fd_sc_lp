* File: sky130_fd_sc_lp__dlrbn_1.pxi.spice
* Created: Fri Aug 28 10:25:32 2020
* 
x_PM_SKY130_FD_SC_LP__DLRBN_1%GATE_N N_GATE_N_c_192_n N_GATE_N_M1009_g
+ N_GATE_N_M1011_g N_GATE_N_c_198_n GATE_N GATE_N GATE_N GATE_N N_GATE_N_c_195_n
+ PM_SKY130_FD_SC_LP__DLRBN_1%GATE_N
x_PM_SKY130_FD_SC_LP__DLRBN_1%A_112_70# N_A_112_70#_M1009_d N_A_112_70#_M1011_d
+ N_A_112_70#_c_223_n N_A_112_70#_c_224_n N_A_112_70#_M1001_g
+ N_A_112_70#_M1005_g N_A_112_70#_c_233_n N_A_112_70#_c_234_n
+ N_A_112_70#_c_235_n N_A_112_70#_c_236_n N_A_112_70#_M1016_g
+ N_A_112_70#_c_237_n N_A_112_70#_M1000_g N_A_112_70#_c_227_n
+ N_A_112_70#_c_239_n N_A_112_70#_c_240_n N_A_112_70#_c_241_n
+ N_A_112_70#_c_242_n N_A_112_70#_c_243_n N_A_112_70#_c_244_n
+ N_A_112_70#_c_245_n N_A_112_70#_c_228_n N_A_112_70#_c_229_n
+ N_A_112_70#_c_247_n N_A_112_70#_c_230_n N_A_112_70#_c_248_n
+ PM_SKY130_FD_SC_LP__DLRBN_1%A_112_70#
x_PM_SKY130_FD_SC_LP__DLRBN_1%D N_D_c_352_n N_D_M1017_g N_D_M1018_g D D
+ N_D_c_355_n PM_SKY130_FD_SC_LP__DLRBN_1%D
x_PM_SKY130_FD_SC_LP__DLRBN_1%A_207_40# N_A_207_40#_M1001_s N_A_207_40#_M1005_s
+ N_A_207_40#_c_389_n N_A_207_40#_M1007_g N_A_207_40#_c_391_n
+ N_A_207_40#_c_392_n N_A_207_40#_M1013_g N_A_207_40#_c_394_n
+ N_A_207_40#_c_395_n N_A_207_40#_c_399_n N_A_207_40#_c_396_n
+ N_A_207_40#_c_397_n PM_SKY130_FD_SC_LP__DLRBN_1%A_207_40#
x_PM_SKY130_FD_SC_LP__DLRBN_1%A_437_144# N_A_437_144#_M1017_d
+ N_A_437_144#_M1018_d N_A_437_144#_c_470_n N_A_437_144#_c_471_n
+ N_A_437_144#_c_472_n N_A_437_144#_M1015_g N_A_437_144#_c_474_n
+ N_A_437_144#_M1019_g N_A_437_144#_c_475_n N_A_437_144#_c_476_n
+ N_A_437_144#_c_483_n N_A_437_144#_c_484_n N_A_437_144#_c_477_n
+ N_A_437_144#_c_478_n N_A_437_144#_c_479_n N_A_437_144#_c_480_n
+ N_A_437_144#_c_481_n PM_SKY130_FD_SC_LP__DLRBN_1%A_437_144#
x_PM_SKY130_FD_SC_LP__DLRBN_1%A_955_271# N_A_955_271#_M1008_s
+ N_A_955_271#_M1012_d N_A_955_271#_M1004_g N_A_955_271#_M1021_g
+ N_A_955_271#_M1020_g N_A_955_271#_c_564_n N_A_955_271#_M1023_g
+ N_A_955_271#_M1014_g N_A_955_271#_c_566_n N_A_955_271#_M1006_g
+ N_A_955_271#_c_567_n N_A_955_271#_c_568_n N_A_955_271#_c_587_n
+ N_A_955_271#_c_569_n N_A_955_271#_c_570_n N_A_955_271#_c_598_p
+ N_A_955_271#_c_588_n N_A_955_271#_c_610_p N_A_955_271#_c_625_p
+ N_A_955_271#_c_659_p N_A_955_271#_c_571_n N_A_955_271#_c_572_n
+ N_A_955_271#_c_573_n N_A_955_271#_c_574_n N_A_955_271#_c_575_n
+ N_A_955_271#_c_576_n N_A_955_271#_c_577_n N_A_955_271#_c_578_n
+ N_A_955_271#_c_579_n N_A_955_271#_c_580_n N_A_955_271#_c_652_p
+ N_A_955_271#_c_581_n PM_SKY130_FD_SC_LP__DLRBN_1%A_955_271#
x_PM_SKY130_FD_SC_LP__DLRBN_1%A_630_167# N_A_630_167#_M1016_d
+ N_A_630_167#_M1000_d N_A_630_167#_c_740_n N_A_630_167#_c_741_n
+ N_A_630_167#_c_733_n N_A_630_167#_c_734_n N_A_630_167#_c_744_n
+ N_A_630_167#_M1012_g N_A_630_167#_M1008_g N_A_630_167#_c_736_n
+ N_A_630_167#_c_746_n N_A_630_167#_c_737_n N_A_630_167#_c_738_n
+ N_A_630_167#_c_749_n N_A_630_167#_c_750_n N_A_630_167#_c_739_n
+ N_A_630_167#_c_751_n N_A_630_167#_c_752_n N_A_630_167#_c_753_n
+ PM_SKY130_FD_SC_LP__DLRBN_1%A_630_167#
x_PM_SKY130_FD_SC_LP__DLRBN_1%RESET_B N_RESET_B_M1010_g N_RESET_B_M1003_g
+ RESET_B RESET_B N_RESET_B_c_847_n PM_SKY130_FD_SC_LP__DLRBN_1%RESET_B
x_PM_SKY130_FD_SC_LP__DLRBN_1%A_1394_367# N_A_1394_367#_M1023_d
+ N_A_1394_367#_M1020_d N_A_1394_367#_c_885_n N_A_1394_367#_c_886_n
+ N_A_1394_367#_M1002_g N_A_1394_367#_c_893_n N_A_1394_367#_M1022_g
+ N_A_1394_367#_c_888_n N_A_1394_367#_c_889_n N_A_1394_367#_c_895_n
+ N_A_1394_367#_c_896_n N_A_1394_367#_c_890_n
+ PM_SKY130_FD_SC_LP__DLRBN_1%A_1394_367#
x_PM_SKY130_FD_SC_LP__DLRBN_1%VPWR N_VPWR_M1011_s N_VPWR_M1005_d N_VPWR_M1015_d
+ N_VPWR_M1012_s N_VPWR_M1003_d N_VPWR_M1022_d N_VPWR_c_933_n N_VPWR_c_934_n
+ N_VPWR_c_935_n N_VPWR_c_936_n N_VPWR_c_937_n N_VPWR_c_938_n N_VPWR_c_939_n
+ N_VPWR_c_940_n N_VPWR_c_941_n N_VPWR_c_942_n N_VPWR_c_943_n N_VPWR_c_944_n
+ VPWR N_VPWR_c_945_n N_VPWR_c_946_n N_VPWR_c_947_n N_VPWR_c_948_n
+ N_VPWR_c_932_n N_VPWR_c_950_n N_VPWR_c_951_n N_VPWR_c_952_n N_VPWR_c_953_n
+ PM_SKY130_FD_SC_LP__DLRBN_1%VPWR
x_PM_SKY130_FD_SC_LP__DLRBN_1%A_625_377# N_A_625_377#_M1000_s
+ N_A_625_377#_M1004_d N_A_625_377#_c_1051_n N_A_625_377#_c_1052_n
+ N_A_625_377#_c_1053_n PM_SKY130_FD_SC_LP__DLRBN_1%A_625_377#
x_PM_SKY130_FD_SC_LP__DLRBN_1%Q_N N_Q_N_M1002_s N_Q_N_M1022_s Q_N Q_N Q_N Q_N
+ Q_N Q_N N_Q_N_c_1084_n N_Q_N_c_1087_n Q_N PM_SKY130_FD_SC_LP__DLRBN_1%Q_N
x_PM_SKY130_FD_SC_LP__DLRBN_1%Q N_Q_M1006_d N_Q_M1014_d Q Q Q Q Q Q Q
+ N_Q_c_1106_n Q N_Q_c_1110_n PM_SKY130_FD_SC_LP__DLRBN_1%Q
x_PM_SKY130_FD_SC_LP__DLRBN_1%VGND N_VGND_M1009_s N_VGND_M1001_d N_VGND_M1019_d
+ N_VGND_M1010_d N_VGND_M1002_d N_VGND_c_1126_n N_VGND_c_1127_n N_VGND_c_1128_n
+ N_VGND_c_1129_n N_VGND_c_1130_n N_VGND_c_1131_n N_VGND_c_1132_n
+ N_VGND_c_1133_n N_VGND_c_1134_n N_VGND_c_1135_n N_VGND_c_1136_n
+ N_VGND_c_1137_n VGND N_VGND_c_1138_n N_VGND_c_1139_n N_VGND_c_1140_n
+ N_VGND_c_1141_n PM_SKY130_FD_SC_LP__DLRBN_1%VGND
x_PM_SKY130_FD_SC_LP__DLRBN_1%A_547_167# N_A_547_167#_M1016_s
+ N_A_547_167#_M1019_s N_A_547_167#_c_1237_n N_A_547_167#_c_1238_n
+ N_A_547_167#_c_1239_n N_A_547_167#_c_1240_n
+ PM_SKY130_FD_SC_LP__DLRBN_1%A_547_167#
x_PM_SKY130_FD_SC_LP__DLRBN_1%A_716_167# N_A_716_167#_M1007_d
+ N_A_716_167#_M1021_d N_A_716_167#_c_1271_n N_A_716_167#_c_1272_n
+ PM_SKY130_FD_SC_LP__DLRBN_1%A_716_167#
cc_1 VNB N_GATE_N_c_192_n 0.022102f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.698
cc_2 VNB N_GATE_N_M1009_g 0.0445365f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.56
cc_3 VNB GATE_N 0.0352051f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_4 VNB N_GATE_N_c_195_n 0.0247807f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.38
cc_5 VNB N_A_112_70#_c_223_n 0.0189297f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.885
cc_6 VNB N_A_112_70#_c_224_n 0.0164996f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.685
cc_7 VNB N_A_112_70#_M1001_g 0.0309051f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.885
cc_8 VNB N_A_112_70#_M1016_g 0.035836f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.295
cc_9 VNB N_A_112_70#_c_227_n 0.00460666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_112_70#_c_228_n 0.00466966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_112_70#_c_229_n 0.00965323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_112_70#_c_230_n 0.0178332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D_c_352_n 0.0165812f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.402
cc_14 VNB N_D_M1018_g 0.00233236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB D 0.0119524f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.685
cc_16 VNB N_D_c_355_n 0.0399811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_207_40#_c_389_n 0.164319f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.885
cc_18 VNB N_A_207_40#_M1007_g 0.0388819f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_19 VNB N_A_207_40#_c_391_n 0.0296578f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB N_A_207_40#_c_392_n 0.00852207f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_A_207_40#_M1013_g 0.00849196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_207_40#_c_394_n 0.00426883f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.38
cc_23 VNB N_A_207_40#_c_395_n 0.00825676f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.38
cc_24 VNB N_A_207_40#_c_396_n 0.00893918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_207_40#_c_397_n 0.0459997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_437_144#_c_470_n 0.020145f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.685
cc_27 VNB N_A_437_144#_c_471_n 0.00818849f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.685
cc_28 VNB N_A_437_144#_c_472_n 0.00851394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_437_144#_M1015_g 0.0387512f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_A_437_144#_c_474_n 0.0184305f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_31 VNB N_A_437_144#_c_475_n 0.0199386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_437_144#_c_476_n 0.0113835f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.38
cc_33 VNB N_A_437_144#_c_477_n 0.0011428f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.38
cc_34 VNB N_A_437_144#_c_478_n 0.0166005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_437_144#_c_479_n 0.0381256f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=2.035
cc_36 VNB N_A_437_144#_c_480_n 0.00712729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_437_144#_c_481_n 0.0119904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_955_271#_M1021_g 0.0504863f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_39 VNB N_A_955_271#_M1020_g 0.00865726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_955_271#_c_564_n 0.0207247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_955_271#_M1014_g 0.00382998f $X=-0.19 $Y=-0.245 $X2=0.282
+ $Y2=0.925
cc_42 VNB N_A_955_271#_c_566_n 0.0215196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_955_271#_c_567_n 0.00867341f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.38
cc_44 VNB N_A_955_271#_c_568_n 0.0271443f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=2.035
cc_45 VNB N_A_955_271#_c_569_n 0.00746048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_955_271#_c_570_n 0.00760717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_955_271#_c_571_n 0.00285116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_955_271#_c_572_n 0.0382893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_955_271#_c_573_n 0.00508445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_955_271#_c_574_n 0.0278536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_955_271#_c_575_n 0.00316737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_955_271#_c_576_n 0.00119883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_955_271#_c_577_n 0.00140078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_955_271#_c_578_n 0.00781641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_955_271#_c_579_n 0.00647587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_955_271#_c_580_n 0.00182506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_955_271#_c_581_n 0.0407724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_630_167#_c_733_n 0.0142491f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.885
cc_59 VNB N_A_630_167#_c_734_n 0.00645169f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_60 VNB N_A_630_167#_M1008_g 0.0403291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_630_167#_c_736_n 0.00393288f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.38
cc_62 VNB N_A_630_167#_c_737_n 0.0033838f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.215
cc_63 VNB N_A_630_167#_c_738_n 0.00274198f $X=-0.19 $Y=-0.245 $X2=0.282
+ $Y2=0.925
cc_64 VNB N_A_630_167#_c_739_n 0.00570983f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.38
cc_65 VNB N_RESET_B_M1010_g 0.0197179f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.215
cc_66 VNB N_RESET_B_M1003_g 0.0050571f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.885
cc_67 VNB RESET_B 0.0116712f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.885
cc_68 VNB N_RESET_B_c_847_n 0.0288014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1394_367#_c_885_n 0.0199249f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.885
cc_70 VNB N_A_1394_367#_c_886_n 0.0158291f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.685
cc_71 VNB N_A_1394_367#_M1002_g 0.0364127f $X=-0.19 $Y=-0.245 $X2=0.417
+ $Y2=1.885
cc_72 VNB N_A_1394_367#_c_888_n 0.00277644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1394_367#_c_889_n 0.0117223f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.38
cc_74 VNB N_A_1394_367#_c_890_n 0.00544099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VPWR_c_932_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_Q_N_c_1084_n 0.0146502f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.38
cc_77 VNB Q 0.0322008f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.685
cc_78 VNB N_Q_c_1106_n 0.033122f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=0.925
cc_79 VNB Q 0.0122143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1126_n 0.0115566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1127_n 0.0216486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1128_n 0.0121757f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.38
cc_83 VNB N_VGND_c_1129_n 0.00812414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1130_n 0.00737335f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.665
cc_85 VNB N_VGND_c_1131_n 0.0040799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1132_n 0.0370024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1133_n 0.00370274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1134_n 0.0653864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1135_n 0.00452017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1136_n 0.0453329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1137_n 0.00392283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1138_n 0.0402435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1139_n 0.0213558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1140_n 0.503064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1141_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_547_167#_c_1237_n 0.00109937f $X=-0.19 $Y=-0.245 $X2=0.53
+ $Y2=2.685
cc_97 VNB N_A_547_167#_c_1238_n 0.0155274f $X=-0.19 $Y=-0.245 $X2=0.417
+ $Y2=1.885
cc_98 VNB N_A_547_167#_c_1239_n 0.00289297f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=0.84
cc_99 VNB N_A_547_167#_c_1240_n 0.00168833f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_100 VNB N_A_716_167#_c_1271_n 0.034297f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.885
cc_101 VNB N_A_716_167#_c_1272_n 0.0035403f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_102 VPB N_GATE_N_c_192_n 0.00356841f $X=-0.19 $Y=1.655 $X2=0.417 $Y2=1.698
cc_103 VPB N_GATE_N_M1011_g 0.0475085f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.685
cc_104 VPB N_GATE_N_c_198_n 0.02231f $X=-0.19 $Y=1.655 $X2=0.417 $Y2=1.885
cc_105 VPB GATE_N 0.0260762f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_106 VPB N_A_112_70#_c_223_n 0.00991156f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.885
cc_107 VPB N_A_112_70#_M1005_g 0.0222898f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_108 VPB N_A_112_70#_c_233_n 0.0877741f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_112_70#_c_234_n 0.0312511f $X=-0.19 $Y=1.655 $X2=0.417 $Y2=1.38
cc_110 VPB N_A_112_70#_c_235_n 0.0274271f $X=-0.19 $Y=1.655 $X2=0.395 $Y2=1.38
cc_111 VPB N_A_112_70#_c_236_n 0.0380486f $X=-0.19 $Y=1.655 $X2=0.417 $Y2=1.215
cc_112 VPB N_A_112_70#_c_237_n 0.018967f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=1.38
cc_113 VPB N_A_112_70#_c_227_n 0.00179035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_112_70#_c_239_n 0.0334714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_112_70#_c_240_n 0.0057181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_112_70#_c_241_n 0.00157798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_112_70#_c_242_n 0.00228309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_112_70#_c_243_n 0.00418727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_112_70#_c_244_n 0.0185524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_112_70#_c_245_n 0.0452622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_112_70#_c_229_n 3.10815e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_112_70#_c_247_n 0.0458965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_112_70#_c_248_n 0.00423627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_D_M1018_g 0.0220283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_207_40#_M1013_g 0.024507f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_207_40#_c_399_n 0.0156544f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_207_40#_c_396_n 0.0014124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_437_144#_M1015_g 0.0229993f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_129 VPB N_A_437_144#_c_483_n 0.00156215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_437_144#_c_484_n 0.00320112f $X=-0.19 $Y=1.655 $X2=0.282
+ $Y2=1.295
cc_131 VPB N_A_437_144#_c_481_n 0.0034106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_955_271#_M1004_g 0.0240779f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.685
cc_133 VPB N_A_955_271#_M1020_g 0.0274269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_955_271#_M1014_g 0.0240564f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=0.925
cc_135 VPB N_A_955_271#_c_567_n 0.00515678f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=1.38
cc_136 VPB N_A_955_271#_c_568_n 0.00649828f $X=-0.19 $Y=1.655 $X2=0.282
+ $Y2=2.035
cc_137 VPB N_A_955_271#_c_587_n 9.68875e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_955_271#_c_588_n 0.00305352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_630_167#_c_740_n 0.143015f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.885
cc_140 VPB N_A_630_167#_c_741_n 0.0752853f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_630_167#_c_733_n 0.00791211f $X=-0.19 $Y=1.655 $X2=0.417
+ $Y2=1.885
cc_142 VPB N_A_630_167#_c_734_n 0.00242399f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_143 VPB N_A_630_167#_c_744_n 0.0182543f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_144 VPB N_A_630_167#_c_736_n 0.00336318f $X=-0.19 $Y=1.655 $X2=0.417 $Y2=1.38
cc_145 VPB N_A_630_167#_c_746_n 0.00491209f $X=-0.19 $Y=1.655 $X2=0.395 $Y2=1.38
cc_146 VPB N_A_630_167#_c_737_n 0.00268534f $X=-0.19 $Y=1.655 $X2=0.417
+ $Y2=1.215
cc_147 VPB N_A_630_167#_c_738_n 3.3304e-19 $X=-0.19 $Y=1.655 $X2=0.282 $Y2=0.925
cc_148 VPB N_A_630_167#_c_749_n 0.00481963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_630_167#_c_750_n 0.00136352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_630_167#_c_751_n 0.0032639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_630_167#_c_752_n 0.0465026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_630_167#_c_753_n 0.00512984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_M1003_g 0.022415f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.885
cc_154 VPB RESET_B 0.00640611f $X=-0.19 $Y=1.655 $X2=0.417 $Y2=1.885
cc_155 VPB N_A_1394_367#_c_885_n 0.0105465f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.885
cc_156 VPB N_A_1394_367#_c_886_n 0.00422854f $X=-0.19 $Y=1.655 $X2=0.53
+ $Y2=2.685
cc_157 VPB N_A_1394_367#_c_893_n 0.0192638f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_158 VPB N_A_1394_367#_c_888_n 0.00251798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_1394_367#_c_895_n 0.0507882f $X=-0.19 $Y=1.655 $X2=0.395 $Y2=1.38
cc_160 VPB N_A_1394_367#_c_896_n 0.0280602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_933_n 0.0127766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_934_n 0.0354917f $X=-0.19 $Y=1.655 $X2=0.395 $Y2=1.38
cc_163 VPB N_VPWR_c_935_n 0.00314186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_936_n 0.0165005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_937_n 0.0243457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_938_n 0.0124552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_939_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_940_n 0.0268023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_941_n 0.00519757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_942_n 0.00502248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_943_n 0.0260919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_944_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_945_n 0.0340688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_946_n 0.0609364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_947_n 0.0432117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_948_n 0.0286786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_932_n 0.087856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_950_n 0.00601091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_951_n 0.00583335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_952_n 0.00680245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_953_n 0.00382116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_625_377#_c_1051_n 0.0240908f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.885
cc_183 VPB N_A_625_377#_c_1052_n 0.00235746f $X=-0.19 $Y=1.655 $X2=0.53
+ $Y2=2.685
cc_184 VPB N_A_625_377#_c_1053_n 0.00651766f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.58
cc_185 VPB Q_N 9.53061e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_Q_N_c_1084_n 0.00170261f $X=-0.19 $Y=1.655 $X2=0.395 $Y2=1.38
cc_187 VPB N_Q_N_c_1087_n 0.0274747f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=2.035
cc_188 VPB Q 0.0107868f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.685
cc_189 VPB Q 0.0567505f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_190 VPB N_Q_c_1110_n 0.0266415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 N_GATE_N_c_192_n N_A_112_70#_c_224_n 0.0202872f $X=0.417 $Y=1.698 $X2=0
+ $Y2=0
cc_192 GATE_N N_A_112_70#_c_224_n 5.22485e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_193 N_GATE_N_c_198_n N_A_112_70#_c_241_n 0.00490506f $X=0.417 $Y=1.885 $X2=0
+ $Y2=0
cc_194 N_GATE_N_M1011_g N_A_112_70#_c_242_n 0.00162302f $X=0.53 $Y=2.685 $X2=0
+ $Y2=0
cc_195 N_GATE_N_c_192_n N_A_112_70#_c_229_n 0.00490506f $X=0.417 $Y=1.698 $X2=0
+ $Y2=0
cc_196 N_GATE_N_c_198_n N_A_112_70#_c_247_n 0.0202872f $X=0.417 $Y=1.885 $X2=0
+ $Y2=0
cc_197 N_GATE_N_M1009_g N_A_112_70#_c_230_n 0.0135329f $X=0.485 $Y=0.56 $X2=0
+ $Y2=0
cc_198 GATE_N N_A_112_70#_c_230_n 0.100563f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_199 N_GATE_N_c_195_n N_A_112_70#_c_230_n 0.00490506f $X=0.395 $Y=1.38 $X2=0
+ $Y2=0
cc_200 N_GATE_N_M1011_g N_A_112_70#_c_248_n 0.00490506f $X=0.53 $Y=2.685 $X2=0
+ $Y2=0
cc_201 N_GATE_N_M1009_g N_A_207_40#_c_394_n 2.81049e-19 $X=0.485 $Y=0.56 $X2=0
+ $Y2=0
cc_202 N_GATE_N_M1009_g N_A_207_40#_c_397_n 0.00501689f $X=0.485 $Y=0.56 $X2=0
+ $Y2=0
cc_203 N_GATE_N_M1011_g N_VPWR_c_934_n 0.0132876f $X=0.53 $Y=2.685 $X2=0 $Y2=0
cc_204 N_GATE_N_c_198_n N_VPWR_c_934_n 9.38971e-19 $X=0.417 $Y=1.885 $X2=0 $Y2=0
cc_205 GATE_N N_VPWR_c_934_n 0.0305154f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_206 N_GATE_N_M1011_g N_VPWR_c_945_n 0.00414769f $X=0.53 $Y=2.685 $X2=0 $Y2=0
cc_207 N_GATE_N_M1011_g N_VPWR_c_932_n 0.00837493f $X=0.53 $Y=2.685 $X2=0 $Y2=0
cc_208 N_GATE_N_M1009_g N_VGND_c_1127_n 0.00934546f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_209 GATE_N N_VGND_c_1127_n 0.0266999f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_210 N_GATE_N_c_195_n N_VGND_c_1127_n 5.61365e-19 $X=0.395 $Y=1.38 $X2=0 $Y2=0
cc_211 N_GATE_N_M1009_g N_VGND_c_1132_n 0.00396895f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_212 N_GATE_N_M1009_g N_VGND_c_1140_n 0.00645901f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_213 GATE_N N_VGND_c_1140_n 0.00340156f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_214 N_A_112_70#_M1001_g N_D_c_352_n 0.0126027f $X=1.68 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A_112_70#_c_233_n N_D_M1018_g 0.00543798f $X=2.71 $Y=3.03 $X2=0 $Y2=0
cc_216 N_A_112_70#_c_227_n N_D_M1018_g 0.0205907f $X=1.695 $Y=1.58 $X2=0 $Y2=0
cc_217 N_A_112_70#_c_239_n N_D_M1018_g 0.0177037f $X=3.075 $Y=1.735 $X2=0 $Y2=0
cc_218 N_A_112_70#_c_223_n D 0.00187322f $X=1.605 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A_112_70#_M1001_g D 0.0175092f $X=1.68 $Y=0.93 $X2=0 $Y2=0
cc_220 N_A_112_70#_c_227_n D 0.0094504f $X=1.695 $Y=1.58 $X2=0 $Y2=0
cc_221 N_A_112_70#_M1001_g N_D_c_355_n 0.0139513f $X=1.68 $Y=0.93 $X2=0 $Y2=0
cc_222 N_A_112_70#_M1016_g N_D_c_355_n 0.00472031f $X=3.075 $Y=1.045 $X2=0 $Y2=0
cc_223 N_A_112_70#_c_227_n N_D_c_355_n 0.00490114f $X=1.695 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A_112_70#_M1001_g N_A_207_40#_c_389_n 0.00912785f $X=1.68 $Y=0.93 $X2=0
+ $Y2=0
cc_225 N_A_112_70#_M1016_g N_A_207_40#_c_389_n 0.00497235f $X=3.075 $Y=1.045
+ $X2=0 $Y2=0
cc_226 N_A_112_70#_M1016_g N_A_207_40#_M1007_g 0.0192721f $X=3.075 $Y=1.045
+ $X2=0 $Y2=0
cc_227 N_A_112_70#_c_237_n N_A_207_40#_c_392_n 0.00741578f $X=3.465 $Y=2.415
+ $X2=0 $Y2=0
cc_228 N_A_112_70#_c_237_n N_A_207_40#_M1013_g 0.0198677f $X=3.465 $Y=2.415
+ $X2=0 $Y2=0
cc_229 N_A_112_70#_M1001_g N_A_207_40#_c_394_n 0.00306523f $X=1.68 $Y=0.93 $X2=0
+ $Y2=0
cc_230 N_A_112_70#_c_228_n N_A_207_40#_c_394_n 0.0288034f $X=0.7 $Y=0.505 $X2=0
+ $Y2=0
cc_231 N_A_112_70#_c_223_n N_A_207_40#_c_395_n 0.00422331f $X=1.605 $Y=1.58
+ $X2=0 $Y2=0
cc_232 N_A_112_70#_c_224_n N_A_207_40#_c_395_n 0.00645718f $X=1.145 $Y=1.58
+ $X2=0 $Y2=0
cc_233 N_A_112_70#_M1001_g N_A_207_40#_c_395_n 0.00359333f $X=1.68 $Y=0.93 $X2=0
+ $Y2=0
cc_234 N_A_112_70#_c_229_n N_A_207_40#_c_395_n 0.0011917f $X=0.98 $Y=1.67 $X2=0
+ $Y2=0
cc_235 N_A_112_70#_c_230_n N_A_207_40#_c_395_n 0.0201976f $X=0.862 $Y=1.505
+ $X2=0 $Y2=0
cc_236 N_A_112_70#_c_223_n N_A_207_40#_c_399_n 0.005599f $X=1.605 $Y=1.58 $X2=0
+ $Y2=0
cc_237 N_A_112_70#_M1005_g N_A_207_40#_c_399_n 0.00843289f $X=1.71 $Y=2.115
+ $X2=0 $Y2=0
cc_238 N_A_112_70#_c_241_n N_A_207_40#_c_399_n 0.016915f $X=0.862 $Y=1.973 $X2=0
+ $Y2=0
cc_239 N_A_112_70#_c_243_n N_A_207_40#_c_399_n 0.0125699f $X=0.745 $Y=2.52 $X2=0
+ $Y2=0
cc_240 N_A_112_70#_c_244_n N_A_207_40#_c_399_n 0.0221854f $X=1.57 $Y=2.94 $X2=0
+ $Y2=0
cc_241 N_A_112_70#_c_245_n N_A_207_40#_c_399_n 0.00496547f $X=1.57 $Y=2.94 $X2=0
+ $Y2=0
cc_242 N_A_112_70#_c_248_n N_A_207_40#_c_399_n 0.016915f $X=0.862 $Y=2.175 $X2=0
+ $Y2=0
cc_243 N_A_112_70#_c_223_n N_A_207_40#_c_396_n 0.0165891f $X=1.605 $Y=1.58 $X2=0
+ $Y2=0
cc_244 N_A_112_70#_M1001_g N_A_207_40#_c_396_n 0.00553663f $X=1.68 $Y=0.93 $X2=0
+ $Y2=0
cc_245 N_A_112_70#_M1005_g N_A_207_40#_c_396_n 0.00148992f $X=1.71 $Y=2.115
+ $X2=0 $Y2=0
cc_246 N_A_112_70#_c_229_n N_A_207_40#_c_396_n 0.016915f $X=0.98 $Y=1.67 $X2=0
+ $Y2=0
cc_247 N_A_112_70#_c_247_n N_A_207_40#_c_396_n 0.00551148f $X=0.98 $Y=1.67 $X2=0
+ $Y2=0
cc_248 N_A_112_70#_c_230_n N_A_207_40#_c_396_n 0.0190938f $X=0.862 $Y=1.505
+ $X2=0 $Y2=0
cc_249 N_A_112_70#_c_228_n N_A_207_40#_c_397_n 0.00162645f $X=0.7 $Y=0.505 $X2=0
+ $Y2=0
cc_250 N_A_112_70#_c_239_n N_A_437_144#_c_483_n 0.00270435f $X=3.075 $Y=1.735
+ $X2=0 $Y2=0
cc_251 N_A_112_70#_c_233_n N_A_437_144#_c_484_n 0.00569216f $X=2.71 $Y=3.03
+ $X2=0 $Y2=0
cc_252 N_A_112_70#_c_234_n N_A_437_144#_c_484_n 0.00270435f $X=2.785 $Y=2.415
+ $X2=0 $Y2=0
cc_253 N_A_112_70#_M1016_g N_A_437_144#_c_478_n 3.91393e-19 $X=3.075 $Y=1.045
+ $X2=0 $Y2=0
cc_254 N_A_112_70#_M1016_g N_A_437_144#_c_480_n 7.50042e-19 $X=3.075 $Y=1.045
+ $X2=0 $Y2=0
cc_255 N_A_112_70#_M1016_g N_A_437_144#_c_481_n 0.00315604f $X=3.075 $Y=1.045
+ $X2=0 $Y2=0
cc_256 N_A_112_70#_c_239_n N_A_437_144#_c_481_n 9.73048e-19 $X=3.075 $Y=1.735
+ $X2=0 $Y2=0
cc_257 N_A_112_70#_c_234_n N_A_630_167#_c_746_n 0.012425f $X=2.785 $Y=2.415
+ $X2=0 $Y2=0
cc_258 N_A_112_70#_c_236_n N_A_630_167#_c_746_n 7.7907e-19 $X=3.39 $Y=2.49 $X2=0
+ $Y2=0
cc_259 N_A_112_70#_c_237_n N_A_630_167#_c_746_n 0.0037207f $X=3.465 $Y=2.415
+ $X2=0 $Y2=0
cc_260 N_A_112_70#_c_239_n N_A_630_167#_c_746_n 0.00886283f $X=3.075 $Y=1.735
+ $X2=0 $Y2=0
cc_261 N_A_112_70#_M1016_g N_A_630_167#_c_737_n 0.013314f $X=3.075 $Y=1.045
+ $X2=0 $Y2=0
cc_262 N_A_112_70#_c_239_n N_A_630_167#_c_737_n 0.00805465f $X=3.075 $Y=1.735
+ $X2=0 $Y2=0
cc_263 N_A_112_70#_c_239_n N_A_630_167#_c_738_n 0.00352393f $X=3.075 $Y=1.735
+ $X2=0 $Y2=0
cc_264 N_A_112_70#_c_236_n N_A_630_167#_c_749_n 0.015858f $X=3.39 $Y=2.49 $X2=0
+ $Y2=0
cc_265 N_A_112_70#_c_239_n N_A_630_167#_c_749_n 0.00100592f $X=3.075 $Y=1.735
+ $X2=0 $Y2=0
cc_266 N_A_112_70#_c_235_n N_A_630_167#_c_750_n 0.00812943f $X=2.785 $Y=2.955
+ $X2=0 $Y2=0
cc_267 N_A_112_70#_c_236_n N_A_630_167#_c_750_n 0.00311662f $X=3.39 $Y=2.49
+ $X2=0 $Y2=0
cc_268 N_A_112_70#_c_240_n N_A_630_167#_c_750_n 0.00270255f $X=2.785 $Y=2.49
+ $X2=0 $Y2=0
cc_269 N_A_112_70#_M1016_g N_A_630_167#_c_739_n 0.0035367f $X=3.075 $Y=1.045
+ $X2=0 $Y2=0
cc_270 N_A_112_70#_c_235_n N_A_630_167#_c_751_n 0.00349639f $X=2.785 $Y=2.955
+ $X2=0 $Y2=0
cc_271 N_A_112_70#_c_235_n N_A_630_167#_c_752_n 0.0096447f $X=2.785 $Y=2.955
+ $X2=0 $Y2=0
cc_272 N_A_112_70#_c_236_n N_A_630_167#_c_752_n 0.0126758f $X=3.39 $Y=2.49 $X2=0
+ $Y2=0
cc_273 N_A_112_70#_c_236_n N_A_630_167#_c_753_n 0.0106888f $X=3.39 $Y=2.49 $X2=0
+ $Y2=0
cc_274 N_A_112_70#_c_237_n N_A_630_167#_c_753_n 0.00321361f $X=3.465 $Y=2.415
+ $X2=0 $Y2=0
cc_275 N_A_112_70#_c_242_n N_VPWR_c_934_n 0.0138892f $X=0.755 $Y=2.775 $X2=0
+ $Y2=0
cc_276 N_A_112_70#_c_243_n N_VPWR_c_934_n 0.01611f $X=0.745 $Y=2.52 $X2=0 $Y2=0
cc_277 N_A_112_70#_M1005_g N_VPWR_c_935_n 0.00768166f $X=1.71 $Y=2.115 $X2=0
+ $Y2=0
cc_278 N_A_112_70#_c_233_n N_VPWR_c_936_n 0.0285459f $X=2.71 $Y=3.03 $X2=0 $Y2=0
cc_279 N_A_112_70#_c_244_n N_VPWR_c_936_n 0.0245744f $X=1.57 $Y=2.94 $X2=0 $Y2=0
cc_280 N_A_112_70#_c_245_n N_VPWR_c_936_n 0.00132938f $X=1.57 $Y=2.94 $X2=0
+ $Y2=0
cc_281 N_A_112_70#_c_233_n N_VPWR_c_942_n 0.00144467f $X=2.71 $Y=3.03 $X2=0
+ $Y2=0
cc_282 N_A_112_70#_c_235_n N_VPWR_c_942_n 0.00908065f $X=2.785 $Y=2.955 $X2=0
+ $Y2=0
cc_283 N_A_112_70#_c_240_n N_VPWR_c_942_n 4.83768e-19 $X=2.785 $Y=2.49 $X2=0
+ $Y2=0
cc_284 N_A_112_70#_c_242_n N_VPWR_c_945_n 0.0135843f $X=0.755 $Y=2.775 $X2=0
+ $Y2=0
cc_285 N_A_112_70#_c_244_n N_VPWR_c_945_n 0.0582626f $X=1.57 $Y=2.94 $X2=0 $Y2=0
cc_286 N_A_112_70#_c_245_n N_VPWR_c_945_n 0.0100221f $X=1.57 $Y=2.94 $X2=0 $Y2=0
cc_287 N_A_112_70#_c_233_n N_VPWR_c_946_n 0.0173898f $X=2.71 $Y=3.03 $X2=0 $Y2=0
cc_288 N_A_112_70#_c_236_n N_VPWR_c_946_n 0.0015473f $X=3.39 $Y=2.49 $X2=0 $Y2=0
cc_289 N_A_112_70#_M1005_g N_VPWR_c_932_n 2.80608e-19 $X=1.71 $Y=2.115 $X2=0
+ $Y2=0
cc_290 N_A_112_70#_c_233_n N_VPWR_c_932_n 0.0358482f $X=2.71 $Y=3.03 $X2=0 $Y2=0
cc_291 N_A_112_70#_c_242_n N_VPWR_c_932_n 0.00738148f $X=0.755 $Y=2.775 $X2=0
+ $Y2=0
cc_292 N_A_112_70#_c_244_n N_VPWR_c_932_n 0.0321842f $X=1.57 $Y=2.94 $X2=0 $Y2=0
cc_293 N_A_112_70#_c_245_n N_VPWR_c_932_n 0.0077944f $X=1.57 $Y=2.94 $X2=0 $Y2=0
cc_294 N_A_112_70#_c_237_n N_A_625_377#_c_1051_n 0.0117889f $X=3.465 $Y=2.415
+ $X2=0 $Y2=0
cc_295 N_A_112_70#_c_234_n N_A_625_377#_c_1052_n 0.00109986f $X=2.785 $Y=2.415
+ $X2=0 $Y2=0
cc_296 N_A_112_70#_c_236_n N_A_625_377#_c_1052_n 0.0031227f $X=3.39 $Y=2.49
+ $X2=0 $Y2=0
cc_297 N_A_112_70#_c_237_n N_A_625_377#_c_1052_n 4.85854e-19 $X=3.465 $Y=2.415
+ $X2=0 $Y2=0
cc_298 N_A_112_70#_c_239_n N_A_625_377#_c_1052_n 2.10991e-19 $X=3.075 $Y=1.735
+ $X2=0 $Y2=0
cc_299 N_A_112_70#_c_228_n N_VGND_c_1127_n 0.0127357f $X=0.7 $Y=0.505 $X2=0
+ $Y2=0
cc_300 N_A_112_70#_M1001_g N_VGND_c_1128_n 0.00144005f $X=1.68 $Y=0.93 $X2=0
+ $Y2=0
cc_301 N_A_112_70#_c_228_n N_VGND_c_1132_n 0.0102398f $X=0.7 $Y=0.505 $X2=0
+ $Y2=0
cc_302 N_A_112_70#_M1001_g N_VGND_c_1140_n 8.46057e-19 $X=1.68 $Y=0.93 $X2=0
+ $Y2=0
cc_303 N_A_112_70#_c_228_n N_VGND_c_1140_n 0.00823993f $X=0.7 $Y=0.505 $X2=0
+ $Y2=0
cc_304 N_A_112_70#_M1016_g N_A_547_167#_c_1237_n 0.00278796f $X=3.075 $Y=1.045
+ $X2=0 $Y2=0
cc_305 N_A_112_70#_c_239_n N_A_547_167#_c_1237_n 0.00196226f $X=3.075 $Y=1.735
+ $X2=0 $Y2=0
cc_306 N_A_112_70#_M1016_g N_A_547_167#_c_1238_n 0.0108629f $X=3.075 $Y=1.045
+ $X2=0 $Y2=0
cc_307 N_D_c_352_n N_A_207_40#_c_389_n 0.00924127f $X=2.11 $Y=1.25 $X2=0 $Y2=0
cc_308 D N_A_207_40#_c_395_n 0.00269322f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_309 D N_A_207_40#_c_399_n 0.00553005f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_310 D N_A_207_40#_c_396_n 0.0304267f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_311 N_D_c_352_n N_A_437_144#_c_476_n 0.00238045f $X=2.11 $Y=1.25 $X2=0 $Y2=0
cc_312 N_D_M1018_g N_A_437_144#_c_483_n 0.00477618f $X=2.295 $Y=2.115 $X2=0
+ $Y2=0
cc_313 N_D_c_352_n N_A_437_144#_c_480_n 2.12546e-19 $X=2.11 $Y=1.25 $X2=0 $Y2=0
cc_314 D N_A_437_144#_c_480_n 0.00327486f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_315 N_D_c_355_n N_A_437_144#_c_480_n 0.0051934f $X=2.295 $Y=1.415 $X2=0 $Y2=0
cc_316 N_D_c_352_n N_A_437_144#_c_481_n 0.00518717f $X=2.11 $Y=1.25 $X2=0 $Y2=0
cc_317 D N_A_437_144#_c_481_n 0.0295473f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_318 N_D_c_355_n N_A_437_144#_c_481_n 0.00477618f $X=2.295 $Y=1.415 $X2=0
+ $Y2=0
cc_319 N_D_M1018_g N_A_630_167#_c_750_n 3.93277e-19 $X=2.295 $Y=2.115 $X2=0
+ $Y2=0
cc_320 N_D_M1018_g N_VPWR_c_935_n 0.00413371f $X=2.295 $Y=2.115 $X2=0 $Y2=0
cc_321 D N_VPWR_c_935_n 0.0258284f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_322 N_D_c_355_n N_VPWR_c_935_n 0.00438271f $X=2.295 $Y=1.415 $X2=0 $Y2=0
cc_323 N_D_M1018_g N_VPWR_c_942_n 0.0058124f $X=2.295 $Y=2.115 $X2=0 $Y2=0
cc_324 N_D_M1018_g N_VPWR_c_932_n 7.14123e-19 $X=2.295 $Y=2.115 $X2=0 $Y2=0
cc_325 N_D_c_352_n N_VGND_c_1128_n 0.00146441f $X=2.11 $Y=1.25 $X2=0 $Y2=0
cc_326 D N_VGND_c_1128_n 0.0167238f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_327 N_D_c_352_n N_VGND_c_1140_n 8.46057e-19 $X=2.11 $Y=1.25 $X2=0 $Y2=0
cc_328 N_D_c_352_n N_A_547_167#_c_1239_n 2.70816e-19 $X=2.11 $Y=1.25 $X2=0 $Y2=0
cc_329 N_A_207_40#_M1007_g N_A_437_144#_c_470_n 0.0144792f $X=3.505 $Y=1.045
+ $X2=0 $Y2=0
cc_330 N_A_207_40#_c_391_n N_A_437_144#_c_472_n 0.00334519f $X=3.915 $Y=1.44
+ $X2=0 $Y2=0
cc_331 N_A_207_40#_M1007_g N_A_437_144#_M1015_g 0.00411158f $X=3.505 $Y=1.045
+ $X2=0 $Y2=0
cc_332 N_A_207_40#_c_391_n N_A_437_144#_M1015_g 0.0816859f $X=3.915 $Y=1.44
+ $X2=0 $Y2=0
cc_333 N_A_207_40#_c_389_n N_A_437_144#_c_477_n 0.00799522f $X=3.43 $Y=0.275
+ $X2=0 $Y2=0
cc_334 N_A_207_40#_c_389_n N_A_437_144#_c_478_n 0.0270563f $X=3.43 $Y=0.275
+ $X2=0 $Y2=0
cc_335 N_A_207_40#_M1007_g N_A_437_144#_c_478_n 0.00596851f $X=3.505 $Y=1.045
+ $X2=0 $Y2=0
cc_336 N_A_207_40#_c_389_n N_A_437_144#_c_479_n 0.0214373f $X=3.43 $Y=0.275
+ $X2=0 $Y2=0
cc_337 N_A_207_40#_c_389_n N_A_437_144#_c_480_n 0.00509328f $X=3.43 $Y=0.275
+ $X2=0 $Y2=0
cc_338 N_A_207_40#_M1013_g N_A_630_167#_c_740_n 0.00710878f $X=3.99 $Y=2.205
+ $X2=0 $Y2=0
cc_339 N_A_207_40#_M1013_g N_A_630_167#_c_737_n 0.00465922f $X=3.99 $Y=2.205
+ $X2=0 $Y2=0
cc_340 N_A_207_40#_M1007_g N_A_630_167#_c_739_n 0.00683395f $X=3.505 $Y=1.045
+ $X2=0 $Y2=0
cc_341 N_A_207_40#_M1013_g N_A_630_167#_c_753_n 0.0105665f $X=3.99 $Y=2.205
+ $X2=0 $Y2=0
cc_342 N_A_207_40#_c_399_n N_VPWR_c_935_n 0.0136775f $X=1.495 $Y=1.94 $X2=0
+ $Y2=0
cc_343 N_A_207_40#_M1013_g N_VPWR_c_937_n 0.00125133f $X=3.99 $Y=2.205 $X2=0
+ $Y2=0
cc_344 N_A_207_40#_c_399_n N_VPWR_c_942_n 0.0136775f $X=1.495 $Y=1.94 $X2=0
+ $Y2=0
cc_345 N_A_207_40#_M1013_g N_VPWR_c_932_n 6.98653e-19 $X=3.99 $Y=2.205 $X2=0
+ $Y2=0
cc_346 N_A_207_40#_c_392_n N_A_625_377#_c_1051_n 0.0116064f $X=3.58 $Y=1.44
+ $X2=0 $Y2=0
cc_347 N_A_207_40#_M1013_g N_A_625_377#_c_1051_n 0.0182637f $X=3.99 $Y=2.205
+ $X2=0 $Y2=0
cc_348 N_A_207_40#_c_394_n N_VGND_c_1127_n 0.00158623f $X=1.2 $Y=0.365 $X2=0
+ $Y2=0
cc_349 N_A_207_40#_c_397_n N_VGND_c_1127_n 9.20395e-19 $X=1.2 $Y=0.275 $X2=0
+ $Y2=0
cc_350 N_A_207_40#_c_389_n N_VGND_c_1128_n 0.0207771f $X=3.43 $Y=0.275 $X2=0
+ $Y2=0
cc_351 N_A_207_40#_c_394_n N_VGND_c_1128_n 0.0179734f $X=1.2 $Y=0.365 $X2=0
+ $Y2=0
cc_352 N_A_207_40#_c_397_n N_VGND_c_1128_n 0.00335098f $X=1.2 $Y=0.275 $X2=0
+ $Y2=0
cc_353 N_A_207_40#_c_394_n N_VGND_c_1132_n 0.0191905f $X=1.2 $Y=0.365 $X2=0
+ $Y2=0
cc_354 N_A_207_40#_c_395_n N_VGND_c_1132_n 0.00332971f $X=1.33 $Y=0.9 $X2=0
+ $Y2=0
cc_355 N_A_207_40#_c_397_n N_VGND_c_1132_n 0.0168486f $X=1.2 $Y=0.275 $X2=0
+ $Y2=0
cc_356 N_A_207_40#_c_389_n N_VGND_c_1134_n 0.0299964f $X=3.43 $Y=0.275 $X2=0
+ $Y2=0
cc_357 N_A_207_40#_c_389_n N_VGND_c_1140_n 0.0539656f $X=3.43 $Y=0.275 $X2=0
+ $Y2=0
cc_358 N_A_207_40#_c_394_n N_VGND_c_1140_n 0.0110719f $X=1.2 $Y=0.365 $X2=0
+ $Y2=0
cc_359 N_A_207_40#_c_395_n N_VGND_c_1140_n 0.00600796f $X=1.33 $Y=0.9 $X2=0
+ $Y2=0
cc_360 N_A_207_40#_c_397_n N_VGND_c_1140_n 0.0083401f $X=1.2 $Y=0.275 $X2=0
+ $Y2=0
cc_361 N_A_207_40#_c_389_n N_A_547_167#_c_1238_n 0.00206418f $X=3.43 $Y=0.275
+ $X2=0 $Y2=0
cc_362 N_A_207_40#_M1007_g N_A_547_167#_c_1238_n 0.015939f $X=3.505 $Y=1.045
+ $X2=0 $Y2=0
cc_363 N_A_207_40#_c_389_n N_A_547_167#_c_1239_n 0.0014299f $X=3.43 $Y=0.275
+ $X2=0 $Y2=0
cc_364 N_A_207_40#_M1007_g N_A_716_167#_c_1271_n 0.00365144f $X=3.505 $Y=1.045
+ $X2=0 $Y2=0
cc_365 N_A_207_40#_c_391_n N_A_716_167#_c_1271_n 0.0151127f $X=3.915 $Y=1.44
+ $X2=0 $Y2=0
cc_366 N_A_437_144#_M1015_g N_A_955_271#_M1004_g 0.0191257f $X=4.35 $Y=2.205
+ $X2=0 $Y2=0
cc_367 N_A_437_144#_M1015_g N_A_955_271#_M1021_g 0.00768641f $X=4.35 $Y=2.205
+ $X2=0 $Y2=0
cc_368 N_A_437_144#_c_474_n N_A_955_271#_M1021_g 0.0184037f $X=4.6 $Y=0.875
+ $X2=0 $Y2=0
cc_369 N_A_437_144#_M1015_g N_A_955_271#_c_567_n 0.00193568f $X=4.35 $Y=2.205
+ $X2=0 $Y2=0
cc_370 N_A_437_144#_M1015_g N_A_955_271#_c_568_n 0.0103745f $X=4.35 $Y=2.205
+ $X2=0 $Y2=0
cc_371 N_A_437_144#_M1015_g N_A_630_167#_c_740_n 0.00720868f $X=4.35 $Y=2.205
+ $X2=0 $Y2=0
cc_372 N_A_437_144#_c_483_n N_A_630_167#_c_746_n 0.0464588f $X=2.525 $Y=1.875
+ $X2=0 $Y2=0
cc_373 N_A_437_144#_c_481_n N_A_630_167#_c_746_n 0.00563541f $X=2.525 $Y=1.775
+ $X2=0 $Y2=0
cc_374 N_A_437_144#_c_481_n N_A_630_167#_c_738_n 0.0125371f $X=2.525 $Y=1.775
+ $X2=0 $Y2=0
cc_375 N_A_437_144#_c_484_n N_A_630_167#_c_750_n 0.00120602f $X=2.51 $Y=1.94
+ $X2=0 $Y2=0
cc_376 N_A_437_144#_c_481_n N_A_630_167#_c_739_n 0.00931683f $X=2.525 $Y=1.775
+ $X2=0 $Y2=0
cc_377 N_A_437_144#_M1015_g N_A_630_167#_c_753_n 0.0012503f $X=4.35 $Y=2.205
+ $X2=0 $Y2=0
cc_378 N_A_437_144#_c_483_n N_VPWR_c_935_n 0.001132f $X=2.525 $Y=1.875 $X2=0
+ $Y2=0
cc_379 N_A_437_144#_M1015_g N_VPWR_c_937_n 0.0109945f $X=4.35 $Y=2.205 $X2=0
+ $Y2=0
cc_380 N_A_437_144#_c_484_n N_VPWR_c_942_n 7.03867e-19 $X=2.51 $Y=1.94 $X2=0
+ $Y2=0
cc_381 N_A_437_144#_M1015_g N_VPWR_c_932_n 7.04242e-19 $X=4.35 $Y=2.205 $X2=0
+ $Y2=0
cc_382 N_A_437_144#_M1015_g N_A_625_377#_c_1051_n 0.0186725f $X=4.35 $Y=2.205
+ $X2=0 $Y2=0
cc_383 N_A_437_144#_M1015_g N_A_625_377#_c_1053_n 6.85495e-19 $X=4.35 $Y=2.205
+ $X2=0 $Y2=0
cc_384 N_A_437_144#_c_476_n N_VGND_c_1128_n 0.0115517f $X=2.51 $Y=0.71 $X2=0
+ $Y2=0
cc_385 N_A_437_144#_c_477_n N_VGND_c_1128_n 0.00726747f $X=2.595 $Y=0.35 $X2=0
+ $Y2=0
cc_386 N_A_437_144#_c_480_n N_VGND_c_1128_n 6.59308e-19 $X=2.51 $Y=0.875 $X2=0
+ $Y2=0
cc_387 N_A_437_144#_c_474_n N_VGND_c_1129_n 0.00239898f $X=4.6 $Y=0.875 $X2=0
+ $Y2=0
cc_388 N_A_437_144#_c_478_n N_VGND_c_1129_n 0.00326002f $X=3.955 $Y=0.35 $X2=0
+ $Y2=0
cc_389 N_A_437_144#_c_479_n N_VGND_c_1129_n 5.37535e-19 $X=3.955 $Y=0.35 $X2=0
+ $Y2=0
cc_390 N_A_437_144#_c_474_n N_VGND_c_1134_n 0.00482246f $X=4.6 $Y=0.875 $X2=0
+ $Y2=0
cc_391 N_A_437_144#_c_477_n N_VGND_c_1134_n 0.0105537f $X=2.595 $Y=0.35 $X2=0
+ $Y2=0
cc_392 N_A_437_144#_c_478_n N_VGND_c_1134_n 0.0886522f $X=3.955 $Y=0.35 $X2=0
+ $Y2=0
cc_393 N_A_437_144#_c_479_n N_VGND_c_1134_n 0.00651318f $X=3.955 $Y=0.35 $X2=0
+ $Y2=0
cc_394 N_A_437_144#_c_480_n N_VGND_c_1134_n 0.00387311f $X=2.51 $Y=0.875 $X2=0
+ $Y2=0
cc_395 N_A_437_144#_c_474_n N_VGND_c_1140_n 0.00949844f $X=4.6 $Y=0.875 $X2=0
+ $Y2=0
cc_396 N_A_437_144#_c_477_n N_VGND_c_1140_n 0.00572329f $X=2.595 $Y=0.35 $X2=0
+ $Y2=0
cc_397 N_A_437_144#_c_478_n N_VGND_c_1140_n 0.0509374f $X=3.955 $Y=0.35 $X2=0
+ $Y2=0
cc_398 N_A_437_144#_c_479_n N_VGND_c_1140_n 0.0093478f $X=3.955 $Y=0.35 $X2=0
+ $Y2=0
cc_399 N_A_437_144#_c_480_n N_VGND_c_1140_n 0.00561723f $X=2.51 $Y=0.875 $X2=0
+ $Y2=0
cc_400 N_A_437_144#_c_480_n N_A_547_167#_c_1237_n 0.0214807f $X=2.51 $Y=0.875
+ $X2=0 $Y2=0
cc_401 N_A_437_144#_c_481_n N_A_547_167#_c_1237_n 0.0128389f $X=2.525 $Y=1.775
+ $X2=0 $Y2=0
cc_402 N_A_437_144#_c_470_n N_A_547_167#_c_1238_n 0.010692f $X=4.045 $Y=0.875
+ $X2=0 $Y2=0
cc_403 N_A_437_144#_c_471_n N_A_547_167#_c_1238_n 0.00176034f $X=4.275 $Y=0.95
+ $X2=0 $Y2=0
cc_404 N_A_437_144#_c_478_n N_A_547_167#_c_1238_n 0.0773815f $X=3.955 $Y=0.35
+ $X2=0 $Y2=0
cc_405 N_A_437_144#_c_479_n N_A_547_167#_c_1238_n 0.0044365f $X=3.955 $Y=0.35
+ $X2=0 $Y2=0
cc_406 N_A_437_144#_c_476_n N_A_547_167#_c_1239_n 0.00886831f $X=2.51 $Y=0.71
+ $X2=0 $Y2=0
cc_407 N_A_437_144#_c_478_n N_A_547_167#_c_1239_n 0.0176524f $X=3.955 $Y=0.35
+ $X2=0 $Y2=0
cc_408 N_A_437_144#_c_480_n N_A_547_167#_c_1239_n 0.00577175f $X=2.51 $Y=0.875
+ $X2=0 $Y2=0
cc_409 N_A_437_144#_c_470_n N_A_547_167#_c_1240_n 2.29952e-19 $X=4.045 $Y=0.875
+ $X2=0 $Y2=0
cc_410 N_A_437_144#_c_474_n N_A_547_167#_c_1240_n 2.46049e-19 $X=4.6 $Y=0.875
+ $X2=0 $Y2=0
cc_411 N_A_437_144#_c_475_n N_A_547_167#_c_1240_n 0.00411914f $X=4.6 $Y=0.95
+ $X2=0 $Y2=0
cc_412 N_A_437_144#_c_478_n N_A_547_167#_c_1240_n 0.00352722f $X=3.955 $Y=0.35
+ $X2=0 $Y2=0
cc_413 N_A_437_144#_c_479_n N_A_547_167#_c_1240_n 0.00420402f $X=3.955 $Y=0.35
+ $X2=0 $Y2=0
cc_414 N_A_437_144#_c_471_n N_A_716_167#_c_1271_n 0.00547283f $X=4.275 $Y=0.95
+ $X2=0 $Y2=0
cc_415 N_A_437_144#_c_472_n N_A_716_167#_c_1271_n 0.00619596f $X=4.12 $Y=0.95
+ $X2=0 $Y2=0
cc_416 N_A_437_144#_M1015_g N_A_716_167#_c_1271_n 0.014695f $X=4.35 $Y=2.205
+ $X2=0 $Y2=0
cc_417 N_A_437_144#_c_475_n N_A_716_167#_c_1271_n 0.0178292f $X=4.6 $Y=0.95
+ $X2=0 $Y2=0
cc_418 N_A_955_271#_M1004_g N_A_630_167#_c_740_n 0.00480446f $X=4.875 $Y=2.095
+ $X2=0 $Y2=0
cc_419 N_A_955_271#_c_587_n N_A_630_167#_c_741_n 0.00627282f $X=5.58 $Y=1.93
+ $X2=0 $Y2=0
cc_420 N_A_955_271#_c_588_n N_A_630_167#_c_741_n 0.00839601f $X=5.735 $Y=2.015
+ $X2=0 $Y2=0
cc_421 N_A_955_271#_c_587_n N_A_630_167#_c_733_n 0.00455615f $X=5.58 $Y=1.93
+ $X2=0 $Y2=0
cc_422 N_A_955_271#_c_598_p N_A_630_167#_c_733_n 0.00130209f $X=6.06 $Y=2.015
+ $X2=0 $Y2=0
cc_423 N_A_955_271#_c_579_n N_A_630_167#_c_733_n 0.0095756f $X=5.58 $Y=1.52
+ $X2=0 $Y2=0
cc_424 N_A_955_271#_c_580_n N_A_630_167#_c_733_n 0.00428463f $X=5.735 $Y=0.915
+ $X2=0 $Y2=0
cc_425 N_A_955_271#_M1004_g N_A_630_167#_c_734_n 0.0149874f $X=4.875 $Y=2.095
+ $X2=0 $Y2=0
cc_426 N_A_955_271#_c_567_n N_A_630_167#_c_734_n 0.00720111f $X=5.425 $Y=1.52
+ $X2=0 $Y2=0
cc_427 N_A_955_271#_c_568_n N_A_630_167#_c_734_n 0.00608898f $X=4.94 $Y=1.52
+ $X2=0 $Y2=0
cc_428 N_A_955_271#_c_587_n N_A_630_167#_c_734_n 9.07068e-19 $X=5.58 $Y=1.93
+ $X2=0 $Y2=0
cc_429 N_A_955_271#_c_579_n N_A_630_167#_c_734_n 0.00203851f $X=5.58 $Y=1.52
+ $X2=0 $Y2=0
cc_430 N_A_955_271#_c_587_n N_A_630_167#_c_744_n 0.00456773f $X=5.58 $Y=1.93
+ $X2=0 $Y2=0
cc_431 N_A_955_271#_c_598_p N_A_630_167#_c_744_n 0.0138274f $X=6.06 $Y=2.015
+ $X2=0 $Y2=0
cc_432 N_A_955_271#_c_569_n N_A_630_167#_M1008_g 0.0120473f $X=5.765 $Y=0.39
+ $X2=0 $Y2=0
cc_433 N_A_955_271#_c_570_n N_A_630_167#_M1008_g 0.00599024f $X=5.637 $Y=1.355
+ $X2=0 $Y2=0
cc_434 N_A_955_271#_c_610_p N_A_630_167#_M1008_g 0.00812227f $X=6.82 $Y=0.915
+ $X2=0 $Y2=0
cc_435 N_A_955_271#_c_579_n N_A_630_167#_M1008_g 0.00175768f $X=5.58 $Y=1.52
+ $X2=0 $Y2=0
cc_436 N_A_955_271#_c_580_n N_A_630_167#_M1008_g 7.32094e-19 $X=5.735 $Y=0.915
+ $X2=0 $Y2=0
cc_437 N_A_955_271#_c_564_n N_RESET_B_M1010_g 0.00717333f $X=7.105 $Y=1.185
+ $X2=0 $Y2=0
cc_438 N_A_955_271#_c_569_n N_RESET_B_M1010_g 0.0019482f $X=5.765 $Y=0.39 $X2=0
+ $Y2=0
cc_439 N_A_955_271#_c_610_p N_RESET_B_M1010_g 0.0125465f $X=6.82 $Y=0.915 $X2=0
+ $Y2=0
cc_440 N_A_955_271#_c_571_n N_RESET_B_M1010_g 0.00332434f $X=6.985 $Y=1.35 $X2=0
+ $Y2=0
cc_441 N_A_955_271#_c_572_n N_RESET_B_M1010_g 6.2477e-19 $X=6.985 $Y=1.35 $X2=0
+ $Y2=0
cc_442 N_A_955_271#_c_573_n N_RESET_B_M1010_g 0.00248953f $X=6.99 $Y=0.83 $X2=0
+ $Y2=0
cc_443 N_A_955_271#_c_575_n N_RESET_B_M1010_g 5.20073e-19 $X=7.08 $Y=0.34 $X2=0
+ $Y2=0
cc_444 N_A_955_271#_M1020_g N_RESET_B_M1003_g 0.0187196f $X=6.895 $Y=2.155 $X2=0
+ $Y2=0
cc_445 N_A_955_271#_c_587_n RESET_B 0.00593875f $X=5.58 $Y=1.93 $X2=0 $Y2=0
cc_446 N_A_955_271#_c_570_n RESET_B 0.0148125f $X=5.637 $Y=1.355 $X2=0 $Y2=0
cc_447 N_A_955_271#_c_598_p RESET_B 0.0102503f $X=6.06 $Y=2.015 $X2=0 $Y2=0
cc_448 N_A_955_271#_c_610_p RESET_B 0.0507408f $X=6.82 $Y=0.915 $X2=0 $Y2=0
cc_449 N_A_955_271#_c_625_p RESET_B 0.0177203f $X=6.172 $Y=2.1 $X2=0 $Y2=0
cc_450 N_A_955_271#_c_571_n RESET_B 0.0286013f $X=6.985 $Y=1.35 $X2=0 $Y2=0
cc_451 N_A_955_271#_c_572_n RESET_B 0.00907317f $X=6.985 $Y=1.35 $X2=0 $Y2=0
cc_452 N_A_955_271#_c_579_n RESET_B 0.0288833f $X=5.58 $Y=1.52 $X2=0 $Y2=0
cc_453 N_A_955_271#_c_580_n RESET_B 0.00204104f $X=5.735 $Y=0.915 $X2=0 $Y2=0
cc_454 N_A_955_271#_c_610_p N_RESET_B_c_847_n 0.00101866f $X=6.82 $Y=0.915 $X2=0
+ $Y2=0
cc_455 N_A_955_271#_c_571_n N_RESET_B_c_847_n 3.44632e-19 $X=6.985 $Y=1.35 $X2=0
+ $Y2=0
cc_456 N_A_955_271#_c_572_n N_RESET_B_c_847_n 0.0188319f $X=6.985 $Y=1.35 $X2=0
+ $Y2=0
cc_457 N_A_955_271#_M1020_g N_A_1394_367#_c_886_n 0.0134608f $X=6.895 $Y=2.155
+ $X2=0 $Y2=0
cc_458 N_A_955_271#_c_566_n N_A_1394_367#_M1002_g 0.0124449f $X=8.905 $Y=1.26
+ $X2=0 $Y2=0
cc_459 N_A_955_271#_c_574_n N_A_1394_367#_M1002_g 0.0144315f $X=8.265 $Y=0.34
+ $X2=0 $Y2=0
cc_460 N_A_955_271#_c_576_n N_A_1394_367#_M1002_g 0.0242002f $X=8.35 $Y=1.26
+ $X2=0 $Y2=0
cc_461 N_A_955_271#_c_577_n N_A_1394_367#_M1002_g 0.00725746f $X=8.435 $Y=1.425
+ $X2=0 $Y2=0
cc_462 N_A_955_271#_c_581_n N_A_1394_367#_M1002_g 0.0204045f $X=8.905 $Y=1.425
+ $X2=0 $Y2=0
cc_463 N_A_955_271#_M1014_g N_A_1394_367#_c_888_n 0.0204045f $X=8.655 $Y=2.465
+ $X2=0 $Y2=0
cc_464 N_A_955_271#_c_577_n N_A_1394_367#_c_888_n 0.0017562f $X=8.435 $Y=1.425
+ $X2=0 $Y2=0
cc_465 N_A_955_271#_M1020_g N_A_1394_367#_c_889_n 0.00300056f $X=6.895 $Y=2.155
+ $X2=0 $Y2=0
cc_466 N_A_955_271#_c_564_n N_A_1394_367#_c_889_n 0.00651829f $X=7.105 $Y=1.185
+ $X2=0 $Y2=0
cc_467 N_A_955_271#_c_571_n N_A_1394_367#_c_889_n 0.023142f $X=6.985 $Y=1.35
+ $X2=0 $Y2=0
cc_468 N_A_955_271#_c_572_n N_A_1394_367#_c_889_n 0.00402314f $X=6.985 $Y=1.35
+ $X2=0 $Y2=0
cc_469 N_A_955_271#_M1020_g N_A_1394_367#_c_896_n 8.53352e-19 $X=6.895 $Y=2.155
+ $X2=0 $Y2=0
cc_470 N_A_955_271#_c_571_n N_A_1394_367#_c_896_n 0.00574113f $X=6.985 $Y=1.35
+ $X2=0 $Y2=0
cc_471 N_A_955_271#_c_572_n N_A_1394_367#_c_896_n 0.00471987f $X=6.985 $Y=1.35
+ $X2=0 $Y2=0
cc_472 N_A_955_271#_c_564_n N_A_1394_367#_c_890_n 0.00726555f $X=7.105 $Y=1.185
+ $X2=0 $Y2=0
cc_473 N_A_955_271#_c_571_n N_A_1394_367#_c_890_n 0.0026176f $X=6.985 $Y=1.35
+ $X2=0 $Y2=0
cc_474 N_A_955_271#_c_573_n N_A_1394_367#_c_890_n 0.00939723f $X=6.99 $Y=0.83
+ $X2=0 $Y2=0
cc_475 N_A_955_271#_c_574_n N_A_1394_367#_c_890_n 0.0202398f $X=8.265 $Y=0.34
+ $X2=0 $Y2=0
cc_476 N_A_955_271#_c_652_p N_A_1394_367#_c_890_n 0.0143173f $X=6.95 $Y=0.915
+ $X2=0 $Y2=0
cc_477 N_A_955_271#_c_587_n N_VPWR_M1012_s 0.00114434f $X=5.58 $Y=1.93 $X2=0
+ $Y2=0
cc_478 N_A_955_271#_c_598_p N_VPWR_M1012_s 0.00248817f $X=6.06 $Y=2.015 $X2=0
+ $Y2=0
cc_479 N_A_955_271#_c_588_n N_VPWR_M1012_s 0.00157697f $X=5.735 $Y=2.015 $X2=0
+ $Y2=0
cc_480 N_A_955_271#_M1004_g N_VPWR_c_937_n 0.00543343f $X=4.875 $Y=2.095 $X2=0
+ $Y2=0
cc_481 N_A_955_271#_c_598_p N_VPWR_c_938_n 0.00768878f $X=6.06 $Y=2.015 $X2=0
+ $Y2=0
cc_482 N_A_955_271#_c_588_n N_VPWR_c_938_n 0.015781f $X=5.735 $Y=2.015 $X2=0
+ $Y2=0
cc_483 N_A_955_271#_c_659_p N_VPWR_c_939_n 0.0136943f $X=6.155 $Y=2.91 $X2=0
+ $Y2=0
cc_484 N_A_955_271#_M1020_g N_VPWR_c_940_n 0.00533578f $X=6.895 $Y=2.155 $X2=0
+ $Y2=0
cc_485 N_A_955_271#_M1014_g N_VPWR_c_941_n 0.00394937f $X=8.655 $Y=2.465 $X2=0
+ $Y2=0
cc_486 N_A_955_271#_c_577_n N_VPWR_c_941_n 0.0113208f $X=8.435 $Y=1.425 $X2=0
+ $Y2=0
cc_487 N_A_955_271#_c_578_n N_VPWR_c_941_n 0.00788372f $X=8.745 $Y=1.425 $X2=0
+ $Y2=0
cc_488 N_A_955_271#_M1020_g N_VPWR_c_947_n 0.00312414f $X=6.895 $Y=2.155 $X2=0
+ $Y2=0
cc_489 N_A_955_271#_M1014_g N_VPWR_c_948_n 0.00585385f $X=8.655 $Y=2.465 $X2=0
+ $Y2=0
cc_490 N_A_955_271#_M1012_d N_VPWR_c_932_n 0.0041489f $X=6.015 $Y=1.835 $X2=0
+ $Y2=0
cc_491 N_A_955_271#_M1020_g N_VPWR_c_932_n 0.00410284f $X=6.895 $Y=2.155 $X2=0
+ $Y2=0
cc_492 N_A_955_271#_M1014_g N_VPWR_c_932_n 0.0119158f $X=8.655 $Y=2.465 $X2=0
+ $Y2=0
cc_493 N_A_955_271#_c_659_p N_VPWR_c_932_n 0.00866972f $X=6.155 $Y=2.91 $X2=0
+ $Y2=0
cc_494 N_A_955_271#_M1004_g N_A_625_377#_c_1051_n 0.0117873f $X=4.875 $Y=2.095
+ $X2=0 $Y2=0
cc_495 N_A_955_271#_c_567_n N_A_625_377#_c_1051_n 0.0108055f $X=5.425 $Y=1.52
+ $X2=0 $Y2=0
cc_496 N_A_955_271#_c_568_n N_A_625_377#_c_1051_n 5.60514e-19 $X=4.94 $Y=1.52
+ $X2=0 $Y2=0
cc_497 N_A_955_271#_M1004_g N_A_625_377#_c_1053_n 0.00636232f $X=4.875 $Y=2.095
+ $X2=0 $Y2=0
cc_498 N_A_955_271#_c_567_n N_A_625_377#_c_1053_n 0.0270287f $X=5.425 $Y=1.52
+ $X2=0 $Y2=0
cc_499 N_A_955_271#_c_568_n N_A_625_377#_c_1053_n 0.00414436f $X=4.94 $Y=1.52
+ $X2=0 $Y2=0
cc_500 N_A_955_271#_c_587_n N_A_625_377#_c_1053_n 0.00587084f $X=5.58 $Y=1.93
+ $X2=0 $Y2=0
cc_501 N_A_955_271#_c_588_n N_A_625_377#_c_1053_n 0.0142642f $X=5.735 $Y=2.015
+ $X2=0 $Y2=0
cc_502 N_A_955_271#_c_574_n N_Q_N_M1002_s 0.00274742f $X=8.265 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_503 N_A_955_271#_c_564_n N_Q_N_c_1084_n 0.00308197f $X=7.105 $Y=1.185 $X2=0
+ $Y2=0
cc_504 N_A_955_271#_c_574_n N_Q_N_c_1084_n 0.0197029f $X=8.265 $Y=0.34 $X2=0
+ $Y2=0
cc_505 N_A_955_271#_c_576_n N_Q_N_c_1084_n 0.0268773f $X=8.35 $Y=1.26 $X2=0
+ $Y2=0
cc_506 N_A_955_271#_c_577_n N_Q_N_c_1084_n 0.026906f $X=8.435 $Y=1.425 $X2=0
+ $Y2=0
cc_507 N_A_955_271#_c_581_n N_Q_N_c_1084_n 5.80764e-19 $X=8.905 $Y=1.425 $X2=0
+ $Y2=0
cc_508 N_A_955_271#_M1014_g Q 0.00734739f $X=8.655 $Y=2.465 $X2=0 $Y2=0
cc_509 N_A_955_271#_c_566_n Q 0.0121166f $X=8.905 $Y=1.26 $X2=0 $Y2=0
cc_510 N_A_955_271#_c_576_n Q 0.00386273f $X=8.35 $Y=1.26 $X2=0 $Y2=0
cc_511 N_A_955_271#_c_578_n Q 0.0280336f $X=8.745 $Y=1.425 $X2=0 $Y2=0
cc_512 N_A_955_271#_c_566_n N_Q_c_1106_n 0.00302508f $X=8.905 $Y=1.26 $X2=0
+ $Y2=0
cc_513 N_A_955_271#_M1014_g N_Q_c_1110_n 0.00342589f $X=8.655 $Y=2.465 $X2=0
+ $Y2=0
cc_514 N_A_955_271#_c_578_n N_Q_c_1110_n 0.00813773f $X=8.745 $Y=1.425 $X2=0
+ $Y2=0
cc_515 N_A_955_271#_c_581_n N_Q_c_1110_n 0.00722975f $X=8.905 $Y=1.425 $X2=0
+ $Y2=0
cc_516 N_A_955_271#_c_610_p N_VGND_M1010_d 0.0147429f $X=6.82 $Y=0.915 $X2=0
+ $Y2=0
cc_517 N_A_955_271#_c_571_n N_VGND_M1010_d 0.00110183f $X=6.985 $Y=1.35 $X2=0
+ $Y2=0
cc_518 N_A_955_271#_c_573_n N_VGND_M1010_d 0.00263528f $X=6.99 $Y=0.83 $X2=0
+ $Y2=0
cc_519 N_A_955_271#_c_652_p N_VGND_M1010_d 0.00214409f $X=6.95 $Y=0.915 $X2=0
+ $Y2=0
cc_520 N_A_955_271#_c_574_n N_VGND_M1002_d 0.00109296f $X=8.265 $Y=0.34 $X2=0
+ $Y2=0
cc_521 N_A_955_271#_c_576_n N_VGND_M1002_d 0.00699673f $X=8.35 $Y=1.26 $X2=0
+ $Y2=0
cc_522 N_A_955_271#_M1021_g N_VGND_c_1129_n 0.00220654f $X=5.03 $Y=0.555 $X2=0
+ $Y2=0
cc_523 N_A_955_271#_c_569_n N_VGND_c_1129_n 0.00373821f $X=5.765 $Y=0.39 $X2=0
+ $Y2=0
cc_524 N_A_955_271#_c_564_n N_VGND_c_1130_n 4.3603e-19 $X=7.105 $Y=1.185 $X2=0
+ $Y2=0
cc_525 N_A_955_271#_c_569_n N_VGND_c_1130_n 0.0137257f $X=5.765 $Y=0.39 $X2=0
+ $Y2=0
cc_526 N_A_955_271#_c_610_p N_VGND_c_1130_n 0.0213827f $X=6.82 $Y=0.915 $X2=0
+ $Y2=0
cc_527 N_A_955_271#_c_573_n N_VGND_c_1130_n 0.0179184f $X=6.99 $Y=0.83 $X2=0
+ $Y2=0
cc_528 N_A_955_271#_c_575_n N_VGND_c_1130_n 0.0144409f $X=7.08 $Y=0.34 $X2=0
+ $Y2=0
cc_529 N_A_955_271#_c_566_n N_VGND_c_1131_n 0.0139907f $X=8.905 $Y=1.26 $X2=0
+ $Y2=0
cc_530 N_A_955_271#_c_574_n N_VGND_c_1131_n 0.0143144f $X=8.265 $Y=0.34 $X2=0
+ $Y2=0
cc_531 N_A_955_271#_c_576_n N_VGND_c_1131_n 0.0494649f $X=8.35 $Y=1.26 $X2=0
+ $Y2=0
cc_532 N_A_955_271#_c_578_n N_VGND_c_1131_n 0.0166162f $X=8.745 $Y=1.425 $X2=0
+ $Y2=0
cc_533 N_A_955_271#_c_581_n N_VGND_c_1131_n 0.00553362f $X=8.905 $Y=1.425 $X2=0
+ $Y2=0
cc_534 N_A_955_271#_c_564_n N_VGND_c_1136_n 2.69083e-19 $X=7.105 $Y=1.185 $X2=0
+ $Y2=0
cc_535 N_A_955_271#_c_574_n N_VGND_c_1136_n 0.0880093f $X=8.265 $Y=0.34 $X2=0
+ $Y2=0
cc_536 N_A_955_271#_c_575_n N_VGND_c_1136_n 0.0129036f $X=7.08 $Y=0.34 $X2=0
+ $Y2=0
cc_537 N_A_955_271#_M1021_g N_VGND_c_1138_n 0.00482246f $X=5.03 $Y=0.555 $X2=0
+ $Y2=0
cc_538 N_A_955_271#_c_569_n N_VGND_c_1138_n 0.0253479f $X=5.765 $Y=0.39 $X2=0
+ $Y2=0
cc_539 N_A_955_271#_c_566_n N_VGND_c_1139_n 0.00477169f $X=8.905 $Y=1.26 $X2=0
+ $Y2=0
cc_540 N_A_955_271#_M1008_s N_VGND_c_1140_n 0.00215158f $X=5.64 $Y=0.235 $X2=0
+ $Y2=0
cc_541 N_A_955_271#_M1021_g N_VGND_c_1140_n 0.00976497f $X=5.03 $Y=0.555 $X2=0
+ $Y2=0
cc_542 N_A_955_271#_c_566_n N_VGND_c_1140_n 0.00944487f $X=8.905 $Y=1.26 $X2=0
+ $Y2=0
cc_543 N_A_955_271#_c_569_n N_VGND_c_1140_n 0.0149015f $X=5.765 $Y=0.39 $X2=0
+ $Y2=0
cc_544 N_A_955_271#_c_610_p N_VGND_c_1140_n 0.0188204f $X=6.82 $Y=0.915 $X2=0
+ $Y2=0
cc_545 N_A_955_271#_c_574_n N_VGND_c_1140_n 0.0504717f $X=8.265 $Y=0.34 $X2=0
+ $Y2=0
cc_546 N_A_955_271#_c_575_n N_VGND_c_1140_n 0.00699798f $X=7.08 $Y=0.34 $X2=0
+ $Y2=0
cc_547 N_A_955_271#_c_652_p N_VGND_c_1140_n 0.00318449f $X=6.95 $Y=0.915 $X2=0
+ $Y2=0
cc_548 N_A_955_271#_M1021_g N_A_716_167#_c_1271_n 0.0203186f $X=5.03 $Y=0.555
+ $X2=0 $Y2=0
cc_549 N_A_955_271#_c_567_n N_A_716_167#_c_1271_n 0.0459515f $X=5.425 $Y=1.52
+ $X2=0 $Y2=0
cc_550 N_A_955_271#_c_568_n N_A_716_167#_c_1271_n 0.00462387f $X=4.94 $Y=1.52
+ $X2=0 $Y2=0
cc_551 N_A_955_271#_c_570_n N_A_716_167#_c_1271_n 0.0148811f $X=5.637 $Y=1.355
+ $X2=0 $Y2=0
cc_552 N_A_955_271#_c_580_n N_A_716_167#_c_1271_n 0.00515325f $X=5.735 $Y=0.915
+ $X2=0 $Y2=0
cc_553 N_A_955_271#_M1021_g N_A_716_167#_c_1272_n 0.00754356f $X=5.03 $Y=0.555
+ $X2=0 $Y2=0
cc_554 N_A_955_271#_c_569_n N_A_716_167#_c_1272_n 0.0355566f $X=5.765 $Y=0.39
+ $X2=0 $Y2=0
cc_555 N_A_955_271#_c_580_n N_A_716_167#_c_1272_n 0.00987742f $X=5.735 $Y=0.915
+ $X2=0 $Y2=0
cc_556 N_A_955_271#_c_610_p A_1211_47# 0.00293659f $X=6.82 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_557 N_A_630_167#_M1008_g N_RESET_B_M1010_g 0.0891896f $X=5.98 $Y=0.655 $X2=0
+ $Y2=0
cc_558 N_A_630_167#_c_744_n N_RESET_B_M1003_g 0.0158965f $X=5.94 $Y=1.725 $X2=0
+ $Y2=0
cc_559 N_A_630_167#_M1008_g N_RESET_B_M1003_g 0.0101049f $X=5.98 $Y=0.655 $X2=0
+ $Y2=0
cc_560 N_A_630_167#_c_744_n RESET_B 0.00250228f $X=5.94 $Y=1.725 $X2=0 $Y2=0
cc_561 N_A_630_167#_M1008_g RESET_B 0.0115099f $X=5.98 $Y=0.655 $X2=0 $Y2=0
cc_562 N_A_630_167#_c_736_n RESET_B 0.00642303f $X=5.96 $Y=1.65 $X2=0 $Y2=0
cc_563 N_A_630_167#_c_740_n N_VPWR_c_937_n 0.0322782f $X=5.345 $Y=3.03 $X2=0
+ $Y2=0
cc_564 N_A_630_167#_c_741_n N_VPWR_c_937_n 0.0125149f $X=5.42 $Y=2.955 $X2=0
+ $Y2=0
cc_565 N_A_630_167#_c_753_n N_VPWR_c_937_n 0.0180825f $X=3.51 $Y=2.452 $X2=0
+ $Y2=0
cc_566 N_A_630_167#_c_741_n N_VPWR_c_938_n 0.0234873f $X=5.42 $Y=2.955 $X2=0
+ $Y2=0
cc_567 N_A_630_167#_c_733_n N_VPWR_c_938_n 6.22796e-19 $X=5.865 $Y=1.65 $X2=0
+ $Y2=0
cc_568 N_A_630_167#_c_744_n N_VPWR_c_938_n 0.0158362f $X=5.94 $Y=1.725 $X2=0
+ $Y2=0
cc_569 N_A_630_167#_c_744_n N_VPWR_c_939_n 0.00486043f $X=5.94 $Y=1.725 $X2=0
+ $Y2=0
cc_570 N_A_630_167#_c_750_n N_VPWR_c_942_n 0.00869323f $X=2.965 $Y=2.57 $X2=0
+ $Y2=0
cc_571 N_A_630_167#_c_740_n N_VPWR_c_943_n 0.0222812f $X=5.345 $Y=3.03 $X2=0
+ $Y2=0
cc_572 N_A_630_167#_c_749_n N_VPWR_c_946_n 0.00739538f $X=3.345 $Y=2.57 $X2=0
+ $Y2=0
cc_573 N_A_630_167#_c_750_n N_VPWR_c_946_n 0.00340038f $X=2.965 $Y=2.57 $X2=0
+ $Y2=0
cc_574 N_A_630_167#_c_751_n N_VPWR_c_946_n 0.0222914f $X=3.51 $Y=2.94 $X2=0
+ $Y2=0
cc_575 N_A_630_167#_c_752_n N_VPWR_c_946_n 0.0240237f $X=3.51 $Y=2.94 $X2=0
+ $Y2=0
cc_576 N_A_630_167#_c_753_n N_VPWR_c_946_n 0.00534322f $X=3.51 $Y=2.452 $X2=0
+ $Y2=0
cc_577 N_A_630_167#_c_740_n N_VPWR_c_932_n 0.0688333f $X=5.345 $Y=3.03 $X2=0
+ $Y2=0
cc_578 N_A_630_167#_c_744_n N_VPWR_c_932_n 0.0082726f $X=5.94 $Y=1.725 $X2=0
+ $Y2=0
cc_579 N_A_630_167#_c_749_n N_VPWR_c_932_n 0.0111918f $X=3.345 $Y=2.57 $X2=0
+ $Y2=0
cc_580 N_A_630_167#_c_750_n N_VPWR_c_932_n 0.00488203f $X=2.965 $Y=2.57 $X2=0
+ $Y2=0
cc_581 N_A_630_167#_c_751_n N_VPWR_c_932_n 0.0112369f $X=3.51 $Y=2.94 $X2=0
+ $Y2=0
cc_582 N_A_630_167#_c_752_n N_VPWR_c_932_n 0.00763827f $X=3.51 $Y=2.94 $X2=0
+ $Y2=0
cc_583 N_A_630_167#_c_753_n N_VPWR_c_932_n 0.00693204f $X=3.51 $Y=2.452 $X2=0
+ $Y2=0
cc_584 N_A_630_167#_M1000_d N_A_625_377#_c_1051_n 0.00296136f $X=3.54 $Y=1.885
+ $X2=0 $Y2=0
cc_585 N_A_630_167#_c_737_n N_A_625_377#_c_1051_n 0.00253381f $X=3.16 $Y=1.6
+ $X2=0 $Y2=0
cc_586 N_A_630_167#_c_753_n N_A_625_377#_c_1051_n 0.0299989f $X=3.51 $Y=2.452
+ $X2=0 $Y2=0
cc_587 N_A_630_167#_c_746_n N_A_625_377#_c_1052_n 0.0305776f $X=2.88 $Y=2.43
+ $X2=0 $Y2=0
cc_588 N_A_630_167#_c_737_n N_A_625_377#_c_1052_n 0.0193484f $X=3.16 $Y=1.6
+ $X2=0 $Y2=0
cc_589 N_A_630_167#_c_749_n N_A_625_377#_c_1052_n 0.0158341f $X=3.345 $Y=2.57
+ $X2=0 $Y2=0
cc_590 N_A_630_167#_c_740_n N_A_625_377#_c_1053_n 0.00614689f $X=5.345 $Y=3.03
+ $X2=0 $Y2=0
cc_591 N_A_630_167#_c_741_n N_A_625_377#_c_1053_n 0.00639547f $X=5.42 $Y=2.955
+ $X2=0 $Y2=0
cc_592 N_A_630_167#_M1008_g N_VGND_c_1130_n 0.00233418f $X=5.98 $Y=0.655 $X2=0
+ $Y2=0
cc_593 N_A_630_167#_M1008_g N_VGND_c_1138_n 0.0054895f $X=5.98 $Y=0.655 $X2=0
+ $Y2=0
cc_594 N_A_630_167#_M1008_g N_VGND_c_1140_n 0.0073794f $X=5.98 $Y=0.655 $X2=0
+ $Y2=0
cc_595 N_A_630_167#_c_738_n N_A_547_167#_c_1237_n 0.00954069f $X=2.965 $Y=1.6
+ $X2=0 $Y2=0
cc_596 N_A_630_167#_c_739_n N_A_547_167#_c_1238_n 0.0158815f $X=3.29 $Y=1.11
+ $X2=0 $Y2=0
cc_597 N_A_630_167#_M1008_g N_A_716_167#_c_1272_n 9.18385e-19 $X=5.98 $Y=0.655
+ $X2=0 $Y2=0
cc_598 N_RESET_B_M1003_g N_VPWR_c_938_n 6.91881e-19 $X=6.37 $Y=2.465 $X2=0 $Y2=0
cc_599 N_RESET_B_M1003_g N_VPWR_c_939_n 0.00585385f $X=6.37 $Y=2.465 $X2=0 $Y2=0
cc_600 N_RESET_B_M1003_g N_VPWR_c_940_n 0.00699015f $X=6.37 $Y=2.465 $X2=0 $Y2=0
cc_601 RESET_B N_VPWR_c_940_n 0.0154975f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_602 N_RESET_B_c_847_n N_VPWR_c_940_n 5.76405e-19 $X=6.43 $Y=1.375 $X2=0 $Y2=0
cc_603 N_RESET_B_M1003_g N_VPWR_c_932_n 0.0118474f $X=6.37 $Y=2.465 $X2=0 $Y2=0
cc_604 N_RESET_B_M1010_g N_VGND_c_1130_n 0.0152611f $X=6.34 $Y=0.655 $X2=0 $Y2=0
cc_605 N_RESET_B_M1010_g N_VGND_c_1138_n 0.00486043f $X=6.34 $Y=0.655 $X2=0
+ $Y2=0
cc_606 N_RESET_B_M1010_g N_VGND_c_1140_n 0.00443044f $X=6.34 $Y=0.655 $X2=0
+ $Y2=0
cc_607 N_A_1394_367#_c_896_n N_VPWR_c_940_n 7.11296e-19 $X=7.53 $Y=2.15 $X2=0
+ $Y2=0
cc_608 N_A_1394_367#_c_893_n N_VPWR_c_941_n 0.0194399f $X=8.225 $Y=1.725 $X2=0
+ $Y2=0
cc_609 N_A_1394_367#_c_893_n N_VPWR_c_947_n 0.00525069f $X=8.225 $Y=1.725 $X2=0
+ $Y2=0
cc_610 N_A_1394_367#_c_893_n N_VPWR_c_932_n 0.0101648f $X=8.225 $Y=1.725 $X2=0
+ $Y2=0
cc_611 N_A_1394_367#_c_896_n N_VPWR_c_932_n 0.0268204f $X=7.53 $Y=2.15 $X2=0
+ $Y2=0
cc_612 N_A_1394_367#_c_885_n N_Q_N_c_1084_n 0.0198922f $X=8.15 $Y=1.65 $X2=0
+ $Y2=0
cc_613 N_A_1394_367#_M1002_g N_Q_N_c_1084_n 0.013151f $X=8.225 $Y=0.73 $X2=0
+ $Y2=0
cc_614 N_A_1394_367#_c_893_n N_Q_N_c_1084_n 0.00267058f $X=8.225 $Y=1.725 $X2=0
+ $Y2=0
cc_615 N_A_1394_367#_c_889_n N_Q_N_c_1084_n 0.0612306f $X=7.56 $Y=1.74 $X2=0
+ $Y2=0
cc_616 N_A_1394_367#_c_895_n N_Q_N_c_1084_n 0.0047936f $X=7.56 $Y=1.74 $X2=0
+ $Y2=0
cc_617 N_A_1394_367#_c_896_n N_Q_N_c_1084_n 0.0563892f $X=7.53 $Y=2.15 $X2=0
+ $Y2=0
cc_618 N_A_1394_367#_c_890_n N_Q_N_c_1084_n 0.027434f $X=7.53 $Y=0.87 $X2=0
+ $Y2=0
cc_619 N_A_1394_367#_M1002_g N_VGND_c_1131_n 0.00355002f $X=8.225 $Y=0.73 $X2=0
+ $Y2=0
cc_620 N_A_1394_367#_M1002_g N_VGND_c_1136_n 0.00311022f $X=8.225 $Y=0.73 $X2=0
+ $Y2=0
cc_621 N_A_1394_367#_M1002_g N_VGND_c_1140_n 0.00549582f $X=8.225 $Y=0.73 $X2=0
+ $Y2=0
cc_622 N_VPWR_M1015_d N_A_625_377#_c_1051_n 0.00327524f $X=4.425 $Y=1.885 $X2=0
+ $Y2=0
cc_623 N_VPWR_c_937_n N_A_625_377#_c_1051_n 0.0218816f $X=4.565 $Y=2.31 $X2=0
+ $Y2=0
cc_624 N_VPWR_c_937_n N_A_625_377#_c_1053_n 0.00453955f $X=4.565 $Y=2.31 $X2=0
+ $Y2=0
cc_625 N_VPWR_c_932_n N_Q_N_M1022_s 0.00336915f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_626 N_VPWR_c_941_n N_Q_N_c_1084_n 0.00186321f $X=8.44 $Y=1.98 $X2=0 $Y2=0
cc_627 N_VPWR_c_947_n N_Q_N_c_1087_n 0.0188828f $X=8.285 $Y=3.33 $X2=0 $Y2=0
cc_628 N_VPWR_c_932_n N_Q_N_c_1087_n 0.0107922f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_629 N_VPWR_c_932_n N_Q_M1014_d 0.00336915f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_630 N_VPWR_c_948_n Q 0.0525755f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_631 N_VPWR_c_932_n Q 0.0290805f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_632 N_VPWR_c_941_n N_Q_c_1110_n 0.00137233f $X=8.44 $Y=1.98 $X2=0 $Y2=0
cc_633 N_A_625_377#_c_1051_n A_813_377# 0.00366293f $X=4.925 $Y=1.94 $X2=-0.19
+ $Y2=1.655
cc_634 N_Q_c_1106_n N_VGND_c_1131_n 0.0293387f $X=9.12 $Y=0.455 $X2=0 $Y2=0
cc_635 N_Q_c_1106_n N_VGND_c_1139_n 0.0295076f $X=9.12 $Y=0.455 $X2=0 $Y2=0
cc_636 N_Q_c_1106_n N_VGND_c_1140_n 0.0192182f $X=9.12 $Y=0.455 $X2=0 $Y2=0
cc_637 N_VGND_c_1134_n N_A_547_167#_c_1238_n 0.00328473f $X=4.685 $Y=0 $X2=0
+ $Y2=0
cc_638 N_VGND_c_1140_n N_A_547_167#_c_1238_n 0.00719115f $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_639 N_VGND_c_1134_n N_A_547_167#_c_1240_n 0.00726672f $X=4.685 $Y=0 $X2=0
+ $Y2=0
cc_640 N_VGND_c_1140_n N_A_547_167#_c_1240_n 0.00787534f $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_641 N_VGND_c_1129_n N_A_716_167#_c_1271_n 0.013624f $X=4.815 $Y=0.555 $X2=0
+ $Y2=0
cc_642 N_VGND_c_1138_n N_A_716_167#_c_1272_n 0.00813734f $X=6.39 $Y=0 $X2=0
+ $Y2=0
cc_643 N_VGND_c_1140_n N_A_716_167#_c_1272_n 0.00821462f $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_644 N_VGND_c_1140_n A_1211_47# 0.00305025f $X=9.36 $Y=0 $X2=-0.19 $Y2=-0.245
cc_645 N_A_547_167#_c_1238_n N_A_716_167#_c_1271_n 0.051986f $X=4.29 $Y=0.69
+ $X2=0 $Y2=0
cc_646 N_A_547_167#_c_1240_n N_A_716_167#_c_1271_n 0.0175016f $X=4.385 $Y=0.555
+ $X2=0 $Y2=0
cc_647 N_A_547_167#_c_1240_n N_A_716_167#_c_1272_n 2.80781e-19 $X=4.385 $Y=0.555
+ $X2=0 $Y2=0
