* File: sky130_fd_sc_lp__o32ai_4.pex.spice
* Created: Wed Sep  2 10:26:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32AI_4%B2 3 7 11 15 19 23 27 31 33 34 35 36 55 56
c86 55 0 9.07802e-20 $X=1.69 $Y=1.46
r87 54 56 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.69 $Y=1.46 $X2=1.78
+ $Y2=1.46
r88 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.46 $X2=1.69 $Y2=1.46
r89 51 54 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.35 $Y=1.46
+ $X2=1.69 $Y2=1.46
r90 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=1.46 $X2=1.35 $Y2=1.46
r91 49 51 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.92 $Y=1.46
+ $X2=1.35 $Y2=1.46
r92 47 49 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.67 $Y=1.46
+ $X2=0.92 $Y2=1.46
r93 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.46 $X2=0.67 $Y2=1.46
r94 45 47 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.49 $Y=1.46 $X2=0.67
+ $Y2=1.46
r95 43 48 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.33 $Y=1.567
+ $X2=0.67 $Y2=1.567
r96 42 45 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.33 $Y=1.46
+ $X2=0.49 $Y2=1.46
r97 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.33
+ $Y=1.46 $X2=0.33 $Y2=1.46
r98 36 55 0.299336 $w=3.83e-07 $l=1e-08 $layer=LI1_cond $X=1.68 $Y=1.567
+ $X2=1.69 $Y2=1.567
r99 36 52 9.87808 $w=3.83e-07 $l=3.3e-07 $layer=LI1_cond $X=1.68 $Y=1.567
+ $X2=1.35 $Y2=1.567
r100 35 52 4.49004 $w=3.83e-07 $l=1.5e-07 $layer=LI1_cond $X=1.2 $Y=1.567
+ $X2=1.35 $Y2=1.567
r101 34 35 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.567
+ $X2=1.2 $Y2=1.567
r102 34 48 1.49668 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=0.72 $Y=1.567
+ $X2=0.67 $Y2=1.567
r103 33 43 2.69402 $w=3.83e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=1.567
+ $X2=0.33 $Y2=1.567
r104 29 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.625
+ $X2=1.78 $Y2=1.46
r105 29 31 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.78 $Y=1.625
+ $X2=1.78 $Y2=2.465
r106 25 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.295
+ $X2=1.78 $Y2=1.46
r107 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.78 $Y=1.295
+ $X2=1.78 $Y2=0.655
r108 21 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.625
+ $X2=1.35 $Y2=1.46
r109 21 23 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.35 $Y=1.625
+ $X2=1.35 $Y2=2.465
r110 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.295
+ $X2=1.35 $Y2=1.46
r111 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.35 $Y=1.295
+ $X2=1.35 $Y2=0.655
r112 13 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.625
+ $X2=0.92 $Y2=1.46
r113 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.92 $Y=1.625
+ $X2=0.92 $Y2=2.465
r114 9 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.295
+ $X2=0.92 $Y2=1.46
r115 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.92 $Y=1.295
+ $X2=0.92 $Y2=0.655
r116 5 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.625
+ $X2=0.49 $Y2=1.46
r117 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.49 $Y=1.625
+ $X2=0.49 $Y2=2.465
r118 1 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.295
+ $X2=0.49 $Y2=1.46
r119 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.49 $Y=1.295 $X2=0.49
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%B1 3 7 11 15 19 23 27 31 33 34 35 36 63
c89 36 0 1.97252e-19 $X=3.6 $Y=1.665
c90 27 0 4.86632e-20 $X=3.5 $Y=0.655
c91 7 0 9.07802e-20 $X=2.245 $Y=2.465
c92 3 0 5.86634e-20 $X=2.21 $Y=0.655
r93 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.59
+ $Y=1.51 $X2=3.59 $Y2=1.51
r94 61 63 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.535 $Y=1.51
+ $X2=3.59 $Y2=1.51
r95 60 61 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.5 $Y=1.51
+ $X2=3.535 $Y2=1.51
r96 59 64 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=3.25 $Y=1.592
+ $X2=3.59 $Y2=1.592
r97 58 60 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.25 $Y=1.51 $X2=3.5
+ $Y2=1.51
r98 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.51 $X2=3.25 $Y2=1.51
r99 56 58 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.105 $Y=1.51
+ $X2=3.25 $Y2=1.51
r100 55 56 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.07 $Y=1.51
+ $X2=3.105 $Y2=1.51
r101 53 55 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.91 $Y=1.51
+ $X2=3.07 $Y2=1.51
r102 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.51 $X2=2.91 $Y2=1.51
r103 51 53 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=2.675 $Y=1.51
+ $X2=2.91 $Y2=1.51
r104 50 51 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.64 $Y=1.51
+ $X2=2.675 $Y2=1.51
r105 48 50 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.57 $Y=1.51 $X2=2.64
+ $Y2=1.51
r106 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.51 $X2=2.57 $Y2=1.51
r107 46 48 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=2.245 $Y=1.51
+ $X2=2.57 $Y2=1.51
r108 45 49 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.23 $Y=1.592
+ $X2=2.57 $Y2=1.592
r109 44 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.23 $Y=1.51
+ $X2=2.245 $Y2=1.51
r110 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.51 $X2=2.23 $Y2=1.51
r111 41 44 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.21 $Y=1.51 $X2=2.23
+ $Y2=1.51
r112 36 64 0.344013 $w=3.33e-07 $l=1e-08 $layer=LI1_cond $X=3.6 $Y=1.592
+ $X2=3.59 $Y2=1.592
r113 35 59 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.592
+ $X2=3.25 $Y2=1.592
r114 35 54 7.22427 $w=3.33e-07 $l=2.1e-07 $layer=LI1_cond $X=3.12 $Y=1.592
+ $X2=2.91 $Y2=1.592
r115 34 54 9.28835 $w=3.33e-07 $l=2.7e-07 $layer=LI1_cond $X=2.64 $Y=1.592
+ $X2=2.91 $Y2=1.592
r116 34 49 2.40809 $w=3.33e-07 $l=7e-08 $layer=LI1_cond $X=2.64 $Y=1.592
+ $X2=2.57 $Y2=1.592
r117 33 45 2.40809 $w=3.33e-07 $l=7e-08 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=2.23 $Y2=1.592
r118 29 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.675
+ $X2=3.535 $Y2=1.51
r119 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.535 $Y=1.675
+ $X2=3.535 $Y2=2.465
r120 25 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.5 $Y=1.345
+ $X2=3.5 $Y2=1.51
r121 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.5 $Y=1.345
+ $X2=3.5 $Y2=0.655
r122 21 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.675
+ $X2=3.105 $Y2=1.51
r123 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.105 $Y=1.675
+ $X2=3.105 $Y2=2.465
r124 17 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.345
+ $X2=3.07 $Y2=1.51
r125 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.07 $Y=1.345
+ $X2=3.07 $Y2=0.655
r126 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.675
+ $X2=2.675 $Y2=1.51
r127 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.675 $Y=1.675
+ $X2=2.675 $Y2=2.465
r128 9 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=1.345
+ $X2=2.64 $Y2=1.51
r129 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.64 $Y=1.345
+ $X2=2.64 $Y2=0.655
r130 5 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.245 $Y=1.675
+ $X2=2.245 $Y2=1.51
r131 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.245 $Y=1.675
+ $X2=2.245 $Y2=2.465
r132 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.345
+ $X2=2.21 $Y2=1.51
r133 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.21 $Y=1.345
+ $X2=2.21 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%A3 3 7 11 15 19 23 27 31 33 34 35 36 60
c90 60 0 1.97252e-19 $X=5.775 $Y=1.42
c91 36 0 4.86632e-20 $X=5.52 $Y=1.665
c92 23 0 6.32785e-20 $X=5.345 $Y=2.375
r93 58 60 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=5.49 $Y=1.42
+ $X2=5.775 $Y2=1.42
r94 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.49
+ $Y=1.42 $X2=5.49 $Y2=1.42
r95 56 58 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.47 $Y=1.42 $X2=5.49
+ $Y2=1.42
r96 55 56 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.345 $Y=1.42
+ $X2=5.47 $Y2=1.42
r97 54 59 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=5.15 $Y=1.547
+ $X2=5.49 $Y2=1.547
r98 53 55 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.15 $Y=1.42
+ $X2=5.345 $Y2=1.42
r99 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.15
+ $Y=1.42 $X2=5.15 $Y2=1.42
r100 51 53 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.97 $Y=1.42
+ $X2=5.15 $Y2=1.42
r101 50 51 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=4.915 $Y=1.42
+ $X2=4.97 $Y2=1.42
r102 48 50 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=4.81 $Y=1.42
+ $X2=4.915 $Y2=1.42
r103 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.81
+ $Y=1.42 $X2=4.81 $Y2=1.42
r104 46 48 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=4.485 $Y=1.42
+ $X2=4.81 $Y2=1.42
r105 44 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.47 $Y=1.42
+ $X2=4.485 $Y2=1.42
r106 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.47
+ $Y=1.42 $X2=4.47 $Y2=1.42
r107 41 44 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.04 $Y=1.42
+ $X2=4.47 $Y2=1.42
r108 36 59 0.813489 $w=4.23e-07 $l=3e-08 $layer=LI1_cond $X=5.52 $Y=1.547
+ $X2=5.49 $Y2=1.547
r109 35 54 2.98279 $w=4.23e-07 $l=1.1e-07 $layer=LI1_cond $X=5.04 $Y=1.547
+ $X2=5.15 $Y2=1.547
r110 35 49 6.23675 $w=4.23e-07 $l=2.3e-07 $layer=LI1_cond $X=5.04 $Y=1.547
+ $X2=4.81 $Y2=1.547
r111 34 49 6.77908 $w=4.23e-07 $l=2.5e-07 $layer=LI1_cond $X=4.56 $Y=1.547
+ $X2=4.81 $Y2=1.547
r112 34 45 2.44047 $w=4.23e-07 $l=9e-08 $layer=LI1_cond $X=4.56 $Y=1.547
+ $X2=4.47 $Y2=1.547
r113 33 45 10.5754 $w=4.23e-07 $l=3.9e-07 $layer=LI1_cond $X=4.08 $Y=1.547
+ $X2=4.47 $Y2=1.547
r114 29 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.775 $Y=1.585
+ $X2=5.775 $Y2=1.42
r115 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.775 $Y=1.585
+ $X2=5.775 $Y2=2.375
r116 25 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.47 $Y=1.255
+ $X2=5.47 $Y2=1.42
r117 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.47 $Y=1.255 $X2=5.47
+ $Y2=0.655
r118 21 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.345 $Y=1.585
+ $X2=5.345 $Y2=1.42
r119 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.345 $Y=1.585
+ $X2=5.345 $Y2=2.375
r120 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.97 $Y=1.255
+ $X2=4.97 $Y2=1.42
r121 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.97 $Y=1.255 $X2=4.97
+ $Y2=0.655
r122 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.915 $Y=1.585
+ $X2=4.915 $Y2=1.42
r123 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.915 $Y=1.585
+ $X2=4.915 $Y2=2.375
r124 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.485 $Y=1.585
+ $X2=4.485 $Y2=1.42
r125 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.485 $Y=1.585
+ $X2=4.485 $Y2=2.375
r126 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.47 $Y=1.255
+ $X2=4.47 $Y2=1.42
r127 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.47 $Y=1.255 $X2=4.47
+ $Y2=0.655
r128 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.04 $Y=1.255
+ $X2=4.04 $Y2=1.42
r129 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.04 $Y=1.255 $X2=4.04
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%A2 3 5 7 10 12 14 17 19 21 24 26 27 28 30 31
+ 32 33 34 52
r84 51 52 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=8.05
+ $Y=1.35 $X2=8.05 $Y2=1.35
r85 48 49 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=7.225 $Y=1.35
+ $X2=7.495 $Y2=1.35
r86 47 48 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=7.065 $Y=1.35
+ $X2=7.225 $Y2=1.35
r87 46 47 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=6.795 $Y=1.35
+ $X2=7.065 $Y2=1.35
r88 45 46 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.635 $Y=1.35
+ $X2=6.795 $Y2=1.35
r89 44 45 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=6.365 $Y=1.35
+ $X2=6.635 $Y2=1.35
r90 42 44 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.35 $Y=1.35
+ $X2=6.365 $Y2=1.35
r91 42 43 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=6.35
+ $Y=1.35 $X2=6.35 $Y2=1.35
r92 39 42 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=6.205 $Y=1.35
+ $X2=6.35 $Y2=1.35
r93 34 52 5.25676 $w=2.83e-07 $l=1.3e-07 $layer=LI1_cond $X=7.92 $Y=1.352
+ $X2=8.05 $Y2=1.352
r94 33 34 19.4096 $w=2.83e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.352
+ $X2=7.92 $Y2=1.352
r95 32 33 19.4096 $w=2.83e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.352
+ $X2=7.44 $Y2=1.352
r96 31 32 19.4096 $w=2.83e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.352
+ $X2=6.96 $Y2=1.352
r97 31 43 5.25676 $w=2.83e-07 $l=1.3e-07 $layer=LI1_cond $X=6.48 $Y=1.352
+ $X2=6.35 $Y2=1.352
r98 28 51 20.1791 $w=1.5e-07 $l=1.9139e-07 $layer=POLY_cond $X=8.025 $Y=1.185
+ $X2=8.082 $Y2=1.35
r99 28 30 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.025 $Y=1.185
+ $X2=8.025 $Y2=0.655
r100 27 49 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.57 $Y=1.35
+ $X2=7.495 $Y2=1.35
r101 26 51 11.9984 $w=3.3e-07 $l=1.32e-07 $layer=POLY_cond $X=7.95 $Y=1.35
+ $X2=8.082 $Y2=1.35
r102 26 27 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=7.95 $Y=1.35
+ $X2=7.57 $Y2=1.35
r103 22 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.495 $Y=1.515
+ $X2=7.495 $Y2=1.35
r104 22 24 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.495 $Y=1.515
+ $X2=7.495 $Y2=2.375
r105 19 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.225 $Y=1.185
+ $X2=7.225 $Y2=1.35
r106 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.225 $Y=1.185
+ $X2=7.225 $Y2=0.655
r107 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.065 $Y=1.515
+ $X2=7.065 $Y2=1.35
r108 15 17 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.065 $Y=1.515
+ $X2=7.065 $Y2=2.375
r109 12 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.185
+ $X2=6.795 $Y2=1.35
r110 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.795 $Y=1.185
+ $X2=6.795 $Y2=0.655
r111 8 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.635 $Y=1.515
+ $X2=6.635 $Y2=1.35
r112 8 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.635 $Y=1.515
+ $X2=6.635 $Y2=2.375
r113 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.185
+ $X2=6.365 $Y2=1.35
r114 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.365 $Y=1.185
+ $X2=6.365 $Y2=0.655
r115 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.515
+ $X2=6.205 $Y2=1.35
r116 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.205 $Y=1.515
+ $X2=6.205 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 39 50
r69 49 50 13.628 $w=4.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.79 $Y=1.425
+ $X2=9.865 $Y2=1.425
r70 48 49 47.9297 $w=4.8e-07 $l=4.3e-07 $layer=POLY_cond $X=9.36 $Y=1.425
+ $X2=9.79 $Y2=1.425
r71 47 48 47.9297 $w=4.8e-07 $l=4.3e-07 $layer=POLY_cond $X=8.93 $Y=1.425
+ $X2=9.36 $Y2=1.425
r72 45 47 37.8979 $w=4.8e-07 $l=3.4e-07 $layer=POLY_cond $X=8.59 $Y=1.425
+ $X2=8.93 $Y2=1.425
r73 45 46 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=8.59
+ $Y=1.35 $X2=8.59 $Y2=1.35
r74 42 45 10.0318 $w=4.8e-07 $l=9e-08 $layer=POLY_cond $X=8.5 $Y=1.425 $X2=8.59
+ $Y2=1.425
r75 39 50 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=10.29 $Y=1.35
+ $X2=9.865 $Y2=1.35
r76 32 39 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=10.29
+ $Y=1.35 $X2=10.29 $Y2=1.35
r77 31 32 18.1965 $w=2.83e-07 $l=4.5e-07 $layer=LI1_cond $X=9.84 $Y=1.352
+ $X2=10.29 $Y2=1.352
r78 30 31 19.4096 $w=2.83e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.352
+ $X2=9.84 $Y2=1.352
r79 29 30 19.4096 $w=2.83e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.352
+ $X2=9.36 $Y2=1.352
r80 29 46 11.7266 $w=2.83e-07 $l=2.9e-07 $layer=LI1_cond $X=8.88 $Y=1.352
+ $X2=8.59 $Y2=1.352
r81 25 49 30.3798 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.79 $Y=1.665
+ $X2=9.79 $Y2=1.425
r82 25 27 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=9.79 $Y=1.665 $X2=9.79
+ $Y2=2.465
r83 22 49 30.3798 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.79 $Y=1.185
+ $X2=9.79 $Y2=1.425
r84 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.79 $Y=1.185
+ $X2=9.79 $Y2=0.655
r85 18 48 30.3798 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.36 $Y=1.665
+ $X2=9.36 $Y2=1.425
r86 18 20 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=9.36 $Y=1.665 $X2=9.36
+ $Y2=2.465
r87 15 48 30.3798 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.36 $Y=1.185
+ $X2=9.36 $Y2=1.425
r88 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.36 $Y=1.185
+ $X2=9.36 $Y2=0.655
r89 11 47 30.3798 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.93 $Y=1.665
+ $X2=8.93 $Y2=1.425
r90 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=8.93 $Y=1.665 $X2=8.93
+ $Y2=2.465
r91 8 47 30.3798 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.93 $Y=1.185
+ $X2=8.93 $Y2=1.425
r92 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.93 $Y=1.185
+ $X2=8.93 $Y2=0.655
r93 4 42 30.3798 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.5 $Y=1.665 $X2=8.5
+ $Y2=1.425
r94 4 6 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=8.5 $Y=1.665 $X2=8.5
+ $Y2=2.465
r95 1 42 30.3798 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.5 $Y=1.185 $X2=8.5
+ $Y2=1.425
r96 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.5 $Y=1.185 $X2=8.5
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%A_30_367# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 34 40 44 46
r54 35 44 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.985 $Y=2.36
+ $X2=2.89 $Y2=2.36
r55 34 46 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=3.655 $Y=2.36
+ $X2=3.785 $Y2=2.36
r56 34 35 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.655 $Y=2.36
+ $X2=2.985 $Y2=2.36
r57 31 42 3.50369 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.125 $Y=2.36
+ $X2=2.03 $Y2=2.36
r58 30 44 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.795 $Y=2.36
+ $X2=2.89 $Y2=2.36
r59 30 31 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.795 $Y=2.36
+ $X2=2.125 $Y2=2.36
r60 28 42 3.31928 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=2.03 $Y=2.45 $X2=2.03
+ $Y2=2.36
r61 28 29 26.5598 $w=1.88e-07 $l=4.55e-07 $layer=LI1_cond $X=2.03 $Y=2.45
+ $X2=2.03 $Y2=2.905
r62 27 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.23 $Y=2.99
+ $X2=1.135 $Y2=2.99
r63 26 29 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.935 $Y=2.99
+ $X2=2.03 $Y2=2.905
r64 26 27 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.935 $Y=2.99
+ $X2=1.23 $Y2=2.99
r65 22 40 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=2.905
+ $X2=1.135 $Y2=2.99
r66 22 24 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=1.135 $Y=2.905
+ $X2=1.135 $Y2=2.435
r67 21 39 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.37 $Y=2.99 $X2=0.24
+ $Y2=2.99
r68 20 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.04 $Y=2.99
+ $X2=1.135 $Y2=2.99
r69 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.04 $Y=2.99
+ $X2=0.37 $Y2=2.99
r70 16 39 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.905
+ $X2=0.24 $Y2=2.99
r71 16 18 35.4598 $w=2.58e-07 $l=8e-07 $layer=LI1_cond $X=0.24 $Y=2.905 $X2=0.24
+ $Y2=2.105
r72 5 46 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=3.61
+ $Y=1.835 $X2=3.75 $Y2=2.435
r73 4 44 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=2.75
+ $Y=1.835 $X2=2.89 $Y2=2.435
r74 3 42 300 $w=1.7e-07 $l=6.81909e-07 $layer=licon1_PDIFF $count=2 $X=1.855
+ $Y=1.835 $X2=2.03 $Y2=2.435
r75 2 24 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.435
r76 1 39 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.91
r77 1 18 400 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%Y 1 2 3 4 5 6 7 8 29 31 32 33 37 39 43 45 49
+ 51 55 57 60 62 63 64 65 66 68 71 73 74
c160 71 0 6.32785e-20 $X=5.92 $Y=2.015
r161 73 79 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.582 $Y=2.015
+ $X2=1.582 $Y2=2.1
r162 73 74 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.582 $Y=2.11
+ $X2=1.582 $Y2=2.405
r163 73 79 0.315738 $w=3.63e-07 $l=1e-08 $layer=LI1_cond $X=1.582 $Y=2.11
+ $X2=1.582 $Y2=2.1
r164 66 73 102.368 $w=3.18e-07 $l=2.805e-06 $layer=LI1_cond $X=4.57 $Y=2.015
+ $X2=1.765 $Y2=2.015
r165 66 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.57 $Y=2.015
+ $X2=4.695 $Y2=2.015
r166 60 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=1.93
+ $X2=5.92 $Y2=2.015
r167 59 60 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.92 $Y=1.165
+ $X2=5.92 $Y2=1.93
r168 57 71 24.3348 $w=1.68e-07 $l=3.73e-07 $layer=LI1_cond $X=5.547 $Y=2.015
+ $X2=5.92 $Y2=2.015
r169 56 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.82 $Y=2.015
+ $X2=4.695 $Y2=2.015
r170 55 57 8.61176 $w=1.68e-07 $l=1.32e-07 $layer=LI1_cond $X=5.415 $Y=2.015
+ $X2=5.547 $Y2=2.015
r171 55 56 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.415 $Y=2.015
+ $X2=4.82 $Y2=2.015
r172 52 65 5.66127 $w=1.7e-07 $l=1.12472e-07 $layer=LI1_cond $X=3.41 $Y=1.08
+ $X2=3.3 $Y2=1.085
r173 51 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.835 $Y=1.08
+ $X2=5.92 $Y2=1.165
r174 51 52 158.209 $w=1.68e-07 $l=2.425e-06 $layer=LI1_cond $X=5.835 $Y=1.08
+ $X2=3.41 $Y2=1.08
r175 47 65 0.945268 $w=1.9e-07 $l=9.72111e-08 $layer=LI1_cond $X=3.285 $Y=0.995
+ $X2=3.3 $Y2=1.085
r176 47 49 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=3.285 $Y=0.995
+ $X2=3.285 $Y2=0.78
r177 46 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.52 $Y=1.09
+ $X2=2.425 $Y2=1.09
r178 45 65 5.66127 $w=1.7e-07 $l=1.12472e-07 $layer=LI1_cond $X=3.19 $Y=1.09
+ $X2=3.3 $Y2=1.085
r179 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.19 $Y=1.09
+ $X2=2.52 $Y2=1.09
r180 41 64 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=1.005
+ $X2=2.425 $Y2=1.09
r181 41 43 14.3014 $w=1.88e-07 $l=2.45e-07 $layer=LI1_cond $X=2.425 $Y=1.005
+ $X2=2.425 $Y2=0.76
r182 40 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.66 $Y=1.09
+ $X2=1.565 $Y2=1.09
r183 39 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.33 $Y=1.09
+ $X2=2.425 $Y2=1.09
r184 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.33 $Y=1.09
+ $X2=1.66 $Y2=1.09
r185 35 63 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=1.005
+ $X2=1.565 $Y2=1.09
r186 35 37 14.3014 $w=1.88e-07 $l=2.45e-07 $layer=LI1_cond $X=1.565 $Y=1.005
+ $X2=1.565 $Y2=0.76
r187 34 62 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=2.015
+ $X2=0.705 $Y2=2.015
r188 33 73 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.4 $Y=2.015
+ $X2=1.582 $Y2=2.015
r189 33 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.4 $Y=2.015
+ $X2=0.87 $Y2=2.015
r190 31 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.47 $Y=1.09
+ $X2=1.565 $Y2=1.09
r191 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.47 $Y=1.09
+ $X2=0.8 $Y2=1.09
r192 27 32 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.685 $Y=1.005
+ $X2=0.8 $Y2=1.09
r193 27 29 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.685 $Y=1.005
+ $X2=0.685 $Y2=0.76
r194 8 57 300 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=2 $X=5.42
+ $Y=1.745 $X2=5.56 $Y2=2.095
r195 7 68 300 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=2 $X=4.56
+ $Y=1.745 $X2=4.7 $Y2=2.095
r196 6 73 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=2.095
r197 5 62 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.095
r198 4 49 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.235 $X2=3.285 $Y2=0.78
r199 3 43 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.285
+ $Y=0.235 $X2=2.425 $Y2=0.76
r200 2 37 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=1.425
+ $Y=0.235 $X2=1.565 $Y2=0.76
r201 1 29 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.705 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%VPWR 1 2 3 4 5 18 22 26 32 38 43 44 46 47 49
+ 50 52 53 55 56 57 82 83
r127 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r128 80 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r129 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r130 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r131 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r132 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r133 73 74 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 70 73 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r135 70 71 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r136 68 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r137 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r138 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r139 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r140 61 65 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r141 60 64 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 60 61 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r143 57 74 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=7.92 $Y2=3.33
r144 57 71 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=3.6 $Y2=3.33
r145 55 79 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=9.88 $Y=3.33 $X2=9.84
+ $Y2=3.33
r146 55 56 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.88 $Y=3.33
+ $X2=10.025 $Y2=3.33
r147 54 82 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=10.17 $Y=3.33
+ $X2=10.32 $Y2=3.33
r148 54 56 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.17 $Y=3.33
+ $X2=10.025 $Y2=3.33
r149 52 76 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=8.98 $Y=3.33 $X2=8.88
+ $Y2=3.33
r150 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.98 $Y=3.33
+ $X2=9.145 $Y2=3.33
r151 51 79 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=9.31 $Y=3.33
+ $X2=9.84 $Y2=3.33
r152 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.31 $Y=3.33
+ $X2=9.145 $Y2=3.33
r153 49 73 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=8.12 $Y=3.33 $X2=7.92
+ $Y2=3.33
r154 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.12 $Y=3.33
+ $X2=8.285 $Y2=3.33
r155 48 76 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.45 $Y=3.33
+ $X2=8.88 $Y2=3.33
r156 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.45 $Y=3.33
+ $X2=8.285 $Y2=3.33
r157 46 67 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.12 $Y2=3.33
r158 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.32 $Y2=3.33
r159 45 70 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.6 $Y2=3.33
r160 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.32 $Y2=3.33
r161 43 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.16 $Y2=3.33
r162 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.46 $Y2=3.33
r163 42 67 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=3.12 $Y2=3.33
r164 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.46 $Y2=3.33
r165 38 41 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=10.025 $Y=1.98
+ $X2=10.025 $Y2=2.95
r166 36 56 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=10.025 $Y=3.245
+ $X2=10.025 $Y2=3.33
r167 36 41 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=10.025 $Y=3.245
+ $X2=10.025 $Y2=2.95
r168 32 35 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=9.145 $Y=2.09
+ $X2=9.145 $Y2=2.95
r169 30 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=3.33
r170 30 35 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=2.95
r171 26 29 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=8.285 $Y=2.09
+ $X2=8.285 $Y2=2.95
r172 24 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.285 $Y=3.245
+ $X2=8.285 $Y2=3.33
r173 24 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.285 $Y=3.245
+ $X2=8.285 $Y2=2.95
r174 20 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=3.245
+ $X2=3.32 $Y2=3.33
r175 20 22 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=3.32 $Y=3.245
+ $X2=3.32 $Y2=2.755
r176 16 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=3.245
+ $X2=2.46 $Y2=3.33
r177 16 18 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.46 $Y=3.245
+ $X2=2.46 $Y2=2.755
r178 5 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.865
+ $Y=1.835 $X2=10.005 $Y2=2.95
r179 5 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.865
+ $Y=1.835 $X2=10.005 $Y2=1.98
r180 4 35 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.005
+ $Y=1.835 $X2=9.145 $Y2=2.95
r181 4 32 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=9.005
+ $Y=1.835 $X2=9.145 $Y2=2.09
r182 3 29 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=8.16
+ $Y=1.835 $X2=8.285 $Y2=2.95
r183 3 26 400 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=8.16
+ $Y=1.835 $X2=8.285 $Y2=2.09
r184 2 22 600 $w=1.7e-07 $l=9.87522e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.835 $X2=3.32 $Y2=2.755
r185 1 18 600 $w=1.7e-07 $l=9.87522e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.835 $X2=2.46 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%A_829_349# 1 2 3 4 5 18 20 21 24 26 30 32 36
+ 40 44 48 49 50
r62 44 47 26.9554 $w=2.93e-07 $l=6.9e-07 $layer=LI1_cond $X=7.727 $Y=2.17
+ $X2=7.727 $Y2=2.86
r63 42 47 1.75796 $w=2.93e-07 $l=4.5e-08 $layer=LI1_cond $X=7.727 $Y=2.905
+ $X2=7.727 $Y2=2.86
r64 41 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.975 $Y=2.99
+ $X2=6.845 $Y2=2.99
r65 40 42 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=7.58 $Y=2.99
+ $X2=7.727 $Y2=2.905
r66 40 41 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.58 $Y=2.99
+ $X2=6.975 $Y2=2.99
r67 36 39 30.5841 $w=2.58e-07 $l=6.9e-07 $layer=LI1_cond $X=6.845 $Y=2.17
+ $X2=6.845 $Y2=2.86
r68 34 50 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=2.905
+ $X2=6.845 $Y2=2.99
r69 34 39 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=6.845 $Y=2.905
+ $X2=6.845 $Y2=2.86
r70 33 49 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.12 $Y=2.99
+ $X2=5.985 $Y2=2.99
r71 32 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.715 $Y=2.99
+ $X2=6.845 $Y2=2.99
r72 32 33 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.715 $Y=2.99
+ $X2=6.12 $Y2=2.99
r73 28 49 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=2.905
+ $X2=5.985 $Y2=2.99
r74 28 30 20.061 $w=2.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.985 $Y=2.905
+ $X2=5.985 $Y2=2.435
r75 27 48 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.245 $Y=2.99
+ $X2=5.117 $Y2=2.99
r76 26 49 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.85 $Y=2.99
+ $X2=5.985 $Y2=2.99
r77 26 27 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.85 $Y=2.99
+ $X2=5.245 $Y2=2.99
r78 22 48 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.117 $Y=2.905
+ $X2=5.117 $Y2=2.99
r79 22 24 21.2411 $w=2.53e-07 $l=4.7e-07 $layer=LI1_cond $X=5.117 $Y=2.905
+ $X2=5.117 $Y2=2.435
r80 20 48 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.99 $Y=2.99
+ $X2=5.117 $Y2=2.99
r81 20 21 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.99 $Y=2.99
+ $X2=4.375 $Y2=2.99
r82 16 21 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.24 $Y=2.905
+ $X2=4.375 $Y2=2.99
r83 16 18 20.061 $w=2.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.24 $Y=2.905
+ $X2=4.24 $Y2=2.435
r84 5 47 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.57
+ $Y=1.745 $X2=7.71 $Y2=2.86
r85 5 44 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=7.57
+ $Y=1.745 $X2=7.71 $Y2=2.17
r86 4 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.71
+ $Y=1.745 $X2=6.85 $Y2=2.86
r87 4 36 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=6.71
+ $Y=1.745 $X2=6.85 $Y2=2.17
r88 3 30 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=5.85
+ $Y=1.745 $X2=5.99 $Y2=2.435
r89 2 24 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=1.745 $X2=5.13 $Y2=2.435
r90 1 18 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=4.145
+ $Y=1.745 $X2=4.27 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%A_1256_349# 1 2 3 4 15 19 20 23 27 31 35 39
+ 43 44
r45 39 41 46.5988 $w=2.28e-07 $l=9.3e-07 $layer=LI1_cond $X=9.595 $Y=1.98
+ $X2=9.595 $Y2=2.91
r46 37 39 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=9.595 $Y=1.835
+ $X2=9.595 $Y2=1.98
r47 36 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.81 $Y=1.75
+ $X2=8.715 $Y2=1.75
r48 35 37 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=9.48 $Y=1.75
+ $X2=9.595 $Y2=1.835
r49 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.48 $Y=1.75
+ $X2=8.81 $Y2=1.75
r50 31 33 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=8.715 $Y=1.98
+ $X2=8.715 $Y2=2.91
r51 29 44 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.715 $Y=1.835
+ $X2=8.715 $Y2=1.75
r52 29 31 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=8.715 $Y=1.835
+ $X2=8.715 $Y2=1.98
r53 28 43 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=7.41 $Y=1.75
+ $X2=7.277 $Y2=1.75
r54 27 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.62 $Y=1.75
+ $X2=8.715 $Y2=1.75
r55 27 28 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=8.62 $Y=1.75
+ $X2=7.41 $Y2=1.75
r56 23 25 30.4419 $w=2.63e-07 $l=7e-07 $layer=LI1_cond $X=7.277 $Y=1.87
+ $X2=7.277 $Y2=2.57
r57 21 43 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.277 $Y=1.835
+ $X2=7.277 $Y2=1.75
r58 21 23 1.52209 $w=2.63e-07 $l=3.5e-08 $layer=LI1_cond $X=7.277 $Y=1.835
+ $X2=7.277 $Y2=1.87
r59 19 43 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.145 $Y=1.75
+ $X2=7.277 $Y2=1.75
r60 19 20 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.145 $Y=1.75
+ $X2=6.545 $Y2=1.75
r61 15 17 31.1838 $w=2.53e-07 $l=6.9e-07 $layer=LI1_cond $X=6.417 $Y=1.87
+ $X2=6.417 $Y2=2.56
r62 13 20 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=6.417 $Y=1.835
+ $X2=6.545 $Y2=1.75
r63 13 15 1.58178 $w=2.53e-07 $l=3.5e-08 $layer=LI1_cond $X=6.417 $Y=1.835
+ $X2=6.417 $Y2=1.87
r64 4 41 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.435
+ $Y=1.835 $X2=9.575 $Y2=2.91
r65 4 39 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.435
+ $Y=1.835 $X2=9.575 $Y2=1.98
r66 3 33 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.835 $X2=8.715 $Y2=2.91
r67 3 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.835 $X2=8.715 $Y2=1.98
r68 2 25 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=7.14
+ $Y=1.745 $X2=7.28 $Y2=2.57
r69 2 23 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.14
+ $Y=1.745 $X2=7.28 $Y2=1.87
r70 1 17 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.745 $X2=6.42 $Y2=2.56
r71 1 15 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.745 $X2=6.42 $Y2=1.87
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%A_30_47# 1 2 3 4 5 6 7 8 9 10 11 36 38 39 42
+ 46 50 52 53 54 55 58 62 63 66 70 72 76 78 82 84 88 91 93 95 99 102 103 104 105
c164 95 0 5.86634e-20 $X=2.855 $Y=0.38
r165 101 102 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=0.54
+ $X2=5.59 $Y2=0.54
r166 86 88 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=10.04 $Y=0.87
+ $X2=10.04 $Y2=0.42
r167 85 105 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.24 $Y=0.955
+ $X2=9.145 $Y2=0.955
r168 84 86 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.91 $Y=0.955
+ $X2=10.04 $Y2=0.87
r169 84 85 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.91 $Y=0.955
+ $X2=9.24 $Y2=0.955
r170 80 105 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=0.87
+ $X2=9.145 $Y2=0.955
r171 80 82 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=9.145 $Y=0.87
+ $X2=9.145 $Y2=0.42
r172 79 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.38 $Y=0.955
+ $X2=8.245 $Y2=0.955
r173 78 105 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.05 $Y=0.955
+ $X2=9.145 $Y2=0.955
r174 78 79 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.05 $Y=0.955
+ $X2=8.38 $Y2=0.955
r175 74 104 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.245 $Y=0.87
+ $X2=8.245 $Y2=0.955
r176 74 76 19.2074 $w=2.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.245 $Y=0.87
+ $X2=8.245 $Y2=0.42
r177 73 103 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=7.14 $Y=0.955
+ $X2=7.027 $Y2=0.955
r178 72 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.11 $Y=0.955
+ $X2=8.245 $Y2=0.955
r179 72 73 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=8.11 $Y=0.955
+ $X2=7.14 $Y2=0.955
r180 68 103 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=7.027 $Y=0.87
+ $X2=7.027 $Y2=0.955
r181 68 70 23.0489 $w=2.23e-07 $l=4.5e-07 $layer=LI1_cond $X=7.027 $Y=0.87
+ $X2=7.027 $Y2=0.42
r182 66 103 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=6.915 $Y=0.955
+ $X2=7.027 $Y2=0.955
r183 66 67 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.915 $Y=0.955
+ $X2=6.345 $Y2=0.955
r184 63 101 2.51806 $w=5.68e-07 $l=1.2e-07 $layer=LI1_cond $X=5.875 $Y=0.54
+ $X2=5.755 $Y2=0.54
r185 63 65 4.61644 $w=5.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.875 $Y=0.54
+ $X2=6.095 $Y2=0.54
r186 62 67 3.8985 $w=5.32e-07 $l=4.92722e-07 $layer=LI1_cond $X=6.175 $Y=0.54
+ $X2=6.345 $Y2=0.955
r187 62 65 1.67871 $w=5.68e-07 $l=8e-08 $layer=LI1_cond $X=6.175 $Y=0.54
+ $X2=6.095 $Y2=0.54
r188 61 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.92 $Y=0.74
+ $X2=4.755 $Y2=0.74
r189 61 102 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.92 $Y=0.74
+ $X2=5.59 $Y2=0.74
r190 56 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=0.655
+ $X2=4.755 $Y2=0.74
r191 56 58 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.755 $Y=0.655
+ $X2=4.755 $Y2=0.375
r192 54 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=0.74
+ $X2=4.755 $Y2=0.74
r193 54 55 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.59 $Y=0.74
+ $X2=3.88 $Y2=0.74
r194 53 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.715 $Y=0.655
+ $X2=3.88 $Y2=0.74
r195 52 97 2.73294 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.715 $Y=0.445
+ $X2=3.715 $Y2=0.35
r196 52 53 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.715 $Y=0.445
+ $X2=3.715 $Y2=0.655
r197 51 95 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0.35
+ $X2=2.855 $Y2=0.35
r198 50 97 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=0.35
+ $X2=3.715 $Y2=0.35
r199 50 51 30.9378 $w=1.88e-07 $l=5.3e-07 $layer=LI1_cond $X=3.55 $Y=0.35
+ $X2=3.02 $Y2=0.35
r200 47 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=0.34
+ $X2=1.995 $Y2=0.34
r201 46 95 8.26956 $w=1.8e-07 $l=1.69926e-07 $layer=LI1_cond $X=2.69 $Y=0.34
+ $X2=2.855 $Y2=0.35
r202 46 47 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.69 $Y=0.34
+ $X2=2.16 $Y2=0.34
r203 43 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=0.34
+ $X2=1.135 $Y2=0.34
r204 42 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=0.34
+ $X2=1.995 $Y2=0.34
r205 42 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.83 $Y=0.34
+ $X2=1.3 $Y2=0.34
r206 38 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0.34
+ $X2=1.135 $Y2=0.34
r207 38 39 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.97 $Y=0.34
+ $X2=0.4 $Y2=0.34
r208 34 39 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=0.255 $Y=0.425
+ $X2=0.4 $Y2=0.34
r209 34 36 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=0.255 $Y=0.425
+ $X2=0.255 $Y2=0.44
r210 11 88 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.865
+ $Y=0.235 $X2=10.005 $Y2=0.42
r211 10 82 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.005
+ $Y=0.235 $X2=9.145 $Y2=0.42
r212 9 76 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.1
+ $Y=0.235 $X2=8.24 $Y2=0.42
r213 8 70 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.87
+ $Y=0.235 $X2=7.01 $Y2=0.42
r214 7 101 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=5.545
+ $Y=0.235 $X2=5.755 $Y2=0.36
r215 7 65 182 $w=1.7e-07 $l=6.89746e-07 $layer=licon1_NDIFF $count=1 $X=5.545
+ $Y=0.235 $X2=6.095 $Y2=0.55
r216 6 99 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=4.545
+ $Y=0.235 $X2=4.685 $Y2=0.74
r217 6 58 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.545
+ $Y=0.235 $X2=4.755 $Y2=0.375
r218 5 97 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.575
+ $Y=0.235 $X2=3.715 $Y2=0.36
r219 4 95 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.715
+ $Y=0.235 $X2=2.855 $Y2=0.38
r220 3 93 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.855
+ $Y=0.235 $X2=1.995 $Y2=0.38
r221 2 91 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.995
+ $Y=0.235 $X2=1.135 $Y2=0.38
r222 1 36 91 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_4%VGND 1 2 3 4 5 6 21 25 29 33 37 40 41 43 44
+ 46 47 49 50 51 63 67 80 81 84 88
r146 88 91 10.1572 $w=6.28e-07 $l=5.35e-07 $layer=LI1_cond $X=7.625 $Y=0
+ $X2=7.625 $Y2=0.535
r147 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r148 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r149 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r150 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.32 $Y2=0
r151 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r152 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r153 75 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r154 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r155 72 88 8.63246 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=7.94 $Y=0 $X2=7.625
+ $Y2=0
r156 72 74 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.94 $Y=0 $X2=8.4
+ $Y2=0
r157 71 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r158 71 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r159 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r160 68 84 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.745 $Y=0 $X2=6.575
+ $Y2=0
r161 68 70 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.96 $Y2=0
r162 67 88 8.63246 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=7.31 $Y=0 $X2=7.625
+ $Y2=0
r163 67 70 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.31 $Y=0 $X2=6.96
+ $Y2=0
r164 66 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r165 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r166 63 84 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.405 $Y=0 $X2=6.575
+ $Y2=0
r167 63 65 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=6.405 $Y=0 $X2=5.52
+ $Y2=0
r168 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r169 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r170 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r171 55 59 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r172 54 58 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r173 54 55 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r174 51 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.52 $Y2=0
r175 51 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.04 $Y2=0
r176 49 77 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=9.41 $Y=0 $X2=9.36
+ $Y2=0
r177 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.41 $Y=0 $X2=9.575
+ $Y2=0
r178 48 80 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=9.74 $Y=0 $X2=10.32
+ $Y2=0
r179 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.74 $Y=0 $X2=9.575
+ $Y2=0
r180 46 74 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.55 $Y=0 $X2=8.4
+ $Y2=0
r181 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.55 $Y=0 $X2=8.715
+ $Y2=0
r182 45 77 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r183 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=8.715
+ $Y2=0
r184 43 61 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=5.09 $Y=0 $X2=5.04
+ $Y2=0
r185 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.09 $Y=0 $X2=5.255
+ $Y2=0
r186 42 65 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.42 $Y=0 $X2=5.52
+ $Y2=0
r187 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.42 $Y=0 $X2=5.255
+ $Y2=0
r188 40 58 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.08
+ $Y2=0
r189 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.255
+ $Y2=0
r190 39 61 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=5.04
+ $Y2=0
r191 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.255
+ $Y2=0
r192 35 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.575 $Y=0.085
+ $X2=9.575 $Y2=0
r193 35 37 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=9.575 $Y=0.085
+ $X2=9.575 $Y2=0.535
r194 31 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.715 $Y=0.085
+ $X2=8.715 $Y2=0
r195 31 33 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.715 $Y=0.085
+ $X2=8.715 $Y2=0.535
r196 27 84 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.575 $Y=0.085
+ $X2=6.575 $Y2=0
r197 27 29 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=6.575 $Y=0.085
+ $X2=6.575 $Y2=0.36
r198 23 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.255 $Y=0.085
+ $X2=5.255 $Y2=0
r199 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.255 $Y=0.085
+ $X2=5.255 $Y2=0.36
r200 19 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0
r201 19 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0.36
r202 6 37 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=9.435
+ $Y=0.235 $X2=9.575 $Y2=0.535
r203 5 33 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=8.575
+ $Y=0.235 $X2=8.715 $Y2=0.535
r204 4 91 91 $w=1.7e-07 $l=6.42729e-07 $layer=licon1_NDIFF $count=2 $X=7.3
+ $Y=0.235 $X2=7.81 $Y2=0.535
r205 3 29 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=6.44
+ $Y=0.235 $X2=6.58 $Y2=0.36
r206 2 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.235 $X2=5.255 $Y2=0.36
r207 1 21 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.115
+ $Y=0.235 $X2=4.255 $Y2=0.36
.ends

