* File: sky130_fd_sc_lp__a41oi_lp.pex.spice
* Created: Wed Sep  2 09:29:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41OI_LP%A4 3 7 9 10 18
r27 16 18 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.585 $Y=0.975
+ $X2=0.775 $Y2=0.975
r28 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=0.975 $X2=0.585 $Y2=0.975
r29 13 16 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.545 $Y=0.975
+ $X2=0.585 $Y2=0.975
r30 10 17 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=0.975
+ $X2=0.585 $Y2=0.975
r31 9 17 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=0.975
+ $X2=0.585 $Y2=0.975
r32 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.775 $Y=0.81
+ $X2=0.775 $Y2=0.975
r33 5 7 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.775 $Y=0.81
+ $X2=0.775 $Y2=0.445
r34 1 13 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.14
+ $X2=0.545 $Y2=0.975
r35 1 3 349.077 $w=2.5e-07 $l=1.405e-06 $layer=POLY_cond $X=0.545 $Y=1.14
+ $X2=0.545 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_LP%A3 3 7 9 10 14 15
c39 3 0 6.44805e-20 $X=1.075 $Y=2.545
r40 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.615
+ $X2=1.075 $Y2=1.45
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.075
+ $Y=1.615 $X2=1.075 $Y2=1.615
r42 10 15 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=1.075 $Y2=1.615
r43 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.72 $Y2=1.615
r44 7 16 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.165 $Y=0.445
+ $X2=1.165 $Y2=1.45
r45 1 14 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.78
+ $X2=1.075 $Y2=1.615
r46 1 3 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.075 $Y=1.78
+ $X2=1.075 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_LP%A2 3 7 11 12 13 14 15 16 22
c46 13 0 6.44805e-20 $X=1.68 $Y=0.555
c47 3 0 1.60092e-19 $X=1.555 $Y=0.445
r48 15 16 12.6936 $w=3.43e-07 $l=3.8e-07 $layer=LI1_cond $X=1.622 $Y=1.285
+ $X2=1.622 $Y2=1.665
r49 15 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.615
+ $Y=1.285 $X2=1.615 $Y2=1.285
r50 14 15 12.0255 $w=3.43e-07 $l=3.6e-07 $layer=LI1_cond $X=1.622 $Y=0.925
+ $X2=1.622 $Y2=1.285
r51 13 14 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.622 $Y=0.555
+ $X2=1.622 $Y2=0.925
r52 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.615 $Y=1.625
+ $X2=1.615 $Y2=1.285
r53 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.625
+ $X2=1.615 $Y2=1.79
r54 10 22 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.12
+ $X2=1.615 $Y2=1.285
r55 7 12 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.605 $Y=2.545
+ $X2=1.605 $Y2=1.79
r56 3 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.555 $Y=0.445
+ $X2=1.555 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_LP%A1 3 5 7 11 12 13 17
r40 12 13 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.155 $Y=1.285
+ $X2=2.155 $Y2=1.665
r41 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.155
+ $Y=1.285 $X2=2.155 $Y2=1.285
r42 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.155 $Y=1.625
+ $X2=2.155 $Y2=1.285
r43 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.12
+ $X2=2.155 $Y2=1.285
r44 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.79
+ $X2=2.155 $Y2=1.625
r45 5 7 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.155 $Y=1.79
+ $X2=2.155 $Y2=2.545
r46 3 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.065 $Y=0.445
+ $X2=2.065 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_LP%B1 1 3 5 8 10 11 12 14 17 18 19 20 24 26
r53 24 26 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.285
+ $X2=2.745 $Y2=1.12
r54 19 20 11.998 $w=3.63e-07 $l=3.8e-07 $layer=LI1_cond $X=2.707 $Y=1.285
+ $X2=2.707 $Y2=1.665
r55 19 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.725
+ $Y=1.285 $X2=2.725 $Y2=1.285
r56 15 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.855 $Y=0.88
+ $X2=2.855 $Y2=0.805
r57 15 26 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.855 $Y=0.88
+ $X2=2.855 $Y2=1.12
r58 12 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.855 $Y=0.73
+ $X2=2.855 $Y2=0.805
r59 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.855 $Y=0.73
+ $X2=2.855 $Y2=0.445
r60 10 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.78 $Y=0.805
+ $X2=2.855 $Y2=0.805
r61 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.78 $Y=0.805
+ $X2=2.57 $Y2=0.805
r62 8 17 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.685 $Y=2.545
+ $X2=2.685 $Y2=1.79
r63 5 17 34.9505 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.745 $Y=1.605
+ $X2=2.745 $Y2=1.79
r64 4 24 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=2.745 $Y=1.305
+ $X2=2.745 $Y2=1.285
r65 4 5 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=2.745 $Y=1.305 $X2=2.745
+ $Y2=1.605
r66 1 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.495 $Y=0.73
+ $X2=2.57 $Y2=0.805
r67 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.495 $Y=0.73 $X2=2.495
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_LP%A_27_409# 1 2 3 12 16 17 20 24 28 32
r53 28 30 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.42 $Y=2.19 $X2=2.42
+ $Y2=2.9
r54 26 28 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.42 $Y=2.14 $X2=2.42
+ $Y2=2.19
r55 25 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=2.055
+ $X2=1.34 $Y2=2.055
r56 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.255 $Y=2.055
+ $X2=2.42 $Y2=2.14
r57 24 25 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.255 $Y=2.055
+ $X2=1.505 $Y2=2.055
r58 20 22 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.34 $Y=2.19 $X2=1.34
+ $Y2=2.9
r59 18 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.34 $Y=2.14 $X2=1.34
+ $Y2=2.055
r60 18 20 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.34 $Y=2.14 $X2=1.34
+ $Y2=2.19
r61 16 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=2.055
+ $X2=1.34 $Y2=2.055
r62 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.175 $Y=2.055
+ $X2=0.445 $Y2=2.055
r63 12 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.19 $X2=0.28
+ $Y2=2.9
r64 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.14
+ $X2=0.445 $Y2=2.055
r65 10 12 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.28 $Y=2.14 $X2=0.28
+ $Y2=2.19
r66 3 30 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=2.045 $X2=2.42 $Y2=2.9
r67 3 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=2.045 $X2=2.42 $Y2=2.19
r68 2 22 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.045 $X2=1.34 $Y2=2.9
r69 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.045 $X2=1.34 $Y2=2.19
r70 1 14 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r71 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_LP%VPWR 1 2 11 15 18 19 20 30 31 34
r41 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r45 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r47 22 24 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 20 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 20 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 20 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 18 24 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.87 $Y2=3.33
r53 17 27 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.87 $Y2=3.33
r55 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=3.33
r56 13 15 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=2.485
r57 9 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245 $X2=0.81
+ $Y2=3.33
r58 9 11 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.485
r59 2 15 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=1.73
+ $Y=2.045 $X2=1.87 $Y2=2.485
r60 1 11 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_LP%Y 1 2 7 8 11 17 18 19 22
c42 8 0 1.60092e-19 $X=2.445 $Y=0.855
r43 19 22 2.44894 $w=3.98e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0.555
+ $X2=2.245 $Y2=0.47
r44 17 18 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.012 $Y=2.19
+ $X2=3.012 $Y2=2.025
r45 15 19 6.19438 $w=3.98e-07 $l=2.15e-07 $layer=LI1_cond $X=2.245 $Y=0.77
+ $X2=2.245 $Y2=0.555
r46 13 18 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.155 $Y=0.94
+ $X2=3.155 $Y2=2.025
r47 9 17 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=3.012 $Y=2.252
+ $X2=3.012 $Y2=2.19
r48 9 11 17.0343 $w=4.53e-07 $l=6.48e-07 $layer=LI1_cond $X=3.012 $Y=2.252
+ $X2=3.012 $Y2=2.9
r49 8 15 8.37092 $w=1.7e-07 $l=2.38747e-07 $layer=LI1_cond $X=2.445 $Y=0.855
+ $X2=2.245 $Y2=0.77
r50 7 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.07 $Y=0.855
+ $X2=3.155 $Y2=0.94
r51 7 8 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.07 $Y=0.855
+ $X2=2.445 $Y2=0.855
r52 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.045 $X2=2.95 $Y2=2.19
r53 2 11 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.045 $X2=2.95 $Y2=2.9
r54 1 22 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.235 $X2=2.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_LP%VGND 1 2 9 11 13 15 17 22 28 32
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r43 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.56
+ $Y2=0
r45 23 25 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=0.725 $Y=0
+ $X2=2.64 $Y2=0
r46 22 31 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.132
+ $Y2=0
r47 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.64
+ $Y2=0
r48 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r49 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.56
+ $Y2=0
r51 17 19 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.24
+ $Y2=0
r52 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r53 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r54 11 31 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.132 $Y2=0
r55 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0.4
r56 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.56 $Y=0.085 $X2=0.56
+ $Y2=0
r57 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.56 $Y=0.085 $X2=0.56
+ $Y2=0.42
r58 2 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.235 $X2=3.07 $Y2=0.4
r59 1 9 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.415
+ $Y=0.235 $X2=0.56 $Y2=0.42
.ends

