* NGSPICE file created from sky130_fd_sc_lp__a2111oi_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2111oi_m A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_155_533# D1 Y VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.058e+11p ps=1.82e+06u
M1001 Y B1 VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=4.515e+11p ps=4.67e+06u
M1002 VGND A2 a_443_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1003 VGND C1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_299_533# VPB phighvt w=420000u l=150000u
+  ad=2.1e+11p pd=1.84e+06u as=2.289e+11p ps=2.77e+06u
M1005 a_443_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_299_533# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_227_533# C1 a_155_533# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 a_299_533# B1 a_227_533# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y D1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

