* File: sky130_fd_sc_lp__clkbuf_8.pxi.spice
* Created: Wed Sep  2 09:38:39 2020
* 
x_PM_SKY130_FD_SC_LP__CLKBUF_8%A N_A_M1005_g N_A_M1006_g N_A_M1011_g N_A_M1018_g
+ A A N_A_c_103_n PM_SKY130_FD_SC_LP__CLKBUF_8%A
x_PM_SKY130_FD_SC_LP__CLKBUF_8%A_110_47# N_A_110_47#_M1005_d N_A_110_47#_M1006_s
+ N_A_110_47#_M1003_g N_A_110_47#_M1000_g N_A_110_47#_M1008_g
+ N_A_110_47#_M1001_g N_A_110_47#_M1009_g N_A_110_47#_M1002_g
+ N_A_110_47#_M1010_g N_A_110_47#_M1004_g N_A_110_47#_M1014_g
+ N_A_110_47#_M1007_g N_A_110_47#_M1015_g N_A_110_47#_M1012_g
+ N_A_110_47#_M1017_g N_A_110_47#_M1013_g N_A_110_47#_M1019_g
+ N_A_110_47#_M1016_g N_A_110_47#_c_153_n N_A_110_47#_c_154_n
+ N_A_110_47#_c_155_n N_A_110_47#_c_177_n N_A_110_47#_c_156_n
+ PM_SKY130_FD_SC_LP__CLKBUF_8%A_110_47#
x_PM_SKY130_FD_SC_LP__CLKBUF_8%VPWR N_VPWR_M1006_d N_VPWR_M1018_d N_VPWR_M1001_s
+ N_VPWR_M1004_s N_VPWR_M1012_s N_VPWR_M1016_s N_VPWR_c_294_n N_VPWR_c_295_n
+ N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n N_VPWR_c_299_n N_VPWR_c_300_n
+ N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_305_n
+ N_VPWR_c_306_n N_VPWR_c_307_n VPWR N_VPWR_c_308_n N_VPWR_c_309_n
+ N_VPWR_c_293_n N_VPWR_c_311_n N_VPWR_c_312_n PM_SKY130_FD_SC_LP__CLKBUF_8%VPWR
x_PM_SKY130_FD_SC_LP__CLKBUF_8%X N_X_M1003_s N_X_M1009_s N_X_M1014_s N_X_M1017_s
+ N_X_M1000_d N_X_M1002_d N_X_M1007_d N_X_M1013_d N_X_c_371_n N_X_c_453_n
+ N_X_c_372_n N_X_c_373_n N_X_c_385_n N_X_c_374_n N_X_c_375_n N_X_c_457_n
+ N_X_c_376_n N_X_c_387_n N_X_c_377_n N_X_c_461_n N_X_c_378_n N_X_c_388_n
+ N_X_c_379_n N_X_c_465_n N_X_c_380_n N_X_c_381_n N_X_c_382_n N_X_c_383_n X X X
+ PM_SKY130_FD_SC_LP__CLKBUF_8%X
x_PM_SKY130_FD_SC_LP__CLKBUF_8%VGND N_VGND_M1005_s N_VGND_M1011_s N_VGND_M1008_d
+ N_VGND_M1010_d N_VGND_M1015_d N_VGND_M1019_d N_VGND_c_498_n N_VGND_c_499_n
+ N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n N_VGND_c_503_n N_VGND_c_504_n
+ N_VGND_c_505_n N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n N_VGND_c_509_n
+ N_VGND_c_510_n N_VGND_c_511_n VGND N_VGND_c_512_n N_VGND_c_513_n
+ N_VGND_c_514_n N_VGND_c_515_n N_VGND_c_516_n PM_SKY130_FD_SC_LP__CLKBUF_8%VGND
cc_1 VNB N_A_M1005_g 0.029779f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_M1006_g 0.00673252f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_A_M1011_g 0.0234436f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.445
cc_4 VNB N_A_M1018_g 0.00438735f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_5 VNB A 0.0377278f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A_c_103_n 0.115007f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.235
cc_7 VNB N_A_110_47#_M1003_g 0.0368045f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.9
cc_8 VNB N_A_110_47#_M1000_g 0.00887124f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.57
cc_9 VNB N_A_110_47#_M1008_g 0.0339835f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_10 VNB N_A_110_47#_M1001_g 0.00859472f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.235
cc_11 VNB N_A_110_47#_M1009_g 0.0339835f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.235
cc_12 VNB N_A_110_47#_M1002_g 0.00859472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_110_47#_M1010_g 0.0339835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_110_47#_M1004_g 0.00859472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_110_47#_M1014_g 0.0339634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_110_47#_M1007_g 0.00859221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_110_47#_M1015_g 0.0339274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_110_47#_M1012_g 0.0085582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_110_47#_M1017_g 0.0324784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_110_47#_M1013_g 0.00715497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_110_47#_M1019_g 0.0439172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_110_47#_M1016_g 0.00973407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_110_47#_c_153_n 0.00469476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_110_47#_c_154_n 0.00160831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_110_47#_c_155_n 0.00895475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_110_47#_c_156_n 0.159246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_293_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_371_n 0.00160391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_372_n 0.00524232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_373_n 0.00518582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_374_n 0.00211646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_375_n 0.00126237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_376_n 0.00524232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_377_n 0.00126237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_378_n 0.00573294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_379_n 0.0013724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_380_n 0.00214133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_381_n 0.00211646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_382_n 0.00214133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_383_n 0.00211646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB X 0.0496065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_498_n 0.0115134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_499_n 0.00454665f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.235
cc_44 VNB N_VGND_c_500_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.235
cc_45 VNB N_VGND_c_501_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_502_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_503_n 0.0154623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_504_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_505_n 0.0176102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_506_n 0.0167416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_507_n 0.00497572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_508_n 0.0160902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_509_n 0.00497395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_510_n 0.0154623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_511_n 0.00497395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_512_n 0.0154599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_513_n 0.0196454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_514_n 0.286305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_515_n 0.00497395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_516_n 0.00574315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VPB N_A_M1006_g 0.0277366f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_62 VPB N_A_M1018_g 0.020105f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_63 VPB N_A_110_47#_M1000_g 0.020105f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.57
cc_64 VPB N_A_110_47#_M1001_g 0.018242f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.235
cc_65 VPB N_A_110_47#_M1002_g 0.018242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_110_47#_M1004_g 0.018242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_110_47#_M1007_g 0.018242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_110_47#_M1012_g 0.018242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_110_47#_M1013_g 0.0182686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_110_47#_M1016_g 0.0236642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_110_47#_c_154_n 0.0041076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_294_n 0.0108797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_295_n 0.0515407f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.235
cc_74 VPB N_VPWR_c_296_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_297_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_298_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_299_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_300_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_301_n 0.0443002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_302_n 0.0166965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_303_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_304_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_305_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_306_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_307_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_308_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_309_n 0.0198045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_293_n 0.0628638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_311_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_312_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_X_c_385_n 0.00243419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_X_c_374_n 0.00435877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_X_c_387_n 0.00243419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_X_c_388_n 0.00383483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_X_c_381_n 0.00211646f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_X_c_383_n 0.00211646f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB X 0.0113498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 N_A_M1011_g N_A_110_47#_M1003_g 0.0238708f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_M1018_g N_A_110_47#_M1000_g 0.0238708f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_M1005_g N_A_110_47#_c_153_n 0.00433433f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A_M1011_g N_A_110_47#_c_153_n 0.00356184f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_102 A N_A_110_47#_c_153_n 0.0283784f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_103 N_A_c_103_n N_A_110_47#_c_153_n 0.0160208f $X=0.905 $Y=1.235 $X2=0 $Y2=0
cc_104 N_A_M1006_g N_A_110_47#_c_154_n 0.00745249f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A_M1018_g N_A_110_47#_c_154_n 0.00524359f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_106 A N_A_110_47#_c_154_n 0.00618736f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_107 N_A_c_103_n N_A_110_47#_c_154_n 0.00700563f $X=0.905 $Y=1.235 $X2=0 $Y2=0
cc_108 N_A_c_103_n N_A_110_47#_c_155_n 0.0240189f $X=0.905 $Y=1.235 $X2=0 $Y2=0
cc_109 A N_A_110_47#_c_177_n 0.0262538f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_110 N_A_c_103_n N_A_110_47#_c_177_n 0.0125522f $X=0.905 $Y=1.235 $X2=0 $Y2=0
cc_111 N_A_c_103_n N_A_110_47#_c_156_n 0.0238708f $X=0.905 $Y=1.235 $X2=0 $Y2=0
cc_112 N_A_M1006_g N_VPWR_c_295_n 0.00502529f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_113 A N_VPWR_c_295_n 0.0150693f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_114 N_A_c_103_n N_VPWR_c_295_n 0.00189058f $X=0.905 $Y=1.235 $X2=0 $Y2=0
cc_115 N_A_M1018_g N_VPWR_c_296_n 0.00199892f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_M1006_g N_VPWR_c_302_n 0.00585385f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_M1018_g N_VPWR_c_302_n 0.00585385f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_M1006_g N_VPWR_c_293_n 0.0116496f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_M1018_g N_VPWR_c_293_n 0.0106725f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A_M1005_g N_VGND_c_499_n 0.00369134f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_121 A N_VGND_c_499_n 0.0196051f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_122 N_A_c_103_n N_VGND_c_499_n 0.00130063f $X=0.905 $Y=1.235 $X2=0 $Y2=0
cc_123 N_A_M1011_g N_VGND_c_500_n 0.0016983f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A_M1005_g N_VGND_c_506_n 0.00585385f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_M1011_g N_VGND_c_506_n 0.00585385f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_M1005_g N_VGND_c_514_n 0.0117419f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_127 N_A_M1011_g N_VGND_c_514_n 0.0107648f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_128 A N_VGND_c_514_n 0.00383899f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_129 N_A_110_47#_M1000_g N_VPWR_c_296_n 0.00199892f $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_A_110_47#_c_155_n N_VPWR_c_296_n 0.0100979f $X=3.245 $Y=1.32 $X2=0
+ $Y2=0
cc_131 N_A_110_47#_M1001_g N_VPWR_c_297_n 0.0016342f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_A_110_47#_M1002_g N_VPWR_c_297_n 0.0016342f $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_110_47#_M1004_g N_VPWR_c_298_n 0.0016342f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_110_47#_M1007_g N_VPWR_c_298_n 0.0016342f $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_110_47#_M1007_g N_VPWR_c_299_n 0.00585385f $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A_110_47#_M1012_g N_VPWR_c_299_n 0.00585385f $X=3.485 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A_110_47#_M1012_g N_VPWR_c_300_n 0.0016342f $X=3.485 $Y=2.465 $X2=0
+ $Y2=0
cc_138 N_A_110_47#_M1013_g N_VPWR_c_300_n 0.0016342f $X=3.915 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_110_47#_M1016_g N_VPWR_c_301_n 0.00343774f $X=4.345 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_110_47#_c_154_n N_VPWR_c_302_n 0.0145813f $X=0.69 $Y=2.04 $X2=0 $Y2=0
cc_141 N_A_110_47#_M1000_g N_VPWR_c_304_n 0.00585385f $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_110_47#_M1001_g N_VPWR_c_304_n 0.00585385f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_110_47#_M1002_g N_VPWR_c_306_n 0.00585385f $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_110_47#_M1004_g N_VPWR_c_306_n 0.00585385f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_110_47#_M1013_g N_VPWR_c_308_n 0.00585385f $X=3.915 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_110_47#_M1016_g N_VPWR_c_308_n 0.00585385f $X=4.345 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_110_47#_M1006_s N_VPWR_c_293_n 0.00327921f $X=0.55 $Y=1.835 $X2=0
+ $Y2=0
cc_148 N_A_110_47#_M1000_g N_VPWR_c_293_n 0.0106725f $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_110_47#_M1001_g N_VPWR_c_293_n 0.010584f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_110_47#_M1002_g N_VPWR_c_293_n 0.010584f $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_110_47#_M1004_g N_VPWR_c_293_n 0.010584f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_110_47#_M1007_g N_VPWR_c_293_n 0.010584f $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A_110_47#_M1012_g N_VPWR_c_293_n 0.010584f $X=3.485 $Y=2.465 $X2=0
+ $Y2=0
cc_154 N_A_110_47#_M1013_g N_VPWR_c_293_n 0.010584f $X=3.915 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_110_47#_M1016_g N_VPWR_c_293_n 0.0118837f $X=4.345 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_110_47#_c_154_n N_VPWR_c_293_n 0.00964167f $X=0.69 $Y=2.04 $X2=0
+ $Y2=0
cc_157 N_A_110_47#_M1003_g N_X_c_371_n 0.00120255f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_110_47#_M1008_g N_X_c_371_n 0.00120255f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_110_47#_c_153_n N_X_c_371_n 0.00257148f $X=0.69 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_110_47#_M1008_g N_X_c_372_n 0.0145447f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_110_47#_M1009_g N_X_c_372_n 0.0149644f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_110_47#_c_155_n N_X_c_372_n 0.0430995f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_163 N_A_110_47#_c_156_n N_X_c_372_n 0.0022464f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_164 N_A_110_47#_M1003_g N_X_c_373_n 0.00408223f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_110_47#_c_153_n N_X_c_373_n 0.00821626f $X=0.69 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A_110_47#_c_155_n N_X_c_373_n 0.0210442f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_167 N_A_110_47#_c_156_n N_X_c_373_n 0.00231555f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_168 N_A_110_47#_M1001_g N_X_c_385_n 0.0170144f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_110_47#_M1002_g N_X_c_385_n 0.0173341f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_110_47#_c_155_n N_X_c_385_n 0.0450553f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_171 N_A_110_47#_c_156_n N_X_c_385_n 0.0022602f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_172 N_A_110_47#_M1000_g N_X_c_374_n 0.00309564f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A_110_47#_c_154_n N_X_c_374_n 0.00633313f $X=0.69 $Y=2.04 $X2=0 $Y2=0
cc_174 N_A_110_47#_c_155_n N_X_c_374_n 0.0219298f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_175 N_A_110_47#_c_156_n N_X_c_374_n 0.00232957f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_176 N_A_110_47#_M1009_g N_X_c_375_n 0.00120255f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_177 N_A_110_47#_M1010_g N_X_c_375_n 0.00120255f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A_110_47#_M1010_g N_X_c_376_n 0.0150303f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_179 N_A_110_47#_M1014_g N_X_c_376_n 0.0150303f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_180 N_A_110_47#_c_155_n N_X_c_376_n 0.0430995f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_181 N_A_110_47#_c_156_n N_X_c_376_n 0.0022464f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_182 N_A_110_47#_M1004_g N_X_c_387_n 0.0174f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_110_47#_M1007_g N_X_c_387_n 0.0174f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_110_47#_c_155_n N_X_c_387_n 0.0450553f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_185 N_A_110_47#_c_156_n N_X_c_387_n 0.0022602f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_186 N_A_110_47#_M1014_g N_X_c_377_n 0.00120255f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A_110_47#_M1015_g N_X_c_377_n 0.00120255f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A_110_47#_M1015_g N_X_c_378_n 0.0150303f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_110_47#_c_155_n N_X_c_378_n 0.0134162f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_190 N_A_110_47#_c_156_n N_X_c_378_n 0.00385814f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_191 N_A_110_47#_M1012_g N_X_c_388_n 0.0174f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A_110_47#_c_155_n N_X_c_388_n 0.0140368f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_193 N_A_110_47#_c_156_n N_X_c_388_n 0.00390002f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_194 N_A_110_47#_M1017_g N_X_c_379_n 0.00120255f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_195 N_A_110_47#_M1019_g N_X_c_379_n 0.00221636f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_196 N_A_110_47#_c_155_n N_X_c_380_n 0.0210442f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_197 N_A_110_47#_c_156_n N_X_c_380_n 0.00231555f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_198 N_A_110_47#_c_155_n N_X_c_381_n 0.0219298f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_199 N_A_110_47#_c_156_n N_X_c_381_n 0.00232957f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_200 N_A_110_47#_c_155_n N_X_c_382_n 0.0210442f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_201 N_A_110_47#_c_156_n N_X_c_382_n 0.00231555f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_202 N_A_110_47#_c_155_n N_X_c_383_n 0.0219298f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_203 N_A_110_47#_c_156_n N_X_c_383_n 0.00232957f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_204 N_A_110_47#_M1015_g X 0.0047522f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A_110_47#_M1012_g X 0.00448672f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A_110_47#_M1017_g X 0.0185727f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_207 N_A_110_47#_M1013_g X 0.0053012f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A_110_47#_M1019_g X 0.0231544f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_209 N_A_110_47#_M1016_g X 0.00773738f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A_110_47#_c_155_n X 0.0276335f $X=3.245 $Y=1.32 $X2=0 $Y2=0
cc_211 N_A_110_47#_c_156_n X 0.036842f $X=4.345 $Y=1.32 $X2=0 $Y2=0
cc_212 N_A_110_47#_M1013_g X 0.0162565f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A_110_47#_M1016_g X 0.018257f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A_110_47#_M1003_g N_VGND_c_500_n 0.0016983f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_215 N_A_110_47#_c_155_n N_VGND_c_500_n 0.00793117f $X=3.245 $Y=1.32 $X2=0
+ $Y2=0
cc_216 N_A_110_47#_M1008_g N_VGND_c_501_n 0.0016342f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_217 N_A_110_47#_M1009_g N_VGND_c_501_n 0.0016342f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_A_110_47#_M1010_g N_VGND_c_502_n 0.0016342f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_219 N_A_110_47#_M1014_g N_VGND_c_502_n 0.0016342f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_220 N_A_110_47#_M1014_g N_VGND_c_503_n 0.00439206f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_110_47#_M1015_g N_VGND_c_503_n 0.00439206f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_222 N_A_110_47#_M1015_g N_VGND_c_504_n 0.0016342f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_223 N_A_110_47#_M1017_g N_VGND_c_504_n 0.0016342f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_A_110_47#_M1019_g N_VGND_c_505_n 0.00344007f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_225 N_A_110_47#_c_153_n N_VGND_c_506_n 0.0137139f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_226 N_A_110_47#_M1003_g N_VGND_c_508_n 0.00585385f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_227 N_A_110_47#_M1008_g N_VGND_c_508_n 0.00439206f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_228 N_A_110_47#_M1009_g N_VGND_c_510_n 0.00439206f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_229 N_A_110_47#_M1010_g N_VGND_c_510_n 0.00439206f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_230 N_A_110_47#_M1017_g N_VGND_c_512_n 0.00439071f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_231 N_A_110_47#_M1019_g N_VGND_c_512_n 0.00439071f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_232 N_A_110_47#_M1005_d N_VGND_c_514_n 0.0033672f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_233 N_A_110_47#_M1003_g N_VGND_c_514_n 0.0107648f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_234 N_A_110_47#_M1008_g N_VGND_c_514_n 0.0059518f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_235 N_A_110_47#_M1009_g N_VGND_c_514_n 0.0059518f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_236 N_A_110_47#_M1010_g N_VGND_c_514_n 0.0059518f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_237 N_A_110_47#_M1014_g N_VGND_c_514_n 0.0059518f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_238 N_A_110_47#_M1015_g N_VGND_c_514_n 0.0059518f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_239 N_A_110_47#_M1017_g N_VGND_c_514_n 0.00594932f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_240 N_A_110_47#_M1019_g N_VGND_c_514_n 0.00724901f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_241 N_A_110_47#_c_153_n N_VGND_c_514_n 0.0095959f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_293_n N_X_M1000_d 0.00293134f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_243 N_VPWR_c_293_n N_X_M1002_d 0.00293134f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_293_n N_X_M1007_d 0.00293134f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_c_293_n N_X_M1013_d 0.00293134f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_246 N_VPWR_c_304_n N_X_c_453_n 0.0149362f $X=1.85 $Y=3.33 $X2=0 $Y2=0
cc_247 N_VPWR_c_293_n N_X_c_453_n 0.0100304f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_248 N_VPWR_M1001_s N_X_c_385_n 0.00178346f $X=1.84 $Y=1.835 $X2=0 $Y2=0
cc_249 N_VPWR_c_297_n N_X_c_385_n 0.0138265f $X=1.98 $Y=2.23 $X2=0 $Y2=0
cc_250 N_VPWR_c_306_n N_X_c_457_n 0.0149362f $X=2.71 $Y=3.33 $X2=0 $Y2=0
cc_251 N_VPWR_c_293_n N_X_c_457_n 0.0100304f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_M1004_s N_X_c_387_n 0.00178346f $X=2.7 $Y=1.835 $X2=0 $Y2=0
cc_253 N_VPWR_c_298_n N_X_c_387_n 0.0138265f $X=2.84 $Y=2.23 $X2=0 $Y2=0
cc_254 N_VPWR_c_299_n N_X_c_461_n 0.0149362f $X=3.57 $Y=3.33 $X2=0 $Y2=0
cc_255 N_VPWR_c_293_n N_X_c_461_n 0.0100304f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_M1012_s N_X_c_388_n 0.00152561f $X=3.56 $Y=1.835 $X2=0 $Y2=0
cc_257 N_VPWR_c_300_n N_X_c_388_n 0.0118724f $X=3.7 $Y=2.23 $X2=0 $Y2=0
cc_258 N_VPWR_c_308_n N_X_c_465_n 0.0149362f $X=4.43 $Y=3.33 $X2=0 $Y2=0
cc_259 N_VPWR_c_293_n N_X_c_465_n 0.0100304f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_260 N_VPWR_M1012_s X 2.54524e-19 $X=3.56 $Y=1.835 $X2=0 $Y2=0
cc_261 N_VPWR_M1016_s X 0.00258406f $X=4.42 $Y=1.835 $X2=0 $Y2=0
cc_262 N_VPWR_c_300_n X 0.00207372f $X=3.7 $Y=2.23 $X2=0 $Y2=0
cc_263 N_VPWR_c_301_n X 0.0224079f $X=4.56 $Y=2.23 $X2=0 $Y2=0
cc_264 N_X_c_372_n N_VGND_c_501_n 0.0169367f $X=2.28 $Y=0.855 $X2=0 $Y2=0
cc_265 N_X_c_376_n N_VGND_c_502_n 0.0169367f $X=3.14 $Y=0.855 $X2=0 $Y2=0
cc_266 N_X_c_376_n N_VGND_c_503_n 0.00229795f $X=3.14 $Y=0.855 $X2=0 $Y2=0
cc_267 N_X_c_377_n N_VGND_c_503_n 0.0129148f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_268 N_X_c_378_n N_VGND_c_503_n 0.00229795f $X=3.76 $Y=0.855 $X2=0 $Y2=0
cc_269 N_X_c_378_n N_VGND_c_504_n 0.013324f $X=3.76 $Y=0.855 $X2=0 $Y2=0
cc_270 X N_VGND_c_504_n 0.00403165f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_271 X N_VGND_c_505_n 0.0243168f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_272 N_X_c_371_n N_VGND_c_508_n 0.0129148f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_273 N_X_c_372_n N_VGND_c_508_n 0.00229795f $X=2.28 $Y=0.855 $X2=0 $Y2=0
cc_274 N_X_c_372_n N_VGND_c_510_n 0.00229795f $X=2.28 $Y=0.855 $X2=0 $Y2=0
cc_275 N_X_c_375_n N_VGND_c_510_n 0.0129148f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_276 N_X_c_376_n N_VGND_c_510_n 0.00229795f $X=3.14 $Y=0.855 $X2=0 $Y2=0
cc_277 N_X_c_379_n N_VGND_c_512_n 0.0128989f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_278 X N_VGND_c_512_n 0.004977f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_279 N_X_M1003_s N_VGND_c_514_n 0.00268594f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_280 N_X_M1009_s N_VGND_c_514_n 0.00234583f $X=2.27 $Y=0.235 $X2=0 $Y2=0
cc_281 N_X_M1014_s N_VGND_c_514_n 0.00234583f $X=3.13 $Y=0.235 $X2=0 $Y2=0
cc_282 N_X_M1017_s N_VGND_c_514_n 0.00234553f $X=3.99 $Y=0.235 $X2=0 $Y2=0
cc_283 N_X_c_371_n N_VGND_c_514_n 0.00991486f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_284 N_X_c_372_n N_VGND_c_514_n 0.00851977f $X=2.28 $Y=0.855 $X2=0 $Y2=0
cc_285 N_X_c_375_n N_VGND_c_514_n 0.00991486f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_286 N_X_c_376_n N_VGND_c_514_n 0.00851977f $X=3.14 $Y=0.855 $X2=0 $Y2=0
cc_287 N_X_c_377_n N_VGND_c_514_n 0.00991486f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_288 N_X_c_378_n N_VGND_c_514_n 0.00449126f $X=3.76 $Y=0.855 $X2=0 $Y2=0
cc_289 N_X_c_379_n N_VGND_c_514_n 0.00990863f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_290 X N_VGND_c_514_n 0.00953214f $X=3.995 $Y=0.84 $X2=0 $Y2=0
