# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand4b_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nand4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.035000 0.435000 1.625000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 1.415000 2.735000 1.750000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.425000 4.715000 1.750000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.885000 1.425000 5.605000 1.750000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.659000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.595000 1.805000 1.075000 ;
        RECT 1.475000 1.075000 3.215000 1.245000 ;
        RECT 1.505000 1.920000 5.075000 2.090000 ;
        RECT 1.505000 2.090000 1.770000 3.075000 ;
        RECT 2.440000 2.090000 4.215000 2.120000 ;
        RECT 2.440000 2.120000 2.675000 3.075000 ;
        RECT 2.905000 1.245000 3.215000 1.920000 ;
        RECT 4.025000 2.120000 4.215000 3.075000 ;
        RECT 4.885000 2.090000 5.075000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.155000  0.300000 0.345000 0.695000 ;
      RECT 0.155000  0.695000 0.785000 0.865000 ;
      RECT 0.420000  1.895000 0.785000 2.225000 ;
      RECT 0.525000  0.085000 0.855000 0.525000 ;
      RECT 0.605000  0.865000 0.785000 1.415000 ;
      RECT 0.605000  1.415000 1.755000 1.645000 ;
      RECT 0.605000  1.645000 0.785000 1.895000 ;
      RECT 0.955000  1.815000 1.335000 3.245000 ;
      RECT 1.045000  0.255000 2.305000 0.425000 ;
      RECT 1.045000  0.425000 1.305000 1.185000 ;
      RECT 1.940000  2.260000 2.270000 3.245000 ;
      RECT 1.975000  0.425000 2.305000 0.725000 ;
      RECT 1.975000  0.725000 3.235000 0.905000 ;
      RECT 2.475000  0.255000 4.285000 0.425000 ;
      RECT 2.475000  0.425000 2.805000 0.555000 ;
      RECT 2.845000  2.290000 3.855000 3.245000 ;
      RECT 2.975000  0.645000 3.235000 0.725000 ;
      RECT 3.445000  0.595000 3.775000 1.085000 ;
      RECT 3.445000  1.085000 5.605000 1.255000 ;
      RECT 3.955000  0.425000 4.285000 0.915000 ;
      RECT 4.385000  2.260000 4.715000 3.245000 ;
      RECT 4.455000  0.325000 4.655000 1.085000 ;
      RECT 4.825000  0.085000 5.155000 0.915000 ;
      RECT 5.245000  1.920000 5.575000 3.245000 ;
      RECT 5.325000  0.325000 5.605000 1.085000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__nand4b_2
END LIBRARY
