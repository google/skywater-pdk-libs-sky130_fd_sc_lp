* File: sky130_fd_sc_lp__sleep_pargate_plv_21.spice
* Created: Fri Aug 28 11:32:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sleep_pargate_plv_21.pex.spice"
.subckt sky130_fd_sc_lp__sleep_pargate_plv_21  VPB SLEEP VPWR VIRTPWR
* 
* VIRTPWR	VIRTPWR
* VPWR	VPWR
* SLEEP	SLEEP
* VPB	VPB
MM1000 N_VIRTPWR_M1000_d N_SLEEP_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=7
+ AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 M=1 R=46.6667 SA=75000.2
+ SB=75001.1 A=1.05 P=14.3 MULT=1
MM1001 N_VIRTPWR_M1000_d N_SLEEP_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=7
+ AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 M=1 R=46.6667 SA=75000.6
+ SB=75000.6 A=1.05 P=14.3 MULT=1
MM1002 N_VIRTPWR_M1002_d N_SLEEP_M1002_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=7
+ AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 M=1 R=46.6667 SA=75001.1
+ SB=75000.2 A=1.05 P=14.3 MULT=1
DX3_noxref noxref_1 VPB NWDIODE A=20.4407 P=23.47
c_36 VPB 0 8.20372e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sleep_pargate_plv_21.pxi.spice"
*
.ends
*
*
