* File: sky130_fd_sc_lp__sdfxbp_lp.pxi.spice
* Created: Wed Sep  2 10:36:24 2020
* 
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_27_409# N_A_27_409#_M1037_s
+ N_A_27_409#_M1017_s N_A_27_409#_c_267_n N_A_27_409#_M1036_g
+ N_A_27_409#_M1015_g N_A_27_409#_c_259_n N_A_27_409#_c_260_n
+ N_A_27_409#_c_261_n N_A_27_409#_c_262_n N_A_27_409#_c_263_n
+ N_A_27_409#_c_264_n N_A_27_409#_c_265_n N_A_27_409#_c_266_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%D N_D_M1003_g N_D_M1019_g N_D_c_321_n
+ N_D_c_326_n D N_D_c_322_n N_D_c_323_n PM_SKY130_FD_SC_LP__SDFXBP_LP%D
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%SCE N_SCE_M1017_g N_SCE_M1037_g N_SCE_M1008_g
+ N_SCE_c_363_n N_SCE_c_364_n N_SCE_M1020_g N_SCE_c_366_n N_SCE_M1006_g SCE
+ N_SCE_c_367_n PM_SKY130_FD_SC_LP__SDFXBP_LP%SCE
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%SCD N_SCD_M1012_g N_SCD_c_438_n N_SCD_M1040_g
+ N_SCD_c_435_n SCD N_SCD_c_436_n N_SCD_c_437_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%SCD
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%CLK N_CLK_M1035_g N_CLK_M1005_g N_CLK_M1021_g
+ CLK CLK N_CLK_c_480_n PM_SKY130_FD_SC_LP__SDFXBP_LP%CLK
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1530_231# N_A_1530_231#_M1018_d
+ N_A_1530_231#_M1022_d N_A_1530_231#_M1013_d N_A_1530_231#_M1007_g
+ N_A_1530_231#_M1009_g N_A_1530_231#_c_518_n N_A_1530_231#_c_519_n
+ N_A_1530_231#_c_520_n N_A_1530_231#_c_521_n N_A_1530_231#_c_522_n
+ N_A_1530_231#_c_523_n N_A_1530_231#_c_524_n N_A_1530_231#_c_538_p
+ N_A_1530_231#_c_525_n PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1530_231#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1278_155# N_A_1278_155#_M1014_d
+ N_A_1278_155#_M1010_d N_A_1278_155#_M1028_g N_A_1278_155#_M1013_g
+ N_A_1278_155#_M1018_g N_A_1278_155#_c_613_n N_A_1278_155#_c_618_n
+ N_A_1278_155#_c_619_n N_A_1278_155#_c_614_n N_A_1278_155#_c_615_n
+ N_A_1278_155#_c_616_n PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1278_155#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_706_66# N_A_706_66#_M1035_s
+ N_A_706_66#_M1005_s N_A_706_66#_c_690_n N_A_706_66#_M1004_g
+ N_A_706_66#_M1030_g N_A_706_66#_M1039_g N_A_706_66#_c_693_n
+ N_A_706_66#_c_694_n N_A_706_66#_M1041_g N_A_706_66#_c_696_n
+ N_A_706_66#_c_697_n N_A_706_66#_M1038_g N_A_706_66#_c_699_n
+ N_A_706_66#_c_700_n N_A_706_66#_M1024_g N_A_706_66#_c_702_n
+ N_A_706_66#_M1042_g N_A_706_66#_c_703_n N_A_706_66#_c_704_n
+ N_A_706_66#_c_705_n N_A_706_66#_c_706_n N_A_706_66#_c_707_n
+ N_A_706_66#_c_715_n N_A_706_66#_c_708_n N_A_706_66#_c_709_n
+ N_A_706_66#_c_710_n N_A_706_66#_c_711_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%A_706_66#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_975_347# N_A_975_347#_M1039_d
+ N_A_975_347#_M1030_d N_A_975_347#_c_857_n N_A_975_347#_c_847_n
+ N_A_975_347#_c_848_n N_A_975_347#_c_858_n N_A_975_347#_c_859_n
+ N_A_975_347#_c_849_n N_A_975_347#_M1014_g N_A_975_347#_M1010_g
+ N_A_975_347#_c_861_n N_A_975_347#_M1033_g N_A_975_347#_M1022_g
+ N_A_975_347#_c_863_n N_A_975_347#_c_864_n N_A_975_347#_c_852_n
+ N_A_975_347#_c_865_n N_A_975_347#_c_853_n N_A_975_347#_c_854_n
+ N_A_975_347#_c_855_n N_A_975_347#_c_856_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%A_975_347#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_2089_254# N_A_2089_254#_M1002_d
+ N_A_2089_254#_M1000_d N_A_2089_254#_M1034_g N_A_2089_254#_c_949_n
+ N_A_2089_254#_c_950_n N_A_2089_254#_c_951_n N_A_2089_254#_M1001_g
+ N_A_2089_254#_M1032_g N_A_2089_254#_M1043_g N_A_2089_254#_M1025_g
+ N_A_2089_254#_M1011_g N_A_2089_254#_M1029_g N_A_2089_254#_M1023_g
+ N_A_2089_254#_c_957_n N_A_2089_254#_c_958_n N_A_2089_254#_c_959_n
+ N_A_2089_254#_c_960_n N_A_2089_254#_c_961_n N_A_2089_254#_c_962_n
+ N_A_2089_254#_c_963_n N_A_2089_254#_c_964_n N_A_2089_254#_c_965_n
+ N_A_2089_254#_c_976_n N_A_2089_254#_c_977_n N_A_2089_254#_c_966_n
+ N_A_2089_254#_c_967_n N_A_2089_254#_c_968_n N_A_2089_254#_c_969_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%A_2089_254#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1902_347# N_A_1902_347#_M1042_d
+ N_A_1902_347#_M1024_d N_A_1902_347#_M1000_g N_A_1902_347#_c_1119_n
+ N_A_1902_347#_M1016_g N_A_1902_347#_c_1120_n N_A_1902_347#_c_1121_n
+ N_A_1902_347#_c_1122_n N_A_1902_347#_M1002_g N_A_1902_347#_c_1123_n
+ N_A_1902_347#_c_1128_n N_A_1902_347#_c_1124_n N_A_1902_347#_c_1130_n
+ N_A_1902_347#_c_1125_n N_A_1902_347#_c_1132_n N_A_1902_347#_c_1126_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1902_347#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_2714_401# N_A_2714_401#_M1023_d
+ N_A_2714_401#_M1011_d N_A_2714_401#_M1027_g N_A_2714_401#_M1031_g
+ N_A_2714_401#_c_1212_n N_A_2714_401#_M1026_g N_A_2714_401#_c_1220_n
+ N_A_2714_401#_c_1221_n N_A_2714_401#_c_1222_n N_A_2714_401#_c_1214_n
+ N_A_2714_401#_c_1215_n N_A_2714_401#_c_1216_n N_A_2714_401#_c_1217_n
+ N_A_2714_401#_c_1218_n PM_SKY130_FD_SC_LP__SDFXBP_LP%A_2714_401#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%VPWR N_VPWR_M1017_d N_VPWR_M1006_d
+ N_VPWR_M1005_d N_VPWR_M1007_d N_VPWR_M1034_d N_VPWR_M1032_d N_VPWR_M1027_s
+ N_VPWR_c_1275_n N_VPWR_c_1276_n N_VPWR_c_1277_n N_VPWR_c_1278_n
+ N_VPWR_c_1279_n N_VPWR_c_1280_n N_VPWR_c_1281_n N_VPWR_c_1282_n
+ N_VPWR_c_1283_n N_VPWR_c_1284_n N_VPWR_c_1285_n VPWR N_VPWR_c_1286_n
+ N_VPWR_c_1287_n N_VPWR_c_1288_n N_VPWR_c_1289_n N_VPWR_c_1290_n
+ N_VPWR_c_1291_n N_VPWR_c_1274_n N_VPWR_c_1293_n N_VPWR_c_1294_n
+ N_VPWR_c_1295_n N_VPWR_c_1296_n N_VPWR_c_1297_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%VPWR
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_239_417# N_A_239_417#_M1036_s
+ N_A_239_417#_M1040_d N_A_239_417#_c_1407_n N_A_239_417#_c_1408_n
+ N_A_239_417#_c_1409_n N_A_239_417#_c_1410_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%A_239_417#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_343_417# N_A_343_417#_M1003_d
+ N_A_343_417#_M1041_d N_A_343_417#_M1036_d N_A_343_417#_M1010_s
+ N_A_343_417#_c_1454_n N_A_343_417#_c_1448_n N_A_343_417#_c_1456_n
+ N_A_343_417#_c_1449_n N_A_343_417#_c_1450_n N_A_343_417#_c_1451_n
+ N_A_343_417#_c_1452_n N_A_343_417#_c_1476_n N_A_343_417#_c_1457_n
+ N_A_343_417#_c_1453_n PM_SKY130_FD_SC_LP__SDFXBP_LP%A_343_417#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%Q N_Q_M1043_s N_Q_M1032_s N_Q_c_1552_n
+ N_Q_c_1553_n N_Q_c_1554_n Q Q N_Q_c_1556_n N_Q_c_1555_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%Q
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%Q_N N_Q_N_M1026_d N_Q_N_M1027_d N_Q_N_c_1587_n
+ Q_N Q_N Q_N PM_SKY130_FD_SC_LP__SDFXBP_LP%Q_N
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%VGND N_VGND_M1008_d N_VGND_M1012_d
+ N_VGND_M1021_d N_VGND_M1009_d N_VGND_M1001_d N_VGND_M1025_d N_VGND_M1031_s
+ N_VGND_c_1608_n N_VGND_c_1609_n N_VGND_c_1610_n N_VGND_c_1611_n
+ N_VGND_c_1612_n N_VGND_c_1613_n N_VGND_c_1614_n N_VGND_c_1615_n
+ N_VGND_c_1616_n N_VGND_c_1617_n VGND N_VGND_c_1618_n N_VGND_c_1619_n
+ N_VGND_c_1620_n N_VGND_c_1621_n N_VGND_c_1622_n N_VGND_c_1623_n
+ N_VGND_c_1624_n N_VGND_c_1625_n N_VGND_c_1626_n N_VGND_c_1627_n
+ N_VGND_c_1628_n N_VGND_c_1629_n N_VGND_c_1630_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%VGND
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1127_155# N_A_1127_155#_M1014_s
+ N_A_1127_155#_M1009_s N_A_1127_155#_c_1766_n N_A_1127_155#_c_1767_n
+ N_A_1127_155#_c_1768_n N_A_1127_155#_c_1769_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1127_155#
x_PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1859_155# N_A_1859_155#_M1042_s
+ N_A_1859_155#_M1001_s N_A_1859_155#_c_1800_n N_A_1859_155#_c_1801_n
+ N_A_1859_155#_c_1802_n N_A_1859_155#_c_1803_n
+ PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1859_155#
cc_1 VNB N_A_27_409#_c_259_n 0.0171345f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.165
cc_2 VNB N_A_27_409#_c_260_n 0.0230544f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.67
cc_3 VNB N_A_27_409#_c_261_n 0.031625f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.835
cc_4 VNB N_A_27_409#_c_262_n 0.0170869f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=2.19
cc_5 VNB N_A_27_409#_c_263_n 0.0251419f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.25
cc_6 VNB N_A_27_409#_c_264_n 0.0124808f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.25
cc_7 VNB N_A_27_409#_c_265_n 0.00486937f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_8 VNB N_A_27_409#_c_266_n 0.0148905f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_9 VNB N_D_M1003_g 0.0196163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_D_c_321_n 0.0172743f $X=-0.19 $Y=-0.245 $X2=1.61 $Y2=0.835
cc_11 VNB N_D_c_322_n 0.0155394f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.165
cc_12 VNB N_D_c_323_n 0.00729552f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.835
cc_13 VNB N_SCE_M1037_g 0.040928f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.96
cc_14 VNB N_SCE_M1008_g 0.0497964f $X=-0.19 $Y=-0.245 $X2=1.61 $Y2=0.835
cc_15 VNB N_SCE_c_363_n 0.115894f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_16 VNB N_SCE_c_364_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.165
cc_17 VNB N_SCE_M1020_g 0.0518047f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.835
cc_18 VNB N_SCE_c_366_n 0.00637503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_SCE_c_367_n 0.0218048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_SCD_M1012_g 0.0266427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_SCD_c_435_n 0.0298615f $X=-0.19 $Y=-0.245 $X2=1.61 $Y2=0.835
cc_22 VNB N_SCD_c_436_n 0.0250082f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.165
cc_23 VNB N_SCD_c_437_n 0.00310789f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.835
cc_24 VNB N_CLK_M1035_g 0.039376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_CLK_M1005_g 0.00416164f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.96
cc_26 VNB N_CLK_M1021_g 0.0298691f $X=-0.19 $Y=-0.245 $X2=1.61 $Y2=0.835
cc_27 VNB CLK 0.0125182f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.165
cc_28 VNB N_CLK_c_480_n 0.042149f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=2.9
cc_29 VNB N_A_1530_231#_M1007_g 0.00449428f $X=-0.19 $Y=-0.245 $X2=1.61
+ $Y2=0.835
cc_30 VNB N_A_1530_231#_c_518_n 0.00643702f $X=-0.19 $Y=-0.245 $X2=0.34
+ $Y2=0.835
cc_31 VNB N_A_1530_231#_c_519_n 8.91202e-19 $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=2.19
cc_32 VNB N_A_1530_231#_c_520_n 0.00312419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1530_231#_c_521_n 0.00488395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_1530_231#_c_522_n 0.0252031f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.25
cc_35 VNB N_A_1530_231#_c_523_n 0.00815663f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_36 VNB N_A_1530_231#_c_524_n 0.0270611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1530_231#_c_525_n 0.0165137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1278_155#_M1028_g 0.0195583f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.585
cc_39 VNB N_A_1278_155#_M1018_g 0.0184905f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.835
cc_40 VNB N_A_1278_155#_c_613_n 9.21676e-19 $X=-0.19 $Y=-0.245 $X2=0.225
+ $Y2=2.19
cc_41 VNB N_A_1278_155#_c_614_n 0.00673279f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.25
cc_42 VNB N_A_1278_155#_c_615_n 2.86565e-19 $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_43 VNB N_A_1278_155#_c_616_n 0.0310401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_706_66#_c_690_n 0.0155037f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.96
cc_45 VNB N_A_706_66#_M1030_g 0.00170344f $X=-0.19 $Y=-0.245 $X2=1.61 $Y2=0.835
cc_46 VNB N_A_706_66#_M1039_g 0.0101514f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.835
cc_47 VNB N_A_706_66#_c_693_n 0.113741f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.835
cc_48 VNB N_A_706_66#_c_694_n 0.0113293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_706_66#_M1041_g 0.0427494f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=2.19
cc_50 VNB N_A_706_66#_c_696_n 0.0202261f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=2.9
cc_51 VNB N_A_706_66#_c_697_n 0.0126912f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.25
cc_52 VNB N_A_706_66#_M1038_g 0.0115928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_706_66#_c_699_n 0.136318f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_54 VNB N_A_706_66#_c_700_n 0.0617025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_706_66#_M1024_g 0.0102955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_706_66#_c_702_n 0.014578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_706_66#_c_703_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_706_66#_c_704_n 0.0578274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_706_66#_c_705_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_706_66#_c_706_n 0.0369316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_706_66#_c_707_n 0.00795882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_706_66#_c_708_n 0.0199106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_706_66#_c_709_n 0.00504083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_706_66#_c_710_n 4.36532e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_706_66#_c_711_n 0.0675331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_975_347#_c_847_n 0.061175f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.585
cc_67 VNB N_A_975_347#_c_848_n 0.0163946f $X=-0.19 $Y=-0.245 $X2=1.61 $Y2=1.165
cc_68 VNB N_A_975_347#_c_849_n 0.0156413f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_69 VNB N_A_975_347#_M1033_g 0.00101233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_975_347#_M1022_g 0.0228161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_975_347#_c_852_n 0.012524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_975_347#_c_853_n 0.00558143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_975_347#_c_854_n 0.0105631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_975_347#_c_855_n 0.00507957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_975_347#_c_856_n 0.0140198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_2089_254#_c_949_n 0.0123891f $X=-0.19 $Y=-0.245 $X2=1.61 $Y2=0.835
cc_77 VNB N_A_2089_254#_c_950_n 0.0192196f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_78 VNB N_A_2089_254#_c_951_n 0.00968387f $X=-0.19 $Y=-0.245 $X2=1.52
+ $Y2=1.165
cc_79 VNB N_A_2089_254#_M1001_g 0.0301483f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.835
cc_80 VNB N_A_2089_254#_M1043_g 0.0318019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_2089_254#_M1025_g 0.0300914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_2089_254#_M1029_g 0.0301672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2089_254#_M1023_g 0.0341771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2089_254#_c_957_n 0.0013253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2089_254#_c_958_n 0.0144532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2089_254#_c_959_n 0.00341713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2089_254#_c_960_n 0.0103183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_2089_254#_c_961_n 0.0040442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2089_254#_c_962_n 0.0227961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2089_254#_c_963_n 0.00257414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2089_254#_c_964_n 0.00619014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2089_254#_c_965_n 0.001214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2089_254#_c_966_n 0.0186423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2089_254#_c_967_n 0.00171403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2089_254#_c_968_n 0.0356517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2089_254#_c_969_n 0.0568098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1902_347#_c_1119_n 0.0138266f $X=-0.19 $Y=-0.245 $X2=1.61
+ $Y2=0.835
cc_98 VNB N_A_1902_347#_c_1120_n 0.0241429f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.67
cc_99 VNB N_A_1902_347#_c_1121_n 0.0207919f $X=-0.19 $Y=-0.245 $X2=0.34
+ $Y2=1.165
cc_100 VNB N_A_1902_347#_c_1122_n 0.0173306f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=0.835
cc_101 VNB N_A_1902_347#_c_1123_n 0.00536562f $X=-0.19 $Y=-0.245 $X2=0.225
+ $Y2=2.19
cc_102 VNB N_A_1902_347#_c_1124_n 0.00386945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1902_347#_c_1125_n 0.00271625f $X=-0.19 $Y=-0.245 $X2=1.52
+ $Y2=1.33
cc_104 VNB N_A_1902_347#_c_1126_n 0.0354118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2714_401#_M1027_g 0.0059088f $X=-0.19 $Y=-0.245 $X2=1.59
+ $Y2=2.585
cc_106 VNB N_A_2714_401#_M1031_g 0.0238391f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_107 VNB N_A_2714_401#_c_1212_n 0.0302927f $X=-0.19 $Y=-0.245 $X2=1.52
+ $Y2=1.67
cc_108 VNB N_A_2714_401#_M1026_g 0.0249044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2714_401#_c_1214_n 0.025065f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.25
cc_110 VNB N_A_2714_401#_c_1215_n 0.00294153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2714_401#_c_1216_n 4.84214e-19 $X=-0.19 $Y=-0.245 $X2=0.34
+ $Y2=1.25
cc_112 VNB N_A_2714_401#_c_1217_n 0.00325948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2714_401#_c_1218_n 0.0894996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VPWR_c_1274_n 0.661241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_343_417#_c_1448_n 0.00969607f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=0.835
cc_116 VNB N_A_343_417#_c_1449_n 0.00713917f $X=-0.19 $Y=-0.245 $X2=0.225
+ $Y2=2.9
cc_117 VNB N_A_343_417#_c_1450_n 0.00278398f $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=2.9
cc_118 VNB N_A_343_417#_c_1451_n 0.00668443f $X=-0.19 $Y=-0.245 $X2=0.58
+ $Y2=1.25
cc_119 VNB N_A_343_417#_c_1452_n 0.00351648f $X=-0.19 $Y=-0.245 $X2=1.52
+ $Y2=1.33
cc_120 VNB N_A_343_417#_c_1453_n 0.00456775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_Q_c_1552_n 0.0185493f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.585
cc_122 VNB N_Q_c_1553_n 0.00402868f $X=-0.19 $Y=-0.245 $X2=1.61 $Y2=1.165
cc_123 VNB N_Q_c_1554_n 0.0094263f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_124 VNB N_Q_c_1555_n 0.00828106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_Q_N_c_1587_n 0.0689518f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.585
cc_126 VNB N_VGND_c_1608_n 0.0166303f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=2.9
cc_127 VNB N_VGND_c_1609_n 0.020796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1610_n 0.00293489f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_129 VNB N_VGND_c_1611_n 0.080284f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.33
cc_130 VNB N_VGND_c_1612_n 0.00881541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1613_n 0.00355527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1614_n 0.0230967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1615_n 0.0189585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1616_n 0.0452185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1617_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1618_n 0.0354332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1619_n 0.0434751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1620_n 0.0285659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1621_n 0.0763689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1622_n 0.0299115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1623_n 0.0267212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1624_n 0.822542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1625_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1626_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_1627_n 0.00555411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_1628_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_1629_n 0.00394875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_1630_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_A_1127_155#_c_1766_n 0.016681f $X=-0.19 $Y=-0.245 $X2=1.59
+ $Y2=2.585
cc_150 VNB N_A_1127_155#_c_1767_n 0.0311854f $X=-0.19 $Y=-0.245 $X2=1.61
+ $Y2=0.835
cc_151 VNB N_A_1127_155#_c_1768_n 0.00437116f $X=-0.19 $Y=-0.245 $X2=1.61
+ $Y2=0.835
cc_152 VNB N_A_1127_155#_c_1769_n 0.00720319f $X=-0.19 $Y=-0.245 $X2=1.52
+ $Y2=1.67
cc_153 VNB N_A_1859_155#_c_1800_n 0.00865773f $X=-0.19 $Y=-0.245 $X2=1.59
+ $Y2=2.585
cc_154 VNB N_A_1859_155#_c_1801_n 0.0148285f $X=-0.19 $Y=-0.245 $X2=1.61
+ $Y2=0.835
cc_155 VNB N_A_1859_155#_c_1802_n 0.00388015f $X=-0.19 $Y=-0.245 $X2=1.61
+ $Y2=0.835
cc_156 VNB N_A_1859_155#_c_1803_n 0.0110898f $X=-0.19 $Y=-0.245 $X2=1.52
+ $Y2=1.67
cc_157 VPB N_A_27_409#_c_267_n 0.0286324f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.96
cc_158 VPB N_A_27_409#_c_260_n 0.030407f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.67
cc_159 VPB N_A_27_409#_c_262_n 0.060749f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=2.19
cc_160 VPB N_A_27_409#_c_265_n 0.00114046f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.33
cc_161 VPB N_D_M1019_g 0.0274258f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.96
cc_162 VPB N_D_c_321_n 0.00403486f $X=-0.19 $Y=1.655 $X2=1.61 $Y2=0.835
cc_163 VPB N_D_c_326_n 0.0126013f $X=-0.19 $Y=1.655 $X2=1.61 $Y2=0.835
cc_164 VPB N_D_c_323_n 0.00237492f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=0.835
cc_165 VPB N_SCE_M1017_g 0.0391252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_SCE_c_366_n 0.00571439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_SCE_M1006_g 0.0329616f $X=-0.19 $Y=1.655 $X2=0.225 $Y2=2.19
cc_168 VPB SCE 0.00196975f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=2.9
cc_169 VPB N_SCE_c_367_n 0.0335097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_SCD_c_438_n 0.0160231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_SCD_M1040_g 0.032948f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.96
cc_172 VPB N_SCD_c_436_n 0.00910116f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.165
cc_173 VPB N_SCD_c_437_n 8.31394e-19 $X=-0.19 $Y=1.655 $X2=0.34 $Y2=0.835
cc_174 VPB N_CLK_M1005_g 0.033216f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.96
cc_175 VPB N_A_1530_231#_M1007_g 0.0248415f $X=-0.19 $Y=1.655 $X2=1.61 $Y2=0.835
cc_176 VPB N_A_1530_231#_c_520_n 0.00515973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_1278_155#_M1013_g 0.0257288f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.33
cc_178 VPB N_A_1278_155#_c_618_n 0.00264581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_1278_155#_c_619_n 0.0125306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_1278_155#_c_614_n 0.00526516f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.25
cc_181 VPB N_A_1278_155#_c_615_n 0.00104849f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.33
cc_182 VPB N_A_1278_155#_c_616_n 0.0105298f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_706_66#_M1030_g 0.0293033f $X=-0.19 $Y=1.655 $X2=1.61 $Y2=0.835
cc_184 VPB N_A_706_66#_M1038_g 0.0230911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_706_66#_M1024_g 0.0281744f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_706_66#_c_715_n 0.00680377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_706_66#_c_710_n 0.00289202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_975_347#_c_857_n 0.0848446f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=2.585
cc_189 VPB N_A_975_347#_c_858_n 0.0733613f $X=-0.19 $Y=1.655 $X2=1.61 $Y2=0.835
cc_190 VPB N_A_975_347#_c_859_n 0.012806f $X=-0.19 $Y=1.655 $X2=1.61 $Y2=0.835
cc_191 VPB N_A_975_347#_M1010_g 0.0525101f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.835
cc_192 VPB N_A_975_347#_c_861_n 0.250196f $X=-0.19 $Y=1.655 $X2=0.225 $Y2=1.335
cc_193 VPB N_A_975_347#_M1033_g 0.0414114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_975_347#_c_863_n 0.018623f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.33
cc_195 VPB N_A_975_347#_c_864_n 0.0124845f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.33
cc_196 VPB N_A_975_347#_c_865_n 0.008218f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_975_347#_c_854_n 0.00529233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_975_347#_c_855_n 0.0207885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_2089_254#_M1034_g 0.0274152f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=2.585
cc_200 VPB N_A_2089_254#_M1032_g 0.0332093f $X=-0.19 $Y=1.655 $X2=0.225 $Y2=2.19
cc_201 VPB N_A_2089_254#_M1011_g 0.0357371f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.33
cc_202 VPB N_A_2089_254#_c_957_n 0.00190329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_2089_254#_c_960_n 0.0127137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_2089_254#_c_965_n 0.00101054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_2089_254#_c_976_n 0.0110466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_2089_254#_c_977_n 0.0130119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_2089_254#_c_967_n 0.00142676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_2089_254#_c_968_n 0.00736443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_2089_254#_c_969_n 0.0591776f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_1902_347#_M1000_g 0.032209f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=2.585
cc_211 VPB N_A_1902_347#_c_1128_n 0.00354194f $X=-0.19 $Y=1.655 $X2=0.265
+ $Y2=2.9
cc_212 VPB N_A_1902_347#_c_1124_n 0.00235803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_1902_347#_c_1130_n 0.00147494f $X=-0.19 $Y=1.655 $X2=0.34
+ $Y2=1.25
cc_214 VPB N_A_1902_347#_c_1125_n 0.00126953f $X=-0.19 $Y=1.655 $X2=1.52
+ $Y2=1.33
cc_215 VPB N_A_1902_347#_c_1132_n 0.00393493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_1902_347#_c_1126_n 0.0148428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_2714_401#_M1027_g 0.0517939f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=2.585
cc_218 VPB N_A_2714_401#_c_1220_n 0.00211757f $X=-0.19 $Y=1.655 $X2=0.225
+ $Y2=2.19
cc_219 VPB N_A_2714_401#_c_1221_n 0.0123719f $X=-0.19 $Y=1.655 $X2=0.225 $Y2=2.9
cc_220 VPB N_A_2714_401#_c_1222_n 0.0210243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_2714_401#_c_1216_n 0.00709691f $X=-0.19 $Y=1.655 $X2=0.34
+ $Y2=1.25
cc_222 VPB N_VPWR_c_1275_n 0.0162937f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=2.9
cc_223 VPB N_VPWR_c_1276_n 7.46595e-19 $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.25
cc_224 VPB N_VPWR_c_1277_n 0.0229058f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.33
cc_225 VPB N_VPWR_c_1278_n 0.0183667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1279_n 0.020364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1280_n 0.00515606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1281_n 0.0119679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1282_n 0.0458493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1283_n 0.0044842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1284_n 0.0234142f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1285_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1286_n 0.0191856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1287_n 0.0364355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1288_n 0.0967214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1289_n 0.0765034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1290_n 0.0531282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1291_n 0.034152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1274_n 0.188888f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1293_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1294_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1295_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1296_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1297_n 0.00546719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_239_417#_c_1407_n 0.0126786f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=2.585
cc_246 VPB N_A_239_417#_c_1408_n 0.00299582f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.33
cc_247 VPB N_A_239_417#_c_1409_n 0.0106052f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=0.835
cc_248 VPB N_A_239_417#_c_1410_n 0.00525261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_343_417#_c_1454_n 0.0148191f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.33
cc_250 VPB N_A_343_417#_c_1448_n 0.0031944f $X=-0.19 $Y=1.655 $X2=0.415
+ $Y2=0.835
cc_251 VPB N_A_343_417#_c_1456_n 0.0575745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_343_417#_c_1457_n 0.0296642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_343_417#_c_1453_n 0.0046872f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_Q_c_1556_n 0.0480818f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=2.9
cc_255 VPB N_Q_c_1555_n 0.0085848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_Q_N_c_1587_n 0.0172849f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=2.585
cc_257 VPB Q_N 0.102509f $X=-0.19 $Y=1.655 $X2=1.61 $Y2=0.835
cc_258 N_A_27_409#_c_259_n N_D_M1003_g 0.0233528f $X=1.52 $Y=1.165 $X2=0 $Y2=0
cc_259 N_A_27_409#_c_265_n N_D_M1003_g 7.58678e-19 $X=1.52 $Y=1.33 $X2=0 $Y2=0
cc_260 N_A_27_409#_c_260_n N_D_M1019_g 0.0495707f $X=1.52 $Y=1.67 $X2=0 $Y2=0
cc_261 N_A_27_409#_c_260_n N_D_c_321_n 0.0233528f $X=1.52 $Y=1.67 $X2=0 $Y2=0
cc_262 N_A_27_409#_c_260_n N_D_c_326_n 0.00331853f $X=1.52 $Y=1.67 $X2=0 $Y2=0
cc_263 N_A_27_409#_c_265_n N_D_c_322_n 0.00183338f $X=1.52 $Y=1.33 $X2=0 $Y2=0
cc_264 N_A_27_409#_c_266_n N_D_c_322_n 0.0233528f $X=1.52 $Y=1.33 $X2=0 $Y2=0
cc_265 N_A_27_409#_c_260_n N_D_c_323_n 0.00218366f $X=1.52 $Y=1.67 $X2=0 $Y2=0
cc_266 N_A_27_409#_c_265_n N_D_c_323_n 0.0357605f $X=1.52 $Y=1.33 $X2=0 $Y2=0
cc_267 N_A_27_409#_c_261_n N_SCE_M1037_g 0.0142128f $X=0.415 $Y=0.835 $X2=0
+ $Y2=0
cc_268 N_A_27_409#_c_262_n N_SCE_M1037_g 0.00617929f $X=0.265 $Y=2.19 $X2=0
+ $Y2=0
cc_269 N_A_27_409#_c_263_n N_SCE_M1037_g 0.0107743f $X=1.355 $Y=1.25 $X2=0 $Y2=0
cc_270 N_A_27_409#_c_264_n N_SCE_M1037_g 0.00452984f $X=0.34 $Y=1.25 $X2=0 $Y2=0
cc_271 N_A_27_409#_c_259_n N_SCE_M1008_g 0.0146973f $X=1.52 $Y=1.165 $X2=0 $Y2=0
cc_272 N_A_27_409#_c_261_n N_SCE_M1008_g 0.00199825f $X=0.415 $Y=0.835 $X2=0
+ $Y2=0
cc_273 N_A_27_409#_c_263_n N_SCE_M1008_g 0.0186426f $X=1.355 $Y=1.25 $X2=0 $Y2=0
cc_274 N_A_27_409#_c_265_n N_SCE_M1008_g 0.00187033f $X=1.52 $Y=1.33 $X2=0 $Y2=0
cc_275 N_A_27_409#_c_266_n N_SCE_M1008_g 0.0127446f $X=1.52 $Y=1.33 $X2=0 $Y2=0
cc_276 N_A_27_409#_c_259_n N_SCE_c_363_n 0.00907339f $X=1.52 $Y=1.165 $X2=0
+ $Y2=0
cc_277 N_A_27_409#_c_260_n SCE 0.00116801f $X=1.52 $Y=1.67 $X2=0 $Y2=0
cc_278 N_A_27_409#_c_262_n SCE 0.024436f $X=0.265 $Y=2.19 $X2=0 $Y2=0
cc_279 N_A_27_409#_c_263_n SCE 0.0196541f $X=1.355 $Y=1.25 $X2=0 $Y2=0
cc_280 N_A_27_409#_c_264_n SCE 0.0039252f $X=0.34 $Y=1.25 $X2=0 $Y2=0
cc_281 N_A_27_409#_c_265_n SCE 0.0100245f $X=1.52 $Y=1.33 $X2=0 $Y2=0
cc_282 N_A_27_409#_c_260_n N_SCE_c_367_n 0.0164041f $X=1.52 $Y=1.67 $X2=0 $Y2=0
cc_283 N_A_27_409#_c_262_n N_SCE_c_367_n 0.0183587f $X=0.265 $Y=2.19 $X2=0 $Y2=0
cc_284 N_A_27_409#_c_263_n N_SCE_c_367_n 0.00133659f $X=1.355 $Y=1.25 $X2=0
+ $Y2=0
cc_285 N_A_27_409#_c_264_n N_SCE_c_367_n 0.00666029f $X=0.34 $Y=1.25 $X2=0 $Y2=0
cc_286 N_A_27_409#_c_267_n N_VPWR_c_1275_n 0.00579437f $X=1.59 $Y=1.96 $X2=0
+ $Y2=0
cc_287 N_A_27_409#_c_262_n N_VPWR_c_1275_n 0.0272606f $X=0.265 $Y=2.19 $X2=0
+ $Y2=0
cc_288 N_A_27_409#_c_267_n N_VPWR_c_1282_n 0.00689754f $X=1.59 $Y=1.96 $X2=0
+ $Y2=0
cc_289 N_A_27_409#_c_262_n N_VPWR_c_1286_n 0.0167213f $X=0.265 $Y=2.19 $X2=0
+ $Y2=0
cc_290 N_A_27_409#_c_267_n N_VPWR_c_1274_n 0.0101052f $X=1.59 $Y=1.96 $X2=0
+ $Y2=0
cc_291 N_A_27_409#_c_262_n N_VPWR_c_1274_n 0.0095959f $X=0.265 $Y=2.19 $X2=0
+ $Y2=0
cc_292 N_A_27_409#_c_267_n N_A_239_417#_c_1407_n 0.0103575f $X=1.59 $Y=1.96
+ $X2=0 $Y2=0
cc_293 N_A_27_409#_c_260_n N_A_239_417#_c_1407_n 8.23522e-19 $X=1.52 $Y=1.67
+ $X2=0 $Y2=0
cc_294 N_A_27_409#_c_265_n N_A_239_417#_c_1407_n 0.00931822f $X=1.52 $Y=1.33
+ $X2=0 $Y2=0
cc_295 N_A_27_409#_c_267_n N_A_239_417#_c_1408_n 0.0168883f $X=1.59 $Y=1.96
+ $X2=0 $Y2=0
cc_296 N_A_27_409#_c_265_n N_A_239_417#_c_1408_n 0.00466377f $X=1.52 $Y=1.33
+ $X2=0 $Y2=0
cc_297 N_A_27_409#_c_267_n N_A_239_417#_c_1410_n 0.0125111f $X=1.59 $Y=1.96
+ $X2=0 $Y2=0
cc_298 N_A_27_409#_c_267_n N_A_343_417#_c_1454_n 0.00624708f $X=1.59 $Y=1.96
+ $X2=0 $Y2=0
cc_299 N_A_27_409#_c_259_n N_VGND_c_1608_n 0.00598409f $X=1.52 $Y=1.165 $X2=0
+ $Y2=0
cc_300 N_A_27_409#_c_261_n N_VGND_c_1608_n 0.00590801f $X=0.415 $Y=0.835 $X2=0
+ $Y2=0
cc_301 N_A_27_409#_c_263_n N_VGND_c_1608_n 0.0160998f $X=1.355 $Y=1.25 $X2=0
+ $Y2=0
cc_302 N_A_27_409#_c_265_n N_VGND_c_1608_n 0.0103105f $X=1.52 $Y=1.33 $X2=0
+ $Y2=0
cc_303 N_A_27_409#_c_266_n N_VGND_c_1608_n 9.60587e-19 $X=1.52 $Y=1.33 $X2=0
+ $Y2=0
cc_304 N_A_27_409#_c_261_n N_VGND_c_1618_n 0.0102582f $X=0.415 $Y=0.835 $X2=0
+ $Y2=0
cc_305 N_A_27_409#_c_259_n N_VGND_c_1624_n 9.49986e-19 $X=1.52 $Y=1.165 $X2=0
+ $Y2=0
cc_306 N_A_27_409#_c_261_n N_VGND_c_1624_n 0.0148003f $X=0.415 $Y=0.835 $X2=0
+ $Y2=0
cc_307 N_D_M1003_g N_SCE_c_363_n 0.00907339f $X=2 $Y=0.835 $X2=0 $Y2=0
cc_308 N_D_M1003_g N_SCE_M1020_g 0.0141983f $X=2 $Y=0.835 $X2=0 $Y2=0
cc_309 N_D_c_322_n N_SCE_M1020_g 0.0144038f $X=2.09 $Y=1.38 $X2=0 $Y2=0
cc_310 N_D_c_323_n N_SCE_M1020_g 0.00222056f $X=2.09 $Y=1.38 $X2=0 $Y2=0
cc_311 N_D_c_321_n N_SCE_c_366_n 0.0144038f $X=2.09 $Y=1.72 $X2=0 $Y2=0
cc_312 N_D_M1019_g N_SCE_M1006_g 0.0847292f $X=2.12 $Y=2.585 $X2=0 $Y2=0
cc_313 N_D_c_326_n N_SCE_M1006_g 0.0144038f $X=2.09 $Y=1.885 $X2=0 $Y2=0
cc_314 N_D_M1019_g N_VPWR_c_1276_n 0.00189839f $X=2.12 $Y=2.585 $X2=0 $Y2=0
cc_315 N_D_M1019_g N_VPWR_c_1282_n 0.00699368f $X=2.12 $Y=2.585 $X2=0 $Y2=0
cc_316 N_D_M1019_g N_VPWR_c_1274_n 0.00878302f $X=2.12 $Y=2.585 $X2=0 $Y2=0
cc_317 N_D_M1019_g N_A_239_417#_c_1407_n 6.31982e-19 $X=2.12 $Y=2.585 $X2=0
+ $Y2=0
cc_318 N_D_M1019_g N_A_239_417#_c_1408_n 0.0168827f $X=2.12 $Y=2.585 $X2=0 $Y2=0
cc_319 N_D_M1019_g N_A_239_417#_c_1410_n 0.00167569f $X=2.12 $Y=2.585 $X2=0
+ $Y2=0
cc_320 N_D_M1019_g N_A_343_417#_c_1454_n 0.0158567f $X=2.12 $Y=2.585 $X2=0 $Y2=0
cc_321 N_D_c_326_n N_A_343_417#_c_1454_n 5.6123e-19 $X=2.09 $Y=1.885 $X2=0 $Y2=0
cc_322 N_D_c_323_n N_A_343_417#_c_1454_n 0.026525f $X=2.09 $Y=1.38 $X2=0 $Y2=0
cc_323 N_D_M1003_g N_A_343_417#_c_1448_n 0.00288917f $X=2 $Y=0.835 $X2=0 $Y2=0
cc_324 N_D_M1019_g N_A_343_417#_c_1448_n 0.00347224f $X=2.12 $Y=2.585 $X2=0
+ $Y2=0
cc_325 N_D_c_322_n N_A_343_417#_c_1448_n 0.00189779f $X=2.09 $Y=1.38 $X2=0 $Y2=0
cc_326 N_D_c_323_n N_A_343_417#_c_1448_n 0.0512418f $X=2.09 $Y=1.38 $X2=0 $Y2=0
cc_327 N_D_M1003_g N_A_343_417#_c_1452_n 0.0125397f $X=2 $Y=0.835 $X2=0 $Y2=0
cc_328 N_D_c_322_n N_A_343_417#_c_1452_n 7.03802e-19 $X=2.09 $Y=1.38 $X2=0 $Y2=0
cc_329 N_D_c_323_n N_A_343_417#_c_1452_n 0.00923904f $X=2.09 $Y=1.38 $X2=0 $Y2=0
cc_330 N_D_M1003_g N_VGND_c_1624_n 9.49986e-19 $X=2 $Y=0.835 $X2=0 $Y2=0
cc_331 N_SCE_M1020_g N_SCD_M1012_g 0.0541821f $X=2.54 $Y=0.835 $X2=0 $Y2=0
cc_332 N_SCE_M1006_g N_SCD_c_438_n 0.00721431f $X=2.59 $Y=2.585 $X2=0 $Y2=0
cc_333 N_SCE_M1006_g N_SCD_M1040_g 0.0464232f $X=2.59 $Y=2.585 $X2=0 $Y2=0
cc_334 N_SCE_M1020_g N_SCD_c_436_n 0.00818216f $X=2.54 $Y=0.835 $X2=0 $Y2=0
cc_335 N_SCE_c_366_n N_SCD_c_436_n 0.00721431f $X=2.59 $Y=1.76 $X2=0 $Y2=0
cc_336 N_SCE_M1020_g N_SCD_c_437_n 4.59768e-19 $X=2.54 $Y=0.835 $X2=0 $Y2=0
cc_337 N_SCE_c_366_n N_SCD_c_437_n 0.0010341f $X=2.59 $Y=1.76 $X2=0 $Y2=0
cc_338 N_SCE_M1017_g N_VPWR_c_1275_n 0.0231789f $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_339 SCE N_VPWR_c_1275_n 0.0183894f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_340 N_SCE_c_367_n N_VPWR_c_1275_n 0.00923211f $X=0.695 $Y=1.68 $X2=0 $Y2=0
cc_341 N_SCE_M1006_g N_VPWR_c_1276_n 0.00974128f $X=2.59 $Y=2.585 $X2=0 $Y2=0
cc_342 N_SCE_M1006_g N_VPWR_c_1282_n 0.00628722f $X=2.59 $Y=2.585 $X2=0 $Y2=0
cc_343 N_SCE_M1017_g N_VPWR_c_1286_n 0.00802402f $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_344 N_SCE_M1017_g N_VPWR_c_1274_n 0.0149648f $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_345 N_SCE_M1006_g N_VPWR_c_1274_n 0.00697167f $X=2.59 $Y=2.585 $X2=0 $Y2=0
cc_346 N_SCE_M1006_g N_A_239_417#_c_1408_n 0.0166118f $X=2.59 $Y=2.585 $X2=0
+ $Y2=0
cc_347 N_SCE_M1006_g N_A_239_417#_c_1409_n 5.47451e-19 $X=2.59 $Y=2.585 $X2=0
+ $Y2=0
cc_348 N_SCE_M1017_g N_A_239_417#_c_1410_n 6.6939e-19 $X=0.53 $Y=2.545 $X2=0
+ $Y2=0
cc_349 N_SCE_M1020_g N_A_343_417#_c_1448_n 0.0120665f $X=2.54 $Y=0.835 $X2=0
+ $Y2=0
cc_350 N_SCE_c_366_n N_A_343_417#_c_1448_n 0.00356178f $X=2.59 $Y=1.76 $X2=0
+ $Y2=0
cc_351 N_SCE_M1006_g N_A_343_417#_c_1448_n 0.00874271f $X=2.59 $Y=2.585 $X2=0
+ $Y2=0
cc_352 N_SCE_M1006_g N_A_343_417#_c_1456_n 0.0083692f $X=2.59 $Y=2.585 $X2=0
+ $Y2=0
cc_353 N_SCE_c_363_n N_A_343_417#_c_1452_n 0.00412283f $X=2.465 $Y=0.18 $X2=0
+ $Y2=0
cc_354 N_SCE_M1020_g N_A_343_417#_c_1452_n 0.0108615f $X=2.54 $Y=0.835 $X2=0
+ $Y2=0
cc_355 N_SCE_M1006_g N_A_343_417#_c_1476_n 0.010259f $X=2.59 $Y=2.585 $X2=0
+ $Y2=0
cc_356 N_SCE_M1008_g N_VGND_c_1608_n 0.0157955f $X=1.02 $Y=0.835 $X2=0 $Y2=0
cc_357 N_SCE_c_363_n N_VGND_c_1608_n 0.0248025f $X=2.465 $Y=0.18 $X2=0 $Y2=0
cc_358 N_SCE_c_363_n N_VGND_c_1609_n 0.011085f $X=2.465 $Y=0.18 $X2=0 $Y2=0
cc_359 N_SCE_M1020_g N_VGND_c_1609_n 0.0010356f $X=2.54 $Y=0.835 $X2=0 $Y2=0
cc_360 N_SCE_M1037_g N_VGND_c_1618_n 0.00399929f $X=0.63 $Y=0.835 $X2=0 $Y2=0
cc_361 N_SCE_c_364_n N_VGND_c_1618_n 0.00796123f $X=1.095 $Y=0.18 $X2=0 $Y2=0
cc_362 N_SCE_c_363_n N_VGND_c_1619_n 0.0359211f $X=2.465 $Y=0.18 $X2=0 $Y2=0
cc_363 N_SCE_M1037_g N_VGND_c_1624_n 0.00469432f $X=0.63 $Y=0.835 $X2=0 $Y2=0
cc_364 N_SCE_c_363_n N_VGND_c_1624_n 0.0483377f $X=2.465 $Y=0.18 $X2=0 $Y2=0
cc_365 N_SCE_c_364_n N_VGND_c_1624_n 0.0114838f $X=1.095 $Y=0.18 $X2=0 $Y2=0
cc_366 N_SCD_M1012_g CLK 0.00182718f $X=2.9 $Y=0.835 $X2=0 $Y2=0
cc_367 N_SCD_c_435_n CLK 0.00261831f $X=3.055 $Y=1.395 $X2=0 $Y2=0
cc_368 N_SCD_c_437_n CLK 0.0197462f $X=3.12 $Y=1.41 $X2=0 $Y2=0
cc_369 N_SCD_c_435_n N_CLK_c_480_n 0.00477175f $X=3.055 $Y=1.395 $X2=0 $Y2=0
cc_370 N_SCD_c_437_n N_CLK_c_480_n 2.17668e-19 $X=3.12 $Y=1.41 $X2=0 $Y2=0
cc_371 N_SCD_M1012_g N_A_706_66#_c_707_n 8.7948e-19 $X=2.9 $Y=0.835 $X2=0 $Y2=0
cc_372 N_SCD_M1040_g N_A_706_66#_c_715_n 0.00171015f $X=3.12 $Y=2.585 $X2=0
+ $Y2=0
cc_373 N_SCD_c_436_n N_A_706_66#_c_715_n 0.00370034f $X=3.12 $Y=1.41 $X2=0 $Y2=0
cc_374 N_SCD_c_437_n N_A_706_66#_c_715_n 0.00741569f $X=3.12 $Y=1.41 $X2=0 $Y2=0
cc_375 N_SCD_M1040_g N_VPWR_c_1276_n 0.0098582f $X=3.12 $Y=2.585 $X2=0 $Y2=0
cc_376 N_SCD_M1040_g N_VPWR_c_1287_n 0.00619108f $X=3.12 $Y=2.585 $X2=0 $Y2=0
cc_377 N_SCD_M1040_g N_VPWR_c_1274_n 0.00830296f $X=3.12 $Y=2.585 $X2=0 $Y2=0
cc_378 N_SCD_M1040_g N_A_239_417#_c_1408_n 0.0161244f $X=3.12 $Y=2.585 $X2=0
+ $Y2=0
cc_379 N_SCD_M1040_g N_A_239_417#_c_1409_n 0.00908033f $X=3.12 $Y=2.585 $X2=0
+ $Y2=0
cc_380 N_SCD_M1012_g N_A_343_417#_c_1448_n 0.00463317f $X=2.9 $Y=0.835 $X2=0
+ $Y2=0
cc_381 N_SCD_M1040_g N_A_343_417#_c_1448_n 8.26219e-19 $X=3.12 $Y=2.585 $X2=0
+ $Y2=0
cc_382 N_SCD_c_436_n N_A_343_417#_c_1448_n 0.00244943f $X=3.12 $Y=1.41 $X2=0
+ $Y2=0
cc_383 N_SCD_c_437_n N_A_343_417#_c_1448_n 0.0295579f $X=3.12 $Y=1.41 $X2=0
+ $Y2=0
cc_384 N_SCD_M1040_g N_A_343_417#_c_1456_n 0.0176591f $X=3.12 $Y=2.585 $X2=0
+ $Y2=0
cc_385 N_SCD_c_437_n N_A_343_417#_c_1456_n 0.0169044f $X=3.12 $Y=1.41 $X2=0
+ $Y2=0
cc_386 N_SCD_M1012_g N_A_343_417#_c_1452_n 0.00112422f $X=2.9 $Y=0.835 $X2=0
+ $Y2=0
cc_387 N_SCD_M1040_g N_A_343_417#_c_1476_n 4.90465e-19 $X=3.12 $Y=2.585 $X2=0
+ $Y2=0
cc_388 N_SCD_M1012_g N_VGND_c_1609_n 0.0127779f $X=2.9 $Y=0.835 $X2=0 $Y2=0
cc_389 N_SCD_c_435_n N_VGND_c_1609_n 0.00236087f $X=3.055 $Y=1.395 $X2=0 $Y2=0
cc_390 N_SCD_c_437_n N_VGND_c_1609_n 0.0274564f $X=3.12 $Y=1.41 $X2=0 $Y2=0
cc_391 N_SCD_M1012_g N_VGND_c_1619_n 0.00345209f $X=2.9 $Y=0.835 $X2=0 $Y2=0
cc_392 N_SCD_M1012_g N_VGND_c_1624_n 0.00394323f $X=2.9 $Y=0.835 $X2=0 $Y2=0
cc_393 N_CLK_M1021_g N_A_706_66#_c_690_n 0.0286345f $X=4.23 $Y=0.54 $X2=0 $Y2=0
cc_394 N_CLK_M1005_g N_A_706_66#_M1030_g 0.0451124f $X=4.22 $Y=2.235 $X2=0 $Y2=0
cc_395 N_CLK_M1035_g N_A_706_66#_c_707_n 0.0113373f $X=3.87 $Y=0.54 $X2=0 $Y2=0
cc_396 N_CLK_M1021_g N_A_706_66#_c_707_n 0.0018251f $X=4.23 $Y=0.54 $X2=0 $Y2=0
cc_397 N_CLK_M1005_g N_A_706_66#_c_715_n 0.0206107f $X=4.22 $Y=2.235 $X2=0 $Y2=0
cc_398 CLK N_A_706_66#_c_715_n 0.0269535f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_399 N_CLK_c_480_n N_A_706_66#_c_715_n 0.00767252f $X=4.23 $Y=1.345 $X2=0
+ $Y2=0
cc_400 N_CLK_M1035_g N_A_706_66#_c_708_n 0.00806747f $X=3.87 $Y=0.54 $X2=0 $Y2=0
cc_401 N_CLK_M1021_g N_A_706_66#_c_708_n 0.0189993f $X=4.23 $Y=0.54 $X2=0 $Y2=0
cc_402 CLK N_A_706_66#_c_708_n 0.0537786f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_403 N_CLK_c_480_n N_A_706_66#_c_708_n 0.00646481f $X=4.23 $Y=1.345 $X2=0
+ $Y2=0
cc_404 N_CLK_M1035_g N_A_706_66#_c_709_n 0.00419338f $X=3.87 $Y=0.54 $X2=0 $Y2=0
cc_405 CLK N_A_706_66#_c_709_n 0.0278467f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_406 N_CLK_M1005_g N_A_706_66#_c_710_n 0.00415409f $X=4.22 $Y=2.235 $X2=0
+ $Y2=0
cc_407 CLK N_A_706_66#_c_711_n 2.30698e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_408 N_CLK_c_480_n N_A_706_66#_c_711_n 0.0188053f $X=4.23 $Y=1.345 $X2=0 $Y2=0
cc_409 N_CLK_M1005_g N_VPWR_c_1277_n 0.0184641f $X=4.22 $Y=2.235 $X2=0 $Y2=0
cc_410 N_CLK_M1005_g N_VPWR_c_1287_n 0.00646289f $X=4.22 $Y=2.235 $X2=0 $Y2=0
cc_411 N_CLK_M1005_g N_VPWR_c_1274_n 0.00719887f $X=4.22 $Y=2.235 $X2=0 $Y2=0
cc_412 N_CLK_M1005_g N_A_239_417#_c_1408_n 0.00496458f $X=4.22 $Y=2.235 $X2=0
+ $Y2=0
cc_413 N_CLK_M1005_g N_A_239_417#_c_1409_n 0.00501972f $X=4.22 $Y=2.235 $X2=0
+ $Y2=0
cc_414 N_CLK_M1005_g N_A_343_417#_c_1456_n 0.0234019f $X=4.22 $Y=2.235 $X2=0
+ $Y2=0
cc_415 CLK N_A_343_417#_c_1456_n 0.0094748f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_416 N_CLK_M1035_g N_VGND_c_1609_n 0.00587929f $X=3.87 $Y=0.54 $X2=0 $Y2=0
cc_417 N_CLK_M1035_g N_VGND_c_1610_n 0.00163126f $X=3.87 $Y=0.54 $X2=0 $Y2=0
cc_418 N_CLK_M1021_g N_VGND_c_1610_n 0.00983975f $X=4.23 $Y=0.54 $X2=0 $Y2=0
cc_419 N_CLK_M1035_g N_VGND_c_1620_n 0.0046526f $X=3.87 $Y=0.54 $X2=0 $Y2=0
cc_420 N_CLK_M1021_g N_VGND_c_1620_n 0.00411131f $X=4.23 $Y=0.54 $X2=0 $Y2=0
cc_421 N_CLK_M1035_g N_VGND_c_1624_n 0.00553875f $X=3.87 $Y=0.54 $X2=0 $Y2=0
cc_422 N_CLK_M1021_g N_VGND_c_1624_n 0.00401821f $X=4.23 $Y=0.54 $X2=0 $Y2=0
cc_423 N_A_1530_231#_c_518_n N_A_1278_155#_M1028_g 0.011542f $X=8.705 $Y=0.98
+ $X2=0 $Y2=0
cc_424 N_A_1530_231#_c_519_n N_A_1278_155#_M1028_g 0.001518f $X=8.87 $Y=0.835
+ $X2=0 $Y2=0
cc_425 N_A_1530_231#_c_523_n N_A_1278_155#_M1028_g 0.0033783f $X=7.815 $Y=0.98
+ $X2=0 $Y2=0
cc_426 N_A_1530_231#_c_524_n N_A_1278_155#_M1028_g 0.0178275f $X=7.815 $Y=1.32
+ $X2=0 $Y2=0
cc_427 N_A_1530_231#_c_525_n N_A_1278_155#_M1028_g 0.0166686f $X=7.815 $Y=1.155
+ $X2=0 $Y2=0
cc_428 N_A_1530_231#_M1007_g N_A_1278_155#_M1013_g 0.0139706f $X=7.775 $Y=2.235
+ $X2=0 $Y2=0
cc_429 N_A_1530_231#_c_520_n N_A_1278_155#_M1013_g 0.0315506f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_430 N_A_1530_231#_c_518_n N_A_1278_155#_M1018_g 0.0113997f $X=8.705 $Y=0.98
+ $X2=0 $Y2=0
cc_431 N_A_1530_231#_c_519_n N_A_1278_155#_M1018_g 0.00905777f $X=8.87 $Y=0.835
+ $X2=0 $Y2=0
cc_432 N_A_1530_231#_c_520_n N_A_1278_155#_M1018_g 0.00525241f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_433 N_A_1530_231#_c_538_p N_A_1278_155#_M1018_g 0.00211036f $X=8.89 $Y=0.98
+ $X2=0 $Y2=0
cc_434 N_A_1530_231#_M1007_g N_A_1278_155#_c_618_n 0.00397468f $X=7.775 $Y=2.235
+ $X2=0 $Y2=0
cc_435 N_A_1530_231#_M1007_g N_A_1278_155#_c_619_n 0.022849f $X=7.775 $Y=2.235
+ $X2=0 $Y2=0
cc_436 N_A_1530_231#_c_518_n N_A_1278_155#_c_619_n 0.007489f $X=8.705 $Y=0.98
+ $X2=0 $Y2=0
cc_437 N_A_1530_231#_c_520_n N_A_1278_155#_c_619_n 0.0121506f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_438 N_A_1530_231#_c_523_n N_A_1278_155#_c_619_n 0.0234901f $X=7.815 $Y=0.98
+ $X2=0 $Y2=0
cc_439 N_A_1530_231#_c_524_n N_A_1278_155#_c_619_n 5.56982e-19 $X=7.815 $Y=1.32
+ $X2=0 $Y2=0
cc_440 N_A_1530_231#_M1007_g N_A_1278_155#_c_614_n 7.73787e-19 $X=7.775 $Y=2.235
+ $X2=0 $Y2=0
cc_441 N_A_1530_231#_c_523_n N_A_1278_155#_c_614_n 0.00315266f $X=7.815 $Y=0.98
+ $X2=0 $Y2=0
cc_442 N_A_1530_231#_M1007_g N_A_1278_155#_c_615_n 0.00261188f $X=7.775 $Y=2.235
+ $X2=0 $Y2=0
cc_443 N_A_1530_231#_c_518_n N_A_1278_155#_c_615_n 0.0242553f $X=8.705 $Y=0.98
+ $X2=0 $Y2=0
cc_444 N_A_1530_231#_c_520_n N_A_1278_155#_c_615_n 0.0281386f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_445 N_A_1530_231#_c_523_n N_A_1278_155#_c_615_n 0.0137249f $X=7.815 $Y=0.98
+ $X2=0 $Y2=0
cc_446 N_A_1530_231#_c_524_n N_A_1278_155#_c_615_n 3.0694e-19 $X=7.815 $Y=1.32
+ $X2=0 $Y2=0
cc_447 N_A_1530_231#_M1007_g N_A_1278_155#_c_616_n 0.00401762f $X=7.775 $Y=2.235
+ $X2=0 $Y2=0
cc_448 N_A_1530_231#_c_518_n N_A_1278_155#_c_616_n 2.08868e-19 $X=8.705 $Y=0.98
+ $X2=0 $Y2=0
cc_449 N_A_1530_231#_c_520_n N_A_1278_155#_c_616_n 0.0107888f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_450 N_A_1530_231#_c_538_p N_A_1278_155#_c_616_n 7.17987e-19 $X=8.89 $Y=0.98
+ $X2=0 $Y2=0
cc_451 N_A_1530_231#_c_523_n N_A_706_66#_c_697_n 0.00120856f $X=7.815 $Y=0.98
+ $X2=0 $Y2=0
cc_452 N_A_1530_231#_c_524_n N_A_706_66#_c_697_n 0.0442265f $X=7.815 $Y=1.32
+ $X2=0 $Y2=0
cc_453 N_A_1530_231#_M1007_g N_A_706_66#_M1038_g 0.0442265f $X=7.775 $Y=2.235
+ $X2=0 $Y2=0
cc_454 N_A_1530_231#_c_518_n N_A_706_66#_c_699_n 0.00460578f $X=8.705 $Y=0.98
+ $X2=0 $Y2=0
cc_455 N_A_1530_231#_c_521_n N_A_706_66#_c_699_n 0.00637147f $X=9.075 $Y=0.35
+ $X2=0 $Y2=0
cc_456 N_A_1530_231#_c_523_n N_A_706_66#_c_699_n 3.87137e-19 $X=7.815 $Y=0.98
+ $X2=0 $Y2=0
cc_457 N_A_1530_231#_c_525_n N_A_706_66#_c_699_n 0.00907339f $X=7.815 $Y=1.155
+ $X2=0 $Y2=0
cc_458 N_A_1530_231#_c_519_n N_A_706_66#_c_700_n 0.0168164f $X=8.87 $Y=0.835
+ $X2=0 $Y2=0
cc_459 N_A_1530_231#_c_520_n N_A_706_66#_c_700_n 0.00483785f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_460 N_A_1530_231#_c_521_n N_A_706_66#_c_700_n 0.00370441f $X=9.075 $Y=0.35
+ $X2=0 $Y2=0
cc_461 N_A_1530_231#_c_522_n N_A_706_66#_c_700_n 0.0139997f $X=10.41 $Y=0.35
+ $X2=0 $Y2=0
cc_462 N_A_1530_231#_c_538_p N_A_706_66#_c_700_n 0.00388024f $X=8.89 $Y=0.98
+ $X2=0 $Y2=0
cc_463 N_A_1530_231#_c_520_n N_A_706_66#_M1024_g 0.0168469f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_464 N_A_1530_231#_c_522_n N_A_706_66#_c_702_n 9.5131e-19 $X=10.41 $Y=0.35
+ $X2=0 $Y2=0
cc_465 N_A_1530_231#_c_523_n N_A_706_66#_c_704_n 0.00111924f $X=7.815 $Y=0.98
+ $X2=0 $Y2=0
cc_466 N_A_1530_231#_c_524_n N_A_706_66#_c_704_n 0.0038775f $X=7.815 $Y=1.32
+ $X2=0 $Y2=0
cc_467 N_A_1530_231#_c_525_n N_A_706_66#_c_704_n 0.0137309f $X=7.815 $Y=1.155
+ $X2=0 $Y2=0
cc_468 N_A_1530_231#_c_520_n N_A_706_66#_c_706_n 0.00600173f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_469 N_A_1530_231#_M1007_g N_A_975_347#_c_861_n 0.0172549f $X=7.775 $Y=2.235
+ $X2=0 $Y2=0
cc_470 N_A_1530_231#_c_520_n N_A_975_347#_c_861_n 0.00624358f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_471 N_A_1530_231#_c_522_n N_A_975_347#_M1022_g 9.5131e-19 $X=10.41 $Y=0.35
+ $X2=0 $Y2=0
cc_472 N_A_1530_231#_c_522_n N_A_2089_254#_M1001_g 3.95743e-19 $X=10.41 $Y=0.35
+ $X2=0 $Y2=0
cc_473 N_A_1530_231#_c_520_n N_A_1902_347#_c_1128_n 0.0151161f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_474 N_A_1530_231#_c_520_n N_A_1902_347#_c_1124_n 0.0148342f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_475 N_A_1530_231#_c_520_n N_A_1902_347#_c_1132_n 0.00467678f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_476 N_A_1530_231#_M1007_g N_VPWR_c_1278_n 0.0196874f $X=7.775 $Y=2.235 $X2=0
+ $Y2=0
cc_477 N_A_1530_231#_c_520_n N_VPWR_c_1278_n 0.0233457f $X=8.91 $Y=1.88 $X2=0
+ $Y2=0
cc_478 N_A_1530_231#_c_520_n N_VPWR_c_1289_n 0.00749462f $X=8.91 $Y=1.88 $X2=0
+ $Y2=0
cc_479 N_A_1530_231#_M1007_g N_VPWR_c_1274_n 0.00141512f $X=7.775 $Y=2.235 $X2=0
+ $Y2=0
cc_480 N_A_1530_231#_c_520_n N_VPWR_c_1274_n 0.00907254f $X=8.91 $Y=1.88 $X2=0
+ $Y2=0
cc_481 N_A_1530_231#_c_523_n N_A_343_417#_c_1451_n 0.00684186f $X=7.815 $Y=0.98
+ $X2=0 $Y2=0
cc_482 N_A_1530_231#_c_518_n N_VGND_M1009_d 0.00208561f $X=8.705 $Y=0.98 $X2=0
+ $Y2=0
cc_483 N_A_1530_231#_c_523_n N_VGND_M1009_d 0.00167665f $X=7.815 $Y=0.98 $X2=0
+ $Y2=0
cc_484 N_A_1530_231#_c_518_n N_VGND_c_1612_n 0.0142305f $X=8.705 $Y=0.98 $X2=0
+ $Y2=0
cc_485 N_A_1530_231#_c_519_n N_VGND_c_1612_n 0.00805647f $X=8.87 $Y=0.835 $X2=0
+ $Y2=0
cc_486 N_A_1530_231#_c_521_n N_VGND_c_1612_n 0.00686833f $X=9.075 $Y=0.35 $X2=0
+ $Y2=0
cc_487 N_A_1530_231#_c_523_n N_VGND_c_1612_n 0.00965762f $X=7.815 $Y=0.98 $X2=0
+ $Y2=0
cc_488 N_A_1530_231#_c_524_n N_VGND_c_1612_n 5.43878e-19 $X=7.815 $Y=1.32 $X2=0
+ $Y2=0
cc_489 N_A_1530_231#_c_525_n N_VGND_c_1612_n 0.0019223f $X=7.815 $Y=1.155 $X2=0
+ $Y2=0
cc_490 N_A_1530_231#_c_521_n N_VGND_c_1621_n 0.024922f $X=9.075 $Y=0.35 $X2=0
+ $Y2=0
cc_491 N_A_1530_231#_c_522_n N_VGND_c_1621_n 0.0902505f $X=10.41 $Y=0.35 $X2=0
+ $Y2=0
cc_492 N_A_1530_231#_M1022_d N_VGND_c_1624_n 0.00239627f $X=10.205 $Y=0.775
+ $X2=0 $Y2=0
cc_493 N_A_1530_231#_c_521_n N_VGND_c_1624_n 0.0128084f $X=9.075 $Y=0.35 $X2=0
+ $Y2=0
cc_494 N_A_1530_231#_c_522_n N_VGND_c_1624_n 0.0553923f $X=10.41 $Y=0.35 $X2=0
+ $Y2=0
cc_495 N_A_1530_231#_c_525_n N_VGND_c_1624_n 9.49986e-19 $X=7.815 $Y=1.155 $X2=0
+ $Y2=0
cc_496 N_A_1530_231#_c_525_n N_A_1127_155#_c_1769_n 0.00119246f $X=7.815
+ $Y=1.155 $X2=0 $Y2=0
cc_497 N_A_1530_231#_c_518_n A_1674_125# 0.00166171f $X=8.705 $Y=0.98 $X2=-0.19
+ $Y2=-0.245
cc_498 N_A_1530_231#_c_519_n N_A_1859_155#_c_1800_n 0.00815185f $X=8.87 $Y=0.835
+ $X2=0 $Y2=0
cc_499 N_A_1530_231#_c_520_n N_A_1859_155#_c_1800_n 0.0110873f $X=8.91 $Y=1.88
+ $X2=0 $Y2=0
cc_500 N_A_1530_231#_c_538_p N_A_1859_155#_c_1800_n 0.0133773f $X=8.89 $Y=0.98
+ $X2=0 $Y2=0
cc_501 N_A_1530_231#_M1022_d N_A_1859_155#_c_1801_n 0.0124064f $X=10.205
+ $Y=0.775 $X2=0 $Y2=0
cc_502 N_A_1530_231#_c_522_n N_A_1859_155#_c_1801_n 0.0718716f $X=10.41 $Y=0.35
+ $X2=0 $Y2=0
cc_503 N_A_1530_231#_c_519_n N_A_1859_155#_c_1802_n 0.0138381f $X=8.87 $Y=0.835
+ $X2=0 $Y2=0
cc_504 N_A_1530_231#_c_522_n N_A_1859_155#_c_1802_n 0.0187075f $X=10.41 $Y=0.35
+ $X2=0 $Y2=0
cc_505 N_A_1530_231#_c_522_n N_A_1859_155#_c_1803_n 0.0134878f $X=10.41 $Y=0.35
+ $X2=0 $Y2=0
cc_506 N_A_1278_155#_c_613_n N_A_706_66#_M1041_g 0.00683629f $X=6.54 $Y=1.05
+ $X2=0 $Y2=0
cc_507 N_A_1278_155#_c_614_n N_A_706_66#_M1041_g 0.00173358f $X=7.185 $Y=1.75
+ $X2=0 $Y2=0
cc_508 N_A_1278_155#_c_613_n N_A_706_66#_c_697_n 0.00229469f $X=6.54 $Y=1.05
+ $X2=0 $Y2=0
cc_509 N_A_1278_155#_c_614_n N_A_706_66#_c_697_n 0.00122688f $X=7.185 $Y=1.75
+ $X2=0 $Y2=0
cc_510 N_A_1278_155#_c_618_n N_A_706_66#_M1038_g 0.0186025f $X=7.02 $Y=1.88
+ $X2=0 $Y2=0
cc_511 N_A_1278_155#_c_619_n N_A_706_66#_M1038_g 0.024785f $X=8.22 $Y=1.75 $X2=0
+ $Y2=0
cc_512 N_A_1278_155#_c_614_n N_A_706_66#_M1038_g 0.0122003f $X=7.185 $Y=1.75
+ $X2=0 $Y2=0
cc_513 N_A_1278_155#_M1028_g N_A_706_66#_c_699_n 0.00868355f $X=8.295 $Y=0.835
+ $X2=0 $Y2=0
cc_514 N_A_1278_155#_M1018_g N_A_706_66#_c_699_n 0.00847339f $X=8.655 $Y=0.835
+ $X2=0 $Y2=0
cc_515 N_A_1278_155#_M1018_g N_A_706_66#_c_700_n 0.0185804f $X=8.655 $Y=0.835
+ $X2=0 $Y2=0
cc_516 N_A_1278_155#_c_616_n N_A_706_66#_c_700_n 0.00728703f $X=8.655 $Y=1.41
+ $X2=0 $Y2=0
cc_517 N_A_1278_155#_c_616_n N_A_706_66#_M1024_g 0.01826f $X=8.655 $Y=1.41 $X2=0
+ $Y2=0
cc_518 N_A_1278_155#_c_613_n N_A_706_66#_c_704_n 3.22591e-19 $X=6.54 $Y=1.05
+ $X2=0 $Y2=0
cc_519 N_A_1278_155#_c_613_n N_A_975_347#_c_847_n 0.00305853f $X=6.54 $Y=1.05
+ $X2=0 $Y2=0
cc_520 N_A_1278_155#_c_614_n N_A_975_347#_c_847_n 0.00273606f $X=7.185 $Y=1.75
+ $X2=0 $Y2=0
cc_521 N_A_1278_155#_c_613_n N_A_975_347#_c_849_n 0.00496621f $X=6.54 $Y=1.05
+ $X2=0 $Y2=0
cc_522 N_A_1278_155#_c_618_n N_A_975_347#_M1010_g 0.0168151f $X=7.02 $Y=1.88
+ $X2=0 $Y2=0
cc_523 N_A_1278_155#_c_614_n N_A_975_347#_M1010_g 0.0145147f $X=7.185 $Y=1.75
+ $X2=0 $Y2=0
cc_524 N_A_1278_155#_M1013_g N_A_975_347#_c_861_n 0.0172445f $X=8.645 $Y=2.235
+ $X2=0 $Y2=0
cc_525 N_A_1278_155#_c_618_n N_A_975_347#_c_861_n 0.00392786f $X=7.02 $Y=1.88
+ $X2=0 $Y2=0
cc_526 N_A_1278_155#_c_619_n N_VPWR_M1007_d 0.0151336f $X=8.22 $Y=1.75 $X2=0
+ $Y2=0
cc_527 N_A_1278_155#_M1013_g N_VPWR_c_1278_n 0.0106985f $X=8.645 $Y=2.235 $X2=0
+ $Y2=0
cc_528 N_A_1278_155#_c_619_n N_VPWR_c_1278_n 0.0209601f $X=8.22 $Y=1.75 $X2=0
+ $Y2=0
cc_529 N_A_1278_155#_c_618_n N_VPWR_c_1288_n 0.0074415f $X=7.02 $Y=1.88 $X2=0
+ $Y2=0
cc_530 N_A_1278_155#_M1013_g N_VPWR_c_1274_n 0.0015654f $X=8.645 $Y=2.235 $X2=0
+ $Y2=0
cc_531 N_A_1278_155#_c_618_n N_VPWR_c_1274_n 0.00902447f $X=7.02 $Y=1.88 $X2=0
+ $Y2=0
cc_532 N_A_1278_155#_M1014_d N_A_343_417#_c_1449_n 0.00191634f $X=6.39 $Y=0.775
+ $X2=0 $Y2=0
cc_533 N_A_1278_155#_c_613_n N_A_343_417#_c_1449_n 0.0162371f $X=6.54 $Y=1.05
+ $X2=0 $Y2=0
cc_534 N_A_1278_155#_c_614_n N_A_343_417#_c_1449_n 0.00434265f $X=7.185 $Y=1.75
+ $X2=0 $Y2=0
cc_535 N_A_1278_155#_c_613_n N_A_343_417#_c_1451_n 0.0096883f $X=6.54 $Y=1.05
+ $X2=0 $Y2=0
cc_536 N_A_1278_155#_c_614_n N_A_343_417#_c_1451_n 0.0221003f $X=7.185 $Y=1.75
+ $X2=0 $Y2=0
cc_537 N_A_1278_155#_c_618_n N_A_343_417#_c_1457_n 0.0637354f $X=7.02 $Y=1.88
+ $X2=0 $Y2=0
cc_538 N_A_1278_155#_c_614_n N_A_343_417#_c_1457_n 0.0284065f $X=7.185 $Y=1.75
+ $X2=0 $Y2=0
cc_539 N_A_1278_155#_c_613_n N_A_343_417#_c_1453_n 0.0221922f $X=6.54 $Y=1.05
+ $X2=0 $Y2=0
cc_540 N_A_1278_155#_c_614_n N_A_343_417#_c_1453_n 0.0183529f $X=7.185 $Y=1.75
+ $X2=0 $Y2=0
cc_541 N_A_1278_155#_c_619_n A_1482_347# 0.0048076f $X=8.22 $Y=1.75 $X2=-0.19
+ $Y2=-0.245
cc_542 N_A_1278_155#_M1028_g N_VGND_c_1612_n 0.00245827f $X=8.295 $Y=0.835 $X2=0
+ $Y2=0
cc_543 N_A_1278_155#_M1028_g N_VGND_c_1624_n 9.49986e-19 $X=8.295 $Y=0.835 $X2=0
+ $Y2=0
cc_544 N_A_1278_155#_M1018_g N_VGND_c_1624_n 7.94319e-19 $X=8.655 $Y=0.835 $X2=0
+ $Y2=0
cc_545 N_A_706_66#_M1030_g N_A_975_347#_c_857_n 0.0184245f $X=4.75 $Y=2.235
+ $X2=0 $Y2=0
cc_546 N_A_706_66#_c_711_n N_A_975_347#_c_848_n 0.012193f $X=4.75 $Y=1.025 $X2=0
+ $Y2=0
cc_547 N_A_706_66#_c_693_n N_A_975_347#_c_849_n 0.00378063f $X=6.68 $Y=0.18
+ $X2=0 $Y2=0
cc_548 N_A_706_66#_M1041_g N_A_975_347#_c_849_n 0.014427f $X=6.755 $Y=0.985
+ $X2=0 $Y2=0
cc_549 N_A_706_66#_M1041_g N_A_975_347#_M1010_g 0.00667326f $X=6.755 $Y=0.985
+ $X2=0 $Y2=0
cc_550 N_A_706_66#_M1038_g N_A_975_347#_M1010_g 0.0128253f $X=7.285 $Y=2.235
+ $X2=0 $Y2=0
cc_551 N_A_706_66#_M1038_g N_A_975_347#_c_861_n 0.0172445f $X=7.285 $Y=2.235
+ $X2=0 $Y2=0
cc_552 N_A_706_66#_M1024_g N_A_975_347#_c_861_n 0.0173606f $X=9.385 $Y=2.235
+ $X2=0 $Y2=0
cc_553 N_A_706_66#_c_702_n N_A_975_347#_M1022_g 0.0192025f $X=9.635 $Y=1.27
+ $X2=0 $Y2=0
cc_554 N_A_706_66#_M1024_g N_A_975_347#_c_852_n 0.0305763f $X=9.385 $Y=2.235
+ $X2=0 $Y2=0
cc_555 N_A_706_66#_c_706_n N_A_975_347#_c_852_n 0.00108809f $X=9.635 $Y=1.345
+ $X2=0 $Y2=0
cc_556 N_A_706_66#_M1030_g N_A_975_347#_c_865_n 0.00498895f $X=4.75 $Y=2.235
+ $X2=0 $Y2=0
cc_557 N_A_706_66#_c_715_n N_A_975_347#_c_865_n 0.0138037f $X=4.375 $Y=1.845
+ $X2=0 $Y2=0
cc_558 N_A_706_66#_c_708_n N_A_975_347#_c_865_n 0.00447141f $X=4.375 $Y=0.915
+ $X2=0 $Y2=0
cc_559 N_A_706_66#_c_711_n N_A_975_347#_c_865_n 0.00816274f $X=4.75 $Y=1.025
+ $X2=0 $Y2=0
cc_560 N_A_706_66#_c_690_n N_A_975_347#_c_853_n 9.25422e-19 $X=4.66 $Y=0.86
+ $X2=0 $Y2=0
cc_561 N_A_706_66#_M1039_g N_A_975_347#_c_853_n 0.00716517f $X=5.02 $Y=0.54
+ $X2=0 $Y2=0
cc_562 N_A_706_66#_c_693_n N_A_975_347#_c_853_n 0.00513458f $X=6.68 $Y=0.18
+ $X2=0 $Y2=0
cc_563 N_A_706_66#_M1030_g N_A_975_347#_c_854_n 0.00405892f $X=4.75 $Y=2.235
+ $X2=0 $Y2=0
cc_564 N_A_706_66#_c_711_n N_A_975_347#_c_854_n 0.0104153f $X=4.75 $Y=1.025
+ $X2=0 $Y2=0
cc_565 N_A_706_66#_M1030_g N_A_975_347#_c_855_n 0.00711187f $X=4.75 $Y=2.235
+ $X2=0 $Y2=0
cc_566 N_A_706_66#_M1039_g N_A_975_347#_c_856_n 0.0104153f $X=5.02 $Y=0.54 $X2=0
+ $Y2=0
cc_567 N_A_706_66#_c_708_n N_A_975_347#_c_856_n 0.0349414f $X=4.375 $Y=0.915
+ $X2=0 $Y2=0
cc_568 N_A_706_66#_M1024_g N_A_1902_347#_c_1128_n 0.00649345f $X=9.385 $Y=2.235
+ $X2=0 $Y2=0
cc_569 N_A_706_66#_M1024_g N_A_1902_347#_c_1124_n 0.00360165f $X=9.385 $Y=2.235
+ $X2=0 $Y2=0
cc_570 N_A_706_66#_c_702_n N_A_1902_347#_c_1124_n 0.00489605f $X=9.635 $Y=1.27
+ $X2=0 $Y2=0
cc_571 N_A_706_66#_M1024_g N_A_1902_347#_c_1132_n 0.00178373f $X=9.385 $Y=2.235
+ $X2=0 $Y2=0
cc_572 N_A_706_66#_c_706_n N_A_1902_347#_c_1132_n 0.00543608f $X=9.635 $Y=1.345
+ $X2=0 $Y2=0
cc_573 N_A_706_66#_c_715_n N_VPWR_M1005_d 0.00446866f $X=4.375 $Y=1.845 $X2=0
+ $Y2=0
cc_574 N_A_706_66#_M1030_g N_VPWR_c_1277_n 0.0184641f $X=4.75 $Y=2.235 $X2=0
+ $Y2=0
cc_575 N_A_706_66#_M1038_g N_VPWR_c_1278_n 0.0036745f $X=7.285 $Y=2.235 $X2=0
+ $Y2=0
cc_576 N_A_706_66#_M1030_g N_VPWR_c_1288_n 0.00646289f $X=4.75 $Y=2.235 $X2=0
+ $Y2=0
cc_577 N_A_706_66#_M1030_g N_VPWR_c_1274_n 0.00719887f $X=4.75 $Y=2.235 $X2=0
+ $Y2=0
cc_578 N_A_706_66#_M1038_g N_VPWR_c_1274_n 0.0015654f $X=7.285 $Y=2.235 $X2=0
+ $Y2=0
cc_579 N_A_706_66#_M1024_g N_VPWR_c_1274_n 0.0015654f $X=9.385 $Y=2.235 $X2=0
+ $Y2=0
cc_580 N_A_706_66#_M1005_s N_A_343_417#_c_1456_n 0.0119732f $X=3.81 $Y=1.735
+ $X2=0 $Y2=0
cc_581 N_A_706_66#_M1030_g N_A_343_417#_c_1456_n 0.0257642f $X=4.75 $Y=2.235
+ $X2=0 $Y2=0
cc_582 N_A_706_66#_c_715_n N_A_343_417#_c_1456_n 0.0457322f $X=4.375 $Y=1.845
+ $X2=0 $Y2=0
cc_583 N_A_706_66#_c_708_n N_A_343_417#_c_1456_n 0.00745327f $X=4.375 $Y=0.915
+ $X2=0 $Y2=0
cc_584 N_A_706_66#_M1041_g N_A_343_417#_c_1449_n 0.0122763f $X=6.755 $Y=0.985
+ $X2=0 $Y2=0
cc_585 N_A_706_66#_c_704_n N_A_343_417#_c_1449_n 0.00175014f $X=7.285 $Y=1.27
+ $X2=0 $Y2=0
cc_586 N_A_706_66#_M1041_g N_A_343_417#_c_1451_n 2.60089e-19 $X=6.755 $Y=0.985
+ $X2=0 $Y2=0
cc_587 N_A_706_66#_c_704_n N_A_343_417#_c_1451_n 0.00529114f $X=7.285 $Y=1.27
+ $X2=0 $Y2=0
cc_588 N_A_706_66#_M1038_g N_A_343_417#_c_1457_n 2.60115e-19 $X=7.285 $Y=2.235
+ $X2=0 $Y2=0
cc_589 N_A_706_66#_c_707_n N_VGND_c_1609_n 0.0373045f $X=3.655 $Y=0.54 $X2=0
+ $Y2=0
cc_590 N_A_706_66#_c_709_n N_VGND_c_1609_n 0.0129575f $X=3.82 $Y=0.915 $X2=0
+ $Y2=0
cc_591 N_A_706_66#_c_690_n N_VGND_c_1610_n 0.00983875f $X=4.66 $Y=0.86 $X2=0
+ $Y2=0
cc_592 N_A_706_66#_c_694_n N_VGND_c_1610_n 0.0038616f $X=5.095 $Y=0.18 $X2=0
+ $Y2=0
cc_593 N_A_706_66#_c_707_n N_VGND_c_1610_n 0.0113755f $X=3.655 $Y=0.54 $X2=0
+ $Y2=0
cc_594 N_A_706_66#_c_708_n N_VGND_c_1610_n 0.0218683f $X=4.375 $Y=0.915 $X2=0
+ $Y2=0
cc_595 N_A_706_66#_c_690_n N_VGND_c_1611_n 0.00411131f $X=4.66 $Y=0.86 $X2=0
+ $Y2=0
cc_596 N_A_706_66#_c_694_n N_VGND_c_1611_n 0.0708265f $X=5.095 $Y=0.18 $X2=0
+ $Y2=0
cc_597 N_A_706_66#_c_699_n N_VGND_c_1612_n 0.0255216f $X=9.07 $Y=0.18 $X2=0
+ $Y2=0
cc_598 N_A_706_66#_c_704_n N_VGND_c_1612_n 0.00106263f $X=7.285 $Y=1.27 $X2=0
+ $Y2=0
cc_599 N_A_706_66#_c_707_n N_VGND_c_1620_n 0.0173629f $X=3.655 $Y=0.54 $X2=0
+ $Y2=0
cc_600 N_A_706_66#_c_699_n N_VGND_c_1621_n 0.0298216f $X=9.07 $Y=0.18 $X2=0
+ $Y2=0
cc_601 N_A_706_66#_c_690_n N_VGND_c_1624_n 0.00401612f $X=4.66 $Y=0.86 $X2=0
+ $Y2=0
cc_602 N_A_706_66#_c_693_n N_VGND_c_1624_n 0.0433171f $X=6.68 $Y=0.18 $X2=0
+ $Y2=0
cc_603 N_A_706_66#_c_694_n N_VGND_c_1624_n 0.0101746f $X=5.095 $Y=0.18 $X2=0
+ $Y2=0
cc_604 N_A_706_66#_c_696_n N_VGND_c_1624_n 0.00813257f $X=7.17 $Y=0.18 $X2=0
+ $Y2=0
cc_605 N_A_706_66#_c_699_n N_VGND_c_1624_n 0.0537286f $X=9.07 $Y=0.18 $X2=0
+ $Y2=0
cc_606 N_A_706_66#_c_703_n N_VGND_c_1624_n 0.00371014f $X=6.755 $Y=0.18 $X2=0
+ $Y2=0
cc_607 N_A_706_66#_c_705_n N_VGND_c_1624_n 0.00371014f $X=7.245 $Y=0.18 $X2=0
+ $Y2=0
cc_608 N_A_706_66#_c_707_n N_VGND_c_1624_n 0.0122896f $X=3.655 $Y=0.54 $X2=0
+ $Y2=0
cc_609 N_A_706_66#_c_708_n N_VGND_c_1624_n 0.0264313f $X=4.375 $Y=0.915 $X2=0
+ $Y2=0
cc_610 N_A_706_66#_c_693_n N_A_1127_155#_c_1767_n 0.0152969f $X=6.68 $Y=0.18
+ $X2=0 $Y2=0
cc_611 N_A_706_66#_M1041_g N_A_1127_155#_c_1767_n 0.0122426f $X=6.755 $Y=0.985
+ $X2=0 $Y2=0
cc_612 N_A_706_66#_c_696_n N_A_1127_155#_c_1767_n 0.00373676f $X=7.17 $Y=0.18
+ $X2=0 $Y2=0
cc_613 N_A_706_66#_c_699_n N_A_1127_155#_c_1767_n 0.00480075f $X=9.07 $Y=0.18
+ $X2=0 $Y2=0
cc_614 N_A_706_66#_c_704_n N_A_1127_155#_c_1767_n 0.0160569f $X=7.285 $Y=1.27
+ $X2=0 $Y2=0
cc_615 N_A_706_66#_M1039_g N_A_1127_155#_c_1768_n 0.00159081f $X=5.02 $Y=0.54
+ $X2=0 $Y2=0
cc_616 N_A_706_66#_c_693_n N_A_1127_155#_c_1768_n 0.00615835f $X=6.68 $Y=0.18
+ $X2=0 $Y2=0
cc_617 N_A_706_66#_c_697_n N_A_1127_155#_c_1769_n 0.00228233f $X=7.285 $Y=1.395
+ $X2=0 $Y2=0
cc_618 N_A_706_66#_c_704_n N_A_1127_155#_c_1769_n 0.00903572f $X=7.285 $Y=1.27
+ $X2=0 $Y2=0
cc_619 N_A_706_66#_c_700_n N_A_1859_155#_c_1800_n 0.0036617f $X=9.145 $Y=1.27
+ $X2=0 $Y2=0
cc_620 N_A_706_66#_c_702_n N_A_1859_155#_c_1800_n 2.79531e-19 $X=9.635 $Y=1.27
+ $X2=0 $Y2=0
cc_621 N_A_706_66#_c_706_n N_A_1859_155#_c_1800_n 0.00859761f $X=9.635 $Y=1.345
+ $X2=0 $Y2=0
cc_622 N_A_706_66#_c_702_n N_A_1859_155#_c_1801_n 0.0140961f $X=9.635 $Y=1.27
+ $X2=0 $Y2=0
cc_623 N_A_706_66#_c_700_n N_A_1859_155#_c_1802_n 0.00203807f $X=9.145 $Y=1.27
+ $X2=0 $Y2=0
cc_624 N_A_975_347#_M1022_g N_A_2089_254#_c_951_n 0.0060673f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_625 N_A_975_347#_M1022_g N_A_2089_254#_c_957_n 0.00200781f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_626 N_A_975_347#_M1022_g N_A_2089_254#_c_959_n 0.00163469f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_627 N_A_975_347#_M1033_g N_A_2089_254#_c_968_n 0.0743485f $X=10.075 $Y=2.26
+ $X2=0 $Y2=0
cc_628 N_A_975_347#_M1022_g N_A_2089_254#_c_968_n 0.015059f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_629 N_A_975_347#_c_861_n N_A_1902_347#_c_1128_n 0.00608619f $X=9.95 $Y=3.15
+ $X2=0 $Y2=0
cc_630 N_A_975_347#_M1033_g N_A_1902_347#_c_1128_n 0.00620234f $X=10.075 $Y=2.26
+ $X2=0 $Y2=0
cc_631 N_A_975_347#_M1033_g N_A_1902_347#_c_1124_n 0.00675518f $X=10.075 $Y=2.26
+ $X2=0 $Y2=0
cc_632 N_A_975_347#_M1022_g N_A_1902_347#_c_1124_n 0.0102815f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_633 N_A_975_347#_c_852_n N_A_1902_347#_c_1124_n 0.00794476f $X=10.077 $Y=1.55
+ $X2=0 $Y2=0
cc_634 N_A_975_347#_M1033_g N_A_1902_347#_c_1130_n 0.014166f $X=10.075 $Y=2.26
+ $X2=0 $Y2=0
cc_635 N_A_975_347#_M1033_g N_A_1902_347#_c_1132_n 0.0136777f $X=10.075 $Y=2.26
+ $X2=0 $Y2=0
cc_636 N_A_975_347#_c_861_n N_VPWR_c_1278_n 0.025796f $X=9.95 $Y=3.15 $X2=0
+ $Y2=0
cc_637 N_A_975_347#_M1033_g N_VPWR_c_1279_n 0.00866561f $X=10.075 $Y=2.26 $X2=0
+ $Y2=0
cc_638 N_A_975_347#_c_859_n N_VPWR_c_1288_n 0.0749139f $X=5.665 $Y=3.15 $X2=0
+ $Y2=0
cc_639 N_A_975_347#_c_861_n N_VPWR_c_1289_n 0.0641473f $X=9.95 $Y=3.15 $X2=0
+ $Y2=0
cc_640 N_A_975_347#_c_858_n N_VPWR_c_1274_n 0.0360637f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_641 N_A_975_347#_c_859_n N_VPWR_c_1274_n 0.0116041f $X=5.665 $Y=3.15 $X2=0
+ $Y2=0
cc_642 N_A_975_347#_c_861_n N_VPWR_c_1274_n 0.119485f $X=9.95 $Y=3.15 $X2=0
+ $Y2=0
cc_643 N_A_975_347#_c_864_n N_VPWR_c_1274_n 0.0138136f $X=6.755 $Y=3.15 $X2=0
+ $Y2=0
cc_644 N_A_975_347#_M1030_d N_A_343_417#_c_1456_n 0.0120199f $X=4.875 $Y=1.735
+ $X2=0 $Y2=0
cc_645 N_A_975_347#_c_857_n N_A_343_417#_c_1456_n 0.0181654f $X=5.59 $Y=3.075
+ $X2=0 $Y2=0
cc_646 N_A_975_347#_c_863_n N_A_343_417#_c_1456_n 0.00123832f $X=5.5 $Y=1.975
+ $X2=0 $Y2=0
cc_647 N_A_975_347#_c_865_n N_A_343_417#_c_1456_n 0.023263f $X=5.23 $Y=1.845
+ $X2=0 $Y2=0
cc_648 N_A_975_347#_c_854_n N_A_343_417#_c_1456_n 0.0326591f $X=5.5 $Y=1.47
+ $X2=0 $Y2=0
cc_649 N_A_975_347#_c_849_n N_A_343_417#_c_1449_n 0.0131405f $X=6.315 $Y=1.305
+ $X2=0 $Y2=0
cc_650 N_A_975_347#_c_857_n N_A_343_417#_c_1457_n 0.014713f $X=5.59 $Y=3.075
+ $X2=0 $Y2=0
cc_651 N_A_975_347#_c_847_n N_A_343_417#_c_1457_n 0.00744664f $X=6.24 $Y=1.38
+ $X2=0 $Y2=0
cc_652 N_A_975_347#_c_858_n N_A_343_417#_c_1457_n 0.0104411f $X=6.63 $Y=3.15
+ $X2=0 $Y2=0
cc_653 N_A_975_347#_M1010_g N_A_343_417#_c_1457_n 0.0184865f $X=6.755 $Y=2.235
+ $X2=0 $Y2=0
cc_654 N_A_975_347#_c_863_n N_A_343_417#_c_1457_n 0.00730077f $X=5.5 $Y=1.975
+ $X2=0 $Y2=0
cc_655 N_A_975_347#_c_847_n N_A_343_417#_c_1453_n 0.0156266f $X=6.24 $Y=1.38
+ $X2=0 $Y2=0
cc_656 N_A_975_347#_c_849_n N_A_343_417#_c_1453_n 0.0103775f $X=6.315 $Y=1.305
+ $X2=0 $Y2=0
cc_657 N_A_975_347#_M1010_g N_A_343_417#_c_1453_n 0.00248252f $X=6.755 $Y=2.235
+ $X2=0 $Y2=0
cc_658 N_A_975_347#_c_854_n N_A_343_417#_c_1453_n 0.029516f $X=5.5 $Y=1.47 $X2=0
+ $Y2=0
cc_659 N_A_975_347#_c_855_n N_A_343_417#_c_1453_n 0.00730077f $X=5.5 $Y=1.47
+ $X2=0 $Y2=0
cc_660 N_A_975_347#_c_856_n N_A_343_417#_c_1453_n 0.00535296f $X=5.445 $Y=1.305
+ $X2=0 $Y2=0
cc_661 N_A_975_347#_c_853_n N_VGND_c_1610_n 0.0113755f $X=5.235 $Y=0.48 $X2=0
+ $Y2=0
cc_662 N_A_975_347#_c_853_n N_VGND_c_1611_n 0.0169315f $X=5.235 $Y=0.48 $X2=0
+ $Y2=0
cc_663 N_A_975_347#_c_853_n N_VGND_c_1624_n 0.0109178f $X=5.235 $Y=0.48 $X2=0
+ $Y2=0
cc_664 N_A_975_347#_c_848_n N_A_1127_155#_c_1766_n 0.00803894f $X=5.665 $Y=1.38
+ $X2=0 $Y2=0
cc_665 N_A_975_347#_c_849_n N_A_1127_155#_c_1766_n 0.00119826f $X=6.315 $Y=1.305
+ $X2=0 $Y2=0
cc_666 N_A_975_347#_c_853_n N_A_1127_155#_c_1766_n 0.0493124f $X=5.235 $Y=0.48
+ $X2=0 $Y2=0
cc_667 N_A_975_347#_c_854_n N_A_1127_155#_c_1766_n 0.00532952f $X=5.5 $Y=1.47
+ $X2=0 $Y2=0
cc_668 N_A_975_347#_c_849_n N_A_1127_155#_c_1767_n 4.81812e-19 $X=6.315 $Y=1.305
+ $X2=0 $Y2=0
cc_669 N_A_975_347#_c_853_n N_A_1127_155#_c_1768_n 0.0100356f $X=5.235 $Y=0.48
+ $X2=0 $Y2=0
cc_670 N_A_975_347#_M1022_g N_A_1859_155#_c_1801_n 0.0153104f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_671 N_A_975_347#_c_852_n N_A_1859_155#_c_1801_n 2.43383e-19 $X=10.077 $Y=1.55
+ $X2=0 $Y2=0
cc_672 N_A_2089_254#_c_960_n N_A_1902_347#_M1000_g 0.00641062f $X=11.815 $Y=2.13
+ $X2=0 $Y2=0
cc_673 N_A_2089_254#_c_976_n N_A_1902_347#_M1000_g 0.00882313f $X=11.525
+ $Y=2.295 $X2=0 $Y2=0
cc_674 N_A_2089_254#_c_977_n N_A_1902_347#_M1000_g 0.00305221f $X=11.815
+ $Y=2.215 $X2=0 $Y2=0
cc_675 N_A_2089_254#_M1001_g N_A_1902_347#_c_1119_n 0.0136879f $X=11.15 $Y=0.495
+ $X2=0 $Y2=0
cc_676 N_A_2089_254#_c_961_n N_A_1902_347#_c_1119_n 0.00133433f $X=12.155
+ $Y=0.495 $X2=0 $Y2=0
cc_677 N_A_2089_254#_c_963_n N_A_1902_347#_c_1119_n 4.60652e-19 $X=12.32 $Y=0.35
+ $X2=0 $Y2=0
cc_678 N_A_2089_254#_c_949_n N_A_1902_347#_c_1120_n 0.00444378f $X=10.82 $Y=1.27
+ $X2=0 $Y2=0
cc_679 N_A_2089_254#_c_957_n N_A_1902_347#_c_1120_n 8.84011e-19 $X=10.73
+ $Y=1.435 $X2=0 $Y2=0
cc_680 N_A_2089_254#_c_958_n N_A_1902_347#_c_1120_n 0.0191506f $X=11.73 $Y=1.05
+ $X2=0 $Y2=0
cc_681 N_A_2089_254#_c_960_n N_A_1902_347#_c_1120_n 0.0159339f $X=11.815 $Y=2.13
+ $X2=0 $Y2=0
cc_682 N_A_2089_254#_c_966_n N_A_1902_347#_c_1120_n 0.00140844f $X=11.815
+ $Y=0.945 $X2=0 $Y2=0
cc_683 N_A_2089_254#_c_958_n N_A_1902_347#_c_1121_n 0.00355951f $X=11.73 $Y=1.05
+ $X2=0 $Y2=0
cc_684 N_A_2089_254#_c_966_n N_A_1902_347#_c_1121_n 0.0162007f $X=11.815
+ $Y=0.945 $X2=0 $Y2=0
cc_685 N_A_2089_254#_c_961_n N_A_1902_347#_c_1122_n 0.00732971f $X=12.155
+ $Y=0.495 $X2=0 $Y2=0
cc_686 N_A_2089_254#_c_963_n N_A_1902_347#_c_1122_n 0.0037573f $X=12.32 $Y=0.35
+ $X2=0 $Y2=0
cc_687 N_A_2089_254#_c_966_n N_A_1902_347#_c_1122_n 0.00291995f $X=11.815
+ $Y=0.945 $X2=0 $Y2=0
cc_688 N_A_2089_254#_c_950_n N_A_1902_347#_c_1123_n 0.0136879f $X=11.075 $Y=1
+ $X2=0 $Y2=0
cc_689 N_A_2089_254#_c_951_n N_A_1902_347#_c_1124_n 2.55335e-19 $X=10.895 $Y=1
+ $X2=0 $Y2=0
cc_690 N_A_2089_254#_c_957_n N_A_1902_347#_c_1124_n 0.0153704f $X=10.73 $Y=1.435
+ $X2=0 $Y2=0
cc_691 N_A_2089_254#_c_959_n N_A_1902_347#_c_1124_n 0.0065444f $X=10.895 $Y=1.05
+ $X2=0 $Y2=0
cc_692 N_A_2089_254#_c_968_n N_A_1902_347#_c_1124_n 0.00172326f $X=10.82
+ $Y=1.435 $X2=0 $Y2=0
cc_693 N_A_2089_254#_M1000_d N_A_1902_347#_c_1130_n 0.00286131f $X=11.385
+ $Y=1.805 $X2=0 $Y2=0
cc_694 N_A_2089_254#_M1034_g N_A_1902_347#_c_1130_n 0.0264034f $X=10.57 $Y=2.26
+ $X2=0 $Y2=0
cc_695 N_A_2089_254#_c_957_n N_A_1902_347#_c_1130_n 0.0222146f $X=10.73 $Y=1.435
+ $X2=0 $Y2=0
cc_696 N_A_2089_254#_c_958_n N_A_1902_347#_c_1130_n 0.00904887f $X=11.73 $Y=1.05
+ $X2=0 $Y2=0
cc_697 N_A_2089_254#_c_960_n N_A_1902_347#_c_1130_n 0.0135268f $X=11.815 $Y=2.13
+ $X2=0 $Y2=0
cc_698 N_A_2089_254#_c_977_n N_A_1902_347#_c_1130_n 0.0101481f $X=11.815
+ $Y=2.215 $X2=0 $Y2=0
cc_699 N_A_2089_254#_c_968_n N_A_1902_347#_c_1130_n 0.00124448f $X=10.82
+ $Y=1.435 $X2=0 $Y2=0
cc_700 N_A_2089_254#_M1034_g N_A_1902_347#_c_1125_n 9.19697e-19 $X=10.57 $Y=2.26
+ $X2=0 $Y2=0
cc_701 N_A_2089_254#_c_957_n N_A_1902_347#_c_1125_n 0.0127287f $X=10.73 $Y=1.435
+ $X2=0 $Y2=0
cc_702 N_A_2089_254#_c_958_n N_A_1902_347#_c_1125_n 0.0247942f $X=11.73 $Y=1.05
+ $X2=0 $Y2=0
cc_703 N_A_2089_254#_c_960_n N_A_1902_347#_c_1125_n 0.033993f $X=11.815 $Y=2.13
+ $X2=0 $Y2=0
cc_704 N_A_2089_254#_c_968_n N_A_1902_347#_c_1125_n 9.75898e-19 $X=10.82
+ $Y=1.435 $X2=0 $Y2=0
cc_705 N_A_2089_254#_M1034_g N_A_1902_347#_c_1132_n 3.34489e-19 $X=10.57 $Y=2.26
+ $X2=0 $Y2=0
cc_706 N_A_2089_254#_M1034_g N_A_1902_347#_c_1126_n 0.0307373f $X=10.57 $Y=2.26
+ $X2=0 $Y2=0
cc_707 N_A_2089_254#_c_950_n N_A_1902_347#_c_1126_n 0.00505209f $X=11.075 $Y=1
+ $X2=0 $Y2=0
cc_708 N_A_2089_254#_c_957_n N_A_1902_347#_c_1126_n 0.00120089f $X=10.73
+ $Y=1.435 $X2=0 $Y2=0
cc_709 N_A_2089_254#_c_958_n N_A_1902_347#_c_1126_n 0.0028919f $X=11.73 $Y=1.05
+ $X2=0 $Y2=0
cc_710 N_A_2089_254#_c_977_n N_A_1902_347#_c_1126_n 0.0036686f $X=11.815
+ $Y=2.215 $X2=0 $Y2=0
cc_711 N_A_2089_254#_c_968_n N_A_1902_347#_c_1126_n 0.0159182f $X=10.82 $Y=1.435
+ $X2=0 $Y2=0
cc_712 N_A_2089_254#_M1011_g N_A_2714_401#_c_1220_n 0.00377468f $X=13.445
+ $Y=2.505 $X2=0 $Y2=0
cc_713 N_A_2089_254#_c_965_n N_A_2714_401#_c_1220_n 0.0265437f $X=14 $Y=1.64
+ $X2=0 $Y2=0
cc_714 N_A_2089_254#_c_969_n N_A_2714_401#_c_1220_n 0.00814315f $X=14.04 $Y=1.64
+ $X2=0 $Y2=0
cc_715 N_A_2089_254#_M1032_g N_A_2714_401#_c_1221_n 2.28436e-19 $X=12.915
+ $Y=2.505 $X2=0 $Y2=0
cc_716 N_A_2089_254#_M1011_g N_A_2714_401#_c_1221_n 0.015148f $X=13.445 $Y=2.505
+ $X2=0 $Y2=0
cc_717 N_A_2089_254#_c_965_n N_A_2714_401#_c_1222_n 0.0208405f $X=14 $Y=1.64
+ $X2=0 $Y2=0
cc_718 N_A_2089_254#_c_969_n N_A_2714_401#_c_1222_n 0.00739336f $X=14.04 $Y=1.64
+ $X2=0 $Y2=0
cc_719 N_A_2089_254#_M1029_g N_A_2714_401#_c_1214_n 0.0012512f $X=13.68 $Y=0.845
+ $X2=0 $Y2=0
cc_720 N_A_2089_254#_M1023_g N_A_2714_401#_c_1214_n 0.00954654f $X=14.04
+ $Y=0.845 $X2=0 $Y2=0
cc_721 N_A_2089_254#_c_965_n N_A_2714_401#_c_1214_n 0.00312582f $X=14 $Y=1.64
+ $X2=0 $Y2=0
cc_722 N_A_2089_254#_c_969_n N_A_2714_401#_c_1214_n 9.88065e-19 $X=14.04 $Y=1.64
+ $X2=0 $Y2=0
cc_723 N_A_2089_254#_M1023_g N_A_2714_401#_c_1215_n 0.00974994f $X=14.04
+ $Y=0.845 $X2=0 $Y2=0
cc_724 N_A_2089_254#_c_965_n N_A_2714_401#_c_1217_n 0.0256723f $X=14 $Y=1.64
+ $X2=0 $Y2=0
cc_725 N_A_2089_254#_c_969_n N_A_2714_401#_c_1217_n 0.00113627f $X=14.04 $Y=1.64
+ $X2=0 $Y2=0
cc_726 N_A_2089_254#_M1023_g N_A_2714_401#_c_1218_n 0.0142038f $X=14.04 $Y=0.845
+ $X2=0 $Y2=0
cc_727 N_A_2089_254#_c_965_n N_A_2714_401#_c_1218_n 3.29687e-19 $X=14 $Y=1.64
+ $X2=0 $Y2=0
cc_728 N_A_2089_254#_c_969_n N_A_2714_401#_c_1218_n 0.0123908f $X=14.04 $Y=1.64
+ $X2=0 $Y2=0
cc_729 N_A_2089_254#_M1034_g N_VPWR_c_1279_n 0.0082347f $X=10.57 $Y=2.26 $X2=0
+ $Y2=0
cc_730 N_A_2089_254#_c_976_n N_VPWR_c_1279_n 0.0137792f $X=11.525 $Y=2.295 $X2=0
+ $Y2=0
cc_731 N_A_2089_254#_M1032_g N_VPWR_c_1280_n 0.0237779f $X=12.915 $Y=2.505 $X2=0
+ $Y2=0
cc_732 N_A_2089_254#_M1011_g N_VPWR_c_1280_n 0.0246323f $X=13.445 $Y=2.505 $X2=0
+ $Y2=0
cc_733 N_A_2089_254#_c_965_n N_VPWR_c_1280_n 0.0187596f $X=14 $Y=1.64 $X2=0
+ $Y2=0
cc_734 N_A_2089_254#_c_967_n N_VPWR_c_1280_n 0.00791636f $X=12.98 $Y=1.64 $X2=0
+ $Y2=0
cc_735 N_A_2089_254#_c_969_n N_VPWR_c_1280_n 0.00270827f $X=14.04 $Y=1.64 $X2=0
+ $Y2=0
cc_736 N_A_2089_254#_M1011_g N_VPWR_c_1281_n 0.00356684f $X=13.445 $Y=2.505
+ $X2=0 $Y2=0
cc_737 N_A_2089_254#_M1011_g N_VPWR_c_1284_n 0.00717535f $X=13.445 $Y=2.505
+ $X2=0 $Y2=0
cc_738 N_A_2089_254#_M1034_g N_VPWR_c_1289_n 0.00742524f $X=10.57 $Y=2.26 $X2=0
+ $Y2=0
cc_739 N_A_2089_254#_M1032_g N_VPWR_c_1290_n 0.00692317f $X=12.915 $Y=2.505
+ $X2=0 $Y2=0
cc_740 N_A_2089_254#_c_976_n N_VPWR_c_1290_n 0.00872995f $X=11.525 $Y=2.295
+ $X2=0 $Y2=0
cc_741 N_A_2089_254#_M1034_g N_VPWR_c_1274_n 0.00808164f $X=10.57 $Y=2.26 $X2=0
+ $Y2=0
cc_742 N_A_2089_254#_M1032_g N_VPWR_c_1274_n 0.0129547f $X=12.915 $Y=2.505 $X2=0
+ $Y2=0
cc_743 N_A_2089_254#_M1011_g N_VPWR_c_1274_n 0.0136934f $X=13.445 $Y=2.505 $X2=0
+ $Y2=0
cc_744 N_A_2089_254#_c_976_n N_VPWR_c_1274_n 0.0107923f $X=11.525 $Y=2.295 $X2=0
+ $Y2=0
cc_745 N_A_2089_254#_M1043_g N_Q_c_1552_n 0.00393197f $X=12.89 $Y=0.845 $X2=0
+ $Y2=0
cc_746 N_A_2089_254#_c_964_n N_Q_c_1552_n 0.0130598f $X=13.025 $Y=1.475 $X2=0
+ $Y2=0
cc_747 N_A_2089_254#_c_966_n N_Q_c_1552_n 0.00199132f $X=11.815 $Y=0.945 $X2=0
+ $Y2=0
cc_748 N_A_2089_254#_c_967_n N_Q_c_1552_n 0.0226786f $X=12.98 $Y=1.64 $X2=0
+ $Y2=0
cc_749 N_A_2089_254#_c_969_n N_Q_c_1552_n 0.0065625f $X=14.04 $Y=1.64 $X2=0
+ $Y2=0
cc_750 N_A_2089_254#_c_960_n N_Q_c_1553_n 0.0110029f $X=11.815 $Y=2.13 $X2=0
+ $Y2=0
cc_751 N_A_2089_254#_c_966_n N_Q_c_1553_n 0.0160566f $X=11.815 $Y=0.945 $X2=0
+ $Y2=0
cc_752 N_A_2089_254#_M1043_g N_Q_c_1554_n 0.00257696f $X=12.89 $Y=0.845 $X2=0
+ $Y2=0
cc_753 N_A_2089_254#_c_961_n N_Q_c_1554_n 0.0120283f $X=12.155 $Y=0.495 $X2=0
+ $Y2=0
cc_754 N_A_2089_254#_c_962_n N_Q_c_1554_n 0.0187378f $X=12.94 $Y=0.35 $X2=0
+ $Y2=0
cc_755 N_A_2089_254#_c_964_n N_Q_c_1554_n 0.019843f $X=13.025 $Y=1.475 $X2=0
+ $Y2=0
cc_756 N_A_2089_254#_c_966_n N_Q_c_1554_n 0.0197866f $X=11.815 $Y=0.945 $X2=0
+ $Y2=0
cc_757 N_A_2089_254#_M1032_g N_Q_c_1556_n 0.0209683f $X=12.915 $Y=2.505 $X2=0
+ $Y2=0
cc_758 N_A_2089_254#_M1011_g N_Q_c_1556_n 2.6212e-19 $X=13.445 $Y=2.505 $X2=0
+ $Y2=0
cc_759 N_A_2089_254#_c_976_n N_Q_c_1556_n 0.0242444f $X=11.525 $Y=2.295 $X2=0
+ $Y2=0
cc_760 N_A_2089_254#_c_977_n N_Q_c_1556_n 0.0126921f $X=11.815 $Y=2.215 $X2=0
+ $Y2=0
cc_761 N_A_2089_254#_c_967_n N_Q_c_1556_n 0.0287998f $X=12.98 $Y=1.64 $X2=0
+ $Y2=0
cc_762 N_A_2089_254#_c_969_n N_Q_c_1556_n 0.00730196f $X=14.04 $Y=1.64 $X2=0
+ $Y2=0
cc_763 N_A_2089_254#_M1032_g N_Q_c_1555_n 0.00462368f $X=12.915 $Y=2.505 $X2=0
+ $Y2=0
cc_764 N_A_2089_254#_M1043_g N_Q_c_1555_n 0.00277607f $X=12.89 $Y=0.845 $X2=0
+ $Y2=0
cc_765 N_A_2089_254#_c_960_n N_Q_c_1555_n 0.0527095f $X=11.815 $Y=2.13 $X2=0
+ $Y2=0
cc_766 N_A_2089_254#_c_964_n N_Q_c_1555_n 0.00465229f $X=13.025 $Y=1.475 $X2=0
+ $Y2=0
cc_767 N_A_2089_254#_c_967_n N_Q_c_1555_n 0.025097f $X=12.98 $Y=1.64 $X2=0 $Y2=0
cc_768 N_A_2089_254#_c_969_n N_Q_c_1555_n 0.00225377f $X=14.04 $Y=1.64 $X2=0
+ $Y2=0
cc_769 N_A_2089_254#_M1001_g N_VGND_c_1613_n 0.00256223f $X=11.15 $Y=0.495 $X2=0
+ $Y2=0
cc_770 N_A_2089_254#_c_958_n N_VGND_c_1613_n 0.0100858f $X=11.73 $Y=1.05 $X2=0
+ $Y2=0
cc_771 N_A_2089_254#_c_961_n N_VGND_c_1613_n 0.00522496f $X=12.155 $Y=0.495
+ $X2=0 $Y2=0
cc_772 N_A_2089_254#_c_963_n N_VGND_c_1613_n 0.00591401f $X=12.32 $Y=0.35 $X2=0
+ $Y2=0
cc_773 N_A_2089_254#_M1043_g N_VGND_c_1614_n 4.59707e-19 $X=12.89 $Y=0.845 $X2=0
+ $Y2=0
cc_774 N_A_2089_254#_M1025_g N_VGND_c_1614_n 0.00922403f $X=13.25 $Y=0.845 $X2=0
+ $Y2=0
cc_775 N_A_2089_254#_M1029_g N_VGND_c_1614_n 0.0124989f $X=13.68 $Y=0.845 $X2=0
+ $Y2=0
cc_776 N_A_2089_254#_M1023_g N_VGND_c_1614_n 0.00180305f $X=14.04 $Y=0.845 $X2=0
+ $Y2=0
cc_777 N_A_2089_254#_c_962_n N_VGND_c_1614_n 0.0139003f $X=12.94 $Y=0.35 $X2=0
+ $Y2=0
cc_778 N_A_2089_254#_c_964_n N_VGND_c_1614_n 0.0439228f $X=13.025 $Y=1.475 $X2=0
+ $Y2=0
cc_779 N_A_2089_254#_c_965_n N_VGND_c_1614_n 0.0144149f $X=14 $Y=1.64 $X2=0
+ $Y2=0
cc_780 N_A_2089_254#_c_969_n N_VGND_c_1614_n 0.00232715f $X=14.04 $Y=1.64 $X2=0
+ $Y2=0
cc_781 N_A_2089_254#_M1023_g N_VGND_c_1615_n 0.00312861f $X=14.04 $Y=0.845 $X2=0
+ $Y2=0
cc_782 N_A_2089_254#_M1043_g N_VGND_c_1616_n 2.23678e-19 $X=12.89 $Y=0.845 $X2=0
+ $Y2=0
cc_783 N_A_2089_254#_M1025_g N_VGND_c_1616_n 0.00340865f $X=13.25 $Y=0.845 $X2=0
+ $Y2=0
cc_784 N_A_2089_254#_c_962_n N_VGND_c_1616_n 0.049001f $X=12.94 $Y=0.35 $X2=0
+ $Y2=0
cc_785 N_A_2089_254#_c_963_n N_VGND_c_1616_n 0.0221635f $X=12.32 $Y=0.35 $X2=0
+ $Y2=0
cc_786 N_A_2089_254#_M1001_g N_VGND_c_1621_n 0.00502664f $X=11.15 $Y=0.495 $X2=0
+ $Y2=0
cc_787 N_A_2089_254#_M1029_g N_VGND_c_1622_n 0.00340865f $X=13.68 $Y=0.845 $X2=0
+ $Y2=0
cc_788 N_A_2089_254#_M1023_g N_VGND_c_1622_n 0.00394394f $X=14.04 $Y=0.845 $X2=0
+ $Y2=0
cc_789 N_A_2089_254#_M1001_g N_VGND_c_1624_n 0.0103357f $X=11.15 $Y=0.495 $X2=0
+ $Y2=0
cc_790 N_A_2089_254#_M1025_g N_VGND_c_1624_n 0.00392009f $X=13.25 $Y=0.845 $X2=0
+ $Y2=0
cc_791 N_A_2089_254#_M1029_g N_VGND_c_1624_n 0.00392009f $X=13.68 $Y=0.845 $X2=0
+ $Y2=0
cc_792 N_A_2089_254#_M1023_g N_VGND_c_1624_n 0.00466677f $X=14.04 $Y=0.845 $X2=0
+ $Y2=0
cc_793 N_A_2089_254#_c_962_n N_VGND_c_1624_n 0.0297409f $X=12.94 $Y=0.35 $X2=0
+ $Y2=0
cc_794 N_A_2089_254#_c_963_n N_VGND_c_1624_n 0.0126536f $X=12.32 $Y=0.35 $X2=0
+ $Y2=0
cc_795 N_A_2089_254#_c_966_n N_VGND_c_1624_n 0.00947202f $X=11.815 $Y=0.945
+ $X2=0 $Y2=0
cc_796 N_A_2089_254#_c_951_n N_A_1859_155#_c_1801_n 0.00782685f $X=10.895 $Y=1
+ $X2=0 $Y2=0
cc_797 N_A_2089_254#_M1001_g N_A_1859_155#_c_1801_n 0.00600547f $X=11.15
+ $Y=0.495 $X2=0 $Y2=0
cc_798 N_A_2089_254#_c_958_n N_A_1859_155#_c_1801_n 0.0153085f $X=11.73 $Y=1.05
+ $X2=0 $Y2=0
cc_799 N_A_2089_254#_c_959_n N_A_1859_155#_c_1801_n 0.0267801f $X=10.895 $Y=1.05
+ $X2=0 $Y2=0
cc_800 N_A_2089_254#_c_966_n N_A_1859_155#_c_1801_n 3.00621e-19 $X=11.815
+ $Y=0.945 $X2=0 $Y2=0
cc_801 N_A_2089_254#_c_968_n N_A_1859_155#_c_1801_n 0.0042396f $X=10.82 $Y=1.435
+ $X2=0 $Y2=0
cc_802 N_A_2089_254#_M1001_g N_A_1859_155#_c_1803_n 0.00463537f $X=11.15
+ $Y=0.495 $X2=0 $Y2=0
cc_803 N_A_2089_254#_c_964_n A_2593_127# 0.00356941f $X=13.025 $Y=1.475
+ $X2=-0.19 $Y2=-0.245
cc_804 N_A_1902_347#_c_1130_n N_VPWR_M1034_d 0.00892257f $X=11.22 $Y=1.865 $X2=0
+ $Y2=0
cc_805 N_A_1902_347#_M1000_g N_VPWR_c_1279_n 0.00886434f $X=11.26 $Y=2.305 $X2=0
+ $Y2=0
cc_806 N_A_1902_347#_c_1130_n N_VPWR_c_1279_n 0.0254128f $X=11.22 $Y=1.865 $X2=0
+ $Y2=0
cc_807 N_A_1902_347#_c_1128_n N_VPWR_c_1289_n 0.0080024f $X=9.73 $Y=2.615 $X2=0
+ $Y2=0
cc_808 N_A_1902_347#_M1000_g N_VPWR_c_1290_n 0.00767722f $X=11.26 $Y=2.305 $X2=0
+ $Y2=0
cc_809 N_A_1902_347#_M1000_g N_VPWR_c_1274_n 0.00829933f $X=11.26 $Y=2.305 $X2=0
+ $Y2=0
cc_810 N_A_1902_347#_c_1128_n N_VPWR_c_1274_n 0.00928628f $X=9.73 $Y=2.615 $X2=0
+ $Y2=0
cc_811 N_A_1902_347#_c_1130_n A_2040_352# 0.00999675f $X=11.22 $Y=1.865
+ $X2=-0.19 $Y2=-0.245
cc_812 N_A_1902_347#_c_1120_n N_Q_c_1553_n 4.08969e-19 $X=11.58 $Y=1.315 $X2=0
+ $Y2=0
cc_813 N_A_1902_347#_c_1122_n N_Q_c_1554_n 0.001018f $X=11.94 $Y=0.78 $X2=0
+ $Y2=0
cc_814 N_A_1902_347#_c_1119_n N_VGND_c_1613_n 0.00966784f $X=11.58 $Y=0.78 $X2=0
+ $Y2=0
cc_815 N_A_1902_347#_c_1122_n N_VGND_c_1613_n 0.00174445f $X=11.94 $Y=0.78 $X2=0
+ $Y2=0
cc_816 N_A_1902_347#_c_1119_n N_VGND_c_1616_n 0.00445056f $X=11.58 $Y=0.78 $X2=0
+ $Y2=0
cc_817 N_A_1902_347#_c_1121_n N_VGND_c_1616_n 2.13211e-19 $X=11.865 $Y=0.855
+ $X2=0 $Y2=0
cc_818 N_A_1902_347#_c_1122_n N_VGND_c_1616_n 0.00501274f $X=11.94 $Y=0.78 $X2=0
+ $Y2=0
cc_819 N_A_1902_347#_c_1119_n N_VGND_c_1624_n 0.00796275f $X=11.58 $Y=0.78 $X2=0
+ $Y2=0
cc_820 N_A_1902_347#_c_1122_n N_VGND_c_1624_n 0.00642239f $X=11.94 $Y=0.78 $X2=0
+ $Y2=0
cc_821 N_A_1902_347#_c_1124_n N_A_1859_155#_c_1800_n 0.00119908f $X=9.915
+ $Y=1.05 $X2=0 $Y2=0
cc_822 N_A_1902_347#_M1042_d N_A_1859_155#_c_1801_n 0.0024717f $X=9.71 $Y=0.775
+ $X2=0 $Y2=0
cc_823 N_A_1902_347#_c_1119_n N_A_1859_155#_c_1801_n 7.8335e-19 $X=11.58 $Y=0.78
+ $X2=0 $Y2=0
cc_824 N_A_1902_347#_c_1124_n N_A_1859_155#_c_1801_n 0.0197128f $X=9.915 $Y=1.05
+ $X2=0 $Y2=0
cc_825 N_A_2714_401#_c_1222_n N_VPWR_M1027_s 0.00314466f $X=14.345 $Y=2.07 $X2=0
+ $Y2=0
cc_826 N_A_2714_401#_c_1220_n N_VPWR_c_1280_n 0.0119061f $X=13.71 $Y=2.155 $X2=0
+ $Y2=0
cc_827 N_A_2714_401#_c_1221_n N_VPWR_c_1280_n 0.0572919f $X=13.71 $Y=2.86 $X2=0
+ $Y2=0
cc_828 N_A_2714_401#_M1027_g N_VPWR_c_1281_n 0.0193529f $X=14.615 $Y=2.545 $X2=0
+ $Y2=0
cc_829 N_A_2714_401#_c_1221_n N_VPWR_c_1281_n 0.037892f $X=13.71 $Y=2.86 $X2=0
+ $Y2=0
cc_830 N_A_2714_401#_c_1222_n N_VPWR_c_1281_n 0.0219188f $X=14.345 $Y=2.07 $X2=0
+ $Y2=0
cc_831 N_A_2714_401#_c_1221_n N_VPWR_c_1284_n 0.0177662f $X=13.71 $Y=2.86 $X2=0
+ $Y2=0
cc_832 N_A_2714_401#_M1027_g N_VPWR_c_1291_n 0.00769046f $X=14.615 $Y=2.545
+ $X2=0 $Y2=0
cc_833 N_A_2714_401#_M1027_g N_VPWR_c_1274_n 0.0143431f $X=14.615 $Y=2.545 $X2=0
+ $Y2=0
cc_834 N_A_2714_401#_c_1221_n N_VPWR_c_1274_n 0.0123184f $X=13.71 $Y=2.86 $X2=0
+ $Y2=0
cc_835 N_A_2714_401#_M1027_g N_Q_N_c_1587_n 0.00805208f $X=14.615 $Y=2.545 $X2=0
+ $Y2=0
cc_836 N_A_2714_401#_M1031_g N_Q_N_c_1587_n 0.00214984f $X=15 $Y=0.495 $X2=0
+ $Y2=0
cc_837 N_A_2714_401#_c_1212_n N_Q_N_c_1587_n 0.00813286f $X=15.285 $Y=0.98 $X2=0
+ $Y2=0
cc_838 N_A_2714_401#_M1026_g N_Q_N_c_1587_n 0.0156561f $X=15.36 $Y=0.495 $X2=0
+ $Y2=0
cc_839 N_A_2714_401#_c_1214_n N_Q_N_c_1587_n 0.00495922f $X=14.585 $Y=1.075
+ $X2=0 $Y2=0
cc_840 N_A_2714_401#_c_1215_n N_Q_N_c_1587_n 0.015914f $X=14.585 $Y=1.335 $X2=0
+ $Y2=0
cc_841 N_A_2714_401#_c_1218_n N_Q_N_c_1587_n 0.0129438f $X=14.782 $Y=0.98 $X2=0
+ $Y2=0
cc_842 N_A_2714_401#_M1027_g Q_N 0.0302573f $X=14.615 $Y=2.545 $X2=0 $Y2=0
cc_843 N_A_2714_401#_c_1222_n Q_N 0.0125659f $X=14.345 $Y=2.07 $X2=0 $Y2=0
cc_844 N_A_2714_401#_c_1216_n Q_N 0.00429711f $X=14.43 $Y=1.985 $X2=0 $Y2=0
cc_845 N_A_2714_401#_c_1217_n Q_N 0.00554623f $X=14.585 $Y=1.575 $X2=0 $Y2=0
cc_846 N_A_2714_401#_c_1218_n Q_N 0.0106509f $X=14.782 $Y=0.98 $X2=0 $Y2=0
cc_847 N_A_2714_401#_c_1214_n N_VGND_c_1614_n 0.015758f $X=14.585 $Y=1.075 $X2=0
+ $Y2=0
cc_848 N_A_2714_401#_M1031_g N_VGND_c_1615_n 0.0149551f $X=15 $Y=0.495 $X2=0
+ $Y2=0
cc_849 N_A_2714_401#_M1026_g N_VGND_c_1615_n 0.002112f $X=15.36 $Y=0.495 $X2=0
+ $Y2=0
cc_850 N_A_2714_401#_c_1214_n N_VGND_c_1615_n 0.0255999f $X=14.585 $Y=1.075
+ $X2=0 $Y2=0
cc_851 N_A_2714_401#_c_1218_n N_VGND_c_1615_n 0.00633228f $X=14.782 $Y=0.98
+ $X2=0 $Y2=0
cc_852 N_A_2714_401#_c_1214_n N_VGND_c_1622_n 0.00675757f $X=14.585 $Y=1.075
+ $X2=0 $Y2=0
cc_853 N_A_2714_401#_M1031_g N_VGND_c_1623_n 0.00445056f $X=15 $Y=0.495 $X2=0
+ $Y2=0
cc_854 N_A_2714_401#_M1026_g N_VGND_c_1623_n 0.00502664f $X=15.36 $Y=0.495 $X2=0
+ $Y2=0
cc_855 N_A_2714_401#_M1031_g N_VGND_c_1624_n 0.00796275f $X=15 $Y=0.495 $X2=0
+ $Y2=0
cc_856 N_A_2714_401#_M1026_g N_VGND_c_1624_n 0.0100521f $X=15.36 $Y=0.495 $X2=0
+ $Y2=0
cc_857 N_A_2714_401#_c_1214_n N_VGND_c_1624_n 0.00999618f $X=14.585 $Y=1.075
+ $X2=0 $Y2=0
cc_858 N_VPWR_c_1274_n N_A_239_417#_M1036_s 0.00216573f $X=15.6 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_859 N_VPWR_c_1274_n N_A_239_417#_M1040_d 0.00229455f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_860 N_VPWR_c_1275_n N_A_239_417#_c_1407_n 0.0326506f $X=0.795 $Y=2.19 $X2=0
+ $Y2=0
cc_861 N_VPWR_M1006_d N_A_239_417#_c_1408_n 0.00355361f $X=2.715 $Y=2.085 $X2=0
+ $Y2=0
cc_862 N_VPWR_c_1276_n N_A_239_417#_c_1408_n 0.0152929f $X=2.855 $Y=2.94 $X2=0
+ $Y2=0
cc_863 N_VPWR_c_1282_n N_A_239_417#_c_1408_n 0.0175661f $X=2.69 $Y=3.33 $X2=0
+ $Y2=0
cc_864 N_VPWR_c_1287_n N_A_239_417#_c_1408_n 0.00310358f $X=4.32 $Y=3.33 $X2=0
+ $Y2=0
cc_865 N_VPWR_c_1274_n N_A_239_417#_c_1408_n 0.0363714f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_866 N_VPWR_c_1276_n N_A_239_417#_c_1409_n 0.013837f $X=2.855 $Y=2.94 $X2=0
+ $Y2=0
cc_867 N_VPWR_c_1287_n N_A_239_417#_c_1409_n 0.0195379f $X=4.32 $Y=3.33 $X2=0
+ $Y2=0
cc_868 N_VPWR_c_1274_n N_A_239_417#_c_1409_n 0.0125146f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_869 N_VPWR_c_1275_n N_A_239_417#_c_1410_n 0.0423439f $X=0.795 $Y=2.19 $X2=0
+ $Y2=0
cc_870 N_VPWR_c_1282_n N_A_239_417#_c_1410_n 0.0197784f $X=2.69 $Y=3.33 $X2=0
+ $Y2=0
cc_871 N_VPWR_c_1274_n N_A_239_417#_c_1410_n 0.012508f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_872 N_VPWR_c_1274_n N_A_343_417#_M1036_d 0.00333718f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_873 N_VPWR_M1006_d N_A_343_417#_c_1456_n 0.00814554f $X=2.715 $Y=2.085 $X2=0
+ $Y2=0
cc_874 N_VPWR_M1005_d N_A_343_417#_c_1456_n 0.003832f $X=4.345 $Y=1.735 $X2=0
+ $Y2=0
cc_875 N_VPWR_c_1277_n N_A_343_417#_c_1456_n 0.0163515f $X=4.485 $Y=2.59 $X2=0
+ $Y2=0
cc_876 N_VPWR_c_1288_n N_A_343_417#_c_1457_n 0.0144048f $X=7.875 $Y=3.33 $X2=0
+ $Y2=0
cc_877 N_VPWR_c_1274_n N_A_343_417#_c_1457_n 0.0173755f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_878 N_VPWR_c_1274_n A_449_417# 0.00262207f $X=15.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_879 N_VPWR_c_1280_n N_Q_c_1556_n 0.0791802f $X=13.18 $Y=2.15 $X2=0 $Y2=0
cc_880 N_VPWR_c_1290_n N_Q_c_1556_n 0.0383742f $X=13.015 $Y=3.33 $X2=0 $Y2=0
cc_881 N_VPWR_c_1274_n N_Q_c_1556_n 0.0266265f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_882 N_VPWR_c_1281_n Q_N 0.0509221f $X=14.35 $Y=2.5 $X2=0 $Y2=0
cc_883 N_VPWR_c_1291_n Q_N 0.0688921f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_884 N_VPWR_c_1274_n Q_N 0.0394726f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_885 N_A_239_417#_c_1408_n N_A_343_417#_M1036_d 0.00475803f $X=3.22 $Y=2.59
+ $X2=0 $Y2=0
cc_886 N_A_239_417#_c_1407_n N_A_343_417#_c_1454_n 0.0180693f $X=1.325 $Y=2.23
+ $X2=0 $Y2=0
cc_887 N_A_239_417#_c_1408_n N_A_343_417#_c_1454_n 0.0378922f $X=3.22 $Y=2.59
+ $X2=0 $Y2=0
cc_888 N_A_239_417#_M1040_d N_A_343_417#_c_1456_n 0.0113722f $X=3.245 $Y=2.085
+ $X2=0 $Y2=0
cc_889 N_A_239_417#_c_1408_n N_A_343_417#_c_1456_n 0.0527682f $X=3.22 $Y=2.59
+ $X2=0 $Y2=0
cc_890 N_A_239_417#_c_1408_n N_A_343_417#_c_1476_n 0.0115986f $X=3.22 $Y=2.59
+ $X2=0 $Y2=0
cc_891 N_A_239_417#_c_1408_n A_449_417# 0.00304514f $X=3.22 $Y=2.59 $X2=-0.19
+ $Y2=1.655
cc_892 N_A_343_417#_c_1454_n A_449_417# 0.00117218f $X=2.455 $Y=2.195 $X2=-0.19
+ $Y2=-0.245
cc_893 N_A_343_417#_c_1448_n N_VGND_c_1609_n 0.00112583f $X=2.54 $Y=2.065 $X2=0
+ $Y2=0
cc_894 N_A_343_417#_c_1452_n N_VGND_c_1609_n 0.0100863f $X=2.54 $Y=0.82 $X2=0
+ $Y2=0
cc_895 N_A_343_417#_c_1452_n N_VGND_c_1619_n 0.00933263f $X=2.54 $Y=0.82 $X2=0
+ $Y2=0
cc_896 N_A_343_417#_c_1452_n N_VGND_c_1624_n 0.012132f $X=2.54 $Y=0.82 $X2=0
+ $Y2=0
cc_897 N_A_343_417#_c_1453_n N_A_1127_155#_M1014_s 0.00685799f $X=6.34 $Y=1.745
+ $X2=-0.19 $Y2=-0.245
cc_898 N_A_343_417#_c_1450_n N_A_1127_155#_c_1766_n 0.0141271f $X=6.195 $Y=0.7
+ $X2=0 $Y2=0
cc_899 N_A_343_417#_c_1453_n N_A_1127_155#_c_1766_n 0.0243368f $X=6.34 $Y=1.745
+ $X2=0 $Y2=0
cc_900 N_A_343_417#_c_1449_n N_A_1127_155#_c_1767_n 0.0643627f $X=6.885 $Y=0.7
+ $X2=0 $Y2=0
cc_901 N_A_343_417#_c_1450_n N_A_1127_155#_c_1767_n 0.0128438f $X=6.195 $Y=0.7
+ $X2=0 $Y2=0
cc_902 N_A_343_417#_c_1449_n N_A_1127_155#_c_1769_n 0.0122839f $X=6.885 $Y=0.7
+ $X2=0 $Y2=0
cc_903 N_A_343_417#_c_1451_n N_A_1127_155#_c_1769_n 0.0126165f $X=6.97 $Y=0.985
+ $X2=0 $Y2=0
cc_904 N_Q_N_c_1587_n N_VGND_c_1615_n 0.0153904f $X=15.575 $Y=0.495 $X2=0 $Y2=0
cc_905 N_Q_N_c_1587_n N_VGND_c_1623_n 0.0220321f $X=15.575 $Y=0.495 $X2=0 $Y2=0
cc_906 N_Q_N_c_1587_n N_VGND_c_1624_n 0.0125808f $X=15.575 $Y=0.495 $X2=0 $Y2=0
cc_907 N_VGND_c_1611_n N_A_1127_155#_c_1767_n 0.107529f $X=7.85 $Y=0 $X2=0 $Y2=0
cc_908 N_VGND_c_1612_n N_A_1127_155#_c_1767_n 0.0116405f $X=8.015 $Y=0.55 $X2=0
+ $Y2=0
cc_909 N_VGND_c_1624_n N_A_1127_155#_c_1767_n 0.0587956f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_910 N_VGND_c_1611_n N_A_1127_155#_c_1768_n 0.0168491f $X=7.85 $Y=0 $X2=0
+ $Y2=0
cc_911 N_VGND_c_1624_n N_A_1127_155#_c_1768_n 0.00867615f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_912 N_VGND_c_1612_n N_A_1127_155#_c_1769_n 0.011903f $X=8.015 $Y=0.55 $X2=0
+ $Y2=0
cc_913 N_VGND_c_1621_n N_A_1859_155#_c_1801_n 0.00370328f $X=11.28 $Y=0 $X2=0
+ $Y2=0
cc_914 N_VGND_c_1624_n N_A_1859_155#_c_1801_n 0.00794602f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_915 N_VGND_c_1613_n N_A_1859_155#_c_1803_n 0.0125556f $X=11.365 $Y=0.43 $X2=0
+ $Y2=0
cc_916 N_VGND_c_1621_n N_A_1859_155#_c_1803_n 0.0215952f $X=11.28 $Y=0 $X2=0
+ $Y2=0
cc_917 N_VGND_c_1624_n N_A_1859_155#_c_1803_n 0.01249f $X=15.6 $Y=0 $X2=0 $Y2=0
