* File: sky130_fd_sc_lp__or4b_lp.pxi.spice
* Created: Wed Sep  2 10:32:49 2020
* 
x_PM_SKY130_FD_SC_LP__OR4B_LP%D_N N_D_N_M1016_g N_D_N_M1006_g N_D_N_M1011_g
+ N_D_N_c_102_n N_D_N_c_106_n D_N D_N N_D_N_c_104_n
+ PM_SKY130_FD_SC_LP__OR4B_LP%D_N
x_PM_SKY130_FD_SC_LP__OR4B_LP%A_27_57# N_A_27_57#_M1016_s N_A_27_57#_M1006_s
+ N_A_27_57#_c_139_n N_A_27_57#_M1017_g N_A_27_57#_c_140_n N_A_27_57#_M1000_g
+ N_A_27_57#_M1005_g N_A_27_57#_c_142_n N_A_27_57#_c_149_n N_A_27_57#_c_143_n
+ N_A_27_57#_c_144_n N_A_27_57#_c_150_n N_A_27_57#_c_145_n N_A_27_57#_c_146_n
+ N_A_27_57#_c_147_n PM_SKY130_FD_SC_LP__OR4B_LP%A_27_57#
x_PM_SKY130_FD_SC_LP__OR4B_LP%C N_C_c_208_n N_C_M1007_g N_C_c_209_n N_C_c_210_n
+ N_C_c_211_n N_C_M1001_g N_C_M1010_g N_C_c_212_n N_C_c_213_n N_C_c_214_n
+ N_C_c_219_n C C C C N_C_c_215_n N_C_c_216_n PM_SKY130_FD_SC_LP__OR4B_LP%C
x_PM_SKY130_FD_SC_LP__OR4B_LP%B N_B_c_269_n N_B_M1012_g N_B_c_270_n N_B_M1008_g
+ N_B_c_271_n N_B_M1013_g N_B_c_272_n N_B_c_278_n B B B B N_B_c_273_n
+ N_B_c_274_n N_B_c_275_n PM_SKY130_FD_SC_LP__OR4B_LP%B
x_PM_SKY130_FD_SC_LP__OR4B_LP%A N_A_M1015_g N_A_c_325_n N_A_M1002_g N_A_c_326_n
+ N_A_c_327_n N_A_M1014_g N_A_c_328_n N_A_c_329_n N_A_c_335_n N_A_c_330_n A A
+ N_A_c_332_n PM_SKY130_FD_SC_LP__OR4B_LP%A
x_PM_SKY130_FD_SC_LP__OR4B_LP%A_311_417# N_A_311_417#_M1000_d
+ N_A_311_417#_M1013_d N_A_311_417#_M1005_s N_A_311_417#_c_399_n
+ N_A_311_417#_M1009_g N_A_311_417#_M1003_g N_A_311_417#_M1004_g
+ N_A_311_417#_c_388_n N_A_311_417#_c_389_n N_A_311_417#_c_401_n
+ N_A_311_417#_c_390_n N_A_311_417#_c_391_n N_A_311_417#_c_392_n
+ N_A_311_417#_c_393_n N_A_311_417#_c_394_n N_A_311_417#_c_395_n
+ N_A_311_417#_c_396_n N_A_311_417#_c_397_n N_A_311_417#_c_398_n
+ PM_SKY130_FD_SC_LP__OR4B_LP%A_311_417#
x_PM_SKY130_FD_SC_LP__OR4B_LP%VPWR N_VPWR_M1006_d N_VPWR_M1015_d N_VPWR_c_498_n
+ N_VPWR_c_499_n VPWR N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_497_n
+ N_VPWR_c_503_n N_VPWR_c_504_n PM_SKY130_FD_SC_LP__OR4B_LP%VPWR
x_PM_SKY130_FD_SC_LP__OR4B_LP%X N_X_M1004_d N_X_M1009_d X X X X X X X X
+ PM_SKY130_FD_SC_LP__OR4B_LP%X
x_PM_SKY130_FD_SC_LP__OR4B_LP%VGND N_VGND_M1011_d N_VGND_M1001_d N_VGND_M1014_d
+ N_VGND_c_573_n N_VGND_c_574_n N_VGND_c_575_n VGND N_VGND_c_576_n
+ N_VGND_c_577_n N_VGND_c_578_n N_VGND_c_579_n N_VGND_c_580_n N_VGND_c_581_n
+ N_VGND_c_582_n N_VGND_c_583_n PM_SKY130_FD_SC_LP__OR4B_LP%VGND
cc_1 VNB N_D_N_M1016_g 0.0400904f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.495
cc_2 VNB N_D_N_M1011_g 0.0313015f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.495
cc_3 VNB N_D_N_c_102_n 0.0201284f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.325
cc_4 VNB D_N 0.00779872f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_D_N_c_104_n 0.0284895f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.34
cc_6 VNB N_A_27_57#_c_139_n 0.0161159f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_7 VNB N_A_27_57#_c_140_n 0.0157384f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.495
cc_8 VNB N_A_27_57#_M1005_g 0.0106128f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.325
cc_9 VNB N_A_27_57#_c_142_n 0.0241735f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_10 VNB N_A_27_57#_c_143_n 0.0164123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_57#_c_144_n 0.0132078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_57#_c_145_n 0.0308667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_57#_c_146_n 0.0141549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_57#_c_147_n 0.102522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C_c_208_n 0.0137701f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.175
cc_16 VNB N_C_c_209_n 0.0102086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_c_210_n 0.00736545f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.845
cc_18 VNB N_C_c_211_n 0.0137578f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_19 VNB N_C_c_212_n 0.00520908f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.325
cc_20 VNB N_C_c_213_n 0.0206661f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.845
cc_21 VNB N_C_c_214_n 0.0136235f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_22 VNB N_C_c_215_n 0.0157593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_c_216_n 0.00761015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_269_n 0.0137578f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.175
cc_25 VNB N_B_c_270_n 0.0166315f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_26 VNB N_B_c_271_n 0.0137701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_c_272_n 0.0216801f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_28 VNB N_B_c_273_n 0.0155054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B_c_274_n 0.00131573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_c_275_n 0.0156712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_c_325_n 0.0137701f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.845
cc_32 VNB N_A_c_326_n 0.0178225f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.495
cc_33 VNB N_A_c_327_n 0.0137578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_c_328_n 0.0237886f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.658
cc_35 VNB N_A_c_329_n 0.0152048f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.845
cc_36 VNB N_A_c_330_n 0.00437176f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_37 VNB A 0.0104474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_c_332_n 0.0143974f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.295
cc_39 VNB N_A_311_417#_M1003_g 0.033346f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.325
cc_40 VNB N_A_311_417#_M1004_g 0.0372181f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_41 VNB N_A_311_417#_c_388_n 0.00408314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_311_417#_c_389_n 0.0302373f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.34
cc_43 VNB N_A_311_417#_c_390_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_311_417#_c_391_n 0.01427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_311_417#_c_392_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_311_417#_c_393_n 0.0185921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_311_417#_c_394_n 5.94059e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_311_417#_c_395_n 0.0282903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_311_417#_c_396_n 0.00846899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_311_417#_c_397_n 0.00184485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_311_417#_c_398_n 0.00964198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VPWR_c_497_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB X 0.022163f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_54 VNB X 0.0477412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_573_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_574_n 0.00409534f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.658
cc_57 VNB N_VGND_c_575_n 0.00420151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_576_n 0.0268803f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.34
cc_59 VNB N_VGND_c_577_n 0.0352526f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.665
cc_60 VNB N_VGND_c_578_n 0.0352526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_579_n 0.0268803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_580_n 0.31529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_581_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_582_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_583_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VPB N_D_N_M1006_g 0.0407681f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_67 VPB N_D_N_c_106_n 0.0208269f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.845
cc_68 VPB D_N 0.00877136f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_69 VPB N_A_27_57#_M1005_g 0.0465616f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.325
cc_70 VPB N_A_27_57#_c_149_n 0.0358412f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.295
cc_71 VPB N_A_27_57#_c_150_n 0.0122316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_27_57#_c_145_n 0.0174289f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_C_M1010_g 0.0239114f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.325
cc_74 VPB N_C_c_214_n 0.00605488f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_75 VPB N_C_c_219_n 0.0118898f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_76 VPB N_C_c_216_n 0.00268803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_B_c_270_n 0.00710684f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_78 VPB N_B_M1008_g 0.0261778f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.495
cc_79 VPB N_B_c_278_n 0.0152661f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_B_c_274_n 0.00179447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_M1015_g 0.0274613f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.495
cc_82 VPB N_A_c_329_n 0.00675768f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.845
cc_83 VPB N_A_c_335_n 0.0124853f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_84 VPB A 0.00963721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A_311_417#_c_399_n 0.0279838f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.495
cc_86 VPB N_A_311_417#_c_388_n 0.0401506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_311_417#_c_401_n 0.018895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_311_417#_c_394_n 0.00315434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_311_417#_c_396_n 0.0141499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_498_n 0.0273066f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.495
cc_91 VPB N_VPWR_c_499_n 0.00314922f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.845
cc_92 VPB N_VPWR_c_500_n 0.0775982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_501_n 0.0328085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_497_n 0.075268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_503_n 0.0243201f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_504_n 0.00518424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB X 0.0228095f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB X 0.07361f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.495
cc_99 N_D_N_M1011_g N_A_27_57#_c_139_n 0.0147173f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_100 N_D_N_M1016_g N_A_27_57#_c_142_n 0.01276f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_101 N_D_N_M1011_g N_A_27_57#_c_142_n 0.00193397f $X=0.845 $Y=0.495 $X2=0
+ $Y2=0
cc_102 N_D_N_M1006_g N_A_27_57#_c_149_n 0.0158047f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_103 N_D_N_M1016_g N_A_27_57#_c_143_n 0.0086968f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_104 N_D_N_M1011_g N_A_27_57#_c_143_n 0.0132923f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_105 N_D_N_c_102_n N_A_27_57#_c_143_n 2.0622e-19 $X=0.665 $Y=1.325 $X2=0 $Y2=0
cc_106 D_N N_A_27_57#_c_143_n 0.0282577f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_107 N_D_N_M1016_g N_A_27_57#_c_144_n 0.00513266f $X=0.485 $Y=0.495 $X2=0
+ $Y2=0
cc_108 N_D_N_M1006_g N_A_27_57#_c_150_n 0.00461335f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_109 N_D_N_c_106_n N_A_27_57#_c_150_n 4.78658e-19 $X=0.597 $Y=1.845 $X2=0
+ $Y2=0
cc_110 N_D_N_M1016_g N_A_27_57#_c_145_n 0.0209089f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_111 N_D_N_M1006_g N_A_27_57#_c_145_n 0.00483231f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_112 D_N N_A_27_57#_c_145_n 0.0486798f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_113 N_D_N_M1011_g N_A_27_57#_c_146_n 0.00178692f $X=0.845 $Y=0.495 $X2=0
+ $Y2=0
cc_114 D_N N_A_27_57#_c_146_n 0.0146608f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_115 N_D_N_M1011_g N_A_27_57#_c_147_n 0.026393f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_116 D_N N_A_27_57#_c_147_n 0.00193857f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_117 N_D_N_c_104_n N_A_27_57#_c_147_n 0.00508474f $X=0.62 $Y=1.34 $X2=0 $Y2=0
cc_118 N_D_N_M1006_g N_VPWR_c_498_n 0.0249766f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_119 N_D_N_c_102_n N_VPWR_c_498_n 0.00255475f $X=0.665 $Y=1.325 $X2=0 $Y2=0
cc_120 N_D_N_c_106_n N_VPWR_c_498_n 8.93004e-19 $X=0.597 $Y=1.845 $X2=0 $Y2=0
cc_121 D_N N_VPWR_c_498_n 0.0161464f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_122 N_D_N_M1006_g N_VPWR_c_497_n 0.014085f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_123 N_D_N_M1006_g N_VPWR_c_503_n 0.00769046f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_124 N_D_N_M1016_g N_VGND_c_573_n 0.00189426f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_125 N_D_N_M1011_g N_VGND_c_573_n 0.0106455f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_126 N_D_N_M1016_g N_VGND_c_576_n 0.00502664f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_127 N_D_N_M1011_g N_VGND_c_576_n 0.00445056f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_128 N_D_N_M1016_g N_VGND_c_580_n 0.00627191f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_129 N_D_N_M1011_g N_VGND_c_580_n 0.0041956f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_130 N_A_27_57#_c_140_n N_C_c_208_n 0.00898204f $X=1.635 $Y=0.825 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_27_57#_c_147_n N_C_c_210_n 0.0121959f $X=1.635 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_27_57#_c_147_n N_C_c_213_n 0.0050162f $X=1.635 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_27_57#_M1005_g N_C_c_219_n 0.0520878f $X=1.985 $Y=2.585 $X2=0 $Y2=0
cc_134 N_A_27_57#_c_147_n N_C_c_215_n 0.0520878f $X=1.635 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_27_57#_M1005_g N_C_c_216_n 0.0446497f $X=1.985 $Y=2.585 $X2=0 $Y2=0
cc_136 N_A_27_57#_c_147_n N_C_c_216_n 0.00557638f $X=1.635 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_27_57#_M1005_g N_A_311_417#_c_401_n 0.0209189f $X=1.985 $Y=2.585
+ $X2=0 $Y2=0
cc_138 N_A_27_57#_c_147_n N_A_311_417#_c_401_n 0.0047532f $X=1.635 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_27_57#_c_139_n N_A_311_417#_c_390_n 0.00193209f $X=1.275 $Y=0.825
+ $X2=0 $Y2=0
cc_140 N_A_27_57#_c_140_n N_A_311_417#_c_390_n 0.0113199f $X=1.635 $Y=0.825
+ $X2=0 $Y2=0
cc_141 N_A_27_57#_c_146_n N_A_311_417#_c_390_n 0.0060622f $X=1.34 $Y=0.99 $X2=0
+ $Y2=0
cc_142 N_A_27_57#_c_147_n N_A_311_417#_c_390_n 0.00226187f $X=1.635 $Y=1.16
+ $X2=0 $Y2=0
cc_143 N_A_27_57#_c_147_n N_A_311_417#_c_391_n 8.20583e-19 $X=1.635 $Y=1.16
+ $X2=0 $Y2=0
cc_144 N_A_27_57#_M1005_g N_A_311_417#_c_396_n 0.0179823f $X=1.985 $Y=2.585
+ $X2=0 $Y2=0
cc_145 N_A_27_57#_c_146_n N_A_311_417#_c_396_n 0.028737f $X=1.34 $Y=0.99 $X2=0
+ $Y2=0
cc_146 N_A_27_57#_c_147_n N_A_311_417#_c_396_n 0.022513f $X=1.635 $Y=1.16 $X2=0
+ $Y2=0
cc_147 N_A_27_57#_c_146_n N_A_311_417#_c_397_n 0.0133354f $X=1.34 $Y=0.99 $X2=0
+ $Y2=0
cc_148 N_A_27_57#_c_147_n N_A_311_417#_c_397_n 0.0122956f $X=1.635 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_27_57#_c_150_n N_VPWR_c_498_n 0.0686502f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_150 N_A_27_57#_M1005_g N_VPWR_c_500_n 0.0087188f $X=1.985 $Y=2.585 $X2=0
+ $Y2=0
cc_151 N_A_27_57#_M1005_g N_VPWR_c_497_n 0.0158312f $X=1.985 $Y=2.585 $X2=0
+ $Y2=0
cc_152 N_A_27_57#_c_149_n N_VPWR_c_497_n 0.0129677f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_153 N_A_27_57#_c_149_n N_VPWR_c_503_n 0.0227064f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_154 N_A_27_57#_c_139_n N_VGND_c_573_n 0.0106445f $X=1.275 $Y=0.825 $X2=0
+ $Y2=0
cc_155 N_A_27_57#_c_140_n N_VGND_c_573_n 0.00189426f $X=1.635 $Y=0.825 $X2=0
+ $Y2=0
cc_156 N_A_27_57#_c_142_n N_VGND_c_573_n 0.0127138f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_157 N_A_27_57#_c_143_n N_VGND_c_573_n 0.0174563f $X=1.175 $Y=0.91 $X2=0 $Y2=0
cc_158 N_A_27_57#_c_146_n N_VGND_c_573_n 0.00278596f $X=1.34 $Y=0.99 $X2=0 $Y2=0
cc_159 N_A_27_57#_c_142_n N_VGND_c_576_n 0.0220321f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_160 N_A_27_57#_c_139_n N_VGND_c_577_n 0.00445056f $X=1.275 $Y=0.825 $X2=0
+ $Y2=0
cc_161 N_A_27_57#_c_140_n N_VGND_c_577_n 0.00502664f $X=1.635 $Y=0.825 $X2=0
+ $Y2=0
cc_162 N_A_27_57#_c_139_n N_VGND_c_580_n 0.0041935f $X=1.275 $Y=0.825 $X2=0
+ $Y2=0
cc_163 N_A_27_57#_c_140_n N_VGND_c_580_n 0.00942073f $X=1.635 $Y=0.825 $X2=0
+ $Y2=0
cc_164 N_A_27_57#_c_142_n N_VGND_c_580_n 0.0125808f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_165 N_A_27_57#_c_143_n N_VGND_c_580_n 0.0152512f $X=1.175 $Y=0.91 $X2=0 $Y2=0
cc_166 N_A_27_57#_c_146_n N_VGND_c_580_n 0.00979814f $X=1.34 $Y=0.99 $X2=0 $Y2=0
cc_167 N_C_c_211_n N_B_c_269_n 0.00982147f $X=2.425 $Y=0.78 $X2=-0.19 $Y2=-0.245
cc_168 N_C_c_214_n N_B_c_270_n 0.0117599f $X=2.515 $Y=1.76 $X2=0 $Y2=0
cc_169 N_C_M1010_g N_B_M1008_g 0.0490778f $X=2.475 $Y=2.585 $X2=0 $Y2=0
cc_170 N_C_c_212_n N_B_c_272_n 0.00982147f $X=2.425 $Y=0.855 $X2=0 $Y2=0
cc_171 N_C_c_219_n N_B_c_278_n 0.0117599f $X=2.515 $Y=1.925 $X2=0 $Y2=0
cc_172 N_C_c_215_n N_B_c_273_n 0.0117599f $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_173 N_C_c_216_n N_B_c_273_n 0.011785f $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_174 N_C_M1010_g N_B_c_274_n 9.4381e-19 $X=2.475 $Y=2.585 $X2=0 $Y2=0
cc_175 N_C_c_215_n N_B_c_274_n 7.18039e-19 $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_176 N_C_c_216_n N_B_c_274_n 0.130418f $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_177 N_C_c_213_n N_B_c_275_n 0.0104403f $X=2.515 $Y=1.255 $X2=0 $Y2=0
cc_178 N_C_M1010_g N_A_311_417#_c_401_n 7.3032e-19 $X=2.475 $Y=2.585 $X2=0 $Y2=0
cc_179 N_C_c_214_n N_A_311_417#_c_401_n 2.87951e-19 $X=2.515 $Y=1.76 $X2=0 $Y2=0
cc_180 N_C_c_219_n N_A_311_417#_c_401_n 2.87951e-19 $X=2.515 $Y=1.925 $X2=0
+ $Y2=0
cc_181 N_C_c_208_n N_A_311_417#_c_390_n 0.00990299f $X=2.065 $Y=0.78 $X2=0 $Y2=0
cc_182 N_C_c_210_n N_A_311_417#_c_390_n 0.00731877f $X=2.14 $Y=0.855 $X2=0 $Y2=0
cc_183 N_C_c_211_n N_A_311_417#_c_390_n 0.00152289f $X=2.425 $Y=0.78 $X2=0 $Y2=0
cc_184 N_C_c_209_n N_A_311_417#_c_391_n 0.0130706f $X=2.35 $Y=0.855 $X2=0 $Y2=0
cc_185 N_C_c_210_n N_A_311_417#_c_391_n 0.00722414f $X=2.14 $Y=0.855 $X2=0 $Y2=0
cc_186 N_C_c_212_n N_A_311_417#_c_391_n 0.0065347f $X=2.425 $Y=0.855 $X2=0 $Y2=0
cc_187 N_C_c_213_n N_A_311_417#_c_391_n 0.00923322f $X=2.515 $Y=1.255 $X2=0
+ $Y2=0
cc_188 N_C_c_215_n N_A_311_417#_c_391_n 0.00123749f $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_189 N_C_c_216_n N_A_311_417#_c_391_n 0.0553395f $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_190 N_C_c_213_n N_A_311_417#_c_396_n 0.00295336f $X=2.515 $Y=1.255 $X2=0
+ $Y2=0
cc_191 N_C_c_215_n N_A_311_417#_c_396_n 4.72993e-19 $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_192 N_C_c_216_n N_A_311_417#_c_396_n 0.122518f $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_193 N_C_c_210_n N_A_311_417#_c_397_n 6.07461e-19 $X=2.14 $Y=0.855 $X2=0 $Y2=0
cc_194 N_C_M1010_g N_VPWR_c_500_n 0.00642983f $X=2.475 $Y=2.585 $X2=0 $Y2=0
cc_195 N_C_c_216_n N_VPWR_c_500_n 0.0193843f $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_196 N_C_M1010_g N_VPWR_c_497_n 0.00814968f $X=2.475 $Y=2.585 $X2=0 $Y2=0
cc_197 N_C_c_216_n N_VPWR_c_497_n 0.0231209f $X=2.515 $Y=1.42 $X2=0 $Y2=0
cc_198 N_C_c_216_n A_422_417# 0.00175001f $X=2.515 $Y=1.42 $X2=-0.19 $Y2=-0.245
cc_199 N_C_c_216_n A_520_417# 0.0085293f $X=2.515 $Y=1.42 $X2=-0.19 $Y2=-0.245
cc_200 N_C_c_208_n N_VGND_c_574_n 0.002112f $X=2.065 $Y=0.78 $X2=0 $Y2=0
cc_201 N_C_c_211_n N_VGND_c_574_n 0.0125337f $X=2.425 $Y=0.78 $X2=0 $Y2=0
cc_202 N_C_c_208_n N_VGND_c_577_n 0.00502664f $X=2.065 $Y=0.78 $X2=0 $Y2=0
cc_203 N_C_c_209_n N_VGND_c_577_n 4.57848e-19 $X=2.35 $Y=0.855 $X2=0 $Y2=0
cc_204 N_C_c_211_n N_VGND_c_577_n 0.00445056f $X=2.425 $Y=0.78 $X2=0 $Y2=0
cc_205 N_C_c_208_n N_VGND_c_580_n 0.00942073f $X=2.065 $Y=0.78 $X2=0 $Y2=0
cc_206 N_C_c_209_n N_VGND_c_580_n 6.33118e-19 $X=2.35 $Y=0.855 $X2=0 $Y2=0
cc_207 N_C_c_211_n N_VGND_c_580_n 0.00796275f $X=2.425 $Y=0.78 $X2=0 $Y2=0
cc_208 N_B_M1008_g N_A_M1015_g 0.0419737f $X=3.045 $Y=2.585 $X2=0 $Y2=0
cc_209 N_B_c_274_n N_A_M1015_g 0.0113269f $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_210 N_B_c_271_n N_A_c_325_n 0.00899044f $X=3.215 $Y=0.78 $X2=0 $Y2=0
cc_211 N_B_c_275_n N_A_c_328_n 0.00375791f $X=3.092 $Y=1.255 $X2=0 $Y2=0
cc_212 N_B_c_270_n N_A_c_329_n 0.0104548f $X=3.092 $Y=1.753 $X2=0 $Y2=0
cc_213 N_B_c_278_n N_A_c_335_n 0.0104548f $X=3.092 $Y=1.925 $X2=0 $Y2=0
cc_214 N_B_c_272_n N_A_c_330_n 0.00899044f $X=3.215 $Y=0.855 $X2=0 $Y2=0
cc_215 N_B_c_273_n A 0.00466156f $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_216 N_B_c_274_n A 0.0465573f $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_217 N_B_c_273_n N_A_c_332_n 0.0104548f $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_218 N_B_c_274_n N_A_c_332_n 7.88709e-19 $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_219 N_B_c_272_n N_A_311_417#_c_391_n 0.0258968f $X=3.215 $Y=0.855 $X2=0 $Y2=0
cc_220 N_B_c_273_n N_A_311_417#_c_391_n 6.37993e-19 $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_221 N_B_c_274_n N_A_311_417#_c_391_n 0.0245914f $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_222 N_B_c_275_n N_A_311_417#_c_391_n 0.00785554f $X=3.092 $Y=1.255 $X2=0
+ $Y2=0
cc_223 N_B_c_269_n N_A_311_417#_c_392_n 0.00152289f $X=2.855 $Y=0.78 $X2=0 $Y2=0
cc_224 N_B_c_271_n N_A_311_417#_c_392_n 0.00990299f $X=3.215 $Y=0.78 $X2=0 $Y2=0
cc_225 N_B_c_272_n N_A_311_417#_c_392_n 0.00731877f $X=3.215 $Y=0.855 $X2=0
+ $Y2=0
cc_226 N_B_c_272_n N_A_311_417#_c_398_n 7.87572e-19 $X=3.215 $Y=0.855 $X2=0
+ $Y2=0
cc_227 N_B_M1008_g N_VPWR_c_499_n 0.00223744f $X=3.045 $Y=2.585 $X2=0 $Y2=0
cc_228 N_B_c_274_n N_VPWR_c_499_n 0.0267958f $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_229 N_B_M1008_g N_VPWR_c_500_n 0.00663182f $X=3.045 $Y=2.585 $X2=0 $Y2=0
cc_230 N_B_c_274_n N_VPWR_c_500_n 0.00916748f $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_231 N_B_M1008_g N_VPWR_c_497_n 0.00900661f $X=3.045 $Y=2.585 $X2=0 $Y2=0
cc_232 N_B_c_274_n N_VPWR_c_497_n 0.0102702f $X=3.1 $Y=1.42 $X2=0 $Y2=0
cc_233 N_B_c_274_n A_634_417# 0.0116888f $X=3.1 $Y=1.42 $X2=-0.19 $Y2=-0.245
cc_234 N_B_c_269_n N_VGND_c_574_n 0.0125337f $X=2.855 $Y=0.78 $X2=0 $Y2=0
cc_235 N_B_c_271_n N_VGND_c_574_n 0.002112f $X=3.215 $Y=0.78 $X2=0 $Y2=0
cc_236 N_B_c_269_n N_VGND_c_578_n 0.00445056f $X=2.855 $Y=0.78 $X2=0 $Y2=0
cc_237 N_B_c_271_n N_VGND_c_578_n 0.00502664f $X=3.215 $Y=0.78 $X2=0 $Y2=0
cc_238 N_B_c_272_n N_VGND_c_578_n 5.84996e-19 $X=3.215 $Y=0.855 $X2=0 $Y2=0
cc_239 N_B_c_269_n N_VGND_c_580_n 0.00796275f $X=2.855 $Y=0.78 $X2=0 $Y2=0
cc_240 N_B_c_271_n N_VGND_c_580_n 0.00942073f $X=3.215 $Y=0.78 $X2=0 $Y2=0
cc_241 N_B_c_272_n N_VGND_c_580_n 7.94744e-19 $X=3.215 $Y=0.855 $X2=0 $Y2=0
cc_242 N_A_c_327_n N_A_311_417#_M1003_g 0.0190109f $X=4.005 $Y=0.78 $X2=0 $Y2=0
cc_243 N_A_c_328_n N_A_311_417#_M1003_g 0.00351016f $X=3.695 $Y=1.255 $X2=0
+ $Y2=0
cc_244 N_A_M1015_g N_A_311_417#_c_388_n 0.028198f $X=3.655 $Y=2.585 $X2=0 $Y2=0
cc_245 N_A_c_335_n N_A_311_417#_c_388_n 0.00897783f $X=3.695 $Y=1.925 $X2=0
+ $Y2=0
cc_246 A N_A_311_417#_c_388_n 0.00861881f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_247 N_A_c_328_n N_A_311_417#_c_389_n 0.00229379f $X=3.695 $Y=1.255 $X2=0
+ $Y2=0
cc_248 A N_A_311_417#_c_389_n 0.006606f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_249 N_A_c_332_n N_A_311_417#_c_389_n 0.0052829f $X=3.695 $Y=1.42 $X2=0 $Y2=0
cc_250 N_A_c_325_n N_A_311_417#_c_392_n 0.00990299f $X=3.645 $Y=0.78 $X2=0 $Y2=0
cc_251 N_A_c_327_n N_A_311_417#_c_392_n 0.00152289f $X=4.005 $Y=0.78 $X2=0 $Y2=0
cc_252 N_A_c_330_n N_A_311_417#_c_392_n 0.00731877f $X=3.645 $Y=0.855 $X2=0
+ $Y2=0
cc_253 N_A_c_326_n N_A_311_417#_c_393_n 0.0209454f $X=3.93 $Y=0.855 $X2=0 $Y2=0
cc_254 N_A_c_328_n N_A_311_417#_c_393_n 0.00626283f $X=3.695 $Y=1.255 $X2=0
+ $Y2=0
cc_255 N_A_c_330_n N_A_311_417#_c_393_n 0.00576469f $X=3.645 $Y=0.855 $X2=0
+ $Y2=0
cc_256 A N_A_311_417#_c_393_n 0.046681f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_257 N_A_c_332_n N_A_311_417#_c_393_n 0.00105893f $X=3.695 $Y=1.42 $X2=0 $Y2=0
cc_258 N_A_c_328_n N_A_311_417#_c_394_n 8.08207e-19 $X=3.695 $Y=1.255 $X2=0
+ $Y2=0
cc_259 A N_A_311_417#_c_394_n 0.0472654f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_260 N_A_c_332_n N_A_311_417#_c_394_n 3.95399e-19 $X=3.695 $Y=1.42 $X2=0 $Y2=0
cc_261 N_A_c_329_n N_A_311_417#_c_395_n 0.0052829f $X=3.695 $Y=1.76 $X2=0 $Y2=0
cc_262 N_A_c_328_n N_A_311_417#_c_398_n 0.00382264f $X=3.695 $Y=1.255 $X2=0
+ $Y2=0
cc_263 N_A_c_330_n N_A_311_417#_c_398_n 3.5619e-19 $X=3.645 $Y=0.855 $X2=0 $Y2=0
cc_264 A N_A_311_417#_c_398_n 0.00943096f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_265 N_A_c_332_n N_A_311_417#_c_398_n 0.00108331f $X=3.695 $Y=1.42 $X2=0 $Y2=0
cc_266 N_A_M1015_g N_VPWR_c_499_n 0.0283968f $X=3.655 $Y=2.585 $X2=0 $Y2=0
cc_267 N_A_c_335_n N_VPWR_c_499_n 0.0019559f $X=3.695 $Y=1.925 $X2=0 $Y2=0
cc_268 A N_VPWR_c_499_n 0.0257274f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_269 N_A_M1015_g N_VPWR_c_500_n 0.00860995f $X=3.655 $Y=2.585 $X2=0 $Y2=0
cc_270 N_A_M1015_g N_VPWR_c_497_n 0.0147029f $X=3.655 $Y=2.585 $X2=0 $Y2=0
cc_271 N_A_M1015_g X 4.97498e-19 $X=3.655 $Y=2.585 $X2=0 $Y2=0
cc_272 N_A_c_325_n N_VGND_c_575_n 0.002112f $X=3.645 $Y=0.78 $X2=0 $Y2=0
cc_273 N_A_c_327_n N_VGND_c_575_n 0.0125337f $X=4.005 $Y=0.78 $X2=0 $Y2=0
cc_274 N_A_c_325_n N_VGND_c_578_n 0.00502664f $X=3.645 $Y=0.78 $X2=0 $Y2=0
cc_275 N_A_c_326_n N_VGND_c_578_n 4.57848e-19 $X=3.93 $Y=0.855 $X2=0 $Y2=0
cc_276 N_A_c_327_n N_VGND_c_578_n 0.00445056f $X=4.005 $Y=0.78 $X2=0 $Y2=0
cc_277 N_A_c_325_n N_VGND_c_580_n 0.00942073f $X=3.645 $Y=0.78 $X2=0 $Y2=0
cc_278 N_A_c_326_n N_VGND_c_580_n 6.33118e-19 $X=3.93 $Y=0.855 $X2=0 $Y2=0
cc_279 N_A_c_327_n N_VGND_c_580_n 0.00796275f $X=4.005 $Y=0.78 $X2=0 $Y2=0
cc_280 N_A_311_417#_c_401_n N_VPWR_c_498_n 0.0364033f $X=1.7 $Y=2.23 $X2=0 $Y2=0
cc_281 N_A_311_417#_c_399_n N_VPWR_c_499_n 0.0140772f $X=4.275 $Y=1.965 $X2=0
+ $Y2=0
cc_282 N_A_311_417#_c_401_n N_VPWR_c_500_n 0.0198001f $X=1.7 $Y=2.23 $X2=0 $Y2=0
cc_283 N_A_311_417#_c_399_n N_VPWR_c_501_n 0.00923064f $X=4.275 $Y=1.965 $X2=0
+ $Y2=0
cc_284 N_A_311_417#_M1005_s N_VPWR_c_497_n 0.00244752f $X=1.555 $Y=2.085 $X2=0
+ $Y2=0
cc_285 N_A_311_417#_c_399_n N_VPWR_c_497_n 0.0176229f $X=4.275 $Y=1.965 $X2=0
+ $Y2=0
cc_286 N_A_311_417#_c_401_n N_VPWR_c_497_n 0.0126002f $X=1.7 $Y=2.23 $X2=0 $Y2=0
cc_287 N_A_311_417#_M1003_g X 0.00125204f $X=4.435 $Y=0.495 $X2=0 $Y2=0
cc_288 N_A_311_417#_M1004_g X 0.0100682f $X=4.795 $Y=0.495 $X2=0 $Y2=0
cc_289 N_A_311_417#_M1004_g X 0.0179112f $X=4.795 $Y=0.495 $X2=0 $Y2=0
cc_290 N_A_311_417#_c_388_n X 0.00586193f $X=4.477 $Y=1.613 $X2=0 $Y2=0
cc_291 N_A_311_417#_c_393_n X 0.012284f $X=4.375 $Y=0.99 $X2=0 $Y2=0
cc_292 N_A_311_417#_c_394_n X 0.0491383f $X=4.54 $Y=1.335 $X2=0 $Y2=0
cc_293 N_A_311_417#_c_395_n X 0.0121155f $X=4.54 $Y=1.335 $X2=0 $Y2=0
cc_294 N_A_311_417#_c_399_n X 0.02367f $X=4.275 $Y=1.965 $X2=0 $Y2=0
cc_295 N_A_311_417#_c_388_n X 0.00230048f $X=4.477 $Y=1.613 $X2=0 $Y2=0
cc_296 N_A_311_417#_c_394_n X 0.0235551f $X=4.54 $Y=1.335 $X2=0 $Y2=0
cc_297 N_A_311_417#_c_390_n N_VGND_c_573_n 0.0127138f $X=1.85 $Y=0.495 $X2=0
+ $Y2=0
cc_298 N_A_311_417#_c_390_n N_VGND_c_574_n 0.0153904f $X=1.85 $Y=0.495 $X2=0
+ $Y2=0
cc_299 N_A_311_417#_c_391_n N_VGND_c_574_n 0.026201f $X=3.265 $Y=0.99 $X2=0
+ $Y2=0
cc_300 N_A_311_417#_c_392_n N_VGND_c_574_n 0.0153904f $X=3.43 $Y=0.495 $X2=0
+ $Y2=0
cc_301 N_A_311_417#_M1003_g N_VGND_c_575_n 0.0125333f $X=4.435 $Y=0.495 $X2=0
+ $Y2=0
cc_302 N_A_311_417#_M1004_g N_VGND_c_575_n 0.002112f $X=4.795 $Y=0.495 $X2=0
+ $Y2=0
cc_303 N_A_311_417#_c_392_n N_VGND_c_575_n 0.0153904f $X=3.43 $Y=0.495 $X2=0
+ $Y2=0
cc_304 N_A_311_417#_c_393_n N_VGND_c_575_n 0.026241f $X=4.375 $Y=0.99 $X2=0
+ $Y2=0
cc_305 N_A_311_417#_c_390_n N_VGND_c_577_n 0.021949f $X=1.85 $Y=0.495 $X2=0
+ $Y2=0
cc_306 N_A_311_417#_c_392_n N_VGND_c_578_n 0.021949f $X=3.43 $Y=0.495 $X2=0
+ $Y2=0
cc_307 N_A_311_417#_M1003_g N_VGND_c_579_n 0.00445056f $X=4.435 $Y=0.495 $X2=0
+ $Y2=0
cc_308 N_A_311_417#_M1004_g N_VGND_c_579_n 0.00502664f $X=4.795 $Y=0.495 $X2=0
+ $Y2=0
cc_309 N_A_311_417#_M1003_g N_VGND_c_580_n 0.00796275f $X=4.435 $Y=0.495 $X2=0
+ $Y2=0
cc_310 N_A_311_417#_M1004_g N_VGND_c_580_n 0.0100553f $X=4.795 $Y=0.495 $X2=0
+ $Y2=0
cc_311 N_A_311_417#_c_390_n N_VGND_c_580_n 0.0124703f $X=1.85 $Y=0.495 $X2=0
+ $Y2=0
cc_312 N_A_311_417#_c_392_n N_VGND_c_580_n 0.0124703f $X=3.43 $Y=0.495 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_497_n A_422_417# 0.00219029f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_314 N_VPWR_c_497_n A_520_417# 0.00851508f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_315 N_VPWR_c_497_n A_634_417# 0.0122504f $X=5.04 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_316 N_VPWR_c_497_n N_X_M1009_d 0.0022865f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_317 N_VPWR_c_499_n X 0.0522413f $X=3.92 $Y=2.27 $X2=0 $Y2=0
cc_318 N_VPWR_c_501_n X 0.0514475f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_319 N_VPWR_c_497_n X 0.0306938f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_320 X N_VGND_c_575_n 0.0153904f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_321 X N_VGND_c_579_n 0.0218834f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_322 X N_VGND_c_580_n 0.0125494f $X=4.955 $Y=0.47 $X2=0 $Y2=0
