* File: sky130_fd_sc_lp__a211o_m.pex.spice
* Created: Wed Sep  2 09:17:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211O_M%A2 3 7 8 11 13
r27 11 14 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.42
+ $X2=1.43 $Y2=1.585
r28 11 13 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.42
+ $X2=1.43 $Y2=1.255
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.415
+ $Y=1.42 $X2=1.415 $Y2=1.42
r30 8 12 8.14393 $w=3.73e-07 $l=2.65e-07 $layer=LI1_cond $X=1.68 $Y=1.397
+ $X2=1.415 $Y2=1.397
r31 7 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.535 $Y=0.935
+ $X2=1.535 $Y2=1.255
r32 3 14 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.465 $Y=2.155
+ $X2=1.465 $Y2=1.585
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_M%A1 1 5 7 13 16 17 20
c39 5 0 9.50458e-20 $X=1.895 $Y=0.935
r40 16 17 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.555 $X2=1.2
+ $Y2=0.925
r41 14 16 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.2 $Y=0.435 $X2=1.2
+ $Y2=0.555
r42 13 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.35 $X2=1.2
+ $Y2=0.435
r43 11 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.085 $Y=0.35
+ $X2=1.085 $Y2=0.26
r44 10 13 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.085 $Y=0.35
+ $X2=1.2 $Y2=0.35
r45 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=0.35 $X2=1.085 $Y2=0.35
r46 5 7 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=1.895 $Y=0.935
+ $X2=1.895 $Y2=2.155
r47 3 5 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.895 $Y=0.335 $X2=1.895
+ $Y2=0.935
r48 2 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=0.26
+ $X2=1.085 $Y2=0.26
r49 1 3 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.82 $Y=0.26
+ $X2=1.895 $Y2=0.335
r50 1 2 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.82 $Y=0.26 $X2=1.25
+ $Y2=0.26
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_M%A_82_483# 1 2 3 10 12 15 17 20 21 22 23 24
+ 30 32 33 34 37 41 46 47
c85 46 0 2.4567e-19 $X=2.48 $Y=2.095
c86 17 0 1.99932e-19 $X=0.9 $Y=2.49
r87 39 41 9.63158 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=1.165
+ $X2=3.06 $Y2=1
r88 35 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=2.095
+ $X2=2.48 $Y2=2.095
r89 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.565 $Y=2.095
+ $X2=2.9 $Y2=2.095
r90 33 39 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.965 $Y=1.25
+ $X2=3.06 $Y2=1.165
r91 33 34 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.965 $Y=1.25
+ $X2=2.565 $Y2=1.25
r92 31 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=2.26
+ $X2=2.48 $Y2=2.095
r93 31 32 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.48 $Y=2.26
+ $X2=2.48 $Y2=2.735
r94 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=1.93
+ $X2=2.48 $Y2=2.095
r95 29 34 5.75414 $w=3.03e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.48 $Y=1.335
+ $X2=2.565 $Y2=1.25
r96 29 44 14.8977 $w=3.03e-07 $l=4.63249e-07 $layer=LI1_cond $X=2.48 $Y=1.335
+ $X2=2.11 $Y2=1.125
r97 29 30 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.48 $Y=1.335
+ $X2=2.48 $Y2=1.93
r98 27 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.11 $Y=2.9 $X2=2.11
+ $Y2=2.81
r99 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=2.9 $X2=2.11 $Y2=2.9
r100 24 32 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.395 $Y=2.9
+ $X2=2.48 $Y2=2.735
r101 24 26 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.395 $Y=2.9
+ $X2=2.11 $Y2=2.9
r102 21 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.945 $Y=2.81
+ $X2=2.11 $Y2=2.81
r103 21 22 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=1.945 $Y=2.81
+ $X2=1.05 $Y2=2.81
r104 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.975 $Y=2.735
+ $X2=1.05 $Y2=2.81
r105 19 20 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.975 $Y=2.565
+ $X2=0.975 $Y2=2.735
r106 18 23 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=0.595 $Y=2.49
+ $X2=0.502 $Y2=2.49
r107 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.9 $Y=2.49
+ $X2=0.975 $Y2=2.565
r108 17 18 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=0.9 $Y=2.49
+ $X2=0.595 $Y2=2.49
r109 13 23 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=0.52 $Y=2.415
+ $X2=0.502 $Y2=2.49
r110 13 15 758.894 $w=1.5e-07 $l=1.48e-06 $layer=POLY_cond $X=0.52 $Y=2.415
+ $X2=0.52 $Y2=0.935
r111 10 23 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=0.485 $Y=2.565
+ $X2=0.502 $Y2=2.49
r112 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.485 $Y=2.565
+ $X2=0.485 $Y2=2.885
r113 3 37 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=1.945 $X2=2.9 $Y2=2.095
r114 2 41 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.91
+ $Y=0.725 $X2=3.05 $Y2=1
r115 1 44 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.725 $X2=2.11 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_M%B1 3 5 7 8 12 16
c37 3 0 2.29908e-19 $X=2.325 $Y=0.935
r38 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.345 $Y=0.43
+ $X2=2.345 $Y2=0.595
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.345
+ $Y=0.43 $X2=2.345 $Y2=0.43
r40 8 13 6.41193 $w=3.52e-07 $l=1.85e-07 $layer=LI1_cond $X=2.16 $Y=0.452
+ $X2=2.345 $Y2=0.452
r41 8 16 3.37992 $w=3.75e-07 $l=1.02e-07 $layer=LI1_cond $X=2.16 $Y=0.452
+ $X2=2.058 $Y2=0.452
r42 7 16 11.6166 $w=3.73e-07 $l=3.78e-07 $layer=LI1_cond $X=1.68 $Y=0.452
+ $X2=2.058 $Y2=0.452
r43 3 5 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.325 $Y=0.935
+ $X2=2.325 $Y2=2.155
r44 3 15 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.325 $Y=0.935
+ $X2=2.325 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_M%C1 3 7 9 15
c25 9 0 1.61086e-19 $X=3.12 $Y=1.665
r26 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.925
+ $Y=1.62 $X2=2.925 $Y2=1.62
r27 13 15 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.835 $Y=1.62
+ $X2=2.925 $Y2=1.62
r28 11 13 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.685 $Y=1.62
+ $X2=2.835 $Y2=1.62
r29 9 16 10.4524 $w=2.13e-07 $l=1.95e-07 $layer=LI1_cond $X=3.12 $Y=1.642
+ $X2=2.925 $Y2=1.642
r30 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.455
+ $X2=2.835 $Y2=1.62
r31 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.835 $Y=1.455
+ $X2=2.835 $Y2=0.935
r32 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.685 $Y=1.785
+ $X2=2.685 $Y2=1.62
r33 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.685 $Y=1.785
+ $X2=2.685 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_M%X 1 2 7 8 9 10 11 12 13
r10 12 13 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.272 $Y=2.405
+ $X2=0.272 $Y2=2.775
r11 11 12 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.272 $Y=2.035
+ $X2=0.272 $Y2=2.405
r12 10 11 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.272 $Y=1.665
+ $X2=0.272 $Y2=2.035
r13 9 10 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.272 $Y=1.295
+ $X2=0.272 $Y2=1.665
r14 8 9 20.8421 $w=2.33e-07 $l=4.25e-07 $layer=LI1_cond $X=0.272 $Y=0.87
+ $X2=0.272 $Y2=1.295
r15 7 8 15.4476 $w=2.33e-07 $l=3.15e-07 $layer=LI1_cond $X=0.272 $Y=0.555
+ $X2=0.272 $Y2=0.87
r16 2 13 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=2.675 $X2=0.27 $Y2=2.82
r17 1 8 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.725 $X2=0.305 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_M%VPWR 1 2 9 13 15 17 22 32 33 36 39
c34 33 0 1.27732e-19 $X=3.12 $Y=3.33
c35 22 0 7.22003e-20 $X=1.515 $Y=3.33
c36 13 0 1.50624e-19 $X=1.68 $Y=2.22
r37 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r41 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 23 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.7 $Y2=3.33
r47 23 25 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 22 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 17 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.7 $Y2=3.33
r53 17 19 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 15 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 15 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=3.33
r58 11 13 35.7956 $w=3.28e-07 $l=1.025e-06 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=2.22
r59 7 36 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=3.33
r60 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=2.95
r61 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.945 $X2=1.68 $Y2=2.22
r62 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=2.675 $X2=0.7 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_M%A_225_389# 1 2 9 11 12 15
c22 15 0 2.09983e-19 $X=2.11 $Y=2.09
r23 13 15 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.12 $Y=1.935
+ $X2=2.12 $Y2=2.09
r24 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.025 $Y=1.85
+ $X2=2.12 $Y2=1.935
r25 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.025 $Y=1.85
+ $X2=1.335 $Y2=1.85
r26 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.24 $Y=1.935
+ $X2=1.335 $Y2=1.85
r27 7 9 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.24 $Y=1.935
+ $X2=1.24 $Y2=2.09
r28 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.945 $X2=2.11 $Y2=2.09
r29 1 9 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.945 $X2=1.25 $Y2=2.09
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_M%VGND 1 2 8 9 12 16 21 23 25 32 33 36 39
r44 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r45 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r47 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 30 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=0 $X2=2.7
+ $Y2=0
r49 30 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.785 $Y=0 $X2=3.12
+ $Y2=0
r50 28 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r51 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 25 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.655
+ $Y2=0
r53 25 27 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.24
+ $Y2=0
r54 23 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r55 23 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r56 19 21 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=2.62 $Y=0.88 $X2=2.7
+ $Y2=0.88
r57 13 16 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=0.655 $Y=0.87
+ $X2=0.735 $Y2=0.87
r58 12 21 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.7 $Y=0.775 $X2=2.7
+ $Y2=0.88
r59 11 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=0.085 $X2=2.7
+ $Y2=0
r60 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.7 $Y=0.085 $X2=2.7
+ $Y2=0.775
r61 10 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.655
+ $Y2=0
r62 9 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.7
+ $Y2=0
r63 9 10 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=2.615 $Y=0 $X2=0.74
+ $Y2=0
r64 8 13 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.655 $Y=0.765
+ $X2=0.655 $Y2=0.87
r65 7 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.655 $Y=0.085
+ $X2=0.655 $Y2=0
r66 7 8 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.655 $Y=0.085
+ $X2=0.655 $Y2=0.765
r67 2 19 182 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.725 $X2=2.62 $Y2=0.88
r68 1 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.725 $X2=0.735 $Y2=0.87
.ends

