* File: sky130_fd_sc_lp__or4_0.pex.spice
* Created: Wed Sep  2 10:31:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4_0%D 3 5 7 9 10 11 12
c29 5 0 1.51728e-19 $X=0.61 $Y=1.51
r30 11 12 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=2.035
r31 10 11 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r32 9 10 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r33 9 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r34 5 18 73.2939 $w=5.41e-07 $l=6.02993e-07 $layer=POLY_cond $X=0.61 $Y=1.51
+ $X2=0.395 $Y2=1.005
r35 5 7 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.61 $Y=1.51 $X2=0.61
+ $Y2=2.62
r36 1 18 43.0019 $w=5.41e-07 $l=2.29783e-07 $layer=POLY_cond $X=0.55 $Y=0.84
+ $X2=0.395 $Y2=1.005
r37 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.55 $Y=0.84 $X2=0.55
+ $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_0%C 3 5 7 11 12 13 17
c34 7 0 4.6452e-20 $X=1.06 $Y=2.62
c35 5 0 1.2302e-19 $X=1.06 $Y=2.17
r36 12 13 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.095 $Y=1.665
+ $X2=1.095 $Y2=2.035
r37 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.06
+ $Y=1.665 $X2=1.06 $Y2=1.665
r38 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.06 $Y=2.005
+ $X2=1.06 $Y2=1.665
r39 10 17 44.4756 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.5
+ $X2=1.06 $Y2=1.665
r40 5 11 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=2.17
+ $X2=1.06 $Y2=2.005
r41 5 7 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.06 $Y=2.17 $X2=1.06
+ $Y2=2.62
r42 3 10 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=0.98 $Y=0.47
+ $X2=0.98 $Y2=1.5
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_0%B 2 5 9 10 11 12 16 18
r46 16 18 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=0.955
+ $X2=1.63 $Y2=0.79
r47 11 12 12.7875 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=1.647 $Y=0.925
+ $X2=1.647 $Y2=1.295
r48 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=0.955 $X2=1.63 $Y2=0.955
r49 9 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.75 $Y=0.47 $X2=1.75
+ $Y2=0.79
r50 5 10 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=1.51 $Y=2.62
+ $X2=1.51 $Y2=1.46
r51 2 10 49.7341 $w=3.9e-07 $l=1.95e-07 $layer=POLY_cond $X=1.63 $Y=1.265
+ $X2=1.63 $Y2=1.46
r52 1 16 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=1.63 $Y=0.985 $X2=1.63
+ $Y2=0.955
r53 1 2 39.929 $w=3.9e-07 $l=2.8e-07 $layer=POLY_cond $X=1.63 $Y=0.985 $X2=1.63
+ $Y2=1.265
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_0%A 3 7 12 16 17 21
r49 16 17 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.142 $Y=1.295
+ $X2=2.142 $Y2=1.665
r50 16 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.2
+ $Y=1.375 $X2=2.2 $Y2=1.375
r51 15 21 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.21 $X2=2.2
+ $Y2=1.375
r52 12 21 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.2 $Y=1.73 $X2=2.2
+ $Y2=1.375
r53 9 12 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.87 $Y=1.805 $X2=2.2
+ $Y2=1.805
r54 7 15 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.18 $Y=0.47 $X2=2.18
+ $Y2=1.21
r55 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.87 $Y=1.88 $X2=1.87
+ $Y2=1.805
r56 1 3 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.87 $Y=1.88 $X2=1.87
+ $Y2=2.62
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_0%A_54_482# 1 2 3 12 16 20 21 22 27 30 32 35 36
+ 37 39 40 41 42 43 45 47 48 52 56 57
c115 37 0 1.69472e-19 $X=1.635 $Y=2.135
r116 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.77
+ $Y=1.025 $X2=2.77 $Y2=1.025
r117 50 52 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.965 $Y=0.47
+ $X2=2.06 $Y2=0.47
r118 46 47 8.91524 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.717 $Y=1.23
+ $X2=0.717 $Y2=1.4
r119 45 57 20.3142 $w=2.93e-07 $l=5.2e-07 $layer=LI1_cond $X=2.612 $Y=2.05
+ $X2=2.612 $Y2=1.53
r120 43 57 6.47318 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.66 $Y=1.335
+ $X2=2.66 $Y2=1.53
r121 42 55 2.51472 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=1.03
+ $X2=2.66 $Y2=0.945
r122 42 43 9.0127 $w=3.88e-07 $l=3.05e-07 $layer=LI1_cond $X=2.66 $Y=1.03
+ $X2=2.66 $Y2=1.335
r123 40 55 5.76906 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.465 $Y=0.945
+ $X2=2.66 $Y2=0.945
r124 40 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.465 $Y=0.945
+ $X2=2.145 $Y2=0.945
r125 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=0.86
+ $X2=2.145 $Y2=0.945
r126 38 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=0.635
+ $X2=2.06 $Y2=0.47
r127 38 39 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.06 $Y=0.635
+ $X2=2.06 $Y2=0.86
r128 36 45 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=2.465 $Y=2.135
+ $X2=2.612 $Y2=2.05
r129 36 37 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.465 $Y=2.135
+ $X2=1.635 $Y2=2.135
r130 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.55 $Y=2.22
+ $X2=1.635 $Y2=2.135
r131 34 35 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.55 $Y=2.22
+ $X2=1.55 $Y2=2.43
r132 33 48 2.79095 $w=3.42e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.607
+ $X2=0.62 $Y2=2.607
r133 32 35 7.97992 $w=3.55e-07 $l=2.15346e-07 $layer=LI1_cond $X=1.465 $Y=2.607
+ $X2=1.55 $Y2=2.43
r134 32 33 24.672 $w=3.53e-07 $l=7.6e-07 $layer=LI1_cond $X=1.465 $Y=2.607
+ $X2=0.705 $Y2=2.607
r135 30 46 33.6868 $w=2.58e-07 $l=7.6e-07 $layer=LI1_cond $X=0.77 $Y=0.47
+ $X2=0.77 $Y2=1.23
r136 27 48 3.95098 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=0.62 $Y=2.43
+ $X2=0.62 $Y2=2.607
r137 27 47 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.62 $Y=2.43
+ $X2=0.62 $Y2=1.4
r138 22 48 2.79095 $w=3.42e-07 $l=9.12688e-08 $layer=LI1_cond $X=0.535 $Y=2.62
+ $X2=0.62 $Y2=2.607
r139 22 24 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.535 $Y=2.62
+ $X2=0.395 $Y2=2.62
r140 20 56 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.77 $Y=1.365
+ $X2=2.77 $Y2=1.025
r141 20 21 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.365
+ $X2=2.77 $Y2=1.53
r142 19 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=0.86
+ $X2=2.77 $Y2=1.025
r143 16 21 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=2.705 $Y=2.73
+ $X2=2.705 $Y2=1.53
r144 12 19 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.68 $Y=0.47
+ $X2=2.68 $Y2=0.86
r145 3 24 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.27
+ $Y=2.41 $X2=0.395 $Y2=2.62
r146 2 50 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.26 $X2=1.965 $Y2=0.47
r147 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.26 $X2=0.765 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_0%VPWR 1 6 8 10 20 21 24
r30 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r33 18 24 13.5049 $w=1.7e-07 $l=3.43e-07 $layer=LI1_cond $X=2.605 $Y=3.33
+ $X2=2.262 $Y2=3.33
r34 18 20 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.605 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 10 24 13.5049 $w=1.7e-07 $l=3.42e-07 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=2.262 $Y2=3.33
r38 10 16 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 8 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 4 24 2.81621 $w=6.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.262 $Y=3.245
+ $X2=2.262 $Y2=3.33
r43 4 6 12.0481 $w=6.83e-07 $l=6.9e-07 $layer=LI1_cond $X=2.262 $Y=3.245
+ $X2=2.262 $Y2=2.555
r44 1 6 200 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_PDIFF $count=3 $X=1.945
+ $Y=2.41 $X2=2.47 $Y2=2.555
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_0%X 1 2 7 8 9 10 11 12 13 40 43
r19 43 44 3.34702 $w=4.98e-07 $l=1.5e-08 $layer=LI1_cond $X=3.025 $Y=2.405
+ $X2=3.025 $Y2=2.39
r20 23 40 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=0.635
+ $X2=3.15 $Y2=0.47
r21 13 47 5.26274 $w=4.98e-07 $l=2.2e-07 $layer=LI1_cond $X=3.025 $Y=2.775
+ $X2=3.025 $Y2=2.555
r22 12 47 2.75098 $w=4.98e-07 $l=1.15e-07 $layer=LI1_cond $X=3.025 $Y=2.44
+ $X2=3.025 $Y2=2.555
r23 12 43 0.837255 $w=4.98e-07 $l=3.5e-08 $layer=LI1_cond $X=3.025 $Y=2.44
+ $X2=3.025 $Y2=2.405
r24 12 44 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=3.15 $Y=2.355
+ $X2=3.15 $Y2=2.39
r25 11 12 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=3.15 $Y=2.035
+ $X2=3.15 $Y2=2.355
r26 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.15 $Y=1.665
+ $X2=3.15 $Y2=2.035
r27 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.15 $Y=1.295
+ $X2=3.15 $Y2=1.665
r28 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.15 $Y=0.925 $X2=3.15
+ $Y2=1.295
r29 7 40 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=3.12 $Y=0.47 $X2=3.15
+ $Y2=0.47
r30 7 36 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.12 $Y=0.47
+ $X2=2.895 $Y2=0.47
r31 7 8 13.2761 $w=2.48e-07 $l=2.88e-07 $layer=LI1_cond $X=3.15 $Y=0.637
+ $X2=3.15 $Y2=0.925
r32 7 23 0.0921954 $w=2.48e-07 $l=2e-09 $layer=LI1_cond $X=3.15 $Y=0.637
+ $X2=3.15 $Y2=0.635
r33 2 47 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.78
+ $Y=2.41 $X2=2.92 $Y2=2.555
r34 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.26 $X2=2.895 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_0%VGND 1 2 3 10 12 16 19 20 21 23 33 34
c40 34 0 1.51728e-19 $X=3.12 $Y=0
r41 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r42 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r45 28 30 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.665 $Y=0 $X2=2.16
+ $Y2=0
r46 27 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r47 27 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r48 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 24 37 4.36211 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.235
+ $Y2=0
r50 24 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.72
+ $Y2=0
r51 23 44 9.60952 $w=5.83e-07 $l=4.7e-07 $layer=LI1_cond $X=1.372 $Y=0 $X2=1.372
+ $Y2=0.47
r52 23 28 8.15384 $w=1.7e-07 $l=2.93e-07 $layer=LI1_cond $X=1.372 $Y=0 $X2=1.665
+ $Y2=0
r53 23 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 23 26 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=0.72
+ $Y2=0
r55 21 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r56 21 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r57 19 30 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.16
+ $Y2=0
r58 19 20 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.452
+ $Y2=0
r59 18 33 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=3.12
+ $Y2=0
r60 18 20 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.452
+ $Y2=0
r61 14 20 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.452 $Y=0.085
+ $X2=2.452 $Y2=0
r62 14 16 16.1342 $w=2.73e-07 $l=3.85e-07 $layer=LI1_cond $X=2.452 $Y=0.085
+ $X2=2.452 $Y2=0.47
r63 10 37 3.15557 $w=3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.235 $Y2=0
r64 10 12 14.7897 $w=2.98e-07 $l=3.85e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.32 $Y2=0.47
r65 3 16 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=2.255
+ $Y=0.26 $X2=2.44 $Y2=0.47
r66 2 44 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=1.055
+ $Y=0.26 $X2=1.535 $Y2=0.47
r67 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.21
+ $Y=0.26 $X2=0.335 $Y2=0.47
.ends

