* File: sky130_fd_sc_lp__o311a_lp.spice
* Created: Wed Sep  2 10:23:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o311a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o311a_lp  VNB VPB A1 A2 A3 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1001 A_114_141# N_A_84_115#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_84_115#_M1011_g A_114_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.05985 AS=0.0441 PD=0.705 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1006 N_A_273_141#_M1006_d N_A1_M1006_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.05985 PD=0.7 PS=0.705 NRD=0 NRS=1.428 M=1 R=2.8 SA=75001
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_273_141#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.0588 PD=0.86 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_273_141#_M1007_d N_A3_M1007_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0924 PD=0.7 PS=0.86 NRD=0 NRS=22.848 M=1 R=2.8 SA=75002
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_563_141# N_B1_M1008_g N_A_273_141#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_84_115#_M1004_d N_C1_M1004_g A_563_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_84_115#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.25 W=1
+ AD=0.1775 AS=0.285 PD=1.355 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1012 A_258_419# N_A1_M1012_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.1775 PD=1.24 PS=1.355 NRD=12.7853 NRS=14.7553 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1003 A_356_419# N_A2_M1003_g A_258_419# VPB PHIGHVT L=0.25 W=1 AD=0.145
+ AS=0.12 PD=1.29 PS=1.24 NRD=17.7103 NRS=12.7853 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1010 N_A_84_115#_M1010_d N_A3_M1010_g A_356_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0 NRS=17.7103 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_A_84_115#_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0 NRS=1.9503 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1005 N_A_84_115#_M1005_d N_C1_M1005_g N_VPWR_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.145 PD=2.57 PS=1.29 NRD=0 NRS=1.9503 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o311a_lp.pxi.spice"
*
.ends
*
*
