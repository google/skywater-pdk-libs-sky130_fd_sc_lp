* NGSPICE file created from sky130_fd_sc_lp__a2111oi_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2111oi_lp A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_289_57# B1 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.444e+11p ps=4.16e+06u
M1001 a_553_47# C1 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1002 a_711_47# D1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.507e+11p ps=4.19e+06u
M1003 VGND D1 a_711_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_539_409# B1 a_131_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=5.65e+11p ps=5.13e+06u
M1005 VGND A2 a_125_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_131_409# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.55e+11p ps=5.11e+06u
M1007 a_637_409# C1 a_539_409# VPB phighvt w=1e+06u l=250000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
M1008 a_125_57# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_289_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C1 a_553_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y D1 a_637_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1012 VPWR A2 a_131_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

