* File: sky130_fd_sc_lp__a21oi_1.spice
* Created: Fri Aug 28 09:51:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a21oi_1  VNB VPB A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1002 A_110_69# N_A2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.2226 PD=1.08 PS=2.21 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2 SB=75001.1
+ A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g A_110_69# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.1008 PD=1.23 PS=1.08 NRD=9.996 NRS=9.276 M=1 R=5.6 SA=75000.6 SB=75000.8
+ A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2436 AS=0.1638 PD=2.26 PS=1.23 NRD=3.564 NRS=5.712 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_27_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.3339 PD=1.61 PS=3.05 NRD=5.4569 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_A_27_367#_M1004_d N_A1_M1004_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2205 PD=1.54 PS=1.61 NRD=0 NRS=5.4569 M=1 R=8.4 SA=75000.7
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_27_367#_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.2895 P=8.33
*
.include "sky130_fd_sc_lp__a21oi_1.pxi.spice"
*
.ends
*
*
