* NGSPICE file created from sky130_fd_sc_lp__a211o_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_303_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.497e+11p pd=6.23e+06u as=1.1592e+12p ps=9.4e+06u
M1001 a_80_21# C1 VGND VNB nshort w=840000u l=150000u
+  ad=6.426e+11p pd=4.89e+06u as=1.1298e+12p ps=7.73e+06u
M1002 X a_80_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1003 VPWR a_80_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1004 VGND a_80_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_386_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1006 a_80_21# C1 a_590_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=3.402e+11p ps=3.06e+06u
M1007 a_80_21# A1 a_386_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_590_367# B1 a_303_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_303_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B1 a_80_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_80_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

