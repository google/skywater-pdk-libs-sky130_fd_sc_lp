* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__srsdfxtp_1 CLK D SCD SCE SLEEP_B KAPWR VGND VNB VPB VPWR
+ Q
X0 a_786_139# a_540_21# a_1010_530# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1010_530# a_914_245# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_786_139# a_914_245# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_1247_69# a_570_47# a_1319_69# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 VGND a_2504_57# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_210_47# D a_282_477# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_282_477# SCE a_396_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 KAPWR SLEEP_B a_540_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_914_245# a_540_21# a_1372_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_1372_379# a_540_21# a_1319_69# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 a_786_139# a_570_47# a_872_139# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND a_31_477# a_210_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1704_125# a_1319_69# a_1493_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_2504_57# a_1319_69# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_368_477# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 VPWR a_540_21# a_570_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_2321_178# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_282_477# a_31_477# a_368_477# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_204_477# D a_282_477# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 VGND a_1319_69# a_1704_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 KAPWR a_1319_69# a_1493_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 a_872_139# a_914_245# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR a_786_139# a_914_245# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 a_1319_69# a_540_21# a_1451_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_540_21# CLK KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_2243_178# SLEEP_B a_2321_178# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1523_113# a_1493_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_31_477# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 VGND a_540_21# a_570_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1319_69# a_570_47# a_1858_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X30 a_282_477# a_570_47# a_786_139# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_540_21# CLK a_2243_178# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VPWR SCE a_204_477# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 a_396_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1451_113# a_1493_21# a_1523_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1858_419# a_1493_21# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X36 a_31_477# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_282_477# a_540_21# a_786_139# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_914_245# a_570_47# a_1247_69# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X39 VPWR a_2504_57# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X40 a_2504_57# a_1319_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
