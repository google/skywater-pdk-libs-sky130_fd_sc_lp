* File: sky130_fd_sc_lp__sdfsbp_1.spice
* Created: Wed Sep  2 10:35:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfsbp_1.pex.spice"
.subckt sky130_fd_sc_lp__sdfsbp_1  VNB VPB SCE D SCD CLK SET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_SCE_M1013_g N_A_34_481#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1032 A_252_47# N_A_34_481#_M1032_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1014 N_A_275_481#_M1014_d N_D_M1014_g A_252_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0441 PD=1.04 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 A_478_47# N_SCE_M1006_g N_A_275_481#_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.1302 PD=0.695 PS=1.04 NRD=23.568 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_SCD_M1036_g A_478_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.05775 PD=0.7 PS=0.695 NRD=0 NRS=23.568 M=1 R=2.8 SA=75002.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1023 N_A_640_481#_M1023_d N_CLK_M1023_g N_VGND_M1036_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 N_A_901_441#_M1026_d N_A_640_481#_M1026_g N_VGND_M1026_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_A_1146_463#_M1024_d N_A_640_481#_M1024_g N_A_275_481#_M1024_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1025 A_1245_119# N_A_901_441#_M1025_g N_A_1146_463#_M1024_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_1274_401#_M1015_g A_1245_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_1575_119# N_A_1146_463#_M1005_g N_A_1274_401#_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1041 N_VGND_M1041_d N_SET_B_M1041_g A_1575_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.167128 AS=0.0441 PD=1.18472 PS=0.63 NRD=164.28 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1029 A_1848_119# N_A_1146_463#_M1029_g N_VGND_M1041_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.254672 PD=0.85 PS=1.80528 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1038 N_A_1920_119#_M1038_d N_A_901_441#_M1038_g A_1848_119# VNB NSHORT L=0.15
+ W=0.64 AD=0.130717 AS=0.0672 PD=1.2317 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75001.5 SB=75001 A=0.096 P=1.58 MULT=1
MM1030 A_2025_118# N_A_640_481#_M1030_g N_A_1920_119#_M1038_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.085783 PD=0.63 PS=0.808302 NRD=14.28 NRS=27.132 M=1
+ R=2.8 SA=75002.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1035 A_2097_118# N_A_2067_92#_M1035_g A_2025_118# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75002.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_SET_B_M1028_g A_2097_118# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_A_1920_119#_M1033_g N_A_2067_92#_M1033_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1827 AS=0.1113 PD=1.29 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_2582_150#_M1002_d N_A_1920_119#_M1002_g N_VGND_M1033_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1827 PD=1.37 PS=1.29 NRD=0 NRS=71.424 M=1 R=2.8
+ SA=75001.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_2582_150#_M1020_g N_Q_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.20075 AS=0.2394 PD=1.39 PS=2.25 NRD=12.132 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1021 N_Q_N_M1021_d N_A_1920_119#_M1021_g N_VGND_M1020_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.20075 PD=2.21 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 N_VPWR_M1022_d N_SCE_M1022_g N_A_34_481#_M1022_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1034 A_203_481# N_SCE_M1034_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1039 N_A_275_481#_M1039_d N_D_M1039_g A_203_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=33.8446 NRS=15.3857 M=1 R=4.26667
+ SA=75001 SB=75002 A=0.096 P=1.58 MULT=1
MM1008 A_383_481# N_A_34_481#_M1008_g N_A_275_481#_M1039_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0672 AS=0.1248 PD=0.85 PS=1.03 NRD=15.3857 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1011_d N_SCD_M1011_g A_383_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.248 AS=0.0672 PD=1.415 PS=0.85 NRD=47.6937 NRS=15.3857 M=1 R=4.26667
+ SA=75001.9 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_A_640_481#_M1009_d N_CLK_M1009_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.248 PD=1.81 PS=1.415 NRD=0 NRS=104.646 M=1 R=4.26667
+ SA=75002.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_901_441#_M1017_d N_A_640_481#_M1017_g N_VPWR_M1017_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.3179 PD=1.81 PS=2.7 NRD=0 NRS=135.95 M=1
+ R=4.26667 SA=75000.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_A_1146_463#_M1018_d N_A_901_441#_M1018_g N_A_275_481#_M1018_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75005.3 A=0.063 P=1.14 MULT=1
MM1000 A_1232_463# N_A_640_481#_M1000_g N_A_1146_463#_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75004.9 A=0.063 P=1.14 MULT=1
MM1031 N_VPWR_M1031_d N_A_1274_401#_M1031_g A_1232_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.10605 AS=0.0441 PD=0.925 PS=0.63 NRD=4.6886 NRS=23.443 M=1 R=2.8
+ SA=75001 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1004 N_A_1274_401#_M1004_d N_A_1146_463#_M1004_g N_VPWR_M1031_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.10605 PD=0.7 PS=0.925 NRD=0 NRS=100.844 M=1 R=2.8
+ SA=75001.6 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_SET_B_M1010_g N_A_1274_401#_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.271275 AS=0.0588 PD=1.53333 PS=0.7 NRD=39.8531 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1019 A_1818_379# N_A_1146_463#_M1019_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.15995 AS=0.54255 PD=1.325 PS=3.06667 NRD=31.7564 NRS=19.9167 M=1
+ R=5.6 SA=75001.9 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1040 N_A_1920_119#_M1040_d N_A_640_481#_M1040_g A_1818_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1792 AS=0.15995 PD=1.62 PS=1.325 NRD=5.8509 NRS=31.7564 M=1 R=5.6
+ SA=75002.3 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1012 A_2025_488# N_A_901_441#_M1012_g N_A_1920_119#_M1040_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0896 PD=0.63 PS=0.81 NRD=23.443 NRS=21.0987 M=1 R=2.8
+ SA=75003.4 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_2067_92#_M1001_g A_2025_488# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.15015 AS=0.0441 PD=1.135 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75003.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_A_1920_119#_M1003_d N_SET_B_M1003_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.15015 PD=1.37 PS=1.135 NRD=0 NRS=0 M=1 R=2.8 SA=75004.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_VPWR_M1016_d N_A_1920_119#_M1016_g N_A_2067_92#_M1016_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.126277 AS=0.1113 PD=0.998491 PS=1.37 NRD=160.634 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1037 N_A_2582_150#_M1037_d N_A_1920_119#_M1037_g N_VPWR_M1016_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.192423 PD=1.81 PS=1.52151 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1027 N_VPWR_M1027_d N_A_2582_150#_M1027_g N_Q_M1027_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1007 N_Q_N_M1007_d N_A_1920_119#_M1007_g N_VPWR_M1027_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX42_noxref VNB VPB NWDIODE A=29.3551 P=35.21
c_146 VNB 0 2.12464e-19 $X=0 $Y=0
c_284 VPB 0 1.71354e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfsbp_1.pxi.spice"
*
.ends
*
*
