* File: sky130_fd_sc_lp__a41o_m.pex.spice
* Created: Wed Sep  2 09:29:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41O_M%A_80_153# 1 2 10 13 15 17 20 22 26 27 28 29
+ 30 31 34 38 41
r69 36 38 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=1.32 $Y=0.775
+ $X2=1.32 $Y2=0.51
r70 32 34 6.33766 $w=2.08e-07 $l=1.2e-07 $layer=LI1_cond $X=1.21 $Y=2.565
+ $X2=1.21 $Y2=2.685
r71 30 32 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.105 $Y=2.48
+ $X2=1.21 $Y2=2.565
r72 30 31 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.105 $Y=2.48
+ $X2=0.695 $Y2=2.48
r73 28 36 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.225 $Y=0.86
+ $X2=1.32 $Y2=0.775
r74 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.225 $Y=0.86
+ $X2=0.695 $Y2=0.86
r75 27 41 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=2.01
+ $X2=0.587 $Y2=1.845
r76 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=2.01 $X2=0.61 $Y2=2.01
r77 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=2.395
+ $X2=0.695 $Y2=2.48
r78 24 26 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.61 $Y=2.395
+ $X2=0.61 $Y2=2.01
r79 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.945
+ $X2=0.695 $Y2=0.86
r80 23 26 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=0.61 $Y=0.945
+ $X2=0.61 $Y2=2.01
r81 18 20 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.475 $Y=0.84
+ $X2=0.685 $Y2=0.84
r82 15 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.685 $Y=0.765
+ $X2=0.685 $Y2=0.84
r83 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.685 $Y=0.765
+ $X2=0.685 $Y2=0.445
r84 13 22 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.475 $Y=2.885
+ $X2=0.475 $Y2=2.515
r85 10 22 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.587 $Y=2.328
+ $X2=0.587 $Y2=2.515
r86 9 27 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.587 $Y=2.032
+ $X2=0.587 $Y2=2.01
r87 9 10 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.587 $Y=2.032
+ $X2=0.587 $Y2=2.328
r88 7 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=0.915
+ $X2=0.475 $Y2=0.84
r89 7 41 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=0.475 $Y=0.915
+ $X2=0.475 $Y2=1.845
r90 2 34 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=2.54 $X2=1.21 $Y2=2.685
r91 1 38 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.19
+ $Y=0.235 $X2=1.33 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_M%B1 3 7 12 14 16 17 18 23
r50 17 18 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.665
+ $X2=1.175 $Y2=2.035
r51 17 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.71 $X2=1.15 $Y2=1.71
r52 16 17 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.295
+ $X2=1.175 $Y2=1.665
r53 12 23 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.15 $Y=2.065
+ $X2=1.15 $Y2=1.71
r54 12 14 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=1.15 $Y=2.14
+ $X2=1.425 $Y2=2.14
r55 10 23 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.545
+ $X2=1.15 $Y2=1.71
r56 5 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=2.215
+ $X2=1.425 $Y2=2.14
r57 5 7 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.425 $Y=2.215
+ $X2=1.425 $Y2=2.75
r58 3 10 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=1.115 $Y=0.445
+ $X2=1.115 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_M%A1 3 7 12 13 14 15 16 17 18 25
r52 17 18 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=2.035
r53 16 17 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.295
+ $X2=1.685 $Y2=1.665
r54 16 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.32 $X2=1.69 $Y2=1.32
r55 15 16 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=0.925
+ $X2=1.685 $Y2=1.295
r56 14 15 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=0.555
+ $X2=1.685 $Y2=0.925
r57 12 25 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.69 $Y=1.675
+ $X2=1.69 $Y2=1.32
r58 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.727 $Y=1.675
+ $X2=1.727 $Y2=1.825
r59 10 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.155
+ $X2=1.69 $Y2=1.32
r60 7 13 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.855 $Y=2.75
+ $X2=1.855 $Y2=1.825
r61 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.6 $Y=0.445 $X2=1.6
+ $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_M%A2 3 6 9 10 11 12 13 14 15 16 23
r45 15 16 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=2.035
r46 14 15 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=1.295
+ $X2=2.195 $Y2=1.665
r47 13 14 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=0.925
+ $X2=2.195 $Y2=1.295
r48 13 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23
+ $Y=0.93 $X2=2.23 $Y2=0.93
r49 12 13 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=0.555
+ $X2=2.195 $Y2=0.925
r50 10 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.23 $Y=1.27
+ $X2=2.23 $Y2=0.93
r51 10 11 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.27
+ $X2=2.23 $Y2=1.435
r52 9 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=0.765
+ $X2=2.23 $Y2=0.93
r53 6 11 674.287 $w=1.5e-07 $l=1.315e-06 $layer=POLY_cond $X=2.285 $Y=2.75
+ $X2=2.285 $Y2=1.435
r54 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.14 $Y=0.445 $X2=2.14
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_M%A3 3 7 11 12 13 14 15 16 22
r46 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.77
+ $Y=1.395 $X2=2.77 $Y2=1.395
r47 15 16 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.705 $Y=1.665
+ $X2=2.705 $Y2=2.035
r48 15 23 10.372 $w=2.98e-07 $l=2.7e-07 $layer=LI1_cond $X=2.705 $Y=1.665
+ $X2=2.705 $Y2=1.395
r49 14 23 3.84148 $w=2.98e-07 $l=1e-07 $layer=LI1_cond $X=2.705 $Y=1.295
+ $X2=2.705 $Y2=1.395
r50 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.705 $Y=0.925
+ $X2=2.705 $Y2=1.295
r51 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.77 $Y=1.735
+ $X2=2.77 $Y2=1.395
r52 11 12 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.735
+ $X2=2.77 $Y2=1.9
r53 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.23
+ $X2=2.77 $Y2=1.395
r54 7 12 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=2.715 $Y=2.75
+ $X2=2.715 $Y2=1.9
r55 3 10 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.68 $Y=0.445
+ $X2=2.68 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_M%A4 3 7 10 14 18 21 22 23 24 25 31
r37 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.43
+ $Y=1.005 $X2=3.43 $Y2=1.005
r38 24 25 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.515 $Y=1.665
+ $X2=3.515 $Y2=2.035
r39 23 24 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.515 $Y=1.295
+ $X2=3.515 $Y2=1.665
r40 23 32 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=3.515 $Y=1.295
+ $X2=3.515 $Y2=1.005
r41 22 32 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=3.515 $Y=0.925
+ $X2=3.515 $Y2=1.005
r42 20 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.43 $Y=1.345
+ $X2=3.43 $Y2=1.005
r43 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.345
+ $X2=3.43 $Y2=1.51
r44 16 18 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.145 $Y=2.215
+ $X2=3.34 $Y2=2.215
r45 14 31 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.43 $Y=0.99
+ $X2=3.43 $Y2=1.005
r46 11 14 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.04 $Y=0.915
+ $X2=3.43 $Y2=0.915
r47 10 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.34 $Y=2.14
+ $X2=3.34 $Y2=2.215
r48 10 21 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.34 $Y=2.14
+ $X2=3.34 $Y2=1.51
r49 5 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.145 $Y=2.29
+ $X2=3.145 $Y2=2.215
r50 5 7 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.145 $Y=2.29
+ $X2=3.145 $Y2=2.75
r51 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.04 $Y=0.84 $X2=3.04
+ $Y2=0.915
r52 1 3 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.04 $Y=0.84 $X2=3.04
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_M%X 1 2 7 8 9 10 11 12 13 43
r16 41 43 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.25 $Y=0.43
+ $X2=0.47 $Y2=0.43
r17 22 41 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.25 $Y=0.595
+ $X2=0.25 $Y2=0.43
r18 12 13 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=2.405
+ $X2=0.25 $Y2=2.775
r19 11 12 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=2.035
+ $X2=0.25 $Y2=2.405
r20 10 11 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.665
+ $X2=0.25 $Y2=2.035
r21 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.665
r22 8 9 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=0.925 $X2=0.25
+ $Y2=1.295
r23 7 41 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=0.43 $X2=0.25
+ $Y2=0.43
r24 7 8 17.9789 $w=1.88e-07 $l=3.08e-07 $layer=LI1_cond $X=0.25 $Y=0.617
+ $X2=0.25 $Y2=0.925
r25 7 22 1.28421 $w=1.88e-07 $l=2.2e-08 $layer=LI1_cond $X=0.25 $Y=0.617
+ $X2=0.25 $Y2=0.595
r26 2 13 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.675 $X2=0.26 $Y2=2.82
r27 1 43 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.345
+ $Y=0.235 $X2=0.47 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_M%VPWR 1 2 3 12 16 20 23 24 26 27 28 30 43 44
+ 47
r53 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 38 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 35 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r60 35 37 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 33 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 30 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r64 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r65 28 41 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 28 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 26 40 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 26 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.93 $Y2=3.33
r69 25 43 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=3.6 $Y2=3.33
r70 25 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=2.93 $Y2=3.33
r71 23 37 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.07 $Y2=3.33
r73 22 40 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.64 $Y2=3.33
r74 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.07 $Y2=3.33
r75 18 27 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=3.245
+ $X2=2.93 $Y2=3.33
r76 18 20 22.71 $w=2.08e-07 $l=4.3e-07 $layer=LI1_cond $X=2.93 $Y=3.245 $X2=2.93
+ $Y2=2.815
r77 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=3.33
r78 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=2.815
r79 10 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r80 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.95
r81 3 20 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=2.54 $X2=2.93 $Y2=2.815
r82 2 16 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=2.54 $X2=2.07 $Y2=2.815
r83 1 12 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.675 $X2=0.69 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_M%A_300_508# 1 2 3 12 14 15 18 20 24 26
r39 22 24 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=3.36 $Y=2.47
+ $X2=3.36 $Y2=2.685
r40 21 26 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.605 $Y=2.385
+ $X2=2.51 $Y2=2.385
r41 20 22 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.255 $Y=2.385
+ $X2=3.36 $Y2=2.47
r42 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.255 $Y=2.385
+ $X2=2.605 $Y2=2.385
r43 16 26 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=2.47
+ $X2=2.51 $Y2=2.385
r44 16 18 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=2.51 $Y=2.47
+ $X2=2.51 $Y2=2.685
r45 14 26 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.415 $Y=2.385
+ $X2=2.51 $Y2=2.385
r46 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.415 $Y=2.385
+ $X2=1.725 $Y2=2.385
r47 10 15 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.63 $Y=2.47
+ $X2=1.725 $Y2=2.385
r48 10 12 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=1.63 $Y=2.47
+ $X2=1.63 $Y2=2.685
r49 3 24 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.22
+ $Y=2.54 $X2=3.36 $Y2=2.685
r50 2 18 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=2.54 $X2=2.5 $Y2=2.685
r51 1 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=2.54 $X2=1.64 $Y2=2.685
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_M%VGND 1 2 9 13 16 17 18 24 30 31 34
r48 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r50 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.255
+ $Y2=0
r52 28 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.6
+ $Y2=0
r53 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=3.255
+ $Y2=0
r55 24 26 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=3.09 $Y=0 $X2=1.2
+ $Y2=0
r56 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r57 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 18 35 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r59 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r60 16 21 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.72
+ $Y2=0
r61 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.9
+ $Y2=0
r62 15 26 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.2
+ $Y2=0
r63 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.9
+ $Y2=0
r64 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.255 $Y=0.085
+ $X2=3.255 $Y2=0
r65 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.255 $Y=0.085
+ $X2=3.255 $Y2=0.38
r66 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=0.085 $X2=0.9
+ $Y2=0
r67 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.9 $Y=0.085 $X2=0.9
+ $Y2=0.38
r68 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.235 $X2=3.255 $Y2=0.38
r69 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.76
+ $Y=0.235 $X2=0.9 $Y2=0.38
.ends

