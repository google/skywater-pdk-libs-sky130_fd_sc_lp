* File: sky130_fd_sc_lp__a2111oi_0.spice
* Created: Fri Aug 28 09:46:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111oi_0.pex.spice"
.subckt sky130_fd_sc_lp__a2111oi_0  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_D1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_C1_M1008_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1000 A_432_47# N_A1_M1000_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g A_432_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.9 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 A_174_483# N_D1_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.1888 PD=0.85 PS=1.87 NRD=15.3857 NRS=9.2196 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1004 A_246_483# N_C1_M1004_g A_174_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.0672 PD=0.85 PS=0.85 NRD=15.3857 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1009 N_A_318_483#_M1009_d N_B1_M1009_g A_246_483# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.9
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_318_483#_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1216 AS=0.0896 PD=1.02 PS=0.92 NRD=13.8491 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1001 N_A_318_483#_M1001_d N_A2_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1216 PD=1.81 PS=1.02 NRD=0 NRS=16.9223 M=1 R=4.26667
+ SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a2111oi_0.pxi.spice"
*
.ends
*
*
