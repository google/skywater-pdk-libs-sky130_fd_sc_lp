* File: sky130_fd_sc_lp__nor4bb_2.spice
* Created: Wed Sep  2 10:11:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4bb_2.pex.spice"
.subckt sky130_fd_sc_lp__nor4bb_2  VNB VPB C_N D_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_C_N_M1006_g N_A_45_164#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1491 AS=0.1113 PD=1.13 PS=1.37 NRD=2.856 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_A_286_512#_M1007_d N_D_N_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1491 PD=1.37 PS=1.13 NRD=0 NRS=120 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_Y_M1012_d N_A_286_512#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.7 A=0.126 P=1.98 MULT=1
MM1015 N_Y_M1012_d N_A_286_512#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_A_45_164#_M1000_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1010 N_Y_M1000_d N_A_45_164#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3192 PD=1.12 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5 SB=75002.4
+ A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.3192 PD=1.12 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4 SB=75001.5 A=0.126
+ P=1.98 MULT=1
MM1008 N_Y_M1002_d N_B_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8 SB=75001.1 A=0.126
+ P=1.98 MULT=1
MM1004 N_VGND_M1008_s N_A_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2 SB=75000.6 A=0.126
+ P=1.98 MULT=1
MM1018 N_VGND_M1018_d N_A_M1018_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.7 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1014 N_VPWR_M1014_d N_C_N_M1014_g N_A_45_164#_M1014_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1302 AS=0.1113 PD=1.04 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1011 N_A_286_512#_M1011_d N_D_N_M1011_g N_VPWR_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1449 AS=0.1302 PD=1.53 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_A_286_512#_M1005_g N_A_463_355#_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1016 N_Y_M1005_d N_A_286_512#_M1016_g N_A_463_355#_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1001 N_A_718_355#_M1001_d N_A_45_164#_M1001_g N_A_463_355#_M1016_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1017 N_A_718_355#_M1001_d N_A_45_164#_M1017_g N_A_463_355#_M1017_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.2016 AS=0.3339 PD=1.58 PS=3.05 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1009 N_A_718_355#_M1009_d N_B_M1009_g N_A_919_367#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1019 N_A_718_355#_M1009_d N_B_M1019_g N_A_919_367#_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 N_A_919_367#_M1019_s N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_A_919_367#_M1013_d N_A_M1013_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=13.3837 P=18.05
*
.include "sky130_fd_sc_lp__nor4bb_2.pxi.spice"
*
.ends
*
*
