* File: sky130_fd_sc_lp__a31oi_1.pxi.spice
* Created: Wed Sep  2 09:26:56 2020
* 
x_PM_SKY130_FD_SC_LP__A31OI_1%A3 N_A3_M1003_g N_A3_M1000_g A3 A3 N_A3_c_47_n
+ PM_SKY130_FD_SC_LP__A31OI_1%A3
x_PM_SKY130_FD_SC_LP__A31OI_1%A2 N_A2_M1006_g N_A2_M1005_g A2 A2 N_A2_c_75_n
+ N_A2_c_76_n PM_SKY130_FD_SC_LP__A31OI_1%A2
x_PM_SKY130_FD_SC_LP__A31OI_1%A1 N_A1_M1007_g N_A1_M1001_g A1 N_A1_c_111_n
+ N_A1_c_112_n PM_SKY130_FD_SC_LP__A31OI_1%A1
x_PM_SKY130_FD_SC_LP__A31OI_1%B1 N_B1_c_144_n N_B1_M1002_g N_B1_M1004_g
+ N_B1_c_146_n B1 N_B1_c_148_n PM_SKY130_FD_SC_LP__A31OI_1%B1
x_PM_SKY130_FD_SC_LP__A31OI_1%VPWR N_VPWR_M1000_s N_VPWR_M1005_d N_VPWR_c_169_n
+ N_VPWR_c_170_n N_VPWR_c_171_n N_VPWR_c_172_n N_VPWR_c_173_n N_VPWR_c_174_n
+ VPWR N_VPWR_c_175_n N_VPWR_c_168_n PM_SKY130_FD_SC_LP__A31OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A31OI_1%A_151_367# N_A_151_367#_M1000_d
+ N_A_151_367#_M1001_d N_A_151_367#_c_202_n N_A_151_367#_c_203_n
+ N_A_151_367#_c_206_n N_A_151_367#_c_210_n N_A_151_367#_c_207_n
+ PM_SKY130_FD_SC_LP__A31OI_1%A_151_367#
x_PM_SKY130_FD_SC_LP__A31OI_1%Y N_Y_M1007_d N_Y_M1004_d N_Y_c_229_n N_Y_c_243_n
+ N_Y_c_237_n N_Y_c_231_n N_Y_c_238_n N_Y_c_249_n Y Y Y N_Y_c_232_n
+ PM_SKY130_FD_SC_LP__A31OI_1%Y
x_PM_SKY130_FD_SC_LP__A31OI_1%VGND N_VGND_M1003_s N_VGND_M1002_d N_VGND_c_286_n
+ N_VGND_c_287_n N_VGND_c_288_n N_VGND_c_289_n N_VGND_c_290_n N_VGND_c_291_n
+ VGND N_VGND_c_292_n N_VGND_c_293_n PM_SKY130_FD_SC_LP__A31OI_1%VGND
cc_1 VNB N_A3_M1003_g 0.0227684f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.655
cc_2 VNB N_A3_M1000_g 0.00576589f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.465
cc_3 VNB A3 0.0292683f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A3_c_47_n 0.0490987f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.375
cc_5 VNB N_A2_M1005_g 0.00827039f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.465
cc_6 VNB A2 0.00460928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A2_c_75_n 0.0314162f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.375
cc_8 VNB N_A2_c_76_n 0.016325f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.375
cc_9 VNB N_A1_M1001_g 0.00830966f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.465
cc_10 VNB A1 0.00330794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_111_n 0.0326602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_c_112_n 0.0185809f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.375
cc_13 VNB N_B1_c_144_n 0.0223944f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.21
cc_14 VNB N_B1_M1004_g 0.0114223f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.465
cc_15 VNB N_B1_c_146_n 0.0085837f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB B1 0.0204929f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_B1_c_148_n 0.0584173f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.375
cc_18 VNB N_VPWR_c_168_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_229_n 0.00388667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_286_n 0.0350191f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_21 VNB N_VGND_c_287_n 0.033023f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.375
cc_22 VNB N_VGND_c_288_n 0.0116899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_289_n 0.00470882f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.375
cc_24 VNB N_VGND_c_290_n 0.0383484f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.295
cc_25 VNB N_VGND_c_291_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_292_n 0.0139174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_293_n 0.187335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A3_M1000_g 0.0238541f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.465
cc_29 VPB A3 0.0174886f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_30 VPB N_A2_M1005_g 0.0204119f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.465
cc_31 VPB N_A1_M1001_g 0.0204395f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.465
cc_32 VPB N_B1_M1004_g 0.0244821f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.465
cc_33 VPB N_VPWR_c_169_n 0.0483272f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_34 VPB N_VPWR_c_170_n 0.00561774f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.375
cc_35 VPB N_VPWR_c_171_n 0.0116899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_172_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=1.295
cc_37 VPB N_VPWR_c_173_n 0.0185493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_174_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=1.375
cc_39 VPB N_VPWR_c_175_n 0.0356957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_168_n 0.0539702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_Y_c_229_n 2.74761e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_Y_c_231_n 0.0280147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_Y_c_232_n 0.0610829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 N_A3_c_47_n N_A2_M1005_g 0.0267895f $X=0.68 $Y=1.375 $X2=0 $Y2=0
cc_45 N_A3_M1003_g A2 6.50599e-19 $X=0.68 $Y=0.655 $X2=0 $Y2=0
cc_46 N_A3_c_47_n N_A2_c_75_n 0.0432999f $X=0.68 $Y=1.375 $X2=0 $Y2=0
cc_47 N_A3_M1003_g N_A2_c_76_n 0.0432999f $X=0.68 $Y=0.655 $X2=0 $Y2=0
cc_48 N_A3_M1000_g N_VPWR_c_169_n 0.00565666f $X=0.68 $Y=2.465 $X2=0 $Y2=0
cc_49 A3 N_VPWR_c_169_n 0.0221097f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_50 N_A3_c_47_n N_VPWR_c_169_n 0.00143386f $X=0.68 $Y=1.375 $X2=0 $Y2=0
cc_51 N_A3_M1000_g N_VPWR_c_173_n 0.00549284f $X=0.68 $Y=2.465 $X2=0 $Y2=0
cc_52 N_A3_M1000_g N_VPWR_c_168_n 0.0108686f $X=0.68 $Y=2.465 $X2=0 $Y2=0
cc_53 N_A3_M1000_g N_A_151_367#_c_202_n 0.00216508f $X=0.68 $Y=2.465 $X2=0 $Y2=0
cc_54 N_A3_M1000_g N_A_151_367#_c_203_n 0.0101703f $X=0.68 $Y=2.465 $X2=0 $Y2=0
cc_55 N_A3_M1003_g N_Y_c_229_n 0.0164968f $X=0.68 $Y=0.655 $X2=0 $Y2=0
cc_56 N_A3_M1000_g N_Y_c_229_n 0.0026683f $X=0.68 $Y=2.465 $X2=0 $Y2=0
cc_57 A3 N_Y_c_229_n 0.0354012f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_58 N_A3_c_47_n N_Y_c_229_n 0.00746582f $X=0.68 $Y=1.375 $X2=0 $Y2=0
cc_59 N_A3_M1003_g N_Y_c_237_n 0.00605394f $X=0.68 $Y=0.655 $X2=0 $Y2=0
cc_60 N_A3_M1000_g N_Y_c_238_n 0.0078215f $X=0.68 $Y=2.465 $X2=0 $Y2=0
cc_61 A3 N_Y_c_238_n 0.00817525f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A3_M1003_g N_VGND_c_286_n 0.00910611f $X=0.68 $Y=0.655 $X2=0 $Y2=0
cc_63 A3 N_VGND_c_286_n 0.0210263f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A3_c_47_n N_VGND_c_286_n 0.00192328f $X=0.68 $Y=1.375 $X2=0 $Y2=0
cc_65 N_A3_M1003_g N_VGND_c_290_n 0.0052466f $X=0.68 $Y=0.655 $X2=0 $Y2=0
cc_66 N_A3_M1003_g N_VGND_c_293_n 0.0101938f $X=0.68 $Y=0.655 $X2=0 $Y2=0
cc_67 N_A2_M1005_g N_A1_M1001_g 0.0404761f $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_68 A2 A1 0.02585f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_69 N_A2_c_75_n A1 3.80526e-19 $X=1.14 $Y=1.35 $X2=0 $Y2=0
cc_70 N_A2_c_75_n N_A1_c_111_n 0.0206327f $X=1.14 $Y=1.35 $X2=0 $Y2=0
cc_71 A2 N_A1_c_112_n 0.00821384f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_72 N_A2_c_76_n N_A1_c_112_n 0.0293133f $X=1.135 $Y=1.185 $X2=0 $Y2=0
cc_73 N_A2_M1005_g N_VPWR_c_170_n 0.00763749f $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_74 N_A2_M1005_g N_VPWR_c_173_n 0.00549284f $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_75 N_A2_M1005_g N_VPWR_c_168_n 0.0103164f $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_76 N_A2_M1005_g N_A_151_367#_c_202_n 7.32094e-19 $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A2_M1005_g N_A_151_367#_c_203_n 0.0118094f $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A2_M1005_g N_A_151_367#_c_206_n 0.0118785f $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A2_M1005_g N_A_151_367#_c_207_n 9.05717e-19 $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A2_M1005_g N_Y_c_229_n 0.00358154f $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_81 A2 N_Y_c_229_n 0.0564627f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_82 N_A2_c_76_n N_Y_c_229_n 0.00945139f $X=1.135 $Y=1.185 $X2=0 $Y2=0
cc_83 A2 N_Y_c_243_n 0.0146619f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A2_c_75_n N_Y_c_243_n 5.07257e-19 $X=1.14 $Y=1.35 $X2=0 $Y2=0
cc_85 N_A2_c_76_n N_Y_c_243_n 0.0169681f $X=1.135 $Y=1.185 $X2=0 $Y2=0
cc_86 N_A2_M1005_g N_Y_c_231_n 0.0118095f $X=1.11 $Y=2.465 $X2=0 $Y2=0
cc_87 A2 N_Y_c_231_n 0.0227105f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A2_c_75_n N_Y_c_231_n 0.00375137f $X=1.14 $Y=1.35 $X2=0 $Y2=0
cc_89 A2 N_Y_c_249_n 0.0136523f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_90 N_A2_c_76_n N_Y_c_249_n 0.00123497f $X=1.135 $Y=1.185 $X2=0 $Y2=0
cc_91 N_A2_c_76_n N_VGND_c_290_n 0.00357877f $X=1.135 $Y=1.185 $X2=0 $Y2=0
cc_92 N_A2_c_76_n N_VGND_c_293_n 0.00556329f $X=1.135 $Y=1.185 $X2=0 $Y2=0
cc_93 A2 A_223_47# 0.00631717f $X=1.115 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_94 N_A1_c_112_n N_B1_c_144_n 0.0198942f $X=1.68 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_95 N_A1_M1001_g N_B1_M1004_g 0.0282691f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_96 A1 N_B1_c_146_n 3.73807e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A1_c_111_n N_B1_c_146_n 0.0207362f $X=1.68 $Y=1.35 $X2=0 $Y2=0
cc_98 A1 B1 0.0276613f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A1_c_111_n B1 0.00201148f $X=1.68 $Y=1.35 $X2=0 $Y2=0
cc_100 N_A1_M1001_g N_VPWR_c_170_n 0.00763749f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A1_M1001_g N_VPWR_c_175_n 0.00549284f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A1_M1001_g N_VPWR_c_168_n 0.0103164f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A1_M1001_g N_A_151_367#_c_203_n 9.05717e-19 $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A1_M1001_g N_A_151_367#_c_206_n 0.0118785f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A1_M1001_g N_A_151_367#_c_210_n 7.32094e-19 $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A1_M1001_g N_A_151_367#_c_207_n 0.0118094f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_107 A1 N_Y_c_243_n 0.00285319f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_108 N_A1_c_112_n N_Y_c_243_n 0.0117041f $X=1.68 $Y=1.185 $X2=0 $Y2=0
cc_109 N_A1_M1001_g N_Y_c_231_n 0.0111672f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_110 A1 N_Y_c_231_n 0.0242118f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_111 N_A1_c_111_n N_Y_c_231_n 0.00124454f $X=1.68 $Y=1.35 $X2=0 $Y2=0
cc_112 A1 N_Y_c_249_n 0.0145712f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_113 N_A1_c_111_n N_Y_c_249_n 0.00123361f $X=1.68 $Y=1.35 $X2=0 $Y2=0
cc_114 N_A1_c_112_n N_Y_c_249_n 0.011119f $X=1.68 $Y=1.185 $X2=0 $Y2=0
cc_115 N_A1_c_112_n N_VGND_c_287_n 0.0011553f $X=1.68 $Y=1.185 $X2=0 $Y2=0
cc_116 N_A1_c_112_n N_VGND_c_290_n 0.00357835f $X=1.68 $Y=1.185 $X2=0 $Y2=0
cc_117 N_A1_c_112_n N_VGND_c_293_n 0.00592798f $X=1.68 $Y=1.185 $X2=0 $Y2=0
cc_118 N_B1_M1004_g N_VPWR_c_175_n 0.00549284f $X=2.13 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B1_M1004_g N_VPWR_c_168_n 0.0110478f $X=2.13 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B1_M1004_g N_A_151_367#_c_210_n 0.00216614f $X=2.13 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_B1_M1004_g N_A_151_367#_c_207_n 0.0101703f $X=2.13 $Y=2.465 $X2=0 $Y2=0
cc_122 N_B1_M1004_g N_Y_c_231_n 0.0156445f $X=2.13 $Y=2.465 $X2=0 $Y2=0
cc_123 B1 N_Y_c_231_n 0.0634408f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_124 N_B1_c_148_n N_Y_c_231_n 0.0120519f $X=2.56 $Y=1.35 $X2=0 $Y2=0
cc_125 N_B1_c_144_n N_VGND_c_287_n 0.0176364f $X=2.13 $Y=1.185 $X2=0 $Y2=0
cc_126 B1 N_VGND_c_287_n 0.0244507f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B1_c_148_n N_VGND_c_287_n 0.00688795f $X=2.56 $Y=1.35 $X2=0 $Y2=0
cc_128 N_B1_c_144_n N_VGND_c_290_n 0.00486043f $X=2.13 $Y=1.185 $X2=0 $Y2=0
cc_129 N_B1_c_144_n N_VGND_c_293_n 0.00864313f $X=2.13 $Y=1.185 $X2=0 $Y2=0
cc_130 N_VPWR_c_168_n N_A_151_367#_M1000_d 0.00223819f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_131 N_VPWR_c_168_n N_A_151_367#_M1001_d 0.00223819f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_132 N_VPWR_c_173_n N_A_151_367#_c_203_n 0.0177952f $X=1.24 $Y=3.33 $X2=0
+ $Y2=0
cc_133 N_VPWR_c_168_n N_A_151_367#_c_203_n 0.0123247f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_134 N_VPWR_M1005_d N_A_151_367#_c_206_n 0.0075503f $X=1.185 $Y=1.835 $X2=0
+ $Y2=0
cc_135 N_VPWR_c_170_n N_A_151_367#_c_206_n 0.0265229f $X=1.405 $Y=2.45 $X2=0
+ $Y2=0
cc_136 N_VPWR_c_175_n N_A_151_367#_c_207_n 0.0177952f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_137 N_VPWR_c_168_n N_A_151_367#_c_207_n 0.0123247f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_138 N_VPWR_c_168_n N_Y_M1004_d 0.00438725f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_139 N_VPWR_M1005_d N_Y_c_231_n 0.00355802f $X=1.185 $Y=1.835 $X2=0 $Y2=0
cc_140 N_VPWR_c_175_n N_Y_c_232_n 0.0381319f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_141 N_VPWR_c_168_n N_Y_c_232_n 0.0211106f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_142 N_A_151_367#_M1000_d N_Y_c_231_n 9.77978e-19 $X=0.755 $Y=1.835 $X2=0
+ $Y2=0
cc_143 N_A_151_367#_M1001_d N_Y_c_231_n 0.00176461f $X=1.775 $Y=1.835 $X2=0
+ $Y2=0
cc_144 N_A_151_367#_c_202_n N_Y_c_231_n 0.00939213f $X=0.895 $Y=2.195 $X2=0
+ $Y2=0
cc_145 N_A_151_367#_c_206_n N_Y_c_231_n 0.0405558f $X=1.75 $Y=2.11 $X2=0 $Y2=0
cc_146 N_A_151_367#_c_210_n N_Y_c_231_n 0.01723f $X=1.915 $Y=2.195 $X2=0 $Y2=0
cc_147 N_A_151_367#_M1000_d N_Y_c_238_n 8.07836e-19 $X=0.755 $Y=1.835 $X2=0
+ $Y2=0
cc_148 N_A_151_367#_c_202_n N_Y_c_238_n 0.00865576f $X=0.895 $Y=2.195 $X2=0
+ $Y2=0
cc_149 N_Y_c_229_n N_VGND_c_286_n 0.0368122f $X=0.8 $Y=1.685 $X2=0 $Y2=0
cc_150 N_Y_c_237_n N_VGND_c_286_n 0.0221788f $X=0.885 $Y=0.392 $X2=0 $Y2=0
cc_151 N_Y_c_243_n N_VGND_c_290_n 0.0433579f $X=1.635 $Y=0.392 $X2=0 $Y2=0
cc_152 N_Y_c_237_n N_VGND_c_290_n 0.00988214f $X=0.885 $Y=0.392 $X2=0 $Y2=0
cc_153 N_Y_c_249_n N_VGND_c_290_n 0.0238669f $X=1.845 $Y=0.42 $X2=0 $Y2=0
cc_154 N_Y_M1007_d N_VGND_c_293_n 0.00470374f $X=1.665 $Y=0.235 $X2=0 $Y2=0
cc_155 N_Y_c_243_n N_VGND_c_293_n 0.0272577f $X=1.635 $Y=0.392 $X2=0 $Y2=0
cc_156 N_Y_c_237_n N_VGND_c_293_n 0.00642618f $X=0.885 $Y=0.392 $X2=0 $Y2=0
cc_157 N_Y_c_249_n N_VGND_c_293_n 0.0143687f $X=1.845 $Y=0.42 $X2=0 $Y2=0
cc_158 N_Y_c_229_n A_151_47# 0.00507911f $X=0.8 $Y=1.685 $X2=-0.19 $Y2=-0.245
cc_159 N_Y_c_243_n A_151_47# 0.00109935f $X=1.635 $Y=0.392 $X2=-0.19 $Y2=-0.245
cc_160 N_Y_c_237_n A_151_47# 7.13792e-19 $X=0.885 $Y=0.392 $X2=-0.19 $Y2=-0.245
cc_161 N_Y_c_243_n A_223_47# 0.00989114f $X=1.635 $Y=0.392 $X2=-0.19 $Y2=-0.245
cc_162 N_VGND_c_293_n A_151_47# 0.00168881f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_163 N_VGND_c_293_n A_223_47# 0.00323039f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
