* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VGND a_102_53# X VNB nshort w=840000u l=150000u
+  ad=1.0962e+12p pd=9.33e+06u as=2.352e+11p ps=2.24e+06u
M1001 a_753_367# A2 a_645_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.914e+11p pd=3.3e+06u as=4.914e+11p ps=3.3e+06u
M1002 a_465_49# A1 VGND VNB nshort w=840000u l=150000u
+  ad=7.308e+11p pd=6.78e+06u as=0p ps=0u
M1003 VPWR a_102_53# X VPB phighvt w=1.26e+06u l=150000u
+  ad=1.7514e+12p pd=1.034e+07u as=3.528e+11p ps=3.08e+06u
M1004 a_465_49# B1 a_102_53# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1005 VPWR A1 a_753_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_465_49# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_102_53# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.812e+11p pd=3.76e+06u as=0p ps=0u
M1008 a_573_367# A4 a_102_53# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1009 a_645_367# A3 a_573_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A4 a_465_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_102_53# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_465_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_102_53# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
