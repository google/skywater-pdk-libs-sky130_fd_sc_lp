* File: sky130_fd_sc_lp__nor3b_1.pxi.spice
* Created: Wed Sep  2 10:09:34 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3B_1%C_N N_C_N_c_52_n N_C_N_M1000_g N_C_N_c_53_n
+ N_C_N_M1004_g C_N C_N PM_SKY130_FD_SC_LP__NOR3B_1%C_N
x_PM_SKY130_FD_SC_LP__NOR3B_1%A N_A_M1002_g N_A_M1006_g A A N_A_c_80_n
+ PM_SKY130_FD_SC_LP__NOR3B_1%A
x_PM_SKY130_FD_SC_LP__NOR3B_1%B N_B_M1007_g N_B_M1003_g B N_B_c_113_n
+ N_B_c_114_n PM_SKY130_FD_SC_LP__NOR3B_1%B
x_PM_SKY130_FD_SC_LP__NOR3B_1%A_82_131# N_A_82_131#_M1000_s N_A_82_131#_M1004_s
+ N_A_82_131#_M1005_g N_A_82_131#_M1001_g N_A_82_131#_c_150_n
+ N_A_82_131#_c_156_n N_A_82_131#_c_157_n N_A_82_131#_c_158_n
+ N_A_82_131#_c_151_n N_A_82_131#_c_152_n N_A_82_131#_c_153_n
+ PM_SKY130_FD_SC_LP__NOR3B_1%A_82_131#
x_PM_SKY130_FD_SC_LP__NOR3B_1%VPWR N_VPWR_M1004_d N_VPWR_c_211_n VPWR
+ N_VPWR_c_212_n N_VPWR_c_213_n N_VPWR_c_210_n N_VPWR_c_215_n
+ PM_SKY130_FD_SC_LP__NOR3B_1%VPWR
x_PM_SKY130_FD_SC_LP__NOR3B_1%Y N_Y_M1002_d N_Y_M1005_d N_Y_M1001_d N_Y_c_245_n
+ N_Y_c_237_n N_Y_c_238_n Y Y Y Y Y Y Y N_Y_c_241_n Y N_Y_c_244_n Y
+ PM_SKY130_FD_SC_LP__NOR3B_1%Y
x_PM_SKY130_FD_SC_LP__NOR3B_1%VGND N_VGND_M1000_d N_VGND_M1003_d N_VGND_c_280_n
+ N_VGND_c_281_n N_VGND_c_282_n N_VGND_c_283_n N_VGND_c_284_n N_VGND_c_285_n
+ VGND N_VGND_c_286_n N_VGND_c_287_n PM_SKY130_FD_SC_LP__NOR3B_1%VGND
cc_1 VNB N_C_N_c_52_n 0.0220963f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.185
cc_2 VNB N_C_N_c_53_n 0.0453423f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.725
cc_3 VNB C_N 0.00419604f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_M1002_g 0.0204782f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.865
cc_5 VNB N_A_M1006_g 0.00569683f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB A 0.00489625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_c_80_n 0.0324012f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.295
cc_8 VNB N_B_M1003_g 0.0244978f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_9 VNB N_B_c_113_n 0.0239515f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.375
cc_10 VNB N_B_c_114_n 0.00335852f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.375
cc_11 VNB N_A_82_131#_M1005_g 0.0298329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_82_131#_c_150_n 0.0324482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_82_131#_c_151_n 0.0261008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_82_131#_c_152_n 0.00294532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_82_131#_c_153_n 0.0258962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_210_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.665
cc_17 VNB N_Y_c_237_n 0.0054084f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.295
cc_18 VNB N_Y_c_238_n 0.00515006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB Y 0.0113625f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.375
cc_20 VNB Y 0.0248189f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.665
cc_21 VNB N_Y_c_241_n 0.0378672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_280_n 0.0150429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_281_n 4.05231e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_282_n 0.0254736f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.665
cc_25 VNB N_VGND_c_283_n 0.00744248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_284_n 0.0140536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_285_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_286_n 0.0199888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_287_n 0.179791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_C_N_c_53_n 0.0318927f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.725
cc_31 VPB C_N 0.00386745f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_32 VPB N_A_M1006_g 0.021489f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_33 VPB A 0.00249576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_B_M1007_g 0.0187219f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.865
cc_35 VPB N_B_c_113_n 0.00612452f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.375
cc_36 VPB N_B_c_114_n 0.00255697f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.375
cc_37 VPB N_A_82_131#_M1001_g 0.0242036f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.375
cc_38 VPB N_A_82_131#_c_150_n 0.0145882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_82_131#_c_156_n 0.00813385f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.375
cc_40 VPB N_A_82_131#_c_157_n 0.0191401f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.665
cc_41 VPB N_A_82_131#_c_158_n 0.00170512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_82_131#_c_152_n 4.22419e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_82_131#_c_153_n 0.00727464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_211_n 0.0312973f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.045
cc_45 VPB N_VPWR_c_212_n 0.0314195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_213_n 0.0487517f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.375
cc_47 VPB N_VPWR_c_210_n 0.0796963f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.665
cc_48 VPB N_VPWR_c_215_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB Y 0.00949366f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.665
cc_50 VPB Y 0.0497105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_Y_c_244_n 0.0106954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 N_C_N_c_52_n N_A_M1002_g 0.0135375f $X=0.75 $Y=1.185 $X2=0 $Y2=0
cc_53 N_C_N_c_53_n N_A_M1006_g 0.0234138f $X=0.75 $Y=1.725 $X2=0 $Y2=0
cc_54 C_N N_A_M1006_g 5.5391e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_55 N_C_N_c_52_n A 6.99187e-19 $X=0.75 $Y=1.185 $X2=0 $Y2=0
cc_56 N_C_N_c_53_n A 0.00172616f $X=0.75 $Y=1.725 $X2=0 $Y2=0
cc_57 C_N A 0.0463327f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_58 N_C_N_c_53_n N_A_c_80_n 0.0193932f $X=0.75 $Y=1.725 $X2=0 $Y2=0
cc_59 C_N N_A_c_80_n 0.00111883f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_60 N_C_N_c_52_n N_A_82_131#_c_150_n 0.004001f $X=0.75 $Y=1.185 $X2=0 $Y2=0
cc_61 N_C_N_c_53_n N_A_82_131#_c_150_n 0.013228f $X=0.75 $Y=1.725 $X2=0 $Y2=0
cc_62 C_N N_A_82_131#_c_150_n 0.0435819f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_63 N_C_N_c_53_n N_A_82_131#_c_156_n 0.0152038f $X=0.75 $Y=1.725 $X2=0 $Y2=0
cc_64 C_N N_A_82_131#_c_156_n 0.0272342f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_C_N_c_53_n N_A_82_131#_c_151_n 0.00406694f $X=0.75 $Y=1.725 $X2=0 $Y2=0
cc_66 C_N N_A_82_131#_c_151_n 0.0114783f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_C_N_c_53_n N_VPWR_c_211_n 0.00203938f $X=0.75 $Y=1.725 $X2=0 $Y2=0
cc_68 N_C_N_c_52_n N_VGND_c_280_n 0.0144733f $X=0.75 $Y=1.185 $X2=0 $Y2=0
cc_69 C_N N_VGND_c_280_n 0.00309041f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_C_N_c_52_n N_VGND_c_282_n 0.00332367f $X=0.75 $Y=1.185 $X2=0 $Y2=0
cc_71 N_C_N_c_52_n N_VGND_c_287_n 0.00387424f $X=0.75 $Y=1.185 $X2=0 $Y2=0
cc_72 N_A_M1006_g N_B_M1007_g 0.0589271f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A_M1002_g N_B_M1003_g 0.0199485f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_74 A N_B_M1003_g 8.39466e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_75 A N_B_c_113_n 4.47495e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_76 N_A_c_80_n N_B_c_113_n 0.0589271f $X=1.2 $Y=1.375 $X2=0 $Y2=0
cc_77 A N_B_c_114_n 0.0323644f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_c_80_n N_B_c_114_n 0.00224464f $X=1.2 $Y=1.375 $X2=0 $Y2=0
cc_79 N_A_M1006_g N_A_82_131#_c_156_n 0.0165645f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_80 A N_A_82_131#_c_156_n 0.0242298f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_c_80_n N_A_82_131#_c_156_n 7.32358e-19 $X=1.2 $Y=1.375 $X2=0 $Y2=0
cc_82 N_A_M1006_g N_VPWR_c_211_n 0.0227301f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_VPWR_c_213_n 0.00486043f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_84 N_A_M1006_g N_VPWR_c_210_n 0.00818711f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_M1002_g N_Y_c_245_n 0.00291841f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_86 N_A_M1002_g N_Y_c_238_n 0.00473475f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_VGND_c_280_n 0.0206559f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_88 A N_VGND_c_280_n 0.0171479f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_c_80_n N_VGND_c_280_n 0.00122182f $X=1.2 $Y=1.375 $X2=0 $Y2=0
cc_90 N_A_M1002_g N_VGND_c_281_n 5.9376e-19 $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_VGND_c_284_n 0.00486043f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_92 N_A_M1002_g N_VGND_c_287_n 0.00835496f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_93 N_B_M1003_g N_A_82_131#_M1005_g 0.0243592f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_94 N_B_M1007_g N_A_82_131#_M1001_g 0.0491277f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_95 N_B_c_114_n N_A_82_131#_M1001_g 2.31147e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_96 N_B_M1007_g N_A_82_131#_c_156_n 0.0168252f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_97 N_B_c_113_n N_A_82_131#_c_156_n 0.0033148f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_98 N_B_c_114_n N_A_82_131#_c_156_n 0.0188971f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_99 N_B_M1007_g N_A_82_131#_c_158_n 0.0035253f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_100 N_B_c_114_n N_A_82_131#_c_158_n 0.00667571f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_101 N_B_c_113_n N_A_82_131#_c_152_n 0.00217947f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_102 N_B_c_114_n N_A_82_131#_c_152_n 0.0259089f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_103 N_B_c_113_n N_A_82_131#_c_153_n 0.0204013f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_104 N_B_c_114_n N_A_82_131#_c_153_n 2.82575e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B_M1007_g N_VPWR_c_211_n 0.00506879f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_106 N_B_M1007_g N_VPWR_c_213_n 0.00585385f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_107 N_B_M1007_g N_VPWR_c_210_n 0.011101f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_108 N_B_M1003_g N_Y_c_237_n 0.0133931f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_109 N_B_c_113_n N_Y_c_237_n 0.00311113f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_110 N_B_c_114_n N_Y_c_237_n 0.0136199f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_111 N_B_c_113_n N_Y_c_238_n 4.67499e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_112 N_B_c_114_n N_Y_c_238_n 0.00982317f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_113 N_B_M1003_g N_VGND_c_280_n 6.79764e-19 $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_114 N_B_M1003_g N_VGND_c_281_n 0.0102296f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_115 N_B_M1003_g N_VGND_c_284_n 0.00486043f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_116 N_B_M1003_g N_VGND_c_287_n 0.00835496f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_117 N_A_82_131#_c_156_n N_VPWR_M1004_d 0.0116941f $X=2.005 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_82_131#_c_156_n N_VPWR_c_211_n 0.0222677f $X=2.005 $Y=2.035 $X2=0
+ $Y2=0
cc_119 N_A_82_131#_M1001_g N_VPWR_c_213_n 0.00585385f $X=2.2 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_82_131#_M1001_g N_VPWR_c_210_n 0.0122384f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_82_131#_c_156_n A_275_367# 0.00751567f $X=2.005 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_82_131#_c_156_n A_347_367# 0.0162f $X=2.005 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_82_131#_c_158_n A_347_367# 0.00117769f $X=2.09 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_82_131#_M1005_g N_Y_c_237_n 0.0145281f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_125 N_A_82_131#_c_152_n N_Y_c_237_n 0.0231948f $X=2.29 $Y=1.505 $X2=0 $Y2=0
cc_126 N_A_82_131#_c_153_n N_Y_c_237_n 8.94628e-19 $X=2.29 $Y=1.505 $X2=0 $Y2=0
cc_127 N_A_82_131#_c_152_n Y 0.00590333f $X=2.29 $Y=1.505 $X2=0 $Y2=0
cc_128 N_A_82_131#_c_153_n Y 0.00374225f $X=2.29 $Y=1.505 $X2=0 $Y2=0
cc_129 N_A_82_131#_M1005_g Y 0.00379002f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_130 N_A_82_131#_M1001_g Y 0.00226322f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A_82_131#_c_158_n Y 0.00483787f $X=2.09 $Y=1.93 $X2=0 $Y2=0
cc_132 N_A_82_131#_c_152_n Y 0.0257056f $X=2.29 $Y=1.505 $X2=0 $Y2=0
cc_133 N_A_82_131#_c_153_n Y 0.00813609f $X=2.29 $Y=1.505 $X2=0 $Y2=0
cc_134 N_A_82_131#_M1001_g N_Y_c_244_n 0.0259698f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_82_131#_c_156_n N_Y_c_244_n 0.0176628f $X=2.005 $Y=2.035 $X2=0 $Y2=0
cc_136 N_A_82_131#_c_158_n N_Y_c_244_n 0.00679624f $X=2.09 $Y=1.93 $X2=0 $Y2=0
cc_137 N_A_82_131#_c_152_n N_Y_c_244_n 0.00322064f $X=2.29 $Y=1.505 $X2=0 $Y2=0
cc_138 N_A_82_131#_c_153_n N_Y_c_244_n 0.00302008f $X=2.29 $Y=1.505 $X2=0 $Y2=0
cc_139 N_A_82_131#_M1005_g N_VGND_c_281_n 0.0114527f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_140 N_A_82_131#_c_151_n N_VGND_c_282_n 0.00886477f $X=0.535 $Y=0.865 $X2=0
+ $Y2=0
cc_141 N_A_82_131#_M1005_g N_VGND_c_286_n 0.00505556f $X=2.2 $Y=0.655 $X2=0
+ $Y2=0
cc_142 N_A_82_131#_M1005_g N_VGND_c_287_n 0.00963349f $X=2.2 $Y=0.655 $X2=0
+ $Y2=0
cc_143 N_A_82_131#_c_151_n N_VGND_c_287_n 0.0152263f $X=0.535 $Y=0.865 $X2=0
+ $Y2=0
cc_144 N_VPWR_c_210_n A_275_367# 0.00899413f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_145 N_VPWR_c_210_n A_347_367# 0.0167135f $X=2.64 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_146 N_VPWR_c_210_n N_Y_M1001_d 0.00471238f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_147 N_VPWR_c_213_n Y 0.0317922f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_148 N_VPWR_c_210_n Y 0.0174119f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_149 N_Y_c_237_n N_VGND_M1003_d 0.00181776f $X=2.315 $Y=1.085 $X2=0 $Y2=0
cc_150 N_Y_c_245_n N_VGND_c_280_n 0.0491485f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_151 N_Y_c_238_n N_VGND_c_280_n 7.30395e-19 $X=1.645 $Y=1.085 $X2=0 $Y2=0
cc_152 N_Y_c_237_n N_VGND_c_281_n 0.0171036f $X=2.315 $Y=1.085 $X2=0 $Y2=0
cc_153 N_Y_c_245_n N_VGND_c_284_n 0.0128356f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_154 N_Y_c_241_n N_VGND_c_286_n 0.0334011f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_155 N_Y_M1002_d N_VGND_c_287_n 0.00686549f $X=1.375 $Y=0.235 $X2=0 $Y2=0
cc_156 N_Y_M1005_d N_VGND_c_287_n 0.00354308f $X=2.275 $Y=0.235 $X2=0 $Y2=0
cc_157 N_Y_c_245_n N_VGND_c_287_n 0.00730901f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_158 N_Y_c_241_n N_VGND_c_287_n 0.0185835f $X=2.415 $Y=0.42 $X2=0 $Y2=0
