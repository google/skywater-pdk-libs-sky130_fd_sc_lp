* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 X a_100_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR a_100_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR A4 a_495_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_667_47# A2 a_922_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VPWR A1 a_495_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_495_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VPWR a_100_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_667_47# A1 a_100_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 X a_100_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VGND a_100_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_922_47# A2 a_667_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_1115_47# A3 a_922_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VPWR A3 a_495_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_922_47# A3 a_1115_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_495_367# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR A2 a_495_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_1115_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_100_23# A1 a_667_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_495_367# B1 a_100_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VGND a_100_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 X a_100_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 X a_100_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 VGND B1 a_100_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_100_23# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_495_367# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VGND A4 a_1115_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_100_23# B1 a_495_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 a_495_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
