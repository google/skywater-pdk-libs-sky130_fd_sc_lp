* File: sky130_fd_sc_lp__a2bb2oi_0.spice
* Created: Fri Aug 28 09:56:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2oi_0.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2oi_0  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1003 N_A_110_47#_M1003_d N_A1_N_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A2_N_M1006_g N_A_110_47#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.17745 AS=0.0588 PD=1.265 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_A_110_47#_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.17745 PD=0.7 PS=1.265 NRD=0 NRS=64.284 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 A_481_47# N_B2_M1000_g N_Y_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0798
+ AS=0.0588 PD=0.8 PS=0.7 NRD=38.568 NRS=0 M=1 R=2.8 SA=75002 SB=75000.7 A=0.063
+ P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g A_481_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0798 PD=1.37 PS=0.8 NRD=0 NRS=38.568 M=1 R=2.8 SA=75002.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1007 A_110_427# N_A1_N_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1005 N_A_110_47#_M1005_d N_A2_N_M1005_g A_110_427# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_A_420_387#_M1009_d N_A_110_47#_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1004_d N_B2_M1004_g N_A_420_387#_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_420_387#_M1001_d N_B1_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a2bb2oi_0.pxi.spice"
*
.ends
*
*
