* File: sky130_fd_sc_lp__einvp_1.spice
* Created: Wed Sep  2 09:52:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvp_1.pex.spice"
.subckt sky130_fd_sc_lp__einvp_1  VNB VPB A TE Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* TE	TE
* A	A
* VPB	VPB
* VNB	VNB
MM1003 A_128_47# N_A_M1003_g N_Z_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.2226 PD=1.08 PS=2.21 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2 SB=75001
+ A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_TE_M1001_g A_128_47# VNB NSHORT L=0.15 W=0.84 AD=0.2898
+ AS=0.1008 PD=2.14667 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75000.6 SB=75000.7
+ A=0.126 P=1.98 MULT=1
MM1004 N_A_207_302#_M1004_d N_TE_M1004_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1449 PD=1.41 PS=1.07333 NRD=5.712 NRS=82.848 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_161_400# N_A_M1005_g N_Z_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.115
+ AS=0.285 PD=1.23 PS=2.57 NRD=11.8003 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75000.8
+ A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_207_302#_M1002_g A_161_400# VPB PHIGHVT L=0.15 W=1
+ AD=0.223592 AS=0.115 PD=1.95775 PS=1.23 NRD=2.6201 NRS=11.8003 M=1 R=6.66667
+ SA=75000.6 SB=75000.4 A=0.15 P=2.3 MULT=1
MM1000 N_A_207_302#_M1000_d N_TE_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0939085 PD=1.37 PS=0.822254 NRD=0 NRS=43.3794 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__einvp_1.pxi.spice"
*
.ends
*
*
