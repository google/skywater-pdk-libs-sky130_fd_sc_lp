* File: sky130_fd_sc_lp__decap_3.pex.spice
* Created: Wed Sep  2 09:41:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAP_3%VGND 1 7 9 10 13 14 16 19 23 26 36
r27 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r28 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 27 32 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.25
+ $Y2=0
r30 27 29 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.72
+ $Y2=0
r31 26 35 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.195
+ $Y2=0
r32 26 29 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.72
+ $Y2=0
r33 23 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r34 23 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r35 23 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 19 21 5.30815 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.415 $Y=1.77
+ $X2=0.415 $Y2=1.605
r37 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.77 $X2=0.575 $Y2=1.77
r38 14 35 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.195 $Y2=0
r39 14 16 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.46
r40 13 21 39.2878 $w=3.28e-07 $l=1.125e-06 $layer=LI1_cond $X=0.335 $Y=0.48
+ $X2=0.335 $Y2=1.605
r41 10 32 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.25 $Y2=0
r42 10 13 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.48
r43 7 20 36.8902 $w=5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.66 $Y=2.135 $X2=0.66
+ $Y2=1.77
r44 7 9 44.344 $w=5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.66 $Y=2.135 $X2=0.66
+ $Y2=2.595
r45 1 16 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.235 $X2=1.115 $Y2=0.46
r46 1 13 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.235 $X2=0.335 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__DECAP_3%VPWR 1 7 9 10 12 17 19 26 28 31 41
r27 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r28 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 32 37 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r30 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 31 40 4.53846 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.162 $Y2=3.33
r32 31 34 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r34 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 28 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 23 26 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.755 $Y=1.042
+ $X2=1.05 $Y2=1.042
r37 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.06 $X2=0.755 $Y2=1.06
r38 19 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.05 $Y=2.29
+ $X2=1.05 $Y2=2.97
r39 17 40 3.22771 $w=3.3e-07 $l=1.4854e-07 $layer=LI1_cond $X=1.05 $Y=3.245
+ $X2=1.162 $Y2=3.33
r40 17 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.05 $Y=3.245
+ $X2=1.05 $Y2=2.97
r41 16 26 1.32393 $w=3.3e-07 $l=1.83e-07 $layer=LI1_cond $X=1.05 $Y=1.225
+ $X2=1.05 $Y2=1.042
r42 16 19 37.1925 $w=3.28e-07 $l=1.065e-06 $layer=LI1_cond $X=1.05 $Y=1.225
+ $X2=1.05 $Y2=2.29
r43 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.27
+ $X2=0.26 $Y2=2.95
r44 10 37 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r45 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r46 7 24 39.9593 $w=5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.725 $Y=0.665
+ $X2=0.725 $Y2=1.06
r47 7 9 14.942 $w=5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.725 $Y=0.665 $X2=0.725
+ $Y2=0.51
r48 1 21 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.095 $X2=1.05 $Y2=2.97
r49 1 19 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.095 $X2=1.05 $Y2=2.29
r50 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.095 $X2=0.26 $Y2=2.95
r51 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.095 $X2=0.26 $Y2=2.27
.ends

