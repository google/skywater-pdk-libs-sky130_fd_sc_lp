* File: sky130_fd_sc_lp__a32oi_4.pex.spice
* Created: Wed Sep  2 09:28:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32OI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 49
r83 49 50 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=1.77 $Y=1.35 $X2=1.84
+ $Y2=1.35
r84 47 49 13.472 $w=3.22e-07 $l=9e-08 $layer=POLY_cond $X=1.68 $Y=1.35 $X2=1.77
+ $Y2=1.35
r85 45 47 40.4161 $w=3.22e-07 $l=2.7e-07 $layer=POLY_cond $X=1.41 $Y=1.35
+ $X2=1.68 $Y2=1.35
r86 44 45 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=1.34 $Y=1.35 $X2=1.41
+ $Y2=1.35
r87 43 44 53.8882 $w=3.22e-07 $l=3.6e-07 $layer=POLY_cond $X=0.98 $Y=1.35
+ $X2=1.34 $Y2=1.35
r88 42 43 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=0.91 $Y=1.35 $X2=0.98
+ $Y2=1.35
r89 41 42 53.8882 $w=3.22e-07 $l=3.6e-07 $layer=POLY_cond $X=0.55 $Y=1.35
+ $X2=0.91 $Y2=1.35
r90 40 41 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=0.48 $Y=1.35 $X2=0.55
+ $Y2=1.35
r91 38 40 23.9503 $w=3.22e-07 $l=1.6e-07 $layer=POLY_cond $X=0.32 $Y=1.35
+ $X2=0.48 $Y2=1.35
r92 32 47 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=1.35 $X2=1.68 $Y2=1.35
r93 31 32 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.322
+ $X2=1.68 $Y2=1.322
r94 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.322
+ $X2=1.2 $Y2=1.322
r95 29 30 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.322
+ $X2=0.72 $Y2=1.322
r96 29 38 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.32
+ $Y=1.35 $X2=0.32 $Y2=1.35
r97 25 50 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=1.515
+ $X2=1.84 $Y2=1.35
r98 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.84 $Y=1.515
+ $X2=1.84 $Y2=2.465
r99 22 49 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.185
+ $X2=1.77 $Y2=1.35
r100 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.77 $Y=1.185
+ $X2=1.77 $Y2=0.655
r101 18 45 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.515
+ $X2=1.41 $Y2=1.35
r102 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.41 $Y=1.515
+ $X2=1.41 $Y2=2.465
r103 15 44 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.185
+ $X2=1.34 $Y2=1.35
r104 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.34 $Y=1.185
+ $X2=1.34 $Y2=0.655
r105 11 43 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.515
+ $X2=0.98 $Y2=1.35
r106 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.98 $Y=1.515
+ $X2=0.98 $Y2=2.465
r107 8 42 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.185
+ $X2=0.91 $Y2=1.35
r108 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.91 $Y=1.185
+ $X2=0.91 $Y2=0.655
r109 4 41 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.515
+ $X2=0.55 $Y2=1.35
r110 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.55 $Y=1.515
+ $X2=0.55 $Y2=2.465
r111 1 40 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.185
+ $X2=0.48 $Y2=1.35
r112 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.48 $Y=1.185
+ $X2=0.48 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 50
r83 48 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.56 $Y=1.35 $X2=3.65
+ $Y2=1.35
r84 47 48 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.49 $Y=1.35 $X2=3.56
+ $Y2=1.35
r85 46 47 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.13 $Y=1.35
+ $X2=3.49 $Y2=1.35
r86 45 46 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.06 $Y=1.35 $X2=3.13
+ $Y2=1.35
r87 44 45 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.7 $Y=1.35 $X2=3.06
+ $Y2=1.35
r88 43 44 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.63 $Y=1.35 $X2=2.7
+ $Y2=1.35
r89 41 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.29 $Y=1.35
+ $X2=2.63 $Y2=1.35
r90 41 42 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.35 $X2=2.29 $Y2=1.35
r91 39 41 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.27 $Y=1.35 $X2=2.29
+ $Y2=1.35
r92 37 39 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.2 $Y=1.35 $X2=2.27
+ $Y2=1.35
r93 32 50 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.65
+ $Y=1.35 $X2=3.65 $Y2=1.35
r94 31 32 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.322
+ $X2=3.6 $Y2=1.322
r95 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.322
+ $X2=3.12 $Y2=1.322
r96 30 42 17.9269 $w=2.23e-07 $l=3.5e-07 $layer=LI1_cond $X=2.64 $Y=1.322
+ $X2=2.29 $Y2=1.322
r97 29 42 6.65856 $w=2.23e-07 $l=1.3e-07 $layer=LI1_cond $X=2.16 $Y=1.322
+ $X2=2.29 $Y2=1.322
r98 25 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=1.515
+ $X2=3.56 $Y2=1.35
r99 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.56 $Y=1.515
+ $X2=3.56 $Y2=2.465
r100 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=1.185
+ $X2=3.49 $Y2=1.35
r101 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.49 $Y=1.185
+ $X2=3.49 $Y2=0.655
r102 18 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.13 $Y=1.515
+ $X2=3.13 $Y2=1.35
r103 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.13 $Y=1.515
+ $X2=3.13 $Y2=2.465
r104 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.185
+ $X2=3.06 $Y2=1.35
r105 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.06 $Y=1.185
+ $X2=3.06 $Y2=0.655
r106 11 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.515
+ $X2=2.7 $Y2=1.35
r107 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.7 $Y=1.515
+ $X2=2.7 $Y2=2.465
r108 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.63 $Y=1.185
+ $X2=2.63 $Y2=1.35
r109 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.63 $Y=1.185
+ $X2=2.63 $Y2=0.655
r110 4 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.515
+ $X2=2.27 $Y2=1.35
r111 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.27 $Y=1.515
+ $X2=2.27 $Y2=2.465
r112 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.185
+ $X2=2.2 $Y2=1.35
r113 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.2 $Y=1.185 $X2=2.2
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%A1 3 7 9 11 14 16 18 19 21 24 26 28 29 30 31
+ 32 49
c72 49 0 1.00341e-19 $X=5.73 $Y=1.425
r73 47 49 18.7792 $w=4.62e-07 $l=1.8e-07 $layer=POLY_cond $X=5.55 $Y=1.425
+ $X2=5.73 $Y2=1.425
r74 45 47 15.6494 $w=4.62e-07 $l=1.5e-07 $layer=POLY_cond $X=5.4 $Y=1.425
+ $X2=5.55 $Y2=1.425
r75 44 45 44.8615 $w=4.62e-07 $l=4.3e-07 $layer=POLY_cond $X=4.97 $Y=1.425
+ $X2=5.4 $Y2=1.425
r76 43 44 1.04329 $w=4.62e-07 $l=1e-08 $layer=POLY_cond $X=4.96 $Y=1.425
+ $X2=4.97 $Y2=1.425
r77 42 43 43.8182 $w=4.62e-07 $l=4.2e-07 $layer=POLY_cond $X=4.54 $Y=1.425
+ $X2=4.96 $Y2=1.425
r78 41 42 1.04329 $w=4.62e-07 $l=1e-08 $layer=POLY_cond $X=4.53 $Y=1.425
+ $X2=4.54 $Y2=1.425
r79 39 41 35.4719 $w=4.62e-07 $l=3.4e-07 $layer=POLY_cond $X=4.19 $Y=1.425
+ $X2=4.53 $Y2=1.425
r80 39 40 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.19
+ $Y=1.35 $X2=4.19 $Y2=1.35
r81 37 39 9.38961 $w=4.62e-07 $l=9e-08 $layer=POLY_cond $X=4.1 $Y=1.425 $X2=4.19
+ $Y2=1.425
r82 32 47 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.55
+ $Y=1.35 $X2=5.55 $Y2=1.35
r83 31 32 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.322
+ $X2=5.52 $Y2=1.322
r84 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.322
+ $X2=5.04 $Y2=1.322
r85 30 40 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=4.56 $Y=1.322
+ $X2=4.19 $Y2=1.322
r86 29 40 5.63417 $w=2.23e-07 $l=1.1e-07 $layer=LI1_cond $X=4.08 $Y=1.322
+ $X2=4.19 $Y2=1.322
r87 26 49 10.4329 $w=4.62e-07 $l=2.85657e-07 $layer=POLY_cond $X=5.83 $Y=1.185
+ $X2=5.73 $Y2=1.425
r88 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.83 $Y=1.185
+ $X2=5.83 $Y2=0.655
r89 22 49 29.4226 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.73 $Y=1.665
+ $X2=5.73 $Y2=1.425
r90 22 24 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.73 $Y=1.665 $X2=5.73
+ $Y2=2.465
r91 19 45 29.4226 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.4 $Y=1.185 $X2=5.4
+ $Y2=1.425
r92 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.4 $Y=1.185 $X2=5.4
+ $Y2=0.655
r93 16 44 29.4226 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.97 $Y=1.185
+ $X2=4.97 $Y2=1.425
r94 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.97 $Y=1.185
+ $X2=4.97 $Y2=0.655
r95 12 43 29.4226 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.96 $Y=1.665
+ $X2=4.96 $Y2=1.425
r96 12 14 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.96 $Y=1.665 $X2=4.96
+ $Y2=2.465
r97 9 42 29.4226 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.54 $Y=1.185
+ $X2=4.54 $Y2=1.425
r98 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.54 $Y=1.185
+ $X2=4.54 $Y2=0.655
r99 5 41 29.4226 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.53 $Y=1.665
+ $X2=4.53 $Y2=1.425
r100 5 7 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.53 $Y=1.665 $X2=4.53
+ $Y2=2.465
r101 1 37 29.4226 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.1 $Y=1.665 $X2=4.1
+ $Y2=1.425
r102 1 3 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.1 $Y=1.665 $X2=4.1
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%A2 1 3 4 6 7 9 12 14 16 19 21 23 26 28 29 30
+ 31 47
c81 31 0 1.00341e-19 $X=7.92 $Y=1.295
r82 47 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=7.79
+ $Y=1.35 $X2=7.79 $Y2=1.35
r83 45 47 34.3264 $w=3.37e-07 $l=2.4e-07 $layer=POLY_cond $X=7.55 $Y=1.455
+ $X2=7.79 $Y2=1.455
r84 39 41 37.1869 $w=3.37e-07 $l=2.6e-07 $layer=POLY_cond $X=6.43 $Y=1.455
+ $X2=6.69 $Y2=1.455
r85 37 39 24.3145 $w=3.37e-07 $l=1.7e-07 $layer=POLY_cond $X=6.26 $Y=1.455
+ $X2=6.43 $Y2=1.455
r86 31 48 6.65856 $w=2.23e-07 $l=1.3e-07 $layer=LI1_cond $X=7.92 $Y=1.322
+ $X2=7.79 $Y2=1.322
r87 30 48 17.9269 $w=2.23e-07 $l=3.5e-07 $layer=LI1_cond $X=7.44 $Y=1.322
+ $X2=7.79 $Y2=1.322
r88 29 30 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.322
+ $X2=7.44 $Y2=1.322
r89 28 29 27.1464 $w=2.23e-07 $l=5.3e-07 $layer=LI1_cond $X=6.43 $Y=1.322
+ $X2=6.96 $Y2=1.322
r90 28 39 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.43
+ $Y=1.35 $X2=6.43 $Y2=1.35
r91 24 47 2.86053 $w=3.37e-07 $l=2e-08 $layer=POLY_cond $X=7.81 $Y=1.455
+ $X2=7.79 $Y2=1.455
r92 24 26 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.81 $Y=1.515
+ $X2=7.81 $Y2=2.465
r93 21 45 21.7231 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.55 $Y=1.185
+ $X2=7.55 $Y2=1.455
r94 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.55 $Y=1.185
+ $X2=7.55 $Y2=0.655
r95 17 45 24.3145 $w=3.37e-07 $l=1.7e-07 $layer=POLY_cond $X=7.38 $Y=1.455
+ $X2=7.55 $Y2=1.455
r96 17 43 37.1869 $w=3.37e-07 $l=2.6e-07 $layer=POLY_cond $X=7.38 $Y=1.455
+ $X2=7.12 $Y2=1.455
r97 17 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.38 $Y=1.515
+ $X2=7.38 $Y2=2.465
r98 14 43 21.7231 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.12 $Y=1.185
+ $X2=7.12 $Y2=1.455
r99 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.12 $Y=1.185
+ $X2=7.12 $Y2=0.655
r100 10 43 24.3145 $w=3.37e-07 $l=1.7e-07 $layer=POLY_cond $X=6.95 $Y=1.455
+ $X2=7.12 $Y2=1.455
r101 10 41 37.1869 $w=3.37e-07 $l=2.6e-07 $layer=POLY_cond $X=6.95 $Y=1.455
+ $X2=6.69 $Y2=1.455
r102 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.95 $Y=1.515
+ $X2=6.95 $Y2=2.465
r103 7 41 21.7231 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.69 $Y=1.185
+ $X2=6.69 $Y2=1.455
r104 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.69 $Y=1.185
+ $X2=6.69 $Y2=0.655
r105 4 37 21.7231 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.26 $Y=1.185
+ $X2=6.26 $Y2=1.455
r106 4 6 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.26 $Y=1.185
+ $X2=6.26 $Y2=0.655
r107 1 37 14.3027 $w=3.37e-07 $l=3.1607e-07 $layer=POLY_cond $X=6.16 $Y=1.725
+ $X2=6.26 $Y2=1.455
r108 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.16 $Y=1.725
+ $X2=6.16 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%A3 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 33 39 41
r76 53 54 30.867 $w=4.06e-07 $l=2.6e-07 $layer=POLY_cond $X=9.53 $Y=1.425
+ $X2=9.79 $Y2=1.425
r77 52 53 20.1823 $w=4.06e-07 $l=1.7e-07 $layer=POLY_cond $X=9.36 $Y=1.425
+ $X2=9.53 $Y2=1.425
r78 51 52 30.867 $w=4.06e-07 $l=2.6e-07 $layer=POLY_cond $X=9.1 $Y=1.425
+ $X2=9.36 $Y2=1.425
r79 50 51 20.1823 $w=4.06e-07 $l=1.7e-07 $layer=POLY_cond $X=8.93 $Y=1.425
+ $X2=9.1 $Y2=1.425
r80 49 50 30.867 $w=4.06e-07 $l=2.6e-07 $layer=POLY_cond $X=8.67 $Y=1.425
+ $X2=8.93 $Y2=1.425
r81 47 49 9.49754 $w=4.06e-07 $l=8e-08 $layer=POLY_cond $X=8.59 $Y=1.425
+ $X2=8.67 $Y2=1.425
r82 47 48 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=8.59
+ $Y=1.35 $X2=8.59 $Y2=1.35
r83 45 47 10.6847 $w=4.06e-07 $l=9e-08 $layer=POLY_cond $X=8.5 $Y=1.425 $X2=8.59
+ $Y2=1.425
r84 39 54 10.7347 $w=4.06e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.865 $Y=1.35
+ $X2=9.79 $Y2=1.425
r85 39 41 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=9.865 $Y=1.35
+ $X2=10.29 $Y2=1.35
r86 33 41 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=10.29
+ $Y=1.35 $X2=10.29 $Y2=1.35
r87 32 33 23.0489 $w=2.23e-07 $l=4.5e-07 $layer=LI1_cond $X=9.84 $Y=1.322
+ $X2=10.29 $Y2=1.322
r88 31 32 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.322
+ $X2=9.84 $Y2=1.322
r89 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.322
+ $X2=9.36 $Y2=1.322
r90 30 48 14.8537 $w=2.23e-07 $l=2.9e-07 $layer=LI1_cond $X=8.88 $Y=1.322
+ $X2=8.59 $Y2=1.322
r91 29 48 9.73174 $w=2.23e-07 $l=1.9e-07 $layer=LI1_cond $X=8.4 $Y=1.322
+ $X2=8.59 $Y2=1.322
r92 26 54 26.2263 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.79 $Y=1.185
+ $X2=9.79 $Y2=1.425
r93 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.79 $Y=1.185
+ $X2=9.79 $Y2=0.655
r94 22 53 26.2263 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.53 $Y=1.665
+ $X2=9.53 $Y2=1.425
r95 22 24 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=9.53 $Y=1.665 $X2=9.53
+ $Y2=2.465
r96 19 52 26.2263 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.36 $Y=1.185
+ $X2=9.36 $Y2=1.425
r97 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.36 $Y=1.185
+ $X2=9.36 $Y2=0.655
r98 15 51 26.2263 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.1 $Y=1.665 $X2=9.1
+ $Y2=1.425
r99 15 17 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=9.1 $Y=1.665 $X2=9.1
+ $Y2=2.465
r100 12 50 26.2263 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.93 $Y=1.185
+ $X2=8.93 $Y2=1.425
r101 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.93 $Y=1.185
+ $X2=8.93 $Y2=0.655
r102 8 49 26.2263 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.67 $Y=1.665
+ $X2=8.67 $Y2=1.425
r103 8 10 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=8.67 $Y=1.665 $X2=8.67
+ $Y2=2.465
r104 5 45 26.2263 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.5 $Y=1.185 $X2=8.5
+ $Y2=1.425
r105 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.5 $Y=1.185 $X2=8.5
+ $Y2=0.655
r106 1 45 30.867 $w=4.06e-07 $l=3.60555e-07 $layer=POLY_cond $X=8.24 $Y=1.665
+ $X2=8.5 $Y2=1.425
r107 1 3 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=8.24 $Y=1.665 $X2=8.24
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%A_42_367# 1 2 3 4 5 6 7 8 9 10 11 34 36 38
+ 42 44 48 50 54 56 58 59 60 64 66 70 72 77 80 82 83 86 90 94 98 102 109 111 113
+ 119 121 122 123 124
r139 102 104 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=9.78 $Y=1.98
+ $X2=9.78 $Y2=2.91
r140 100 102 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=9.78 $Y=1.775
+ $X2=9.78 $Y2=1.98
r141 99 124 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.98 $Y=1.69
+ $X2=8.885 $Y2=1.69
r142 98 100 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.65 $Y=1.69
+ $X2=9.78 $Y2=1.775
r143 98 99 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.65 $Y=1.69
+ $X2=8.98 $Y2=1.69
r144 94 96 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=8.885 $Y=1.98
+ $X2=8.885 $Y2=2.91
r145 92 124 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=1.775
+ $X2=8.885 $Y2=1.69
r146 92 94 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=8.885 $Y=1.775
+ $X2=8.885 $Y2=1.98
r147 91 123 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.12 $Y=1.69
+ $X2=8.025 $Y2=1.69
r148 90 124 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.79 $Y=1.69
+ $X2=8.885 $Y2=1.69
r149 90 91 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.79 $Y=1.69
+ $X2=8.12 $Y2=1.69
r150 86 88 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=8.025 $Y=1.96
+ $X2=8.025 $Y2=2.91
r151 84 123 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.025 $Y=1.775
+ $X2=8.025 $Y2=1.69
r152 84 86 10.799 $w=1.88e-07 $l=1.85e-07 $layer=LI1_cond $X=8.025 $Y=1.775
+ $X2=8.025 $Y2=1.96
r153 82 123 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.93 $Y=1.69
+ $X2=8.025 $Y2=1.69
r154 82 83 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.93 $Y=1.69
+ $X2=7.26 $Y2=1.69
r155 78 122 4.27425 $w=2.25e-07 $l=1.06066e-07 $layer=LI1_cond $X=7.165 $Y=2.225
+ $X2=7.13 $Y2=2.135
r156 78 80 14.0096 $w=1.88e-07 $l=2.4e-07 $layer=LI1_cond $X=7.165 $Y=2.225
+ $X2=7.165 $Y2=2.465
r157 75 122 4.27425 $w=2.25e-07 $l=9e-08 $layer=LI1_cond $X=7.13 $Y=2.045
+ $X2=7.13 $Y2=2.135
r158 75 77 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=7.13 $Y=2.045
+ $X2=7.13 $Y2=1.96
r159 74 83 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.13 $Y=1.775
+ $X2=7.26 $Y2=1.69
r160 74 77 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=7.13 $Y=1.775
+ $X2=7.13 $Y2=1.96
r161 73 121 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.04 $Y=2.135
+ $X2=5.945 $Y2=2.135
r162 72 122 2.15711 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=7 $Y=2.135 $X2=7.13
+ $Y2=2.135
r163 72 73 59.1515 $w=1.78e-07 $l=9.6e-07 $layer=LI1_cond $X=7 $Y=2.135 $X2=6.04
+ $Y2=2.135
r164 68 121 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=5.945 $Y=2.225
+ $X2=5.945 $Y2=2.135
r165 68 70 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=5.945 $Y=2.225
+ $X2=5.945 $Y2=2.91
r166 67 119 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.84 $Y=2.135
+ $X2=4.745 $Y2=2.135
r167 66 121 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.85 $Y=2.135
+ $X2=5.945 $Y2=2.135
r168 66 67 62.2323 $w=1.78e-07 $l=1.01e-06 $layer=LI1_cond $X=5.85 $Y=2.135
+ $X2=4.84 $Y2=2.135
r169 62 119 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=4.745 $Y=2.225
+ $X2=4.745 $Y2=2.135
r170 62 64 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=4.745 $Y=2.225
+ $X2=4.745 $Y2=2.91
r171 61 115 4.61608 $w=1.8e-07 $l=1.5e-07 $layer=LI1_cond $X=3.98 $Y=2.135
+ $X2=3.83 $Y2=2.135
r172 60 119 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.65 $Y=2.135
+ $X2=4.745 $Y2=2.135
r173 60 61 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.65 $Y=2.135
+ $X2=3.98 $Y2=2.135
r174 59 117 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.83 $Y=2.905
+ $X2=3.83 $Y2=2.99
r175 58 115 2.76965 $w=3e-07 $l=9e-08 $layer=LI1_cond $X=3.83 $Y=2.225 $X2=3.83
+ $Y2=2.135
r176 58 59 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=3.83 $Y=2.225
+ $X2=3.83 $Y2=2.905
r177 57 113 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.01 $Y=2.99
+ $X2=2.915 $Y2=2.99
r178 56 117 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.68 $Y=2.99
+ $X2=3.83 $Y2=2.99
r179 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.68 $Y=2.99
+ $X2=3.01 $Y2=2.99
r180 52 113 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=2.905
+ $X2=2.915 $Y2=2.99
r181 52 54 40.5694 $w=1.88e-07 $l=6.95e-07 $layer=LI1_cond $X=2.915 $Y=2.905
+ $X2=2.915 $Y2=2.21
r182 51 111 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.15 $Y=2.99
+ $X2=2.055 $Y2=2.99
r183 50 113 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.82 $Y=2.99
+ $X2=2.915 $Y2=2.99
r184 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.82 $Y=2.99
+ $X2=2.15 $Y2=2.99
r185 46 111 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.905
+ $X2=2.055 $Y2=2.99
r186 46 48 40.5694 $w=1.88e-07 $l=6.95e-07 $layer=LI1_cond $X=2.055 $Y=2.905
+ $X2=2.055 $Y2=2.21
r187 45 109 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.29 $Y=2.99
+ $X2=1.195 $Y2=2.99
r188 44 111 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.96 $Y=2.99
+ $X2=2.055 $Y2=2.99
r189 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.96 $Y=2.99
+ $X2=1.29 $Y2=2.99
r190 40 109 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=2.905
+ $X2=1.195 $Y2=2.99
r191 40 42 40.5694 $w=1.88e-07 $l=6.95e-07 $layer=LI1_cond $X=1.195 $Y=2.905
+ $X2=1.195 $Y2=2.21
r192 39 107 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.43 $Y=2.99
+ $X2=0.3 $Y2=2.99
r193 38 109 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.1 $Y=2.99
+ $X2=1.195 $Y2=2.99
r194 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.1 $Y=2.99
+ $X2=0.43 $Y2=2.99
r195 34 107 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.3 $Y=2.905
+ $X2=0.3 $Y2=2.99
r196 34 36 40.5571 $w=2.58e-07 $l=9.15e-07 $layer=LI1_cond $X=0.3 $Y=2.905
+ $X2=0.3 $Y2=1.99
r197 11 104 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.605
+ $Y=1.835 $X2=9.745 $Y2=2.91
r198 11 102 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.605
+ $Y=1.835 $X2=9.745 $Y2=1.98
r199 10 96 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.835 $X2=8.885 $Y2=2.91
r200 10 94 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.835 $X2=8.885 $Y2=1.98
r201 9 88 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.835 $X2=8.025 $Y2=2.91
r202 9 86 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.835 $X2=8.025 $Y2=1.96
r203 8 80 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=7.025
+ $Y=1.835 $X2=7.165 $Y2=2.465
r204 8 77 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=1.835 $X2=7.165 $Y2=1.96
r205 7 121 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.835 $X2=5.945 $Y2=2.21
r206 7 70 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.835 $X2=5.945 $Y2=2.91
r207 6 119 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=4.605
+ $Y=1.835 $X2=4.745 $Y2=2.21
r208 6 64 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.605
+ $Y=1.835 $X2=4.745 $Y2=2.91
r209 5 117 400 $w=1.7e-07 $l=1.16844e-06 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.835 $X2=3.83 $Y2=2.91
r210 5 115 400 $w=1.7e-07 $l=4.62331e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.835 $X2=3.83 $Y2=2.21
r211 4 113 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.915 $Y2=2.91
r212 4 54 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.915 $Y2=2.21
r213 3 111 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.91
r214 3 48 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.21
r215 2 109 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.835 $X2=1.195 $Y2=2.91
r216 2 42 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.835 $X2=1.195 $Y2=2.21
r217 1 107 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=1.835 $X2=0.335 $Y2=2.91
r218 1 36 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=1.835 $X2=0.335 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%Y 1 2 3 4 5 6 7 8 27 31 32 35 39 43 47 51 55
+ 57 58 59 60 61 62 63 64 65 66 72
c136 55 0 1.99728e-19 $X=5.885 $Y=1.74
r137 74 77 36.04 $w=2.73e-07 $l=8.6e-07 $layer=LI1_cond $X=2.415 $Y=0.902
+ $X2=3.275 $Y2=0.902
r138 72 89 11.3149 $w=2.73e-07 $l=2.7e-07 $layer=LI1_cond $X=5.885 $Y=0.902
+ $X2=5.615 $Y2=0.902
r139 66 72 3.01473 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=5.99 $Y=0.902
+ $X2=5.885 $Y2=0.902
r140 65 89 3.98117 $w=2.73e-07 $l=9.5e-08 $layer=LI1_cond $X=5.52 $Y=0.902
+ $X2=5.615 $Y2=0.902
r141 64 65 20.1154 $w=2.73e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=0.902
+ $X2=5.52 $Y2=0.902
r142 64 83 11.9435 $w=2.73e-07 $l=2.85e-07 $layer=LI1_cond $X=5.04 $Y=0.902
+ $X2=4.755 $Y2=0.902
r143 63 83 8.17187 $w=2.73e-07 $l=1.95e-07 $layer=LI1_cond $X=4.56 $Y=0.902
+ $X2=4.755 $Y2=0.902
r144 62 63 20.1154 $w=2.73e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=0.902
+ $X2=4.56 $Y2=0.902
r145 62 77 33.7351 $w=2.73e-07 $l=8.05e-07 $layer=LI1_cond $X=4.08 $Y=0.902
+ $X2=3.275 $Y2=0.902
r146 57 66 3.96222 $w=2.1e-07 $l=1.38e-07 $layer=LI1_cond $X=5.99 $Y=1.04
+ $X2=5.99 $Y2=0.902
r147 57 58 29.8398 $w=2.08e-07 $l=5.65e-07 $layer=LI1_cond $X=5.99 $Y=1.04
+ $X2=5.99 $Y2=1.605
r148 56 61 6.08426 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.51 $Y=1.74
+ $X2=3.345 $Y2=1.74
r149 55 58 6.95594 $w=2.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.885 $Y=1.74
+ $X2=5.99 $Y2=1.605
r150 55 56 101.372 $w=2.68e-07 $l=2.375e-06 $layer=LI1_cond $X=5.885 $Y=1.74
+ $X2=3.51 $Y2=1.74
r151 51 53 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.345 $Y=1.97
+ $X2=3.345 $Y2=2.65
r152 49 61 0.630948 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=3.345 $Y=1.875
+ $X2=3.345 $Y2=1.74
r153 49 51 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.345 $Y=1.875
+ $X2=3.345 $Y2=1.97
r154 48 60 6.08426 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=1.74
+ $X2=2.485 $Y2=1.74
r155 47 61 6.08426 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=1.74
+ $X2=3.345 $Y2=1.74
r156 47 48 22.622 $w=2.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.18 $Y=1.74
+ $X2=2.65 $Y2=1.74
r157 43 45 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.485 $Y=1.97
+ $X2=2.485 $Y2=2.65
r158 41 60 0.630948 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=2.485 $Y=1.875
+ $X2=2.485 $Y2=1.74
r159 41 43 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.485 $Y=1.875
+ $X2=2.485 $Y2=1.97
r160 40 59 6.08426 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=1.74
+ $X2=1.625 $Y2=1.74
r161 39 60 6.08426 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=1.74
+ $X2=2.485 $Y2=1.74
r162 39 40 22.622 $w=2.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.32 $Y=1.74
+ $X2=1.79 $Y2=1.74
r163 35 37 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.625 $Y=1.97
+ $X2=1.625 $Y2=2.65
r164 33 59 0.630948 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=1.625 $Y=1.875
+ $X2=1.625 $Y2=1.74
r165 33 35 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.625 $Y=1.875
+ $X2=1.625 $Y2=1.97
r166 31 59 6.08426 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=1.74
+ $X2=1.625 $Y2=1.74
r167 31 32 22.622 $w=2.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.46 $Y=1.74
+ $X2=0.93 $Y2=1.74
r168 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.765 $Y=1.97
+ $X2=0.765 $Y2=2.65
r169 25 32 6.90553 $w=2.7e-07 $l=2.22486e-07 $layer=LI1_cond $X=0.765 $Y=1.875
+ $X2=0.93 $Y2=1.74
r170 25 27 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.765 $Y=1.875
+ $X2=0.765 $Y2=1.97
r171 8 53 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.835 $X2=3.345 $Y2=2.65
r172 8 51 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.835 $X2=3.345 $Y2=1.97
r173 7 45 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.835 $X2=2.485 $Y2=2.65
r174 7 43 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.835 $X2=2.485 $Y2=1.97
r175 6 37 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=2.65
r176 6 35 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=1.97
r177 5 29 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.835 $X2=0.765 $Y2=2.65
r178 5 27 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.835 $X2=0.765 $Y2=1.97
r179 4 89 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=5.475
+ $Y=0.235 $X2=5.615 $Y2=0.925
r180 3 83 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.235 $X2=4.755 $Y2=0.925
r181 2 77 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=3.135
+ $Y=0.235 $X2=3.275 $Y2=0.925
r182 1 74 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.235 $X2=2.415 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%VPWR 1 2 3 4 5 6 21 23 27 31 33 37 43 49 53
+ 54 55 64 69 74 81 82 85 90 93 96 99
r142 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r143 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r144 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r145 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r146 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r147 85 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r148 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r149 82 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.36 $Y2=3.33
r150 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r151 79 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.48 $Y=3.33
+ $X2=9.315 $Y2=3.33
r152 79 81 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=9.48 $Y=3.33
+ $X2=10.32 $Y2=3.33
r153 78 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r154 78 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r156 75 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=3.33
+ $X2=8.455 $Y2=3.33
r157 75 77 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.62 $Y=3.33
+ $X2=8.88 $Y2=3.33
r158 74 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.15 $Y=3.33
+ $X2=9.315 $Y2=3.33
r159 74 77 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.15 $Y=3.33
+ $X2=8.88 $Y2=3.33
r160 73 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r161 73 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r162 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r163 70 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=3.33
+ $X2=7.595 $Y2=3.33
r164 70 72 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=3.33
+ $X2=7.92 $Y2=3.33
r165 69 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.29 $Y=3.33
+ $X2=8.455 $Y2=3.33
r166 69 72 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.29 $Y=3.33
+ $X2=7.92 $Y2=3.33
r167 68 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r168 68 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r169 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r170 65 85 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=5.68 $Y=3.33
+ $X2=5.345 $Y2=3.33
r171 65 67 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.68 $Y=3.33 $X2=6
+ $Y2=3.33
r172 64 90 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=6.21 $Y=3.33
+ $X2=6.555 $Y2=3.33
r173 64 67 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.21 $Y=3.33 $X2=6
+ $Y2=3.33
r174 63 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r175 62 63 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r176 59 63 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r177 58 62 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r178 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r179 55 86 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r180 55 88 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r181 53 62 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.15 $Y=3.33 $X2=4.08
+ $Y2=3.33
r182 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=4.315 $Y2=3.33
r183 49 52 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=9.315 $Y=2.03
+ $X2=9.315 $Y2=2.95
r184 47 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.315 $Y=3.245
+ $X2=9.315 $Y2=3.33
r185 47 52 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.315 $Y=3.245
+ $X2=9.315 $Y2=2.95
r186 43 46 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=8.455 $Y=2.03
+ $X2=8.455 $Y2=2.95
r187 41 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.455 $Y=3.245
+ $X2=8.455 $Y2=3.33
r188 41 46 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.455 $Y=3.245
+ $X2=8.455 $Y2=2.95
r189 37 40 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=7.595 $Y=2.03
+ $X2=7.595 $Y2=2.95
r190 35 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.595 $Y=3.245
+ $X2=7.595 $Y2=3.33
r191 35 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.595 $Y=3.245
+ $X2=7.595 $Y2=2.95
r192 34 90 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=6.9 $Y=3.33
+ $X2=6.555 $Y2=3.33
r193 33 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=3.33
+ $X2=7.595 $Y2=3.33
r194 33 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.43 $Y=3.33
+ $X2=6.9 $Y2=3.33
r195 29 90 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=3.245
+ $X2=6.555 $Y2=3.33
r196 29 31 12.9142 $w=6.88e-07 $l=7.45e-07 $layer=LI1_cond $X=6.555 $Y=3.245
+ $X2=6.555 $Y2=2.5
r197 25 85 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=3.245
+ $X2=5.345 $Y2=3.33
r198 25 27 12.4963 $w=6.68e-07 $l=7e-07 $layer=LI1_cond $X=5.345 $Y=3.245
+ $X2=5.345 $Y2=2.545
r199 24 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.48 $Y=3.33
+ $X2=4.315 $Y2=3.33
r200 23 85 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=5.345 $Y2=3.33
r201 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=4.48 $Y2=3.33
r202 19 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=3.245
+ $X2=4.315 $Y2=3.33
r203 19 21 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.315 $Y=3.245
+ $X2=4.315 $Y2=2.5
r204 6 52 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.835 $X2=9.315 $Y2=2.95
r205 6 49 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.835 $X2=9.315 $Y2=2.03
r206 5 46 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.315
+ $Y=1.835 $X2=8.455 $Y2=2.95
r207 5 43 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=8.315
+ $Y=1.835 $X2=8.455 $Y2=2.03
r208 4 40 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.455
+ $Y=1.835 $X2=7.595 $Y2=2.95
r209 4 37 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=7.455
+ $Y=1.835 $X2=7.595 $Y2=2.03
r210 3 31 150 $w=1.7e-07 $l=8.80185e-07 $layer=licon1_PDIFF $count=4 $X=6.235
+ $Y=1.835 $X2=6.735 $Y2=2.5
r211 2 27 150 $w=1.7e-07 $l=9.19184e-07 $layer=licon1_PDIFF $count=4 $X=5.035
+ $Y=1.835 $X2=5.515 $Y2=2.545
r212 1 21 300 $w=1.7e-07 $l=7.31659e-07 $layer=licon1_PDIFF $count=2 $X=4.175
+ $Y=1.835 $X2=4.315 $Y2=2.5
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%A_28_47# 1 2 3 4 5 18 20 21 24 26 28 29 34
+ 36
r45 32 34 29.15 $w=3.38e-07 $l=8.6e-07 $layer=LI1_cond $X=2.845 $Y=0.425
+ $X2=3.705 $Y2=0.425
r46 30 38 2.70725 $w=3.4e-07 $l=9.5e-08 $layer=LI1_cond $X=2.08 $Y=0.425
+ $X2=1.985 $Y2=0.425
r47 30 32 25.93 $w=3.38e-07 $l=7.65e-07 $layer=LI1_cond $X=2.08 $Y=0.425
+ $X2=2.845 $Y2=0.425
r48 29 40 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.87
+ $X2=1.985 $Y2=0.955
r49 28 38 4.84456 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=1.985 $Y=0.595
+ $X2=1.985 $Y2=0.425
r50 28 29 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=1.985 $Y=0.595
+ $X2=1.985 $Y2=0.87
r51 27 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.22 $Y=0.955
+ $X2=1.125 $Y2=0.955
r52 26 40 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.89 $Y=0.955
+ $X2=1.985 $Y2=0.955
r53 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.89 $Y=0.955
+ $X2=1.22 $Y2=0.955
r54 22 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.87
+ $X2=1.125 $Y2=0.955
r55 22 24 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=1.125 $Y=0.87
+ $X2=1.125 $Y2=0.42
r56 20 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.03 $Y=0.955
+ $X2=1.125 $Y2=0.955
r57 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.03 $Y=0.955
+ $X2=0.36 $Y2=0.955
r58 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.23 $Y=0.87
+ $X2=0.36 $Y2=0.955
r59 16 18 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=0.23 $Y=0.87
+ $X2=0.23 $Y2=0.42
r60 5 34 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=3.565
+ $Y=0.235 $X2=3.705 $Y2=0.43
r61 4 32 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.705
+ $Y=0.235 $X2=2.845 $Y2=0.43
r62 3 40 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.235 $X2=1.985 $Y2=0.875
r63 3 38 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.235 $X2=1.985 $Y2=0.42
r64 2 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.235 $X2=1.125 $Y2=0.42
r65 1 18 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%VGND 1 2 3 4 5 18 22 26 30 32 36 39 40 41 42
+ 43 45 50 64 65 68 71 74
r119 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r120 71 72 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r121 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r122 65 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r123 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r124 62 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.17 $Y=0
+ $X2=10.005 $Y2=0
r125 62 64 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=10.17 $Y=0 $X2=10.32
+ $Y2=0
r126 61 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r127 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r128 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r129 57 58 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r130 55 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=0 $X2=1.555
+ $Y2=0
r131 55 57 404.492 $w=1.68e-07 $l=6.2e-06 $layer=LI1_cond $X=1.72 $Y=0 $X2=7.92
+ $Y2=0
r132 54 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r133 54 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r134 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r135 51 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=0.695
+ $Y2=0
r136 51 53 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=1.2
+ $Y2=0
r137 50 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.555
+ $Y2=0
r138 50 53 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.2
+ $Y2=0
r139 48 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r140 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r141 45 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.695
+ $Y2=0
r142 45 47 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.24
+ $Y2=0
r143 43 58 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=7.92
+ $Y2=0
r144 43 72 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=1.68
+ $Y2=0
r145 41 60 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=8.98 $Y=0 $X2=8.88
+ $Y2=0
r146 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.98 $Y=0 $X2=9.145
+ $Y2=0
r147 39 57 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=8.12 $Y=0 $X2=7.92
+ $Y2=0
r148 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.12 $Y=0 $X2=8.285
+ $Y2=0
r149 38 60 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.45 $Y=0 $X2=8.88
+ $Y2=0
r150 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.45 $Y=0 $X2=8.285
+ $Y2=0
r151 34 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.005 $Y=0.085
+ $X2=10.005 $Y2=0
r152 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.005 $Y=0.085
+ $X2=10.005 $Y2=0.38
r153 33 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.31 $Y=0 $X2=9.145
+ $Y2=0
r154 32 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.84 $Y=0
+ $X2=10.005 $Y2=0
r155 32 33 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=9.84 $Y=0 $X2=9.31
+ $Y2=0
r156 28 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=0.085
+ $X2=9.145 $Y2=0
r157 28 30 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=9.145 $Y=0.085
+ $X2=9.145 $Y2=0.465
r158 24 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.285 $Y=0.085
+ $X2=8.285 $Y2=0
r159 24 26 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=8.285 $Y=0.085
+ $X2=8.285 $Y2=0.465
r160 20 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=0.085
+ $X2=1.555 $Y2=0
r161 20 22 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.555 $Y=0.085
+ $X2=1.555 $Y2=0.56
r162 16 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0
r163 16 18 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0.56
r164 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.865
+ $Y=0.235 $X2=10.005 $Y2=0.38
r165 4 30 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=9.005
+ $Y=0.235 $X2=9.145 $Y2=0.465
r166 3 26 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=8.16
+ $Y=0.235 $X2=8.285 $Y2=0.465
r167 2 22 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.235 $X2=1.555 $Y2=0.56
r168 1 18 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.235 $X2=0.695 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%A_840_47# 1 2 3 4 5 26
r33 24 26 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=6.905 $Y=0.43
+ $X2=7.765 $Y2=0.43
r34 22 24 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=6.045 $Y=0.43
+ $X2=6.905 $Y2=0.43
r35 20 22 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.185 $Y=0.43
+ $X2=6.045 $Y2=0.43
r36 17 20 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.325 $Y=0.43
+ $X2=5.185 $Y2=0.43
r37 5 26 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=7.625
+ $Y=0.235 $X2=7.765 $Y2=0.43
r38 4 24 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=6.765
+ $Y=0.235 $X2=6.905 $Y2=0.43
r39 3 22 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.235 $X2=6.045 $Y2=0.43
r40 2 20 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.235 $X2=5.185 $Y2=0.43
r41 1 17 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.235 $X2=4.325 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_4%A_1267_47# 1 2 3 4 13 21 23 27 30
r39 25 27 23.0574 $w=1.88e-07 $l=3.95e-07 $layer=LI1_cond $X=9.575 $Y=0.815
+ $X2=9.575 $Y2=0.42
r40 24 30 4.08801 $w=2.5e-07 $l=1.06771e-07 $layer=LI1_cond $X=8.81 $Y=0.927
+ $X2=8.715 $Y2=0.902
r41 23 25 6.87974 $w=2.25e-07 $l=1.52263e-07 $layer=LI1_cond $X=9.48 $Y=0.927
+ $X2=9.575 $Y2=0.815
r42 23 24 34.3172 $w=2.23e-07 $l=6.7e-07 $layer=LI1_cond $X=9.48 $Y=0.927
+ $X2=8.81 $Y2=0.927
r43 19 30 2.34704 $w=1.9e-07 $l=1.37e-07 $layer=LI1_cond $X=8.715 $Y=0.765
+ $X2=8.715 $Y2=0.902
r44 19 21 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=8.715 $Y=0.765
+ $X2=8.715 $Y2=0.42
r45 15 18 36.04 $w=2.73e-07 $l=8.6e-07 $layer=LI1_cond $X=6.475 $Y=0.902
+ $X2=7.335 $Y2=0.902
r46 13 30 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=8.62 $Y=0.902
+ $X2=8.715 $Y2=0.902
r47 13 18 53.8505 $w=2.73e-07 $l=1.285e-06 $layer=LI1_cond $X=8.62 $Y=0.902
+ $X2=7.335 $Y2=0.902
r48 4 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.435
+ $Y=0.235 $X2=9.575 $Y2=0.42
r49 3 30 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=8.575
+ $Y=0.235 $X2=8.715 $Y2=0.875
r50 3 21 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=8.575
+ $Y=0.235 $X2=8.715 $Y2=0.42
r51 2 18 182 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_NDIFF $count=1 $X=7.195
+ $Y=0.235 $X2=7.335 $Y2=0.88
r52 1 15 182 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.235 $X2=6.475 $Y2=0.88
.ends

