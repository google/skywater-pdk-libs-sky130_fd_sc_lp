# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfrbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.570000 0.840000 1.805000 1.495000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.575000 0.255000 13.810000 3.075000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.650000 0.255000 11.915000 3.075000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.325000 1.920000  3.695000 2.200000 ;
        RECT  7.300000 1.825000  7.605000 2.155000 ;
        RECT 10.125000 1.940000 10.505000 2.300000 ;
      LAYER mcon ;
        RECT  3.515000 1.950000  3.685000 2.120000 ;
        RECT  7.355000 1.950000  7.525000 2.120000 ;
        RECT 10.205000 1.950000 10.375000 2.120000 ;
      LAYER met1 ;
        RECT  3.455000 1.920000  3.745000 1.965000 ;
        RECT  3.455000 1.965000 10.435000 2.105000 ;
        RECT  3.455000 2.105000  3.745000 2.150000 ;
        RECT  7.295000 1.920000  7.585000 1.965000 ;
        RECT  7.295000 2.105000  7.585000 2.150000 ;
        RECT 10.145000 1.920000 10.435000 1.965000 ;
        RECT 10.145000 2.105000 10.435000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.565000 2.805000 2.275000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.515000 1.345000 1.675000 ;
        RECT 0.535000 1.675000 2.355000 1.845000 ;
        RECT 2.185000 1.135000 2.515000 1.395000 ;
        RECT 2.185000 1.395000 2.355000 1.675000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.210000 4.175000 1.750000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.400000 0.085000 ;
        RECT  0.525000  0.085000  0.855000 0.765000 ;
        RECT  3.350000  0.085000  3.610000 0.780000 ;
        RECT  4.260000  0.085000  4.590000 0.690000 ;
        RECT  5.260000  0.085000  5.430000 0.905000 ;
        RECT  7.595000  0.085000  7.925000 0.550000 ;
        RECT  9.880000  0.085000 10.210000 0.670000 ;
        RECT 11.190000  0.085000 11.480000 0.900000 ;
        RECT 12.085000  0.085000 12.405000 1.095000 ;
        RECT 13.095000  0.085000 13.405000 1.060000 ;
        RECT 13.980000  0.085000 14.285000 1.140000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 14.400000 3.415000 ;
        RECT  1.050000 2.435000  1.310000 3.245000 ;
        RECT  2.670000 2.835000  3.000000 3.245000 ;
        RECT  4.215000 2.825000  4.545000 3.245000 ;
        RECT  6.690000 2.675000  7.020000 3.245000 ;
        RECT  7.775000 2.085000  8.025000 3.245000 ;
        RECT  9.710000 2.850000 10.455000 3.245000 ;
        RECT 10.105000 2.525000 10.455000 2.850000 ;
        RECT 11.150000 2.280000 11.480000 3.245000 ;
        RECT 12.085000 1.795000 12.405000 3.245000 ;
        RECT 13.095000 1.815000 13.405000 3.245000 ;
        RECT 13.980000 1.815000 14.285000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.095000 0.465000  0.355000 0.935000 ;
      RECT  0.095000 0.935000  1.255000 1.265000 ;
      RECT  0.095000 1.265000  0.365000 2.015000 ;
      RECT  0.095000 2.015000  2.335000 2.195000 ;
      RECT  0.530000 2.195000  2.335000 2.265000 ;
      RECT  0.530000 2.265000  0.880000 3.075000 ;
      RECT  1.115000 0.265000  3.180000 0.435000 ;
      RECT  1.115000 0.435000  1.490000 0.685000 ;
      RECT  1.115000 0.685000  1.415000 0.765000 ;
      RECT  1.770000 2.445000  3.145000 2.485000 ;
      RECT  1.770000 2.485000  5.625000 2.655000 ;
      RECT  1.770000 2.655000  2.100000 3.075000 ;
      RECT  1.975000 0.605000  2.305000 0.795000 ;
      RECT  1.975000 0.795000  3.145000 0.965000 ;
      RECT  2.850000 0.435000  3.180000 0.625000 ;
      RECT  2.975000 0.965000  3.145000 2.445000 ;
      RECT  3.210000 2.655000  3.540000 3.075000 ;
      RECT  3.800000 0.595000  4.060000 0.860000 ;
      RECT  3.800000 0.860000  4.515000 1.040000 ;
      RECT  3.865000 1.930000  4.515000 2.100000 ;
      RECT  3.865000 2.100000  4.115000 2.315000 ;
      RECT  4.345000 1.040000  4.515000 1.280000 ;
      RECT  4.345000 1.280000  4.780000 1.610000 ;
      RECT  4.345000 1.610000  4.515000 1.930000 ;
      RECT  4.685000 1.815000  5.120000 2.145000 ;
      RECT  4.685000 2.145000  5.085000 2.315000 ;
      RECT  4.770000 0.595000  5.090000 1.050000 ;
      RECT  4.770000 1.050000  5.120000 1.075000 ;
      RECT  4.770000 1.075000  5.770000 1.110000 ;
      RECT  4.905000 1.110000  5.770000 1.155000 ;
      RECT  4.950000 1.155000  5.770000 1.780000 ;
      RECT  4.950000 1.780000  5.120000 1.815000 ;
      RECT  5.355000 2.325000  5.625000 2.485000 ;
      RECT  5.390000 1.950000  6.110000 2.120000 ;
      RECT  5.390000 2.120000  5.625000 2.325000 ;
      RECT  5.600000 0.310000  7.425000 0.480000 ;
      RECT  5.600000 0.480000  5.770000 1.075000 ;
      RECT  5.795000 2.290000  6.450000 2.335000 ;
      RECT  5.795000 2.335000  7.565000 2.505000 ;
      RECT  5.795000 2.505000  6.520000 2.695000 ;
      RECT  5.940000 0.650000  6.110000 1.950000 ;
      RECT  6.280000 0.650000  6.620000 0.890000 ;
      RECT  6.280000 0.890000  6.450000 2.290000 ;
      RECT  6.620000 1.060000  8.560000 1.235000 ;
      RECT  6.620000 1.235000  6.790000 2.155000 ;
      RECT  6.960000 1.405000  8.140000 1.645000 ;
      RECT  6.960000 1.645000  7.130000 2.335000 ;
      RECT  7.190000 2.505000  7.565000 2.695000 ;
      RECT  7.245000 0.480000  7.425000 0.720000 ;
      RECT  7.245000 0.720000  8.850000 0.775000 ;
      RECT  7.245000 0.775000  8.900000 0.820000 ;
      RECT  7.245000 0.820000  9.070000 0.890000 ;
      RECT  7.965000 1.645000  8.140000 1.735000 ;
      RECT  8.310000 1.235000  8.560000 2.080000 ;
      RECT  8.310000 2.080000  8.630000 2.910000 ;
      RECT  8.670000 0.890000  9.070000 0.930000 ;
      RECT  8.705000 0.930000  9.070000 0.965000 ;
      RECT  8.730000 0.965000  9.070000 1.700000 ;
      RECT  8.730000 1.700000  9.515000 1.900000 ;
      RECT  8.825000 2.080000  9.105000 2.490000 ;
      RECT  8.825000 2.490000  9.935000 2.670000 ;
      RECT  8.825000 2.670000  9.155000 2.910000 ;
      RECT  9.020000 0.255000  9.445000 0.650000 ;
      RECT  9.240000 0.650000  9.445000 1.360000 ;
      RECT  9.240000 1.360000  9.955000 1.430000 ;
      RECT  9.240000 1.430000 10.875000 1.530000 ;
      RECT  9.275000 1.900000  9.515000 1.990000 ;
      RECT  9.275000 1.990000  9.595000 2.320000 ;
      RECT  9.615000 0.860000 11.000000 1.070000 ;
      RECT  9.615000 1.070000 11.235000 1.190000 ;
      RECT  9.765000 1.530000 10.875000 1.760000 ;
      RECT  9.765000 1.760000  9.935000 2.490000 ;
      RECT 10.125000 1.190000 11.235000 1.260000 ;
      RECT 10.625000 2.470000 10.895000 2.855000 ;
      RECT 10.670000 0.330000 11.000000 0.860000 ;
      RECT 10.675000 1.940000 11.235000 2.110000 ;
      RECT 10.675000 2.110000 10.895000 2.470000 ;
      RECT 11.065000 1.260000 11.235000 1.940000 ;
      RECT 12.575000 0.285000 12.905000 1.230000 ;
      RECT 12.575000 1.230000 13.405000 1.560000 ;
      RECT 12.575000 1.560000 12.885000 2.495000 ;
  END
END sky130_fd_sc_lp__sdfrbp_2
