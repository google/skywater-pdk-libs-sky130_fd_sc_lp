* File: sky130_fd_sc_lp__iso1n_lp.spice
* Created: Fri Aug 28 10:41:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__iso1n_lp.pex.spice"
.subckt sky130_fd_sc_lp__iso1n_lp  VNB VPB SLEEP_B A VPWR X KAGND VGND
* 
* KAGND	KAGND
* X	X
* VPWR	VPWR
* A	A
* SLEEP_B	SLEEP_B
* VPB	VPB
* VNB	VNB
MM1006 A_110_93# N_SLEEP_B_M1006_g N_A_27_93#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1001 N_KAGND_M1001_d N_SLEEP_B_M1001_g A_110_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1011 A_268_93# N_A_27_93#_M1011_g N_KAGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_340_93#_M1007_d N_A_27_93#_M1007_g A_268_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.0714 AS=0.0441 PD=0.76 PS=0.63 NRD=17.136 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1002 A_438_93# N_A_M1002_g N_A_340_93#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0714 PD=0.63 PS=0.76 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_KAGND_M1012_d N_A_M1012_g A_438_93# VNB NSHORT L=0.15 W=0.42 AD=0.0651
+ AS=0.0441 PD=0.73 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1003 A_602_93# N_A_340_93#_M1003_g N_KAGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0651 PD=0.63 PS=0.73 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75002.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_340_93#_M1005_g A_602_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_154_489# N_SLEEP_B_M1004_g N_A_27_93#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1113 PD=0.66 PS=1.37 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_SLEEP_B_M1009_g A_154_489# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=25.7873 NRS=30.4759 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 A_340_489# N_A_27_93#_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=25.7873 M=1 R=2.8
+ SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_340_93#_M1013_d N_A_M1013_g A_340_489# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 A_602_367# N_A_340_93#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_X_M1010_d N_A_340_93#_M1010_g A_602_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.91692 P=12.22
c_29 VNB 0 8.05229e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__iso1n_lp.pxi.spice"
*
.ends
*
*
