* File: sky130_fd_sc_lp__sdlclkp_lp.spice
* Created: Wed Sep  2 10:37:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdlclkp_lp.pex.spice"
.subckt sky130_fd_sc_lp__sdlclkp_lp  VNB VPB GATE SCE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1011 A_114_101# N_GATE_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1027 N_A_93_376#_M1027_d N_GATE_M1027_g A_114_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1019 A_278_101# N_SCE_M1019_g N_A_93_376#_M1027_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_SCE_M1023_g A_278_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1015 A_436_101# N_A_356_278#_M1015_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_447_376#_M1009_d N_A_356_278#_M1009_g A_436_101# VNB NSHORT L=0.15
+ W=0.42 AD=0.1533 AS=0.0441 PD=1.57 PS=0.63 NRD=22.848 NRS=14.28 M=1 R=2.8
+ SA=75002.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1013 N_A_698_405#_M1013_d N_A_356_278#_M1013_g N_A_93_376#_M1013_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1026 A_812_47# N_A_447_376#_M1026_g N_A_698_405#_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_860_21#_M1024_g A_812_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1008 AS=0.0504 PD=0.9 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1014 A_1016_47# N_A_698_405#_M1014_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1008 PD=0.66 PS=0.9 NRD=18.564 NRS=57.132 M=1 R=2.8 SA=75001.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_860_21#_M1004_d N_A_698_405#_M1004_g A_1016_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75002.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 A_1234_192# N_CLK_M1017_g N_A_356_278#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_CLK_M1012_g A_1234_192# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1016 A_1392_192# N_CLK_M1016_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_1384_416#_M1001_d N_A_860_21#_M1001_g A_1392_192# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 A_1548_48# N_A_1384_416#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1281 PD=0.63 PS=1.45 NRD=14.28 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_GCLK_M1005_d N_A_1384_416#_M1005_g A_1548_48# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 A_200_376# N_GATE_M1018_g N_A_93_376#_M1018_s VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_SCE_M1000_g A_200_376# VPB PHIGHVT L=0.25 W=1
+ AD=0.293175 AS=0.12 PD=1.81 PS=1.24 NRD=46.9057 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1006 N_A_447_376#_M1006_d N_A_356_278#_M1006_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.39545 AS=0.293175 PD=2.94 PS=1.81 NRD=16.7253 NRS=46.9057 M=1
+ R=4 SA=125001 SB=125000 A=0.25 P=2.5 MULT=1
MM1002 N_A_698_405#_M1002_d N_A_447_376#_M1002_g N_A_93_376#_M1002_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1021 A_804_405# N_A_356_278#_M1021_g N_A_698_405#_M1002_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=16.7253 NRS=0 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_A_860_21#_M1008_g A_804_405# VPB PHIGHVT L=0.25 W=1
+ AD=0.1575 AS=0.14 PD=1.315 PS=1.28 NRD=0 NRS=16.7253 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1003 N_A_860_21#_M1003_d N_A_698_405#_M1003_g N_VPWR_M1008_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.1575 PD=2.57 PS=1.315 NRD=0 NRS=6.8753 M=1 R=4
+ SA=125002 SB=125000 A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_CLK_M1007_g N_A_356_278#_M1007_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1025 N_A_1384_416#_M1025_d N_CLK_M1025_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1010 N_VPWR_M1010_d N_A_860_21#_M1010_g N_A_1384_416#_M1025_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.23015 AS=0.14 PD=1.51 PS=1.28 NRD=16.7253 NRS=0 M=1 R=4
+ SA=125001 SB=125001 A=0.25 P=2.5 MULT=1
MM1022 N_GCLK_M1022_d N_A_1384_416#_M1022_g N_VPWR_M1010_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.23015 PD=2.57 PS=1.51 NRD=0 NRS=16.7253 M=1 R=4 SA=125002
+ SB=125000 A=0.25 P=2.5 MULT=1
DX28_noxref VNB VPB NWDIODE A=16.8619 P=22.02
*
.include "sky130_fd_sc_lp__sdlclkp_lp.pxi.spice"
*
.ends
*
*
