* File: sky130_fd_sc_lp__o32ai_lp.pex.spice
* Created: Wed Sep  2 10:27:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32AI_LP%B1 3 7 9 12 13
r28 12 15 30.6934 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.472 $Y=1.68
+ $X2=0.472 $Y2=1.845
r29 12 14 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.472 $Y=1.68
+ $X2=0.472 $Y2=1.515
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.44
+ $Y=1.68 $X2=0.44 $Y2=1.68
r31 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.24 $Y=1.68 $X2=0.44
+ $Y2=1.68
r32 7 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.575 $Y=1.105
+ $X2=0.575 $Y2=1.515
r33 3 15 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.545 $Y=2.595
+ $X2=0.545 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_LP%B2 3 6 8 9 12 14 15
c44 3 0 1.36103e-20 $X=1.035 $Y=2.595
r45 14 15 16.4348 $w=2.28e-07 $l=3.28e-07 $layer=LI1_cond $X=1.68 $Y=0.597
+ $X2=1.68 $Y2=0.925
r46 12 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=0.41
+ $X2=1.095 $Y2=0.575
r47 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=0.41 $X2=1.095 $Y2=0.41
r48 9 14 3.06749 $w=2.9e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=0.41
+ $X2=1.68 $Y2=0.41
r49 9 11 18.6775 $w=2.88e-07 $l=4.7e-07 $layer=LI1_cond $X=1.565 $Y=0.41
+ $X2=1.095 $Y2=0.41
r50 8 21 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.005 $Y=1.105
+ $X2=1.005 $Y2=0.575
r51 6 8 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.005 $Y=1.39
+ $X2=1.005 $Y2=1.105
r52 1 6 55.4603 $w=2.39e-07 $l=2.89612e-07 $layer=POLY_cond $X=1.035 $Y=1.665
+ $X2=1.005 $Y2=1.39
r53 1 3 231.062 $w=2.5e-07 $l=9.3e-07 $layer=POLY_cond $X=1.035 $Y=1.665
+ $X2=1.035 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_LP%A3 3 7 11 12 15 16 17
c41 11 0 1.36103e-20 $X=1.66 $Y=1.77
c42 7 0 1.44789e-19 $X=1.595 $Y=0.975
r43 16 17 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=2.405
+ $X2=1.695 $Y2=2.775
r44 15 16 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=2.035
+ $X2=1.695 $Y2=2.405
r45 14 15 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=1.695 $Y=1.935
+ $X2=1.695 $Y2=2.035
r46 12 23 30.6629 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.632 $Y=1.77
+ $X2=1.632 $Y2=1.935
r47 12 22 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.632 $Y=1.77
+ $X2=1.632 $Y2=1.605
r48 11 14 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=1.77
+ $X2=1.66 $Y2=1.935
r49 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=1.77 $X2=1.66 $Y2=1.77
r50 7 22 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.595 $Y=0.975
+ $X2=1.595 $Y2=1.605
r51 3 23 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.565 $Y=2.595
+ $X2=1.565 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_LP%A2 1 3 7 9 10 11 17
r37 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.77 $X2=2.23 $Y2=1.77
r38 10 11 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.22 $Y=2.405
+ $X2=2.22 $Y2=2.775
r39 9 10 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.22 $Y=2.035 $X2=2.22
+ $Y2=2.405
r40 9 17 8.72564 $w=3.48e-07 $l=2.65e-07 $layer=LI1_cond $X=2.22 $Y=2.035
+ $X2=2.22 $Y2=1.77
r41 5 16 46.4372 $w=3.43e-07 $l=2.68626e-07 $layer=POLY_cond $X=2.355 $Y=1.55
+ $X2=2.247 $Y2=1.77
r42 5 7 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.355 $Y=1.55
+ $X2=2.355 $Y2=0.975
r43 1 16 26.8176 $w=3.43e-07 $l=1.9139e-07 $layer=POLY_cond $X=2.19 $Y=1.935
+ $X2=2.247 $Y2=1.77
r44 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.19 $Y=1.935 $X2=2.19
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_LP%A1 1 3 4 6 8 9 14 15
r31 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.08
+ $Y=1.46 $X2=3.08 $Y2=1.46
r32 11 14 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=2.785 $Y=1.46
+ $X2=3.08 $Y2=1.46
r33 9 15 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.08 $Y=1.665
+ $X2=3.08 $Y2=1.46
r34 7 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.625
+ $X2=2.785 $Y2=1.46
r35 7 8 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.785 $Y=1.625
+ $X2=2.785 $Y2=1.94
r36 4 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.295
+ $X2=2.785 $Y2=1.46
r37 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.785 $Y=1.295
+ $X2=2.785 $Y2=0.975
r38 1 8 29.5102 $w=2.45e-07 $l=1.62019e-07 $layer=POLY_cond $X=2.76 $Y=2.09
+ $X2=2.785 $Y2=1.94
r39 1 3 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.76 $Y=2.09 $X2=2.76
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_LP%VPWR 1 2 7 9 13 15 19 21 34
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 25 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 24 27 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 22 30 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r47 22 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 21 33 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.86 $Y=3.33 $X2=3.11
+ $Y2=3.33
r49 21 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.86 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 19 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 19 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.025 $Y=2.24
+ $X2=3.025 $Y2=2.95
r53 13 33 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.025 $Y=3.245
+ $X2=3.11 $Y2=3.33
r54 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.025 $Y=3.245
+ $X2=3.025 $Y2=2.95
r55 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.24 $X2=0.28
+ $Y2=2.95
r56 7 30 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r57 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.95
r58 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.885
+ $Y=2.095 $X2=3.025 $Y2=2.95
r59 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.885
+ $Y=2.095 $X2=3.025 $Y2=2.24
r60 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.95
r61 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_LP%Y 1 2 8 10 13 14 15 21
c33 10 0 1.44789e-19 $X=0.79 $Y=1.17
r34 19 21 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.235 $Y=2.265
+ $X2=1.235 $Y2=2.28
r35 14 15 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.235 $Y=2.405
+ $X2=1.235 $Y2=2.775
r36 14 21 4.80185 $w=2.98e-07 $l=1.25e-07 $layer=LI1_cond $X=1.235 $Y=2.405
+ $X2=1.235 $Y2=2.28
r37 13 19 1.82479 $w=2.34e-07 $l=3.5e-08 $layer=LI1_cond $X=1.2 $Y=2.092
+ $X2=1.235 $Y2=2.092
r38 10 12 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=1.17
+ $X2=0.79 $Y2=1.335
r39 8 13 17.2051 $w=2.34e-07 $l=4.07014e-07 $layer=LI1_cond $X=0.87 $Y=1.92
+ $X2=1.2 $Y2=2.092
r40 8 12 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=0.87 $Y=1.92
+ $X2=0.87 $Y2=1.335
r41 2 21 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=1.16
+ $Y=2.095 $X2=1.3 $Y2=2.28
r42 1 10 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.895 $X2=0.79 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_LP%A_27_179# 1 2 3 12 14 15 19 20 21 24
r48 22 24 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.57 $Y=1.255
+ $X2=2.57 $Y2=0.975
r49 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.405 $Y=1.34
+ $X2=2.57 $Y2=1.255
r50 20 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.405 $Y=1.34
+ $X2=1.385 $Y2=1.34
r51 17 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.26 $Y=1.255
+ $X2=1.385 $Y2=1.34
r52 17 19 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.26 $Y=1.255
+ $X2=1.26 $Y2=1.04
r53 16 19 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=1.26 $Y=0.905
+ $X2=1.26 $Y2=1.04
r54 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.135 $Y=0.82
+ $X2=1.26 $Y2=0.905
r55 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.135 $Y=0.82
+ $X2=0.445 $Y2=0.82
r56 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.905
+ $X2=0.445 $Y2=0.82
r57 10 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.28 $Y=0.905 $X2=0.28
+ $Y2=1.105
r58 3 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.765 $X2=2.57 $Y2=0.975
r59 2 19 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.895 $X2=1.3 $Y2=1.04
r60 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.895 $X2=0.28 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_LP%VGND 1 2 9 11 13 16 17 18 27 33
r36 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r37 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 27 32 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r40 27 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r41 21 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r42 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r43 18 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r44 18 22 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r45 18 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r46 16 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.68
+ $Y2=0
r47 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.1
+ $Y2=0
r48 15 29 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.64
+ $Y2=0
r49 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.1
+ $Y2=0
r50 11 32 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r51 11 13 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.93
r52 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=0.085
+ $X2=2.1 $Y2=0
r53 7 9 38.0306 $w=2.48e-07 $l=8.25e-07 $layer=LI1_cond $X=2.1 $Y=0.085 $X2=2.1
+ $Y2=0.91
r54 2 13 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=2.86
+ $Y=0.765 $X2=3.08 $Y2=0.93
r55 1 9 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.765 $X2=2.06 $Y2=0.91
.ends

