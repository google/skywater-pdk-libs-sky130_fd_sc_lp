* File: sky130_fd_sc_lp__o221ai_4.pex.spice
* Created: Wed Sep  2 10:19:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221AI_4%C1 3 7 11 15 19 23 27 31 33 34 35 36 37 66
r84 64 66 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.115 $Y=1.51
+ $X2=2.455 $Y2=1.51
r85 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=1.51 $X2=2.115 $Y2=1.51
r86 62 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.025 $Y=1.51
+ $X2=2.115 $Y2=1.51
r87 61 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.935 $Y=1.51
+ $X2=2.025 $Y2=1.51
r88 60 65 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.775 $Y=1.587
+ $X2=2.115 $Y2=1.587
r89 59 61 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.775 $Y=1.51
+ $X2=1.935 $Y2=1.51
r90 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.775
+ $Y=1.51 $X2=1.775 $Y2=1.51
r91 57 59 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.595 $Y=1.51
+ $X2=1.775 $Y2=1.51
r92 55 57 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.435 $Y=1.51
+ $X2=1.595 $Y2=1.51
r93 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.435
+ $Y=1.51 $X2=1.435 $Y2=1.51
r94 53 55 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.425 $Y=1.51
+ $X2=1.435 $Y2=1.51
r95 52 53 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.165 $Y=1.51
+ $X2=1.425 $Y2=1.51
r96 50 52 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.095 $Y=1.51
+ $X2=1.165 $Y2=1.51
r97 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.51 $X2=1.095 $Y2=1.51
r98 48 50 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.915 $Y=1.51
+ $X2=1.095 $Y2=1.51
r99 47 48 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.485 $Y=1.51
+ $X2=0.915 $Y2=1.51
r100 44 47 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.415 $Y=1.51
+ $X2=0.485 $Y2=1.51
r101 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=1.51 $X2=0.415 $Y2=1.51
r102 37 65 1.59569 $w=3.23e-07 $l=4.5e-08 $layer=LI1_cond $X=2.16 $Y=1.587
+ $X2=2.115 $Y2=1.587
r103 36 60 3.36868 $w=3.23e-07 $l=9.5e-08 $layer=LI1_cond $X=1.68 $Y=1.587
+ $X2=1.775 $Y2=1.587
r104 36 56 8.68765 $w=3.23e-07 $l=2.45e-07 $layer=LI1_cond $X=1.68 $Y=1.587
+ $X2=1.435 $Y2=1.587
r105 35 56 8.33305 $w=3.23e-07 $l=2.35e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.435 $Y2=1.587
r106 35 51 3.72328 $w=3.23e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.095 $Y2=1.587
r107 34 51 13.2974 $w=3.23e-07 $l=3.75e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=1.095 $Y2=1.587
r108 34 45 10.8152 $w=3.23e-07 $l=3.05e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=0.415 $Y2=1.587
r109 33 45 6.20546 $w=3.23e-07 $l=1.75e-07 $layer=LI1_cond $X=0.24 $Y=1.587
+ $X2=0.415 $Y2=1.587
r110 29 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.455 $Y=1.675
+ $X2=2.455 $Y2=1.51
r111 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.455 $Y=1.675
+ $X2=2.455 $Y2=2.465
r112 25 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.025 $Y=1.675
+ $X2=2.025 $Y2=1.51
r113 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.025 $Y=1.675
+ $X2=2.025 $Y2=2.465
r114 21 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.345
+ $X2=1.935 $Y2=1.51
r115 21 23 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.935 $Y=1.345
+ $X2=1.935 $Y2=0.745
r116 17 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.675
+ $X2=1.595 $Y2=1.51
r117 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.595 $Y=1.675
+ $X2=1.595 $Y2=2.465
r118 13 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=1.51
r119 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=0.745
r120 9 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.165 $Y=1.675
+ $X2=1.165 $Y2=1.51
r121 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.165 $Y=1.675
+ $X2=1.165 $Y2=2.465
r122 5 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.345
+ $X2=0.915 $Y2=1.51
r123 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.915 $Y=1.345 $X2=0.915
+ $Y2=0.745
r124 1 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.345
+ $X2=0.485 $Y2=1.51
r125 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.485 $Y=1.345 $X2=0.485
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%B1 3 7 11 15 19 23 27 31 33 38 43 44 50 53
+ 54
c126 50 0 4.50227e-20 $X=3.745 $Y=1.51
c127 23 0 4.83235e-20 $X=3.745 $Y=2.465
c128 3 0 1.66203e-19 $X=2.885 $Y=0.655
r129 53 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.46
+ $X2=5.95 $Y2=1.625
r130 53 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.46
+ $X2=5.95 $Y2=1.295
r131 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.46 $X2=5.95 $Y2=1.46
r132 44 61 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=5.98 $Y=1.665
+ $X2=5.98 $Y2=1.7
r133 44 54 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.98 $Y=1.665
+ $X2=5.98 $Y2=1.46
r134 42 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.655 $Y=1.51
+ $X2=3.745 $Y2=1.51
r135 41 43 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.655 $Y=1.592
+ $X2=3.82 $Y2=1.592
r136 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=1.51 $X2=3.655 $Y2=1.51
r137 38 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=1.7
+ $X2=5.98 $Y2=1.7
r138 38 43 130.155 $w=1.68e-07 $l=1.995e-06 $layer=LI1_cond $X=5.815 $Y=1.7
+ $X2=3.82 $Y2=1.7
r139 36 42 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.315 $Y=1.51
+ $X2=3.655 $Y2=1.51
r140 36 46 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.315 $Y=1.51
+ $X2=2.885 $Y2=1.51
r141 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.315
+ $Y=1.51 $X2=3.315 $Y2=1.51
r142 33 41 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=3.628 $Y=1.592
+ $X2=3.655 $Y2=1.592
r143 33 35 9.36921 $w=3.83e-07 $l=3.13e-07 $layer=LI1_cond $X=3.628 $Y=1.592
+ $X2=3.315 $Y2=1.592
r144 31 56 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.895 $Y=2.465
+ $X2=5.895 $Y2=1.625
r145 27 55 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.895 $Y=0.655
+ $X2=5.895 $Y2=1.295
r146 21 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.745 $Y=1.675
+ $X2=3.745 $Y2=1.51
r147 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.745 $Y=1.675
+ $X2=3.745 $Y2=2.465
r148 17 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.745 $Y=1.345
+ $X2=3.745 $Y2=1.51
r149 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.745 $Y=1.345
+ $X2=3.745 $Y2=0.655
r150 13 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=1.675
+ $X2=3.315 $Y2=1.51
r151 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.315 $Y=1.675
+ $X2=3.315 $Y2=2.465
r152 9 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=1.345
+ $X2=3.315 $Y2=1.51
r153 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.315 $Y=1.345
+ $X2=3.315 $Y2=0.655
r154 5 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.675
+ $X2=2.885 $Y2=1.51
r155 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.885 $Y=1.675
+ $X2=2.885 $Y2=2.465
r156 1 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.345
+ $X2=2.885 $Y2=1.51
r157 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.885 $Y=1.345
+ $X2=2.885 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 45
c84 31 0 4.50227e-20 $X=5.52 $Y=1.295
c85 1 0 1.20142e-19 $X=4.175 $Y=1.185
r86 43 45 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=5.41 $Y=1.35
+ $X2=5.465 $Y2=1.35
r87 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.41
+ $Y=1.35 $X2=5.41 $Y2=1.35
r88 41 43 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=5.035 $Y=1.35
+ $X2=5.41 $Y2=1.35
r89 40 41 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.605 $Y=1.35
+ $X2=5.035 $Y2=1.35
r90 38 40 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.39 $Y=1.35
+ $X2=4.605 $Y2=1.35
r91 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.39
+ $Y=1.35 $X2=4.39 $Y2=1.35
r92 35 38 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.175 $Y=1.35
+ $X2=4.39 $Y2=1.35
r93 31 44 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=5.52 $Y=1.32
+ $X2=5.41 $Y2=1.32
r94 30 44 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=5.04 $Y=1.32
+ $X2=5.41 $Y2=1.32
r95 29 30 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.32
+ $X2=5.04 $Y2=1.32
r96 29 39 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=4.56 $Y=1.32
+ $X2=4.39 $Y2=1.32
r97 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.465 $Y=1.515
+ $X2=5.465 $Y2=1.35
r98 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.465 $Y=1.515
+ $X2=5.465 $Y2=2.465
r99 22 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.465 $Y=1.185
+ $X2=5.465 $Y2=1.35
r100 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.465 $Y=1.185
+ $X2=5.465 $Y2=0.655
r101 18 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.035 $Y=1.515
+ $X2=5.035 $Y2=1.35
r102 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.035 $Y=1.515
+ $X2=5.035 $Y2=2.465
r103 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.035 $Y=1.185
+ $X2=5.035 $Y2=1.35
r104 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.035 $Y=1.185
+ $X2=5.035 $Y2=0.655
r105 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.605 $Y=1.515
+ $X2=4.605 $Y2=1.35
r106 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.605 $Y=1.515
+ $X2=4.605 $Y2=2.465
r107 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.605 $Y=1.185
+ $X2=4.605 $Y2=1.35
r108 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.605 $Y=1.185
+ $X2=4.605 $Y2=0.655
r109 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.175 $Y=1.515
+ $X2=4.175 $Y2=1.35
r110 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.175 $Y=1.515
+ $X2=4.175 $Y2=2.465
r111 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.175 $Y=1.185
+ $X2=4.175 $Y2=1.35
r112 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.175 $Y=1.185
+ $X2=4.175 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%A1 3 6 8 10 13 15 17 20 22 24 27 31 35 38
+ 39 40 41 42 47 60
c111 60 0 6.98577e-20 $X=9.77 $Y=1.35
c112 31 0 1.01656e-19 $X=6.53 $Y=1.16
r113 58 60 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=9.555 $Y=1.35
+ $X2=9.77 $Y2=1.35
r114 57 58 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=9.52 $Y=1.35
+ $X2=9.555 $Y2=1.35
r115 56 57 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=9.125 $Y=1.35
+ $X2=9.52 $Y2=1.35
r116 55 56 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=9.09 $Y=1.35
+ $X2=9.125 $Y2=1.35
r117 53 55 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.75 $Y=1.35
+ $X2=9.09 $Y2=1.35
r118 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.75
+ $Y=1.35 $X2=8.75 $Y2=1.35
r119 51 53 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=8.695 $Y=1.35
+ $X2=8.75 $Y2=1.35
r120 49 51 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=8.66 $Y=1.35
+ $X2=8.695 $Y2=1.35
r121 42 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.77
+ $Y=1.35 $X2=9.77 $Y2=1.35
r122 41 42 15.242 $w=3.08e-07 $l=4.1e-07 $layer=LI1_cond $X=9.36 $Y=1.365
+ $X2=9.77 $Y2=1.365
r123 40 41 17.8443 $w=3.08e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=9.36 $Y2=1.365
r124 40 54 4.83283 $w=3.08e-07 $l=1.3e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=8.75 $Y2=1.365
r125 39 54 5.94809 $w=3.08e-07 $l=1.6e-07 $layer=LI1_cond $X=8.59 $Y=1.365
+ $X2=8.75 $Y2=1.365
r126 38 39 9.95431 $w=3.08e-07 $l=2.05e-07 $layer=LI1_cond $X=8.385 $Y=1.297
+ $X2=8.59 $Y2=1.297
r127 35 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.49 $Y=1.35
+ $X2=6.49 $Y2=1.515
r128 35 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.49 $Y=1.35
+ $X2=6.49 $Y2=1.185
r129 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.49
+ $Y=1.35 $X2=6.49 $Y2=1.35
r130 31 34 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=6.53 $Y=1.16
+ $X2=6.53 $Y2=1.35
r131 30 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.655 $Y=1.16
+ $X2=6.53 $Y2=1.16
r132 30 38 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=6.655 $Y=1.16
+ $X2=8.385 $Y2=1.16
r133 25 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.555 $Y=1.515
+ $X2=9.555 $Y2=1.35
r134 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.555 $Y=1.515
+ $X2=9.555 $Y2=2.465
r135 22 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.52 $Y=1.185
+ $X2=9.52 $Y2=1.35
r136 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.52 $Y=1.185
+ $X2=9.52 $Y2=0.655
r137 18 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.125 $Y=1.515
+ $X2=9.125 $Y2=1.35
r138 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.125 $Y=1.515
+ $X2=9.125 $Y2=2.465
r139 15 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.09 $Y=1.185
+ $X2=9.09 $Y2=1.35
r140 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.09 $Y=1.185
+ $X2=9.09 $Y2=0.655
r141 11 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.695 $Y=1.515
+ $X2=8.695 $Y2=1.35
r142 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.695 $Y=1.515
+ $X2=8.695 $Y2=2.465
r143 8 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.66 $Y=1.185
+ $X2=8.66 $Y2=1.35
r144 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.66 $Y=1.185
+ $X2=8.66 $Y2=0.655
r145 6 48 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.51 $Y=2.465
+ $X2=6.51 $Y2=1.515
r146 3 47 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.51 $Y=0.655
+ $X2=6.51 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%A2 3 7 11 15 19 23 27 31 33 34 35 50 51
c82 51 0 1.01656e-19 $X=8.23 $Y=1.51
c83 50 0 6.98577e-20 $X=8.05 $Y=1.51
c84 23 0 4.10644e-20 $X=7.8 $Y=2.465
r85 49 51 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=8.05 $Y=1.51 $X2=8.23
+ $Y2=1.51
r86 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.05
+ $Y=1.51 $X2=8.05 $Y2=1.51
r87 47 49 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=7.8 $Y=1.51 $X2=8.05
+ $Y2=1.51
r88 45 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.71 $Y=1.51 $X2=7.8
+ $Y2=1.51
r89 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.71
+ $Y=1.51 $X2=7.71 $Y2=1.51
r90 42 45 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.37 $Y=1.51
+ $X2=7.71 $Y2=1.51
r91 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.37
+ $Y=1.51 $X2=7.37 $Y2=1.51
r92 39 42 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.94 $Y=1.51
+ $X2=7.37 $Y2=1.51
r93 35 50 4.60977 $w=3.23e-07 $l=1.3e-07 $layer=LI1_cond $X=7.92 $Y=1.587
+ $X2=8.05 $Y2=1.587
r94 35 46 7.44655 $w=3.23e-07 $l=2.1e-07 $layer=LI1_cond $X=7.92 $Y=1.587
+ $X2=7.71 $Y2=1.587
r95 34 46 9.57414 $w=3.23e-07 $l=2.7e-07 $layer=LI1_cond $X=7.44 $Y=1.587
+ $X2=7.71 $Y2=1.587
r96 34 43 2.48218 $w=3.23e-07 $l=7e-08 $layer=LI1_cond $X=7.44 $Y=1.587 $X2=7.37
+ $Y2=1.587
r97 33 43 14.5385 $w=3.23e-07 $l=4.1e-07 $layer=LI1_cond $X=6.96 $Y=1.587
+ $X2=7.37 $Y2=1.587
r98 29 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=1.675
+ $X2=8.23 $Y2=1.51
r99 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.23 $Y=1.675
+ $X2=8.23 $Y2=2.465
r100 25 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=1.345
+ $X2=8.23 $Y2=1.51
r101 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.23 $Y=1.345
+ $X2=8.23 $Y2=0.655
r102 21 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.8 $Y=1.675
+ $X2=7.8 $Y2=1.51
r103 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.8 $Y=1.675
+ $X2=7.8 $Y2=2.465
r104 17 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.8 $Y=1.345
+ $X2=7.8 $Y2=1.51
r105 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.8 $Y=1.345
+ $X2=7.8 $Y2=0.655
r106 13 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.37 $Y=1.675
+ $X2=7.37 $Y2=1.51
r107 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.37 $Y=1.675
+ $X2=7.37 $Y2=2.465
r108 9 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.37 $Y=1.345
+ $X2=7.37 $Y2=1.51
r109 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.37 $Y=1.345
+ $X2=7.37 $Y2=0.655
r110 5 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.94 $Y=1.675
+ $X2=6.94 $Y2=1.51
r111 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.94 $Y=1.675
+ $X2=6.94 $Y2=2.465
r112 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.94 $Y=1.345
+ $X2=6.94 $Y2=1.51
r113 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.94 $Y=1.345
+ $X2=6.94 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 48 52
+ 54 58 59 61 62 63 69 74 86 93 99 102 105 108 112
r144 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r145 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r146 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r147 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r148 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r149 97 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r150 97 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r151 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r152 94 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.075 $Y=3.33
+ $X2=8.91 $Y2=3.33
r153 94 96 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.075 $Y=3.33
+ $X2=9.36 $Y2=3.33
r154 93 111 4.352 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=9.64 $Y=3.33 $X2=9.86
+ $Y2=3.33
r155 93 96 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=9.64 $Y=3.33
+ $X2=9.36 $Y2=3.33
r156 92 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r157 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r158 89 92 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r159 88 91 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r160 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r161 86 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.745 $Y=3.33
+ $X2=8.91 $Y2=3.33
r162 86 91 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.745 $Y=3.33
+ $X2=8.4 $Y2=3.33
r163 85 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r164 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r165 82 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r166 81 84 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r167 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r168 79 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=3.33
+ $X2=3.53 $Y2=3.33
r169 79 81 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.695 $Y=3.33
+ $X2=4.08 $Y2=3.33
r170 78 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r171 78 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r172 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r173 75 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.67 $Y2=3.33
r174 75 77 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.12 $Y2=3.33
r175 74 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.53 $Y2=3.33
r176 74 77 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.12 $Y2=3.33
r177 73 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r178 73 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r179 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r180 70 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=1.81 $Y2=3.33
r181 70 72 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=2.16 $Y2=3.33
r182 69 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.67 $Y2=3.33
r183 69 72 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r184 67 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r185 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r186 63 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r187 63 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r188 61 84 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.05 $Y=3.33 $X2=6
+ $Y2=3.33
r189 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.05 $Y=3.33
+ $X2=6.215 $Y2=3.33
r190 60 88 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.38 $Y=3.33 $X2=6.48
+ $Y2=3.33
r191 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.38 $Y=3.33
+ $X2=6.215 $Y2=3.33
r192 58 66 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.72 $Y2=3.33
r193 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.95 $Y2=3.33
r194 54 57 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=9.787 $Y=1.98
+ $X2=9.787 $Y2=2.95
r195 52 111 3.12553 $w=2.95e-07 $l=1.15888e-07 $layer=LI1_cond $X=9.787 $Y=3.245
+ $X2=9.86 $Y2=3.33
r196 52 57 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=9.787 $Y=3.245
+ $X2=9.787 $Y2=2.95
r197 48 51 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=8.91 $Y=2.115
+ $X2=8.91 $Y2=2.95
r198 46 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=3.245
+ $X2=8.91 $Y2=3.33
r199 46 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.91 $Y=3.245
+ $X2=8.91 $Y2=2.95
r200 42 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.215 $Y=3.245
+ $X2=6.215 $Y2=3.33
r201 42 44 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=6.215 $Y=3.245
+ $X2=6.215 $Y2=2.435
r202 38 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=3.245
+ $X2=3.53 $Y2=3.33
r203 38 40 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.53 $Y=3.245
+ $X2=3.53 $Y2=2.75
r204 34 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=3.33
r205 34 36 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=2.42
r206 30 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=3.245
+ $X2=1.81 $Y2=3.33
r207 30 32 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=1.81 $Y=3.245
+ $X2=1.81 $Y2=2.38
r208 29 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.95 $Y2=3.33
r209 28 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=1.81 $Y2=3.33
r210 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=1.115 $Y2=3.33
r211 24 27 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.95 $Y=2.005
+ $X2=0.95 $Y2=2.95
r212 22 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.95 $Y=3.245
+ $X2=0.95 $Y2=3.33
r213 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.95 $Y=3.245
+ $X2=0.95 $Y2=2.95
r214 7 57 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.63
+ $Y=1.835 $X2=9.77 $Y2=2.95
r215 7 54 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.63
+ $Y=1.835 $X2=9.77 $Y2=1.98
r216 6 51 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.835 $X2=8.91 $Y2=2.95
r217 6 48 400 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.835 $X2=8.91 $Y2=2.115
r218 5 44 300 $w=1.7e-07 $l=7.12039e-07 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=1.835 $X2=6.215 $Y2=2.435
r219 4 40 600 $w=1.7e-07 $l=9.8251e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.835 $X2=3.53 $Y2=2.75
r220 3 36 300 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_PDIFF $count=2 $X=2.53
+ $Y=1.835 $X2=2.67 $Y2=2.42
r221 2 32 300 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=2 $X=1.67
+ $Y=1.835 $X2=1.81 $Y2=2.38
r222 1 27 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.825
+ $Y=1.835 $X2=0.95 $Y2=2.95
r223 1 24 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.825
+ $Y=1.835 $X2=0.95 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%Y 1 2 3 4 5 6 7 8 27 29 30 31 33 39 41 45
+ 48 49 53 59 65 68 70 72 75 77 78 79 91 92
c141 92 0 4.10644e-20 $X=7.32 $Y=2.042
c142 72 0 4.83235e-20 $X=4.39 $Y=2.04
r143 91 92 9.98442 $w=1.83e-07 $l=1.65e-07 $layer=LI1_cond $X=7.155 $Y=2.042
+ $X2=7.32 $Y2=2.042
r144 79 91 11.6904 $w=1.83e-07 $l=1.95e-07 $layer=LI1_cond $X=6.96 $Y=2.042
+ $X2=7.155 $Y2=2.042
r145 78 79 28.7764 $w=1.83e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=2.042
+ $X2=6.96 $Y2=2.042
r146 73 78 34.1196 $w=3.43e-07 $l=9.8e-07 $layer=LI1_cond $X=5.415 $Y=2.045
+ $X2=6.395 $Y2=2.045
r147 73 75 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.415 $Y=2.045
+ $X2=5.25 $Y2=2.045
r148 67 68 5.49576 $w=2.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.24 $Y=2.022
+ $X2=2.145 $Y2=2.022
r149 59 77 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.85 $Y=2.035
+ $X2=8.015 $Y2=2.035
r150 59 92 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.85 $Y=2.035
+ $X2=7.32 $Y2=2.035
r151 54 72 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=4.555 $Y=2.045
+ $X2=4.39 $Y2=2.045
r152 53 75 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.085 $Y=2.045
+ $X2=5.25 $Y2=2.045
r153 53 54 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=5.085 $Y=2.045
+ $X2=4.555 $Y2=2.045
r154 49 72 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.225 $Y=2.04
+ $X2=4.39 $Y2=2.045
r155 49 70 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=4.225 $Y=2.04
+ $X2=2.64 $Y2=2.04
r156 48 70 5.22525 $w=2.03e-07 $l=9e-08 $layer=LI1_cond $X=2.55 $Y=2.022
+ $X2=2.64 $Y2=2.022
r157 48 67 16.7716 $w=2.03e-07 $l=3.1e-07 $layer=LI1_cond $X=2.55 $Y=2.022
+ $X2=2.24 $Y2=2.022
r158 47 48 40.9747 $w=1.78e-07 $l=6.65e-07 $layer=LI1_cond $X=2.55 $Y=1.255
+ $X2=2.55 $Y2=1.92
r159 43 67 1.17563 $w=1.9e-07 $l=1.03e-07 $layer=LI1_cond $X=2.24 $Y=2.125
+ $X2=2.24 $Y2=2.022
r160 43 45 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=2.24 $Y=2.125
+ $X2=2.24 $Y2=2.48
r161 42 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=1.17
+ $X2=1.7 $Y2=1.17
r162 41 47 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.46 $Y=1.17
+ $X2=2.55 $Y2=1.255
r163 41 42 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.46 $Y=1.17
+ $X2=1.865 $Y2=1.17
r164 37 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=1.085 $X2=1.7
+ $Y2=1.17
r165 37 39 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.7 $Y=1.085
+ $X2=1.7 $Y2=0.7
r166 36 64 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.465 $Y=2.005
+ $X2=1.375 $Y2=2.005
r167 36 68 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.465 $Y=2.005
+ $X2=2.145 $Y2=2.005
r168 31 64 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=2.09
+ $X2=1.375 $Y2=2.005
r169 31 33 50.5253 $w=1.78e-07 $l=8.2e-07 $layer=LI1_cond $X=1.375 $Y=2.09
+ $X2=1.375 $Y2=2.91
r170 29 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=1.17
+ $X2=1.7 $Y2=1.17
r171 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=1.17
+ $X2=0.865 $Y2=1.17
r172 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.7 $Y=1.085
+ $X2=0.865 $Y2=1.17
r173 25 27 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.7 $Y=1.085
+ $X2=0.7 $Y2=0.7
r174 8 77 300 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=2 $X=7.875
+ $Y=1.835 $X2=8.015 $Y2=2.035
r175 7 91 300 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=2 $X=7.015
+ $Y=1.835 $X2=7.155 $Y2=2.035
r176 6 75 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=5.11
+ $Y=1.835 $X2=5.25 $Y2=2.04
r177 5 72 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=4.25
+ $Y=1.835 $X2=4.39 $Y2=2.04
r178 4 67 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.835 $X2=2.24 $Y2=2.005
r179 4 45 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=2.1
+ $Y=1.835 $X2=2.24 $Y2=2.48
r180 3 64 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.24
+ $Y=1.835 $X2=1.38 $Y2=2.085
r181 3 33 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.24
+ $Y=1.835 $X2=1.38 $Y2=2.91
r182 2 39 91 $w=1.7e-07 $l=4.64354e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.325 $X2=1.7 $Y2=0.7
r183 1 27 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.325 $X2=0.7 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%A_592_367# 1 2 3 4 15 17 19 20 23 25 29 32
+ 35
r39 27 29 19.2813 $w=2.58e-07 $l=4.35e-07 $layer=LI1_cond $X=5.715 $Y=2.905
+ $X2=5.715 $Y2=2.47
r40 26 35 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.915 $Y=2.99
+ $X2=4.82 $Y2=2.99
r41 25 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.585 $Y=2.99
+ $X2=5.715 $Y2=2.905
r42 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.585 $Y=2.99
+ $X2=4.915 $Y2=2.99
r43 21 35 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.82 $Y=2.905
+ $X2=4.82 $Y2=2.99
r44 21 23 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=4.82 $Y=2.905
+ $X2=4.82 $Y2=2.48
r45 19 35 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.725 $Y=2.99
+ $X2=4.82 $Y2=2.99
r46 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.725 $Y=2.99
+ $X2=4.055 $Y2=2.99
r47 18 20 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.96 $Y=2.905
+ $X2=4.055 $Y2=2.99
r48 17 34 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=2.465
+ $X2=3.96 $Y2=2.38
r49 17 18 25.6842 $w=1.88e-07 $l=4.4e-07 $layer=LI1_cond $X=3.96 $Y=2.465
+ $X2=3.96 $Y2=2.905
r50 16 32 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.195 $Y=2.38 $X2=3.1
+ $Y2=2.38
r51 15 34 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.865 $Y=2.38
+ $X2=3.96 $Y2=2.38
r52 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.865 $Y=2.38
+ $X2=3.195 $Y2=2.38
r53 4 29 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=5.54
+ $Y=1.835 $X2=5.68 $Y2=2.47
r54 3 23 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=4.68
+ $Y=1.835 $X2=4.82 $Y2=2.48
r55 2 34 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=3.82
+ $Y=1.835 $X2=3.96 $Y2=2.46
r56 1 32 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%A_1317_367# 1 2 3 4 15 17 18 21 23 26 28 29
+ 30 33 37
r46 33 35 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=9.357 $Y=1.98
+ $X2=9.357 $Y2=2.91
r47 31 33 6.14636 $w=2.23e-07 $l=1.2e-07 $layer=LI1_cond $X=9.357 $Y=1.86
+ $X2=9.357 $Y2=1.98
r48 29 31 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=9.245 $Y=1.775
+ $X2=9.357 $Y2=1.86
r49 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.245 $Y=1.775
+ $X2=8.575 $Y2=1.775
r50 26 39 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.48 $Y=2.905
+ $X2=8.48 $Y2=2.99
r51 26 28 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=8.48 $Y=2.905
+ $X2=8.48 $Y2=1.98
r52 25 30 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.48 $Y=1.86
+ $X2=8.575 $Y2=1.775
r53 25 28 7.00478 $w=1.88e-07 $l=1.2e-07 $layer=LI1_cond $X=8.48 $Y=1.86
+ $X2=8.48 $Y2=1.98
r54 24 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.68 $Y=2.99
+ $X2=7.585 $Y2=2.99
r55 23 39 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.385 $Y=2.99
+ $X2=8.48 $Y2=2.99
r56 23 24 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=8.385 $Y=2.99
+ $X2=7.68 $Y2=2.99
r57 19 37 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.585 $Y=2.905
+ $X2=7.585 $Y2=2.99
r58 19 21 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=7.585 $Y=2.905
+ $X2=7.585 $Y2=2.455
r59 17 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.49 $Y=2.99
+ $X2=7.585 $Y2=2.99
r60 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.49 $Y=2.99
+ $X2=6.82 $Y2=2.99
r61 13 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.69 $Y=2.905
+ $X2=6.82 $Y2=2.99
r62 13 15 19.2813 $w=2.58e-07 $l=4.35e-07 $layer=LI1_cond $X=6.69 $Y=2.905
+ $X2=6.69 $Y2=2.47
r63 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.2
+ $Y=1.835 $X2=9.34 $Y2=2.91
r64 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.2
+ $Y=1.835 $X2=9.34 $Y2=1.98
r65 3 39 400 $w=1.7e-07 $l=1.1592e-06 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.835 $X2=8.48 $Y2=2.91
r66 3 28 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.835 $X2=8.48 $Y2=1.98
r67 2 21 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=7.445
+ $Y=1.835 $X2=7.585 $Y2=2.455
r68 1 15 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=6.585
+ $Y=1.835 $X2=6.725 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%A_29_65# 1 2 3 4 5 6 7 24 26 27 30 32 35 36
+ 38 44 55 58 59
c93 38 0 1.66203e-19 $X=3.865 $Y=1.117
r94 58 59 6.36939 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=0.845
+ $X2=5.515 $Y2=0.845
r95 55 56 11.7142 $w=2.26e-07 $l=2.17e-07 $layer=LI1_cond $X=3.99 $Y=0.9
+ $X2=3.99 $Y2=1.117
r96 54 55 6.47788 $w=2.26e-07 $l=1.2e-07 $layer=LI1_cond $X=3.99 $Y=0.78
+ $X2=3.99 $Y2=0.9
r97 50 51 8.89028 $w=3.83e-07 $l=2.97e-07 $layer=LI1_cond $X=3.002 $Y=0.82
+ $X2=3.002 $Y2=1.117
r98 43 59 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=4.82 $Y=0.9
+ $X2=5.515 $Y2=0.9
r99 41 55 0.0912679 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=4.115 $Y=0.9
+ $X2=3.99 $Y2=0.9
r100 41 43 32.4989 $w=2.48e-07 $l=7.05e-07 $layer=LI1_cond $X=4.115 $Y=0.9
+ $X2=4.82 $Y2=0.9
r101 39 51 3.89577 $w=2.25e-07 $l=1.93e-07 $layer=LI1_cond $X=3.195 $Y=1.117
+ $X2=3.002 $Y2=1.117
r102 38 56 0.770517 $w=2.25e-07 $l=1.25e-07 $layer=LI1_cond $X=3.865 $Y=1.117
+ $X2=3.99 $Y2=1.117
r103 38 39 34.3172 $w=2.23e-07 $l=6.7e-07 $layer=LI1_cond $X=3.865 $Y=1.117
+ $X2=3.195 $Y2=1.117
r104 37 46 3.54079 $w=2.6e-07 $l=1.4e-07 $layer=LI1_cond $X=2.315 $Y=0.785
+ $X2=2.175 $Y2=0.785
r105 36 50 1.04768 $w=3.83e-07 $l=3.5e-08 $layer=LI1_cond $X=3.002 $Y=0.785
+ $X2=3.002 $Y2=0.82
r106 36 37 21.9407 $w=2.58e-07 $l=4.95e-07 $layer=LI1_cond $X=2.81 $Y=0.785
+ $X2=2.315 $Y2=0.785
r107 35 46 3.28787 $w=2.8e-07 $l=1.3e-07 $layer=LI1_cond $X=2.175 $Y=0.655
+ $X2=2.175 $Y2=0.785
r108 34 35 9.4665 $w=2.78e-07 $l=2.3e-07 $layer=LI1_cond $X=2.175 $Y=0.425
+ $X2=2.175 $Y2=0.655
r109 33 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0.34
+ $X2=1.2 $Y2=0.34
r110 32 34 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=2.175 $Y2=0.425
r111 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=1.365 $Y2=0.34
r112 28 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.425 $X2=1.2
+ $Y2=0.34
r113 28 30 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.2 $Y=0.425
+ $X2=1.2 $Y2=0.45
r114 26 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0.34
+ $X2=1.2 $Y2=0.34
r115 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.035 $Y=0.34
+ $X2=0.365 $Y2=0.34
r116 22 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.235 $Y=0.425
+ $X2=0.365 $Y2=0.34
r117 22 24 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=0.235 $Y=0.425
+ $X2=0.235 $Y2=0.47
r118 7 58 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.54
+ $Y=0.235 $X2=5.68 $Y2=0.83
r119 6 43 182 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_NDIFF $count=1 $X=4.68
+ $Y=0.235 $X2=4.82 $Y2=0.89
r120 5 54 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=3.82
+ $Y=0.235 $X2=3.96 $Y2=0.78
r121 4 50 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.82
r122 3 46 182 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_NDIFF $count=1 $X=2.01
+ $Y=0.325 $X2=2.15 $Y2=0.75
r123 2 30 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=0.99
+ $Y=0.325 $X2=1.2 $Y2=0.45
r124 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.325 $X2=0.27 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%A_509_47# 1 2 3 4 5 6 7 8 9 28 36 37 38 40
+ 41 42 46 48 52 54 58 60 64 67 70 79 81 82
c106 67 0 1.20142e-19 $X=3.53 $Y=0.38
r107 85 86 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=8.865 $Y=0.875
+ $X2=8.865 $Y2=0.955
r108 82 85 2.90476 $w=2.08e-07 $l=5.5e-08 $layer=LI1_cond $X=8.865 $Y=0.82
+ $X2=8.865 $Y2=0.875
r109 82 83 4.61288 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=8.865 $Y=0.82
+ $X2=8.865 $Y2=0.735
r110 72 73 5.84923 $w=3.48e-07 $l=1.05e-07 $layer=LI1_cond $X=5.25 $Y=0.43
+ $X2=5.355 $Y2=0.43
r111 69 70 5.84923 $w=3.48e-07 $l=1.05e-07 $layer=LI1_cond $X=4.39 $Y=0.43
+ $X2=4.285 $Y2=0.43
r112 62 64 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=9.77 $Y=0.87
+ $X2=9.77 $Y2=0.42
r113 61 86 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.97 $Y=0.955
+ $X2=8.865 $Y2=0.955
r114 60 62 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.64 $Y=0.955
+ $X2=9.77 $Y2=0.87
r115 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.64 $Y=0.955
+ $X2=8.97 $Y2=0.955
r116 58 83 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=8.875 $Y=0.42
+ $X2=8.875 $Y2=0.735
r117 55 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.11 $Y=0.82
+ $X2=8.015 $Y2=0.82
r118 54 82 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.76 $Y=0.82
+ $X2=8.865 $Y2=0.82
r119 54 55 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.76 $Y=0.82
+ $X2=8.11 $Y2=0.82
r120 50 81 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=0.735
+ $X2=8.015 $Y2=0.82
r121 50 52 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=8.015 $Y=0.735
+ $X2=8.015 $Y2=0.42
r122 49 79 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.25 $Y=0.82
+ $X2=7.155 $Y2=0.82
r123 48 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.92 $Y=0.82
+ $X2=8.015 $Y2=0.82
r124 48 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.92 $Y=0.82
+ $X2=7.25 $Y2=0.82
r125 44 79 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.155 $Y=0.735
+ $X2=7.155 $Y2=0.82
r126 44 46 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=7.155 $Y=0.735
+ $X2=7.155 $Y2=0.42
r127 43 77 4.95428 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=6.39 $Y=0.82
+ $X2=6.225 $Y2=0.84
r128 42 79 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.06 $Y=0.82
+ $X2=7.155 $Y2=0.82
r129 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.06 $Y=0.82
+ $X2=6.39 $Y2=0.82
r130 41 77 2.81189 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=6.225 $Y=0.735
+ $X2=6.225 $Y2=0.84
r131 40 75 2.73294 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=6.225 $Y=0.445
+ $X2=6.225 $Y2=0.35
r132 40 41 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=6.225 $Y=0.445
+ $X2=6.225 $Y2=0.735
r133 38 75 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=6.06 $Y=0.35
+ $X2=6.225 $Y2=0.35
r134 38 73 41.1531 $w=1.88e-07 $l=7.05e-07 $layer=LI1_cond $X=6.06 $Y=0.35
+ $X2=5.355 $Y2=0.35
r135 37 69 8.0671 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=4.635 $Y=0.43
+ $X2=4.39 $Y2=0.43
r136 36 72 2.30489 $w=3.48e-07 $l=7e-08 $layer=LI1_cond $X=5.18 $Y=0.43 $X2=5.25
+ $Y2=0.43
r137 36 37 17.9452 $w=3.48e-07 $l=5.45e-07 $layer=LI1_cond $X=5.18 $Y=0.43
+ $X2=4.635 $Y2=0.43
r138 35 67 7.38875 $w=2.1e-07 $l=1.74714e-07 $layer=LI1_cond $X=3.695 $Y=0.35
+ $X2=3.53 $Y2=0.37
r139 35 70 34.4402 $w=1.88e-07 $l=5.9e-07 $layer=LI1_cond $X=3.695 $Y=0.35
+ $X2=4.285 $Y2=0.35
r140 28 67 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0.37
+ $X2=3.53 $Y2=0.37
r141 28 30 34.8238 $w=2.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.365 $Y=0.37
+ $X2=2.67 $Y2=0.37
r142 9 64 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.595
+ $Y=0.235 $X2=9.735 $Y2=0.42
r143 8 85 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.235 $X2=8.875 $Y2=0.875
r144 8 58 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.235 $X2=8.875 $Y2=0.42
r145 7 81 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=7.875
+ $Y=0.235 $X2=8.015 $Y2=0.82
r146 7 52 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=7.875
+ $Y=0.235 $X2=8.015 $Y2=0.42
r147 6 79 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=7.015
+ $Y=0.235 $X2=7.155 $Y2=0.82
r148 6 46 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=7.015
+ $Y=0.235 $X2=7.155 $Y2=0.42
r149 5 77 182 $w=1.7e-07 $l=7.00999e-07 $layer=licon1_NDIFF $count=1 $X=5.97
+ $Y=0.235 $X2=6.225 $Y2=0.82
r150 5 75 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=5.97
+ $Y=0.235 $X2=6.225 $Y2=0.38
r151 4 72 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.11
+ $Y=0.235 $X2=5.25 $Y2=0.44
r152 3 69 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=4.25
+ $Y=0.235 $X2=4.39 $Y2=0.44
r153 2 67 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.39
+ $Y=0.235 $X2=3.53 $Y2=0.38
r154 1 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.235 $X2=2.67 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_4%VGND 1 2 3 4 15 17 21 25 29 31 32 33 42 47
+ 54 55 58 61 64
r127 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r128 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r129 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r130 55 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r131 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r132 52 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.47 $Y=0 $X2=9.305
+ $Y2=0
r133 52 54 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.47 $Y=0 $X2=9.84
+ $Y2=0
r134 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r135 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r136 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r137 48 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.61 $Y=0 $X2=8.445
+ $Y2=0
r138 48 50 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.61 $Y=0 $X2=8.88
+ $Y2=0
r139 47 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.14 $Y=0 $X2=9.305
+ $Y2=0
r140 47 50 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.14 $Y=0 $X2=8.88
+ $Y2=0
r141 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r142 46 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r143 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r144 43 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.75 $Y=0 $X2=7.585
+ $Y2=0
r145 43 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.75 $Y=0 $X2=7.92
+ $Y2=0
r146 42 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=0 $X2=8.445
+ $Y2=0
r147 42 45 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.28 $Y=0 $X2=7.92
+ $Y2=0
r148 41 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r149 40 41 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r150 36 40 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=6.48
+ $Y2=0
r151 36 37 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r152 33 41 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r153 33 37 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=0.24
+ $Y2=0
r154 31 40 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.48
+ $Y2=0
r155 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.725
+ $Y2=0
r156 27 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.305 $Y=0.085
+ $X2=9.305 $Y2=0
r157 27 29 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=9.305 $Y=0.085
+ $X2=9.305 $Y2=0.555
r158 23 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.445 $Y=0.085
+ $X2=8.445 $Y2=0
r159 23 25 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=8.445 $Y=0.085
+ $X2=8.445 $Y2=0.44
r160 19 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.585 $Y=0.085
+ $X2=7.585 $Y2=0
r161 19 21 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=7.585 $Y=0.085
+ $X2=7.585 $Y2=0.44
r162 18 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.89 $Y=0 $X2=6.725
+ $Y2=0
r163 17 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.42 $Y=0 $X2=7.585
+ $Y2=0
r164 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.42 $Y=0 $X2=6.89
+ $Y2=0
r165 13 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.725 $Y=0.085
+ $X2=6.725 $Y2=0
r166 13 15 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=6.725 $Y=0.085
+ $X2=6.725 $Y2=0.44
r167 4 29 182 $w=1.7e-07 $l=3.83667e-07 $layer=licon1_NDIFF $count=1 $X=9.165
+ $Y=0.235 $X2=9.305 $Y2=0.555
r168 3 25 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=8.305
+ $Y=0.235 $X2=8.445 $Y2=0.44
r169 2 21 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=7.445
+ $Y=0.235 $X2=7.585 $Y2=0.44
r170 1 15 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=6.585
+ $Y=0.235 $X2=6.725 $Y2=0.44
.ends

