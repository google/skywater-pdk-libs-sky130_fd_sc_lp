* File: sky130_fd_sc_lp__sdfrtp_4.pex.spice
* Created: Wed Sep  2 10:34:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%A_27_74# 1 2 9 12 16 19 22 23 25 26 29 31
+ 33 34 36 37 42
c82 36 0 1.94921e-19 $X=2.77 $Y=1.935
c83 16 0 9.46857e-21 $X=0.26 $Y=0.58
c84 12 0 8.81054e-20 $X=2.75 $Y=2.635
r85 37 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.935
+ $X2=2.77 $Y2=2.1
r86 36 39 4.24099 $w=2.48e-07 $l=9.2e-08 $layer=LI1_cond $X=2.73 $Y=1.935
+ $X2=2.73 $Y2=2.027
r87 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.935 $X2=2.77 $Y2=1.935
r88 32 34 5.63431 $w=2.7e-07 $l=1.83712e-07 $layer=LI1_cond $X=1.45 $Y=2.027
+ $X2=1.3 $Y2=2.102
r89 31 39 2.2192 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=2.605 $Y=2.027
+ $X2=2.73 $Y2=2.027
r90 31 32 65.6923 $w=1.93e-07 $l=1.155e-06 $layer=LI1_cond $X=2.605 $Y=2.027
+ $X2=1.45 $Y2=2.027
r91 27 34 0.966048 $w=3e-07 $l=1.73e-07 $layer=LI1_cond $X=1.3 $Y=2.275 $X2=1.3
+ $Y2=2.102
r92 27 29 7.10673 $w=2.98e-07 $l=1.85e-07 $layer=LI1_cond $X=1.3 $Y=2.275
+ $X2=1.3 $Y2=2.46
r93 25 34 5.63431 $w=2.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.15 $Y=2.102 $X2=1.3
+ $Y2=2.102
r94 25 26 25.7212 $w=3.43e-07 $l=7.7e-07 $layer=LI1_cond $X=1.15 $Y=2.102
+ $X2=0.38 $Y2=2.102
r95 23 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=0.945
+ $X2=1.335 $Y2=0.78
r96 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.335
+ $Y=0.945 $X2=1.335 $Y2=0.945
r97 20 33 0.982774 $w=2.35e-07 $l=1.13e-07 $layer=LI1_cond $X=0.38 $Y=0.912
+ $X2=0.267 $Y2=0.912
r98 20 22 46.8333 $w=2.33e-07 $l=9.55e-07 $layer=LI1_cond $X=0.38 $Y=0.912
+ $X2=1.335 $Y2=0.912
r99 19 26 7.21695 $w=3.45e-07 $l=2.21405e-07 $layer=LI1_cond $X=0.267 $Y=1.93
+ $X2=0.38 $Y2=2.102
r100 18 33 5.61269 $w=2.12e-07 $l=1.18e-07 $layer=LI1_cond $X=0.267 $Y=1.03
+ $X2=0.267 $Y2=0.912
r101 18 19 46.0977 $w=2.23e-07 $l=9e-07 $layer=LI1_cond $X=0.267 $Y=1.03
+ $X2=0.267 $Y2=1.93
r102 14 33 5.61269 $w=2.12e-07 $l=1.22854e-07 $layer=LI1_cond $X=0.255 $Y=0.795
+ $X2=0.267 $Y2=0.912
r103 14 16 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=0.255 $Y=0.795
+ $X2=0.255 $Y2=0.58
r104 12 46 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.75 $Y=2.635
+ $X2=2.75 $Y2=2.1
r105 9 42 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.425 $Y=0.46
+ $X2=1.425 $Y2=0.78
r106 2 29 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.19
+ $Y=2.315 $X2=1.315 $Y2=2.46
r107 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.26 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%SCE 3 6 7 8 9 11 12 14 16 19 21 26 27 28 29
+ 30 31 43
r82 40 43 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.265 $Y=1.295
+ $X2=2.445 $Y2=1.295
r83 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.265
+ $Y=1.295 $X2=2.265 $Y2=1.295
r84 31 41 21.3287 $w=1.93e-07 $l=3.75e-07 $layer=LI1_cond $X=2.64 $Y=1.302
+ $X2=2.265 $Y2=1.302
r85 30 41 5.97203 $w=1.93e-07 $l=1.05e-07 $layer=LI1_cond $X=2.16 $Y=1.302
+ $X2=2.265 $Y2=1.302
r86 29 30 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.302
+ $X2=2.16 $Y2=1.302
r87 28 29 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.302
+ $X2=1.68 $Y2=1.302
r88 27 38 83.87 $w=4.8e-07 $l=5.05e-07 $layer=POLY_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.8
r89 27 37 45.9721 $w=4.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.13
r90 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.715
+ $Y=1.295 $X2=0.715 $Y2=1.295
r91 24 28 18.2005 $w=1.93e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=1.302
+ $X2=1.2 $Y2=1.302
r92 24 26 4.65494 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=1.302
+ $X2=0.715 $Y2=1.302
r93 17 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=1.13
+ $X2=2.445 $Y2=1.295
r94 17 19 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.445 $Y=1.13
+ $X2=2.445 $Y2=0.615
r95 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.96 $Y=2.205
+ $X2=1.96 $Y2=2.635
r96 13 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.605 $Y=2.13
+ $X2=1.53 $Y2=2.13
r97 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.885 $Y=2.13
+ $X2=1.96 $Y2=2.205
r98 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.885 $Y=2.13
+ $X2=1.605 $Y2=2.13
r99 9 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.53 $Y=2.205
+ $X2=1.53 $Y2=2.13
r100 9 11 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.53 $Y=2.205
+ $X2=1.53 $Y2=2.635
r101 7 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.455 $Y=2.13
+ $X2=1.53 $Y2=2.13
r102 7 8 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.455 $Y=2.13
+ $X2=0.55 $Y2=2.13
r103 6 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=2.055
+ $X2=0.55 $Y2=2.13
r104 6 38 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.475 $Y=2.055
+ $X2=0.475 $Y2=1.8
r105 3 37 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.475 $Y=0.58
+ $X2=0.475 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%D 3 5 9 11 12 13 18
c44 9 0 1.29538e-19 $X=2.32 $Y=2.635
r45 18 21 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.755
r46 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.5
r47 12 13 28.0191 $w=1.88e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=2.16 $Y2=1.665
r48 12 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.695
+ $Y=1.665 $X2=1.695 $Y2=1.665
r49 11 12 28.0191 $w=1.88e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.68 $Y2=1.665
r50 7 9 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=2.32 $Y=1.83 $X2=2.32
+ $Y2=2.635
r51 6 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.86 $Y=1.755
+ $X2=1.695 $Y2=1.755
r52 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.245 $Y=1.755
+ $X2=2.32 $Y2=1.83
r53 5 6 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.245 $Y=1.755
+ $X2=1.86 $Y2=1.755
r54 3 20 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.785 $Y=0.46
+ $X2=1.785 $Y2=1.5
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%SCD 3 5 6 9 13 14 15 19 20
c48 20 0 2.47684e-19 $X=3.31 $Y=1.455
c49 9 0 6.53831e-20 $X=3.22 $Y=2.635
c50 3 0 3.56444e-20 $X=2.805 $Y=0.615
r51 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.31
+ $Y=1.455 $X2=3.31 $Y2=1.455
r52 14 15 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.25 $Y=1.665
+ $X2=3.25 $Y2=2.035
r53 14 20 5.5817 $w=4.48e-07 $l=2.1e-07 $layer=LI1_cond $X=3.25 $Y=1.665
+ $X2=3.25 $Y2=1.455
r54 12 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.31 $Y=1.795
+ $X2=3.31 $Y2=1.455
r55 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.795
+ $X2=3.31 $Y2=1.96
r56 11 19 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.31 $Y=1.44
+ $X2=3.31 $Y2=1.455
r57 9 13 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=1.96
r58 5 11 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.145 $Y=1.365
+ $X2=3.31 $Y2=1.44
r59 5 6 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.145 $Y=1.365
+ $X2=2.88 $Y2=1.365
r60 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.805 $Y=1.29
+ $X2=2.88 $Y2=1.365
r61 1 3 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.805 $Y=1.29
+ $X2=2.805 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%A_851_242# 1 2 9 13 14 16 17 18 21 24 26 27
+ 31 32 36 39 40 41 42 43 44 47 56 57 60 64 65 66 68
c214 65 0 2.69883e-19 $X=5.48 $Y=1.29
c215 42 0 1.62646e-19 $X=5.665 $Y=1.295
c216 40 0 1.4984e-20 $X=4.705 $Y=1.295
c217 32 0 3.68148e-20 $X=8.375 $Y=2.22
c218 26 0 5.89179e-20 $X=8.275 $Y=2.055
r219 68 71 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8 $Y=1.17 $X2=8
+ $Y2=1.26
r220 64 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.48 $Y=1.29
+ $X2=5.48 $Y2=1.125
r221 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.48
+ $Y=1.29 $X2=5.48 $Y2=1.29
r222 57 88 30.9578 $w=2.53e-07 $l=6.85e-07 $layer=LI1_cond $X=10.792 $Y=1.295
+ $X2=10.792 $Y2=1.98
r223 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=1.295
+ $X2=10.8 $Y2=1.295
r224 54 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8 $Y=1.26
+ $X2=8 $Y2=1.26
r225 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.295
+ $X2=7.92 $Y2=1.295
r226 50 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r227 47 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.5
+ $Y=1.375 $X2=4.5 $Y2=1.375
r228 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=1.295
+ $X2=4.56 $Y2=1.295
r229 44 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=1.295
+ $X2=7.92 $Y2=1.295
r230 43 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=1.295
+ $X2=10.8 $Y2=1.295
r231 43 44 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=1.295
+ $X2=8.065 $Y2=1.295
r232 42 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.295
+ $X2=5.52 $Y2=1.295
r233 41 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=1.295
+ $X2=7.92 $Y2=1.295
r234 41 42 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=7.775 $Y=1.295
+ $X2=5.665 $Y2=1.295
r235 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=1.295
+ $X2=4.56 $Y2=1.295
r236 39 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=5.52 $Y2=1.295
r237 39 40 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=4.705 $Y2=1.295
r238 38 57 5.8752 $w=2.53e-07 $l=1.3e-07 $layer=LI1_cond $X=10.792 $Y=1.165
+ $X2=10.792 $Y2=1.295
r239 36 38 4.29215 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=10.83 $Y=1.06
+ $X2=10.83 $Y2=1.165
r240 32 74 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=8.375 $Y=2.22
+ $X2=8.235 $Y2=2.22
r241 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.375
+ $Y=2.22 $X2=8.375 $Y2=2.22
r242 28 31 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=8.275 $Y=2.185
+ $X2=8.375 $Y2=2.185
r243 27 54 14.6075 $w=2.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.19 $Y=1.277
+ $X2=7.92 $Y2=1.277
r244 26 28 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.275 $Y=2.055
+ $X2=8.275 $Y2=2.185
r245 25 27 6.89401 $w=2.05e-07 $l=1.39155e-07 $layer=LI1_cond $X=8.275 $Y=1.38
+ $X2=8.19 $Y2=1.277
r246 25 26 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=8.275 $Y=1.38
+ $X2=8.275 $Y2=2.055
r247 23 60 40.6942 $w=4.1e-07 $l=3e-07 $layer=POLY_cond $X=4.46 $Y=1.675
+ $X2=4.46 $Y2=1.375
r248 23 24 51.3336 $w=4.1e-07 $l=2.05e-07 $layer=POLY_cond $X=4.46 $Y=1.675
+ $X2=4.46 $Y2=1.88
r249 19 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.235 $Y=2.385
+ $X2=8.235 $Y2=2.22
r250 19 21 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=8.235 $Y=2.385
+ $X2=8.235 $Y2=2.875
r251 17 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.835 $Y=1.17
+ $X2=8 $Y2=1.17
r252 17 18 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=7.835 $Y=1.17
+ $X2=7.62 $Y2=1.17
r253 14 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.545 $Y=1.095
+ $X2=7.62 $Y2=1.17
r254 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.545 $Y=1.095
+ $X2=7.545 $Y2=0.665
r255 13 66 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.46 $Y=0.805
+ $X2=5.46 $Y2=1.125
r256 9 24 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.33 $Y=2.525
+ $X2=4.33 $Y2=1.88
r257 2 88 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=10.7
+ $Y=1.835 $X2=10.825 $Y2=1.98
r258 1 36 182 $w=1.7e-07 $l=7.84156e-07 $layer=licon1_NDIFF $count=1 $X=10.685
+ $Y=0.345 $X2=10.83 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%A_1047_369# 1 2 9 11 12 15 22 26 29 30 31
+ 32 36
c102 11 0 1.12934e-19 $X=5.855 $Y=1.74
r103 30 31 8.67671 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=5.87 $Y=1.76
+ $X2=6.04 $Y2=1.76
r104 29 36 9.91637 $w=2.13e-07 $l=1.85e-07 $layer=LI1_cond $X=7.215 $Y=2.007
+ $X2=7.4 $Y2=2.007
r105 28 32 4.40882 $w=2.05e-07 $l=8.74643e-08 $layer=LI1_cond $X=7.215 $Y=1.725
+ $X2=7.21 $Y2=1.64
r106 28 29 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=7.215 $Y=1.725
+ $X2=7.215 $Y2=1.9
r107 24 32 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.21 $Y=1.555
+ $X2=7.21 $Y2=1.64
r108 24 26 55.7186 $w=2.08e-07 $l=1.055e-06 $layer=LI1_cond $X=7.21 $Y=1.555
+ $X2=7.21 $Y2=0.5
r109 22 32 2.0246 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.105 $Y=1.64
+ $X2=7.21 $Y2=1.64
r110 22 31 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=7.105 $Y=1.64
+ $X2=6.04 $Y2=1.64
r111 20 38 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=5.43 $Y=1.83
+ $X2=5.31 $Y2=1.83
r112 19 30 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=5.43 $Y=1.815
+ $X2=5.87 $Y2=1.815
r113 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.43
+ $Y=1.83 $X2=5.43 $Y2=1.83
r114 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.93 $Y=1.665
+ $X2=5.93 $Y2=0.805
r115 12 20 38.5363 $w=3.15e-07 $l=2.05122e-07 $layer=POLY_cond $X=5.595 $Y=1.74
+ $X2=5.43 $Y2=1.83
r116 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.855 $Y=1.74
+ $X2=5.93 $Y2=1.665
r117 11 12 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.855 $Y=1.74
+ $X2=5.595 $Y2=1.74
r118 7 38 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.995
+ $X2=5.31 $Y2=1.83
r119 7 9 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.31 $Y=1.995
+ $X2=5.31 $Y2=2.525
r120 2 36 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.895 $X2=7.4 $Y2=2.02
r121 1 26 91 $w=1.7e-07 $l=3.02738e-07 $layer=licon1_NDIFF $count=2 $X=6.985
+ $Y=0.345 $X2=7.22 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%RESET_B 3 5 6 9 11 13 15 16 17 21 24 28 30
+ 32 33 34 36 37 38 39 41 46 47 51 54 66
c185 47 0 2.58091e-20 $X=9.525 $Y=2.34
c186 3 0 3.04204e-19 $X=3.235 $Y=0.615
r187 54 56 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.382 $Y=1.99
+ $X2=6.382 $Y2=1.825
r188 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.385
+ $Y=1.99 $X2=6.385 $Y2=1.99
r189 51 66 0.735602 $w=2.33e-07 $l=1.5e-08 $layer=LI1_cond $X=6.48 $Y=2.012
+ $X2=6.495 $Y2=2.012
r190 51 55 4.65881 $w=2.33e-07 $l=9.5e-08 $layer=LI1_cond $X=6.48 $Y=2.012
+ $X2=6.385 $Y2=2.012
r191 47 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.525 $Y=2.34
+ $X2=9.525 $Y2=2.505
r192 47 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.525 $Y=2.34
+ $X2=9.525 $Y2=2.175
r193 46 49 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=9.525 $Y=2.34
+ $X2=9.525 $Y2=2.57
r194 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.525
+ $Y=2.34 $X2=9.525 $Y2=2.34
r195 41 43 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.275 $Y=2.57
+ $X2=8.275 $Y2=2.81
r196 40 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=2.57
+ $X2=8.275 $Y2=2.57
r197 39 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.36 $Y=2.57
+ $X2=9.525 $Y2=2.57
r198 39 40 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=9.36 $Y=2.57 $X2=8.36
+ $Y2=2.57
r199 37 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.19 $Y=2.81
+ $X2=8.275 $Y2=2.81
r200 37 38 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=8.19 $Y=2.81
+ $X2=7.37 $Y2=2.81
r201 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.285 $Y=2.725
+ $X2=7.37 $Y2=2.81
r202 35 36 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.285 $Y=2.455
+ $X2=7.285 $Y2=2.725
r203 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.2 $Y=2.37
+ $X2=7.285 $Y2=2.455
r204 33 34 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.2 $Y=2.37
+ $X2=6.58 $Y2=2.37
r205 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.495 $Y=2.285
+ $X2=6.58 $Y2=2.37
r206 31 66 2.6346 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=6.495 $Y=2.13
+ $X2=6.495 $Y2=2.012
r207 31 32 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.495 $Y=2.13
+ $X2=6.495 $Y2=2.285
r208 28 61 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.545 $Y=2.875
+ $X2=9.545 $Y2=2.505
r209 24 60 702.489 $w=1.5e-07 $l=1.37e-06 $layer=POLY_cond $X=9.435 $Y=0.805
+ $X2=9.435 $Y2=2.175
r210 21 56 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=6.29 $Y=0.805
+ $X2=6.29 $Y2=1.825
r211 18 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.29 $Y=0.255
+ $X2=6.29 $Y2=0.805
r212 16 54 24.1152 $w=3.35e-07 $l=1.4e-07 $layer=POLY_cond $X=6.382 $Y=2.13
+ $X2=6.382 $Y2=1.99
r213 16 17 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.215 $Y=2.13
+ $X2=5.985 $Y2=2.13
r214 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.91 $Y=2.205
+ $X2=5.985 $Y2=2.13
r215 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.91 $Y=2.205
+ $X2=5.91 $Y2=2.525
r216 12 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.88 $Y=0.18
+ $X2=3.805 $Y2=0.18
r217 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.215 $Y=0.18
+ $X2=6.29 $Y2=0.255
r218 11 12 1197.31 $w=1.5e-07 $l=2.335e-06 $layer=POLY_cond $X=6.215 $Y=0.18
+ $X2=3.88 $Y2=0.18
r219 7 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.805 $Y=0.255
+ $X2=3.805 $Y2=0.18
r220 7 9 1220.38 $w=1.5e-07 $l=2.38e-06 $layer=POLY_cond $X=3.805 $Y=0.255
+ $X2=3.805 $Y2=2.635
r221 5 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.73 $Y=0.18
+ $X2=3.805 $Y2=0.18
r222 5 6 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.73 $Y=0.18 $X2=3.31
+ $Y2=0.18
r223 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.235 $Y=0.255
+ $X2=3.31 $Y2=0.18
r224 1 3 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.235 $Y=0.255
+ $X2=3.235 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%A_881_463# 1 2 3 12 16 19 20 23 24 25 29 30
+ 32 35 40 46
c141 20 0 1.12934e-19 $X=5.87 $Y=2.22
c142 16 0 7.80833e-20 $X=7.185 $Y=2.315
r143 38 40 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.905 $Y=1.295
+ $X2=5.13 $Y2=1.295
r144 35 37 8.00215 $w=4.65e-07 $l=3.05e-07 $layer=LI1_cond $X=4.7 $Y=2.22
+ $X2=4.7 $Y2=2.525
r145 33 46 26.5669 $w=2.54e-07 $l=1.4e-07 $layer=POLY_cond $X=6.77 $Y=1.29
+ $X2=6.91 $Y2=1.29
r146 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.77
+ $Y=1.29 $X2=6.77 $Y2=1.29
r147 30 32 42.6928 $w=2.18e-07 $l=8.15e-07 $layer=LI1_cond $X=5.955 $Y=1.275
+ $X2=6.77 $Y2=1.275
r148 29 30 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.87 $Y=1.165
+ $X2=5.955 $Y2=1.275
r149 28 29 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.87 $Y=0.955
+ $X2=5.87 $Y2=1.165
r150 25 27 1.09756 $w=3.13e-07 $l=3e-08 $layer=LI1_cond $X=5.215 $Y=0.797
+ $X2=5.245 $Y2=0.797
r151 24 28 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=5.785 $Y=0.797
+ $X2=5.87 $Y2=0.955
r152 24 27 19.7562 $w=3.13e-07 $l=5.4e-07 $layer=LI1_cond $X=5.785 $Y=0.797
+ $X2=5.245 $Y2=0.797
r153 23 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.13 $Y=1.21
+ $X2=5.13 $Y2=1.295
r154 22 25 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=5.13 $Y=0.955
+ $X2=5.215 $Y2=0.797
r155 22 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.13 $Y=0.955
+ $X2=5.13 $Y2=1.21
r156 21 35 6.7035 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.995 $Y=2.22
+ $X2=4.7 $Y2=2.22
r157 20 44 12.9201 $w=2.88e-07 $l=3.86588e-07 $layer=LI1_cond $X=5.87 $Y=2.22
+ $X2=6.055 $Y2=2.525
r158 20 21 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=5.87 $Y=2.22
+ $X2=4.995 $Y2=2.22
r159 19 35 6.99515 $w=4.65e-07 $l=2.43824e-07 $layer=LI1_cond $X=4.905 $Y=2.135
+ $X2=4.7 $Y2=2.22
r160 18 38 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=1.38
+ $X2=4.905 $Y2=1.295
r161 18 19 46.5202 $w=1.78e-07 $l=7.55e-07 $layer=LI1_cond $X=4.905 $Y=1.38
+ $X2=4.905 $Y2=2.135
r162 14 46 52.185 $w=2.54e-07 $l=3.47851e-07 $layer=POLY_cond $X=7.185 $Y=1.455
+ $X2=6.91 $Y2=1.29
r163 14 16 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.185 $Y=1.455
+ $X2=7.185 $Y2=2.315
r164 10 46 15.087 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.91 $Y=1.125
+ $X2=6.91 $Y2=1.29
r165 10 12 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=6.91 $Y=1.125
+ $X2=6.91 $Y2=0.665
r166 3 44 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.985
+ $Y=2.315 $X2=6.125 $Y2=2.525
r167 2 37 600 $w=1.7e-07 $l=3.23381e-07 $layer=licon1_PDIFF $count=1 $X=4.405
+ $Y=2.315 $X2=4.64 $Y2=2.525
r168 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.595 $X2=5.245 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%A_975_255# 1 2 10 13 15 16 20 22 25 29 33
+ 37 39 42 43 44 45 46 47 50 55 57 60 64 66 68 69 72
c203 66 0 1.28163e-19 $X=11.887 $Y=1.51
c204 57 0 9.8418e-20 $X=8.79 $Y=1.65
c205 37 0 3.54913e-19 $X=5.03 $Y=1.35
c206 22 0 5.89179e-20 $X=7.69 $Y=1.74
c207 13 0 4.8898e-21 $X=5.03 $Y=0.805
c208 10 0 8.77104e-20 $X=4.95 $Y=2.525
r209 71 72 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.45 $Y=1.65
+ $X2=8.375 $Y2=1.65
r210 68 69 8.46863 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=11.932 $Y=2.835
+ $X2=11.932 $Y2=2.67
r211 61 64 3.96938 $w=1.88e-07 $l=6.8e-08 $layer=LI1_cond $X=11.887 $Y=1.07
+ $X2=11.955 $Y2=1.07
r212 60 77 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.155 $Y=1.51
+ $X2=11.155 $Y2=1.675
r213 60 76 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.155 $Y=1.51
+ $X2=11.155 $Y2=1.345
r214 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.175
+ $Y=1.51 $X2=11.175 $Y2=1.51
r215 55 71 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=8.625 $Y=1.65
+ $X2=8.45 $Y2=1.65
r216 54 57 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=1.65
+ $X2=8.79 $Y2=1.65
r217 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.625
+ $Y=1.65 $X2=8.625 $Y2=1.65
r218 51 66 8.03064 $w=1.87e-07 $l=1.68953e-07 $layer=LI1_cond $X=11.895 $Y=1.675
+ $X2=11.887 $Y2=1.51
r219 51 69 61.3081 $w=1.78e-07 $l=9.95e-07 $layer=LI1_cond $X=11.895 $Y=1.675
+ $X2=11.895 $Y2=2.67
r220 50 66 8.03064 $w=1.87e-07 $l=1.65e-07 $layer=LI1_cond $X=11.887 $Y=1.345
+ $X2=11.887 $Y2=1.51
r221 49 61 0.589566 $w=1.95e-07 $l=9.5e-08 $layer=LI1_cond $X=11.887 $Y=1.165
+ $X2=11.887 $Y2=1.07
r222 49 50 10.2378 $w=1.93e-07 $l=1.8e-07 $layer=LI1_cond $X=11.887 $Y=1.165
+ $X2=11.887 $Y2=1.345
r223 48 59 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.26 $Y=1.51
+ $X2=11.175 $Y2=1.51
r224 47 66 0.588983 $w=3.3e-07 $l=9.7e-08 $layer=LI1_cond $X=11.79 $Y=1.51
+ $X2=11.887 $Y2=1.51
r225 47 48 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=11.79 $Y=1.51
+ $X2=11.26 $Y2=1.51
r226 45 59 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.175 $Y=1.675
+ $X2=11.175 $Y2=1.51
r227 45 46 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=11.175 $Y=1.675
+ $X2=11.175 $Y2=2.325
r228 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.09 $Y=2.41
+ $X2=11.175 $Y2=2.325
r229 43 44 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=11.09 $Y=2.41
+ $X2=10.39 $Y2=2.41
r230 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.305 $Y=2.325
+ $X2=10.39 $Y2=2.41
r231 41 42 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=10.305 $Y=1.725
+ $X2=10.305 $Y2=2.325
r232 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.22 $Y=1.64
+ $X2=10.305 $Y2=1.725
r233 39 57 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=10.22 $Y=1.64
+ $X2=8.79 $Y2=1.64
r234 35 37 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=4.95 $Y=1.35 $X2=5.03
+ $Y2=1.35
r235 33 77 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.045 $Y=2.465
+ $X2=11.045 $Y2=1.675
r236 29 76 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.045 $Y=0.765
+ $X2=11.045 $Y2=1.345
r237 23 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.45 $Y=1.485
+ $X2=8.45 $Y2=1.65
r238 23 25 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=8.45 $Y=1.485
+ $X2=8.45 $Y2=0.775
r239 22 72 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=7.69 $Y=1.74
+ $X2=8.375 $Y2=1.74
r240 18 20 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.615 $Y=3.075
+ $X2=7.615 $Y2=2.315
r241 17 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.615 $Y=1.815
+ $X2=7.69 $Y2=1.74
r242 17 20 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.615 $Y=1.815
+ $X2=7.615 $Y2=2.315
r243 15 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.54 $Y=3.15
+ $X2=7.615 $Y2=3.075
r244 15 16 1289.61 $w=1.5e-07 $l=2.515e-06 $layer=POLY_cond $X=7.54 $Y=3.15
+ $X2=5.025 $Y2=3.15
r245 11 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.03 $Y=1.275
+ $X2=5.03 $Y2=1.35
r246 11 13 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.03 $Y=1.275 $X2=5.03
+ $Y2=0.805
r247 8 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.95 $Y=3.075
+ $X2=5.025 $Y2=3.15
r248 8 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.95 $Y=3.075
+ $X2=4.95 $Y2=2.525
r249 7 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.95 $Y=1.425
+ $X2=4.95 $Y2=1.35
r250 7 10 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=4.95 $Y=1.425
+ $X2=4.95 $Y2=2.525
r251 2 68 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=11.815
+ $Y=1.835 $X2=11.955 $Y2=2.835
r252 1 64 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=11.815
+ $Y=0.345 $X2=11.955 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%A_1524_69# 1 2 9 12 16 19 22 23 24 29 31 34
+ 36 38 39 40 42 43 44 51 52 53 59 62 65
c185 31 0 7.80833e-20 $X=7.9 $Y=2.04
r186 59 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.025 $Y=1.35
+ $X2=13.025 $Y2=1.515
r187 59 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.025 $Y=1.35
+ $X2=13.025 $Y2=1.185
r188 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.025
+ $Y=1.35 $X2=13.025 $Y2=1.35
r189 51 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.885 $Y=1.29
+ $X2=9.885 $Y2=1.455
r190 51 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.885 $Y=1.29
+ $X2=9.885 $Y2=1.125
r191 50 53 24.7295 $w=2.38e-07 $l=5.15e-07 $layer=LI1_cond $X=9.885 $Y=1.255
+ $X2=10.4 $Y2=1.255
r192 50 52 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=9.885 $Y=1.255
+ $X2=9.72 $Y2=1.255
r193 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.885
+ $Y=1.29 $X2=9.885 $Y2=1.29
r194 43 58 3.35256 $w=2.73e-07 $l=8e-08 $layer=LI1_cond $X=12.997 $Y=1.27
+ $X2=12.997 $Y2=1.35
r195 43 44 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=12.86 $Y=1.27
+ $X2=12.47 $Y2=1.27
r196 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.385 $Y=1.185
+ $X2=12.47 $Y2=1.27
r197 41 42 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=12.385 $Y=0.795
+ $X2=12.385 $Y2=1.185
r198 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.3 $Y=0.71
+ $X2=12.385 $Y2=0.795
r199 39 40 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=12.3 $Y=0.71
+ $X2=10.485 $Y2=0.71
r200 38 53 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=10.4 $Y=1.135
+ $X2=10.4 $Y2=1.255
r201 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.4 $Y=0.795
+ $X2=10.485 $Y2=0.71
r202 37 38 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=10.4 $Y=0.795
+ $X2=10.4 $Y2=1.135
r203 36 52 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=8.71 $Y=1.22
+ $X2=9.72 $Y2=1.22
r204 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.625 $Y=1.135
+ $X2=8.71 $Y2=1.22
r205 33 34 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=8.625 $Y=0.945
+ $X2=8.625 $Y2=1.135
r206 29 45 20.0289 $w=1.68e-07 $l=3.07e-07 $layer=LI1_cond $X=7.877 $Y=1.645
+ $X2=7.57 $Y2=1.645
r207 29 31 12.5353 $w=2.83e-07 $l=3.1e-07 $layer=LI1_cond $X=7.877 $Y=1.73
+ $X2=7.877 $Y2=2.04
r208 26 28 10.3298 $w=5.48e-07 $l=4.75e-07 $layer=LI1_cond $X=7.76 $Y=0.67
+ $X2=8.235 $Y2=0.67
r209 24 26 2.28342 $w=5.48e-07 $l=1.05e-07 $layer=LI1_cond $X=7.655 $Y=0.67
+ $X2=7.76 $Y2=0.67
r210 23 33 9.64472 $w=5.5e-07 $l=3.14643e-07 $layer=LI1_cond $X=8.54 $Y=0.67
+ $X2=8.625 $Y2=0.945
r211 23 28 6.6328 $w=5.48e-07 $l=3.05e-07 $layer=LI1_cond $X=8.54 $Y=0.67
+ $X2=8.235 $Y2=0.67
r212 22 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.57 $Y=1.56
+ $X2=7.57 $Y2=1.645
r213 21 24 9.64472 $w=5.5e-07 $l=3.14643e-07 $layer=LI1_cond $X=7.57 $Y=0.945
+ $X2=7.655 $Y2=0.67
r214 21 22 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=7.57 $Y=0.945
+ $X2=7.57 $Y2=1.56
r215 19 66 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=13.115 $Y=2.465
+ $X2=13.115 $Y2=1.515
r216 16 65 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=13.115 $Y=0.655
+ $X2=13.115 $Y2=1.185
r217 12 63 728.128 $w=1.5e-07 $l=1.42e-06 $layer=POLY_cond $X=9.975 $Y=2.875
+ $X2=9.975 $Y2=1.455
r218 9 62 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.795 $Y=0.805
+ $X2=9.795 $Y2=1.125
r219 2 31 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=1.895 $X2=7.9 $Y2=2.04
r220 1 28 182 $w=1.7e-07 $l=7.97825e-07 $layer=licon1_NDIFF $count=1 $X=7.62
+ $Y=0.345 $X2=8.235 $Y2=0.765
r221 1 26 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=7.62
+ $Y=0.345 $X2=7.76 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%A_1747_21# 1 2 10 13 15 16 18 21 23 25 31
+ 34 35 37 40 47 49
c111 21 0 6.16032e-20 $X=9.075 $Y=1.17
r112 43 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.985 $Y=2.22
+ $X2=9.075 $Y2=2.22
r113 43 44 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=8.985 $Y=2.22
+ $X2=8.825 $Y2=2.22
r114 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.985
+ $Y=2.22 $X2=8.985 $Y2=2.22
r115 40 42 10.3542 $w=2.71e-07 $l=2.3e-07 $layer=LI1_cond $X=8.985 $Y=1.99
+ $X2=8.985 $Y2=2.22
r116 38 49 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=10.41 $Y=0.35
+ $X2=10.41 $Y2=0.18
r117 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.41
+ $Y=0.35 $X2=10.41 $Y2=0.35
r118 35 37 14.6955 $w=1.98e-07 $l=2.65e-07 $layer=LI1_cond $X=10.145 $Y=0.355
+ $X2=10.41 $Y2=0.355
r119 33 34 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=9.955 $Y=2.075
+ $X2=9.955 $Y2=2.825
r120 29 35 7.17723 $w=2e-07 $l=1.93649e-07 $layer=LI1_cond $X=9.995 $Y=0.455
+ $X2=10.145 $Y2=0.355
r121 29 31 13.2531 $w=2.98e-07 $l=3.45e-07 $layer=LI1_cond $X=9.995 $Y=0.455
+ $X2=9.995 $Y2=0.8
r122 25 34 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=9.87 $Y=2.935
+ $X2=9.955 $Y2=2.825
r123 25 27 5.76222 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=9.87 $Y=2.935
+ $X2=9.76 $Y2=2.935
r124 24 40 3.46554 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.15 $Y=1.99
+ $X2=8.985 $Y2=1.99
r125 23 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.87 $Y=1.99
+ $X2=9.955 $Y2=2.075
r126 23 24 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=9.87 $Y=1.99
+ $X2=9.15 $Y2=1.99
r127 19 21 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=8.81 $Y=1.17
+ $X2=9.075 $Y2=1.17
r128 18 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.075 $Y=2.055
+ $X2=9.075 $Y2=2.22
r129 17 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.075 $Y=1.245
+ $X2=9.075 $Y2=1.17
r130 17 18 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.075 $Y=1.245
+ $X2=9.075 $Y2=2.055
r131 15 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.245 $Y=0.18
+ $X2=10.41 $Y2=0.18
r132 15 16 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=10.245 $Y=0.18
+ $X2=8.885 $Y2=0.18
r133 11 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.825 $Y=2.385
+ $X2=8.825 $Y2=2.22
r134 11 13 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=8.825 $Y=2.385
+ $X2=8.825 $Y2=2.875
r135 8 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.81 $Y=1.095
+ $X2=8.81 $Y2=1.17
r136 8 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.81 $Y=1.095
+ $X2=8.81 $Y2=0.775
r137 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.81 $Y=0.255
+ $X2=8.885 $Y2=0.18
r138 7 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=8.81 $Y=0.255
+ $X2=8.81 $Y2=0.775
r139 2 27 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=9.62
+ $Y=2.665 $X2=9.76 $Y2=2.94
r140 1 31 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=9.87
+ $Y=0.595 $X2=10.01 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%CLK 3 7 9 11 13 14 15 20 21
r52 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.405
+ $Y=1.625 $X2=12.405 $Y2=1.625
r53 14 15 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=12.362 $Y=2.035
+ $X2=12.362 $Y2=2.405
r54 13 14 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=12.362 $Y=1.665
+ $X2=12.362 $Y2=2.035
r55 13 21 1.11079 $w=4.13e-07 $l=4e-08 $layer=LI1_cond $X=12.362 $Y=1.665
+ $X2=12.362 $Y2=1.625
r56 12 20 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=12.405 $Y=1.61
+ $X2=12.405 $Y2=1.625
r57 10 11 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.815 $Y=1.535
+ $X2=11.74 $Y2=1.535
r58 9 12 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=12.24 $Y=1.535
+ $X2=12.405 $Y2=1.61
r59 9 10 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=12.24 $Y=1.535
+ $X2=11.815 $Y2=1.535
r60 5 11 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.74 $Y=1.61
+ $X2=11.74 $Y2=1.535
r61 5 7 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=11.74 $Y=1.61
+ $X2=11.74 $Y2=2.465
r62 1 11 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.74 $Y=1.46
+ $X2=11.74 $Y2=1.535
r63 1 3 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=11.74 $Y=1.46
+ $X2=11.74 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%A_2555_47# 1 2 9 13 17 21 25 29 33 37 41 45
+ 49 50 51 52 54 56 62 65 73
r118 70 71 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=14.405 $Y=1.48
+ $X2=14.445 $Y2=1.48
r119 69 70 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=13.975 $Y=1.48
+ $X2=14.405 $Y2=1.48
r120 63 73 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=14.655 $Y=1.48
+ $X2=14.875 $Y2=1.48
r121 63 71 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=14.655 $Y=1.48
+ $X2=14.445 $Y2=1.48
r122 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.655
+ $Y=1.48 $X2=14.655 $Y2=1.48
r123 60 69 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=13.635 $Y=1.48
+ $X2=13.975 $Y2=1.48
r124 60 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=13.635 $Y=1.48
+ $X2=13.545 $Y2=1.48
r125 59 62 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=13.635 $Y=1.48
+ $X2=14.655 $Y2=1.48
r126 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.635
+ $Y=1.48 $X2=13.635 $Y2=1.48
r127 57 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.475 $Y=1.48
+ $X2=13.39 $Y2=1.48
r128 57 59 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=13.475 $Y=1.48
+ $X2=13.635 $Y2=1.48
r129 55 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.39 $Y=1.565
+ $X2=13.39 $Y2=1.48
r130 55 56 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=13.39 $Y=1.565
+ $X2=13.39 $Y2=1.755
r131 54 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.39 $Y=1.395
+ $X2=13.39 $Y2=1.48
r132 53 54 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=13.39 $Y=1.015
+ $X2=13.39 $Y2=1.395
r133 51 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.305 $Y=1.84
+ $X2=13.39 $Y2=1.755
r134 51 52 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=13.305 $Y=1.84
+ $X2=12.995 $Y2=1.84
r135 49 53 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=13.305 $Y=0.925
+ $X2=13.39 $Y2=1.015
r136 49 50 19.101 $w=1.78e-07 $l=3.1e-07 $layer=LI1_cond $X=13.305 $Y=0.925
+ $X2=12.995 $Y2=0.925
r137 45 47 42.0303 $w=2.53e-07 $l=9.3e-07 $layer=LI1_cond $X=12.867 $Y=1.98
+ $X2=12.867 $Y2=2.91
r138 43 52 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=12.867 $Y=1.925
+ $X2=12.995 $Y2=1.84
r139 43 45 2.48566 $w=2.53e-07 $l=5.5e-08 $layer=LI1_cond $X=12.867 $Y=1.925
+ $X2=12.867 $Y2=1.98
r140 39 50 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=12.865 $Y=0.835
+ $X2=12.995 $Y2=0.925
r141 39 41 18.3948 $w=2.58e-07 $l=4.15e-07 $layer=LI1_cond $X=12.865 $Y=0.835
+ $X2=12.865 $Y2=0.42
r142 35 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.875 $Y=1.645
+ $X2=14.875 $Y2=1.48
r143 35 37 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=14.875 $Y=1.645
+ $X2=14.875 $Y2=2.465
r144 31 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.875 $Y=1.315
+ $X2=14.875 $Y2=1.48
r145 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.875 $Y=1.315
+ $X2=14.875 $Y2=0.655
r146 27 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.445 $Y=1.645
+ $X2=14.445 $Y2=1.48
r147 27 29 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=14.445 $Y=1.645
+ $X2=14.445 $Y2=2.465
r148 23 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.405 $Y=1.315
+ $X2=14.405 $Y2=1.48
r149 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.405 $Y=1.315
+ $X2=14.405 $Y2=0.655
r150 19 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.975 $Y=1.645
+ $X2=13.975 $Y2=1.48
r151 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=13.975 $Y=1.645
+ $X2=13.975 $Y2=2.465
r152 15 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.975 $Y=1.315
+ $X2=13.975 $Y2=1.48
r153 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.975 $Y=1.315
+ $X2=13.975 $Y2=0.655
r154 11 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.545 $Y=1.645
+ $X2=13.545 $Y2=1.48
r155 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=13.545 $Y=1.645
+ $X2=13.545 $Y2=2.465
r156 7 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.545 $Y=1.315
+ $X2=13.545 $Y2=1.48
r157 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.545 $Y=1.315
+ $X2=13.545 $Y2=0.655
r158 2 47 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=12.775
+ $Y=1.835 $X2=12.9 $Y2=2.91
r159 2 45 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=12.775
+ $Y=1.835 $X2=12.9 $Y2=1.98
r160 1 41 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=12.775
+ $Y=0.235 $X2=12.9 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 55 58 61 65 71 75 77 82 83 85 87 92 100 108 117 121 126 131 136 142 145 148
+ 151 154 157 160 163 167
c181 167 0 2.58091e-20 $X=15.12 $Y=3.33
r182 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r183 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r184 160 161 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r185 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r186 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r187 151 152 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r188 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r189 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r190 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r191 140 167 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r192 140 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r193 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r194 137 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.375 $Y=3.33
+ $X2=14.21 $Y2=3.33
r195 137 139 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=14.375 $Y=3.33
+ $X2=14.64 $Y2=3.33
r196 136 166 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=14.925 $Y=3.33
+ $X2=15.142 $Y2=3.33
r197 136 139 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=14.925 $Y=3.33
+ $X2=14.64 $Y2=3.33
r198 135 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r199 135 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r200 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r201 132 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.495 $Y=3.33
+ $X2=13.33 $Y2=3.33
r202 132 134 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=13.495 $Y=3.33
+ $X2=13.68 $Y2=3.33
r203 131 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.045 $Y=3.33
+ $X2=14.21 $Y2=3.33
r204 131 134 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=14.045 $Y=3.33
+ $X2=13.68 $Y2=3.33
r205 130 161 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=13.2 $Y2=3.33
r206 130 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r207 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r208 127 157 11.4944 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=11.61 $Y=3.33
+ $X2=11.352 $Y2=3.33
r209 127 129 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=11.61 $Y=3.33
+ $X2=11.76 $Y2=3.33
r210 126 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.165 $Y=3.33
+ $X2=13.33 $Y2=3.33
r211 126 129 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=13.165 $Y=3.33
+ $X2=11.76 $Y2=3.33
r212 125 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r213 125 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r214 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r215 122 154 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=10.41 $Y=3.33
+ $X2=10.31 $Y2=3.33
r216 122 124 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.41 $Y=3.33
+ $X2=10.8 $Y2=3.33
r217 121 157 11.4944 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=11.095 $Y=3.33
+ $X2=11.352 $Y2=3.33
r218 121 124 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.095 $Y=3.33
+ $X2=10.8 $Y2=3.33
r219 120 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r220 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r221 117 154 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=10.21 $Y=3.33
+ $X2=10.31 $Y2=3.33
r222 117 119 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.21 $Y=3.33
+ $X2=9.84 $Y2=3.33
r223 116 120 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r224 115 116 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r225 113 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.02 $Y=3.33
+ $X2=6.855 $Y2=3.33
r226 113 115 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=7.02 $Y=3.33
+ $X2=8.88 $Y2=3.33
r227 112 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r228 112 149 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r229 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r230 109 148 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.7 $Y=3.33
+ $X2=5.53 $Y2=3.33
r231 109 111 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.7 $Y=3.33
+ $X2=6.48 $Y2=3.33
r232 108 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=3.33
+ $X2=6.855 $Y2=3.33
r233 108 111 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.69 $Y=3.33
+ $X2=6.48 $Y2=3.33
r234 107 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r235 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r236 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r237 104 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r238 103 106 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r239 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r240 101 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.52 $Y2=3.33
r241 101 103 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=4.08 $Y2=3.33
r242 100 148 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.36 $Y=3.33
+ $X2=5.53 $Y2=3.33
r243 100 106 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.36 $Y=3.33
+ $X2=5.04 $Y2=3.33
r244 99 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r245 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r246 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r247 96 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r248 95 98 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r249 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r250 93 142 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.91 $Y=3.33
+ $X2=1.765 $Y2=3.33
r251 93 95 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.91 $Y=3.33
+ $X2=2.16 $Y2=3.33
r252 92 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.52 $Y2=3.33
r253 92 98 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.12 $Y2=3.33
r254 90 143 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r255 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r256 87 142 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.62 $Y=3.33
+ $X2=1.765 $Y2=3.33
r257 87 89 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.62 $Y=3.33
+ $X2=0.24 $Y2=3.33
r258 85 116 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=8.88 $Y2=3.33
r259 85 152 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=6.96 $Y2=3.33
r260 82 115 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.005 $Y=3.33
+ $X2=8.88 $Y2=3.33
r261 82 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.005 $Y=3.33
+ $X2=9.17 $Y2=3.33
r262 81 119 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=9.335 $Y=3.33
+ $X2=9.84 $Y2=3.33
r263 81 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.335 $Y=3.33
+ $X2=9.17 $Y2=3.33
r264 77 80 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=15.09 $Y=2.24
+ $X2=15.09 $Y2=2.95
r265 75 166 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=15.09 $Y=3.245
+ $X2=15.142 $Y2=3.33
r266 75 80 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=15.09 $Y=3.245
+ $X2=15.09 $Y2=2.95
r267 71 74 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=14.21 $Y=2.24
+ $X2=14.21 $Y2=2.95
r268 69 163 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.21 $Y=3.245
+ $X2=14.21 $Y2=3.33
r269 69 74 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=14.21 $Y=3.245
+ $X2=14.21 $Y2=2.95
r270 65 68 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=13.33 $Y=2.18
+ $X2=13.33 $Y2=2.95
r271 63 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.33 $Y=3.245
+ $X2=13.33 $Y2=3.33
r272 63 68 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=13.33 $Y=3.245
+ $X2=13.33 $Y2=2.95
r273 61 84 24.3384 $w=1.78e-07 $l=3.95e-07 $layer=LI1_cond $X=11.52 $Y=2.27
+ $X2=11.52 $Y2=2.665
r274 56 157 2.14989 $w=5.15e-07 $l=8.5e-08 $layer=LI1_cond $X=11.352 $Y=3.245
+ $X2=11.352 $Y2=3.33
r275 56 58 6.85132 $w=5.13e-07 $l=2.95e-07 $layer=LI1_cond $X=11.352 $Y=3.245
+ $X2=11.352 $Y2=2.95
r276 55 84 11.3458 $w=5.13e-07 $l=2.57e-07 $layer=LI1_cond $X=11.352 $Y=2.922
+ $X2=11.352 $Y2=2.665
r277 55 58 0.650295 $w=5.13e-07 $l=2.8e-08 $layer=LI1_cond $X=11.352 $Y=2.922
+ $X2=11.352 $Y2=2.95
r278 51 154 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=10.31 $Y=3.245
+ $X2=10.31 $Y2=3.33
r279 51 53 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=10.31 $Y=3.245
+ $X2=10.31 $Y2=2.94
r280 47 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.17 $Y=3.245
+ $X2=9.17 $Y2=3.33
r281 47 49 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=9.17 $Y=3.245
+ $X2=9.17 $Y2=2.94
r282 43 151 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.855 $Y=3.245
+ $X2=6.855 $Y2=3.33
r283 43 45 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=6.855 $Y=3.245
+ $X2=6.855 $Y2=2.72
r284 39 148 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=3.33
r285 39 41 22.2015 $w=3.38e-07 $l=6.55e-07 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=2.59
r286 35 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=3.33
r287 35 37 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=2.77
r288 31 142 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=3.245
+ $X2=1.765 $Y2=3.33
r289 31 33 31.1954 $w=2.88e-07 $l=7.85e-07 $layer=LI1_cond $X=1.765 $Y=3.245
+ $X2=1.765 $Y2=2.46
r290 10 80 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=14.95
+ $Y=1.835 $X2=15.09 $Y2=2.95
r291 10 77 400 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=14.95
+ $Y=1.835 $X2=15.09 $Y2=2.24
r292 9 74 400 $w=1.7e-07 $l=1.19232e-06 $layer=licon1_PDIFF $count=1 $X=14.05
+ $Y=1.835 $X2=14.21 $Y2=2.95
r293 9 71 400 $w=1.7e-07 $l=4.78357e-07 $layer=licon1_PDIFF $count=1 $X=14.05
+ $Y=1.835 $X2=14.21 $Y2=2.24
r294 8 68 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=13.19
+ $Y=1.835 $X2=13.33 $Y2=2.95
r295 8 65 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=13.19
+ $Y=1.835 $X2=13.33 $Y2=2.18
r296 7 61 300 $w=1.7e-07 $l=6.04483e-07 $layer=licon1_PDIFF $count=2 $X=11.12
+ $Y=1.835 $X2=11.525 $Y2=2.27
r297 7 58 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=11.12
+ $Y=1.835 $X2=11.26 $Y2=2.95
r298 6 53 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=10.05
+ $Y=2.665 $X2=10.305 $Y2=2.94
r299 5 49 600 $w=1.7e-07 $l=3.87137e-07 $layer=licon1_PDIFF $count=1 $X=8.9
+ $Y=2.665 $X2=9.17 $Y2=2.94
r300 4 45 600 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.71
+ $Y=1.895 $X2=6.855 $Y2=2.72
r301 3 41 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=2.315 $X2=5.535 $Y2=2.59
r302 2 37 600 $w=1.7e-07 $l=5.56237e-07 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=2.315 $X2=3.52 $Y2=2.77
r303 1 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.605
+ $Y=2.315 $X2=1.745 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%A_372_50# 1 2 3 4 17 19 22 27 30 35 36 37
+ 38 40
r93 36 37 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.905 $Y=0.94
+ $X2=3.075 $Y2=0.94
r94 30 32 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.115 $Y=0.7 $X2=2.115
+ $Y2=0.9
r95 25 38 8.22654 $w=2.5e-07 $l=4.97971e-07 $layer=LI1_cond $X=4.235 $Y=0.805
+ $X2=3.78 $Y2=0.895
r96 25 27 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=4.235 $Y=0.805
+ $X2=4.78 $Y2=0.805
r97 22 40 2.45085 $w=4.17e-07 $l=9e-08 $layer=LI1_cond $X=4.007 $Y=2.295
+ $X2=4.007 $Y2=2.385
r98 21 38 0.695174 $w=4.55e-07 $l=3.00198e-07 $layer=LI1_cond $X=4.007 $Y=1.065
+ $X2=3.78 $Y2=0.895
r99 21 22 32.3335 $w=4.53e-07 $l=1.23e-06 $layer=LI1_cond $X=4.007 $Y=1.065
+ $X2=4.007 $Y2=2.295
r100 19 38 8.22654 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=0.98
+ $X2=3.78 $Y2=0.895
r101 19 37 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.78 $Y=0.98
+ $X2=3.075 $Y2=0.98
r102 18 35 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=2.385
+ $X2=2.535 $Y2=2.385
r103 17 40 4.48849 $w=1.8e-07 $l=2.27e-07 $layer=LI1_cond $X=3.78 $Y=2.385
+ $X2=4.007 $Y2=2.385
r104 17 18 66.5455 $w=1.78e-07 $l=1.08e-06 $layer=LI1_cond $X=3.78 $Y=2.385
+ $X2=2.7 $Y2=2.385
r105 14 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=0.9
+ $X2=2.115 $Y2=0.9
r106 14 36 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.28 $Y=0.9
+ $X2=2.905 $Y2=0.9
r107 4 40 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.88
+ $Y=2.315 $X2=4.02 $Y2=2.46
r108 3 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.395
+ $Y=2.315 $X2=2.535 $Y2=2.46
r109 2 27 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=4.655
+ $Y=0.595 $X2=4.78 $Y2=0.805
r110 1 30 182 $w=1.7e-07 $l=5.6325e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.25 $X2=2.115 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%Q 1 2 3 4 15 17 19 21 22 23 27 29 31 34 38
+ 40 41 44
r57 41 44 21.9616 $w=2.63e-07 $l=5.05e-07 $layer=LI1_cond $X=14.657 $Y=0.925
+ $X2=14.657 $Y2=0.42
r58 37 41 5.21861 $w=2.63e-07 $l=1.2e-07 $layer=LI1_cond $X=14.657 $Y=1.045
+ $X2=14.657 $Y2=0.925
r59 37 38 0.0993765 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=14.657 $Y=1.045
+ $X2=14.657 $Y2=1.135
r60 33 34 22.6056 $w=2.58e-07 $l=5.1e-07 $layer=LI1_cond $X=15.13 $Y=1.225
+ $X2=15.13 $Y2=1.735
r61 32 38 7.18598 $w=1.75e-07 $l=1.35477e-07 $layer=LI1_cond $X=14.79 $Y=1.14
+ $X2=14.657 $Y2=1.135
r62 31 33 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=15 $Y=1.14
+ $X2=15.13 $Y2=1.225
r63 31 32 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=15 $Y=1.14 $X2=14.79
+ $Y2=1.14
r64 30 40 4.27425 $w=2.5e-07 $l=1e-07 $layer=LI1_cond $X=14.745 $Y=1.86
+ $X2=14.645 $Y2=1.86
r65 29 34 6.8199 $w=2.5e-07 $l=1.82071e-07 $layer=LI1_cond $X=15 $Y=1.86
+ $X2=15.13 $Y2=1.735
r66 29 30 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=15 $Y=1.86
+ $X2=14.745 $Y2=1.86
r67 25 40 2.15711 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=14.645 $Y=1.985
+ $X2=14.645 $Y2=1.86
r68 25 27 51.2955 $w=1.98e-07 $l=9.25e-07 $layer=LI1_cond $X=14.645 $Y=1.985
+ $X2=14.645 $Y2=2.91
r69 24 36 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=13.875 $Y=1.86
+ $X2=13.77 $Y2=1.86
r70 23 40 4.27425 $w=2.5e-07 $l=1e-07 $layer=LI1_cond $X=14.545 $Y=1.86
+ $X2=14.645 $Y2=1.86
r71 23 24 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=14.545 $Y=1.86
+ $X2=13.875 $Y2=1.86
r72 21 38 7.18598 $w=1.75e-07 $l=1.32e-07 $layer=LI1_cond $X=14.525 $Y=1.135
+ $X2=14.657 $Y2=1.135
r73 21 22 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=14.525 $Y=1.135
+ $X2=13.855 $Y2=1.135
r74 17 36 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=13.77 $Y=1.985
+ $X2=13.77 $Y2=1.86
r75 17 19 48.8528 $w=2.08e-07 $l=9.25e-07 $layer=LI1_cond $X=13.77 $Y=1.985
+ $X2=13.77 $Y2=2.91
r76 13 22 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=13.76 $Y=1.045
+ $X2=13.855 $Y2=1.135
r77 13 15 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=13.76 $Y=1.045
+ $X2=13.76 $Y2=0.42
r78 4 40 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=1.835 $X2=14.66 $Y2=1.98
r79 4 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=1.835 $X2=14.66 $Y2=2.91
r80 3 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.62
+ $Y=1.835 $X2=13.76 $Y2=1.98
r81 3 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=13.62
+ $Y=1.835 $X2=13.76 $Y2=2.91
r82 2 44 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=14.48
+ $Y=0.235 $X2=14.62 $Y2=0.42
r83 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=13.62
+ $Y=0.235 $X2=13.76 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%VGND 1 2 3 4 5 6 7 8 27 31 33 37 41 45 49
+ 53 55 57 60 61 62 64 69 84 91 96 101 107 110 113 116 119 122 126
c158 126 0 3.56444e-20 $X=15.12 $Y=0
r159 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r160 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r161 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r162 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r163 113 114 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r164 111 114 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=6.48 $Y2=0
r165 110 111 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r166 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r167 105 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r168 105 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=14.16 $Y2=0
r169 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r170 102 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.355 $Y=0
+ $X2=14.19 $Y2=0
r171 102 104 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=14.355 $Y=0
+ $X2=14.64 $Y2=0
r172 101 125 4.42457 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=14.96 $Y=0 $X2=15.16
+ $Y2=0
r173 101 104 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=14.96 $Y=0
+ $X2=14.64 $Y2=0
r174 100 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r175 100 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r176 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r177 97 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.495 $Y=0
+ $X2=13.33 $Y2=0
r178 97 99 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=13.495 $Y=0
+ $X2=13.68 $Y2=0
r179 96 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.025 $Y=0
+ $X2=14.19 $Y2=0
r180 96 99 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=14.025 $Y=0
+ $X2=13.68 $Y2=0
r181 95 120 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r182 95 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r183 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r184 92 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=11.34 $Y2=0
r185 92 94 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=11.76 $Y2=0
r186 91 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.165 $Y=0
+ $X2=13.33 $Y2=0
r187 91 94 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=13.165 $Y=0
+ $X2=11.76 $Y2=0
r188 90 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r189 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r190 87 90 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r191 86 89 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=9.36 $Y=0 $X2=10.8
+ $Y2=0
r192 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r193 84 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.175 $Y=0
+ $X2=11.34 $Y2=0
r194 84 89 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.175 $Y=0
+ $X2=10.8 $Y2=0
r195 83 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r196 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r197 80 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r198 79 82 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=8.88
+ $Y2=0
r199 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r200 77 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=0 $X2=6.6
+ $Y2=0
r201 77 79 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.765 $Y=0
+ $X2=6.96 $Y2=0
r202 76 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r203 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r204 73 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r205 73 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r206 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r207 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r208 70 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0
+ $X2=0.69 $Y2=0
r209 70 72 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r210 69 110 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.355 $Y=0
+ $X2=3.485 $Y2=0
r211 69 75 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=0
+ $X2=3.12 $Y2=0
r212 67 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r213 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r214 64 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.69 $Y2=0
r215 64 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.24 $Y2=0
r216 62 83 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=7.68 $Y=0 $X2=8.88
+ $Y2=0
r217 62 80 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.68 $Y=0 $X2=6.96
+ $Y2=0
r218 60 82 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=8.955 $Y=0 $X2=8.88
+ $Y2=0
r219 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.955 $Y=0 $X2=9.12
+ $Y2=0
r220 59 86 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=9.285 $Y=0 $X2=9.36
+ $Y2=0
r221 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.285 $Y=0 $X2=9.12
+ $Y2=0
r222 55 125 3.05295 $w=2.95e-07 $l=1.08305e-07 $layer=LI1_cond $X=15.107
+ $Y=0.085 $X2=15.16 $Y2=0
r223 55 57 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=15.107 $Y=0.085
+ $X2=15.107 $Y2=0.38
r224 51 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.19 $Y=0.085
+ $X2=14.19 $Y2=0
r225 51 53 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=14.19 $Y=0.085
+ $X2=14.19 $Y2=0.36
r226 47 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.33 $Y=0.085
+ $X2=13.33 $Y2=0
r227 47 49 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=13.33 $Y=0.085
+ $X2=13.33 $Y2=0.535
r228 43 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.34 $Y=0.085
+ $X2=11.34 $Y2=0
r229 43 45 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=11.34 $Y=0.085
+ $X2=11.34 $Y2=0.36
r230 39 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.12 $Y=0.085
+ $X2=9.12 $Y2=0
r231 39 41 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=9.12 $Y=0.085
+ $X2=9.12 $Y2=0.8
r232 35 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.6 $Y=0.085
+ $X2=6.6 $Y2=0
r233 35 37 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6.6 $Y=0.085
+ $X2=6.6 $Y2=0.49
r234 34 110 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.615 $Y=0
+ $X2=3.485 $Y2=0
r235 33 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=0 $X2=6.6
+ $Y2=0
r236 33 34 183.979 $w=1.68e-07 $l=2.82e-06 $layer=LI1_cond $X=6.435 $Y=0
+ $X2=3.615 $Y2=0
r237 29 110 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=0.085
+ $X2=3.485 $Y2=0
r238 29 31 21.0542 $w=2.58e-07 $l=4.75e-07 $layer=LI1_cond $X=3.485 $Y=0.085
+ $X2=3.485 $Y2=0.56
r239 25 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r240 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.525
r241 8 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.95
+ $Y=0.235 $X2=15.09 $Y2=0.38
r242 7 53 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=14.05
+ $Y=0.235 $X2=14.19 $Y2=0.36
r243 6 49 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=13.19
+ $Y=0.235 $X2=13.33 $Y2=0.535
r244 5 45 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=11.12
+ $Y=0.345 $X2=11.34 $Y2=0.36
r245 4 41 182 $w=1.7e-07 $l=3.3234e-07 $layer=licon1_NDIFF $count=1 $X=8.885
+ $Y=0.565 $X2=9.12 $Y2=0.8
r246 3 37 91 $w=1.7e-07 $l=2.82666e-07 $layer=licon1_NDIFF $count=2 $X=6.365
+ $Y=0.595 $X2=6.6 $Y2=0.49
r247 2 31 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.31
+ $Y=0.405 $X2=3.45 $Y2=0.56
r248 1 27 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.37 $X2=0.69 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_4%noxref_24 1 2 7 9 14
c35 7 0 1.44625e-19 $X=2.855 $Y=0.34
r36 14 17 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.02 $Y=0.34
+ $X2=3.02 $Y2=0.53
r37 9 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.21 $Y=0.34 $X2=1.21
+ $Y2=0.46
r38 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.34 $X2=1.21
+ $Y2=0.34
r39 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=0.34
+ $X2=3.02 $Y2=0.34
r40 7 8 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=2.855 $Y=0.34
+ $X2=1.375 $Y2=0.34
r41 2 17 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.88
+ $Y=0.405 $X2=3.02 $Y2=0.53
r42 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.25 $X2=1.21 $Y2=0.46
.ends

