* File: sky130_fd_sc_lp__dlclkp_1.pxi.spice
* Created: Fri Aug 28 10:24:51 2020
* 
x_PM_SKY130_FD_SC_LP__DLCLKP_1%A_80_269# N_A_80_269#_M1016_d N_A_80_269#_M1000_d
+ N_A_80_269#_M1019_g N_A_80_269#_M1008_g N_A_80_269#_c_156_n
+ N_A_80_269#_c_163_p N_A_80_269#_c_182_p N_A_80_269#_c_150_n
+ N_A_80_269#_c_221_p N_A_80_269#_c_184_p N_A_80_269#_c_151_n
+ N_A_80_269#_c_152_n N_A_80_269#_c_153_n N_A_80_269#_c_154_n
+ PM_SKY130_FD_SC_LP__DLCLKP_1%A_80_269#
x_PM_SKY130_FD_SC_LP__DLCLKP_1%GATE N_GATE_M1018_g N_GATE_M1002_g GATE
+ N_GATE_c_244_n PM_SKY130_FD_SC_LP__DLCLKP_1%GATE
x_PM_SKY130_FD_SC_LP__DLCLKP_1%A_315_382# N_A_315_382#_M1012_d
+ N_A_315_382#_M1003_d N_A_315_382#_M1000_g N_A_315_382#_M1010_g
+ N_A_315_382#_c_290_n N_A_315_382#_c_298_n N_A_315_382#_c_291_n
+ N_A_315_382#_c_299_n N_A_315_382#_c_292_n N_A_315_382#_c_301_n
+ N_A_315_382#_c_302_n N_A_315_382#_c_293_n N_A_315_382#_c_294_n
+ N_A_315_382#_c_295_n N_A_315_382#_c_303_n
+ PM_SKY130_FD_SC_LP__DLCLKP_1%A_315_382#
x_PM_SKY130_FD_SC_LP__DLCLKP_1%A_27_367# N_A_27_367#_M1008_s N_A_27_367#_M1019_s
+ N_A_27_367#_M1001_g N_A_27_367#_M1004_g N_A_27_367#_c_435_n
+ N_A_27_367#_c_436_n N_A_27_367#_M1005_g N_A_27_367#_M1017_g
+ N_A_27_367#_c_420_n N_A_27_367#_c_421_n N_A_27_367#_c_439_n
+ N_A_27_367#_c_440_n N_A_27_367#_c_422_n N_A_27_367#_c_441_n
+ N_A_27_367#_c_442_n N_A_27_367#_c_443_n N_A_27_367#_c_475_n
+ N_A_27_367#_c_423_n N_A_27_367#_c_424_n N_A_27_367#_c_444_n
+ N_A_27_367#_c_445_n N_A_27_367#_c_446_n N_A_27_367#_c_425_n
+ N_A_27_367#_c_447_n N_A_27_367#_c_448_n N_A_27_367#_c_426_n
+ N_A_27_367#_c_427_n N_A_27_367#_c_428_n N_A_27_367#_c_429_n
+ N_A_27_367#_c_430_n N_A_27_367#_c_450_n N_A_27_367#_c_431_n
+ N_A_27_367#_c_432_n N_A_27_367#_c_451_n N_A_27_367#_c_452_n
+ N_A_27_367#_c_453_n N_A_27_367#_c_433_n PM_SKY130_FD_SC_LP__DLCLKP_1%A_27_367#
x_PM_SKY130_FD_SC_LP__DLCLKP_1%A_321_55# N_A_321_55#_M1013_s N_A_321_55#_M1011_s
+ N_A_321_55#_M1016_g N_A_321_55#_c_650_n N_A_321_55#_c_651_n
+ N_A_321_55#_M1009_g N_A_321_55#_M1012_g N_A_321_55#_c_664_n
+ N_A_321_55#_M1003_g N_A_321_55#_c_653_n N_A_321_55#_c_654_n
+ N_A_321_55#_c_655_n N_A_321_55#_c_656_n N_A_321_55#_c_699_n
+ N_A_321_55#_c_657_n N_A_321_55#_c_733_n N_A_321_55#_c_658_n
+ N_A_321_55#_c_705_n N_A_321_55#_c_659_n N_A_321_55#_c_660_n
+ PM_SKY130_FD_SC_LP__DLCLKP_1%A_321_55#
x_PM_SKY130_FD_SC_LP__DLCLKP_1%CLK N_CLK_c_756_n N_CLK_M1013_g N_CLK_c_765_n
+ N_CLK_M1011_g N_CLK_c_758_n N_CLK_c_759_n N_CLK_M1007_g N_CLK_c_768_n
+ N_CLK_M1006_g N_CLK_c_761_n CLK N_CLK_c_762_n N_CLK_c_763_n
+ PM_SKY130_FD_SC_LP__DLCLKP_1%CLK
x_PM_SKY130_FD_SC_LP__DLCLKP_1%A_1046_367# N_A_1046_367#_M1005_d
+ N_A_1046_367#_M1006_d N_A_1046_367#_M1014_g N_A_1046_367#_M1015_g
+ N_A_1046_367#_c_839_n N_A_1046_367#_c_832_n N_A_1046_367#_c_833_n
+ N_A_1046_367#_c_834_n N_A_1046_367#_c_835_n N_A_1046_367#_c_836_n
+ N_A_1046_367#_c_837_n PM_SKY130_FD_SC_LP__DLCLKP_1%A_1046_367#
x_PM_SKY130_FD_SC_LP__DLCLKP_1%VPWR N_VPWR_M1019_d N_VPWR_M1001_d N_VPWR_M1011_d
+ N_VPWR_M1017_d N_VPWR_c_890_n N_VPWR_c_891_n N_VPWR_c_892_n N_VPWR_c_893_n
+ N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n N_VPWR_c_897_n VPWR
+ N_VPWR_c_898_n N_VPWR_c_899_n N_VPWR_c_900_n N_VPWR_c_889_n N_VPWR_c_902_n
+ N_VPWR_c_903_n PM_SKY130_FD_SC_LP__DLCLKP_1%VPWR
x_PM_SKY130_FD_SC_LP__DLCLKP_1%GCLK N_GCLK_M1014_d N_GCLK_M1015_d GCLK GCLK GCLK
+ GCLK GCLK N_GCLK_c_982_n PM_SKY130_FD_SC_LP__DLCLKP_1%GCLK
x_PM_SKY130_FD_SC_LP__DLCLKP_1%VGND N_VGND_M1008_d N_VGND_M1004_d N_VGND_M1013_d
+ N_VGND_M1014_s N_VGND_c_992_n N_VGND_c_993_n N_VGND_c_994_n N_VGND_c_995_n
+ N_VGND_c_996_n N_VGND_c_997_n N_VGND_c_998_n N_VGND_c_999_n VGND
+ N_VGND_c_1000_n N_VGND_c_1001_n N_VGND_c_1002_n N_VGND_c_1003_n
+ N_VGND_c_1004_n N_VGND_c_1005_n PM_SKY130_FD_SC_LP__DLCLKP_1%VGND
cc_1 VNB N_A_80_269#_M1008_g 0.0325856f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.655
cc_2 VNB N_A_80_269#_c_150_n 0.00576458f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=1.56
cc_3 VNB N_A_80_269#_c_151_n 0.0013153f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.51
cc_4 VNB N_A_80_269#_c_152_n 0.0334984f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.51
cc_5 VNB N_A_80_269#_c_153_n 0.00468376f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.65
cc_6 VNB N_A_80_269#_c_154_n 0.0063298f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=1.65
cc_7 VNB N_GATE_M1018_g 0.0100018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_GATE_M1002_g 0.0263989f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.675
cc_9 VNB GATE 0.00560014f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_10 VNB N_GATE_c_244_n 0.0297832f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.655
cc_11 VNB N_A_315_382#_M1010_g 0.0176552f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.655
cc_12 VNB N_A_315_382#_c_290_n 0.00858725f $X=-0.19 $Y=-0.245 $X2=0.795
+ $Y2=1.645
cc_13 VNB N_A_315_382#_c_291_n 0.0206201f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.61
cc_14 VNB N_A_315_382#_c_292_n 0.00758956f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=1.56
cc_15 VNB N_A_315_382#_c_293_n 0.00244027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_315_382#_c_294_n 0.0312179f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.65
cc_17 VNB N_A_315_382#_c_295_n 0.0129347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_367#_M1005_g 0.0234292f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.485
cc_19 VNB N_A_27_367#_M1017_g 0.0171376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_367#_c_420_n 0.0274647f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=0.695
cc_21 VNB N_A_27_367#_c_421_n 0.0299901f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.51
cc_22 VNB N_A_27_367#_c_422_n 0.0037121f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.65
cc_23 VNB N_A_27_367#_c_423_n 0.00876632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_367#_c_424_n 0.00234964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_367#_c_425_n 0.00140861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_367#_c_426_n 0.00253085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_367#_c_427_n 0.00346183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_367#_c_428_n 0.0108457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_367#_c_429_n 0.0400353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_367#_c_430_n 0.0162813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_367#_c_431_n 0.00488664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_367#_c_432_n 0.0324184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_367#_c_433_n 0.0169662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_321_55#_M1016_g 0.0397659f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_35 VNB N_A_321_55#_c_650_n 0.0123426f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.345
cc_36 VNB N_A_321_55#_c_651_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.655
cc_37 VNB N_A_321_55#_M1012_g 0.0313385f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.61
cc_38 VNB N_A_321_55#_c_653_n 0.00493328f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=0.695
cc_39 VNB N_A_321_55#_c_654_n 0.035113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_321_55#_c_655_n 0.0345474f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.51
cc_41 VNB N_A_321_55#_c_656_n 0.00797477f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.51
cc_42 VNB N_A_321_55#_c_657_n 0.00292844f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.65
cc_43 VNB N_A_321_55#_c_658_n 0.0174291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_321_55#_c_659_n 0.00950456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_321_55#_c_660_n 0.0172832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_CLK_c_756_n 0.0101314f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=0.405
cc_47 VNB N_CLK_M1013_g 0.0310614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_CLK_c_758_n 0.00583158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_CLK_c_759_n 0.0109921f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.345
cc_50 VNB N_CLK_M1007_g 0.0532229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_CLK_c_761_n 0.010805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_CLK_c_762_n 0.0027696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_CLK_c_763_n 0.0216444f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.51
cc_54 VNB N_A_1046_367#_M1014_g 0.0298984f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=2.465
cc_55 VNB N_A_1046_367#_c_832_n 0.00439781f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=2.61
cc_56 VNB N_A_1046_367#_c_833_n 0.00256254f $X=-0.19 $Y=-0.245 $X2=1.905
+ $Y2=2.61
cc_57 VNB N_A_1046_367#_c_834_n 0.00804482f $X=-0.19 $Y=-0.245 $X2=1.905
+ $Y2=2.61
cc_58 VNB N_A_1046_367#_c_835_n 0.00209518f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=1.56
cc_59 VNB N_A_1046_367#_c_836_n 0.0059763f $X=-0.19 $Y=-0.245 $X2=1.895
+ $Y2=0.695
cc_60 VNB N_A_1046_367#_c_837_n 0.031932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VPWR_c_889_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_GCLK_c_982_n 0.0608596f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.485
cc_63 VNB N_VGND_c_992_n 0.00761256f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.645
cc_64 VNB N_VGND_c_993_n 0.010524f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.61
cc_65 VNB N_VGND_c_994_n 0.0191354f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=0.795
cc_66 VNB N_VGND_c_995_n 0.00729673f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=0.7
cc_67 VNB N_VGND_c_996_n 0.0212313f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.51
cc_68 VNB N_VGND_c_997_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.51
cc_69 VNB N_VGND_c_998_n 0.0415946f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.645
cc_70 VNB N_VGND_c_999_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1000_n 0.0387797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1001_n 0.0318304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1002_n 0.0153759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1003_n 0.389689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1004_n 0.00631736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1005_n 0.00510306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VPB N_A_80_269#_M1019_g 0.0256352f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_78 VPB N_A_80_269#_c_156_n 0.00554581f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=2.485
cc_79 VPB N_A_80_269#_c_151_n 0.00238808f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.51
cc_80 VPB N_A_80_269#_c_152_n 0.00863729f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.51
cc_81 VPB N_A_80_269#_c_153_n 0.00589237f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=1.65
cc_82 VPB N_A_80_269#_c_154_n 0.00522923f $X=-0.19 $Y=1.655 $X2=1.67 $Y2=1.65
cc_83 VPB N_GATE_M1018_g 0.0566578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_315_382#_M1000_g 0.0216934f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_85 VPB N_A_315_382#_c_290_n 0.00443108f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=1.645
cc_86 VPB N_A_315_382#_c_298_n 0.0172888f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=1.74
cc_87 VPB N_A_315_382#_c_299_n 0.00770161f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=2.61
cc_88 VPB N_A_315_382#_c_292_n 7.17385e-19 $X=-0.19 $Y=1.655 $X2=1.67 $Y2=1.56
cc_89 VPB N_A_315_382#_c_301_n 0.0309143f $X=-0.19 $Y=1.655 $X2=1.895 $Y2=0.7
cc_90 VPB N_A_315_382#_c_302_n 0.00433271f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.51
cc_91 VPB N_A_315_382#_c_303_n 0.007441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_27_367#_M1001_g 0.022037f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_93 VPB N_A_27_367#_c_435_n 0.0663742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_27_367#_c_436_n 0.0124856f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=1.645
cc_95 VPB N_A_27_367#_M1017_g 0.0232346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_27_367#_c_421_n 0.0115478f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.51
cc_97 VPB N_A_27_367#_c_439_n 0.0391498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_27_367#_c_440_n 0.0113053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_27_367#_c_441_n 0.00654649f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.51
cc_100 VPB N_A_27_367#_c_442_n 0.0104884f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.345
cc_101 VPB N_A_27_367#_c_443_n 0.00156179f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.675
cc_102 VPB N_A_27_367#_c_444_n 0.00130526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_27_367#_c_445_n 9.50589e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_27_367#_c_446_n 0.00279106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_27_367#_c_447_n 0.00248192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_27_367#_c_448_n 0.0206287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_27_367#_c_426_n 7.01374e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_27_367#_c_450_n 0.00717518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_27_367#_c_451_n 0.00171674f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_27_367#_c_452_n 0.00414843f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_27_367#_c_453_n 0.0629982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_321_55#_c_650_n 0.00948125f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.345
cc_113 VPB N_A_321_55#_c_651_n 0.00245614f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.655
cc_114 VPB N_A_321_55#_M1009_g 0.0463282f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=1.645
cc_115 VPB N_A_321_55#_c_664_n 0.0220346f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=2.61
cc_116 VPB N_A_321_55#_c_653_n 0.00778966f $X=-0.19 $Y=1.655 $X2=1.755 $Y2=0.695
cc_117 VPB N_A_321_55#_c_655_n 0.0335994f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.51
cc_118 VPB N_A_321_55#_c_656_n 0.0169471f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.51
cc_119 VPB N_A_321_55#_c_659_n 0.00887013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_CLK_c_756_n 0.0103311f $X=-0.19 $Y=1.655 $X2=1.755 $Y2=0.405
cc_121 VPB N_CLK_c_765_n 0.0207336f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.675
cc_122 VPB N_CLK_c_758_n 0.00797943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_CLK_c_759_n 0.0105625f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.345
cc_124 VPB N_CLK_c_768_n 0.0180789f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=1.645
cc_125 VPB N_CLK_c_761_n 0.00960089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_CLK_c_762_n 0.00534587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_CLK_c_763_n 0.014517f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.51
cc_128 VPB N_A_1046_367#_M1015_g 0.0258644f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.655
cc_129 VPB N_A_1046_367#_c_839_n 0.00725272f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=1.74
cc_130 VPB N_A_1046_367#_c_832_n 0.00411544f $X=-0.19 $Y=1.655 $X2=1.485
+ $Y2=2.61
cc_131 VPB N_A_1046_367#_c_835_n 0.00210868f $X=-0.19 $Y=1.655 $X2=1.67 $Y2=1.56
cc_132 VPB N_A_1046_367#_c_837_n 0.00718539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_890_n 0.00489893f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=1.645
cc_134 VPB N_VPWR_c_891_n 0.0037814f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.61
cc_135 VPB N_VPWR_c_892_n 0.014738f $X=-0.19 $Y=1.655 $X2=1.67 $Y2=0.795
cc_136 VPB N_VPWR_c_893_n 0.021488f $X=-0.19 $Y=1.655 $X2=1.895 $Y2=0.7
cc_137 VPB N_VPWR_c_894_n 0.0458341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_895_n 0.00479588f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.645
cc_139 VPB N_VPWR_c_896_n 0.0427677f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=1.65
cc_140 VPB N_VPWR_c_897_n 0.00631189f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=1.65
cc_141 VPB N_VPWR_c_898_n 0.0181824f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.51
cc_142 VPB N_VPWR_c_899_n 0.0190152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_900_n 0.0153759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_889_n 0.0793362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_902_n 0.00382106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_903_n 0.00953241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_GCLK_c_982_n 0.056799f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=2.485
cc_148 N_A_80_269#_M1019_g N_GATE_M1018_g 0.0136317f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_80_269#_c_156_n N_GATE_M1018_g 0.0198254f $X=1.4 $Y=2.485 $X2=0 $Y2=0
cc_150 N_A_80_269#_c_163_p N_GATE_M1018_g 0.00605615f $X=1.485 $Y=2.61 $X2=0
+ $Y2=0
cc_151 N_A_80_269#_c_150_n N_GATE_M1018_g 0.00190422f $X=1.67 $Y=1.56 $X2=0
+ $Y2=0
cc_152 N_A_80_269#_c_151_n N_GATE_M1018_g 6.92594e-19 $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_153 N_A_80_269#_c_152_n N_GATE_M1018_g 0.00615769f $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_154 N_A_80_269#_c_153_n N_GATE_M1018_g 0.010081f $X=1.315 $Y=1.65 $X2=0 $Y2=0
cc_155 N_A_80_269#_c_154_n N_GATE_M1018_g 0.00447524f $X=1.67 $Y=1.65 $X2=0
+ $Y2=0
cc_156 N_A_80_269#_M1008_g N_GATE_M1002_g 0.0144066f $X=0.63 $Y=0.655 $X2=0
+ $Y2=0
cc_157 N_A_80_269#_c_150_n N_GATE_M1002_g 0.00381858f $X=1.67 $Y=1.56 $X2=0
+ $Y2=0
cc_158 N_A_80_269#_M1008_g GATE 0.00190077f $X=0.63 $Y=0.655 $X2=0 $Y2=0
cc_159 N_A_80_269#_c_150_n GATE 0.0185761f $X=1.67 $Y=1.56 $X2=0 $Y2=0
cc_160 N_A_80_269#_c_151_n GATE 0.00337269f $X=0.63 $Y=1.51 $X2=0 $Y2=0
cc_161 N_A_80_269#_c_152_n GATE 2.98167e-19 $X=0.63 $Y=1.51 $X2=0 $Y2=0
cc_162 N_A_80_269#_c_153_n GATE 0.0320474f $X=1.315 $Y=1.65 $X2=0 $Y2=0
cc_163 N_A_80_269#_M1008_g N_GATE_c_244_n 0.00674614f $X=0.63 $Y=0.655 $X2=0
+ $Y2=0
cc_164 N_A_80_269#_c_150_n N_GATE_c_244_n 0.00204856f $X=1.67 $Y=1.56 $X2=0
+ $Y2=0
cc_165 N_A_80_269#_c_151_n N_GATE_c_244_n 5.35311e-19 $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_166 N_A_80_269#_c_152_n N_GATE_c_244_n 0.00576524f $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_167 N_A_80_269#_c_153_n N_GATE_c_244_n 0.00365313f $X=1.315 $Y=1.65 $X2=0
+ $Y2=0
cc_168 N_A_80_269#_c_154_n N_GATE_c_244_n 8.59174e-19 $X=1.67 $Y=1.65 $X2=0
+ $Y2=0
cc_169 N_A_80_269#_c_182_p N_A_315_382#_M1000_g 0.0124423f $X=1.905 $Y=2.61
+ $X2=0 $Y2=0
cc_170 N_A_80_269#_c_150_n N_A_315_382#_M1010_g 8.83118e-19 $X=1.67 $Y=1.56
+ $X2=0 $Y2=0
cc_171 N_A_80_269#_c_184_p N_A_315_382#_M1010_g 0.00364692f $X=1.895 $Y=0.7
+ $X2=0 $Y2=0
cc_172 N_A_80_269#_c_156_n N_A_315_382#_c_290_n 0.00663451f $X=1.4 $Y=2.485
+ $X2=0 $Y2=0
cc_173 N_A_80_269#_c_150_n N_A_315_382#_c_290_n 0.0187142f $X=1.67 $Y=1.56 $X2=0
+ $Y2=0
cc_174 N_A_80_269#_c_154_n N_A_315_382#_c_290_n 0.0139798f $X=1.67 $Y=1.65 $X2=0
+ $Y2=0
cc_175 N_A_80_269#_c_156_n N_A_315_382#_c_301_n 0.00742776f $X=1.4 $Y=2.485
+ $X2=0 $Y2=0
cc_176 N_A_80_269#_c_182_p N_A_315_382#_c_301_n 0.00371519f $X=1.905 $Y=2.61
+ $X2=0 $Y2=0
cc_177 N_A_80_269#_c_154_n N_A_315_382#_c_301_n 0.00292163f $X=1.67 $Y=1.65
+ $X2=0 $Y2=0
cc_178 N_A_80_269#_c_156_n N_A_315_382#_c_302_n 0.0257833f $X=1.4 $Y=2.485 $X2=0
+ $Y2=0
cc_179 N_A_80_269#_c_182_p N_A_315_382#_c_302_n 0.0222937f $X=1.905 $Y=2.61
+ $X2=0 $Y2=0
cc_180 N_A_80_269#_c_154_n N_A_315_382#_c_302_n 0.00754852f $X=1.67 $Y=1.65
+ $X2=0 $Y2=0
cc_181 N_A_80_269#_c_150_n N_A_315_382#_c_293_n 0.0250402f $X=1.67 $Y=1.56 $X2=0
+ $Y2=0
cc_182 N_A_80_269#_c_184_p N_A_315_382#_c_293_n 0.00803622f $X=1.895 $Y=0.7
+ $X2=0 $Y2=0
cc_183 N_A_80_269#_c_150_n N_A_315_382#_c_294_n 3.80323e-19 $X=1.67 $Y=1.56
+ $X2=0 $Y2=0
cc_184 N_A_80_269#_c_184_p N_A_315_382#_c_294_n 0.00144548f $X=1.895 $Y=0.7
+ $X2=0 $Y2=0
cc_185 N_A_80_269#_M1008_g N_A_27_367#_c_420_n 0.0102901f $X=0.63 $Y=0.655 $X2=0
+ $Y2=0
cc_186 N_A_80_269#_M1008_g N_A_27_367#_c_421_n 0.00664999f $X=0.63 $Y=0.655
+ $X2=0 $Y2=0
cc_187 N_A_80_269#_c_151_n N_A_27_367#_c_421_n 0.0294303f $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_188 N_A_80_269#_c_152_n N_A_27_367#_c_421_n 0.0147395f $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_189 N_A_80_269#_M1019_g N_A_27_367#_c_439_n 0.0157153f $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_190 N_A_80_269#_M1019_g N_A_27_367#_c_440_n 0.0155848f $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_191 N_A_80_269#_c_156_n N_A_27_367#_c_440_n 0.0137143f $X=1.4 $Y=2.485 $X2=0
+ $Y2=0
cc_192 N_A_80_269#_c_151_n N_A_27_367#_c_440_n 0.0182886f $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_193 N_A_80_269#_c_152_n N_A_27_367#_c_440_n 0.00135631f $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_194 N_A_80_269#_c_153_n N_A_27_367#_c_440_n 0.027848f $X=1.315 $Y=1.65 $X2=0
+ $Y2=0
cc_195 N_A_80_269#_M1008_g N_A_27_367#_c_422_n 0.0105073f $X=0.63 $Y=0.655 $X2=0
+ $Y2=0
cc_196 N_A_80_269#_c_150_n N_A_27_367#_c_422_n 0.0138463f $X=1.67 $Y=1.56 $X2=0
+ $Y2=0
cc_197 N_A_80_269#_c_151_n N_A_27_367#_c_422_n 0.00757838f $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_198 N_A_80_269#_c_152_n N_A_27_367#_c_422_n 3.63634e-19 $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_199 N_A_80_269#_c_153_n N_A_27_367#_c_422_n 0.00558777f $X=1.315 $Y=1.65
+ $X2=0 $Y2=0
cc_200 N_A_80_269#_M1019_g N_A_27_367#_c_441_n 0.00217798f $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_201 N_A_80_269#_c_156_n N_A_27_367#_c_441_n 0.0294959f $X=1.4 $Y=2.485 $X2=0
+ $Y2=0
cc_202 N_A_80_269#_c_163_p N_A_27_367#_c_441_n 0.0196495f $X=1.485 $Y=2.61 $X2=0
+ $Y2=0
cc_203 N_A_80_269#_M1000_d N_A_27_367#_c_442_n 0.00234513f $X=1.725 $Y=2.4 $X2=0
+ $Y2=0
cc_204 N_A_80_269#_c_163_p N_A_27_367#_c_442_n 0.00831808f $X=1.485 $Y=2.61
+ $X2=0 $Y2=0
cc_205 N_A_80_269#_c_182_p N_A_27_367#_c_442_n 0.0320264f $X=1.905 $Y=2.61 $X2=0
+ $Y2=0
cc_206 N_A_80_269#_M1008_g N_A_27_367#_c_475_n 6.86494e-19 $X=0.63 $Y=0.655
+ $X2=0 $Y2=0
cc_207 N_A_80_269#_M1016_d N_A_27_367#_c_423_n 0.001755f $X=1.755 $Y=0.405 $X2=0
+ $Y2=0
cc_208 N_A_80_269#_c_221_p N_A_27_367#_c_423_n 0.0106506f $X=1.755 $Y=0.695
+ $X2=0 $Y2=0
cc_209 N_A_80_269#_c_184_p N_A_27_367#_c_423_n 0.0130599f $X=1.895 $Y=0.7 $X2=0
+ $Y2=0
cc_210 N_A_80_269#_M1008_g N_A_27_367#_c_430_n 0.00380634f $X=0.63 $Y=0.655
+ $X2=0 $Y2=0
cc_211 N_A_80_269#_c_151_n N_A_27_367#_c_430_n 0.00268438f $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_212 N_A_80_269#_c_152_n N_A_27_367#_c_430_n 0.00618141f $X=0.63 $Y=1.51 $X2=0
+ $Y2=0
cc_213 N_A_80_269#_M1019_g N_A_27_367#_c_450_n 0.00156562f $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_214 N_A_80_269#_c_150_n N_A_321_55#_M1016_g 0.0153816f $X=1.67 $Y=1.56 $X2=0
+ $Y2=0
cc_215 N_A_80_269#_c_221_p N_A_321_55#_M1016_g 0.00529199f $X=1.755 $Y=0.695
+ $X2=0 $Y2=0
cc_216 N_A_80_269#_c_150_n N_A_321_55#_c_651_n 0.00209583f $X=1.67 $Y=1.56 $X2=0
+ $Y2=0
cc_217 N_A_80_269#_c_154_n N_A_321_55#_c_651_n 0.00581464f $X=1.67 $Y=1.65 $X2=0
+ $Y2=0
cc_218 N_A_80_269#_c_156_n N_A_321_55#_M1009_g 3.92747e-19 $X=1.4 $Y=2.485 $X2=0
+ $Y2=0
cc_219 N_A_80_269#_M1019_g N_VPWR_c_890_n 0.00507177f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_220 N_A_80_269#_M1019_g N_VPWR_c_898_n 0.0054895f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_221 N_A_80_269#_M1019_g N_VPWR_c_889_n 0.011678f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_222 N_A_80_269#_c_156_n A_273_480# 9.33292e-19 $X=1.4 $Y=2.485 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_80_269#_c_163_p A_273_480# 6.55502e-19 $X=1.485 $Y=2.61 $X2=-0.19
+ $Y2=-0.245
cc_224 N_A_80_269#_c_182_p A_273_480# 0.00160818f $X=1.905 $Y=2.61 $X2=-0.19
+ $Y2=-0.245
cc_225 N_A_80_269#_M1008_g N_VGND_c_992_n 0.00827162f $X=0.63 $Y=0.655 $X2=0
+ $Y2=0
cc_226 N_A_80_269#_M1008_g N_VGND_c_996_n 0.0055654f $X=0.63 $Y=0.655 $X2=0
+ $Y2=0
cc_227 N_A_80_269#_M1008_g N_VGND_c_1003_n 0.00855039f $X=0.63 $Y=0.655 $X2=0
+ $Y2=0
cc_228 N_GATE_M1018_g N_A_315_382#_c_290_n 0.00103642f $X=1.29 $Y=2.72 $X2=0
+ $Y2=0
cc_229 N_GATE_M1018_g N_A_315_382#_c_301_n 0.0787562f $X=1.29 $Y=2.72 $X2=0
+ $Y2=0
cc_230 N_GATE_M1018_g N_A_315_382#_c_302_n 2.88086e-19 $X=1.29 $Y=2.72 $X2=0
+ $Y2=0
cc_231 N_GATE_M1002_g N_A_27_367#_c_420_n 5.45827e-19 $X=1.32 $Y=0.615 $X2=0
+ $Y2=0
cc_232 GATE N_A_27_367#_c_421_n 0.00629024f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_233 N_GATE_M1018_g N_A_27_367#_c_440_n 0.00204747f $X=1.29 $Y=2.72 $X2=0
+ $Y2=0
cc_234 N_GATE_M1002_g N_A_27_367#_c_422_n 0.00799386f $X=1.32 $Y=0.615 $X2=0
+ $Y2=0
cc_235 GATE N_A_27_367#_c_422_n 0.0334567f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_236 N_GATE_c_244_n N_A_27_367#_c_422_n 0.00430025f $X=1.23 $Y=1.295 $X2=0
+ $Y2=0
cc_237 N_GATE_M1018_g N_A_27_367#_c_441_n 0.0119725f $X=1.29 $Y=2.72 $X2=0 $Y2=0
cc_238 N_GATE_M1018_g N_A_27_367#_c_442_n 0.0126857f $X=1.29 $Y=2.72 $X2=0 $Y2=0
cc_239 N_GATE_M1002_g N_A_27_367#_c_475_n 0.00978188f $X=1.32 $Y=0.615 $X2=0
+ $Y2=0
cc_240 N_GATE_M1002_g N_A_27_367#_c_424_n 0.00560041f $X=1.32 $Y=0.615 $X2=0
+ $Y2=0
cc_241 N_GATE_M1002_g N_A_27_367#_c_430_n 4.4685e-19 $X=1.32 $Y=0.615 $X2=0
+ $Y2=0
cc_242 N_GATE_M1018_g N_A_321_55#_M1016_g 0.0118644f $X=1.29 $Y=2.72 $X2=0 $Y2=0
cc_243 N_GATE_M1002_g N_A_321_55#_M1016_g 0.0744462f $X=1.32 $Y=0.615 $X2=0
+ $Y2=0
cc_244 GATE N_A_321_55#_M1016_g 7.55897e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_245 N_GATE_M1018_g N_VPWR_c_890_n 0.00259619f $X=1.29 $Y=2.72 $X2=0 $Y2=0
cc_246 N_GATE_M1018_g N_VPWR_c_894_n 0.00322875f $X=1.29 $Y=2.72 $X2=0 $Y2=0
cc_247 N_GATE_M1018_g N_VPWR_c_889_n 0.00516743f $X=1.29 $Y=2.72 $X2=0 $Y2=0
cc_248 N_GATE_M1002_g N_VGND_c_992_n 0.00252952f $X=1.32 $Y=0.615 $X2=0 $Y2=0
cc_249 N_GATE_M1002_g N_VGND_c_998_n 9.14566e-19 $X=1.32 $Y=0.615 $X2=0 $Y2=0
cc_250 N_A_315_382#_c_298_n N_A_27_367#_M1001_g 0.0013307f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_251 N_A_315_382#_M1000_g N_A_27_367#_c_442_n 0.010671f $X=1.65 $Y=2.72 $X2=0
+ $Y2=0
cc_252 N_A_315_382#_c_302_n N_A_27_367#_c_442_n 7.64704e-19 $X=2.095 $Y=2.075
+ $X2=0 $Y2=0
cc_253 N_A_315_382#_M1010_g N_A_27_367#_c_423_n 0.0114841f $X=2.11 $Y=0.615
+ $X2=0 $Y2=0
cc_254 N_A_315_382#_c_293_n N_A_27_367#_c_423_n 0.00542706f $X=2.13 $Y=1.13
+ $X2=0 $Y2=0
cc_255 N_A_315_382#_c_294_n N_A_27_367#_c_423_n 0.00180888f $X=2.13 $Y=1.13
+ $X2=0 $Y2=0
cc_256 N_A_315_382#_c_298_n N_A_27_367#_c_445_n 0.0525374f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_257 N_A_315_382#_c_298_n N_A_27_367#_c_446_n 0.0143581f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_258 N_A_315_382#_M1010_g N_A_27_367#_c_425_n 0.00359008f $X=2.11 $Y=0.615
+ $X2=0 $Y2=0
cc_259 N_A_315_382#_c_295_n N_A_27_367#_c_425_n 0.0013997f $X=3.335 $Y=0.61
+ $X2=0 $Y2=0
cc_260 N_A_315_382#_M1003_d N_A_27_367#_c_447_n 0.00326506f $X=3.345 $Y=1.975
+ $X2=0 $Y2=0
cc_261 N_A_315_382#_c_298_n N_A_27_367#_c_447_n 0.00570113f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_262 N_A_315_382#_c_303_n N_A_27_367#_c_447_n 0.00150375f $X=3.695 $Y=2.02
+ $X2=0 $Y2=0
cc_263 N_A_315_382#_c_299_n N_A_27_367#_c_448_n 0.0581202f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_264 N_A_315_382#_c_299_n N_A_27_367#_c_426_n 0.0138308f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_265 N_A_315_382#_c_292_n N_A_27_367#_c_426_n 0.0645511f $X=4.67 $Y=2.225
+ $X2=0 $Y2=0
cc_266 N_A_315_382#_c_292_n N_A_27_367#_c_427_n 0.0255711f $X=4.67 $Y=2.225
+ $X2=0 $Y2=0
cc_267 N_A_315_382#_M1010_g N_A_27_367#_c_431_n 3.06083e-19 $X=2.11 $Y=0.615
+ $X2=0 $Y2=0
cc_268 N_A_315_382#_c_293_n N_A_27_367#_c_431_n 0.0242357f $X=2.13 $Y=1.13 $X2=0
+ $Y2=0
cc_269 N_A_315_382#_c_294_n N_A_27_367#_c_431_n 0.00177856f $X=2.13 $Y=1.13
+ $X2=0 $Y2=0
cc_270 N_A_315_382#_c_293_n N_A_27_367#_c_432_n 3.24287e-19 $X=2.13 $Y=1.13
+ $X2=0 $Y2=0
cc_271 N_A_315_382#_c_294_n N_A_27_367#_c_432_n 0.0187224f $X=2.13 $Y=1.13 $X2=0
+ $Y2=0
cc_272 N_A_315_382#_c_298_n N_A_27_367#_c_451_n 0.00879088f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_273 N_A_315_382#_M1003_d N_A_27_367#_c_452_n 0.00250831f $X=3.345 $Y=1.975
+ $X2=0 $Y2=0
cc_274 N_A_315_382#_c_299_n N_A_27_367#_c_452_n 0.00734099f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_275 N_A_315_382#_c_303_n N_A_27_367#_c_452_n 0.0205676f $X=3.695 $Y=2.02
+ $X2=0 $Y2=0
cc_276 N_A_315_382#_c_299_n N_A_27_367#_c_453_n 3.82927e-19 $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_277 N_A_315_382#_c_303_n N_A_27_367#_c_453_n 0.00111382f $X=3.695 $Y=2.02
+ $X2=0 $Y2=0
cc_278 N_A_315_382#_M1010_g N_A_27_367#_c_433_n 0.0243464f $X=2.11 $Y=0.615
+ $X2=0 $Y2=0
cc_279 N_A_315_382#_c_291_n N_A_321_55#_M1013_s 0.00259572f $X=4.585 $Y=0.77
+ $X2=-0.19 $Y2=-0.245
cc_280 N_A_315_382#_c_299_n N_A_321_55#_M1011_s 0.00861385f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_281 N_A_315_382#_M1010_g N_A_321_55#_M1016_g 0.0161138f $X=2.11 $Y=0.615
+ $X2=0 $Y2=0
cc_282 N_A_315_382#_c_290_n N_A_321_55#_M1016_g 0.0039922f $X=2.01 $Y=1.91 $X2=0
+ $Y2=0
cc_283 N_A_315_382#_c_293_n N_A_321_55#_M1016_g 0.001696f $X=2.13 $Y=1.13 $X2=0
+ $Y2=0
cc_284 N_A_315_382#_c_294_n N_A_321_55#_M1016_g 0.0195317f $X=2.13 $Y=1.13 $X2=0
+ $Y2=0
cc_285 N_A_315_382#_c_290_n N_A_321_55#_c_650_n 0.0126942f $X=2.01 $Y=1.91 $X2=0
+ $Y2=0
cc_286 N_A_315_382#_c_298_n N_A_321_55#_c_650_n 4.20204e-19 $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_287 N_A_315_382#_c_302_n N_A_321_55#_c_650_n 0.0025228f $X=2.095 $Y=2.075
+ $X2=0 $Y2=0
cc_288 N_A_315_382#_c_293_n N_A_321_55#_c_650_n 0.00115249f $X=2.13 $Y=1.13
+ $X2=0 $Y2=0
cc_289 N_A_315_382#_c_294_n N_A_321_55#_c_650_n 0.0224321f $X=2.13 $Y=1.13 $X2=0
+ $Y2=0
cc_290 N_A_315_382#_c_301_n N_A_321_55#_c_651_n 0.0186076f $X=1.74 $Y=2.075
+ $X2=0 $Y2=0
cc_291 N_A_315_382#_M1000_g N_A_321_55#_M1009_g 0.0147138f $X=1.65 $Y=2.72 $X2=0
+ $Y2=0
cc_292 N_A_315_382#_c_298_n N_A_321_55#_M1009_g 0.0179904f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_293 N_A_315_382#_c_301_n N_A_321_55#_M1009_g 0.0203408f $X=1.74 $Y=2.075
+ $X2=0 $Y2=0
cc_294 N_A_315_382#_c_302_n N_A_321_55#_M1009_g 0.00458007f $X=2.095 $Y=2.075
+ $X2=0 $Y2=0
cc_295 N_A_315_382#_c_295_n N_A_321_55#_M1012_g 0.00128551f $X=3.335 $Y=0.61
+ $X2=0 $Y2=0
cc_296 N_A_315_382#_c_298_n N_A_321_55#_c_664_n 0.0151832f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_297 N_A_315_382#_c_303_n N_A_321_55#_c_664_n 0.0073256f $X=3.695 $Y=2.02
+ $X2=0 $Y2=0
cc_298 N_A_315_382#_c_290_n N_A_321_55#_c_653_n 0.00921967f $X=2.01 $Y=1.91
+ $X2=0 $Y2=0
cc_299 N_A_315_382#_c_298_n N_A_321_55#_c_655_n 0.0174129f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_300 N_A_315_382#_c_298_n N_A_321_55#_c_656_n 0.00122406f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_301 N_A_315_382#_c_290_n N_A_321_55#_c_699_n 0.0199478f $X=2.01 $Y=1.91 $X2=0
+ $Y2=0
cc_302 N_A_315_382#_c_298_n N_A_321_55#_c_699_n 0.0771009f $X=3.565 $Y=2.02
+ $X2=0 $Y2=0
cc_303 N_A_315_382#_c_293_n N_A_321_55#_c_699_n 9.03003e-19 $X=2.13 $Y=1.13
+ $X2=0 $Y2=0
cc_304 N_A_315_382#_c_295_n N_A_321_55#_c_657_n 0.0075809f $X=3.335 $Y=0.61
+ $X2=0 $Y2=0
cc_305 N_A_315_382#_c_291_n N_A_321_55#_c_658_n 0.0446003f $X=4.585 $Y=0.77
+ $X2=0 $Y2=0
cc_306 N_A_315_382#_c_295_n N_A_321_55#_c_658_n 0.0168275f $X=3.335 $Y=0.61
+ $X2=0 $Y2=0
cc_307 N_A_315_382#_c_291_n N_A_321_55#_c_705_n 0.0189505f $X=4.585 $Y=0.77
+ $X2=0 $Y2=0
cc_308 N_A_315_382#_c_292_n N_A_321_55#_c_705_n 0.00840018f $X=4.67 $Y=2.225
+ $X2=0 $Y2=0
cc_309 N_A_315_382#_c_299_n N_A_321_55#_c_659_n 0.0267445f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_310 N_A_315_382#_c_292_n N_A_321_55#_c_659_n 0.0609824f $X=4.67 $Y=2.225
+ $X2=0 $Y2=0
cc_311 N_A_315_382#_c_303_n N_A_321_55#_c_659_n 0.00730302f $X=3.695 $Y=2.02
+ $X2=0 $Y2=0
cc_312 N_A_315_382#_c_295_n N_A_321_55#_c_660_n 0.00120843f $X=3.335 $Y=0.61
+ $X2=0 $Y2=0
cc_313 N_A_315_382#_c_299_n N_CLK_c_756_n 0.00453651f $X=4.585 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_314 N_A_315_382#_c_291_n N_CLK_M1013_g 0.01263f $X=4.585 $Y=0.77 $X2=0 $Y2=0
cc_315 N_A_315_382#_c_292_n N_CLK_M1013_g 0.0055748f $X=4.67 $Y=2.225 $X2=0
+ $Y2=0
cc_316 N_A_315_382#_c_299_n N_CLK_c_765_n 0.0140779f $X=4.585 $Y=2.31 $X2=0
+ $Y2=0
cc_317 N_A_315_382#_c_292_n N_CLK_c_765_n 0.0162531f $X=4.67 $Y=2.225 $X2=0
+ $Y2=0
cc_318 N_A_315_382#_c_303_n N_CLK_c_765_n 0.00417533f $X=3.695 $Y=2.02 $X2=0
+ $Y2=0
cc_319 N_A_315_382#_c_292_n N_CLK_c_758_n 0.00703249f $X=4.67 $Y=2.225 $X2=0
+ $Y2=0
cc_320 N_A_315_382#_c_299_n N_CLK_c_759_n 0.00145537f $X=4.585 $Y=2.31 $X2=0
+ $Y2=0
cc_321 N_A_315_382#_c_292_n N_CLK_c_759_n 0.00417338f $X=4.67 $Y=2.225 $X2=0
+ $Y2=0
cc_322 N_A_315_382#_c_291_n N_CLK_M1007_g 0.00318195f $X=4.585 $Y=0.77 $X2=0
+ $Y2=0
cc_323 N_A_315_382#_c_292_n N_CLK_M1007_g 0.00848375f $X=4.67 $Y=2.225 $X2=0
+ $Y2=0
cc_324 N_A_315_382#_c_299_n N_CLK_c_768_n 5.29316e-19 $X=4.585 $Y=2.31 $X2=0
+ $Y2=0
cc_325 N_A_315_382#_c_292_n N_CLK_c_768_n 0.00123648f $X=4.67 $Y=2.225 $X2=0
+ $Y2=0
cc_326 N_A_315_382#_c_298_n N_CLK_c_762_n 0.00795663f $X=3.565 $Y=2.02 $X2=0
+ $Y2=0
cc_327 N_A_315_382#_c_299_n N_CLK_c_762_n 0.0035978f $X=4.585 $Y=2.31 $X2=0
+ $Y2=0
cc_328 N_A_315_382#_c_303_n N_CLK_c_762_n 0.0222053f $X=3.695 $Y=2.02 $X2=0
+ $Y2=0
cc_329 N_A_315_382#_c_299_n N_CLK_c_763_n 0.00130879f $X=4.585 $Y=2.31 $X2=0
+ $Y2=0
cc_330 N_A_315_382#_c_303_n N_CLK_c_763_n 0.00152906f $X=3.695 $Y=2.02 $X2=0
+ $Y2=0
cc_331 N_A_315_382#_c_291_n N_A_1046_367#_c_836_n 0.00468066f $X=4.585 $Y=0.77
+ $X2=0 $Y2=0
cc_332 N_A_315_382#_c_298_n N_VPWR_M1001_d 0.00626267f $X=3.565 $Y=2.02 $X2=0
+ $Y2=0
cc_333 N_A_315_382#_c_299_n N_VPWR_M1011_d 0.00220447f $X=4.585 $Y=2.31 $X2=0
+ $Y2=0
cc_334 N_A_315_382#_c_292_n N_VPWR_M1011_d 0.0034563f $X=4.67 $Y=2.225 $X2=0
+ $Y2=0
cc_335 N_A_315_382#_M1000_g N_VPWR_c_894_n 0.00322875f $X=1.65 $Y=2.72 $X2=0
+ $Y2=0
cc_336 N_A_315_382#_M1000_g N_VPWR_c_889_n 0.00556106f $X=1.65 $Y=2.72 $X2=0
+ $Y2=0
cc_337 N_A_315_382#_c_291_n N_VGND_M1013_d 0.0121517f $X=4.585 $Y=0.77 $X2=0
+ $Y2=0
cc_338 N_A_315_382#_c_292_n N_VGND_M1013_d 0.0072819f $X=4.67 $Y=2.225 $X2=0
+ $Y2=0
cc_339 N_A_315_382#_c_291_n N_VGND_c_994_n 0.0256982f $X=4.585 $Y=0.77 $X2=0
+ $Y2=0
cc_340 N_A_315_382#_M1010_g N_VGND_c_998_n 9.15902e-19 $X=2.11 $Y=0.615 $X2=0
+ $Y2=0
cc_341 N_A_315_382#_c_291_n N_VGND_c_1000_n 0.0154511f $X=4.585 $Y=0.77 $X2=0
+ $Y2=0
cc_342 N_A_315_382#_c_295_n N_VGND_c_1000_n 0.00815599f $X=3.335 $Y=0.61 $X2=0
+ $Y2=0
cc_343 N_A_315_382#_c_291_n N_VGND_c_1003_n 0.0272557f $X=4.585 $Y=0.77 $X2=0
+ $Y2=0
cc_344 N_A_315_382#_c_295_n N_VGND_c_1003_n 0.00981596f $X=3.335 $Y=0.61 $X2=0
+ $Y2=0
cc_345 N_A_27_367#_c_422_n N_A_321_55#_M1016_g 5.98939e-19 $X=1.245 $Y=0.905
+ $X2=0 $Y2=0
cc_346 N_A_27_367#_c_423_n N_A_321_55#_M1016_g 0.00935878f $X=2.45 $Y=0.34 $X2=0
+ $Y2=0
cc_347 N_A_27_367#_M1001_g N_A_321_55#_M1009_g 0.0366693f $X=2.55 $Y=2.61 $X2=0
+ $Y2=0
cc_348 N_A_27_367#_c_442_n N_A_321_55#_M1009_g 0.0107162f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_349 N_A_27_367#_c_444_n N_A_321_55#_M1009_g 0.00336109f $X=2.36 $Y=2.905
+ $X2=0 $Y2=0
cc_350 N_A_27_367#_c_446_n N_A_321_55#_M1009_g 0.00418393f $X=2.445 $Y=2.36
+ $X2=0 $Y2=0
cc_351 N_A_27_367#_c_425_n N_A_321_55#_M1012_g 7.83566e-19 $X=2.535 $Y=0.95
+ $X2=0 $Y2=0
cc_352 N_A_27_367#_c_431_n N_A_321_55#_M1012_g 7.76287e-19 $X=2.67 $Y=1.1 $X2=0
+ $Y2=0
cc_353 N_A_27_367#_c_432_n N_A_321_55#_M1012_g 0.0209541f $X=2.67 $Y=1.1 $X2=0
+ $Y2=0
cc_354 N_A_27_367#_c_433_n N_A_321_55#_M1012_g 0.0112139f $X=2.67 $Y=0.935 $X2=0
+ $Y2=0
cc_355 N_A_27_367#_M1001_g N_A_321_55#_c_664_n 0.00789379f $X=2.55 $Y=2.61 $X2=0
+ $Y2=0
cc_356 N_A_27_367#_c_435_n N_A_321_55#_c_664_n 0.00608234f $X=3.585 $Y=3.115
+ $X2=0 $Y2=0
cc_357 N_A_27_367#_c_445_n N_A_321_55#_c_664_n 0.00512953f $X=3.225 $Y=2.36
+ $X2=0 $Y2=0
cc_358 N_A_27_367#_c_447_n N_A_321_55#_c_664_n 0.00168274f $X=3.585 $Y=2.655
+ $X2=0 $Y2=0
cc_359 N_A_27_367#_c_451_n N_A_321_55#_c_664_n 0.018776f $X=3.31 $Y=2.36 $X2=0
+ $Y2=0
cc_360 N_A_27_367#_M1001_g N_A_321_55#_c_655_n 0.00371611f $X=2.55 $Y=2.61 $X2=0
+ $Y2=0
cc_361 N_A_27_367#_c_431_n N_A_321_55#_c_655_n 0.00245418f $X=2.67 $Y=1.1 $X2=0
+ $Y2=0
cc_362 N_A_27_367#_c_432_n N_A_321_55#_c_655_n 0.0176822f $X=2.67 $Y=1.1 $X2=0
+ $Y2=0
cc_363 N_A_27_367#_c_431_n N_A_321_55#_c_699_n 0.0216935f $X=2.67 $Y=1.1 $X2=0
+ $Y2=0
cc_364 N_A_27_367#_c_432_n N_A_321_55#_c_699_n 0.00130494f $X=2.67 $Y=1.1 $X2=0
+ $Y2=0
cc_365 N_A_27_367#_c_431_n N_A_321_55#_c_657_n 0.0153173f $X=2.67 $Y=1.1 $X2=0
+ $Y2=0
cc_366 N_A_27_367#_c_432_n N_A_321_55#_c_657_n 2.80642e-19 $X=2.67 $Y=1.1 $X2=0
+ $Y2=0
cc_367 N_A_27_367#_c_431_n N_A_321_55#_c_733_n 8.52574e-19 $X=2.67 $Y=1.1 $X2=0
+ $Y2=0
cc_368 N_A_27_367#_c_448_n N_CLK_c_765_n 0.00667685f $X=4.925 $Y=2.65 $X2=0
+ $Y2=0
cc_369 N_A_27_367#_c_426_n N_CLK_c_765_n 0.00508919f $X=5.01 $Y=2.565 $X2=0
+ $Y2=0
cc_370 N_A_27_367#_M1005_g N_CLK_M1007_g 0.0546692f $X=5.295 $Y=0.605 $X2=0
+ $Y2=0
cc_371 N_A_27_367#_M1017_g N_CLK_M1007_g 0.00447751f $X=5.585 $Y=2.155 $X2=0
+ $Y2=0
cc_372 N_A_27_367#_c_426_n N_CLK_M1007_g 0.00599029f $X=5.01 $Y=2.565 $X2=0
+ $Y2=0
cc_373 N_A_27_367#_c_427_n N_CLK_M1007_g 0.0126905f $X=5.095 $Y=1.165 $X2=0
+ $Y2=0
cc_374 N_A_27_367#_c_429_n N_CLK_M1007_g 0.00642656f $X=5.51 $Y=1.17 $X2=0 $Y2=0
cc_375 N_A_27_367#_c_448_n N_CLK_c_768_n 0.00160564f $X=4.925 $Y=2.65 $X2=0
+ $Y2=0
cc_376 N_A_27_367#_c_426_n N_CLK_c_768_n 0.017458f $X=5.01 $Y=2.565 $X2=0 $Y2=0
cc_377 N_A_27_367#_M1017_g N_CLK_c_761_n 0.0153595f $X=5.585 $Y=2.155 $X2=0
+ $Y2=0
cc_378 N_A_27_367#_c_426_n N_CLK_c_761_n 0.00919164f $X=5.01 $Y=2.565 $X2=0
+ $Y2=0
cc_379 N_A_27_367#_c_428_n N_CLK_c_761_n 0.00529729f $X=5.51 $Y=1.17 $X2=0 $Y2=0
cc_380 N_A_27_367#_c_429_n N_CLK_c_761_n 2.61989e-19 $X=5.51 $Y=1.17 $X2=0 $Y2=0
cc_381 N_A_27_367#_c_428_n N_A_1046_367#_M1014_g 2.98545e-19 $X=5.51 $Y=1.17
+ $X2=0 $Y2=0
cc_382 N_A_27_367#_c_429_n N_A_1046_367#_M1014_g 0.00647706f $X=5.51 $Y=1.17
+ $X2=0 $Y2=0
cc_383 N_A_27_367#_M1017_g N_A_1046_367#_M1015_g 0.0117393f $X=5.585 $Y=2.155
+ $X2=0 $Y2=0
cc_384 N_A_27_367#_M1017_g N_A_1046_367#_c_839_n 0.00433882f $X=5.585 $Y=2.155
+ $X2=0 $Y2=0
cc_385 N_A_27_367#_c_426_n N_A_1046_367#_c_839_n 0.0353065f $X=5.01 $Y=2.565
+ $X2=0 $Y2=0
cc_386 N_A_27_367#_M1017_g N_A_1046_367#_c_832_n 0.0142306f $X=5.585 $Y=2.155
+ $X2=0 $Y2=0
cc_387 N_A_27_367#_c_428_n N_A_1046_367#_c_832_n 0.0151465f $X=5.51 $Y=1.17
+ $X2=0 $Y2=0
cc_388 N_A_27_367#_c_429_n N_A_1046_367#_c_832_n 0.00135885f $X=5.51 $Y=1.17
+ $X2=0 $Y2=0
cc_389 N_A_27_367#_c_426_n N_A_1046_367#_c_833_n 0.0140162f $X=5.01 $Y=2.565
+ $X2=0 $Y2=0
cc_390 N_A_27_367#_c_428_n N_A_1046_367#_c_833_n 0.0171596f $X=5.51 $Y=1.17
+ $X2=0 $Y2=0
cc_391 N_A_27_367#_c_429_n N_A_1046_367#_c_833_n 0.00334892f $X=5.51 $Y=1.17
+ $X2=0 $Y2=0
cc_392 N_A_27_367#_M1005_g N_A_1046_367#_c_835_n 0.00397467f $X=5.295 $Y=0.605
+ $X2=0 $Y2=0
cc_393 N_A_27_367#_M1017_g N_A_1046_367#_c_835_n 9.96517e-19 $X=5.585 $Y=2.155
+ $X2=0 $Y2=0
cc_394 N_A_27_367#_c_428_n N_A_1046_367#_c_835_n 0.0183533f $X=5.51 $Y=1.17
+ $X2=0 $Y2=0
cc_395 N_A_27_367#_c_429_n N_A_1046_367#_c_835_n 0.00154738f $X=5.51 $Y=1.17
+ $X2=0 $Y2=0
cc_396 N_A_27_367#_M1005_g N_A_1046_367#_c_836_n 0.00830845f $X=5.295 $Y=0.605
+ $X2=0 $Y2=0
cc_397 N_A_27_367#_c_428_n N_A_1046_367#_c_836_n 0.026303f $X=5.51 $Y=1.17 $X2=0
+ $Y2=0
cc_398 N_A_27_367#_c_429_n N_A_1046_367#_c_836_n 0.00755495f $X=5.51 $Y=1.17
+ $X2=0 $Y2=0
cc_399 N_A_27_367#_M1017_g N_A_1046_367#_c_837_n 0.0150761f $X=5.585 $Y=2.155
+ $X2=0 $Y2=0
cc_400 N_A_27_367#_c_440_n N_VPWR_M1019_d 0.00511041f $X=0.975 $Y=1.985
+ $X2=-0.19 $Y2=-0.245
cc_401 N_A_27_367#_c_441_n N_VPWR_M1019_d 0.0126791f $X=1.06 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_402 N_A_27_367#_c_442_n N_VPWR_M1019_d 4.57867e-19 $X=2.275 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_403 N_A_27_367#_c_443_n N_VPWR_M1019_d 0.00174567f $X=1.145 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_404 N_A_27_367#_c_445_n N_VPWR_M1001_d 0.0117532f $X=3.225 $Y=2.36 $X2=0
+ $Y2=0
cc_405 N_A_27_367#_c_448_n N_VPWR_M1011_d 0.0105579f $X=4.925 $Y=2.65 $X2=0
+ $Y2=0
cc_406 N_A_27_367#_c_426_n N_VPWR_M1011_d 0.00703775f $X=5.01 $Y=2.565 $X2=0
+ $Y2=0
cc_407 N_A_27_367#_c_440_n N_VPWR_c_890_n 0.0160276f $X=0.975 $Y=1.985 $X2=0
+ $Y2=0
cc_408 N_A_27_367#_c_441_n N_VPWR_c_890_n 0.0490737f $X=1.06 $Y=2.905 $X2=0
+ $Y2=0
cc_409 N_A_27_367#_c_443_n N_VPWR_c_890_n 0.0140458f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_410 N_A_27_367#_M1001_g N_VPWR_c_891_n 0.00827967f $X=2.55 $Y=2.61 $X2=0
+ $Y2=0
cc_411 N_A_27_367#_c_435_n N_VPWR_c_891_n 0.0249849f $X=3.585 $Y=3.115 $X2=0
+ $Y2=0
cc_412 N_A_27_367#_c_442_n N_VPWR_c_891_n 0.0107161f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_413 N_A_27_367#_c_444_n N_VPWR_c_891_n 0.0106679f $X=2.36 $Y=2.905 $X2=0
+ $Y2=0
cc_414 N_A_27_367#_c_445_n N_VPWR_c_891_n 0.0266856f $X=3.225 $Y=2.36 $X2=0
+ $Y2=0
cc_415 N_A_27_367#_c_451_n N_VPWR_c_891_n 0.00920481f $X=3.31 $Y=2.36 $X2=0
+ $Y2=0
cc_416 N_A_27_367#_c_452_n N_VPWR_c_891_n 0.0105711f $X=3.75 $Y=2.65 $X2=0 $Y2=0
cc_417 N_A_27_367#_c_453_n N_VPWR_c_891_n 0.00461972f $X=3.75 $Y=2.94 $X2=0
+ $Y2=0
cc_418 N_A_27_367#_c_448_n N_VPWR_c_892_n 0.0254965f $X=4.925 $Y=2.65 $X2=0
+ $Y2=0
cc_419 N_A_27_367#_M1017_g N_VPWR_c_893_n 0.0118465f $X=5.585 $Y=2.155 $X2=0
+ $Y2=0
cc_420 N_A_27_367#_c_448_n N_VPWR_c_893_n 0.00663281f $X=4.925 $Y=2.65 $X2=0
+ $Y2=0
cc_421 N_A_27_367#_c_426_n N_VPWR_c_893_n 0.00200972f $X=5.01 $Y=2.565 $X2=0
+ $Y2=0
cc_422 N_A_27_367#_c_436_n N_VPWR_c_894_n 0.00876931f $X=2.625 $Y=3.115 $X2=0
+ $Y2=0
cc_423 N_A_27_367#_c_442_n N_VPWR_c_894_n 0.0840479f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_424 N_A_27_367#_c_443_n N_VPWR_c_894_n 0.0121867f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_425 N_A_27_367#_c_435_n N_VPWR_c_896_n 0.0213306f $X=3.585 $Y=3.115 $X2=0
+ $Y2=0
cc_426 N_A_27_367#_c_447_n N_VPWR_c_896_n 0.00387812f $X=3.585 $Y=2.655 $X2=0
+ $Y2=0
cc_427 N_A_27_367#_c_448_n N_VPWR_c_896_n 0.0155084f $X=4.925 $Y=2.65 $X2=0
+ $Y2=0
cc_428 N_A_27_367#_c_451_n N_VPWR_c_896_n 0.0034135f $X=3.31 $Y=2.36 $X2=0 $Y2=0
cc_429 N_A_27_367#_c_452_n N_VPWR_c_896_n 0.0219012f $X=3.75 $Y=2.65 $X2=0 $Y2=0
cc_430 N_A_27_367#_c_439_n N_VPWR_c_898_n 0.0210467f $X=0.26 $Y=2.91 $X2=0 $Y2=0
cc_431 N_A_27_367#_M1017_g N_VPWR_c_899_n 0.00259749f $X=5.585 $Y=2.155 $X2=0
+ $Y2=0
cc_432 N_A_27_367#_c_448_n N_VPWR_c_899_n 0.00153289f $X=4.925 $Y=2.65 $X2=0
+ $Y2=0
cc_433 N_A_27_367#_M1019_s N_VPWR_c_889_n 0.00215158f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_434 N_A_27_367#_c_435_n N_VPWR_c_889_n 0.0239353f $X=3.585 $Y=3.115 $X2=0
+ $Y2=0
cc_435 N_A_27_367#_c_436_n N_VPWR_c_889_n 0.0110375f $X=2.625 $Y=3.115 $X2=0
+ $Y2=0
cc_436 N_A_27_367#_M1017_g N_VPWR_c_889_n 0.00344639f $X=5.585 $Y=2.155 $X2=0
+ $Y2=0
cc_437 N_A_27_367#_c_439_n N_VPWR_c_889_n 0.0125583f $X=0.26 $Y=2.91 $X2=0 $Y2=0
cc_438 N_A_27_367#_c_442_n N_VPWR_c_889_n 0.0477215f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_439 N_A_27_367#_c_443_n N_VPWR_c_889_n 0.00660921f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_440 N_A_27_367#_c_447_n N_VPWR_c_889_n 0.00488291f $X=3.585 $Y=2.655 $X2=0
+ $Y2=0
cc_441 N_A_27_367#_c_448_n N_VPWR_c_889_n 0.0269115f $X=4.925 $Y=2.65 $X2=0
+ $Y2=0
cc_442 N_A_27_367#_c_451_n N_VPWR_c_889_n 0.0044027f $X=3.31 $Y=2.36 $X2=0 $Y2=0
cc_443 N_A_27_367#_c_452_n N_VPWR_c_889_n 0.0111578f $X=3.75 $Y=2.65 $X2=0 $Y2=0
cc_444 N_A_27_367#_c_453_n N_VPWR_c_889_n 0.00961448f $X=3.75 $Y=2.94 $X2=0
+ $Y2=0
cc_445 N_A_27_367#_c_442_n A_273_480# 0.00101072f $X=2.275 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_446 N_A_27_367#_c_444_n A_453_480# 5.4199e-19 $X=2.36 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_447 N_A_27_367#_c_422_n N_VGND_M1008_d 0.0100754f $X=1.245 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
cc_448 N_A_27_367#_c_422_n N_VGND_c_992_n 0.0247837f $X=1.245 $Y=0.905 $X2=0
+ $Y2=0
cc_449 N_A_27_367#_c_475_n N_VGND_c_992_n 0.0166147f $X=1.33 $Y=0.82 $X2=0 $Y2=0
cc_450 N_A_27_367#_c_424_n N_VGND_c_992_n 0.0143263f $X=1.415 $Y=0.34 $X2=0
+ $Y2=0
cc_451 N_A_27_367#_c_423_n N_VGND_c_993_n 0.014035f $X=2.45 $Y=0.34 $X2=0 $Y2=0
cc_452 N_A_27_367#_c_425_n N_VGND_c_993_n 0.0256554f $X=2.535 $Y=0.95 $X2=0
+ $Y2=0
cc_453 N_A_27_367#_c_431_n N_VGND_c_993_n 0.00362176f $X=2.67 $Y=1.1 $X2=0 $Y2=0
cc_454 N_A_27_367#_c_432_n N_VGND_c_993_n 0.00104367f $X=2.67 $Y=1.1 $X2=0 $Y2=0
cc_455 N_A_27_367#_c_433_n N_VGND_c_993_n 0.00370862f $X=2.67 $Y=0.935 $X2=0
+ $Y2=0
cc_456 N_A_27_367#_M1005_g N_VGND_c_995_n 0.00425581f $X=5.295 $Y=0.605 $X2=0
+ $Y2=0
cc_457 N_A_27_367#_c_420_n N_VGND_c_996_n 0.0318172f $X=0.415 $Y=0.42 $X2=0
+ $Y2=0
cc_458 N_A_27_367#_c_423_n N_VGND_c_998_n 0.0788214f $X=2.45 $Y=0.34 $X2=0 $Y2=0
cc_459 N_A_27_367#_c_424_n N_VGND_c_998_n 0.0121867f $X=1.415 $Y=0.34 $X2=0
+ $Y2=0
cc_460 N_A_27_367#_c_433_n N_VGND_c_998_n 0.00198997f $X=2.67 $Y=0.935 $X2=0
+ $Y2=0
cc_461 N_A_27_367#_M1005_g N_VGND_c_1001_n 0.00535318f $X=5.295 $Y=0.605 $X2=0
+ $Y2=0
cc_462 N_A_27_367#_M1008_s N_VGND_c_1003_n 0.00215158f $X=0.29 $Y=0.235 $X2=0
+ $Y2=0
cc_463 N_A_27_367#_M1005_g N_VGND_c_1003_n 0.00537853f $X=5.295 $Y=0.605 $X2=0
+ $Y2=0
cc_464 N_A_27_367#_c_420_n N_VGND_c_1003_n 0.0184234f $X=0.415 $Y=0.42 $X2=0
+ $Y2=0
cc_465 N_A_27_367#_c_422_n N_VGND_c_1003_n 0.0119678f $X=1.245 $Y=0.905 $X2=0
+ $Y2=0
cc_466 N_A_27_367#_c_423_n N_VGND_c_1003_n 0.0455187f $X=2.45 $Y=0.34 $X2=0
+ $Y2=0
cc_467 N_A_27_367#_c_424_n N_VGND_c_1003_n 0.00660921f $X=1.415 $Y=0.34 $X2=0
+ $Y2=0
cc_468 N_A_27_367#_c_433_n N_VGND_c_1003_n 0.00124755f $X=2.67 $Y=0.935 $X2=0
+ $Y2=0
cc_469 N_A_27_367#_c_423_n A_279_81# 0.00366293f $X=2.45 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_470 N_A_27_367#_c_423_n A_437_81# 0.00668583f $X=2.45 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_471 N_A_321_55#_c_658_n N_CLK_c_756_n 0.00417045f $X=4.085 $Y=1.137 $X2=-0.19
+ $Y2=-0.245
cc_472 N_A_321_55#_c_659_n N_CLK_c_756_n 0.0106356f $X=4.25 $Y=1.96 $X2=-0.19
+ $Y2=-0.245
cc_473 N_A_321_55#_c_705_n N_CLK_M1013_g 0.00701443f $X=4.25 $Y=1.25 $X2=0 $Y2=0
cc_474 N_A_321_55#_c_659_n N_CLK_M1013_g 0.0111295f $X=4.25 $Y=1.96 $X2=0 $Y2=0
cc_475 N_A_321_55#_c_659_n N_CLK_c_765_n 0.00690867f $X=4.25 $Y=1.96 $X2=0 $Y2=0
cc_476 N_A_321_55#_c_659_n N_CLK_c_759_n 0.00832448f $X=4.25 $Y=1.96 $X2=0 $Y2=0
cc_477 N_A_321_55#_c_654_n N_CLK_c_762_n 0.00259386f $X=3.21 $Y=1.505 $X2=0
+ $Y2=0
cc_478 N_A_321_55#_c_656_n N_CLK_c_762_n 3.99748e-19 $X=3.045 $Y=1.505 $X2=0
+ $Y2=0
cc_479 N_A_321_55#_c_699_n N_CLK_c_762_n 0.0223588f $X=3.045 $Y=1.635 $X2=0
+ $Y2=0
cc_480 N_A_321_55#_c_733_n N_CLK_c_762_n 0.00667946f $X=3.17 $Y=1.505 $X2=0
+ $Y2=0
cc_481 N_A_321_55#_c_658_n N_CLK_c_762_n 0.0352956f $X=4.085 $Y=1.137 $X2=0
+ $Y2=0
cc_482 N_A_321_55#_c_659_n N_CLK_c_762_n 0.0273492f $X=4.25 $Y=1.96 $X2=0 $Y2=0
cc_483 N_A_321_55#_c_654_n N_CLK_c_763_n 0.01797f $X=3.21 $Y=1.505 $X2=0 $Y2=0
cc_484 N_A_321_55#_c_699_n N_CLK_c_763_n 2.05464e-19 $X=3.045 $Y=1.635 $X2=0
+ $Y2=0
cc_485 N_A_321_55#_c_658_n N_CLK_c_763_n 0.00793179f $X=4.085 $Y=1.137 $X2=0
+ $Y2=0
cc_486 N_A_321_55#_c_659_n N_CLK_c_763_n 0.00136876f $X=4.25 $Y=1.96 $X2=0 $Y2=0
cc_487 N_A_321_55#_c_664_n N_VPWR_c_891_n 0.00118821f $X=3.27 $Y=1.865 $X2=0
+ $Y2=0
cc_488 N_A_321_55#_M1009_g N_VPWR_c_894_n 6.91459e-19 $X=2.19 $Y=2.61 $X2=0
+ $Y2=0
cc_489 N_A_321_55#_M1012_g N_VGND_c_993_n 0.00382769f $X=3.12 $Y=0.615 $X2=0
+ $Y2=0
cc_490 N_A_321_55#_M1016_g N_VGND_c_998_n 9.15902e-19 $X=1.68 $Y=0.615 $X2=0
+ $Y2=0
cc_491 N_A_321_55#_M1012_g N_VGND_c_1000_n 0.00552345f $X=3.12 $Y=0.615 $X2=0
+ $Y2=0
cc_492 N_A_321_55#_M1012_g N_VGND_c_1003_n 0.00534666f $X=3.12 $Y=0.615 $X2=0
+ $Y2=0
cc_493 N_CLK_c_761_n N_A_1046_367#_c_839_n 0.00150545f $X=5.155 $Y=1.65 $X2=0
+ $Y2=0
cc_494 N_CLK_M1007_g N_A_1046_367#_c_833_n 2.99725e-19 $X=4.935 $Y=0.605 $X2=0
+ $Y2=0
cc_495 N_CLK_c_761_n N_A_1046_367#_c_833_n 9.28488e-19 $X=5.155 $Y=1.65 $X2=0
+ $Y2=0
cc_496 N_CLK_M1007_g N_A_1046_367#_c_836_n 0.00150674f $X=4.935 $Y=0.605 $X2=0
+ $Y2=0
cc_497 N_CLK_c_768_n N_VPWR_c_893_n 5.08223e-19 $X=5.155 $Y=1.725 $X2=0 $Y2=0
cc_498 N_CLK_c_765_n N_VPWR_c_896_n 4.81819e-19 $X=4.565 $Y=1.725 $X2=0 $Y2=0
cc_499 N_CLK_c_768_n N_VPWR_c_899_n 0.00285987f $X=5.155 $Y=1.725 $X2=0 $Y2=0
cc_500 N_CLK_c_768_n N_VPWR_c_889_n 0.00369256f $X=5.155 $Y=1.725 $X2=0 $Y2=0
cc_501 N_CLK_M1007_g N_VGND_c_994_n 0.00910687f $X=4.935 $Y=0.605 $X2=0 $Y2=0
cc_502 N_CLK_M1013_g N_VGND_c_1000_n 5.44798e-19 $X=4.31 $Y=1.035 $X2=0 $Y2=0
cc_503 N_CLK_M1007_g N_VGND_c_1001_n 0.00559701f $X=4.935 $Y=0.605 $X2=0 $Y2=0
cc_504 N_CLK_M1007_g N_VGND_c_1003_n 0.00537853f $X=4.935 $Y=0.605 $X2=0 $Y2=0
cc_505 N_A_1046_367#_M1015_g N_VPWR_c_893_n 0.0311271f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_506 N_A_1046_367#_c_839_n N_VPWR_c_893_n 0.0275831f $X=5.37 $Y=1.96 $X2=0
+ $Y2=0
cc_507 N_A_1046_367#_c_832_n N_VPWR_c_893_n 0.0227566f $X=5.945 $Y=1.58 $X2=0
+ $Y2=0
cc_508 N_A_1046_367#_c_835_n N_VPWR_c_893_n 0.0191281f $X=6.07 $Y=1.495 $X2=0
+ $Y2=0
cc_509 N_A_1046_367#_c_837_n N_VPWR_c_893_n 0.00160808f $X=6.11 $Y=1.5 $X2=0
+ $Y2=0
cc_510 N_A_1046_367#_M1015_g N_VPWR_c_900_n 0.00486043f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_511 N_A_1046_367#_M1015_g N_VPWR_c_889_n 0.00917987f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_512 N_A_1046_367#_c_839_n N_VPWR_c_889_n 0.00784141f $X=5.37 $Y=1.96 $X2=0
+ $Y2=0
cc_513 N_A_1046_367#_M1014_g N_GCLK_c_982_n 0.0269401f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_514 N_A_1046_367#_c_835_n N_GCLK_c_982_n 0.0544518f $X=6.07 $Y=1.495 $X2=0
+ $Y2=0
cc_515 N_A_1046_367#_c_834_n N_VGND_M1014_s 0.00375745f $X=5.945 $Y=0.75 $X2=0
+ $Y2=0
cc_516 N_A_1046_367#_c_835_n N_VGND_M1014_s 0.00422169f $X=6.07 $Y=1.495 $X2=0
+ $Y2=0
cc_517 N_A_1046_367#_c_836_n N_VGND_c_994_n 0.00223361f $X=5.51 $Y=0.605 $X2=0
+ $Y2=0
cc_518 N_A_1046_367#_M1014_g N_VGND_c_995_n 0.00937641f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_519 N_A_1046_367#_c_834_n N_VGND_c_995_n 0.0223095f $X=5.945 $Y=0.75 $X2=0
+ $Y2=0
cc_520 N_A_1046_367#_c_836_n N_VGND_c_995_n 0.00423513f $X=5.51 $Y=0.605 $X2=0
+ $Y2=0
cc_521 N_A_1046_367#_c_834_n N_VGND_c_1001_n 0.00324506f $X=5.945 $Y=0.75 $X2=0
+ $Y2=0
cc_522 N_A_1046_367#_c_836_n N_VGND_c_1001_n 0.00921768f $X=5.51 $Y=0.605 $X2=0
+ $Y2=0
cc_523 N_A_1046_367#_M1014_g N_VGND_c_1002_n 0.00486043f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_524 N_A_1046_367#_M1014_g N_VGND_c_1003_n 0.00917987f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_525 N_A_1046_367#_c_834_n N_VGND_c_1003_n 0.00686771f $X=5.945 $Y=0.75 $X2=0
+ $Y2=0
cc_526 N_A_1046_367#_c_836_n N_VGND_c_1003_n 0.0111687f $X=5.51 $Y=0.605 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_889_n N_GCLK_M1015_d 0.00371702f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_528 N_VPWR_c_900_n N_GCLK_c_982_n 0.0178111f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_529 N_VPWR_c_889_n N_GCLK_c_982_n 0.0100304f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_530 N_GCLK_c_982_n N_VGND_c_1002_n 0.0178111f $X=6.46 $Y=0.42 $X2=0 $Y2=0
cc_531 N_GCLK_M1014_d N_VGND_c_1003_n 0.00371702f $X=6.32 $Y=0.235 $X2=0 $Y2=0
cc_532 N_GCLK_c_982_n N_VGND_c_1003_n 0.0100304f $X=6.46 $Y=0.42 $X2=0 $Y2=0
