* File: sky130_fd_sc_lp__a2bb2o_m.spice
* Created: Fri Aug 28 09:56:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2o_m.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2o_m  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_85_345#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1004 N_A_210_125#_M1004_d N_A1_N_M1004_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.114875 AS=0.0588 PD=1.015 PS=0.7 NRD=62.424 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A2_N_M1001_g N_A_210_125#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.114875 PD=0.7 PS=1.015 NRD=0 NRS=62.424 M=1 R=2.8
+ SA=75001.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1002 N_A_85_345#_M1002_d N_A_210_125#_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.11235 AS=0.0588 PD=0.955 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 A_551_125# N_B2_M1009_g N_A_85_345#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.11235 PD=0.81 PS=0.955 NRD=39.996 NRS=72.852 M=1 R=2.8
+ SA=75002.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_B1_M1010_g A_551_125# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75002.9 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_85_345#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=9.3772 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_223_535# N_A1_N_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_210_125#_M1007_d N_A2_N_M1007_g A_223_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1141 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_479_429#_M1011_d N_A_210_125#_M1011_g N_A_85_345#_M1011_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1141 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_B2_M1005_g N_A_479_429#_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_479_429#_M1008_d N_B1_M1008_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0735 PD=1.37 PS=0.77 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_71 VPB 0 2.80181e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a2bb2o_m.pxi.spice"
*
.ends
*
*
