* File: sky130_fd_sc_lp__bushold0_1.pex.spice
* Created: Wed Sep  2 09:37:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUSHOLD0_1%X 1 2 9 13 17 18 21 22 24 25 28 30 31 32
+ 33 34 35 36 37 46
c80 22 0 1.66928e-19 $X=0.65 $Y=1.69
r81 37 59 4.37134 $w=2.88e-07 $l=1.1e-07 $layer=LI1_cond $X=2.17 $Y=2.775
+ $X2=2.17 $Y2=2.885
r82 37 55 9.53746 $w=2.88e-07 $l=2.4e-07 $layer=LI1_cond $X=2.17 $Y=2.775
+ $X2=2.17 $Y2=2.535
r83 36 47 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.45 $X2=2.17
+ $Y2=2.365
r84 36 55 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.45 $X2=2.17
+ $Y2=2.535
r85 36 47 0.914007 $w=2.88e-07 $l=2.3e-08 $layer=LI1_cond $X=2.17 $Y=2.342
+ $X2=2.17 $Y2=2.365
r86 35 36 12.2 $w=2.88e-07 $l=3.07e-07 $layer=LI1_cond $X=2.17 $Y=2.035 $X2=2.17
+ $Y2=2.342
r87 34 35 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=1.665
+ $X2=2.17 $Y2=2.035
r88 33 34 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=1.295
+ $X2=2.17 $Y2=1.665
r89 33 46 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=2.17 $Y=1.295
+ $X2=2.17 $Y2=1.015
r90 32 46 2.78474 $w=2.9e-07 $l=8.8e-08 $layer=LI1_cond $X=2.17 $Y=0.927
+ $X2=2.17 $Y2=1.015
r91 30 32 4.58849 $w=1.75e-07 $l=1.45e-07 $layer=LI1_cond $X=2.025 $Y=0.927
+ $X2=2.17 $Y2=0.927
r92 30 31 31.6883 $w=1.73e-07 $l=5e-07 $layer=LI1_cond $X=2.025 $Y=0.927
+ $X2=1.525 $Y2=0.927
r93 26 31 7.44913 $w=1.75e-07 $l=1.88547e-07 $layer=LI1_cond $X=1.375 $Y=0.84
+ $X2=1.525 $Y2=0.927
r94 26 28 16.1342 $w=2.98e-07 $l=4.2e-07 $layer=LI1_cond $X=1.375 $Y=0.84
+ $X2=1.375 $Y2=0.42
r95 24 36 3.3199 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.025 $Y=2.45
+ $X2=2.17 $Y2=2.45
r96 24 25 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=2.025 $Y=2.45
+ $X2=0.815 $Y2=2.45
r97 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.65
+ $Y=1.69 $X2=0.65 $Y2=1.69
r98 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.65 $Y=2.365
+ $X2=0.815 $Y2=2.45
r99 19 21 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.65 $Y=2.365
+ $X2=0.65 $Y2=1.69
r100 17 22 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=0.65 $Y=2.065
+ $X2=0.65 $Y2=1.69
r101 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=2.065
+ $X2=0.65 $Y2=2.23
r102 16 22 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=1.525
+ $X2=0.65 $Y2=1.69
r103 13 18 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.74 $Y=2.885
+ $X2=0.74 $Y2=2.23
r104 9 16 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=0.715 $Y=0.445
+ $X2=0.715 $Y2=1.525
r105 2 59 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=2.675 $X2=2.14 $Y2=2.885
r106 1 28 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.22
+ $Y=0.235 $X2=1.36 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUSHOLD0_1%RESET 3 7 11 12 13 14 18
r40 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=1.665
+ $X2=1.19 $Y2=2.035
r41 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.19
+ $Y=1.69 $X2=1.19 $Y2=1.69
r42 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.19 $Y=2.03
+ $X2=1.19 $Y2=1.69
r43 11 12 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=2.03
+ $X2=1.19 $Y2=2.195
r44 10 18 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.525
+ $X2=1.19 $Y2=1.69
r45 7 12 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.215 $Y=2.885
+ $X2=1.215 $Y2=2.195
r46 3 10 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=1.145 $Y=0.445
+ $X2=1.145 $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__BUSHOLD0_1%A_27_535# 1 2 7 9 10 12 14 21 23 25 27 33
+ 35 36 40
c64 23 0 1.66928e-19 $X=1.605 $Y=1.27
r65 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.35 $X2=1.73 $Y2=1.35
r66 35 36 6.80499 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.255 $Y=2.885
+ $X2=0.255 $Y2=2.72
r67 32 33 7.71634 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=0.48 $Y=1.205
+ $X2=0.625 $Y2=1.205
r68 30 32 10.7561 $w=2.98e-07 $l=2.8e-07 $layer=LI1_cond $X=0.2 $Y=1.205
+ $X2=0.48 $Y2=1.205
r69 28 40 86.939 $w=4.35e-07 $l=6.8e-07 $layer=POLY_cond $X=1.782 $Y=2.03
+ $X2=1.782 $Y2=1.35
r70 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=2.03 $X2=1.73 $Y2=2.03
r71 25 39 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=1.355
+ $X2=1.73 $Y2=1.27
r72 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.73 $Y=1.355
+ $X2=1.73 $Y2=2.03
r73 23 39 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.605 $Y=1.27
+ $X2=1.73 $Y2=1.27
r74 23 33 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=1.605 $Y=1.27
+ $X2=0.625 $Y2=1.27
r75 19 32 0.922372 $w=2.9e-07 $l=1.5e-07 $layer=LI1_cond $X=0.48 $Y=1.055
+ $X2=0.48 $Y2=1.205
r76 19 21 25.2345 $w=2.88e-07 $l=6.35e-07 $layer=LI1_cond $X=0.48 $Y=1.055
+ $X2=0.48 $Y2=0.42
r77 17 30 2.29563 $w=2.3e-07 $l=1.5e-07 $layer=LI1_cond $X=0.2 $Y=1.355 $X2=0.2
+ $Y2=1.205
r78 17 36 68.395 $w=2.28e-07 $l=1.365e-06 $layer=LI1_cond $X=0.2 $Y=1.355
+ $X2=0.2 $Y2=2.72
r79 16 28 47.9443 $w=4.35e-07 $l=3.75e-07 $layer=POLY_cond $X=1.782 $Y=2.405
+ $X2=1.782 $Y2=2.03
r80 14 40 47.9443 $w=4.35e-07 $l=3.75e-07 $layer=POLY_cond $X=1.782 $Y=0.975
+ $X2=1.782 $Y2=1.35
r81 10 16 27.7985 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.75 $Y=2.655 $X2=1.75
+ $Y2=2.405
r82 10 12 22.172 $w=5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.75 $Y=2.655 $X2=1.75
+ $Y2=2.885
r83 7 14 27.7985 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.75 $Y=0.725 $X2=1.75
+ $Y2=0.975
r84 7 9 26.992 $w=5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.75 $Y=0.725 $X2=1.75
+ $Y2=0.445
r85 2 35 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.675 $X2=0.26 $Y2=2.885
r86 1 21 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.375
+ $Y=0.235 $X2=0.5 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUSHOLD0_1%VPWR 1 6 9 10 11 21 22 28
r25 22 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.44 $Y2=3.33
r26 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 18 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r28 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 11 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.44 $Y2=3.33
r30 11 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 11 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 9 14 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=3.33 $X2=1
+ $Y2=3.33
r34 8 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.165 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=3.33 $X2=1
+ $Y2=3.33
r36 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=3.33
r37 4 6 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=2.885
r38 1 6 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=0.815
+ $Y=2.675 $X2=1 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__BUSHOLD0_1%VGND 1 2 9 11 13 16 17 18 24 30 35
r28 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r29 27 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r30 27 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.44
+ $Y2=0
r31 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r32 24 29 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.187
+ $Y2=0
r33 24 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.68
+ $Y2=0
r34 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r35 18 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.44
+ $Y2=0
r36 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r37 16 21 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.72
+ $Y2=0
r38 16 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.925
+ $Y2=0
r39 15 26 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.68
+ $Y2=0
r40 15 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.925
+ $Y2=0
r41 11 29 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.187 $Y2=0
r42 11 13 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.445
r43 7 17 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=0.085
+ $X2=0.925 $Y2=0
r44 7 9 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.925 $Y=0.085
+ $X2=0.925 $Y2=0.445
r45 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.235 $X2=2.14 $Y2=0.445
r46 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.79
+ $Y=0.235 $X2=0.93 $Y2=0.445
.ends

