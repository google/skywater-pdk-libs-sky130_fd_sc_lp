* File: sky130_fd_sc_lp__o21ba_4.spice
* Created: Wed Sep  2 10:16:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ba_4.pex.spice"
.subckt sky130_fd_sc_lp__o21ba_4  VNB VPB B1_N A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_B1_N_M1020_g N_A_37_49#_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=2.856 M=1 R=5.6 SA=75000.2
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1020_d N_A_180_23#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_180_23#_M1009_g N_X_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1009_d N_A_180_23#_M1016_g N_X_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1019_d N_A_180_23#_M1019_g N_X_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_575_65#_M1001_d N_A_37_49#_M1001_g N_A_180_23#_M1001_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.2898 AS=0.1176 PD=2.37 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6
+ SA=75000.3 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1013 N_A_575_65#_M1013_d N_A_37_49#_M1013_g N_A_180_23#_M1001_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6
+ SA=75000.7 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A1_M1005_g N_A_575_65#_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1512 PD=1.2 PS=1.2 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1012 N_A_575_65#_M1012_d N_A2_M1012_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=1.428 M=1 R=5.6 SA=75001.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1017 N_A_575_65#_M1012_d N_A2_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1017_s N_A1_M1008_g N_A_575_65#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=2.856 M=1 R=5.6 SA=75002.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_VPWR_M1021_d N_B1_N_M1021_g N_A_37_49#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.3 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1021_d N_A_180_23#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.8 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A_180_23#_M1002_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.17955 AS=0.1764 PD=1.545 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.4 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1002_d N_A_180_23#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.17955 AS=0.1764 PD=1.545 PS=1.54 NRD=0.7683 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75004 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_A_180_23#_M1018_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.41265 AS=0.1764 PD=1.915 PS=1.54 NRD=58.6272 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1006 N_A_180_23#_M1006_d N_A_37_49#_M1006_g N_VPWR_M1018_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.41265 PD=1.54 PS=1.915 NRD=0 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1011 N_A_180_23#_M1006_d N_A_37_49#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3906 PD=1.54 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75003.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1011_s N_A1_M1010_g N_A_878_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3906 AS=0.1764 PD=1.88 PS=1.54 NRD=35.4206 NRS=0 M=1 R=8.4
+ SA=75003.9 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1004 N_A_180_23#_M1004_d N_A2_M1004_g N_A_878_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.4
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1015 N_A_180_23#_M1004_d N_A2_M1015_g N_A_878_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.8
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A1_M1014_g N_A_878_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3969 AS=0.1764 PD=3.15 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75005.2 SB=75000.2 A=0.189 P=2.82 MULT=1
DX22_noxref VNB VPB NWDIODE A=12.3463 P=16.97
*
.include "sky130_fd_sc_lp__o21ba_4.pxi.spice"
*
.ends
*
*
