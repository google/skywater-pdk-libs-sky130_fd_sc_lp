* File: sky130_fd_sc_lp__nand4_4.spice
* Created: Wed Sep  2 10:05:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4_4.pex.spice"
.subckt sky130_fd_sc_lp__nand4_4  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1001 N_A_27_65#_M1001_d N_D_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1011 N_A_27_65#_M1011_d N_D_M1011_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1023 N_A_27_65#_M1011_d N_D_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1031 N_A_27_65#_M1031_d N_D_M1031_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5 SB=75002
+ A=0.126 P=1.98 MULT=1
MM1006 N_A_27_65#_M1031_d N_C_M1006_g N_A_454_65#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1009 N_A_27_65#_M1009_d N_C_M1009_g N_A_454_65#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1018 N_A_27_65#_M1009_d N_C_M1018_g N_A_454_65#_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1030 N_A_27_65#_M1030_d N_C_M1030_g N_A_454_65#_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.3066 AS=0.1176 PD=2.41 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6
+ SA=75003.2 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1013 N_A_454_65#_M1013_d N_B_M1013_g N_A_843_67#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1014 N_A_454_65#_M1013_d N_B_M1014_g N_A_843_67#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1020 N_A_454_65#_M1020_d N_B_M1020_g N_A_843_67#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1026 N_A_454_65#_M1020_d N_B_M1026_g N_A_843_67#_M1026_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1004 N_A_843_67#_M1026_s N_A_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1005 N_A_843_67#_M1005_d N_A_M1005_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1024 N_A_843_67#_M1005_d N_A_M1024_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1025 N_A_843_67#_M1025_d N_A_M1025_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_D_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75007.2 A=0.189 P=2.82 MULT=1
MM1012 N_Y_M1000_d N_D_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75006.8 A=0.189 P=2.82 MULT=1
MM1019 N_Y_M1019_d N_D_M1019_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75006.4 A=0.189 P=2.82 MULT=1
MM1027 N_Y_M1019_d N_D_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2772 PD=1.54 PS=1.7 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75001.5
+ SB=75006 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_C_M1002_g N_VPWR_M1027_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2772 PD=1.54 PS=1.7 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75002.1
+ SB=75005.4 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1002_d N_C_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1016 N_Y_M1016_d N_C_M1016_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1028 N_Y_M1016_d N_C_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.4
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1010_d N_B_M1010_g N_VPWR_M1028_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.8
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1015 N_Y_M1010_d N_B_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1022 N_Y_M1022_d N_B_M1022_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1029 N_Y_M1022_d N_B_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4599 PD=1.54 PS=1.99 NRD=0 NRS=0 M=1 R=8.4 SA=75005.1
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4599 PD=1.54 PS=1.99 NRD=0 NRS=0 M=1 R=8.4 SA=75006 SB=75001.5
+ A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1003_d N_A_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.4
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1017 N_Y_M1017_d N_A_M1017_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1021 N_Y_M1017_d N_A_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75007.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.9271 P=20.81
*
.include "sky130_fd_sc_lp__nand4_4.pxi.spice"
*
.ends
*
*
