* File: sky130_fd_sc_lp__o32ai_lp.pxi.spice
* Created: Wed Sep  2 10:27:04 2020
* 
x_PM_SKY130_FD_SC_LP__O32AI_LP%B1 N_B1_M1008_g N_B1_M1009_g B1 N_B1_c_58_n
+ N_B1_c_59_n PM_SKY130_FD_SC_LP__O32AI_LP%B1
x_PM_SKY130_FD_SC_LP__O32AI_LP%B2 N_B2_M1000_g N_B2_c_85_n N_B2_M1003_g
+ N_B2_c_87_n N_B2_c_88_n B2 B2 PM_SKY130_FD_SC_LP__O32AI_LP%B2
x_PM_SKY130_FD_SC_LP__O32AI_LP%A3 N_A3_M1002_g N_A3_M1005_g N_A3_c_130_n
+ N_A3_c_131_n A3 A3 A3 PM_SKY130_FD_SC_LP__O32AI_LP%A3
x_PM_SKY130_FD_SC_LP__O32AI_LP%A2 N_A2_c_170_n N_A2_M1004_g N_A2_M1006_g A2 A2
+ A2 N_A2_c_172_n PM_SKY130_FD_SC_LP__O32AI_LP%A2
x_PM_SKY130_FD_SC_LP__O32AI_LP%A1 N_A1_c_211_n N_A1_M1001_g N_A1_c_207_n
+ N_A1_M1007_g N_A1_c_208_n A1 N_A1_c_209_n N_A1_c_210_n
+ PM_SKY130_FD_SC_LP__O32AI_LP%A1
x_PM_SKY130_FD_SC_LP__O32AI_LP%VPWR N_VPWR_M1008_s N_VPWR_M1001_d N_VPWR_c_239_n
+ N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n VPWR N_VPWR_c_243_n
+ N_VPWR_c_238_n PM_SKY130_FD_SC_LP__O32AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O32AI_LP%Y N_Y_M1009_d N_Y_M1000_d N_Y_c_278_n N_Y_c_279_n
+ Y Y Y N_Y_c_288_n PM_SKY130_FD_SC_LP__O32AI_LP%Y
x_PM_SKY130_FD_SC_LP__O32AI_LP%A_27_179# N_A_27_179#_M1009_s N_A_27_179#_M1003_d
+ N_A_27_179#_M1006_d N_A_27_179#_c_315_n N_A_27_179#_c_316_n
+ N_A_27_179#_c_317_n N_A_27_179#_c_330_n N_A_27_179#_c_318_n
+ N_A_27_179#_c_319_n N_A_27_179#_c_320_n PM_SKY130_FD_SC_LP__O32AI_LP%A_27_179#
x_PM_SKY130_FD_SC_LP__O32AI_LP%VGND N_VGND_M1005_d N_VGND_M1007_d N_VGND_c_363_n
+ N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n VGND
+ N_VGND_c_368_n N_VGND_c_369_n PM_SKY130_FD_SC_LP__O32AI_LP%VGND
cc_1 VNB N_B1_M1009_g 0.0274037f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.105
cc_2 VNB N_B1_c_58_n 0.019001f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.68
cc_3 VNB N_B1_c_59_n 0.0068445f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.68
cc_4 VNB N_B2_c_85_n 0.0186679f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.105
cc_5 VNB N_B2_M1003_g 0.0261366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_B2_c_87_n 0.021381f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_B2_c_88_n 0.0472993f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.68
cc_8 VNB B2 0.00878649f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.515
cc_9 VNB N_A3_M1005_g 0.0384317f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.105
cc_10 VNB N_A3_c_130_n 0.0017016f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.68
cc_11 VNB N_A3_c_131_n 0.0104816f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.68
cc_12 VNB N_A2_c_170_n 0.0135183f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.845
cc_13 VNB N_A2_M1006_g 0.034055f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.105
cc_14 VNB N_A2_c_172_n 5.20105e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_207_n 0.020629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_208_n 0.00163053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_209_n 0.0651369f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.515
cc_18 VNB N_A1_c_210_n 0.00449722f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.845
cc_19 VNB N_VPWR_c_238_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_278_n 0.00251073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_279_n 0.00434925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_179#_c_315_n 0.019484f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.68
cc_23 VNB N_A_27_179#_c_316_n 0.00943756f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.515
cc_24 VNB N_A_27_179#_c_317_n 0.0130133f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.845
cc_25 VNB N_A_27_179#_c_318_n 0.0379435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_179#_c_319_n 0.00560076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_179#_c_320_n 0.00421379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_363_n 0.0305835f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_VGND_c_364_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.68
cc_30 VNB N_VGND_c_365_n 0.0608511f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.68
cc_31 VNB N_VGND_c_366_n 0.0540508f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.68
cc_32 VNB N_VGND_c_367_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_368_n 0.0207211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_369_n 0.225386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_B1_M1008_g 0.0399526f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_36 VPB N_B1_c_58_n 0.0203941f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.68
cc_37 VPB N_B1_c_59_n 0.00893009f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.68
cc_38 VPB N_B2_M1000_g 0.0389353f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_39 VPB N_B2_c_85_n 5.74677e-19 $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.105
cc_40 VPB N_A3_M1002_g 0.0258996f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_41 VPB N_A3_c_131_n 0.0257837f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.68
cc_42 VPB A3 0.00108113f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.845
cc_43 VPB N_A2_c_170_n 0.0232121f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.845
cc_44 VPB N_A2_M1004_g 0.025337f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_45 VPB N_A2_c_172_n 0.00478701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A1_c_211_n 0.0175754f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.845
cc_47 VPB N_A1_c_208_n 0.03743f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A1_c_210_n 0.0110506f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.845
cc_49 VPB N_VPWR_c_239_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.105
cc_50 VPB N_VPWR_c_240_n 0.0443603f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_51 VPB N_VPWR_c_241_n 0.0127321f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.68
cc_52 VPB N_VPWR_c_242_n 0.0442179f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.845
cc_53 VPB N_VPWR_c_243_n 0.0679766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_238_n 0.0474307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_Y_c_278_n 0.0018251f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB Y 0.0102985f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.68
cc_57 N_B1_M1008_g N_B2_M1000_g 0.0454261f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_58 N_B1_c_58_n N_B2_c_85_n 0.0466158f $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_59 N_B1_c_59_n N_B2_c_85_n 2.98958e-19 $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_60 N_B1_M1009_g N_B2_M1003_g 0.01738f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_61 N_B1_M1008_g N_VPWR_c_240_n 0.0284937f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_62 N_B1_c_58_n N_VPWR_c_240_n 0.00327168f $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_63 N_B1_c_59_n N_VPWR_c_240_n 0.0219892f $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_64 N_B1_M1008_g N_VPWR_c_243_n 0.008763f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_65 N_B1_M1008_g N_VPWR_c_238_n 0.0144563f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_66 N_B1_M1009_g N_Y_c_278_n 0.00386428f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_67 N_B1_c_58_n N_Y_c_278_n 0.00385431f $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_68 N_B1_c_59_n N_Y_c_278_n 0.0244136f $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_69 N_B1_M1009_g N_Y_c_279_n 0.00439122f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_70 N_B1_c_58_n N_Y_c_279_n 8.54694e-19 $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_71 N_B1_M1008_g Y 0.00494099f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_72 N_B1_M1008_g N_Y_c_288_n 0.00236978f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_73 N_B1_M1009_g N_A_27_179#_c_315_n 0.00830146f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_74 N_B1_c_58_n N_A_27_179#_c_315_n 0.00398952f $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_75 N_B1_c_59_n N_A_27_179#_c_315_n 0.0261276f $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_76 N_B1_M1009_g N_A_27_179#_c_316_n 0.0128771f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_77 N_B1_c_59_n N_A_27_179#_c_316_n 0.00331855f $X=0.44 $Y=1.68 $X2=0 $Y2=0
cc_78 N_B1_M1009_g N_VGND_c_366_n 4.9181e-19 $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_79 N_B2_M1000_g N_A3_M1002_g 0.018876f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_80 N_B2_c_85_n N_A3_M1005_g 0.00783666f $X=1.005 $Y=1.39 $X2=0 $Y2=0
cc_81 N_B2_M1003_g N_A3_M1005_g 0.0154301f $X=1.005 $Y=1.105 $X2=0 $Y2=0
cc_82 N_B2_c_87_n N_A3_M1005_g 0.00215099f $X=1.565 $Y=0.41 $X2=0 $Y2=0
cc_83 B2 N_A3_M1005_g 0.0163637f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_84 N_B2_c_85_n N_A3_c_130_n 0.00116738f $X=1.005 $Y=1.39 $X2=0 $Y2=0
cc_85 N_B2_c_85_n N_A3_c_131_n 0.018876f $X=1.005 $Y=1.39 $X2=0 $Y2=0
cc_86 N_B2_M1000_g A3 4.79811e-19 $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_87 N_B2_M1000_g N_VPWR_c_240_n 0.0036637f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_88 N_B2_M1000_g N_VPWR_c_243_n 0.00864331f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_89 N_B2_M1000_g N_VPWR_c_238_n 0.0142996f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_90 N_B2_M1000_g N_Y_c_278_n 0.00692089f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_91 N_B2_c_85_n N_Y_c_278_n 0.00775642f $X=1.005 $Y=1.39 $X2=0 $Y2=0
cc_92 N_B2_M1003_g N_Y_c_278_n 9.49841e-19 $X=1.005 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B2_M1003_g N_Y_c_279_n 0.00320124f $X=1.005 $Y=1.105 $X2=0 $Y2=0
cc_94 N_B2_M1000_g Y 0.0275589f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_95 N_B2_M1000_g N_Y_c_288_n 0.0226292f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_96 N_B2_M1003_g N_A_27_179#_c_316_n 0.015002f $X=1.005 $Y=1.105 $X2=0 $Y2=0
cc_97 N_B2_c_87_n N_A_27_179#_c_316_n 0.0330485f $X=1.565 $Y=0.41 $X2=0 $Y2=0
cc_98 N_B2_c_88_n N_A_27_179#_c_316_n 0.0042163f $X=1.095 $Y=0.41 $X2=0 $Y2=0
cc_99 B2 N_A_27_179#_c_316_n 0.013154f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_100 B2 N_A_27_179#_c_330_n 0.00951906f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_101 B2 N_A_27_179#_c_318_n 0.013058f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_102 N_B2_c_85_n N_A_27_179#_c_319_n 0.00232395f $X=1.005 $Y=1.39 $X2=0 $Y2=0
cc_103 N_B2_M1003_g N_A_27_179#_c_319_n 0.00113138f $X=1.005 $Y=1.105 $X2=0
+ $Y2=0
cc_104 B2 N_VGND_M1005_d 0.00341692f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_105 B2 N_VGND_c_363_n 0.060276f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_106 N_B2_c_87_n N_VGND_c_366_n 0.0389212f $X=1.565 $Y=0.41 $X2=0 $Y2=0
cc_107 N_B2_c_88_n N_VGND_c_366_n 0.00582385f $X=1.095 $Y=0.41 $X2=0 $Y2=0
cc_108 B2 N_VGND_c_366_n 0.0155076f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_109 N_B2_c_87_n N_VGND_c_369_n 0.0225036f $X=1.565 $Y=0.41 $X2=0 $Y2=0
cc_110 N_B2_c_88_n N_VGND_c_369_n 0.0112336f $X=1.095 $Y=0.41 $X2=0 $Y2=0
cc_111 B2 N_VGND_c_369_n 0.00889943f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_112 N_A3_M1005_g N_A2_c_170_n 0.00217489f $X=1.595 $Y=0.975 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A3_c_130_n N_A2_c_170_n 4.06548e-19 $X=1.66 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A3_c_131_n N_A2_c_170_n 0.0177499f $X=1.66 $Y=1.77 $X2=-0.19 $Y2=-0.245
cc_115 N_A3_M1002_g N_A2_M1004_g 0.0417994f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_116 A3 N_A2_M1004_g 0.00346436f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_117 N_A3_M1005_g N_A2_M1006_g 0.0149257f $X=1.595 $Y=0.975 $X2=0 $Y2=0
cc_118 N_A3_M1002_g N_A2_c_172_n 0.00100552f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_119 N_A3_c_130_n N_A2_c_172_n 0.0579764f $X=1.66 $Y=1.77 $X2=0 $Y2=0
cc_120 N_A3_c_131_n N_A2_c_172_n 0.00206081f $X=1.66 $Y=1.77 $X2=0 $Y2=0
cc_121 N_A3_M1002_g N_VPWR_c_243_n 0.00816902f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_122 A3 N_VPWR_c_243_n 0.00712674f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_123 N_A3_M1002_g N_VPWR_c_238_n 0.0128987f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_124 A3 N_VPWR_c_238_n 0.0083777f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_125 N_A3_M1005_g N_Y_c_278_n 7.46202e-19 $X=1.595 $Y=0.975 $X2=0 $Y2=0
cc_126 N_A3_c_130_n N_Y_c_278_n 0.00869001f $X=1.66 $Y=1.77 $X2=0 $Y2=0
cc_127 N_A3_c_131_n N_Y_c_278_n 9.41867e-19 $X=1.66 $Y=1.77 $X2=0 $Y2=0
cc_128 N_A3_c_130_n Y 0.0011869f $X=1.66 $Y=1.77 $X2=0 $Y2=0
cc_129 N_A3_c_131_n Y 0.00154769f $X=1.66 $Y=1.77 $X2=0 $Y2=0
cc_130 A3 Y 0.0108083f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_131 A3 A_338_419# 0.0087259f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_132 N_A3_M1005_g N_A_27_179#_c_316_n 0.00148618f $X=1.595 $Y=0.975 $X2=0
+ $Y2=0
cc_133 N_A3_M1005_g N_A_27_179#_c_330_n 0.0059999f $X=1.595 $Y=0.975 $X2=0 $Y2=0
cc_134 N_A3_M1005_g N_A_27_179#_c_318_n 0.0137851f $X=1.595 $Y=0.975 $X2=0 $Y2=0
cc_135 N_A3_c_130_n N_A_27_179#_c_318_n 0.0242419f $X=1.66 $Y=1.77 $X2=0 $Y2=0
cc_136 N_A3_c_131_n N_A_27_179#_c_318_n 0.00353467f $X=1.66 $Y=1.77 $X2=0 $Y2=0
cc_137 N_A3_M1005_g N_VGND_c_363_n 0.00163842f $X=1.595 $Y=0.975 $X2=0 $Y2=0
cc_138 N_A3_M1005_g N_VGND_c_366_n 3.33119e-19 $X=1.595 $Y=0.975 $X2=0 $Y2=0
cc_139 N_A2_M1006_g N_A1_c_207_n 0.0156621f $X=2.355 $Y=0.975 $X2=0 $Y2=0
cc_140 N_A2_c_170_n N_A1_c_208_n 0.00950193f $X=2.19 $Y=1.935 $X2=0 $Y2=0
cc_141 N_A2_M1004_g N_A1_c_208_n 0.0487487f $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_142 N_A2_c_172_n N_A1_c_208_n 0.0106728f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_143 N_A2_c_170_n N_A1_c_209_n 0.0156621f $X=2.19 $Y=1.935 $X2=0 $Y2=0
cc_144 N_A2_c_172_n N_A1_c_209_n 0.00159981f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_145 N_A2_M1006_g N_A1_c_210_n 9.19382e-19 $X=2.355 $Y=0.975 $X2=0 $Y2=0
cc_146 N_A2_c_172_n N_A1_c_210_n 0.00589673f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_147 N_A2_M1004_g N_VPWR_c_242_n 0.00238619f $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_148 N_A2_c_172_n N_VPWR_c_242_n 0.0291824f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_149 N_A2_M1004_g N_VPWR_c_243_n 0.00655603f $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_150 N_A2_c_172_n N_VPWR_c_243_n 0.00949589f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_151 N_A2_M1004_g N_VPWR_c_238_n 0.00859421f $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_152 N_A2_c_172_n N_VPWR_c_238_n 0.0108878f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_153 N_A2_c_172_n A_463_419# 0.0109985f $X=2.23 $Y=1.77 $X2=-0.19 $Y2=-0.245
cc_154 N_A2_c_170_n N_A_27_179#_c_318_n 0.00599723f $X=2.19 $Y=1.935 $X2=0 $Y2=0
cc_155 N_A2_M1006_g N_A_27_179#_c_318_n 0.0159777f $X=2.355 $Y=0.975 $X2=0 $Y2=0
cc_156 N_A2_c_172_n N_A_27_179#_c_318_n 0.0262831f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_157 N_A2_M1006_g N_A_27_179#_c_320_n 0.0132117f $X=2.355 $Y=0.975 $X2=0 $Y2=0
cc_158 N_A2_M1006_g N_VGND_c_363_n 0.00594303f $X=2.355 $Y=0.975 $X2=0 $Y2=0
cc_159 N_A2_M1006_g N_VGND_c_368_n 0.00337154f $X=2.355 $Y=0.975 $X2=0 $Y2=0
cc_160 N_A2_M1006_g N_VGND_c_369_n 0.00432409f $X=2.355 $Y=0.975 $X2=0 $Y2=0
cc_161 N_A1_c_211_n N_VPWR_c_242_n 0.0254448f $X=2.76 $Y=2.09 $X2=0 $Y2=0
cc_162 N_A1_c_208_n N_VPWR_c_242_n 0.00102331f $X=2.785 $Y=1.94 $X2=0 $Y2=0
cc_163 N_A1_c_209_n N_VPWR_c_242_n 0.00265427f $X=3.08 $Y=1.46 $X2=0 $Y2=0
cc_164 N_A1_c_210_n N_VPWR_c_242_n 0.016956f $X=3.08 $Y=1.46 $X2=0 $Y2=0
cc_165 N_A1_c_211_n N_VPWR_c_243_n 0.008763f $X=2.76 $Y=2.09 $X2=0 $Y2=0
cc_166 N_A1_c_211_n N_VPWR_c_238_n 0.0146671f $X=2.76 $Y=2.09 $X2=0 $Y2=0
cc_167 N_A1_c_207_n N_A_27_179#_c_318_n 0.00229462f $X=2.785 $Y=1.295 $X2=0
+ $Y2=0
cc_168 N_A1_c_208_n N_A_27_179#_c_318_n 0.00251218f $X=2.785 $Y=1.94 $X2=0 $Y2=0
cc_169 N_A1_c_209_n N_A_27_179#_c_318_n 0.00504051f $X=3.08 $Y=1.46 $X2=0 $Y2=0
cc_170 N_A1_c_210_n N_A_27_179#_c_318_n 0.00990958f $X=3.08 $Y=1.46 $X2=0 $Y2=0
cc_171 N_A1_c_207_n N_A_27_179#_c_320_n 0.0119146f $X=2.785 $Y=1.295 $X2=0 $Y2=0
cc_172 N_A1_c_207_n N_VGND_c_365_n 0.011778f $X=2.785 $Y=1.295 $X2=0 $Y2=0
cc_173 N_A1_c_209_n N_VGND_c_365_n 0.00257359f $X=3.08 $Y=1.46 $X2=0 $Y2=0
cc_174 N_A1_c_210_n N_VGND_c_365_n 0.0267429f $X=3.08 $Y=1.46 $X2=0 $Y2=0
cc_175 N_A1_c_207_n N_VGND_c_368_n 0.00337154f $X=2.785 $Y=1.295 $X2=0 $Y2=0
cc_176 N_A1_c_207_n N_VGND_c_369_n 0.00432409f $X=2.785 $Y=1.295 $X2=0 $Y2=0
cc_177 N_VPWR_c_238_n A_134_419# 0.010279f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_178 N_VPWR_c_238_n N_Y_M1000_d 0.00415099f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_179 N_VPWR_c_240_n Y 0.00505797f $X=0.28 $Y=2.24 $X2=0 $Y2=0
cc_180 N_VPWR_c_240_n N_Y_c_288_n 0.0197492f $X=0.28 $Y=2.24 $X2=0 $Y2=0
cc_181 N_VPWR_c_243_n N_Y_c_288_n 0.0176125f $X=2.86 $Y=3.33 $X2=0 $Y2=0
cc_182 N_VPWR_c_238_n N_Y_c_288_n 0.0111115f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_238_n A_338_419# 0.0109044f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_184 N_VPWR_c_238_n A_463_419# 0.0110428f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_185 N_Y_c_279_n N_A_27_179#_c_315_n 0.00971956f $X=0.79 $Y=1.17 $X2=0 $Y2=0
cc_186 N_Y_M1009_d N_A_27_179#_c_316_n 0.00180746f $X=0.65 $Y=0.895 $X2=0 $Y2=0
cc_187 N_Y_c_279_n N_A_27_179#_c_316_n 0.0157582f $X=0.79 $Y=1.17 $X2=0 $Y2=0
cc_188 N_Y_c_279_n N_A_27_179#_c_319_n 0.010462f $X=0.79 $Y=1.17 $X2=0 $Y2=0
cc_189 Y N_A_27_179#_c_319_n 0.00778508f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_190 N_A_27_179#_c_330_n N_VGND_c_363_n 0.00105828f $X=1.3 $Y=1.04 $X2=0 $Y2=0
cc_191 N_A_27_179#_c_318_n N_VGND_c_363_n 0.0196257f $X=2.405 $Y=1.34 $X2=0
+ $Y2=0
cc_192 N_A_27_179#_c_320_n N_VGND_c_363_n 0.0125556f $X=2.57 $Y=0.975 $X2=0
+ $Y2=0
cc_193 N_A_27_179#_c_320_n N_VGND_c_365_n 0.0140205f $X=2.57 $Y=0.975 $X2=0
+ $Y2=0
cc_194 N_A_27_179#_c_316_n N_VGND_c_366_n 0.00722746f $X=1.135 $Y=0.82 $X2=0
+ $Y2=0
cc_195 N_A_27_179#_c_317_n N_VGND_c_366_n 0.00544512f $X=0.445 $Y=0.82 $X2=0
+ $Y2=0
cc_196 N_A_27_179#_c_320_n N_VGND_c_368_n 0.00526067f $X=2.57 $Y=0.975 $X2=0
+ $Y2=0
cc_197 N_A_27_179#_c_316_n N_VGND_c_369_n 0.0131227f $X=1.135 $Y=0.82 $X2=0
+ $Y2=0
cc_198 N_A_27_179#_c_317_n N_VGND_c_369_n 0.00924242f $X=0.445 $Y=0.82 $X2=0
+ $Y2=0
cc_199 N_A_27_179#_c_320_n N_VGND_c_369_n 0.00911247f $X=2.57 $Y=0.975 $X2=0
+ $Y2=0
