* File: sky130_fd_sc_lp__dlrtn_lp.spice
* Created: Wed Sep  2 09:47:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrtn_lp.pex.spice"
.subckt sky130_fd_sc_lp__dlrtn_lp  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1003 A_114_47# N_D_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_D_M1019_g A_114_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1004 A_272_47# N_GATE_N_M1004_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_264_415#_M1005_d N_GATE_N_M1005_g A_272_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 A_554_47# N_A_264_415#_M1018_g N_A_399_415#_M1018_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_264_415#_M1010_g A_554_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1022 A_712_47# N_A_27_47#_M1022_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1020 N_A_744_415#_M1020_d N_A_264_415#_M1020_g A_712_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=31.428 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1007 A_898_47# N_A_399_415#_M1007_g N_A_744_415#_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.0819 PD=0.84 PS=0.81 NRD=44.28 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_949_335#_M1013_g A_898_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1449 AS=0.0882 PD=1.53 PS=0.84 NRD=17.136 NRS=44.28 M=1 R=2.8 SA=75002.5
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1001 A_1222_57# N_A_744_415#_M1001_g N_A_949_335#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_RESET_B_M1006_g A_1222_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1011 A_1380_57# N_A_949_335#_M1011_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_Q_M1014_d N_A_949_335#_M1014_g A_1380_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_27_47#_M1000_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1012 N_A_264_415#_M1012_d N_GATE_N_M1012_g N_VPWR_M1000_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1015 N_VPWR_M1015_d N_A_264_415#_M1015_g N_A_399_415#_M1015_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.225 AS=0.285 PD=1.45 PS=2.57 NRD=33.4703 NRS=0 M=1 R=4
+ SA=125000 SB=125005 A=0.25 P=2.5 MULT=1
MM1016 A_646_415# N_A_27_47#_M1016_g N_VPWR_M1015_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.225 PD=1.24 PS=1.45 NRD=12.7853 NRS=0 M=1 R=4 SA=125001 SB=125004
+ A=0.25 P=2.5 MULT=1
MM1002 N_A_744_415#_M1002_d N_A_399_415#_M1002_g A_646_415# VPB PHIGHVT L=0.25
+ W=1 AD=0.2675 AS=0.12 PD=1.535 PS=1.24 NRD=50.2153 NRS=12.7853 M=1 R=4
+ SA=125001 SB=125003 A=0.25 P=2.5 MULT=1
MM1023 A_901_415# N_A_264_415#_M1023_g N_A_744_415#_M1002_d VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.2675 PD=1.24 PS=1.535 NRD=12.7853 NRS=0 M=1 R=4 SA=125002
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A_949_335#_M1009_g A_901_415# VPB PHIGHVT L=0.25 W=1
+ AD=0.3225 AS=0.12 PD=1.645 PS=1.24 NRD=40.3653 NRS=12.7853 M=1 R=4 SA=125003
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1021 N_A_949_335#_M1021_d N_A_744_415#_M1021_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.3225 PD=1.28 PS=1.645 NRD=0 NRS=31.5003 M=1 R=4
+ SA=125004 SB=125001 A=0.25 P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_RESET_B_M1008_g N_A_949_335#_M1021_d VPB PHIGHVT L=0.25
+ W=1 AD=0.1925 AS=0.14 PD=1.385 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1017 N_Q_M1017_d N_A_949_335#_M1017_g N_VPWR_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.1925 PD=2.57 PS=1.385 NRD=0 NRS=20.685 M=1 R=4 SA=125005
+ SB=125000 A=0.25 P=2.5 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.0319 P=19.85
*
.include "sky130_fd_sc_lp__dlrtn_lp.pxi.spice"
*
.ends
*
*
