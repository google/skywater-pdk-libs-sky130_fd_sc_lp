* File: sky130_fd_sc_lp__a31o_2.spice
* Created: Wed Sep  2 09:26:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a31o_2.pex.spice"
.subckt sky130_fd_sc_lp__a31o_2  VNB VPB A3 A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_85_23#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_85_23#_M1009_g N_X_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1006 A_355_49# N_A3_M1006_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.2604 PD=1.05 PS=1.46 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001.4 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1004 A_427_49# N_A2_M1004_g A_355_49# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75001.7 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1011 N_A_85_23#_M1011_d N_A1_M1011_g A_427_49# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=5.712 NRS=19.992 M=1 R=5.6 SA=75002.3
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_B1_M1000_g N_A_85_23#_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_85_23#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4725 AS=0.1764 PD=3.27 PS=1.54 NRD=17.1981 NRS=0 M=1 R=8.4 SA=75000.3
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A_85_23#_M1007_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=7.0329 NRS=0 M=1 R=8.4 SA=75000.7
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1003 N_A_342_367#_M1003_d N_A3_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2268 PD=1.54 PS=1.62 NRD=0 NRS=5.4569 M=1 R=8.4
+ SA=75001.2 SB=75001.7 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_342_367#_M1003_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.31185 AS=0.1764 PD=1.755 PS=1.54 NRD=17.1981 NRS=0 M=1 R=8.4
+ SA=75001.7 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1001 N_A_342_367#_M1001_d N_A1_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.31185 PD=1.54 PS=1.755 NRD=0 NRS=16.4101 M=1 R=8.4
+ SA=75002.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_A_85_23#_M1010_d N_B1_M1010_g N_A_342_367#_M1001_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a31o_2.pxi.spice"
*
.ends
*
*
