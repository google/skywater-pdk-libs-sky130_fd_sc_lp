* File: sky130_fd_sc_lp__xor3_1.pxi.spice
* Created: Wed Sep  2 10:41:45 2020
* 
x_PM_SKY130_FD_SC_LP__XOR3_1%A_86_305# N_A_86_305#_M1004_d N_A_86_305#_M1021_d
+ N_A_86_305#_M1016_d N_A_86_305#_M1019_d N_A_86_305#_M1000_g
+ N_A_86_305#_M1007_g N_A_86_305#_c_182_n N_A_86_305#_c_183_n
+ N_A_86_305#_c_184_n N_A_86_305#_c_198_p N_A_86_305#_c_176_n
+ N_A_86_305#_c_186_n N_A_86_305#_c_187_n N_A_86_305#_c_177_n
+ N_A_86_305#_c_178_n N_A_86_305#_c_190_n N_A_86_305#_c_179_n
+ N_A_86_305#_c_180_n PM_SKY130_FD_SC_LP__XOR3_1%A_86_305#
x_PM_SKY130_FD_SC_LP__XOR3_1%A N_A_c_278_n N_A_M1004_g N_A_M1016_g A N_A_c_280_n
+ PM_SKY130_FD_SC_LP__XOR3_1%A
x_PM_SKY130_FD_SC_LP__XOR3_1%A_474_313# N_A_474_313#_M1005_s
+ N_A_474_313#_M1006_s N_A_474_313#_M1003_g N_A_474_313#_M1020_g
+ N_A_474_313#_c_318_n N_A_474_313#_c_319_n N_A_474_313#_M1019_g
+ N_A_474_313#_c_320_n N_A_474_313#_M1021_g N_A_474_313#_c_322_n
+ N_A_474_313#_c_323_n N_A_474_313#_c_393_p N_A_474_313#_c_324_n
+ N_A_474_313#_c_325_n N_A_474_313#_c_326_n N_A_474_313#_c_327_n
+ PM_SKY130_FD_SC_LP__XOR3_1%A_474_313#
x_PM_SKY130_FD_SC_LP__XOR3_1%B N_B_M1002_g N_B_M1018_g N_B_c_433_n N_B_c_434_n
+ N_B_c_419_n N_B_c_420_n N_B_M1013_g N_B_c_436_n N_B_M1010_g N_B_c_422_n
+ N_B_c_423_n N_B_c_424_n N_B_c_425_n N_B_M1005_g N_B_M1006_g N_B_c_439_n
+ N_B_c_427_n N_B_c_428_n B N_B_c_430_n N_B_c_431_n PM_SKY130_FD_SC_LP__XOR3_1%B
x_PM_SKY130_FD_SC_LP__XOR3_1%A_1263_295# N_A_1263_295#_M1015_s
+ N_A_1263_295#_M1008_s N_A_1263_295#_M1001_g N_A_1263_295#_M1017_g
+ N_A_1263_295#_c_540_n N_A_1263_295#_c_541_n N_A_1263_295#_c_542_n
+ N_A_1263_295#_c_550_n N_A_1263_295#_c_551_n N_A_1263_295#_c_552_n
+ N_A_1263_295#_c_543_n N_A_1263_295#_c_557_p N_A_1263_295#_c_544_n
+ N_A_1263_295#_c_545_n PM_SKY130_FD_SC_LP__XOR3_1%A_1263_295#
x_PM_SKY130_FD_SC_LP__XOR3_1%C N_C_c_612_n N_C_M1014_g N_C_M1011_g N_C_c_613_n
+ N_C_c_614_n N_C_M1008_g N_C_M1015_g N_C_c_617_n C PM_SKY130_FD_SC_LP__XOR3_1%C
x_PM_SKY130_FD_SC_LP__XOR3_1%A_1363_127# N_A_1363_127#_M1001_d
+ N_A_1363_127#_M1017_d N_A_1363_127#_M1012_g N_A_1363_127#_M1009_g
+ N_A_1363_127#_c_692_n N_A_1363_127#_c_682_n N_A_1363_127#_c_683_n
+ N_A_1363_127#_c_688_n N_A_1363_127#_c_689_n N_A_1363_127#_c_690_n
+ N_A_1363_127#_c_726_p N_A_1363_127#_c_684_n N_A_1363_127#_c_685_n
+ PM_SKY130_FD_SC_LP__XOR3_1%A_1363_127#
x_PM_SKY130_FD_SC_LP__XOR3_1%A_42_411# N_A_42_411#_M1007_s N_A_42_411#_M1020_d
+ N_A_42_411#_M1000_s N_A_42_411#_M1003_d N_A_42_411#_c_768_n
+ N_A_42_411#_c_758_n N_A_42_411#_c_759_n N_A_42_411#_c_760_n
+ N_A_42_411#_c_761_n N_A_42_411#_c_769_n N_A_42_411#_c_762_n
+ N_A_42_411#_c_763_n N_A_42_411#_c_764_n N_A_42_411#_c_770_n
+ N_A_42_411#_c_765_n N_A_42_411#_c_766_n N_A_42_411#_c_767_n
+ PM_SKY130_FD_SC_LP__XOR3_1%A_42_411#
x_PM_SKY130_FD_SC_LP__XOR3_1%VPWR N_VPWR_M1000_d N_VPWR_M1006_d N_VPWR_M1008_d
+ N_VPWR_c_842_n N_VPWR_c_843_n N_VPWR_c_844_n N_VPWR_c_845_n N_VPWR_c_846_n
+ VPWR N_VPWR_c_847_n N_VPWR_c_848_n N_VPWR_c_849_n N_VPWR_c_841_n
+ N_VPWR_c_851_n N_VPWR_c_852_n PM_SKY130_FD_SC_LP__XOR3_1%VPWR
x_PM_SKY130_FD_SC_LP__XOR3_1%A_402_411# N_A_402_411#_M1010_d
+ N_A_402_411#_M1001_s N_A_402_411#_M1002_d N_A_402_411#_M1011_d
+ N_A_402_411#_c_923_n N_A_402_411#_c_924_n N_A_402_411#_c_925_n
+ N_A_402_411#_c_915_n N_A_402_411#_c_916_n N_A_402_411#_c_917_n
+ N_A_402_411#_c_961_n N_A_402_411#_c_918_n N_A_402_411#_c_965_n
+ N_A_402_411#_c_919_n N_A_402_411#_c_920_n N_A_402_411#_c_921_n
+ N_A_402_411#_c_927_n N_A_402_411#_c_922_n N_A_402_411#_c_929_n
+ PM_SKY130_FD_SC_LP__XOR3_1%A_402_411#
x_PM_SKY130_FD_SC_LP__XOR3_1%A_425_117# N_A_425_117#_M1018_d
+ N_A_425_117#_M1014_d N_A_425_117#_M1013_d N_A_425_117#_M1017_s
+ N_A_425_117#_c_1044_n N_A_425_117#_c_1045_n N_A_425_117#_c_1046_n
+ N_A_425_117#_c_1047_n N_A_425_117#_c_1048_n N_A_425_117#_c_1100_n
+ N_A_425_117#_c_1049_n N_A_425_117#_c_1050_n N_A_425_117#_c_1051_n
+ N_A_425_117#_c_1054_n N_A_425_117#_c_1055_n N_A_425_117#_c_1056_n
+ N_A_425_117#_c_1057_n N_A_425_117#_c_1052_n N_A_425_117#_c_1053_n
+ PM_SKY130_FD_SC_LP__XOR3_1%A_425_117#
x_PM_SKY130_FD_SC_LP__XOR3_1%X N_X_M1012_d N_X_M1009_d X X X X X X X
+ N_X_c_1159_n X PM_SKY130_FD_SC_LP__XOR3_1%X
x_PM_SKY130_FD_SC_LP__XOR3_1%VGND N_VGND_M1007_d N_VGND_M1005_d N_VGND_M1015_d
+ N_VGND_c_1175_n N_VGND_c_1176_n N_VGND_c_1177_n N_VGND_c_1178_n
+ N_VGND_c_1179_n N_VGND_c_1180_n N_VGND_c_1181_n N_VGND_c_1182_n VGND
+ N_VGND_c_1183_n N_VGND_c_1184_n PM_SKY130_FD_SC_LP__XOR3_1%VGND
cc_1 VNB N_A_86_305#_M1007_g 0.0353243f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.905
cc_2 VNB N_A_86_305#_c_176_n 0.0103577f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.08
cc_3 VNB N_A_86_305#_c_177_n 0.00472196f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.69
cc_4 VNB N_A_86_305#_c_178_n 0.014133f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.69
cc_5 VNB N_A_86_305#_c_179_n 0.00826721f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=1.905
cc_6 VNB N_A_86_305#_c_180_n 0.00203835f $X=-0.19 $Y=-0.245 $X2=4.405 $Y2=1.05
cc_7 VNB N_A_c_278_n 0.0204237f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.585
cc_8 VNB A 0.00115257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_280_n 0.0402592f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.555
cc_10 VNB N_A_474_313#_M1020_g 0.0344309f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.855
cc_11 VNB N_A_474_313#_c_318_n 0.0260425f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.555
cc_12 VNB N_A_474_313#_c_319_n 0.011317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_474_313#_c_320_n 0.0176312f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.93
cc_14 VNB N_A_474_313#_M1021_g 0.0198876f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.2
cc_15 VNB N_A_474_313#_c_322_n 0.00867197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_474_313#_c_323_n 0.0082541f $X=-0.19 $Y=-0.245 $X2=3.975 $Y2=2.745
cc_17 VNB N_A_474_313#_c_324_n 0.00876201f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.69
cc_18 VNB N_A_474_313#_c_325_n 0.00141616f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=2.07
cc_19 VNB N_A_474_313#_c_326_n 0.0253394f $X=-0.19 $Y=-0.245 $X2=4.055 $Y2=2.07
cc_20 VNB N_A_474_313#_c_327_n 0.00121041f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=1.905
cc_21 VNB N_B_M1018_g 0.0367675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_419_n 0.0740407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_420_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_M1010_g 0.0323889f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.93
cc_25 VNB N_B_c_422_n 0.0965686f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.18
cc_26 VNB N_B_c_423_n 0.0560416f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.2
cc_27 VNB N_B_c_424_n 0.0177059f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.08
cc_28 VNB N_B_c_425_n 0.0216767f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=2.98
cc_29 VNB N_B_M1006_g 0.00589028f $X=-0.19 $Y=-0.245 $X2=4.485 $Y2=1.905
cc_30 VNB N_B_c_427_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.69
cc_31 VNB N_B_c_428_n 0.006715f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.93
cc_32 VNB B 0.0078889f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.93
cc_33 VNB N_B_c_430_n 0.0160093f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=2.07
cc_34 VNB N_B_c_431_n 0.0453933f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=1.905
cc_35 VNB N_A_1263_295#_M1001_g 0.0240691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1263_295#_c_540_n 0.0211268f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.555
cc_37 VNB N_A_1263_295#_c_541_n 0.00827405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1263_295#_c_542_n 0.0031385f $X=-0.19 $Y=-0.245 $X2=0.655
+ $Y2=0.905
cc_39 VNB N_A_1263_295#_c_543_n 0.00329236f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.08
cc_40 VNB N_A_1263_295#_c_544_n 0.00571536f $X=-0.19 $Y=-0.245 $X2=3.975
+ $Y2=2.895
cc_41 VNB N_A_1263_295#_c_545_n 0.00235704f $X=-0.19 $Y=-0.245 $X2=4.485
+ $Y2=1.215
cc_42 VNB N_C_c_612_n 0.018643f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.585
cc_43 VNB N_C_c_613_n 0.0494359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_C_c_614_n 0.0277487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_C_M1008_g 0.0074563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_C_M1015_g 0.0306034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_C_c_617_n 0.0170638f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.905
cc_48 VNB C 0.00194063f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.93
cc_49 VNB N_A_1363_127#_M1012_g 0.0286268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1363_127#_M1009_g 0.00116262f $X=-0.19 $Y=-0.245 $X2=0.57
+ $Y2=1.855
cc_51 VNB N_A_1363_127#_c_682_n 0.00747742f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.93
cc_52 VNB N_A_1363_127#_c_683_n 0.00548183f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.2
cc_53 VNB N_A_1363_127#_c_684_n 2.16116e-19 $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.69
cc_54 VNB N_A_1363_127#_c_685_n 0.0475929f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.98
cc_55 VNB N_A_42_411#_c_758_n 0.00944431f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.905
cc_56 VNB N_A_42_411#_c_759_n 0.00212149f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.93
cc_57 VNB N_A_42_411#_c_760_n 0.0142038f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.18
cc_58 VNB N_A_42_411#_c_761_n 0.00454642f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.895
cc_59 VNB N_A_42_411#_c_762_n 0.00124645f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.08
cc_60 VNB N_A_42_411#_c_763_n 0.00182846f $X=-0.19 $Y=-0.245 $X2=3.975 $Y2=2.745
cc_61 VNB N_A_42_411#_c_764_n 0.0460644f $X=-0.19 $Y=-0.245 $X2=3.975 $Y2=2.895
cc_62 VNB N_A_42_411#_c_765_n 0.0201952f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.93
cc_63 VNB N_A_42_411#_c_766_n 0.0028097f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.98
cc_64 VNB N_A_42_411#_c_767_n 0.00258861f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.9
cc_65 VNB N_VPWR_c_841_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_402_411#_c_915_n 0.00981412f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.93
cc_67 VNB N_A_402_411#_c_916_n 0.022486f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.18
cc_68 VNB N_A_402_411#_c_917_n 0.00291736f $X=-0.19 $Y=-0.245 $X2=1.605
+ $Y2=2.895
cc_69 VNB N_A_402_411#_c_918_n 0.00890163f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.845
cc_70 VNB N_A_402_411#_c_919_n 0.0104525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_402_411#_c_920_n 0.0461014f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=2.98
cc_72 VNB N_A_402_411#_c_921_n 0.00520639f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=2.98
cc_73 VNB N_A_402_411#_c_922_n 0.0248835f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.93
cc_74 VNB N_A_425_117#_c_1044_n 0.0133907f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.555
cc_75 VNB N_A_425_117#_c_1045_n 0.0214775f $X=-0.19 $Y=-0.245 $X2=0.655
+ $Y2=0.905
cc_76 VNB N_A_425_117#_c_1046_n 0.00465802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_425_117#_c_1047_n 0.00869045f $X=-0.19 $Y=-0.245 $X2=1.605
+ $Y2=2.18
cc_78 VNB N_A_425_117#_c_1048_n 0.00533345f $X=-0.19 $Y=-0.245 $X2=1.605
+ $Y2=2.895
cc_79 VNB N_A_425_117#_c_1049_n 0.00233015f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.845
cc_80 VNB N_A_425_117#_c_1050_n 0.00141548f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.08
cc_81 VNB N_A_425_117#_c_1051_n 0.0021309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_425_117#_c_1052_n 0.0105277f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.9
cc_83 VNB N_A_425_117#_c_1053_n 0.00980236f $X=-0.19 $Y=-0.245 $X2=4.405
+ $Y2=1.05
cc_84 VNB X 0.0284043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_X_c_1159_n 0.0303016f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.895
cc_86 VNB X 0.0124797f $X=-0.19 $Y=-0.245 $X2=4.055 $Y2=2.07
cc_87 VNB N_VGND_c_1175_n 0.00987845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1176_n 0.0212331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1177_n 0.0224107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1178_n 0.0235996f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.93
cc_91 VNB N_VGND_c_1179_n 0.110207f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.08
cc_92 VNB N_VGND_c_1180_n 0.0047828f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.08
cc_93 VNB N_VGND_c_1181_n 0.0673221f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=2.98
cc_94 VNB N_VGND_c_1182_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=2.98
cc_95 VNB N_VGND_c_1183_n 0.0216969f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.69
cc_96 VNB N_VGND_c_1184_n 0.50541f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.525
cc_97 VPB N_A_86_305#_M1000_g 0.0284483f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.555
cc_98 VPB N_A_86_305#_c_182_n 0.0236107f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=1.93
cc_99 VPB N_A_86_305#_c_183_n 0.0103524f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=2.18
cc_100 VPB N_A_86_305#_c_184_n 0.0022727f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=2.895
cc_101 VPB N_A_86_305#_c_176_n 0.008255f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.08
cc_102 VPB N_A_86_305#_c_186_n 0.0452957f $X=-0.19 $Y=1.655 $X2=3.89 $Y2=2.98
cc_103 VPB N_A_86_305#_c_187_n 0.00553944f $X=-0.19 $Y=1.655 $X2=3.975 $Y2=2.895
cc_104 VPB N_A_86_305#_c_177_n 0.00607119f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.69
cc_105 VPB N_A_86_305#_c_178_n 0.0210739f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.69
cc_106 VPB N_A_86_305#_c_190_n 0.0299099f $X=-0.19 $Y=1.655 $X2=4.055 $Y2=2.07
cc_107 VPB N_A_86_305#_c_179_n 0.00766464f $X=-0.19 $Y=1.655 $X2=4.23 $Y2=1.905
cc_108 VPB N_A_M1016_g 0.0376181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB A 0.00312254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_c_280_n 0.0107292f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.555
cc_111 VPB N_A_474_313#_M1003_g 0.0356828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_474_313#_c_318_n 0.0183897f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.555
cc_113 VPB N_A_474_313#_c_319_n 0.00693896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_474_313#_M1019_g 0.020111f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=0.905
cc_115 VPB N_A_474_313#_c_320_n 0.0149355f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=1.93
cc_116 VPB N_A_474_313#_c_322_n 0.00228891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_474_313#_c_324_n 0.0167336f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.69
cc_118 VPB N_A_474_313#_c_326_n 0.0140572f $X=-0.19 $Y=1.655 $X2=4.055 $Y2=2.07
cc_119 VPB N_B_M1002_g 0.0224756f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=2.055
cc_120 VPB N_B_c_433_n 0.0515365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_B_c_434_n 0.0107898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_B_M1013_g 0.0358211f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.555
cc_123 VPB N_B_c_436_n 0.12777f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.525
cc_124 VPB N_B_c_424_n 0.0837262f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.08
cc_125 VPB N_B_M1006_g 0.0248475f $X=-0.19 $Y=1.655 $X2=4.485 $Y2=1.905
cc_126 VPB N_B_c_439_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.69
cc_127 VPB N_A_1263_295#_M1017_g 0.0202909f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.855
cc_128 VPB N_A_1263_295#_c_540_n 0.0197844f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.555
cc_129 VPB N_A_1263_295#_c_541_n 0.0078063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_1263_295#_c_542_n 0.00668214f $X=-0.19 $Y=1.655 $X2=0.655
+ $Y2=0.905
cc_131 VPB N_A_1263_295#_c_550_n 0.0341458f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=1.93
cc_132 VPB N_A_1263_295#_c_551_n 0.0106576f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=2.18
cc_133 VPB N_A_1263_295#_c_552_n 0.00694847f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=2.2
cc_134 VPB N_A_1263_295#_c_544_n 0.00230665f $X=-0.19 $Y=1.655 $X2=3.975
+ $Y2=2.895
cc_135 VPB N_C_M1011_g 0.0271558f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_C_c_614_n 0.012742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_C_M1008_g 0.0332899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB C 0.00235782f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=1.93
cc_139 VPB N_A_1363_127#_M1009_g 0.0269448f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.855
cc_140 VPB N_A_1363_127#_c_682_n 0.00444392f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=1.93
cc_141 VPB N_A_1363_127#_c_688_n 0.0046903f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.08
cc_142 VPB N_A_1363_127#_c_689_n 0.00294588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_1363_127#_c_690_n 0.00144208f $X=-0.19 $Y=1.655 $X2=3.975
+ $Y2=2.745
cc_144 VPB N_A_1363_127#_c_684_n 0.00197824f $X=-0.19 $Y=1.655 $X2=0.615
+ $Y2=1.69
cc_145 VPB N_A_42_411#_c_768_n 0.038533f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.525
cc_146 VPB N_A_42_411#_c_769_n 0.00188597f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.845
cc_147 VPB N_A_42_411#_c_770_n 0.014724f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=1.93
cc_148 VPB N_A_42_411#_c_765_n 0.0179523f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=1.93
cc_149 VPB N_VPWR_c_842_n 0.00401817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_843_n 0.0278723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_844_n 0.0119718f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=1.93
cc_152 VPB N_VPWR_c_845_n 0.0714992f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.845
cc_153 VPB N_VPWR_c_846_n 0.00324402f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.08
cc_154 VPB N_VPWR_c_847_n 0.0178789f $X=-0.19 $Y=1.655 $X2=3.89 $Y2=2.98
cc_155 VPB N_VPWR_c_848_n 0.107448f $X=-0.19 $Y=1.655 $X2=4.485 $Y2=1.905
cc_156 VPB N_VPWR_c_849_n 0.0310362f $X=-0.19 $Y=1.655 $X2=4.405 $Y2=1.05
cc_157 VPB N_VPWR_c_841_n 0.119258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_851_n 0.00541171f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.525
cc_159 VPB N_VPWR_c_852_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_402_411#_c_923_n 0.00415815f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.555
cc_161 VPB N_A_402_411#_c_924_n 0.00328617f $X=-0.19 $Y=1.655 $X2=0.655
+ $Y2=1.525
cc_162 VPB N_A_402_411#_c_925_n 3.29996e-19 $X=-0.19 $Y=1.655 $X2=0.655
+ $Y2=0.905
cc_163 VPB N_A_402_411#_c_915_n 0.00562658f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=1.93
cc_164 VPB N_A_402_411#_c_927_n 0.00971891f $X=-0.19 $Y=1.655 $X2=4.485
+ $Y2=1.215
cc_165 VPB N_A_402_411#_c_922_n 0.00507537f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=1.93
cc_166 VPB N_A_402_411#_c_929_n 0.00803929f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=2.98
cc_167 VPB N_A_425_117#_c_1054_n 0.0258977f $X=-0.19 $Y=1.655 $X2=4.485
+ $Y2=1.215
cc_168 VPB N_A_425_117#_c_1055_n 0.0014735f $X=-0.19 $Y=1.655 $X2=4.485
+ $Y2=1.905
cc_169 VPB N_A_425_117#_c_1056_n 0.00320143f $X=-0.19 $Y=1.655 $X2=0.595
+ $Y2=1.69
cc_170 VPB N_A_425_117#_c_1057_n 0.00378903f $X=-0.19 $Y=1.655 $X2=1.605
+ $Y2=2.98
cc_171 VPB N_A_425_117#_c_1052_n 0.0189356f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=2.9
cc_172 VPB N_A_425_117#_c_1053_n 0.00151819f $X=-0.19 $Y=1.655 $X2=4.405
+ $Y2=1.05
cc_173 VPB X 0.0574174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 N_A_86_305#_M1007_g N_A_c_278_n 0.0184123f $X=0.655 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_86_305#_c_176_n N_A_c_278_n 0.00112447f $X=1.565 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A_86_305#_M1000_g N_A_M1016_g 0.0125283f $X=0.57 $Y=2.555 $X2=0 $Y2=0
cc_177 N_A_86_305#_c_182_n N_A_M1016_g 0.0162909f $X=1.44 $Y=1.93 $X2=0 $Y2=0
cc_178 N_A_86_305#_c_183_n N_A_M1016_g 0.0117019f $X=1.605 $Y=2.18 $X2=0 $Y2=0
cc_179 N_A_86_305#_c_184_n N_A_M1016_g 0.00350963f $X=1.605 $Y=2.895 $X2=0 $Y2=0
cc_180 N_A_86_305#_c_198_p N_A_M1016_g 0.0136078f $X=1.605 $Y=2.2 $X2=0 $Y2=0
cc_181 N_A_86_305#_c_177_n N_A_M1016_g 0.0031265f $X=0.595 $Y=1.69 $X2=0 $Y2=0
cc_182 N_A_86_305#_c_178_n N_A_M1016_g 0.00306348f $X=0.595 $Y=1.69 $X2=0 $Y2=0
cc_183 N_A_86_305#_M1007_g A 0.00400595f $X=0.655 $Y=0.905 $X2=0 $Y2=0
cc_184 N_A_86_305#_c_182_n A 0.0244356f $X=1.44 $Y=1.93 $X2=0 $Y2=0
cc_185 N_A_86_305#_c_176_n A 0.03321f $X=1.565 $Y=1.08 $X2=0 $Y2=0
cc_186 N_A_86_305#_c_177_n A 0.0107135f $X=0.595 $Y=1.69 $X2=0 $Y2=0
cc_187 N_A_86_305#_M1007_g N_A_c_280_n 0.010989f $X=0.655 $Y=0.905 $X2=0 $Y2=0
cc_188 N_A_86_305#_c_182_n N_A_c_280_n 0.00293841f $X=1.44 $Y=1.93 $X2=0 $Y2=0
cc_189 N_A_86_305#_c_176_n N_A_c_280_n 0.0166603f $X=1.565 $Y=1.08 $X2=0 $Y2=0
cc_190 N_A_86_305#_c_177_n N_A_c_280_n 8.38617e-19 $X=0.595 $Y=1.69 $X2=0 $Y2=0
cc_191 N_A_86_305#_c_178_n N_A_c_280_n 0.00903084f $X=0.595 $Y=1.69 $X2=0 $Y2=0
cc_192 N_A_86_305#_c_186_n N_A_474_313#_M1003_g 0.00118849f $X=3.89 $Y=2.98
+ $X2=0 $Y2=0
cc_193 N_A_86_305#_c_186_n N_A_474_313#_M1019_g 0.0011735f $X=3.89 $Y=2.98 $X2=0
+ $Y2=0
cc_194 N_A_86_305#_c_190_n N_A_474_313#_M1019_g 0.00597821f $X=4.055 $Y=2.07
+ $X2=0 $Y2=0
cc_195 N_A_86_305#_c_179_n N_A_474_313#_M1021_g 4.91414e-19 $X=4.23 $Y=1.905
+ $X2=0 $Y2=0
cc_196 N_A_86_305#_c_180_n N_A_474_313#_M1021_g 0.00101885f $X=4.405 $Y=1.05
+ $X2=0 $Y2=0
cc_197 N_A_86_305#_M1021_d N_A_474_313#_c_323_n 0.00907757f $X=4.03 $Y=0.625
+ $X2=0 $Y2=0
cc_198 N_A_86_305#_c_180_n N_A_474_313#_c_323_n 0.0246856f $X=4.405 $Y=1.05
+ $X2=0 $Y2=0
cc_199 N_A_86_305#_c_180_n N_A_474_313#_c_324_n 0.106461f $X=4.405 $Y=1.05 $X2=0
+ $Y2=0
cc_200 N_A_86_305#_c_190_n N_A_474_313#_c_325_n 0.0201558f $X=4.055 $Y=2.07
+ $X2=0 $Y2=0
cc_201 N_A_86_305#_c_179_n N_A_474_313#_c_325_n 0.0188763f $X=4.23 $Y=1.905
+ $X2=0 $Y2=0
cc_202 N_A_86_305#_c_190_n N_A_474_313#_c_326_n 0.00835065f $X=4.055 $Y=2.07
+ $X2=0 $Y2=0
cc_203 N_A_86_305#_c_179_n N_A_474_313#_c_326_n 0.00334234f $X=4.23 $Y=1.905
+ $X2=0 $Y2=0
cc_204 N_A_86_305#_c_179_n N_A_474_313#_c_327_n 0.00601149f $X=4.23 $Y=1.905
+ $X2=0 $Y2=0
cc_205 N_A_86_305#_c_183_n N_B_M1002_g 0.00431593f $X=1.605 $Y=2.18 $X2=0 $Y2=0
cc_206 N_A_86_305#_c_198_p N_B_M1002_g 0.00970092f $X=1.605 $Y=2.2 $X2=0 $Y2=0
cc_207 N_A_86_305#_c_186_n N_B_M1002_g 0.0161752f $X=3.89 $Y=2.98 $X2=0 $Y2=0
cc_208 N_A_86_305#_c_176_n N_B_M1018_g 0.00120528f $X=1.565 $Y=1.08 $X2=0 $Y2=0
cc_209 N_A_86_305#_c_186_n N_B_c_433_n 0.0119918f $X=3.89 $Y=2.98 $X2=0 $Y2=0
cc_210 N_A_86_305#_c_186_n N_B_M1013_g 0.013908f $X=3.89 $Y=2.98 $X2=0 $Y2=0
cc_211 N_A_86_305#_c_186_n N_B_c_436_n 0.0218373f $X=3.89 $Y=2.98 $X2=0 $Y2=0
cc_212 N_A_86_305#_c_190_n N_B_c_436_n 0.00969667f $X=4.055 $Y=2.07 $X2=0 $Y2=0
cc_213 N_A_86_305#_c_180_n N_B_c_423_n 0.0111431f $X=4.405 $Y=1.05 $X2=0 $Y2=0
cc_214 N_A_86_305#_c_186_n N_B_c_424_n 0.00217908f $X=3.89 $Y=2.98 $X2=0 $Y2=0
cc_215 N_A_86_305#_c_187_n N_B_c_424_n 0.00338011f $X=3.975 $Y=2.895 $X2=0 $Y2=0
cc_216 N_A_86_305#_c_190_n N_B_c_424_n 0.0111431f $X=4.055 $Y=2.07 $X2=0 $Y2=0
cc_217 N_A_86_305#_c_179_n N_B_c_428_n 0.0111431f $X=4.23 $Y=1.905 $X2=0 $Y2=0
cc_218 N_A_86_305#_M1004_d N_A_42_411#_c_758_n 0.0102533f $X=1.425 $Y=0.585
+ $X2=0 $Y2=0
cc_219 N_A_86_305#_M1007_g N_A_42_411#_c_758_n 0.0130075f $X=0.655 $Y=0.905
+ $X2=0 $Y2=0
cc_220 N_A_86_305#_c_176_n N_A_42_411#_c_758_n 0.0130182f $X=1.565 $Y=1.08 $X2=0
+ $Y2=0
cc_221 N_A_86_305#_M1004_d N_A_42_411#_c_759_n 0.00543658f $X=1.425 $Y=0.585
+ $X2=0 $Y2=0
cc_222 N_A_86_305#_c_176_n N_A_42_411#_c_759_n 0.0360076f $X=1.565 $Y=1.08 $X2=0
+ $Y2=0
cc_223 N_A_86_305#_c_176_n N_A_42_411#_c_761_n 0.0137872f $X=1.565 $Y=1.08 $X2=0
+ $Y2=0
cc_224 N_A_86_305#_M1007_g N_A_42_411#_c_764_n 0.0139396f $X=0.655 $Y=0.905
+ $X2=0 $Y2=0
cc_225 N_A_86_305#_c_177_n N_A_42_411#_c_764_n 0.00945551f $X=0.595 $Y=1.69
+ $X2=0 $Y2=0
cc_226 N_A_86_305#_c_178_n N_A_42_411#_c_764_n 0.00142205f $X=0.595 $Y=1.69
+ $X2=0 $Y2=0
cc_227 N_A_86_305#_M1000_g N_A_42_411#_c_770_n 0.00104673f $X=0.57 $Y=2.555
+ $X2=0 $Y2=0
cc_228 N_A_86_305#_c_178_n N_A_42_411#_c_770_n 3.95676e-19 $X=0.595 $Y=1.69
+ $X2=0 $Y2=0
cc_229 N_A_86_305#_M1000_g N_A_42_411#_c_765_n 0.00252518f $X=0.57 $Y=2.555
+ $X2=0 $Y2=0
cc_230 N_A_86_305#_M1007_g N_A_42_411#_c_765_n 0.00669591f $X=0.655 $Y=0.905
+ $X2=0 $Y2=0
cc_231 N_A_86_305#_c_177_n N_A_42_411#_c_765_n 0.0298935f $X=0.595 $Y=1.69 $X2=0
+ $Y2=0
cc_232 N_A_86_305#_c_178_n N_A_42_411#_c_765_n 0.00743403f $X=0.595 $Y=1.69
+ $X2=0 $Y2=0
cc_233 N_A_86_305#_M1000_g N_VPWR_c_842_n 0.0181462f $X=0.57 $Y=2.555 $X2=0
+ $Y2=0
cc_234 N_A_86_305#_c_182_n N_VPWR_c_842_n 0.0125739f $X=1.44 $Y=1.93 $X2=0 $Y2=0
cc_235 N_A_86_305#_c_184_n N_VPWR_c_842_n 0.00614895f $X=1.605 $Y=2.895 $X2=0
+ $Y2=0
cc_236 N_A_86_305#_c_198_p N_VPWR_c_842_n 0.023891f $X=1.605 $Y=2.2 $X2=0 $Y2=0
cc_237 N_A_86_305#_c_177_n N_VPWR_c_842_n 0.0118601f $X=0.595 $Y=1.69 $X2=0
+ $Y2=0
cc_238 N_A_86_305#_c_178_n N_VPWR_c_842_n 4.86372e-19 $X=0.595 $Y=1.69 $X2=0
+ $Y2=0
cc_239 N_A_86_305#_M1000_g N_VPWR_c_847_n 0.00452967f $X=0.57 $Y=2.555 $X2=0
+ $Y2=0
cc_240 N_A_86_305#_c_184_n N_VPWR_c_848_n 0.0221635f $X=1.605 $Y=2.895 $X2=0
+ $Y2=0
cc_241 N_A_86_305#_c_186_n N_VPWR_c_848_n 0.138471f $X=3.89 $Y=2.98 $X2=0 $Y2=0
cc_242 N_A_86_305#_c_190_n N_VPWR_c_848_n 0.0114579f $X=4.055 $Y=2.07 $X2=0
+ $Y2=0
cc_243 N_A_86_305#_M1000_g N_VPWR_c_841_n 0.0089278f $X=0.57 $Y=2.555 $X2=0
+ $Y2=0
cc_244 N_A_86_305#_c_184_n N_VPWR_c_841_n 0.0126536f $X=1.605 $Y=2.895 $X2=0
+ $Y2=0
cc_245 N_A_86_305#_c_186_n N_VPWR_c_841_n 0.0766555f $X=3.89 $Y=2.98 $X2=0 $Y2=0
cc_246 N_A_86_305#_c_190_n N_VPWR_c_841_n 0.0140075f $X=4.055 $Y=2.07 $X2=0
+ $Y2=0
cc_247 N_A_86_305#_c_183_n N_A_402_411#_c_923_n 0.00946607f $X=1.605 $Y=2.18
+ $X2=0 $Y2=0
cc_248 N_A_86_305#_c_198_p N_A_402_411#_c_923_n 0.0235884f $X=1.605 $Y=2.2 $X2=0
+ $Y2=0
cc_249 N_A_86_305#_M1019_d N_A_402_411#_c_924_n 0.00369473f $X=3.495 $Y=1.885
+ $X2=0 $Y2=0
cc_250 N_A_86_305#_c_186_n N_A_402_411#_c_924_n 0.0895938f $X=3.89 $Y=2.98 $X2=0
+ $Y2=0
cc_251 N_A_86_305#_c_190_n N_A_402_411#_c_924_n 0.014618f $X=4.055 $Y=2.07 $X2=0
+ $Y2=0
cc_252 N_A_86_305#_c_198_p N_A_402_411#_c_925_n 0.0116786f $X=1.605 $Y=2.2 $X2=0
+ $Y2=0
cc_253 N_A_86_305#_c_186_n N_A_402_411#_c_925_n 0.022162f $X=3.89 $Y=2.98 $X2=0
+ $Y2=0
cc_254 N_A_86_305#_M1019_d N_A_402_411#_c_915_n 0.0110792f $X=3.495 $Y=1.885
+ $X2=0 $Y2=0
cc_255 N_A_86_305#_c_190_n N_A_402_411#_c_915_n 0.0479732f $X=4.055 $Y=2.07
+ $X2=0 $Y2=0
cc_256 N_A_86_305#_M1019_d N_A_425_117#_c_1054_n 0.0110348f $X=3.495 $Y=1.885
+ $X2=0 $Y2=0
cc_257 N_A_86_305#_c_190_n N_A_425_117#_c_1054_n 0.0722531f $X=4.055 $Y=2.07
+ $X2=0 $Y2=0
cc_258 N_A_86_305#_M1007_g N_VGND_c_1178_n 0.0033294f $X=0.655 $Y=0.905 $X2=0
+ $Y2=0
cc_259 N_A_86_305#_M1007_g N_VGND_c_1184_n 0.00480627f $X=0.655 $Y=0.905 $X2=0
+ $Y2=0
cc_260 N_A_M1016_g N_B_M1002_g 0.0189679f $X=1.39 $Y=2.555 $X2=0 $Y2=0
cc_261 N_A_c_278_n N_B_M1018_g 0.0124122f $X=1.35 $Y=1.335 $X2=0 $Y2=0
cc_262 N_A_c_280_n N_B_M1018_g 3.50962e-19 $X=1.39 $Y=1.5 $X2=0 $Y2=0
cc_263 N_A_c_278_n N_A_42_411#_c_758_n 0.016958f $X=1.35 $Y=1.335 $X2=0 $Y2=0
cc_264 A N_A_42_411#_c_758_n 0.0104016f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_265 N_A_c_280_n N_A_42_411#_c_758_n 0.00118591f $X=1.39 $Y=1.5 $X2=0 $Y2=0
cc_266 N_A_c_278_n N_A_42_411#_c_759_n 0.00363069f $X=1.35 $Y=1.335 $X2=0 $Y2=0
cc_267 N_A_c_278_n N_A_42_411#_c_764_n 0.00201091f $X=1.35 $Y=1.335 $X2=0 $Y2=0
cc_268 A N_A_42_411#_c_764_n 0.00293182f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_269 N_A_M1016_g N_VPWR_c_842_n 0.0100551f $X=1.39 $Y=2.555 $X2=0 $Y2=0
cc_270 N_A_M1016_g N_VPWR_c_848_n 0.00510245f $X=1.39 $Y=2.555 $X2=0 $Y2=0
cc_271 N_A_M1016_g N_VPWR_c_841_n 0.0103676f $X=1.39 $Y=2.555 $X2=0 $Y2=0
cc_272 A N_VGND_M1007_d 0.00488155f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_273 N_A_c_278_n N_VGND_c_1179_n 0.00332252f $X=1.35 $Y=1.335 $X2=0 $Y2=0
cc_274 N_A_c_278_n N_VGND_c_1184_n 0.00480627f $X=1.35 $Y=1.335 $X2=0 $Y2=0
cc_275 N_A_474_313#_M1003_g N_B_M1002_g 0.0163745f $X=2.445 $Y=2.375 $X2=0 $Y2=0
cc_276 N_A_474_313#_M1020_g N_B_M1018_g 0.00919073f $X=2.595 $Y=1.015 $X2=0
+ $Y2=0
cc_277 N_A_474_313#_M1003_g N_B_c_433_n 0.00737859f $X=2.445 $Y=2.375 $X2=0
+ $Y2=0
cc_278 N_A_474_313#_M1020_g N_B_c_419_n 0.00337775f $X=2.595 $Y=1.015 $X2=0
+ $Y2=0
cc_279 N_A_474_313#_M1003_g N_B_M1013_g 0.026059f $X=2.445 $Y=2.375 $X2=0 $Y2=0
cc_280 N_A_474_313#_c_318_n N_B_M1013_g 0.0106871f $X=3.345 $Y=1.64 $X2=0 $Y2=0
cc_281 N_A_474_313#_M1019_g N_B_M1013_g 0.0212578f $X=3.42 $Y=2.305 $X2=0 $Y2=0
cc_282 N_A_474_313#_M1019_g N_B_c_436_n 0.00882199f $X=3.42 $Y=2.305 $X2=0 $Y2=0
cc_283 N_A_474_313#_M1020_g N_B_M1010_g 0.0109606f $X=2.595 $Y=1.015 $X2=0 $Y2=0
cc_284 N_A_474_313#_c_318_n N_B_M1010_g 0.00995033f $X=3.345 $Y=1.64 $X2=0 $Y2=0
cc_285 N_A_474_313#_M1021_g N_B_M1010_g 0.0125072f $X=3.955 $Y=0.945 $X2=0 $Y2=0
cc_286 N_A_474_313#_M1021_g N_B_c_422_n 0.00737233f $X=3.955 $Y=0.945 $X2=0
+ $Y2=0
cc_287 N_A_474_313#_M1021_g N_B_c_423_n 0.0134764f $X=3.955 $Y=0.945 $X2=0 $Y2=0
cc_288 N_A_474_313#_c_323_n N_B_c_423_n 0.0163773f $X=4.83 $Y=0.7 $X2=0 $Y2=0
cc_289 N_A_474_313#_c_324_n N_B_c_423_n 0.00691194f $X=4.995 $Y=0.855 $X2=0
+ $Y2=0
cc_290 N_A_474_313#_c_327_n N_B_c_423_n 8.36943e-19 $X=4.025 $Y=1.395 $X2=0
+ $Y2=0
cc_291 N_A_474_313#_c_324_n N_B_c_424_n 0.0221731f $X=4.995 $Y=0.855 $X2=0 $Y2=0
cc_292 N_A_474_313#_c_326_n N_B_c_424_n 0.0071705f $X=4.025 $Y=1.56 $X2=0 $Y2=0
cc_293 N_A_474_313#_c_324_n N_B_c_425_n 0.00296946f $X=4.995 $Y=0.855 $X2=0
+ $Y2=0
cc_294 N_A_474_313#_c_324_n B 0.024413f $X=4.995 $Y=0.855 $X2=0 $Y2=0
cc_295 N_A_474_313#_c_324_n N_B_c_430_n 0.016039f $X=4.995 $Y=0.855 $X2=0 $Y2=0
cc_296 N_A_474_313#_c_324_n N_B_c_431_n 0.00998512f $X=4.995 $Y=0.855 $X2=0
+ $Y2=0
cc_297 N_A_474_313#_M1020_g N_A_42_411#_c_759_n 0.00154542f $X=2.595 $Y=1.015
+ $X2=0 $Y2=0
cc_298 N_A_474_313#_c_319_n N_A_42_411#_c_760_n 0.00860924f $X=2.67 $Y=1.64
+ $X2=0 $Y2=0
cc_299 N_A_474_313#_M1003_g N_A_42_411#_c_769_n 0.0207442f $X=2.445 $Y=2.375
+ $X2=0 $Y2=0
cc_300 N_A_474_313#_c_318_n N_A_42_411#_c_769_n 0.00751697f $X=3.345 $Y=1.64
+ $X2=0 $Y2=0
cc_301 N_A_474_313#_c_319_n N_A_42_411#_c_769_n 0.00826294f $X=2.67 $Y=1.64
+ $X2=0 $Y2=0
cc_302 N_A_474_313#_c_322_n N_A_42_411#_c_769_n 9.56406e-19 $X=3.42 $Y=1.655
+ $X2=0 $Y2=0
cc_303 N_A_474_313#_M1020_g N_A_42_411#_c_762_n 0.0106167f $X=2.595 $Y=1.015
+ $X2=0 $Y2=0
cc_304 N_A_474_313#_M1020_g N_A_42_411#_c_763_n 0.00614811f $X=2.595 $Y=1.015
+ $X2=0 $Y2=0
cc_305 N_A_474_313#_M1020_g N_A_42_411#_c_766_n 0.0147015f $X=2.595 $Y=1.015
+ $X2=0 $Y2=0
cc_306 N_A_474_313#_c_318_n N_A_42_411#_c_766_n 0.00480759f $X=3.345 $Y=1.64
+ $X2=0 $Y2=0
cc_307 N_A_474_313#_c_319_n N_A_42_411#_c_766_n 9.23032e-19 $X=2.67 $Y=1.64
+ $X2=0 $Y2=0
cc_308 N_A_474_313#_M1020_g N_A_42_411#_c_767_n 0.00474478f $X=2.595 $Y=1.015
+ $X2=0 $Y2=0
cc_309 N_A_474_313#_c_318_n N_A_42_411#_c_767_n 0.00633169f $X=3.345 $Y=1.64
+ $X2=0 $Y2=0
cc_310 N_A_474_313#_c_324_n N_VPWR_c_843_n 0.0496789f $X=4.995 $Y=0.855 $X2=0
+ $Y2=0
cc_311 N_A_474_313#_c_324_n N_VPWR_c_848_n 0.0167213f $X=4.995 $Y=0.855 $X2=0
+ $Y2=0
cc_312 N_A_474_313#_c_324_n N_VPWR_c_841_n 0.0095959f $X=4.995 $Y=0.855 $X2=0
+ $Y2=0
cc_313 N_A_474_313#_M1003_g N_A_402_411#_c_923_n 0.00273282f $X=2.445 $Y=2.375
+ $X2=0 $Y2=0
cc_314 N_A_474_313#_M1003_g N_A_402_411#_c_924_n 0.0137704f $X=2.445 $Y=2.375
+ $X2=0 $Y2=0
cc_315 N_A_474_313#_M1019_g N_A_402_411#_c_924_n 0.0123318f $X=3.42 $Y=2.305
+ $X2=0 $Y2=0
cc_316 N_A_474_313#_M1019_g N_A_402_411#_c_915_n 0.0157057f $X=3.42 $Y=2.305
+ $X2=0 $Y2=0
cc_317 N_A_474_313#_c_320_n N_A_402_411#_c_915_n 0.0166074f $X=3.86 $Y=1.655
+ $X2=0 $Y2=0
cc_318 N_A_474_313#_M1021_g N_A_402_411#_c_915_n 0.00934298f $X=3.955 $Y=0.945
+ $X2=0 $Y2=0
cc_319 N_A_474_313#_c_393_p N_A_402_411#_c_915_n 0.0127796f $X=4.06 $Y=0.7 $X2=0
+ $Y2=0
cc_320 N_A_474_313#_c_326_n N_A_402_411#_c_915_n 0.00392295f $X=4.025 $Y=1.56
+ $X2=0 $Y2=0
cc_321 N_A_474_313#_c_327_n N_A_402_411#_c_915_n 0.0638805f $X=4.025 $Y=1.395
+ $X2=0 $Y2=0
cc_322 N_A_474_313#_M1005_s N_A_402_411#_c_916_n 0.00467114f $X=4.85 $Y=0.235
+ $X2=0 $Y2=0
cc_323 N_A_474_313#_M1021_g N_A_402_411#_c_916_n 0.00137802f $X=3.955 $Y=0.945
+ $X2=0 $Y2=0
cc_324 N_A_474_313#_c_323_n N_A_402_411#_c_916_n 0.0691523f $X=4.83 $Y=0.7 $X2=0
+ $Y2=0
cc_325 N_A_474_313#_c_393_p N_A_402_411#_c_916_n 0.0122794f $X=4.06 $Y=0.7 $X2=0
+ $Y2=0
cc_326 N_A_474_313#_M1020_g N_A_425_117#_c_1044_n 0.00508076f $X=2.595 $Y=1.015
+ $X2=0 $Y2=0
cc_327 N_A_474_313#_c_319_n N_A_425_117#_c_1044_n 3.301e-19 $X=2.67 $Y=1.64
+ $X2=0 $Y2=0
cc_328 N_A_474_313#_M1020_g N_A_425_117#_c_1045_n 0.00304062f $X=2.595 $Y=1.015
+ $X2=0 $Y2=0
cc_329 N_A_474_313#_M1006_s N_A_425_117#_c_1054_n 0.0040317f $X=4.85 $Y=1.785
+ $X2=0 $Y2=0
cc_330 N_A_474_313#_M1019_g N_A_425_117#_c_1054_n 0.00875945f $X=3.42 $Y=2.305
+ $X2=0 $Y2=0
cc_331 N_A_474_313#_c_320_n N_A_425_117#_c_1054_n 0.00489943f $X=3.86 $Y=1.655
+ $X2=0 $Y2=0
cc_332 N_A_474_313#_c_324_n N_A_425_117#_c_1054_n 0.0296322f $X=4.995 $Y=0.855
+ $X2=0 $Y2=0
cc_333 N_A_474_313#_c_325_n N_A_425_117#_c_1054_n 0.00181318f $X=4.025 $Y=1.56
+ $X2=0 $Y2=0
cc_334 N_A_474_313#_c_318_n N_A_425_117#_c_1055_n 7.06517e-19 $X=3.345 $Y=1.64
+ $X2=0 $Y2=0
cc_335 N_A_474_313#_M1003_g N_A_425_117#_c_1056_n 2.79858e-19 $X=2.445 $Y=2.375
+ $X2=0 $Y2=0
cc_336 N_A_474_313#_c_318_n N_A_425_117#_c_1056_n 0.00736635f $X=3.345 $Y=1.64
+ $X2=0 $Y2=0
cc_337 N_A_474_313#_M1019_g N_A_425_117#_c_1056_n 0.00666869f $X=3.42 $Y=2.305
+ $X2=0 $Y2=0
cc_338 N_A_474_313#_M1003_g N_A_425_117#_c_1053_n 5.34602e-19 $X=2.445 $Y=2.375
+ $X2=0 $Y2=0
cc_339 N_A_474_313#_M1020_g N_A_425_117#_c_1053_n 0.00167137f $X=2.595 $Y=1.015
+ $X2=0 $Y2=0
cc_340 N_A_474_313#_c_318_n N_A_425_117#_c_1053_n 0.00861527f $X=3.345 $Y=1.64
+ $X2=0 $Y2=0
cc_341 N_A_474_313#_M1019_g N_A_425_117#_c_1053_n 0.00327618f $X=3.42 $Y=2.305
+ $X2=0 $Y2=0
cc_342 N_A_474_313#_c_322_n N_A_425_117#_c_1053_n 0.0034267f $X=3.42 $Y=1.655
+ $X2=0 $Y2=0
cc_343 N_A_474_313#_M1005_s N_VGND_c_1184_n 0.00229492f $X=4.85 $Y=0.235 $X2=0
+ $Y2=0
cc_344 N_B_M1018_g N_A_42_411#_c_758_n 0.00551637f $X=2.05 $Y=0.905 $X2=0 $Y2=0
cc_345 N_B_M1018_g N_A_42_411#_c_759_n 0.0154529f $X=2.05 $Y=0.905 $X2=0 $Y2=0
cc_346 N_B_M1018_g N_A_42_411#_c_760_n 0.0056021f $X=2.05 $Y=0.905 $X2=0 $Y2=0
cc_347 N_B_M1002_g N_A_42_411#_c_761_n 0.00515433f $X=1.935 $Y=2.475 $X2=0 $Y2=0
cc_348 N_B_M1002_g N_A_42_411#_c_769_n 6.06703e-19 $X=1.935 $Y=2.475 $X2=0 $Y2=0
cc_349 N_B_M1013_g N_A_42_411#_c_769_n 0.00662908f $X=2.875 $Y=2.375 $X2=0 $Y2=0
cc_350 N_B_M1018_g N_A_42_411#_c_762_n 4.90214e-19 $X=2.05 $Y=0.905 $X2=0 $Y2=0
cc_351 N_B_M1010_g N_A_42_411#_c_762_n 0.00270368f $X=3.295 $Y=0.905 $X2=0 $Y2=0
cc_352 N_B_M1010_g N_A_42_411#_c_763_n 4.06541e-19 $X=3.295 $Y=0.905 $X2=0 $Y2=0
cc_353 N_B_c_436_n N_VPWR_c_843_n 0.0018415f $X=4.625 $Y=3.14 $X2=0 $Y2=0
cc_354 N_B_M1006_g N_VPWR_c_843_n 0.0231912f $X=5.21 $Y=2.415 $X2=0 $Y2=0
cc_355 B N_VPWR_c_843_n 0.0189806f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_356 N_B_c_431_n N_VPWR_c_843_n 0.00677923f $X=5.425 $Y=1.35 $X2=0 $Y2=0
cc_357 N_B_c_434_n N_VPWR_c_848_n 0.0658023f $X=2.01 $Y=3.14 $X2=0 $Y2=0
cc_358 N_B_M1006_g N_VPWR_c_848_n 0.00445056f $X=5.21 $Y=2.415 $X2=0 $Y2=0
cc_359 N_B_c_433_n N_VPWR_c_841_n 0.0186948f $X=2.8 $Y=3.14 $X2=0 $Y2=0
cc_360 N_B_c_434_n N_VPWR_c_841_n 0.00506369f $X=2.01 $Y=3.14 $X2=0 $Y2=0
cc_361 N_B_c_436_n N_VPWR_c_841_n 0.0534722f $X=4.625 $Y=3.14 $X2=0 $Y2=0
cc_362 N_B_M1006_g N_VPWR_c_841_n 0.0082324f $X=5.21 $Y=2.415 $X2=0 $Y2=0
cc_363 N_B_c_439_n N_VPWR_c_841_n 0.00372267f $X=2.875 $Y=3.14 $X2=0 $Y2=0
cc_364 N_B_M1002_g N_A_402_411#_c_923_n 0.00633579f $X=1.935 $Y=2.475 $X2=0
+ $Y2=0
cc_365 N_B_M1013_g N_A_402_411#_c_924_n 0.0146702f $X=2.875 $Y=2.375 $X2=0 $Y2=0
cc_366 N_B_M1002_g N_A_402_411#_c_925_n 0.00227642f $X=1.935 $Y=2.475 $X2=0
+ $Y2=0
cc_367 N_B_M1010_g N_A_402_411#_c_915_n 0.00794051f $X=3.295 $Y=0.905 $X2=0
+ $Y2=0
cc_368 N_B_c_422_n N_A_402_411#_c_916_n 0.0168502f $X=4.625 $Y=0.18 $X2=0 $Y2=0
cc_369 N_B_c_423_n N_A_402_411#_c_916_n 0.0104077f $X=4.7 $Y=1.185 $X2=0 $Y2=0
cc_370 N_B_c_425_n N_A_402_411#_c_916_n 0.0145796f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_371 N_B_M1010_g N_A_402_411#_c_917_n 0.003419f $X=3.295 $Y=0.905 $X2=0 $Y2=0
cc_372 N_B_c_422_n N_A_402_411#_c_917_n 0.00418768f $X=4.625 $Y=0.18 $X2=0 $Y2=0
cc_373 N_B_c_423_n N_A_402_411#_c_961_n 9.66558e-19 $X=4.7 $Y=1.185 $X2=0 $Y2=0
cc_374 N_B_c_425_n N_A_402_411#_c_961_n 0.0107602f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_375 B N_A_402_411#_c_918_n 0.0126577f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_376 N_B_c_431_n N_A_402_411#_c_918_n 0.00103994f $X=5.425 $Y=1.35 $X2=0 $Y2=0
cc_377 N_B_c_425_n N_A_402_411#_c_965_n 0.00632104f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_378 B N_A_402_411#_c_965_n 0.00948731f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_379 N_B_c_431_n N_A_402_411#_c_965_n 8.8406e-19 $X=5.425 $Y=1.35 $X2=0 $Y2=0
cc_380 N_B_M1018_g N_A_425_117#_c_1044_n 0.00587897f $X=2.05 $Y=0.905 $X2=0
+ $Y2=0
cc_381 N_B_c_419_n N_A_425_117#_c_1045_n 0.0143038f $X=3.22 $Y=0.18 $X2=0 $Y2=0
cc_382 N_B_M1010_g N_A_425_117#_c_1045_n 0.0084969f $X=3.295 $Y=0.905 $X2=0
+ $Y2=0
cc_383 N_B_M1018_g N_A_425_117#_c_1046_n 0.00792239f $X=2.05 $Y=0.905 $X2=0
+ $Y2=0
cc_384 N_B_c_419_n N_A_425_117#_c_1046_n 0.00529618f $X=3.22 $Y=0.18 $X2=0 $Y2=0
cc_385 N_B_c_425_n N_A_425_117#_c_1048_n 0.00147308f $X=5.21 $Y=1.185 $X2=0
+ $Y2=0
cc_386 B N_A_425_117#_c_1048_n 0.00779154f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_387 N_B_c_431_n N_A_425_117#_c_1048_n 7.45699e-19 $X=5.425 $Y=1.35 $X2=0
+ $Y2=0
cc_388 N_B_c_424_n N_A_425_117#_c_1054_n 0.0160371f $X=4.7 $Y=3.065 $X2=0 $Y2=0
cc_389 N_B_M1006_g N_A_425_117#_c_1054_n 0.010272f $X=5.21 $Y=2.415 $X2=0 $Y2=0
cc_390 B N_A_425_117#_c_1054_n 0.00328834f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_391 N_B_M1013_g N_A_425_117#_c_1055_n 0.0046644f $X=2.875 $Y=2.375 $X2=0
+ $Y2=0
cc_392 N_B_M1013_g N_A_425_117#_c_1056_n 0.00297146f $X=2.875 $Y=2.375 $X2=0
+ $Y2=0
cc_393 N_B_M1006_g N_A_425_117#_c_1052_n 0.00789799f $X=5.21 $Y=2.415 $X2=0
+ $Y2=0
cc_394 B N_A_425_117#_c_1052_n 0.0137989f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_395 N_B_c_431_n N_A_425_117#_c_1052_n 0.00132729f $X=5.425 $Y=1.35 $X2=0
+ $Y2=0
cc_396 N_B_M1010_g N_A_425_117#_c_1053_n 0.0274531f $X=3.295 $Y=0.905 $X2=0
+ $Y2=0
cc_397 N_B_c_425_n N_VGND_c_1175_n 0.00527444f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_398 N_B_c_420_n N_VGND_c_1179_n 0.0651842f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_399 N_B_c_425_n N_VGND_c_1179_n 0.0035993f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_400 N_B_c_419_n N_VGND_c_1184_n 0.0277331f $X=3.22 $Y=0.18 $X2=0 $Y2=0
cc_401 N_B_c_420_n N_VGND_c_1184_n 0.0107503f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_402 N_B_c_422_n N_VGND_c_1184_n 0.0400359f $X=4.625 $Y=0.18 $X2=0 $Y2=0
cc_403 N_B_c_425_n N_VGND_c_1184_n 0.0070319f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_404 N_B_c_427_n N_VGND_c_1184_n 0.00408042f $X=3.295 $Y=0.18 $X2=0 $Y2=0
cc_405 N_A_1263_295#_M1001_g N_C_c_612_n 0.0266886f $X=6.74 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_406 N_A_1263_295#_M1017_g N_C_M1011_g 0.0139989f $X=6.775 $Y=2.385 $X2=0
+ $Y2=0
cc_407 N_A_1263_295#_c_550_n N_C_M1011_g 0.0103913f $X=7.895 $Y=2.98 $X2=0 $Y2=0
cc_408 N_A_1263_295#_c_557_p N_C_M1011_g 0.00446445f $X=7.98 $Y=2.41 $X2=0 $Y2=0
cc_409 N_A_1263_295#_c_544_n N_C_c_613_n 0.00541671f $X=8.065 $Y=2.245 $X2=0
+ $Y2=0
cc_410 N_A_1263_295#_c_541_n N_C_c_614_n 0.0171317f $X=6.757 $Y=1.64 $X2=0 $Y2=0
cc_411 N_A_1263_295#_c_552_n N_C_M1008_g 0.00956463f $X=8.065 $Y=2.895 $X2=0
+ $Y2=0
cc_412 N_A_1263_295#_c_557_p N_C_M1008_g 0.00297037f $X=7.98 $Y=2.41 $X2=0 $Y2=0
cc_413 N_A_1263_295#_c_544_n N_C_M1008_g 0.0231747f $X=8.065 $Y=2.245 $X2=0
+ $Y2=0
cc_414 N_A_1263_295#_c_543_n N_C_M1015_g 0.0049071f $X=8.15 $Y=0.895 $X2=0 $Y2=0
cc_415 N_A_1263_295#_c_544_n N_C_M1015_g 0.00899398f $X=8.065 $Y=2.245 $X2=0
+ $Y2=0
cc_416 N_A_1263_295#_c_545_n N_C_M1015_g 0.00319949f $X=8.19 $Y=1.125 $X2=0
+ $Y2=0
cc_417 N_A_1263_295#_c_544_n N_C_c_617_n 0.0059599f $X=8.065 $Y=2.245 $X2=0
+ $Y2=0
cc_418 N_A_1263_295#_M1017_g N_A_1363_127#_c_692_n 0.00754181f $X=6.775 $Y=2.385
+ $X2=0 $Y2=0
cc_419 N_A_1263_295#_c_550_n N_A_1363_127#_c_692_n 0.0196019f $X=7.895 $Y=2.98
+ $X2=0 $Y2=0
cc_420 N_A_1263_295#_M1001_g N_A_1363_127#_c_682_n 0.00443107f $X=6.74 $Y=0.955
+ $X2=0 $Y2=0
cc_421 N_A_1263_295#_c_541_n N_A_1363_127#_c_682_n 0.00418522f $X=6.757 $Y=1.64
+ $X2=0 $Y2=0
cc_422 N_A_1263_295#_c_542_n N_A_1363_127#_c_682_n 0.0275507f $X=6.48 $Y=1.64
+ $X2=0 $Y2=0
cc_423 N_A_1263_295#_c_544_n N_A_1363_127#_c_683_n 0.0110868f $X=8.065 $Y=2.245
+ $X2=0 $Y2=0
cc_424 N_A_1263_295#_M1008_s N_A_1363_127#_c_688_n 0.0066702f $X=7.835 $Y=1.915
+ $X2=0 $Y2=0
cc_425 N_A_1263_295#_c_557_p N_A_1363_127#_c_688_n 0.00909304f $X=7.98 $Y=2.41
+ $X2=0 $Y2=0
cc_426 N_A_1263_295#_c_544_n N_A_1363_127#_c_688_n 0.022502f $X=8.065 $Y=2.245
+ $X2=0 $Y2=0
cc_427 N_A_1263_295#_M1017_g N_A_1363_127#_c_689_n 0.0037811f $X=6.775 $Y=2.385
+ $X2=0 $Y2=0
cc_428 N_A_1263_295#_c_542_n N_A_1363_127#_c_689_n 0.00644596f $X=6.48 $Y=1.64
+ $X2=0 $Y2=0
cc_429 N_A_1263_295#_M1017_g N_A_1363_127#_c_690_n 0.00222248f $X=6.775 $Y=2.385
+ $X2=0 $Y2=0
cc_430 N_A_1263_295#_c_542_n N_A_1363_127#_c_690_n 0.028655f $X=6.48 $Y=1.64
+ $X2=0 $Y2=0
cc_431 N_A_1263_295#_c_544_n N_A_1363_127#_c_684_n 0.00538917f $X=8.065 $Y=2.245
+ $X2=0 $Y2=0
cc_432 N_A_1263_295#_c_544_n N_A_1363_127#_c_685_n 8.57467e-19 $X=8.065 $Y=2.245
+ $X2=0 $Y2=0
cc_433 N_A_1263_295#_c_550_n N_VPWR_c_844_n 0.0123439f $X=7.895 $Y=2.98 $X2=0
+ $Y2=0
cc_434 N_A_1263_295#_c_544_n N_VPWR_c_844_n 0.0674604f $X=8.065 $Y=2.245 $X2=0
+ $Y2=0
cc_435 N_A_1263_295#_M1017_g N_VPWR_c_845_n 6.76935e-19 $X=6.775 $Y=2.385 $X2=0
+ $Y2=0
cc_436 N_A_1263_295#_c_550_n N_VPWR_c_845_n 0.0986629f $X=7.895 $Y=2.98 $X2=0
+ $Y2=0
cc_437 N_A_1263_295#_c_551_n N_VPWR_c_845_n 0.0222501f $X=6.645 $Y=2.98 $X2=0
+ $Y2=0
cc_438 N_A_1263_295#_c_550_n N_VPWR_c_841_n 0.0598638f $X=7.895 $Y=2.98 $X2=0
+ $Y2=0
cc_439 N_A_1263_295#_c_551_n N_VPWR_c_841_n 0.0127687f $X=6.645 $Y=2.98 $X2=0
+ $Y2=0
cc_440 N_A_1263_295#_M1001_g N_A_402_411#_c_919_n 0.00513659f $X=6.74 $Y=0.955
+ $X2=0 $Y2=0
cc_441 N_A_1263_295#_M1001_g N_A_402_411#_c_920_n 0.0044673f $X=6.74 $Y=0.955
+ $X2=0 $Y2=0
cc_442 N_A_1263_295#_c_550_n N_A_402_411#_c_927_n 0.0281621f $X=7.895 $Y=2.98
+ $X2=0 $Y2=0
cc_443 N_A_1263_295#_c_557_p N_A_402_411#_c_927_n 0.0375574f $X=7.98 $Y=2.41
+ $X2=0 $Y2=0
cc_444 N_A_1263_295#_c_544_n N_A_402_411#_c_927_n 0.00464118f $X=8.065 $Y=2.245
+ $X2=0 $Y2=0
cc_445 N_A_1263_295#_c_543_n N_A_402_411#_c_922_n 0.0483509f $X=8.15 $Y=0.895
+ $X2=0 $Y2=0
cc_446 N_A_1263_295#_M1008_s N_A_402_411#_c_929_n 0.00220321f $X=7.835 $Y=1.915
+ $X2=0 $Y2=0
cc_447 N_A_1263_295#_c_545_n N_A_402_411#_c_929_n 0.0483509f $X=8.19 $Y=1.125
+ $X2=0 $Y2=0
cc_448 N_A_1263_295#_c_542_n N_A_425_117#_M1017_s 0.0233995f $X=6.48 $Y=1.64
+ $X2=0 $Y2=0
cc_449 N_A_1263_295#_M1001_g N_A_425_117#_c_1047_n 0.00709813f $X=6.74 $Y=0.955
+ $X2=0 $Y2=0
cc_450 N_A_1263_295#_c_540_n N_A_425_117#_c_1047_n 0.00328384f $X=6.665 $Y=1.64
+ $X2=0 $Y2=0
cc_451 N_A_1263_295#_c_542_n N_A_425_117#_c_1047_n 0.0261578f $X=6.48 $Y=1.64
+ $X2=0 $Y2=0
cc_452 N_A_1263_295#_M1001_g N_A_425_117#_c_1100_n 0.0106232f $X=6.74 $Y=0.955
+ $X2=0 $Y2=0
cc_453 N_A_1263_295#_M1001_g N_A_425_117#_c_1049_n 0.0104275f $X=6.74 $Y=0.955
+ $X2=0 $Y2=0
cc_454 N_A_1263_295#_M1001_g N_A_425_117#_c_1050_n 0.00353823f $X=6.74 $Y=0.955
+ $X2=0 $Y2=0
cc_455 N_A_1263_295#_M1001_g N_A_425_117#_c_1051_n 5.58056e-19 $X=6.74 $Y=0.955
+ $X2=0 $Y2=0
cc_456 N_A_1263_295#_c_542_n N_A_425_117#_c_1057_n 0.00736637f $X=6.48 $Y=1.64
+ $X2=0 $Y2=0
cc_457 N_A_1263_295#_M1001_g N_A_425_117#_c_1052_n 0.00440418f $X=6.74 $Y=0.955
+ $X2=0 $Y2=0
cc_458 N_A_1263_295#_c_540_n N_A_425_117#_c_1052_n 0.00819021f $X=6.665 $Y=1.64
+ $X2=0 $Y2=0
cc_459 N_A_1263_295#_c_542_n N_A_425_117#_c_1052_n 0.099006f $X=6.48 $Y=1.64
+ $X2=0 $Y2=0
cc_460 N_A_1263_295#_c_543_n N_VGND_c_1176_n 0.029247f $X=8.15 $Y=0.895 $X2=0
+ $Y2=0
cc_461 N_A_1263_295#_c_543_n N_VGND_c_1181_n 0.00462837f $X=8.15 $Y=0.895 $X2=0
+ $Y2=0
cc_462 N_A_1263_295#_c_543_n N_VGND_c_1184_n 0.00728996f $X=8.15 $Y=0.895 $X2=0
+ $Y2=0
cc_463 N_C_M1015_g N_A_1363_127#_M1012_g 0.0137889f $X=8.365 $Y=0.895 $X2=0
+ $Y2=0
cc_464 N_C_M1008_g N_A_1363_127#_M1009_g 0.00988586f $X=8.195 $Y=2.235 $X2=0
+ $Y2=0
cc_465 N_C_M1011_g N_A_1363_127#_c_692_n 0.00771614f $X=7.205 $Y=2.385 $X2=0
+ $Y2=0
cc_466 N_C_c_612_n N_A_1363_127#_c_682_n 0.00207946f $X=7.17 $Y=1.385 $X2=0
+ $Y2=0
cc_467 N_C_c_614_n N_A_1363_127#_c_682_n 0.00377113f $X=7.54 $Y=1.46 $X2=0 $Y2=0
cc_468 C N_A_1363_127#_c_682_n 0.0348672f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_469 N_C_M1008_g N_A_1363_127#_c_683_n 3.64968e-19 $X=8.195 $Y=2.235 $X2=0
+ $Y2=0
cc_470 N_C_M1015_g N_A_1363_127#_c_683_n 9.99223e-19 $X=8.365 $Y=0.895 $X2=0
+ $Y2=0
cc_471 N_C_M1011_g N_A_1363_127#_c_688_n 0.00845664f $X=7.205 $Y=2.385 $X2=0
+ $Y2=0
cc_472 N_C_c_613_n N_A_1363_127#_c_688_n 0.00330085f $X=8.12 $Y=1.46 $X2=0 $Y2=0
cc_473 N_C_M1008_g N_A_1363_127#_c_688_n 0.00462837f $X=8.195 $Y=2.235 $X2=0
+ $Y2=0
cc_474 N_C_c_617_n N_A_1363_127#_c_688_n 0.00406504f $X=8.365 $Y=1.46 $X2=0
+ $Y2=0
cc_475 C N_A_1363_127#_c_688_n 0.00600197f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_476 N_C_M1011_g N_A_1363_127#_c_690_n 0.00309901f $X=7.205 $Y=2.385 $X2=0
+ $Y2=0
cc_477 N_C_c_614_n N_A_1363_127#_c_690_n 0.00126757f $X=7.54 $Y=1.46 $X2=0 $Y2=0
cc_478 N_C_M1008_g N_A_1363_127#_c_684_n 0.00167029f $X=8.195 $Y=2.235 $X2=0
+ $Y2=0
cc_479 N_C_M1008_g N_A_1363_127#_c_685_n 0.00262646f $X=8.195 $Y=2.235 $X2=0
+ $Y2=0
cc_480 N_C_M1015_g N_A_1363_127#_c_685_n 0.0129883f $X=8.365 $Y=0.895 $X2=0
+ $Y2=0
cc_481 N_C_M1008_g N_VPWR_c_844_n 0.00830447f $X=8.195 $Y=2.235 $X2=0 $Y2=0
cc_482 N_C_M1011_g N_VPWR_c_845_n 6.76935e-19 $X=7.205 $Y=2.385 $X2=0 $Y2=0
cc_483 N_C_M1008_g N_VPWR_c_845_n 0.00112697f $X=8.195 $Y=2.235 $X2=0 $Y2=0
cc_484 N_C_M1008_g N_VPWR_c_841_n 0.00101825f $X=8.195 $Y=2.235 $X2=0 $Y2=0
cc_485 N_C_c_612_n N_A_402_411#_c_920_n 0.00448381f $X=7.17 $Y=1.385 $X2=0 $Y2=0
cc_486 N_C_M1008_g N_A_402_411#_c_927_n 0.0020996f $X=8.195 $Y=2.235 $X2=0 $Y2=0
cc_487 N_C_c_612_n N_A_402_411#_c_922_n 0.00722171f $X=7.17 $Y=1.385 $X2=0 $Y2=0
cc_488 N_C_M1011_g N_A_402_411#_c_922_n 0.00309609f $X=7.205 $Y=2.385 $X2=0
+ $Y2=0
cc_489 N_C_c_613_n N_A_402_411#_c_922_n 0.014475f $X=8.12 $Y=1.46 $X2=0 $Y2=0
cc_490 N_C_c_614_n N_A_402_411#_c_922_n 0.00180051f $X=7.54 $Y=1.46 $X2=0 $Y2=0
cc_491 N_C_M1008_g N_A_402_411#_c_922_n 0.00277518f $X=8.195 $Y=2.235 $X2=0
+ $Y2=0
cc_492 N_C_M1015_g N_A_402_411#_c_922_n 0.00283089f $X=8.365 $Y=0.895 $X2=0
+ $Y2=0
cc_493 C N_A_402_411#_c_922_n 0.0386599f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_494 N_C_M1011_g N_A_402_411#_c_929_n 0.0028137f $X=7.205 $Y=2.385 $X2=0 $Y2=0
cc_495 N_C_c_613_n N_A_402_411#_c_929_n 0.00586467f $X=8.12 $Y=1.46 $X2=0 $Y2=0
cc_496 N_C_c_614_n N_A_402_411#_c_929_n 0.00181925f $X=7.54 $Y=1.46 $X2=0 $Y2=0
cc_497 C N_A_402_411#_c_929_n 0.015293f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_498 C N_A_425_117#_M1014_d 0.00469864f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_499 N_C_c_612_n N_A_425_117#_c_1100_n 5.14907e-19 $X=7.17 $Y=1.385 $X2=0
+ $Y2=0
cc_500 N_C_c_612_n N_A_425_117#_c_1049_n 0.0110254f $X=7.17 $Y=1.385 $X2=0 $Y2=0
cc_501 N_C_c_612_n N_A_425_117#_c_1051_n 0.00526806f $X=7.17 $Y=1.385 $X2=0
+ $Y2=0
cc_502 N_C_c_614_n N_A_425_117#_c_1051_n 6.26524e-19 $X=7.54 $Y=1.46 $X2=0 $Y2=0
cc_503 C N_A_425_117#_c_1051_n 0.0153748f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_504 N_C_M1015_g N_VGND_c_1176_n 0.00624217f $X=8.365 $Y=0.895 $X2=0 $Y2=0
cc_505 N_C_M1015_g N_VGND_c_1181_n 0.00371502f $X=8.365 $Y=0.895 $X2=0 $Y2=0
cc_506 N_C_M1015_g N_VGND_c_1184_n 0.00453162f $X=8.365 $Y=0.895 $X2=0 $Y2=0
cc_507 N_A_1363_127#_c_688_n N_VPWR_M1008_d 0.0173922f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_508 N_A_1363_127#_c_726_p N_VPWR_M1008_d 0.00894451f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_509 N_A_1363_127#_c_684_n N_VPWR_M1008_d 0.00457966f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_510 N_A_1363_127#_M1009_g N_VPWR_c_844_n 0.0159513f $X=9.06 $Y=2.465 $X2=0
+ $Y2=0
cc_511 N_A_1363_127#_c_688_n N_VPWR_c_844_n 0.022078f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_512 N_A_1363_127#_c_726_p N_VPWR_c_844_n 0.00272347f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_513 N_A_1363_127#_c_684_n N_VPWR_c_844_n 0.021984f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_514 N_A_1363_127#_M1009_g N_VPWR_c_849_n 0.00585385f $X=9.06 $Y=2.465 $X2=0
+ $Y2=0
cc_515 N_A_1363_127#_M1009_g N_VPWR_c_841_n 0.0132612f $X=9.06 $Y=2.465 $X2=0
+ $Y2=0
cc_516 N_A_1363_127#_c_688_n N_A_402_411#_M1011_d 0.00247429f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_517 N_A_1363_127#_c_692_n N_A_402_411#_c_927_n 0.0158392f $X=6.99 $Y=2.11
+ $X2=0 $Y2=0
cc_518 N_A_1363_127#_c_688_n N_A_402_411#_c_927_n 0.0229722f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_519 N_A_1363_127#_c_689_n N_A_402_411#_c_927_n 3.16919e-19 $X=7.105 $Y=2.035
+ $X2=0 $Y2=0
cc_520 N_A_1363_127#_c_682_n N_A_402_411#_c_922_n 0.00766772f $X=6.955 $Y=1.13
+ $X2=0 $Y2=0
cc_521 N_A_1363_127#_c_682_n N_A_402_411#_c_929_n 0.00138018f $X=6.955 $Y=1.13
+ $X2=0 $Y2=0
cc_522 N_A_1363_127#_c_688_n N_A_402_411#_c_929_n 0.022643f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_523 N_A_1363_127#_c_689_n N_A_402_411#_c_929_n 3.27782e-19 $X=7.105 $Y=2.035
+ $X2=0 $Y2=0
cc_524 N_A_1363_127#_c_690_n N_A_402_411#_c_929_n 0.0158392f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_525 N_A_1363_127#_c_682_n N_A_425_117#_c_1047_n 0.00752767f $X=6.955 $Y=1.13
+ $X2=0 $Y2=0
cc_526 N_A_1363_127#_M1001_d N_A_425_117#_c_1049_n 0.00180746f $X=6.815 $Y=0.635
+ $X2=0 $Y2=0
cc_527 N_A_1363_127#_c_682_n N_A_425_117#_c_1049_n 0.0129403f $X=6.955 $Y=1.13
+ $X2=0 $Y2=0
cc_528 N_A_1363_127#_M1012_g X 0.00684657f $X=8.99 $Y=0.685 $X2=0 $Y2=0
cc_529 N_A_1363_127#_c_683_n X 0.0490857f $X=8.845 $Y=1.47 $X2=0 $Y2=0
cc_530 N_A_1363_127#_c_726_p X 0.00646375f $X=8.88 $Y=2.035 $X2=0 $Y2=0
cc_531 N_A_1363_127#_c_685_n X 0.0163799f $X=9.06 $Y=1.47 $X2=0 $Y2=0
cc_532 N_A_1363_127#_M1012_g N_X_c_1159_n 0.0101304f $X=8.99 $Y=0.685 $X2=0
+ $Y2=0
cc_533 N_A_1363_127#_M1012_g X 0.00396245f $X=8.99 $Y=0.685 $X2=0 $Y2=0
cc_534 N_A_1363_127#_c_685_n X 0.00335061f $X=9.06 $Y=1.47 $X2=0 $Y2=0
cc_535 N_A_1363_127#_M1012_g N_VGND_c_1176_n 0.0139969f $X=8.99 $Y=0.685 $X2=0
+ $Y2=0
cc_536 N_A_1363_127#_c_683_n N_VGND_c_1176_n 0.0147357f $X=8.845 $Y=1.47 $X2=0
+ $Y2=0
cc_537 N_A_1363_127#_c_685_n N_VGND_c_1176_n 0.00139834f $X=9.06 $Y=1.47 $X2=0
+ $Y2=0
cc_538 N_A_1363_127#_M1012_g N_VGND_c_1183_n 0.00520813f $X=8.99 $Y=0.685 $X2=0
+ $Y2=0
cc_539 N_A_1363_127#_M1012_g N_VGND_c_1184_n 0.0116184f $X=8.99 $Y=0.685 $X2=0
+ $Y2=0
cc_540 N_A_42_411#_c_768_n N_VPWR_c_842_n 0.0315448f $X=0.355 $Y=2.9 $X2=0 $Y2=0
cc_541 N_A_42_411#_c_768_n N_VPWR_c_847_n 0.0234637f $X=0.355 $Y=2.9 $X2=0 $Y2=0
cc_542 N_A_42_411#_c_768_n N_VPWR_c_841_n 0.0134652f $X=0.355 $Y=2.9 $X2=0 $Y2=0
cc_543 N_A_42_411#_c_760_n N_A_402_411#_c_923_n 0.013646f $X=2.495 $Y=1.51 $X2=0
+ $Y2=0
cc_544 N_A_42_411#_c_761_n N_A_402_411#_c_923_n 6.10459e-19 $X=2 $Y=1.51 $X2=0
+ $Y2=0
cc_545 N_A_42_411#_c_769_n N_A_402_411#_c_923_n 0.0125869f $X=2.66 $Y=2.2 $X2=0
+ $Y2=0
cc_546 N_A_42_411#_M1003_d N_A_402_411#_c_924_n 0.00180746f $X=2.52 $Y=2.055
+ $X2=0 $Y2=0
cc_547 N_A_42_411#_c_769_n N_A_402_411#_c_924_n 0.0163515f $X=2.66 $Y=2.2 $X2=0
+ $Y2=0
cc_548 N_A_42_411#_c_758_n N_A_425_117#_c_1044_n 0.00756924f $X=1.83 $Y=0.65
+ $X2=0 $Y2=0
cc_549 N_A_42_411#_c_759_n N_A_425_117#_c_1044_n 0.0172052f $X=1.915 $Y=1.425
+ $X2=0 $Y2=0
cc_550 N_A_42_411#_c_760_n N_A_425_117#_c_1044_n 0.0201137f $X=2.495 $Y=1.51
+ $X2=0 $Y2=0
cc_551 N_A_42_411#_c_762_n N_A_425_117#_c_1044_n 0.0393534f $X=2.832 $Y=1.068
+ $X2=0 $Y2=0
cc_552 N_A_42_411#_c_762_n N_A_425_117#_c_1045_n 0.0262321f $X=2.832 $Y=1.068
+ $X2=0 $Y2=0
cc_553 N_A_42_411#_c_769_n N_A_425_117#_c_1055_n 0.00741212f $X=2.66 $Y=2.2
+ $X2=0 $Y2=0
cc_554 N_A_42_411#_c_769_n N_A_425_117#_c_1056_n 0.0248237f $X=2.66 $Y=2.2 $X2=0
+ $Y2=0
cc_555 N_A_42_411#_c_769_n N_A_425_117#_c_1053_n 0.0116093f $X=2.66 $Y=2.2 $X2=0
+ $Y2=0
cc_556 N_A_42_411#_c_762_n N_A_425_117#_c_1053_n 0.025159f $X=2.832 $Y=1.068
+ $X2=0 $Y2=0
cc_557 N_A_42_411#_c_763_n N_A_425_117#_c_1053_n 0.00794608f $X=2.74 $Y=1.425
+ $X2=0 $Y2=0
cc_558 N_A_42_411#_c_766_n N_A_425_117#_c_1053_n 0.00819057f $X=2.66 $Y=1.51
+ $X2=0 $Y2=0
cc_559 N_A_42_411#_c_758_n N_VGND_M1007_d 0.0154172f $X=1.83 $Y=0.65 $X2=-0.19
+ $Y2=-0.245
cc_560 N_A_42_411#_c_758_n N_VGND_c_1177_n 0.0232826f $X=1.83 $Y=0.65 $X2=0
+ $Y2=0
cc_561 N_A_42_411#_c_758_n N_VGND_c_1178_n 0.0035903f $X=1.83 $Y=0.65 $X2=0
+ $Y2=0
cc_562 N_A_42_411#_c_764_n N_VGND_c_1178_n 0.0120453f $X=0.347 $Y=0.65 $X2=0
+ $Y2=0
cc_563 N_A_42_411#_c_758_n N_VGND_c_1179_n 0.0188844f $X=1.83 $Y=0.65 $X2=0
+ $Y2=0
cc_564 N_A_42_411#_c_758_n N_VGND_c_1184_n 0.0338206f $X=1.83 $Y=0.65 $X2=0
+ $Y2=0
cc_565 N_A_42_411#_c_764_n N_VGND_c_1184_n 0.0163573f $X=0.347 $Y=0.65 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_843_n N_A_425_117#_c_1054_n 0.0314551f $X=5.425 $Y=1.93 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_843_n N_A_425_117#_c_1057_n 0.00251938f $X=5.425 $Y=1.93 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_843_n N_A_425_117#_c_1052_n 0.0555928f $X=5.425 $Y=1.93 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_845_n N_A_425_117#_c_1052_n 0.00677041f $X=8.44 $Y=3.33 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_841_n N_A_425_117#_c_1052_n 0.00826788f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_841_n N_X_M1009_d 0.0042346f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_572 N_VPWR_c_849_n X 0.0187372f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_573 N_VPWR_c_841_n X 0.0109447f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_574 N_A_402_411#_c_924_n N_A_425_117#_M1013_d 0.00496055f $X=3.54 $Y=2.63
+ $X2=0 $Y2=0
cc_575 N_A_402_411#_c_917_n N_A_425_117#_c_1045_n 0.0145115f $X=3.71 $Y=0.35
+ $X2=0 $Y2=0
cc_576 N_A_402_411#_M1001_s N_A_425_117#_c_1047_n 0.0119184f $X=6.11 $Y=0.635
+ $X2=0 $Y2=0
cc_577 N_A_402_411#_c_919_n N_A_425_117#_c_1047_n 0.0159025f $X=6.215 $Y=0.775
+ $X2=0 $Y2=0
cc_578 N_A_402_411#_M1001_s N_A_425_117#_c_1048_n 4.91001e-19 $X=6.11 $Y=0.635
+ $X2=0 $Y2=0
cc_579 N_A_402_411#_c_918_n N_A_425_117#_c_1048_n 0.0165903f $X=6.09 $Y=0.86
+ $X2=0 $Y2=0
cc_580 N_A_402_411#_c_919_n N_A_425_117#_c_1048_n 0.00395819f $X=6.215 $Y=0.775
+ $X2=0 $Y2=0
cc_581 N_A_402_411#_M1001_s N_A_425_117#_c_1100_n 0.00856108f $X=6.11 $Y=0.635
+ $X2=0 $Y2=0
cc_582 N_A_402_411#_c_919_n N_A_425_117#_c_1100_n 0.0124375f $X=6.215 $Y=0.775
+ $X2=0 $Y2=0
cc_583 N_A_402_411#_c_920_n N_A_425_117#_c_1049_n 0.0350745f $X=7.715 $Y=0.35
+ $X2=0 $Y2=0
cc_584 N_A_402_411#_M1001_s N_A_425_117#_c_1050_n 0.00169457f $X=6.11 $Y=0.635
+ $X2=0 $Y2=0
cc_585 N_A_402_411#_c_919_n N_A_425_117#_c_1050_n 0.0137281f $X=6.215 $Y=0.775
+ $X2=0 $Y2=0
cc_586 N_A_402_411#_c_920_n N_A_425_117#_c_1050_n 0.0127436f $X=7.715 $Y=0.35
+ $X2=0 $Y2=0
cc_587 N_A_402_411#_c_920_n N_A_425_117#_c_1051_n 0.0178501f $X=7.715 $Y=0.35
+ $X2=0 $Y2=0
cc_588 N_A_402_411#_c_922_n N_A_425_117#_c_1051_n 0.0225801f $X=7.61 $Y=1.895
+ $X2=0 $Y2=0
cc_589 N_A_402_411#_c_924_n N_A_425_117#_c_1054_n 0.00575441f $X=3.54 $Y=2.63
+ $X2=0 $Y2=0
cc_590 N_A_402_411#_c_915_n N_A_425_117#_c_1054_n 0.0189311f $X=3.625 $Y=0.73
+ $X2=0 $Y2=0
cc_591 N_A_402_411#_c_924_n N_A_425_117#_c_1055_n 0.0023602f $X=3.54 $Y=2.63
+ $X2=0 $Y2=0
cc_592 N_A_402_411#_c_915_n N_A_425_117#_c_1055_n 5.31975e-19 $X=3.625 $Y=0.73
+ $X2=0 $Y2=0
cc_593 N_A_402_411#_c_924_n N_A_425_117#_c_1056_n 0.0214178f $X=3.54 $Y=2.63
+ $X2=0 $Y2=0
cc_594 N_A_402_411#_c_915_n N_A_425_117#_c_1053_n 0.117409f $X=3.625 $Y=0.73
+ $X2=0 $Y2=0
cc_595 N_A_402_411#_c_916_n N_VGND_M1005_d 0.00281172f $X=5.26 $Y=0.35 $X2=0
+ $Y2=0
cc_596 N_A_402_411#_c_961_n N_VGND_M1005_d 0.00528907f $X=5.345 $Y=0.775 $X2=0
+ $Y2=0
cc_597 N_A_402_411#_c_918_n N_VGND_M1005_d 0.0192743f $X=6.09 $Y=0.86 $X2=0
+ $Y2=0
cc_598 N_A_402_411#_c_965_n N_VGND_M1005_d 8.95698e-19 $X=5.43 $Y=0.86 $X2=0
+ $Y2=0
cc_599 N_A_402_411#_c_916_n N_VGND_c_1175_n 0.0136053f $X=5.26 $Y=0.35 $X2=0
+ $Y2=0
cc_600 N_A_402_411#_c_961_n N_VGND_c_1175_n 0.0114341f $X=5.345 $Y=0.775 $X2=0
+ $Y2=0
cc_601 N_A_402_411#_c_918_n N_VGND_c_1175_n 0.0187598f $X=6.09 $Y=0.86 $X2=0
+ $Y2=0
cc_602 N_A_402_411#_c_919_n N_VGND_c_1175_n 0.0103109f $X=6.215 $Y=0.775 $X2=0
+ $Y2=0
cc_603 N_A_402_411#_c_921_n N_VGND_c_1175_n 0.0119254f $X=6.34 $Y=0.35 $X2=0
+ $Y2=0
cc_604 N_A_402_411#_c_920_n N_VGND_c_1176_n 0.00591685f $X=7.715 $Y=0.35 $X2=0
+ $Y2=0
cc_605 N_A_402_411#_c_922_n N_VGND_c_1176_n 0.00714036f $X=7.61 $Y=1.895 $X2=0
+ $Y2=0
cc_606 N_A_402_411#_c_916_n N_VGND_c_1179_n 0.100657f $X=5.26 $Y=0.35 $X2=0
+ $Y2=0
cc_607 N_A_402_411#_c_917_n N_VGND_c_1179_n 0.0114574f $X=3.71 $Y=0.35 $X2=0
+ $Y2=0
cc_608 N_A_402_411#_c_920_n N_VGND_c_1181_n 0.0947801f $X=7.715 $Y=0.35 $X2=0
+ $Y2=0
cc_609 N_A_402_411#_c_921_n N_VGND_c_1181_n 0.0168561f $X=6.34 $Y=0.35 $X2=0
+ $Y2=0
cc_610 N_A_402_411#_c_916_n N_VGND_c_1184_n 0.0594452f $X=5.26 $Y=0.35 $X2=0
+ $Y2=0
cc_611 N_A_402_411#_c_917_n N_VGND_c_1184_n 0.00589978f $X=3.71 $Y=0.35 $X2=0
+ $Y2=0
cc_612 N_A_402_411#_c_918_n N_VGND_c_1184_n 0.0159461f $X=6.09 $Y=0.86 $X2=0
+ $Y2=0
cc_613 N_A_402_411#_c_920_n N_VGND_c_1184_n 0.0579576f $X=7.715 $Y=0.35 $X2=0
+ $Y2=0
cc_614 N_A_402_411#_c_921_n N_VGND_c_1184_n 0.00967329f $X=6.34 $Y=0.35 $X2=0
+ $Y2=0
cc_615 N_A_425_117#_c_1045_n N_VGND_c_1179_n 0.0569889f $X=3.19 $Y=0.35 $X2=0
+ $Y2=0
cc_616 N_A_425_117#_c_1046_n N_VGND_c_1179_n 0.01685f $X=2.43 $Y=0.35 $X2=0
+ $Y2=0
cc_617 N_A_425_117#_c_1045_n N_VGND_c_1184_n 0.0311477f $X=3.19 $Y=0.35 $X2=0
+ $Y2=0
cc_618 N_A_425_117#_c_1046_n N_VGND_c_1184_n 0.00867614f $X=2.43 $Y=0.35 $X2=0
+ $Y2=0
cc_619 N_X_c_1159_n N_VGND_c_1176_n 0.032876f $X=9.205 $Y=0.43 $X2=0 $Y2=0
cc_620 N_X_c_1159_n N_VGND_c_1183_n 0.0268376f $X=9.205 $Y=0.43 $X2=0 $Y2=0
cc_621 N_X_c_1159_n N_VGND_c_1184_n 0.0166333f $X=9.205 $Y=0.43 $X2=0 $Y2=0
