* File: sky130_fd_sc_lp__nor4_0.pex.spice
* Created: Wed Sep  2 10:10:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4_0%A 3 6 9 13 14 17 19 20 24
r39 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.525
+ $Y=1.355 $X2=0.525 $Y2=1.355
r40 20 25 8.71359 $w=4.08e-07 $l=3.1e-07 $layer=LI1_cond $X=0.635 $Y=1.665
+ $X2=0.635 $Y2=1.355
r41 19 25 1.6865 $w=4.08e-07 $l=6e-08 $layer=LI1_cond $X=0.635 $Y=1.295
+ $X2=0.635 $Y2=1.355
r42 15 17 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.615 $Y=2.175
+ $X2=0.795 $Y2=2.175
r43 13 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.525 $Y=1.695
+ $X2=0.525 $Y2=1.355
r44 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.695
+ $X2=0.525 $Y2=1.86
r45 12 24 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.19
+ $X2=0.525 $Y2=1.355
r46 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.795 $Y=2.25
+ $X2=0.795 $Y2=2.175
r47 7 9 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.795 $Y=2.25
+ $X2=0.795 $Y2=2.735
r48 6 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=2.1
+ $X2=0.615 $Y2=2.175
r49 6 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.615 $Y=2.1
+ $X2=0.615 $Y2=1.86
r50 3 12 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.575 $Y=0.56
+ $X2=0.575 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_0%B 3 7 11 12 13 14 18
r38 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.095
+ $Y=1.355 $X2=1.095 $Y2=1.355
r39 14 19 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=1.187 $Y=1.665
+ $X2=1.187 $Y2=1.355
r40 13 19 1.94779 $w=3.53e-07 $l=6e-08 $layer=LI1_cond $X=1.187 $Y=1.295
+ $X2=1.187 $Y2=1.355
r41 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.095 $Y=1.695
+ $X2=1.095 $Y2=1.355
r42 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.695
+ $X2=1.095 $Y2=1.86
r43 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.19
+ $X2=1.095 $Y2=1.355
r44 7 12 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.185 $Y=2.735
+ $X2=1.185 $Y2=1.86
r45 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.005 $Y=0.56
+ $X2=1.005 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_0%C 2 5 9 11 12 13 17
r37 17 19 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.355
+ $X2=1.675 $Y2=1.19
r38 12 13 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.682 $Y=1.295
+ $X2=1.682 $Y2=1.665
r39 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.665
+ $Y=1.355 $X2=1.665 $Y2=1.355
r40 9 19 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.775 $Y=0.56
+ $X2=1.775 $Y2=1.19
r41 5 11 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.575 $Y=2.735
+ $X2=1.575 $Y2=1.86
r42 2 11 48.0802 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.675 $Y=1.685
+ $X2=1.675 $Y2=1.86
r43 1 17 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=1.675 $Y=1.365
+ $X2=1.675 $Y2=1.355
r44 1 2 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.675 $Y=1.365
+ $X2=1.675 $Y2=1.685
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_0%D 3 6 9 14 15 16 17 24 25 26 41
r38 28 41 1.33755 $w=4.63e-07 $l=5.2e-08 $layer=LI1_cond $X=2.562 $Y=1.613
+ $X2=2.562 $Y2=1.665
r39 24 27 73.0393 $w=6e-07 $l=5.05e-07 $layer=POLY_cond $X=2.36 $Y=1.045
+ $X2=2.36 $Y2=1.55
r40 24 26 49.4885 $w=6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.045
+ $X2=2.36 $Y2=0.88
r41 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.495
+ $Y=1.045 $X2=2.495 $Y2=1.045
r42 16 17 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.655 $Y=2.035
+ $X2=2.655 $Y2=2.405
r43 16 43 7.82015 $w=2.78e-07 $l=1.9e-07 $layer=LI1_cond $X=2.655 $Y=2.035
+ $X2=2.655 $Y2=1.845
r44 15 43 6.09719 $w=4.63e-07 $l=1.64e-07 $layer=LI1_cond $X=2.562 $Y=1.681
+ $X2=2.562 $Y2=1.845
r45 15 41 0.411554 $w=4.63e-07 $l=1.6e-08 $layer=LI1_cond $X=2.562 $Y=1.681
+ $X2=2.562 $Y2=1.665
r46 15 28 0.437276 $w=4.63e-07 $l=1.7e-08 $layer=LI1_cond $X=2.562 $Y=1.596
+ $X2=2.562 $Y2=1.613
r47 14 15 7.74236 $w=4.63e-07 $l=3.01e-07 $layer=LI1_cond $X=2.562 $Y=1.295
+ $X2=2.562 $Y2=1.596
r48 14 25 6.43053 $w=4.63e-07 $l=2.5e-07 $layer=LI1_cond $X=2.562 $Y=1.295
+ $X2=2.562 $Y2=1.045
r49 9 26 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.205 $Y=0.56
+ $X2=2.205 $Y2=0.88
r50 6 10 95.8872 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=2.152 $Y=2.175
+ $X2=1.965 $Y2=2.175
r51 6 27 203.183 $w=1.85e-07 $l=5.5e-07 $layer=POLY_cond $X=2.152 $Y=2.1
+ $X2=2.152 $Y2=1.55
r52 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.965 $Y=2.25
+ $X2=1.965 $Y2=2.175
r53 1 3 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.965 $Y=2.25
+ $X2=1.965 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_0%VPWR 1 6 8 10 17 18 21
r22 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r23 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r24 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.58 $Y2=3.33
r25 15 17 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=2.64 $Y2=3.33
r26 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.58 $Y2=3.33
r29 10 12 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 8 18 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 8 22 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.58 $Y=3.245 $X2=0.58
+ $Y2=3.33
r33 4 6 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.58 $Y=3.245
+ $X2=0.58 $Y2=2.57
r34 1 6 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.455
+ $Y=2.415 $X2=0.58 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_0%Y 1 2 3 11 12 13 16 20 22 23 24 25 26 32 41
r63 25 26 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.93 $X2=1.68
+ $Y2=0.93
r64 25 34 19.7172 $w=1.78e-07 $l=3.2e-07 $layer=LI1_cond $X=1.2 $Y=0.93 $X2=0.88
+ $Y2=0.93
r65 24 32 5.28486 $w=1.8e-07 $l=9.2e-08 $layer=LI1_cond $X=0.787 $Y=0.93
+ $X2=0.695 $Y2=0.93
r66 24 34 5.28486 $w=1.8e-07 $l=9.3e-08 $layer=LI1_cond $X=0.787 $Y=0.93
+ $X2=0.88 $Y2=0.93
r67 24 41 12.5325 $w=2.93e-07 $l=2.8e-07 $layer=LI1_cond $X=0.787 $Y=0.84
+ $X2=0.787 $Y2=0.56
r68 24 32 1.84848 $w=1.78e-07 $l=3e-08 $layer=LI1_cond $X=0.665 $Y=0.93
+ $X2=0.695 $Y2=0.93
r69 23 26 13.2475 $w=1.78e-07 $l=2.15e-07 $layer=LI1_cond $X=1.895 $Y=0.93
+ $X2=1.68 $Y2=0.93
r70 22 24 24.9545 $w=1.78e-07 $l=4.05e-07 $layer=LI1_cond $X=0.26 $Y=0.93
+ $X2=0.665 $Y2=0.93
r71 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.18 $Y=2.225
+ $X2=2.18 $Y2=2.56
r72 14 23 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=1.99 $Y=0.84
+ $X2=1.895 $Y2=0.93
r73 14 16 16.3445 $w=1.88e-07 $l=2.8e-07 $layer=LI1_cond $X=1.99 $Y=0.84
+ $X2=1.99 $Y2=0.56
r74 12 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.015 $Y=2.14
+ $X2=2.18 $Y2=2.225
r75 12 13 114.497 $w=1.68e-07 $l=1.755e-06 $layer=LI1_cond $X=2.015 $Y=2.14
+ $X2=0.26 $Y2=2.14
r76 11 13 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.172 $Y=2.055
+ $X2=0.26 $Y2=2.14
r77 10 22 6.81825 $w=1.8e-07 $l=1.2657e-07 $layer=LI1_cond $X=0.172 $Y=1.02
+ $X2=0.26 $Y2=0.93
r78 10 11 65.5948 $w=1.73e-07 $l=1.035e-06 $layer=LI1_cond $X=0.172 $Y=1.02
+ $X2=0.172 $Y2=2.055
r79 3 20 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.04
+ $Y=2.415 $X2=2.18 $Y2=2.56
r80 2 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.85
+ $Y=0.35 $X2=1.99 $Y2=0.56
r81 1 41 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.35 $X2=0.79 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_0%VGND 1 2 3 10 12 16 18 19 20 21 23 34
r35 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r36 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r37 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r38 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 28 30 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.725 $Y=0 $X2=2.16
+ $Y2=0
r40 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r41 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r42 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 24 36 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.262
+ $Y2=0
r44 24 26 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.72
+ $Y2=0
r45 23 43 9.92302 $w=6.73e-07 $l=5.6e-07 $layer=LI1_cond $X=1.387 $Y=0 $X2=1.387
+ $Y2=0.56
r46 23 28 9.08255 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=1.387 $Y=0 $X2=1.725
+ $Y2=0
r47 23 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r48 23 26 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=0.72
+ $Y2=0
r49 21 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r50 21 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r51 19 30 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.16
+ $Y2=0
r52 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.42
+ $Y2=0
r53 18 33 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.64
+ $Y2=0
r54 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.42
+ $Y2=0
r55 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=0.085
+ $X2=2.42 $Y2=0
r56 14 16 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=2.42 $Y=0.085
+ $X2=2.42 $Y2=0.56
r57 10 36 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.262 $Y2=0
r58 10 12 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.36 $Y2=0.56
r59 3 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.35 $X2=2.42 $Y2=0.56
r60 2 43 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=1.08 $Y=0.35
+ $X2=1.56 $Y2=0.56
r61 1 12 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.35 $X2=0.36 $Y2=0.56
.ends

