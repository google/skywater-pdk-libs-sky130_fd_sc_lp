* File: sky130_fd_sc_lp__inv_lp.pex.spice
* Created: Fri Aug 28 10:38:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INV_LP%A 3 7 11 13 15 22
r25 22 24 65.5974 $w=5.4e-07 $l=5.05e-07 $layer=POLY_cond $X=0.74 $Y=1.12
+ $X2=0.74 $Y2=1.625
r26 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.635
+ $Y=1.12 $X2=0.635 $Y2=1.12
r27 15 23 1.23232 $w=8.23e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.367
+ $X2=0.635 $Y2=1.367
r28 13 23 5.72668 $w=8.23e-07 $l=3.95e-07 $layer=LI1_cond $X=0.24 $Y=1.367
+ $X2=0.635 $Y2=1.367
r29 9 22 31.5348 $w=2.7e-07 $l=2.64953e-07 $layer=POLY_cond $X=0.935 $Y=0.955
+ $X2=0.74 $Y2=1.12
r30 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.935 $Y=0.955
+ $X2=0.935 $Y2=0.545
r31 7 24 212.428 $w=2.5e-07 $l=8.55e-07 $layer=POLY_cond $X=0.885 $Y=2.48
+ $X2=0.885 $Y2=1.625
r32 1 22 31.5348 $w=2.7e-07 $l=2.64953e-07 $layer=POLY_cond $X=0.545 $Y=0.955
+ $X2=0.74 $Y2=1.12
r33 1 3 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.545 $Y=0.955
+ $X2=0.545 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__INV_LP%VPWR 1 6 11 12 13 20 21
r14 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r15 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r16 13 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r17 13 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r18 11 16 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.24 $Y2=3.33
r19 11 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.62 $Y2=3.33
r20 10 20 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=1.2 $Y2=3.33
r21 10 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.62 $Y2=3.33
r22 6 9 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.62 $Y=2.125 $X2=0.62
+ $Y2=2.835
r23 4 12 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.62 $Y=3.245 $X2=0.62
+ $Y2=3.33
r24 4 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.62 $Y=3.245 $X2=0.62
+ $Y2=2.835
r25 1 9 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.475
+ $Y=1.98 $X2=0.62 $Y2=2.835
r26 1 6 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.475
+ $Y=1.98 $X2=0.62 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_LP__INV_LP%Y 1 2 7 8 9 10 11 12 13 46
r17 46 47 3.68958 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.15 $Y=2.035
+ $X2=1.15 $Y2=1.96
r18 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=2.405
+ $X2=1.15 $Y2=2.775
r19 12 33 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.15 $Y=2.405
+ $X2=1.15 $Y2=2.125
r20 11 33 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=2.04
+ $X2=1.15 $Y2=2.125
r21 11 46 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=2.04 $X2=1.15
+ $Y2=2.035
r22 11 47 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=1.955 $X2=1.2
+ $Y2=1.96
r23 10 11 14.5308 $w=2.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.2
+ $Y2=1.955
r24 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.665
r25 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.925 $X2=1.2
+ $Y2=1.295
r26 8 44 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.2 $Y=0.925 $X2=1.2
+ $Y2=0.775
r27 7 44 9.10257 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.15 $Y=0.545
+ $X2=1.15 $Y2=0.775
r28 2 13 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.98 $X2=1.15 $Y2=2.835
r29 2 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.98 $X2=1.15 $Y2=2.125
r30 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.335 $X2=1.15 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__INV_LP%VGND 1 4 6 8 12 13
r14 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r15 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r16 10 16 4.62984 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=0.495 $Y=0 $X2=0.247
+ $Y2=0
r17 10 12 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.495 $Y=0 $X2=1.2
+ $Y2=0
r18 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r19 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r20 4 16 3.13634 $w=3.3e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.247 $Y2=0
r21 4 6 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.33 $Y=0.085 $X2=0.33
+ $Y2=0.545
r22 1 6 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.335 $X2=0.33 $Y2=0.545
.ends

