* File: sky130_fd_sc_lp__a221o_0.pex.spice
* Created: Fri Aug 28 09:52:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221O_0%A_72_312# 1 2 3 12 16 20 21 22 24 25 29 30
+ 31 32 35 38 39 40 41 43 47 49
c123 25 0 1.90286e-19 $X=0.525 $Y=1.725
r124 45 47 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=3.585 $Y=2.015
+ $X2=3.585 $Y2=2.29
r125 41 58 21.3337 $w=1.68e-07 $l=3.27e-07 $layer=LI1_cond $X=3.427 $Y=0.73
+ $X2=3.1 $Y2=0.73
r126 41 43 7.81317 $w=2.93e-07 $l=2e-07 $layer=LI1_cond $X=3.427 $Y=0.645
+ $X2=3.427 $Y2=0.445
r127 39 45 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.455 $Y=1.93
+ $X2=3.585 $Y2=2.015
r128 39 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.455 $Y=1.93
+ $X2=3.19 $Y2=1.93
r129 38 40 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.1 $Y=1.845
+ $X2=3.19 $Y2=1.93
r130 37 58 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.815
+ $X2=3.1 $Y2=0.73
r131 37 38 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=3.1 $Y=0.815
+ $X2=3.1 $Y2=1.845
r132 36 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.73
+ $X2=2.525 $Y2=0.73
r133 35 58 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.01 $Y=0.73 $X2=3.1
+ $Y2=0.73
r134 35 36 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.01 $Y=0.73 $X2=2.61
+ $Y2=0.73
r135 32 52 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.285 $Y=0.445
+ $X2=1.285 $Y2=0.81
r136 32 34 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.37 $Y=0.445
+ $X2=2.08 $Y2=0.445
r137 31 56 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.525 $Y=0.445
+ $X2=2.525 $Y2=0.73
r138 31 34 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.44 $Y=0.445
+ $X2=2.08 $Y2=0.445
r139 29 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.81
+ $X2=1.285 $Y2=0.81
r140 29 30 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.2 $Y=0.81
+ $X2=0.675 $Y2=0.81
r141 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.59 $Y=0.895
+ $X2=0.675 $Y2=0.81
r142 27 49 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=0.59 $Y=0.895
+ $X2=0.59 $Y2=1.56
r143 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.525
+ $Y=1.725 $X2=0.525 $Y2=1.725
r144 22 49 6.63891 $w=2.33e-07 $l=1.17e-07 $layer=LI1_cond $X=0.557 $Y=1.677
+ $X2=0.557 $Y2=1.56
r145 22 24 2.35393 $w=2.33e-07 $l=4.8e-08 $layer=LI1_cond $X=0.557 $Y=1.677
+ $X2=0.557 $Y2=1.725
r146 20 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.525 $Y=2.065
+ $X2=0.525 $Y2=1.725
r147 20 21 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=2.065
+ $X2=0.525 $Y2=2.23
r148 19 25 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.56
+ $X2=0.525 $Y2=1.725
r149 16 19 571.734 $w=1.5e-07 $l=1.115e-06 $layer=POLY_cond $X=0.585 $Y=0.445
+ $X2=0.585 $Y2=1.56
r150 12 21 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.555 $Y=2.74
+ $X2=0.555 $Y2=2.23
r151 3 47 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.41
+ $Y=2.145 $X2=3.55 $Y2=2.29
r152 2 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.27
+ $Y=0.235 $X2=3.41 $Y2=0.445
r153 1 34 91 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=2 $X=1.59
+ $Y=0.235 $X2=2.08 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%A2 3 7 11 12 13 16
c45 13 0 1.90286e-19 $X=1.2 $Y=1.295
r46 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.065
+ $Y=1.16 $X2=1.065 $Y2=1.16
r47 13 17 2.93583 $w=5.48e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=1.34
+ $X2=1.065 $Y2=1.34
r48 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.065 $Y=1.5
+ $X2=1.065 $Y2=1.16
r49 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.5
+ $X2=1.065 $Y2=1.665
r50 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=0.995
+ $X2=1.065 $Y2=1.16
r51 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.155 $Y=0.445
+ $X2=1.155 $Y2=0.995
r52 3 12 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=1.005 $Y=2.74
+ $X2=1.005 $Y2=1.665
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%A1 3 7 10 12 15 17 18 19 23
c47 7 0 8.38428e-20 $X=1.515 $Y=0.445
r48 23 25 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.1
+ $X2=1.62 $Y2=0.935
r49 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.635
+ $Y=1.1 $X2=1.635 $Y2=1.1
r50 19 24 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.692 $Y=1.295
+ $X2=1.692 $Y2=1.1
r51 18 24 6.61238 $w=3.03e-07 $l=1.75e-07 $layer=LI1_cond $X=1.692 $Y=0.925
+ $X2=1.692 $Y2=1.1
r52 13 15 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=1.435 $Y=1.98
+ $X2=1.515 $Y2=1.98
r53 12 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.515 $Y=1.905
+ $X2=1.515 $Y2=1.98
r54 12 17 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.515 $Y=1.905
+ $X2=1.515 $Y2=1.605
r55 10 17 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.62 $Y=1.425
+ $X2=1.62 $Y2=1.605
r56 9 23 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.62 $Y=1.115
+ $X2=1.62 $Y2=1.1
r57 9 10 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.62 $Y=1.115
+ $X2=1.62 $Y2=1.425
r58 7 25 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.515 $Y=0.445
+ $X2=1.515 $Y2=0.935
r59 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.435 $Y=2.055
+ $X2=1.435 $Y2=1.98
r60 1 3 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=1.435 $Y=2.055
+ $X2=1.435 $Y2=2.74
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%B1 2 5 9 11 12 16
c36 11 0 1.85865e-19 $X=2.16 $Y=0.925
r37 16 18 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.005
+ $X2=2.19 $Y2=0.84
r38 11 12 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.142 $Y=0.925
+ $X2=2.142 $Y2=1.295
r39 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.175
+ $Y=1.005 $X2=2.175 $Y2=1.005
r40 7 9 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.405 $Y=1.77
+ $X2=2.405 $Y2=2.465
r41 5 18 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.295 $Y=0.445
+ $X2=2.295 $Y2=0.84
r42 2 7 72.8797 $w=2.91e-07 $l=5.36843e-07 $layer=POLY_cond $X=2.19 $Y=1.33
+ $X2=2.405 $Y2=1.77
r43 1 16 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=2.19 $Y=1.02 $X2=2.19
+ $Y2=1.005
r44 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=2.19 $Y=1.02 $X2=2.19
+ $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%B2 3 7 9 12 13
c36 7 0 1.02022e-19 $X=2.835 $Y=2.465
r37 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.215
+ $X2=2.745 $Y2=1.38
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.215
+ $X2=2.745 $Y2=1.05
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.745
+ $Y=1.215 $X2=2.745 $Y2=1.215
r40 9 13 2.34744 $w=5.33e-07 $l=1.05e-07 $layer=LI1_cond $X=2.64 $Y=1.317
+ $X2=2.745 $Y2=1.317
r41 7 15 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=2.835 $Y=2.465
+ $X2=2.835 $Y2=1.38
r42 3 14 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=2.655 $Y=0.445
+ $X2=2.655 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%C1 3 7 9 12
c31 7 0 1.03888e-19 $X=3.335 $Y=2.465
r32 12 15 83.3779 $w=4.9e-07 $l=5.05e-07 $layer=POLY_cond $X=3.365 $Y=1.16
+ $X2=3.365 $Y2=1.665
r33 12 14 46.2534 $w=4.9e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.16
+ $X2=3.365 $Y2=0.995
r34 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.445
+ $Y=1.16 $X2=3.445 $Y2=1.16
r35 9 13 2.76705 $w=6.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.6 $Y=1.33
+ $X2=3.445 $Y2=1.33
r36 7 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.335 $Y=2.465
+ $X2=3.335 $Y2=1.665
r37 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.195 $Y=0.445
+ $X2=3.195 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%X 1 2 12 13 14 15 16 35 38
r25 23 38 1.27004 $w=2.43e-07 $l=2.7e-08 $layer=LI1_cond $X=0.212 $Y=1.268
+ $X2=0.212 $Y2=1.295
r26 16 40 3.9381 $w=2.43e-07 $l=6.6e-08 $layer=LI1_cond $X=0.212 $Y=1.324
+ $X2=0.212 $Y2=1.39
r27 16 38 1.36412 $w=2.43e-07 $l=2.9e-08 $layer=LI1_cond $X=0.212 $Y=1.324
+ $X2=0.212 $Y2=1.295
r28 16 23 1.36412 $w=2.43e-07 $l=2.9e-08 $layer=LI1_cond $X=0.212 $Y=1.239
+ $X2=0.212 $Y2=1.268
r29 15 16 14.7701 $w=2.43e-07 $l=3.14e-07 $layer=LI1_cond $X=0.212 $Y=0.925
+ $X2=0.212 $Y2=1.239
r30 14 35 5.44791 $w=2.73e-07 $l=1.3e-07 $layer=LI1_cond $X=0.24 $Y=0.417
+ $X2=0.37 $Y2=0.417
r31 14 30 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=0.24 $Y=0.417
+ $X2=0.212 $Y2=0.417
r32 14 30 1.43368 $w=2.45e-07 $l=1.38e-07 $layer=LI1_cond $X=0.212 $Y=0.555
+ $X2=0.212 $Y2=0.417
r33 14 15 15.4286 $w=2.43e-07 $l=3.28e-07 $layer=LI1_cond $X=0.212 $Y=0.597
+ $X2=0.212 $Y2=0.925
r34 13 40 62.2323 $w=1.78e-07 $l=1.01e-06 $layer=LI1_cond $X=0.18 $Y=2.4
+ $X2=0.18 $Y2=1.39
r35 12 13 8.22996 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.282 $Y=2.565
+ $X2=0.282 $Y2=2.4
r36 2 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.215
+ $Y=2.42 $X2=0.34 $Y2=2.565
r37 1 35 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%VPWR 1 2 11 15 17 19 29 30 33 36
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 27 30 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r46 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 24 36 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.667 $Y2=3.33
r48 24 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 23 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 20 33 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.785 $Y2=3.33
r53 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 19 36 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=1.52 $Y=3.33
+ $X2=1.667 $Y2=3.33
r55 19 22 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.52 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 17 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 17 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 13 36 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.667 $Y=3.245
+ $X2=1.667 $Y2=3.33
r59 13 15 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=1.667 $Y=3.245
+ $X2=1.667 $Y2=2.565
r60 9 33 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r61 9 11 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.565
r62 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.51
+ $Y=2.42 $X2=1.65 $Y2=2.565
r63 1 11 300 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=2 $X=0.63
+ $Y=2.42 $X2=0.79 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%A_216_484# 1 2 9 11 12 15
c37 11 0 1.03888e-19 $X=2.455 $Y=1.87
r38 13 15 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.62 $Y=1.955
+ $X2=2.62 $Y2=2.27
r39 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.455 $Y=1.87
+ $X2=2.62 $Y2=1.955
r40 11 12 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.455 $Y=1.87
+ $X2=1.35 $Y2=1.87
r41 7 12 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=1.222 $Y=1.955
+ $X2=1.35 $Y2=1.87
r42 7 9 26.6644 $w=2.53e-07 $l=5.9e-07 $layer=LI1_cond $X=1.222 $Y=1.955
+ $X2=1.222 $Y2=2.545
r43 2 15 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=2.145 $X2=2.62 $Y2=2.27
r44 1 9 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=2.42 $X2=1.22 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%A_409_429# 1 2 9 11 12 15
r25 13 15 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=3.12 $Y=2.905
+ $X2=3.12 $Y2=2.3
r26 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=3.12 $Y2=2.905
r27 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=2.285 $Y2=2.99
r28 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.145 $Y=2.905
+ $X2=2.285 $Y2=2.99
r29 7 9 24.901 $w=2.78e-07 $l=6.05e-07 $layer=LI1_cond $X=2.145 $Y=2.905
+ $X2=2.145 $Y2=2.3
r30 2 15 300 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=2.145 $X2=3.12 $Y2=2.3
r31 1 9 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=2.145 $X2=2.17 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_0%VGND 1 2 11 15 18 19 20 30 31 34
r49 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r50 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r52 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r53 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r54 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r55 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r56 22 34 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.872
+ $Y2=0
r57 22 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.2
+ $Y2=0
r58 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r59 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r60 18 27 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.64
+ $Y2=0
r61 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.945
+ $Y2=0
r62 17 30 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.11 $Y=0 $X2=3.6
+ $Y2=0
r63 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=0 $X2=2.945
+ $Y2=0
r64 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0
r65 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0.36
r66 9 34 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.872 $Y=0.085
+ $X2=0.872 $Y2=0
r67 9 11 11.1586 $w=3.13e-07 $l=3.05e-07 $layer=LI1_cond $X=0.872 $Y=0.085
+ $X2=0.872 $Y2=0.39
r68 2 15 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.235 $X2=2.945 $Y2=0.36
r69 1 11 182 $w=1.7e-07 $l=2.71662e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.235 $X2=0.865 $Y2=0.39
.ends

