* File: sky130_fd_sc_lp__a32o_4.pxi.spice
* Created: Wed Sep  2 09:27:48 2020
* 
x_PM_SKY130_FD_SC_LP__A32O_4%A_101_21# N_A_101_21#_M1015_d N_A_101_21#_M1009_d
+ N_A_101_21#_M1024_d N_A_101_21#_M1003_s N_A_101_21#_M1004_g
+ N_A_101_21#_M1000_g N_A_101_21#_M1014_g N_A_101_21#_M1011_g
+ N_A_101_21#_M1017_g N_A_101_21#_M1016_g N_A_101_21#_M1019_g
+ N_A_101_21#_M1021_g N_A_101_21#_c_141_n N_A_101_21#_c_142_n
+ N_A_101_21#_c_143_n N_A_101_21#_c_144_n N_A_101_21#_c_172_p
+ N_A_101_21#_c_145_n N_A_101_21#_c_146_n N_A_101_21#_c_195_p
+ N_A_101_21#_c_198_p N_A_101_21#_c_147_n N_A_101_21#_c_148_n
+ N_A_101_21#_c_149_n N_A_101_21#_c_150_n N_A_101_21#_c_210_p
+ N_A_101_21#_c_199_p N_A_101_21#_c_151_n PM_SKY130_FD_SC_LP__A32O_4%A_101_21#
x_PM_SKY130_FD_SC_LP__A32O_4%A3 N_A3_M1007_g N_A3_M1002_g N_A3_M1026_g
+ N_A3_M1012_g A3 A3 N_A3_c_319_n PM_SKY130_FD_SC_LP__A32O_4%A3
x_PM_SKY130_FD_SC_LP__A32O_4%A2 N_A2_M1001_g N_A2_c_372_n N_A2_M1010_g
+ N_A2_M1008_g N_A2_c_373_n N_A2_M1018_g N_A2_c_369_n N_A2_c_370_n A2 A2
+ PM_SKY130_FD_SC_LP__A32O_4%A2
x_PM_SKY130_FD_SC_LP__A32O_4%A1 N_A1_c_421_n N_A1_M1015_g N_A1_M1006_g
+ N_A1_c_423_n N_A1_M1020_g N_A1_M1023_g A1 A1 N_A1_c_426_n N_A1_c_430_n
+ PM_SKY130_FD_SC_LP__A32O_4%A1
x_PM_SKY130_FD_SC_LP__A32O_4%B1 N_B1_M1024_g N_B1_M1009_g N_B1_M1025_g
+ N_B1_M1027_g B1 N_B1_c_482_n PM_SKY130_FD_SC_LP__A32O_4%B1
x_PM_SKY130_FD_SC_LP__A32O_4%B2 N_B2_M1003_g N_B2_M1005_g N_B2_M1013_g
+ N_B2_M1022_g B2 B2 N_B2_c_540_n PM_SKY130_FD_SC_LP__A32O_4%B2
x_PM_SKY130_FD_SC_LP__A32O_4%VPWR N_VPWR_M1000_d N_VPWR_M1011_d N_VPWR_M1021_d
+ N_VPWR_M1012_d N_VPWR_M1010_s N_VPWR_M1006_s N_VPWR_c_576_n N_VPWR_c_577_n
+ N_VPWR_c_578_n N_VPWR_c_579_n N_VPWR_c_580_n N_VPWR_c_581_n N_VPWR_c_582_n
+ N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n VPWR
+ N_VPWR_c_587_n N_VPWR_c_588_n N_VPWR_c_589_n N_VPWR_c_590_n N_VPWR_c_575_n
+ N_VPWR_c_592_n N_VPWR_c_593_n N_VPWR_c_594_n N_VPWR_c_595_n
+ PM_SKY130_FD_SC_LP__A32O_4%VPWR
x_PM_SKY130_FD_SC_LP__A32O_4%X N_X_M1004_d N_X_M1017_d N_X_M1000_s N_X_M1016_s
+ N_X_c_685_n N_X_c_690_n N_X_c_691_n N_X_c_740_p N_X_c_726_n N_X_c_686_n
+ N_X_c_692_n N_X_c_711_n N_X_c_731_n N_X_c_687_n N_X_c_693_n X X N_X_c_688_n X
+ PM_SKY130_FD_SC_LP__A32O_4%X
x_PM_SKY130_FD_SC_LP__A32O_4%A_511_367# N_A_511_367#_M1002_s
+ N_A_511_367#_M1010_d N_A_511_367#_M1018_d N_A_511_367#_M1023_d
+ N_A_511_367#_M1025_s N_A_511_367#_M1013_d N_A_511_367#_c_764_n
+ N_A_511_367#_c_767_n N_A_511_367#_c_746_n N_A_511_367#_c_747_n
+ N_A_511_367#_c_753_n N_A_511_367#_c_811_n N_A_511_367#_c_755_n
+ N_A_511_367#_c_783_n N_A_511_367#_c_785_n N_A_511_367#_c_756_n
+ N_A_511_367#_c_758_n N_A_511_367#_c_759_n N_A_511_367#_c_748_n
+ N_A_511_367#_c_749_n N_A_511_367#_c_750_n N_A_511_367#_c_762_n
+ N_A_511_367#_c_823_n PM_SKY130_FD_SC_LP__A32O_4%A_511_367#
x_PM_SKY130_FD_SC_LP__A32O_4%VGND N_VGND_M1004_s N_VGND_M1014_s N_VGND_M1019_s
+ N_VGND_M1026_s N_VGND_M1005_d N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n
+ N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n VGND N_VGND_c_832_n
+ N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n
+ N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n
+ PM_SKY130_FD_SC_LP__A32O_4%VGND
x_PM_SKY130_FD_SC_LP__A32O_4%A_511_47# N_A_511_47#_M1007_d N_A_511_47#_M1001_d
+ N_A_511_47#_c_946_n N_A_511_47#_c_939_n N_A_511_47#_c_944_n
+ N_A_511_47#_c_940_n N_A_511_47#_c_941_n N_A_511_47#_c_942_n
+ PM_SKY130_FD_SC_LP__A32O_4%A_511_47#
x_PM_SKY130_FD_SC_LP__A32O_4%A_760_47# N_A_760_47#_M1001_s N_A_760_47#_M1008_s
+ N_A_760_47#_M1020_s N_A_760_47#_c_977_n N_A_760_47#_c_999_n
+ N_A_760_47#_c_982_n N_A_760_47#_c_978_n PM_SKY130_FD_SC_LP__A32O_4%A_760_47#
x_PM_SKY130_FD_SC_LP__A32O_4%A_1208_65# N_A_1208_65#_M1009_s
+ N_A_1208_65#_M1027_s N_A_1208_65#_M1022_s N_A_1208_65#_c_1012_n
+ N_A_1208_65#_c_1013_n N_A_1208_65#_c_1014_n N_A_1208_65#_c_1015_n
+ N_A_1208_65#_c_1016_n N_A_1208_65#_c_1017_n
+ PM_SKY130_FD_SC_LP__A32O_4%A_1208_65#
cc_1 VNB N_A_101_21#_M1004_g 0.0259723f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.655
cc_2 VNB N_A_101_21#_M1000_g 5.27968e-19 $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.465
cc_3 VNB N_A_101_21#_M1014_g 0.0213935f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.655
cc_4 VNB N_A_101_21#_M1011_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=2.465
cc_5 VNB N_A_101_21#_M1017_g 0.0214092f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.655
cc_6 VNB N_A_101_21#_M1016_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.465
cc_7 VNB N_A_101_21#_M1019_g 0.0247122f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.655
cc_8 VNB N_A_101_21#_M1021_g 4.72326e-19 $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=2.465
cc_9 VNB N_A_101_21#_c_141_n 0.00185932f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.485
cc_10 VNB N_A_101_21#_c_142_n 0.0030653f $X=-0.19 $Y=-0.245 $X2=2.11 $Y2=1.385
cc_11 VNB N_A_101_21#_c_143_n 0.00157772f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.16
cc_12 VNB N_A_101_21#_c_144_n 0.00615251f $X=-0.19 $Y=-0.245 $X2=5.065 $Y2=1.18
cc_13 VNB N_A_101_21#_c_145_n 0.0156153f $X=-0.19 $Y=-0.245 $X2=6.255 $Y2=1.09
cc_14 VNB N_A_101_21#_c_146_n 0.00237221f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=1.92
cc_15 VNB N_A_101_21#_c_147_n 0.0406788f $X=-0.19 $Y=-0.245 $X2=4.35 $Y2=1.17
cc_16 VNB N_A_101_21#_c_148_n 0.00359294f $X=-0.19 $Y=-0.245 $X2=4.52 $Y2=1.17
cc_17 VNB N_A_101_21#_c_149_n 6.58869e-19 $X=-0.19 $Y=-0.245 $X2=5.065 $Y2=1.005
cc_18 VNB N_A_101_21#_c_150_n 0.00555694f $X=-0.19 $Y=-0.245 $X2=6.507 $Y2=1.09
cc_19 VNB N_A_101_21#_c_151_n 0.103361f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.48
cc_20 VNB N_A3_M1007_g 0.0251946f $X=-0.19 $Y=-0.245 $X2=6.215 $Y2=1.835
cc_21 VNB N_A3_M1026_g 0.0310724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A3 0.00470788f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.465
cc_23 VNB N_A3_c_319_n 0.0336503f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=2.465
cc_24 VNB N_A2_M1001_g 0.0310686f $X=-0.19 $Y=-0.245 $X2=6.215 $Y2=1.835
cc_25 VNB N_A2_M1008_g 0.0231187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_c_369_n 0.0388304f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.655
cc_27 VNB N_A2_c_370_n 0.0377617f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.465
cc_28 VNB A2 0.00233206f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.315
cc_29 VNB N_A1_c_421_n 0.0154226f $X=-0.19 $Y=-0.245 $X2=5.075 $Y2=0.235
cc_30 VNB N_A1_M1006_g 0.00248417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A1_c_423_n 0.0197633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_M1023_g 0.00219955f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.315
cc_33 VNB A1 0.00218585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A1_c_426_n 0.0758093f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.655
cc_35 VNB N_B1_M1009_g 0.0225971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B1_M1027_g 0.0200387f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.655
cc_37 VNB B1 0.00261634f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.645
cc_38 VNB N_B1_c_482_n 0.048009f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=2.465
cc_39 VNB N_B2_M1005_g 0.0194944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_B2_M1022_g 0.0249241f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.655
cc_41 VNB B2 0.0124118f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.465
cc_42 VNB N_B2_c_540_n 0.03808f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=2.465
cc_43 VNB N_VPWR_c_575_n 0.342803f $X=-0.19 $Y=-0.245 $X2=7.445 $Y2=2.01
cc_44 VNB N_X_c_685_n 0.00264183f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.315
cc_45 VNB N_X_c_686_n 0.00491277f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=2.465
cc_46 VNB N_X_c_687_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=2.465
cc_47 VNB N_X_c_688_n 0.0127231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB X 0.0229484f $X=-0.19 $Y=-0.245 $X2=2.11 $Y2=1.385
cc_49 VNB N_VGND_c_826_n 0.013715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_827_n 0.0276525f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.465
cc_51 VNB N_VGND_c_828_n 3.23981e-19 $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.655
cc_52 VNB N_VGND_c_829_n 0.00505424f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=2.465
cc_53 VNB N_VGND_c_830_n 0.00491137f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.655
cc_54 VNB N_VGND_c_831_n 0.00280617f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.465
cc_55 VNB N_VGND_c_832_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.655
cc_56 VNB N_VGND_c_833_n 0.0160645f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=2.465
cc_57 VNB N_VGND_c_834_n 0.0179543f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.48
cc_58 VNB N_VGND_c_835_n 0.094776f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.16
cc_59 VNB N_VGND_c_836_n 0.0164457f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=1.92
cc_60 VNB N_VGND_c_837_n 0.417458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_838_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=7.28 $Y2=2.01
cc_62 VNB N_VGND_c_839_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_840_n 0.00400911f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.48
cc_64 VNB N_VGND_c_841_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=5.065 $Y2=1.005
cc_65 VNB N_A_511_47#_c_939_n 0.00856246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_511_47#_c_940_n 0.00578081f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.655
cc_67 VNB N_A_511_47#_c_941_n 0.00470309f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.655
cc_68 VNB N_A_511_47#_c_942_n 0.00680243f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.645
cc_69 VNB N_A_760_47#_c_977_n 0.0029187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_760_47#_c_978_n 0.0057213f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.655
cc_71 VNB N_A_1208_65#_c_1012_n 0.00400471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1208_65#_c_1013_n 0.00452996f $X=-0.19 $Y=-0.245 $X2=0.58
+ $Y2=0.655
cc_73 VNB N_A_1208_65#_c_1014_n 0.00362873f $X=-0.19 $Y=-0.245 $X2=0.58
+ $Y2=0.655
cc_74 VNB N_A_1208_65#_c_1015_n 0.0141963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1208_65#_c_1016_n 0.0032521f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.315
cc_76 VNB N_A_1208_65#_c_1017_n 0.0336513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VPB N_A_101_21#_M1000_g 0.0228551f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.465
cc_78 VPB N_A_101_21#_M1011_g 0.018914f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=2.465
cc_79 VPB N_A_101_21#_M1016_g 0.018914f $X=-0.19 $Y=1.655 $X2=1.62 $Y2=2.465
cc_80 VPB N_A_101_21#_M1021_g 0.0201349f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=2.465
cc_81 VPB N_A_101_21#_c_146_n 0.00246378f $X=-0.19 $Y=1.655 $X2=6.345 $Y2=1.92
cc_82 VPB N_A3_M1002_g 0.0187554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A3_M1012_g 0.0231902f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.655
cc_84 VPB A3 0.0060123f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.465
cc_85 VPB N_A3_c_319_n 0.00489857f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=2.465
cc_86 VPB N_A2_c_372_n 0.0212917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A2_c_373_n 0.0162406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A2_c_369_n 0.0217434f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.655
cc_89 VPB N_A2_c_370_n 0.0161134f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.465
cc_90 VPB A2 0.00795006f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=1.315
cc_91 VPB N_A1_M1006_g 0.0203019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A1_M1023_g 0.019961f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.315
cc_93 VPB A1 0.00271665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A1_c_430_n 0.00303762f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=2.465
cc_95 VPB N_B1_M1024_g 0.019461f $X=-0.19 $Y=1.655 $X2=6.215 $Y2=1.835
cc_96 VPB N_B1_M1025_g 0.0209695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB B1 0.00365766f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=1.645
cc_98 VPB N_B1_c_482_n 0.0136721f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=2.465
cc_99 VPB N_B2_M1003_g 0.020497f $X=-0.19 $Y=1.655 $X2=6.215 $Y2=1.835
cc_100 VPB N_B2_M1013_g 0.0244533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB B2 0.0105414f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.465
cc_102 VPB N_B2_c_540_n 0.00530347f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=2.465
cc_103 VPB N_VPWR_c_576_n 0.0415892f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=1.315
cc_104 VPB N_VPWR_c_577_n 3.16049e-19 $X=-0.19 $Y=1.655 $X2=1.19 $Y2=2.465
cc_105 VPB N_VPWR_c_578_n 0.0148832f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=0.655
cc_106 VPB N_VPWR_c_579_n 0.00734048f $X=-0.19 $Y=1.655 $X2=1.62 $Y2=2.465
cc_107 VPB N_VPWR_c_580_n 0.017697f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=1.645
cc_108 VPB N_VPWR_c_581_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=2.025 $Y2=1.485
cc_109 VPB N_VPWR_c_582_n 0.00269298f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_583_n 0.0142356f $X=-0.19 $Y=1.655 $X2=4.35 $Y2=1.16
cc_111 VPB N_VPWR_c_584_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=1.16
cc_112 VPB N_VPWR_c_585_n 0.0129398f $X=-0.19 $Y=1.655 $X2=5.065 $Y2=1.18
cc_113 VPB N_VPWR_c_586_n 0.00436868f $X=-0.19 $Y=1.655 $X2=4.52 $Y2=1.18
cc_114 VPB N_VPWR_c_587_n 0.0152106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_588_n 0.0310212f $X=-0.19 $Y=1.655 $X2=7.28 $Y2=2.01
cc_116 VPB N_VPWR_c_589_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.48
cc_117 VPB N_VPWR_c_590_n 0.061589f $X=-0.19 $Y=1.655 $X2=6.37 $Y2=2.095
cc_118 VPB N_VPWR_c_575_n 0.0830038f $X=-0.19 $Y=1.655 $X2=7.445 $Y2=2.01
cc_119 VPB N_VPWR_c_592_n 0.00439477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_593_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=1.48
cc_121 VPB N_VPWR_c_594_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.62 $Y2=1.48
cc_122 VPB N_VPWR_c_595_n 0.00510472f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=1.48
cc_123 VPB N_X_c_690_n 0.00632202f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.655
cc_124 VPB N_X_c_691_n 0.0178875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_X_c_692_n 0.00586684f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=1.315
cc_126 VPB N_X_c_693_n 0.00144499f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=2.465
cc_127 VPB X 0.00550956f $X=-0.19 $Y=1.655 $X2=2.11 $Y2=1.385
cc_128 VPB N_A_511_367#_c_746_n 0.0300084f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=0.655
cc_129 VPB N_A_511_367#_c_747_n 0.0260196f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=2.465
cc_130 VPB N_A_511_367#_c_748_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.48
cc_131 VPB N_A_511_367#_c_749_n 0.0376742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_511_367#_c_750_n 0.00193743f $X=-0.19 $Y=1.655 $X2=5.065 $Y2=1.18
cc_133 N_A_101_21#_M1019_g N_A3_M1007_g 0.0239473f $X=1.87 $Y=0.655 $X2=0 $Y2=0
cc_134 N_A_101_21#_c_142_n N_A3_M1007_g 0.00197849f $X=2.11 $Y=1.385 $X2=0 $Y2=0
cc_135 N_A_101_21#_c_147_n N_A3_M1007_g 0.0189633f $X=4.35 $Y=1.17 $X2=0 $Y2=0
cc_136 N_A_101_21#_c_151_n N_A3_M1007_g 0.0228008f $X=2.05 $Y=1.48 $X2=0 $Y2=0
cc_137 N_A_101_21#_c_147_n N_A3_M1026_g 0.0125934f $X=4.35 $Y=1.17 $X2=0 $Y2=0
cc_138 N_A_101_21#_M1021_g A3 4.88703e-19 $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_101_21#_c_142_n A3 0.00761478f $X=2.11 $Y=1.385 $X2=0 $Y2=0
cc_140 N_A_101_21#_c_147_n A3 0.0511531f $X=4.35 $Y=1.17 $X2=0 $Y2=0
cc_141 N_A_101_21#_c_151_n A3 5.02134e-19 $X=2.05 $Y=1.48 $X2=0 $Y2=0
cc_142 N_A_101_21#_M1021_g N_A3_c_319_n 0.0217956f $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_101_21#_c_142_n N_A3_c_319_n 9.75998e-19 $X=2.11 $Y=1.385 $X2=0 $Y2=0
cc_144 N_A_101_21#_c_147_n N_A3_c_319_n 0.00244902f $X=4.35 $Y=1.17 $X2=0 $Y2=0
cc_145 N_A_101_21#_c_147_n N_A2_M1001_g 0.0127155f $X=4.35 $Y=1.17 $X2=0 $Y2=0
cc_146 N_A_101_21#_c_148_n N_A2_M1001_g 5.45556e-19 $X=4.52 $Y=1.17 $X2=0 $Y2=0
cc_147 N_A_101_21#_c_144_n N_A2_M1008_g 0.00886608f $X=5.065 $Y=1.18 $X2=0 $Y2=0
cc_148 N_A_101_21#_c_172_p N_A2_M1008_g 3.2364e-19 $X=5.215 $Y=0.78 $X2=0 $Y2=0
cc_149 N_A_101_21#_c_148_n N_A2_M1008_g 0.00396532f $X=4.52 $Y=1.17 $X2=0 $Y2=0
cc_150 N_A_101_21#_c_149_n N_A2_M1008_g 3.88092e-19 $X=5.065 $Y=1.005 $X2=0
+ $Y2=0
cc_151 N_A_101_21#_c_147_n N_A2_c_369_n 0.0141409f $X=4.35 $Y=1.17 $X2=0 $Y2=0
cc_152 N_A_101_21#_c_144_n N_A2_c_370_n 0.00577855f $X=5.065 $Y=1.18 $X2=0 $Y2=0
cc_153 N_A_101_21#_c_147_n N_A2_c_370_n 0.00153185f $X=4.35 $Y=1.17 $X2=0 $Y2=0
cc_154 N_A_101_21#_c_148_n N_A2_c_370_n 0.00193272f $X=4.52 $Y=1.17 $X2=0 $Y2=0
cc_155 N_A_101_21#_c_147_n A2 0.0560529f $X=4.35 $Y=1.17 $X2=0 $Y2=0
cc_156 N_A_101_21#_c_144_n N_A1_c_421_n 0.00613167f $X=5.065 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A_101_21#_c_172_p N_A1_c_421_n 0.00449407f $X=5.215 $Y=0.78 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A_101_21#_c_149_n N_A1_c_421_n 0.00383944f $X=5.065 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A_101_21#_c_145_n N_A1_c_423_n 0.0143692f $X=6.255 $Y=1.09 $X2=0 $Y2=0
cc_160 N_A_101_21#_c_149_n N_A1_c_423_n 2.95668e-19 $X=5.065 $Y=1.005 $X2=0
+ $Y2=0
cc_161 N_A_101_21#_c_145_n A1 0.0347355f $X=6.255 $Y=1.09 $X2=0 $Y2=0
cc_162 N_A_101_21#_c_146_n A1 0.0302761f $X=6.345 $Y=1.92 $X2=0 $Y2=0
cc_163 N_A_101_21#_c_144_n N_A1_c_426_n 0.00454866f $X=5.065 $Y=1.18 $X2=0 $Y2=0
cc_164 N_A_101_21#_c_145_n N_A1_c_426_n 0.0102634f $X=6.255 $Y=1.09 $X2=0 $Y2=0
cc_165 N_A_101_21#_c_146_n N_A1_c_426_n 0.00333612f $X=6.345 $Y=1.92 $X2=0 $Y2=0
cc_166 N_A_101_21#_c_149_n N_A1_c_426_n 0.0114096f $X=5.065 $Y=1.005 $X2=0 $Y2=0
cc_167 N_A_101_21#_c_145_n N_A1_c_430_n 0.0201356f $X=6.255 $Y=1.09 $X2=0 $Y2=0
cc_168 N_A_101_21#_c_149_n N_A1_c_430_n 0.00930273f $X=5.065 $Y=1.005 $X2=0
+ $Y2=0
cc_169 N_A_101_21#_c_146_n N_B1_M1024_g 0.00314347f $X=6.345 $Y=1.92 $X2=0 $Y2=0
cc_170 N_A_101_21#_c_146_n N_B1_M1009_g 0.00502218f $X=6.345 $Y=1.92 $X2=0 $Y2=0
cc_171 N_A_101_21#_c_195_p N_B1_M1009_g 0.0101505f $X=6.595 $Y=0.685 $X2=0 $Y2=0
cc_172 N_A_101_21#_c_150_n N_B1_M1009_g 0.0111181f $X=6.507 $Y=1.09 $X2=0 $Y2=0
cc_173 N_A_101_21#_c_146_n N_B1_M1025_g 0.00323609f $X=6.345 $Y=1.92 $X2=0 $Y2=0
cc_174 N_A_101_21#_c_198_p N_B1_M1025_g 0.0174774f $X=7.28 $Y=2.01 $X2=0 $Y2=0
cc_175 N_A_101_21#_c_199_p N_B1_M1025_g 8.62433e-19 $X=7.445 $Y=2.035 $X2=0
+ $Y2=0
cc_176 N_A_101_21#_c_146_n N_B1_M1027_g 6.71898e-19 $X=6.345 $Y=1.92 $X2=0 $Y2=0
cc_177 N_A_101_21#_c_195_p N_B1_M1027_g 0.00445893f $X=6.595 $Y=0.685 $X2=0
+ $Y2=0
cc_178 N_A_101_21#_c_150_n N_B1_M1027_g 0.00224898f $X=6.507 $Y=1.09 $X2=0 $Y2=0
cc_179 N_A_101_21#_c_146_n B1 0.0229569f $X=6.345 $Y=1.92 $X2=0 $Y2=0
cc_180 N_A_101_21#_c_198_p B1 0.0308046f $X=7.28 $Y=2.01 $X2=0 $Y2=0
cc_181 N_A_101_21#_c_150_n B1 0.00892757f $X=6.507 $Y=1.09 $X2=0 $Y2=0
cc_182 N_A_101_21#_c_145_n N_B1_c_482_n 0.0075683f $X=6.255 $Y=1.09 $X2=0 $Y2=0
cc_183 N_A_101_21#_c_146_n N_B1_c_482_n 0.020985f $X=6.345 $Y=1.92 $X2=0 $Y2=0
cc_184 N_A_101_21#_c_198_p N_B1_c_482_n 0.00115635f $X=7.28 $Y=2.01 $X2=0 $Y2=0
cc_185 N_A_101_21#_c_150_n N_B1_c_482_n 0.00415513f $X=6.507 $Y=1.09 $X2=0 $Y2=0
cc_186 N_A_101_21#_c_210_p N_B1_c_482_n 0.00223208f $X=6.37 $Y=2.095 $X2=0 $Y2=0
cc_187 N_A_101_21#_c_198_p N_B2_M1003_g 0.0140177f $X=7.28 $Y=2.01 $X2=0 $Y2=0
cc_188 N_A_101_21#_c_199_p N_B2_M1003_g 0.012268f $X=7.445 $Y=2.035 $X2=0 $Y2=0
cc_189 N_A_101_21#_c_199_p N_B2_M1013_g 0.011823f $X=7.445 $Y=2.035 $X2=0 $Y2=0
cc_190 N_A_101_21#_c_199_p B2 0.0189955f $X=7.445 $Y=2.035 $X2=0 $Y2=0
cc_191 N_A_101_21#_c_199_p N_B2_c_540_n 6.52238e-19 $X=7.445 $Y=2.035 $X2=0
+ $Y2=0
cc_192 N_A_101_21#_M1000_g N_VPWR_c_576_n 0.0154852f $X=0.76 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_A_101_21#_M1011_g N_VPWR_c_576_n 7.27171e-19 $X=1.19 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_A_101_21#_M1000_g N_VPWR_c_577_n 7.27171e-19 $X=0.76 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_101_21#_M1011_g N_VPWR_c_577_n 0.0143393f $X=1.19 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A_101_21#_M1016_g N_VPWR_c_577_n 0.0144311f $X=1.62 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_A_101_21#_M1021_g N_VPWR_c_577_n 7.43396e-19 $X=2.05 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A_101_21#_M1016_g N_VPWR_c_578_n 0.00486043f $X=1.62 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A_101_21#_M1021_g N_VPWR_c_578_n 0.00585385f $X=2.05 $Y=2.465 $X2=0
+ $Y2=0
cc_200 N_A_101_21#_M1021_g N_VPWR_c_579_n 0.00257804f $X=2.05 $Y=2.465 $X2=0
+ $Y2=0
cc_201 N_A_101_21#_c_142_n N_VPWR_c_579_n 0.0037238f $X=2.11 $Y=1.385 $X2=0
+ $Y2=0
cc_202 N_A_101_21#_c_147_n N_VPWR_c_579_n 0.00631199f $X=4.35 $Y=1.17 $X2=0
+ $Y2=0
cc_203 N_A_101_21#_c_151_n N_VPWR_c_579_n 0.00130979f $X=2.05 $Y=1.48 $X2=0
+ $Y2=0
cc_204 N_A_101_21#_M1000_g N_VPWR_c_585_n 0.00486043f $X=0.76 $Y=2.465 $X2=0
+ $Y2=0
cc_205 N_A_101_21#_M1011_g N_VPWR_c_585_n 0.00486043f $X=1.19 $Y=2.465 $X2=0
+ $Y2=0
cc_206 N_A_101_21#_M1024_d N_VPWR_c_575_n 0.00289524f $X=6.215 $Y=1.835 $X2=0
+ $Y2=0
cc_207 N_A_101_21#_M1003_s N_VPWR_c_575_n 0.00225186f $X=7.305 $Y=1.835 $X2=0
+ $Y2=0
cc_208 N_A_101_21#_M1000_g N_VPWR_c_575_n 0.00824727f $X=0.76 $Y=2.465 $X2=0
+ $Y2=0
cc_209 N_A_101_21#_M1011_g N_VPWR_c_575_n 0.00824727f $X=1.19 $Y=2.465 $X2=0
+ $Y2=0
cc_210 N_A_101_21#_M1016_g N_VPWR_c_575_n 0.00824727f $X=1.62 $Y=2.465 $X2=0
+ $Y2=0
cc_211 N_A_101_21#_M1021_g N_VPWR_c_575_n 0.0105614f $X=2.05 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_A_101_21#_M1004_g N_X_c_685_n 0.0155484f $X=0.58 $Y=0.655 $X2=0 $Y2=0
cc_213 N_A_101_21#_c_141_n N_X_c_685_n 0.013516f $X=2.025 $Y=1.485 $X2=0 $Y2=0
cc_214 N_A_101_21#_M1000_g N_X_c_690_n 0.0150987f $X=0.76 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A_101_21#_c_141_n N_X_c_690_n 0.0265438f $X=2.025 $Y=1.485 $X2=0 $Y2=0
cc_216 N_A_101_21#_c_151_n N_X_c_690_n 0.00508873f $X=2.05 $Y=1.48 $X2=0 $Y2=0
cc_217 N_A_101_21#_M1014_g N_X_c_686_n 0.0139345f $X=1.01 $Y=0.655 $X2=0 $Y2=0
cc_218 N_A_101_21#_M1017_g N_X_c_686_n 0.0143278f $X=1.44 $Y=0.655 $X2=0 $Y2=0
cc_219 N_A_101_21#_M1019_g N_X_c_686_n 0.00465294f $X=1.87 $Y=0.655 $X2=0 $Y2=0
cc_220 N_A_101_21#_c_141_n N_X_c_686_n 0.0683925f $X=2.025 $Y=1.485 $X2=0 $Y2=0
cc_221 N_A_101_21#_c_143_n N_X_c_686_n 0.01083f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_101_21#_c_151_n N_X_c_686_n 0.00582235f $X=2.05 $Y=1.48 $X2=0 $Y2=0
cc_223 N_A_101_21#_M1011_g N_X_c_692_n 0.0131657f $X=1.19 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_101_21#_M1016_g N_X_c_692_n 0.0130597f $X=1.62 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A_101_21#_M1021_g N_X_c_692_n 0.00219544f $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A_101_21#_c_141_n N_X_c_692_n 0.0660589f $X=2.025 $Y=1.485 $X2=0 $Y2=0
cc_227 N_A_101_21#_c_151_n N_X_c_692_n 0.00575333f $X=2.05 $Y=1.48 $X2=0 $Y2=0
cc_228 N_A_101_21#_M1019_g N_X_c_711_n 0.010639f $X=1.87 $Y=0.655 $X2=0 $Y2=0
cc_229 N_A_101_21#_c_141_n N_X_c_687_n 0.0154947f $X=2.025 $Y=1.485 $X2=0 $Y2=0
cc_230 N_A_101_21#_c_151_n N_X_c_687_n 0.00296179f $X=2.05 $Y=1.48 $X2=0 $Y2=0
cc_231 N_A_101_21#_c_141_n N_X_c_693_n 0.0154948f $X=2.025 $Y=1.485 $X2=0 $Y2=0
cc_232 N_A_101_21#_c_151_n N_X_c_693_n 0.00292626f $X=2.05 $Y=1.48 $X2=0 $Y2=0
cc_233 N_A_101_21#_M1004_g X 0.00656472f $X=0.58 $Y=0.655 $X2=0 $Y2=0
cc_234 N_A_101_21#_M1000_g X 0.00320248f $X=0.76 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A_101_21#_c_141_n X 0.0162005f $X=2.025 $Y=1.485 $X2=0 $Y2=0
cc_236 N_A_101_21#_c_151_n X 0.00402444f $X=2.05 $Y=1.48 $X2=0 $Y2=0
cc_237 N_A_101_21#_c_198_p N_A_511_367#_M1025_s 0.0076516f $X=7.28 $Y=2.01 $X2=0
+ $Y2=0
cc_238 N_A_101_21#_c_147_n N_A_511_367#_c_746_n 0.00602555f $X=4.35 $Y=1.17
+ $X2=0 $Y2=0
cc_239 N_A_101_21#_c_147_n N_A_511_367#_c_753_n 0.00223718f $X=4.35 $Y=1.17
+ $X2=0 $Y2=0
cc_240 N_A_101_21#_c_148_n N_A_511_367#_c_753_n 0.0124106f $X=4.52 $Y=1.17 $X2=0
+ $Y2=0
cc_241 N_A_101_21#_c_149_n N_A_511_367#_c_755_n 0.00145776f $X=5.065 $Y=1.005
+ $X2=0 $Y2=0
cc_242 N_A_101_21#_M1024_d N_A_511_367#_c_756_n 0.0049251f $X=6.215 $Y=1.835
+ $X2=0 $Y2=0
cc_243 N_A_101_21#_c_210_p N_A_511_367#_c_756_n 0.0187238f $X=6.37 $Y=2.095
+ $X2=0 $Y2=0
cc_244 N_A_101_21#_c_198_p N_A_511_367#_c_758_n 0.0258086f $X=7.28 $Y=2.01 $X2=0
+ $Y2=0
cc_245 N_A_101_21#_M1003_s N_A_511_367#_c_759_n 0.00332344f $X=7.305 $Y=1.835
+ $X2=0 $Y2=0
cc_246 N_A_101_21#_c_199_p N_A_511_367#_c_759_n 0.0159805f $X=7.445 $Y=2.035
+ $X2=0 $Y2=0
cc_247 N_A_101_21#_c_147_n N_A_511_367#_c_750_n 8.27402e-19 $X=4.35 $Y=1.17
+ $X2=0 $Y2=0
cc_248 N_A_101_21#_c_144_n N_A_511_367#_c_762_n 0.00407135f $X=5.065 $Y=1.18
+ $X2=0 $Y2=0
cc_249 N_A_101_21#_c_149_n N_A_511_367#_c_762_n 8.48097e-19 $X=5.065 $Y=1.005
+ $X2=0 $Y2=0
cc_250 N_A_101_21#_c_143_n N_VGND_M1019_s 0.00186483f $X=2.195 $Y=1.16 $X2=0
+ $Y2=0
cc_251 N_A_101_21#_M1004_g N_VGND_c_827_n 0.0118475f $X=0.58 $Y=0.655 $X2=0
+ $Y2=0
cc_252 N_A_101_21#_M1014_g N_VGND_c_827_n 6.25324e-19 $X=1.01 $Y=0.655 $X2=0
+ $Y2=0
cc_253 N_A_101_21#_M1004_g N_VGND_c_828_n 6.25324e-19 $X=0.58 $Y=0.655 $X2=0
+ $Y2=0
cc_254 N_A_101_21#_M1014_g N_VGND_c_828_n 0.0109423f $X=1.01 $Y=0.655 $X2=0
+ $Y2=0
cc_255 N_A_101_21#_M1017_g N_VGND_c_828_n 0.0111435f $X=1.44 $Y=0.655 $X2=0
+ $Y2=0
cc_256 N_A_101_21#_M1019_g N_VGND_c_828_n 4.85852e-19 $X=1.87 $Y=0.655 $X2=0
+ $Y2=0
cc_257 N_A_101_21#_M1019_g N_VGND_c_829_n 0.00832443f $X=1.87 $Y=0.655 $X2=0
+ $Y2=0
cc_258 N_A_101_21#_c_141_n N_VGND_c_829_n 4.85238e-19 $X=2.025 $Y=1.485 $X2=0
+ $Y2=0
cc_259 N_A_101_21#_c_143_n N_VGND_c_829_n 0.0150074f $X=2.195 $Y=1.16 $X2=0
+ $Y2=0
cc_260 N_A_101_21#_c_147_n N_VGND_c_829_n 0.0118695f $X=4.35 $Y=1.17 $X2=0 $Y2=0
cc_261 N_A_101_21#_c_151_n N_VGND_c_829_n 0.00112419f $X=2.05 $Y=1.48 $X2=0
+ $Y2=0
cc_262 N_A_101_21#_M1004_g N_VGND_c_832_n 0.00486043f $X=0.58 $Y=0.655 $X2=0
+ $Y2=0
cc_263 N_A_101_21#_M1014_g N_VGND_c_832_n 0.00486043f $X=1.01 $Y=0.655 $X2=0
+ $Y2=0
cc_264 N_A_101_21#_M1017_g N_VGND_c_833_n 0.00486043f $X=1.44 $Y=0.655 $X2=0
+ $Y2=0
cc_265 N_A_101_21#_M1019_g N_VGND_c_833_n 0.0054895f $X=1.87 $Y=0.655 $X2=0
+ $Y2=0
cc_266 N_A_101_21#_M1015_d N_VGND_c_837_n 0.00225186f $X=5.075 $Y=0.235 $X2=0
+ $Y2=0
cc_267 N_A_101_21#_M1004_g N_VGND_c_837_n 0.00824727f $X=0.58 $Y=0.655 $X2=0
+ $Y2=0
cc_268 N_A_101_21#_M1014_g N_VGND_c_837_n 0.00824727f $X=1.01 $Y=0.655 $X2=0
+ $Y2=0
cc_269 N_A_101_21#_M1017_g N_VGND_c_837_n 0.00824727f $X=1.44 $Y=0.655 $X2=0
+ $Y2=0
cc_270 N_A_101_21#_M1019_g N_VGND_c_837_n 0.0103565f $X=1.87 $Y=0.655 $X2=0
+ $Y2=0
cc_271 N_A_101_21#_c_147_n N_A_511_47#_c_939_n 0.0522849f $X=4.35 $Y=1.17 $X2=0
+ $Y2=0
cc_272 N_A_101_21#_c_147_n N_A_511_47#_c_944_n 0.0216981f $X=4.35 $Y=1.17 $X2=0
+ $Y2=0
cc_273 N_A_101_21#_c_147_n N_A_511_47#_c_942_n 0.0061084f $X=4.35 $Y=1.17 $X2=0
+ $Y2=0
cc_274 N_A_101_21#_c_145_n N_A_760_47#_M1020_s 0.00253571f $X=6.255 $Y=1.09
+ $X2=0 $Y2=0
cc_275 N_A_101_21#_c_144_n N_A_760_47#_c_977_n 0.0241977f $X=5.065 $Y=1.18 $X2=0
+ $Y2=0
cc_276 N_A_101_21#_c_147_n N_A_760_47#_c_977_n 0.0476369f $X=4.35 $Y=1.17 $X2=0
+ $Y2=0
cc_277 N_A_101_21#_M1015_d N_A_760_47#_c_982_n 0.00333487f $X=5.075 $Y=0.235
+ $X2=0 $Y2=0
cc_278 N_A_101_21#_c_144_n N_A_760_47#_c_982_n 0.00355104f $X=5.065 $Y=1.18
+ $X2=0 $Y2=0
cc_279 N_A_101_21#_c_172_p N_A_760_47#_c_982_n 0.0133188f $X=5.215 $Y=0.78 $X2=0
+ $Y2=0
cc_280 N_A_101_21#_c_145_n N_A_760_47#_c_982_n 0.00319377f $X=6.255 $Y=1.09
+ $X2=0 $Y2=0
cc_281 N_A_101_21#_c_145_n N_A_760_47#_c_978_n 0.0217186f $X=6.255 $Y=1.09 $X2=0
+ $Y2=0
cc_282 N_A_101_21#_c_145_n N_A_1208_65#_M1009_s 0.00295914f $X=6.255 $Y=1.09
+ $X2=-0.19 $Y2=-0.245
cc_283 N_A_101_21#_c_145_n N_A_1208_65#_c_1012_n 0.0199559f $X=6.255 $Y=1.09
+ $X2=0 $Y2=0
cc_284 N_A_101_21#_M1009_d N_A_1208_65#_c_1013_n 0.00176461f $X=6.455 $Y=0.325
+ $X2=0 $Y2=0
cc_285 N_A_101_21#_c_195_p N_A_1208_65#_c_1013_n 0.0157897f $X=6.595 $Y=0.685
+ $X2=0 $Y2=0
cc_286 N_A_101_21#_c_150_n N_A_1208_65#_c_1013_n 0.00345027f $X=6.507 $Y=1.09
+ $X2=0 $Y2=0
cc_287 N_A_101_21#_c_198_p N_A_1208_65#_c_1015_n 0.00319778f $X=7.28 $Y=2.01
+ $X2=0 $Y2=0
cc_288 N_A_101_21#_c_199_p N_A_1208_65#_c_1015_n 0.00126792f $X=7.445 $Y=2.035
+ $X2=0 $Y2=0
cc_289 N_A_101_21#_c_146_n N_A_1208_65#_c_1016_n 7.26297e-19 $X=6.345 $Y=1.92
+ $X2=0 $Y2=0
cc_290 N_A_101_21#_c_198_p N_A_1208_65#_c_1016_n 0.00201842f $X=7.28 $Y=2.01
+ $X2=0 $Y2=0
cc_291 N_A_101_21#_c_150_n N_A_1208_65#_c_1016_n 0.00465389f $X=6.507 $Y=1.09
+ $X2=0 $Y2=0
cc_292 A3 N_A2_c_369_n 0.00127794f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_293 N_A3_c_319_n N_A2_c_369_n 0.00829695f $X=2.91 $Y=1.51 $X2=0 $Y2=0
cc_294 A3 A2 0.0261203f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_295 N_A3_c_319_n A2 0.00115592f $X=2.91 $Y=1.51 $X2=0 $Y2=0
cc_296 N_A3_M1002_g N_VPWR_c_579_n 0.00283131f $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A3_M1002_g N_VPWR_c_580_n 7.25108e-19 $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A3_M1012_g N_VPWR_c_580_n 0.0175037f $X=2.91 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A3_M1002_g N_VPWR_c_587_n 0.00564131f $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A3_M1012_g N_VPWR_c_587_n 0.00486043f $X=2.91 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A3_M1002_g N_VPWR_c_575_n 0.0101343f $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A3_M1012_g N_VPWR_c_575_n 0.00824727f $X=2.91 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A3_M1007_g N_X_c_686_n 2.28684e-19 $X=2.48 $Y=0.655 $X2=0 $Y2=0
cc_304 N_A3_M1007_g N_X_c_711_n 7.56538e-19 $X=2.48 $Y=0.655 $X2=0 $Y2=0
cc_305 N_A3_M1002_g N_A_511_367#_c_764_n 0.00181166f $X=2.48 $Y=2.465 $X2=0
+ $Y2=0
cc_306 A3 N_A_511_367#_c_764_n 0.0184067f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_307 N_A3_c_319_n N_A_511_367#_c_764_n 6.52992e-19 $X=2.91 $Y=1.51 $X2=0 $Y2=0
cc_308 N_A3_M1002_g N_A_511_367#_c_767_n 0.00979812f $X=2.48 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A3_M1012_g N_A_511_367#_c_746_n 0.0143f $X=2.91 $Y=2.465 $X2=0 $Y2=0
cc_310 A3 N_A_511_367#_c_746_n 0.0307065f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_311 N_A3_M1007_g N_VGND_c_829_n 0.00989967f $X=2.48 $Y=0.655 $X2=0 $Y2=0
cc_312 N_A3_M1026_g N_VGND_c_830_n 0.00452846f $X=2.91 $Y=0.655 $X2=0 $Y2=0
cc_313 N_A3_M1007_g N_VGND_c_834_n 0.0054895f $X=2.48 $Y=0.655 $X2=0 $Y2=0
cc_314 N_A3_M1026_g N_VGND_c_834_n 0.00427134f $X=2.91 $Y=0.655 $X2=0 $Y2=0
cc_315 N_A3_M1007_g N_VGND_c_837_n 0.0103565f $X=2.48 $Y=0.655 $X2=0 $Y2=0
cc_316 N_A3_M1026_g N_VGND_c_837_n 0.00712579f $X=2.91 $Y=0.655 $X2=0 $Y2=0
cc_317 N_A3_M1007_g N_A_511_47#_c_946_n 0.00587296f $X=2.48 $Y=0.655 $X2=0 $Y2=0
cc_318 N_A3_M1026_g N_A_511_47#_c_946_n 0.00734598f $X=2.91 $Y=0.655 $X2=0 $Y2=0
cc_319 N_A3_M1026_g N_A_511_47#_c_939_n 0.0107346f $X=2.91 $Y=0.655 $X2=0 $Y2=0
cc_320 N_A3_M1007_g N_A_511_47#_c_944_n 0.00218378f $X=2.48 $Y=0.655 $X2=0 $Y2=0
cc_321 N_A3_M1026_g N_A_511_47#_c_944_n 7.1695e-19 $X=2.91 $Y=0.655 $X2=0 $Y2=0
cc_322 N_A3_M1026_g N_A_511_47#_c_940_n 0.00253083f $X=2.91 $Y=0.655 $X2=0 $Y2=0
cc_323 N_A2_M1008_g N_A1_c_421_n 0.0245583f $X=4.57 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_324 N_A2_c_373_n N_A1_M1006_g 0.0119913f $X=4.79 $Y=1.725 $X2=0 $Y2=0
cc_325 N_A2_M1008_g N_A1_c_426_n 0.00808178f $X=4.57 $Y=0.655 $X2=0 $Y2=0
cc_326 N_A2_c_370_n N_A1_c_426_n 0.0119913f $X=4.57 $Y=1.535 $X2=0 $Y2=0
cc_327 N_A2_c_370_n N_A1_c_430_n 0.00204487f $X=4.57 $Y=1.535 $X2=0 $Y2=0
cc_328 N_A2_c_372_n N_VPWR_c_581_n 0.0166685f $X=4.36 $Y=1.725 $X2=0 $Y2=0
cc_329 N_A2_c_373_n N_VPWR_c_581_n 0.0147787f $X=4.79 $Y=1.725 $X2=0 $Y2=0
cc_330 N_A2_c_373_n N_VPWR_c_582_n 6.80491e-19 $X=4.79 $Y=1.725 $X2=0 $Y2=0
cc_331 N_A2_c_372_n N_VPWR_c_588_n 0.00486043f $X=4.36 $Y=1.725 $X2=0 $Y2=0
cc_332 N_A2_c_373_n N_VPWR_c_589_n 0.00486043f $X=4.79 $Y=1.725 $X2=0 $Y2=0
cc_333 N_A2_c_372_n N_VPWR_c_575_n 0.00954696f $X=4.36 $Y=1.725 $X2=0 $Y2=0
cc_334 N_A2_c_373_n N_VPWR_c_575_n 0.0082726f $X=4.79 $Y=1.725 $X2=0 $Y2=0
cc_335 N_A2_c_369_n N_A_511_367#_c_746_n 0.00239183f $X=4.065 $Y=1.535 $X2=0
+ $Y2=0
cc_336 A2 N_A_511_367#_c_746_n 0.0325033f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_337 N_A2_c_372_n N_A_511_367#_c_753_n 0.0142681f $X=4.36 $Y=1.725 $X2=0 $Y2=0
cc_338 N_A2_c_373_n N_A_511_367#_c_753_n 0.0137805f $X=4.79 $Y=1.725 $X2=0 $Y2=0
cc_339 N_A2_c_370_n N_A_511_367#_c_753_n 0.00302099f $X=4.57 $Y=1.535 $X2=0
+ $Y2=0
cc_340 N_A2_c_369_n N_A_511_367#_c_750_n 0.00249628f $X=4.065 $Y=1.535 $X2=0
+ $Y2=0
cc_341 N_A2_c_370_n N_A_511_367#_c_750_n 0.00104367f $X=4.57 $Y=1.535 $X2=0
+ $Y2=0
cc_342 A2 N_A_511_367#_c_750_n 0.0297788f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_343 N_A2_M1001_g N_VGND_c_835_n 0.00357877f $X=4.14 $Y=0.655 $X2=0 $Y2=0
cc_344 N_A2_M1008_g N_VGND_c_835_n 0.00419907f $X=4.57 $Y=0.655 $X2=0 $Y2=0
cc_345 N_A2_M1001_g N_VGND_c_837_n 0.00675087f $X=4.14 $Y=0.655 $X2=0 $Y2=0
cc_346 N_A2_M1008_g N_VGND_c_837_n 0.00590502f $X=4.57 $Y=0.655 $X2=0 $Y2=0
cc_347 N_A2_M1001_g N_A_511_47#_c_940_n 0.00308861f $X=4.14 $Y=0.655 $X2=0 $Y2=0
cc_348 N_A2_M1001_g N_A_511_47#_c_942_n 0.013065f $X=4.14 $Y=0.655 $X2=0 $Y2=0
cc_349 N_A2_M1008_g N_A_511_47#_c_942_n 0.00314793f $X=4.57 $Y=0.655 $X2=0 $Y2=0
cc_350 N_A2_M1001_g N_A_760_47#_c_977_n 0.00950592f $X=4.14 $Y=0.655 $X2=0 $Y2=0
cc_351 N_A2_M1008_g N_A_760_47#_c_977_n 0.0109752f $X=4.57 $Y=0.655 $X2=0 $Y2=0
cc_352 A1 N_B1_M1024_g 0.00186697f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_353 N_A1_c_426_n N_B1_M1009_g 0.00368882f $X=5.67 $Y=1.44 $X2=0 $Y2=0
cc_354 N_A1_M1023_g N_B1_c_482_n 0.0215482f $X=5.71 $Y=2.465 $X2=0 $Y2=0
cc_355 A1 N_B1_c_482_n 0.00866412f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_356 N_A1_c_426_n N_B1_c_482_n 0.0153333f $X=5.67 $Y=1.44 $X2=0 $Y2=0
cc_357 N_A1_M1006_g N_VPWR_c_581_n 6.80491e-19 $X=5.22 $Y=2.465 $X2=0 $Y2=0
cc_358 N_A1_M1006_g N_VPWR_c_582_n 0.0147329f $X=5.22 $Y=2.465 $X2=0 $Y2=0
cc_359 N_A1_M1023_g N_VPWR_c_582_n 0.00744408f $X=5.71 $Y=2.465 $X2=0 $Y2=0
cc_360 N_A1_M1006_g N_VPWR_c_589_n 0.00486043f $X=5.22 $Y=2.465 $X2=0 $Y2=0
cc_361 N_A1_M1023_g N_VPWR_c_590_n 0.00562613f $X=5.71 $Y=2.465 $X2=0 $Y2=0
cc_362 N_A1_M1006_g N_VPWR_c_575_n 0.0082726f $X=5.22 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A1_M1023_g N_VPWR_c_575_n 0.010364f $X=5.71 $Y=2.465 $X2=0 $Y2=0
cc_364 N_A1_M1006_g N_A_511_367#_c_755_n 0.0131008f $X=5.22 $Y=2.465 $X2=0 $Y2=0
cc_365 N_A1_M1023_g N_A_511_367#_c_755_n 0.0122289f $X=5.71 $Y=2.465 $X2=0 $Y2=0
cc_366 A1 N_A_511_367#_c_755_n 0.0102615f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_367 N_A1_c_426_n N_A_511_367#_c_755_n 7.80219e-19 $X=5.67 $Y=1.44 $X2=0 $Y2=0
cc_368 N_A1_c_430_n N_A_511_367#_c_755_n 0.0303405f $X=5.622 $Y=1.552 $X2=0
+ $Y2=0
cc_369 N_A1_M1023_g N_A_511_367#_c_783_n 4.27055e-19 $X=5.71 $Y=2.465 $X2=0
+ $Y2=0
cc_370 A1 N_A_511_367#_c_783_n 0.0222259f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A1_M1006_g N_A_511_367#_c_785_n 5.7599e-19 $X=5.22 $Y=2.465 $X2=0 $Y2=0
cc_372 N_A1_M1023_g N_A_511_367#_c_785_n 0.0116541f $X=5.71 $Y=2.465 $X2=0 $Y2=0
cc_373 N_A1_c_426_n N_A_511_367#_c_762_n 0.00353709f $X=5.67 $Y=1.44 $X2=0 $Y2=0
cc_374 N_A1_c_421_n N_VGND_c_835_n 0.00357877f $X=5 $Y=1.185 $X2=0 $Y2=0
cc_375 N_A1_c_423_n N_VGND_c_835_n 0.00357842f $X=5.43 $Y=1.185 $X2=0 $Y2=0
cc_376 N_A1_c_421_n N_VGND_c_837_n 0.00537654f $X=5 $Y=1.185 $X2=0 $Y2=0
cc_377 N_A1_c_423_n N_VGND_c_837_n 0.00665087f $X=5.43 $Y=1.185 $X2=0 $Y2=0
cc_378 N_A1_c_421_n N_A_760_47#_c_982_n 0.0102636f $X=5 $Y=1.185 $X2=0 $Y2=0
cc_379 N_A1_c_423_n N_A_760_47#_c_982_n 0.00873689f $X=5.43 $Y=1.185 $X2=0 $Y2=0
cc_380 N_A1_c_421_n N_A_760_47#_c_978_n 4.46139e-19 $X=5 $Y=1.185 $X2=0 $Y2=0
cc_381 N_A1_c_423_n N_A_760_47#_c_978_n 0.00627697f $X=5.43 $Y=1.185 $X2=0 $Y2=0
cc_382 N_B1_M1025_g N_B2_M1003_g 0.0366255f $X=6.65 $Y=2.465 $X2=0 $Y2=0
cc_383 N_B1_M1027_g N_B2_M1005_g 0.0202783f $X=6.81 $Y=0.745 $X2=0 $Y2=0
cc_384 B1 B2 0.0179555f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_385 N_B1_c_482_n B2 2.02182e-19 $X=6.81 $Y=1.51 $X2=0 $Y2=0
cc_386 B1 N_B2_c_540_n 0.00307819f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_387 N_B1_c_482_n N_B2_c_540_n 0.0221969f $X=6.81 $Y=1.51 $X2=0 $Y2=0
cc_388 N_B1_M1024_g N_VPWR_c_590_n 0.00357849f $X=6.14 $Y=2.465 $X2=0 $Y2=0
cc_389 N_B1_M1025_g N_VPWR_c_590_n 0.00357877f $X=6.65 $Y=2.465 $X2=0 $Y2=0
cc_390 N_B1_M1024_g N_VPWR_c_575_n 0.00558517f $X=6.14 $Y=2.465 $X2=0 $Y2=0
cc_391 N_B1_M1025_g N_VPWR_c_575_n 0.00600128f $X=6.65 $Y=2.465 $X2=0 $Y2=0
cc_392 N_B1_M1024_g N_A_511_367#_c_783_n 0.00195231f $X=6.14 $Y=2.465 $X2=0
+ $Y2=0
cc_393 N_B1_M1024_g N_A_511_367#_c_785_n 0.0105661f $X=6.14 $Y=2.465 $X2=0 $Y2=0
cc_394 N_B1_M1025_g N_A_511_367#_c_785_n 9.43705e-19 $X=6.65 $Y=2.465 $X2=0
+ $Y2=0
cc_395 N_B1_M1024_g N_A_511_367#_c_756_n 0.0113075f $X=6.14 $Y=2.465 $X2=0 $Y2=0
cc_396 N_B1_M1025_g N_A_511_367#_c_756_n 0.0154449f $X=6.65 $Y=2.465 $X2=0 $Y2=0
cc_397 N_B1_M1027_g N_VGND_c_831_n 5.15399e-19 $X=6.81 $Y=0.745 $X2=0 $Y2=0
cc_398 N_B1_M1009_g N_VGND_c_835_n 0.00302501f $X=6.38 $Y=0.745 $X2=0 $Y2=0
cc_399 N_B1_M1027_g N_VGND_c_835_n 0.00302501f $X=6.81 $Y=0.745 $X2=0 $Y2=0
cc_400 N_B1_M1009_g N_VGND_c_837_n 0.0048466f $X=6.38 $Y=0.745 $X2=0 $Y2=0
cc_401 N_B1_M1027_g N_VGND_c_837_n 0.00435646f $X=6.81 $Y=0.745 $X2=0 $Y2=0
cc_402 N_B1_M1009_g N_A_760_47#_c_978_n 7.55662e-19 $X=6.38 $Y=0.745 $X2=0 $Y2=0
cc_403 N_B1_c_482_n N_A_1208_65#_c_1012_n 3.00519e-19 $X=6.81 $Y=1.51 $X2=0
+ $Y2=0
cc_404 N_B1_M1009_g N_A_1208_65#_c_1013_n 0.0123522f $X=6.38 $Y=0.745 $X2=0
+ $Y2=0
cc_405 N_B1_M1027_g N_A_1208_65#_c_1013_n 0.0118056f $X=6.81 $Y=0.745 $X2=0
+ $Y2=0
cc_406 N_B1_M1027_g N_A_1208_65#_c_1016_n 0.00196541f $X=6.81 $Y=0.745 $X2=0
+ $Y2=0
cc_407 B1 N_A_1208_65#_c_1016_n 0.00969577f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_408 N_B1_c_482_n N_A_1208_65#_c_1016_n 3.83281e-19 $X=6.81 $Y=1.51 $X2=0
+ $Y2=0
cc_409 N_B2_M1003_g N_VPWR_c_590_n 0.00357877f $X=7.23 $Y=2.465 $X2=0 $Y2=0
cc_410 N_B2_M1013_g N_VPWR_c_590_n 0.00357877f $X=7.66 $Y=2.465 $X2=0 $Y2=0
cc_411 N_B2_M1003_g N_VPWR_c_575_n 0.00579264f $X=7.23 $Y=2.465 $X2=0 $Y2=0
cc_412 N_B2_M1013_g N_VPWR_c_575_n 0.00630663f $X=7.66 $Y=2.465 $X2=0 $Y2=0
cc_413 N_B2_M1003_g N_A_511_367#_c_759_n 0.0142672f $X=7.23 $Y=2.465 $X2=0 $Y2=0
cc_414 N_B2_M1013_g N_A_511_367#_c_759_n 0.0115031f $X=7.66 $Y=2.465 $X2=0 $Y2=0
cc_415 B2 N_A_511_367#_c_749_n 0.0189123f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_416 N_B2_M1005_g N_VGND_c_831_n 0.0101655f $X=7.24 $Y=0.745 $X2=0 $Y2=0
cc_417 N_B2_M1022_g N_VGND_c_831_n 0.0107921f $X=7.67 $Y=0.745 $X2=0 $Y2=0
cc_418 N_B2_M1005_g N_VGND_c_835_n 0.00414769f $X=7.24 $Y=0.745 $X2=0 $Y2=0
cc_419 N_B2_M1022_g N_VGND_c_836_n 0.00414769f $X=7.67 $Y=0.745 $X2=0 $Y2=0
cc_420 N_B2_M1005_g N_VGND_c_837_n 0.0078848f $X=7.24 $Y=0.745 $X2=0 $Y2=0
cc_421 N_B2_M1022_g N_VGND_c_837_n 0.00823909f $X=7.67 $Y=0.745 $X2=0 $Y2=0
cc_422 N_B2_M1005_g N_A_1208_65#_c_1013_n 5.73473e-19 $X=7.24 $Y=0.745 $X2=0
+ $Y2=0
cc_423 N_B2_M1005_g N_A_1208_65#_c_1015_n 0.0152975f $X=7.24 $Y=0.745 $X2=0
+ $Y2=0
cc_424 N_B2_M1022_g N_A_1208_65#_c_1015_n 0.0138712f $X=7.67 $Y=0.745 $X2=0
+ $Y2=0
cc_425 B2 N_A_1208_65#_c_1015_n 0.0491085f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_426 N_B2_c_540_n N_A_1208_65#_c_1015_n 0.00276519f $X=7.66 $Y=1.51 $X2=0
+ $Y2=0
cc_427 N_B2_M1022_g N_A_1208_65#_c_1017_n 0.00467043f $X=7.67 $Y=0.745 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_575_n N_X_M1000_s 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_429 N_VPWR_c_575_n N_X_M1016_s 0.00397496f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_430 N_VPWR_M1000_d N_X_c_690_n 0.00262981f $X=0.42 $Y=1.835 $X2=0 $Y2=0
cc_431 N_VPWR_c_576_n N_X_c_690_n 0.0220026f $X=0.545 $Y=2.18 $X2=0 $Y2=0
cc_432 N_VPWR_c_585_n N_X_c_726_n 0.0124525f $X=1.24 $Y=3.33 $X2=0 $Y2=0
cc_433 N_VPWR_c_575_n N_X_c_726_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_M1011_d N_X_c_692_n 0.00176461f $X=1.265 $Y=1.835 $X2=0 $Y2=0
cc_435 N_VPWR_c_577_n N_X_c_692_n 0.0170777f $X=1.405 $Y=2.18 $X2=0 $Y2=0
cc_436 N_VPWR_c_579_n N_X_c_692_n 0.0016373f $X=2.265 $Y=1.98 $X2=0 $Y2=0
cc_437 N_VPWR_c_578_n N_X_c_731_n 0.0138717f $X=2.14 $Y=3.33 $X2=0 $Y2=0
cc_438 N_VPWR_c_575_n N_X_c_731_n 0.00886411f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_439 N_VPWR_c_575_n N_A_511_367#_M1002_s 0.00380103f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_440 N_VPWR_c_575_n N_A_511_367#_M1010_d 0.00371702f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_575_n N_A_511_367#_M1018_d 0.00536646f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_575_n N_A_511_367#_M1023_d 0.00223559f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_575_n N_A_511_367#_M1025_s 0.00348153f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_575_n N_A_511_367#_M1013_d 0.00215161f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_587_n N_A_511_367#_c_767_n 0.0150063f $X=2.96 $Y=3.33 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_575_n N_A_511_367#_c_767_n 0.00950443f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_447 N_VPWR_M1012_d N_A_511_367#_c_746_n 0.00527061f $X=2.985 $Y=1.835 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_580_n N_A_511_367#_c_746_n 0.0220026f $X=3.125 $Y=2.375 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_580_n N_A_511_367#_c_747_n 0.0294086f $X=3.125 $Y=2.375 $X2=0
+ $Y2=0
cc_450 N_VPWR_c_588_n N_A_511_367#_c_747_n 0.0260551f $X=4.41 $Y=3.33 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_575_n N_A_511_367#_c_747_n 0.0145014f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_452 N_VPWR_M1010_s N_A_511_367#_c_753_n 0.00462128f $X=4.435 $Y=1.835 $X2=0
+ $Y2=0
cc_453 N_VPWR_c_581_n N_A_511_367#_c_753_n 0.0170777f $X=4.575 $Y=2.375 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_589_n N_A_511_367#_c_811_n 0.0124525f $X=5.27 $Y=3.33 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_575_n N_A_511_367#_c_811_n 0.00730901f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_456 N_VPWR_M1006_s N_A_511_367#_c_755_n 0.00451678f $X=5.295 $Y=1.835 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_582_n N_A_511_367#_c_755_n 0.0201731f $X=5.435 $Y=2.375 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_590_n N_A_511_367#_c_785_n 0.0180374f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_575_n N_A_511_367#_c_785_n 0.01194f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_460 N_VPWR_c_590_n N_A_511_367#_c_756_n 0.0385732f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_575_n N_A_511_367#_c_756_n 0.0246608f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_590_n N_A_511_367#_c_759_n 0.0363198f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_575_n N_A_511_367#_c_759_n 0.0239346f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_590_n N_A_511_367#_c_748_n 0.0179183f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_575_n N_A_511_367#_c_748_n 0.0101082f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_590_n N_A_511_367#_c_823_n 0.0227155f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_575_n N_A_511_367#_c_823_n 0.0128296f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_468 N_X_c_685_n N_VGND_M1004_s 0.00119058f $X=0.7 $Y=1.13 $X2=-0.19
+ $Y2=-0.245
cc_469 N_X_c_688_n N_VGND_M1004_s 0.00119244f $X=0.217 $Y=1.215 $X2=-0.19
+ $Y2=-0.245
cc_470 N_X_c_686_n N_VGND_M1014_s 0.00176461f $X=1.56 $Y=1.13 $X2=0 $Y2=0
cc_471 N_X_c_685_n N_VGND_c_827_n 0.0109431f $X=0.7 $Y=1.13 $X2=0 $Y2=0
cc_472 N_X_c_688_n N_VGND_c_827_n 0.0122196f $X=0.217 $Y=1.215 $X2=0 $Y2=0
cc_473 N_X_c_686_n N_VGND_c_828_n 0.0170777f $X=1.56 $Y=1.13 $X2=0 $Y2=0
cc_474 N_X_c_711_n N_VGND_c_829_n 0.0455102f $X=1.655 $Y=0.42 $X2=0 $Y2=0
cc_475 N_X_c_740_p N_VGND_c_832_n 0.0124525f $X=0.795 $Y=0.42 $X2=0 $Y2=0
cc_476 N_X_c_711_n N_VGND_c_833_n 0.015688f $X=1.655 $Y=0.42 $X2=0 $Y2=0
cc_477 N_X_M1004_d N_VGND_c_837_n 0.00536646f $X=0.655 $Y=0.235 $X2=0 $Y2=0
cc_478 N_X_M1017_d N_VGND_c_837_n 0.00380103f $X=1.515 $Y=0.235 $X2=0 $Y2=0
cc_479 N_X_c_740_p N_VGND_c_837_n 0.00730901f $X=0.795 $Y=0.42 $X2=0 $Y2=0
cc_480 N_X_c_711_n N_VGND_c_837_n 0.00984745f $X=1.655 $Y=0.42 $X2=0 $Y2=0
cc_481 N_A_511_367#_c_749_n N_A_1208_65#_c_1015_n 0.00120798f $X=7.875 $Y=2.085
+ $X2=0 $Y2=0
cc_482 N_VGND_c_837_n N_A_511_47#_M1007_d 0.00223559f $X=7.92 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_483 N_VGND_c_837_n N_A_511_47#_M1001_d 0.00223577f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_484 N_VGND_c_829_n N_A_511_47#_c_946_n 0.0341642f $X=2.175 $Y=0.38 $X2=0
+ $Y2=0
cc_485 N_VGND_c_834_n N_A_511_47#_c_946_n 0.0188748f $X=3.03 $Y=0 $X2=0 $Y2=0
cc_486 N_VGND_c_837_n N_A_511_47#_c_946_n 0.012371f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_M1026_s N_A_511_47#_c_939_n 0.00524506f $X=2.985 $Y=0.235 $X2=0
+ $Y2=0
cc_488 N_VGND_c_830_n N_A_511_47#_c_939_n 0.0154494f $X=3.125 $Y=0.4 $X2=0 $Y2=0
cc_489 N_VGND_c_834_n N_A_511_47#_c_939_n 0.00196209f $X=3.03 $Y=0 $X2=0 $Y2=0
cc_490 N_VGND_c_835_n N_A_511_47#_c_939_n 0.00251343f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_491 N_VGND_c_837_n N_A_511_47#_c_939_n 0.00913588f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_492 N_VGND_c_829_n N_A_511_47#_c_944_n 0.0128488f $X=2.175 $Y=0.38 $X2=0
+ $Y2=0
cc_493 N_VGND_c_830_n N_A_511_47#_c_940_n 0.00371907f $X=3.125 $Y=0.4 $X2=0
+ $Y2=0
cc_494 N_VGND_c_830_n N_A_511_47#_c_941_n 0.0219184f $X=3.125 $Y=0.4 $X2=0 $Y2=0
cc_495 N_VGND_c_835_n N_A_511_47#_c_941_n 0.0121451f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_496 N_VGND_c_837_n N_A_511_47#_c_941_n 0.00660136f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_497 N_VGND_c_835_n N_A_511_47#_c_942_n 0.0560141f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_498 N_VGND_c_837_n N_A_511_47#_c_942_n 0.0347267f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_499 N_VGND_c_837_n N_A_760_47#_M1001_s 0.0021598f $X=7.92 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_500 N_VGND_c_837_n N_A_760_47#_M1008_s 0.00242554f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_501 N_VGND_c_837_n N_A_760_47#_M1020_s 0.00215158f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_502 N_VGND_c_835_n N_A_760_47#_c_977_n 0.00222753f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_503 N_VGND_c_837_n N_A_760_47#_c_977_n 0.00539228f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_504 N_VGND_c_835_n N_A_760_47#_c_999_n 0.013043f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_505 N_VGND_c_837_n N_A_760_47#_c_999_n 0.00796681f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_506 N_VGND_c_835_n N_A_760_47#_c_982_n 0.0326653f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_507 N_VGND_c_837_n N_A_760_47#_c_982_n 0.0207161f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_508 N_VGND_c_835_n N_A_760_47#_c_978_n 0.0209663f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_509 N_VGND_c_837_n N_A_760_47#_c_978_n 0.0125896f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_510 N_VGND_c_831_n N_A_1208_65#_c_1013_n 0.00962585f $X=7.455 $Y=0.45 $X2=0
+ $Y2=0
cc_511 N_VGND_c_835_n N_A_1208_65#_c_1013_n 0.0558492f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_512 N_VGND_c_837_n N_A_1208_65#_c_1013_n 0.0312041f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_c_835_n N_A_1208_65#_c_1014_n 0.0184178f $X=7.29 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_837_n N_A_1208_65#_c_1014_n 0.0100667f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_515 N_VGND_M1005_d N_A_1208_65#_c_1015_n 0.00176461f $X=7.315 $Y=0.325 $X2=0
+ $Y2=0
cc_516 N_VGND_c_831_n N_A_1208_65#_c_1015_n 0.0170777f $X=7.455 $Y=0.45 $X2=0
+ $Y2=0
cc_517 N_VGND_c_831_n N_A_1208_65#_c_1017_n 0.0271585f $X=7.455 $Y=0.45 $X2=0
+ $Y2=0
cc_518 N_VGND_c_836_n N_A_1208_65#_c_1017_n 0.0184952f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_837_n N_A_1208_65#_c_1017_n 0.0100304f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_520 N_A_511_47#_c_942_n N_A_760_47#_M1001_s 0.00543849f $X=4.355 $Y=0.375
+ $X2=-0.19 $Y2=-0.245
cc_521 N_A_511_47#_M1001_d N_A_760_47#_c_977_n 0.00340978f $X=4.215 $Y=0.235
+ $X2=0 $Y2=0
cc_522 N_A_511_47#_c_939_n N_A_760_47#_c_977_n 0.0143023f $X=3.41 $Y=0.82 $X2=0
+ $Y2=0
cc_523 N_A_511_47#_c_940_n N_A_760_47#_c_977_n 0.00393781f $X=3.495 $Y=0.735
+ $X2=0 $Y2=0
cc_524 N_A_511_47#_c_942_n N_A_760_47#_c_977_n 0.042109f $X=4.355 $Y=0.375 $X2=0
+ $Y2=0
cc_525 N_A_760_47#_c_978_n N_A_1208_65#_c_1012_n 0.0310308f $X=5.645 $Y=0.38
+ $X2=0 $Y2=0
cc_526 N_A_760_47#_c_978_n N_A_1208_65#_c_1014_n 0.0147157f $X=5.645 $Y=0.38
+ $X2=0 $Y2=0
