* File: sky130_fd_sc_lp__o221a_1.spice
* Created: Wed Sep  2 10:18:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221a_1.pex.spice"
.subckt sky130_fd_sc_lp__o221a_1  VNB VPB C1 B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1002 N_A_179_49#_M1002_d N_C1_M1002_g N_A_96_49#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1344 AS=0.2226 PD=1.16 PS=2.21 NRD=4.284 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1010 N_A_273_49#_M1010_d N_B1_M1010_g N_A_179_49#_M1002_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=1.428 M=1 R=5.6
+ SA=75000.7 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1004 N_A_179_49#_M1004_d N_B2_M1004_g N_A_273_49#_M1010_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_273_49#_M1007_d N_A2_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A1_M1011_g N_A_273_49#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1005 N_X_M1005_d N_A_96_49#_M1005_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1344 PD=2.21 PS=1.16 NRD=0 NRS=5.712 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_C1_M1003_g N_A_96_49#_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.3339 PD=1.65 PS=3.05 NRD=8.5892 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003 A=0.189 P=2.82 MULT=1
MM1006 A_287_367# N_B1_M1006_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.2457 PD=1.5 PS=1.65 NRD=10.1455 NRS=8.5892 M=1 R=8.4 SA=75000.7
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1000 N_A_96_49#_M1000_d N_B2_M1000_g A_287_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4851 AS=0.1512 PD=2.03 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75001.1
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1001 A_549_367# N_A2_M1001_g N_A_96_49#_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.4851 PD=1.47 PS=2.03 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75002
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_549_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.1323 PD=1.685 PS=1.47 NRD=9.3772 NRS=7.8012 M=1 R=8.4
+ SA=75002.4 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1009 N_X_M1009_d N_A_96_49#_M1009_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.26775 PD=3.09 PS=1.685 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75003
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__o221a_1.pxi.spice"
*
.ends
*
*
