* NGSPICE file created from sky130_fd_sc_lp__a211o_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_80_237# C1 a_504_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=3.402e+11p ps=3.06e+06u
M1001 a_80_237# A1 a_294_47# VNB nshort w=840000u l=150000u
+  ad=5.754e+11p pd=4.73e+06u as=2.016e+11p ps=2.16e+06u
M1002 a_294_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=9.156e+11p ps=5.54e+06u
M1003 VPWR A2 a_217_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.875e+11p pd=6.29e+06u as=7.875e+11p ps=6.29e+06u
M1004 a_217_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_504_367# B1 a_217_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B1 a_80_237# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_80_237# C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_80_237# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1009 VGND a_80_237# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
.ends

