* File: sky130_fd_sc_lp__o211ai_lp.pex.spice
* Created: Wed Sep  2 10:14:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211AI_LP%A1 3 7 12 13 14 15 19
r32 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.46
+ $Y=1.335 $X2=0.46 $Y2=1.335
r33 15 20 7.89412 $w=4.98e-07 $l=3.3e-07 $layer=LI1_cond $X=0.375 $Y=1.665
+ $X2=0.375 $Y2=1.335
r34 14 20 0.956863 $w=4.98e-07 $l=4e-08 $layer=LI1_cond $X=0.375 $Y=1.295
+ $X2=0.375 $Y2=1.335
r35 12 19 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.46 $Y=1.69
+ $X2=0.46 $Y2=1.335
r36 12 13 29.7575 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.49 $Y=1.69
+ $X2=0.49 $Y2=1.84
r37 10 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.46 $Y=1.17
+ $X2=0.46 $Y2=1.335
r38 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.55 $Y=0.495
+ $X2=0.55 $Y2=1.17
r39 3 13 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.56 $Y=2.545
+ $X2=0.56 $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_LP%A2 3 7 11 12 13 14 18
r41 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.09
+ $Y=1.335 $X2=1.09 $Y2=1.335
r42 14 19 9.75144 $w=3.88e-07 $l=3.3e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.335
r43 13 19 1.18199 $w=3.88e-07 $l=4e-08 $layer=LI1_cond $X=1.12 $Y=1.295 $X2=1.12
+ $Y2=1.335
r44 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.09 $Y=1.675
+ $X2=1.09 $Y2=1.335
r45 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.675
+ $X2=1.09 $Y2=1.84
r46 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.17
+ $X2=1.09 $Y2=1.335
r47 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.14 $Y=0.495
+ $X2=1.14 $Y2=1.17
r48 3 12 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.05 $Y=2.545
+ $X2=1.05 $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_LP%B1 3 7 11 12 13 14 18
r43 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=1.295
+ $X2=1.66 $Y2=1.665
r44 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.66
+ $Y=1.335 $X2=1.66 $Y2=1.335
r45 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.66 $Y=1.675
+ $X2=1.66 $Y2=1.335
r46 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.675
+ $X2=1.66 $Y2=1.84
r47 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.17
+ $X2=1.66 $Y2=1.335
r48 7 12 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.62 $Y=2.545
+ $X2=1.62 $Y2=1.84
r49 3 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.57 $Y=0.495
+ $X2=1.57 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_LP%C1 1 3 8 12 15 16 17 18 19 23
r45 18 19 12.8415 $w=3.48e-07 $l=3.9e-07 $layer=LI1_cond $X=2.22 $Y=1.275
+ $X2=2.22 $Y2=1.665
r46 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23
+ $Y=1.275 $X2=2.23 $Y2=1.275
r47 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.23 $Y=1.615
+ $X2=2.23 $Y2=1.275
r48 16 17 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.615
+ $X2=2.23 $Y2=1.78
r49 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.11
+ $X2=2.23 $Y2=1.275
r50 10 12 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.96 $Y=0.855
+ $X2=2.14 $Y2=0.855
r51 8 17 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.19 $Y=2.545
+ $X2=2.19 $Y2=1.78
r52 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.14 $Y=0.93 $X2=2.14
+ $Y2=0.855
r53 4 15 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.14 $Y=0.93 $X2=2.14
+ $Y2=1.11
r54 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=0.78 $X2=1.96
+ $Y2=0.855
r55 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.96 $Y=0.78 $X2=1.96
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_LP%VPWR 1 2 7 9 15 18 19 20 30 31
r31 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r37 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 22 34 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=3.33 $X2=0.23
+ $Y2=3.33
r39 22 24 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 20 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 18 27 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r43 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=1.885 $Y2=3.33
r44 17 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.05 $Y=3.33 $X2=2.64
+ $Y2=3.33
r45 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.05 $Y=3.33
+ $X2=1.885 $Y2=3.33
r46 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=3.245
+ $X2=1.885 $Y2=3.33
r47 13 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.885 $Y=3.245
+ $X2=1.885 $Y2=2.535
r48 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.295 $Y=2.19
+ $X2=0.295 $Y2=2.9
r49 7 34 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.23 $Y2=3.33
r50 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.9
r51 2 15 300 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=2 $X=1.745
+ $Y=2.045 $X2=1.885 $Y2=2.535
r52 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.045 $X2=0.295 $Y2=2.9
r53 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.045 $X2=0.295 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_LP%Y 1 2 3 14 16 17 22 24 25 26 27 28 32
r50 28 32 2.39909 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=0.495
+ $X2=2.585 $Y2=0.495
r51 28 32 0.390026 $w=4.58e-07 $l=1.5e-08 $layer=LI1_cond $X=2.57 $Y=0.495
+ $X2=2.585 $Y2=0.495
r52 27 28 10.6607 $w=4.58e-07 $l=4.1e-07 $layer=LI1_cond $X=2.16 $Y=0.495
+ $X2=2.57 $Y2=0.495
r53 25 26 2.99104 $w=3.17e-07 $l=1.85699e-07 $layer=LI1_cond $X=2.67 $Y=2.02
+ $X2=2.522 $Y2=2.105
r54 24 28 6.49166 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.67 $Y=0.725
+ $X2=2.67 $Y2=0.495
r55 24 25 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=2.67 $Y=0.725
+ $X2=2.67 $Y2=2.02
r56 20 26 2.99104 $w=3.17e-07 $l=8.5e-08 $layer=LI1_cond $X=2.522 $Y=2.19
+ $X2=2.522 $Y2=2.105
r57 20 22 18.2627 $w=4.63e-07 $l=7.1e-07 $layer=LI1_cond $X=2.522 $Y=2.19
+ $X2=2.522 $Y2=2.9
r58 16 26 3.66292 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=2.29 $Y=2.105
+ $X2=2.522 $Y2=2.105
r59 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.29 $Y=2.105
+ $X2=1.52 $Y2=2.105
r60 12 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.355 $Y=2.19
+ $X2=1.52 $Y2=2.105
r61 12 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.355 $Y=2.19
+ $X2=1.355 $Y2=2.9
r62 3 22 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=2.045 $X2=2.455 $Y2=2.9
r63 3 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=2.045 $X2=2.455 $Y2=2.19
r64 2 14 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=2.045 $X2=1.355 $Y2=2.9
r65 2 12 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=2.045 $X2=1.355 $Y2=2.19
r66 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.035
+ $Y=0.285 $X2=2.175 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_LP%A_38_57# 1 2 9 11 12 15
r31 13 15 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.355 $Y=0.82
+ $X2=1.355 $Y2=0.495
r32 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.19 $Y=0.905
+ $X2=1.355 $Y2=0.82
r33 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.19 $Y=0.905 $X2=0.5
+ $Y2=0.905
r34 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.335 $Y=0.82
+ $X2=0.5 $Y2=0.905
r35 7 9 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.335 $Y=0.82
+ $X2=0.335 $Y2=0.495
r36 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.285 $X2=1.355 $Y2=0.495
r37 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.285 $X2=0.335 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_LP%VGND 1 8 10 17 18 21
r26 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r27 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r28 15 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r29 14 17 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r30 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r31 12 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.845
+ $Y2=0
r32 12 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.2
+ $Y2=0
r33 10 18 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r34 10 15 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r35 6 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=0.085
+ $X2=0.845 $Y2=0
r36 6 8 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.845 $Y=0.085
+ $X2=0.845 $Y2=0.45
r37 1 8 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.285 $X2=0.845 $Y2=0.45
.ends

