* File: sky130_fd_sc_lp__o32a_1.pex.spice
* Created: Fri Aug 28 11:17:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32A_1%A_88_269# 1 2 9 13 16 17 18 21 25 27 30 33 35
+ 38 39
c87 35 0 5.97642e-20 $X=0.815 $Y=1.495
c88 16 0 1.58015e-19 $X=0.815 $Y=1.93
r89 33 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.51
+ $X2=0.605 $Y2=1.675
r90 33 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.51
+ $X2=0.605 $Y2=1.345
r91 32 35 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=0.605 $Y=1.495
+ $X2=0.815 $Y2=1.495
r92 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.51 $X2=0.605 $Y2=1.51
r93 30 39 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.175 $Y=1.93
+ $X2=3.175 $Y2=1.175
r94 28 38 13.6095 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=2.91 $Y=2.015
+ $X2=2.562 $Y2=2.015
r95 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.09 $Y=2.015
+ $X2=3.175 $Y2=1.93
r96 27 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.09 $Y=2.015
+ $X2=2.91 $Y2=2.015
r97 23 39 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=3.08 $Y=0.995
+ $X2=3.08 $Y2=1.175
r98 23 25 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=3.08 $Y=0.995
+ $X2=3.08 $Y2=0.72
r99 19 38 2.84707 $w=6.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.562 $Y=2.1
+ $X2=2.562 $Y2=2.015
r100 19 21 14.6283 $w=6.93e-07 $l=8.5e-07 $layer=LI1_cond $X=2.562 $Y=2.1
+ $X2=2.562 $Y2=2.95
r101 17 38 13.6095 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=2.215 $Y=2.015
+ $X2=2.562 $Y2=2.015
r102 17 18 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=2.215 $Y=2.015
+ $X2=0.9 $Y2=2.015
r103 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.815 $Y=1.93
+ $X2=0.9 $Y2=2.015
r104 15 35 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.815 $Y=1.645
+ $X2=0.815 $Y2=1.495
r105 15 16 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.815 $Y=1.645
+ $X2=0.815 $Y2=1.93
r106 13 41 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.695 $Y=0.765
+ $X2=0.695 $Y2=1.345
r107 9 42 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.69 $Y=2.465
+ $X2=0.69 $Y2=1.675
r108 2 38 200 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=3 $X=2.25
+ $Y=1.835 $X2=2.39 $Y2=2.015
r109 2 21 200 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=3 $X=2.25
+ $Y=1.835 $X2=2.39 $Y2=2.95
r110 1 25 91 $w=1.7e-07 $l=4.58258e-07 $layer=licon1_NDIFF $count=2 $X=2.88
+ $Y=0.345 $X2=3.065 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_1%A1 3 6 8 9 13 15
c39 6 0 1.13962e-19 $X=1.245 $Y=2.465
r40 13 16 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.46
+ $X2=1.15 $Y2=1.625
r41 13 15 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.46
+ $X2=1.15 $Y2=1.295
r42 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.46 $X2=1.155 $Y2=1.46
r43 9 14 8.2895 $w=2.83e-07 $l=2.05e-07 $layer=LI1_cond $X=1.212 $Y=1.665
+ $X2=1.212 $Y2=1.46
r44 8 14 6.67204 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.212 $Y=1.295
+ $X2=1.212 $Y2=1.46
r45 6 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.245 $Y=2.465
+ $X2=1.245 $Y2=1.625
r46 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.175 $Y=0.765
+ $X2=1.175 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_1%A2 3 6 8 9 13 15
c36 8 0 4.06102e-19 $X=1.68 $Y=1.295
r37 13 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.46
+ $X2=1.71 $Y2=1.625
r38 13 15 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.46
+ $X2=1.71 $Y2=1.295
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.46 $X2=1.725 $Y2=1.46
r40 9 14 7.38284 $w=3.18e-07 $l=2.05e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=1.46
r41 8 14 5.94228 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.295
+ $X2=1.685 $Y2=1.46
r42 6 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.715 $Y=2.465
+ $X2=1.715 $Y2=1.625
r43 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.605 $Y=0.765
+ $X2=1.605 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_1%A3 3 5 7 8 9 17
c39 8 0 1.77524e-19 $X=2.16 $Y=1.295
c40 5 0 1.93889e-19 $X=2.375 $Y=1.295
r41 15 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.285 $Y=1.46
+ $X2=2.375 $Y2=1.46
r42 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.285
+ $Y=1.46 $X2=2.285 $Y2=1.46
r43 12 15 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=2.175 $Y=1.46
+ $X2=2.285 $Y2=1.46
r44 9 16 6.65495 $w=3.53e-07 $l=2.05e-07 $layer=LI1_cond $X=2.192 $Y=1.665
+ $X2=2.192 $Y2=1.46
r45 8 16 5.35643 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.192 $Y=1.295
+ $X2=2.192 $Y2=1.46
r46 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.295
+ $X2=2.375 $Y2=1.46
r47 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.375 $Y=1.295
+ $X2=2.375 $Y2=0.765
r48 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.175 $Y=1.625
+ $X2=2.175 $Y2=1.46
r49 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.175 $Y=1.625
+ $X2=2.175 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_1%B2 3 7 9 12 13
c39 7 0 1.77524e-19 $X=2.945 $Y=2.465
r40 12 15 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.51
+ $X2=2.84 $Y2=1.675
r41 12 14 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.51
+ $X2=2.84 $Y2=1.345
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.825
+ $Y=1.51 $X2=2.825 $Y2=1.51
r43 9 13 5.1374 $w=4.13e-07 $l=1.85e-07 $layer=LI1_cond $X=2.64 $Y=1.552
+ $X2=2.825 $Y2=1.552
r44 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.945 $Y=2.465
+ $X2=2.945 $Y2=1.675
r45 3 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.805 $Y=0.765
+ $X2=2.805 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_1%B1 1 3 6 8 9 10 17
r31 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.525
+ $Y=1.46 $X2=3.525 $Y2=1.46
r32 14 17 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.305 $Y=1.46
+ $X2=3.525 $Y2=1.46
r33 9 10 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.597 $Y=1.665
+ $X2=3.597 $Y2=2.035
r34 9 18 7.50003 $w=3.13e-07 $l=2.05e-07 $layer=LI1_cond $X=3.597 $Y=1.665
+ $X2=3.597 $Y2=1.46
r35 8 18 6.03661 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.597 $Y=1.295
+ $X2=3.597 $Y2=1.46
r36 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.625
+ $X2=3.305 $Y2=1.46
r37 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.305 $Y=1.625
+ $X2=3.305 $Y2=2.465
r38 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.295
+ $X2=3.305 $Y2=1.46
r39 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.305 $Y=1.295
+ $X2=3.305 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_1%X 1 2 11 14 15 16 17 23 29
r24 21 29 0.162574 $w=5.13e-07 $l=7e-09 $layer=LI1_cond $X=0.342 $Y=0.918
+ $X2=0.342 $Y2=0.925
r25 17 31 10.2774 $w=5.13e-07 $l=2.11e-07 $layer=LI1_cond $X=0.342 $Y=0.964
+ $X2=0.342 $Y2=1.175
r26 17 29 0.905768 $w=5.13e-07 $l=3.9e-08 $layer=LI1_cond $X=0.342 $Y=0.964
+ $X2=0.342 $Y2=0.925
r27 17 21 0.905768 $w=5.13e-07 $l=3.9e-08 $layer=LI1_cond $X=0.342 $Y=0.879
+ $X2=0.342 $Y2=0.918
r28 16 17 7.52484 $w=5.13e-07 $l=3.24e-07 $layer=LI1_cond $X=0.342 $Y=0.555
+ $X2=0.342 $Y2=0.879
r29 16 23 1.50961 $w=5.13e-07 $l=6.5e-08 $layer=LI1_cond $X=0.342 $Y=0.555
+ $X2=0.342 $Y2=0.49
r30 15 31 39.4343 $w=1.78e-07 $l=6.4e-07 $layer=LI1_cond $X=0.175 $Y=1.815
+ $X2=0.175 $Y2=1.175
r31 14 15 8.97208 $w=4.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.322 $Y=1.98
+ $X2=0.322 $Y2=1.815
r32 9 14 1.813 $w=4.73e-07 $l=7.2e-08 $layer=LI1_cond $X=0.322 $Y=2.052
+ $X2=0.322 $Y2=1.98
r33 9 11 21.605 $w=4.73e-07 $l=8.58e-07 $layer=LI1_cond $X=0.322 $Y=2.052
+ $X2=0.322 $Y2=2.91
r34 2 14 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=1.835 $X2=0.455 $Y2=1.98
r35 2 11 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=1.835 $X2=0.455 $Y2=2.91
r36 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.335
+ $Y=0.345 $X2=0.48 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_1%VPWR 1 2 9 11 13 16 17 18 24 33
r42 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 26 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 24 32 4.65202 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.597 $Y2=3.33
r48 24 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 18 30 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 16 21 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.8 $Y=3.33 $X2=0.72
+ $Y2=3.33
r54 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.8 $Y=3.33
+ $X2=0.965 $Y2=3.33
r55 15 26 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.13 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.13 $Y=3.33
+ $X2=0.965 $Y2=3.33
r57 11 32 3.11416 $w=3.3e-07 $l=1.17346e-07 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.597 $Y2=3.33
r58 11 13 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=2.4
r59 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=3.245
+ $X2=0.965 $Y2=3.33
r60 7 9 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.965 $Y=3.245
+ $X2=0.965 $Y2=2.395
r61 2 13 300 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=2 $X=3.38
+ $Y=1.835 $X2=3.52 $Y2=2.4
r62 1 9 300 $w=1.7e-07 $l=6.5238e-07 $layer=licon1_PDIFF $count=2 $X=0.765
+ $Y=1.835 $X2=0.965 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_1%VGND 1 2 9 11 13 14 15 26 27 31
r41 31 36 10.3541 $w=6.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.99 $Y=0 $X2=1.99
+ $Y2=0.58
r42 31 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r43 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r44 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 24 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r46 24 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r47 23 26 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r48 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r49 21 31 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=1.99
+ $Y2=0
r50 21 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.64
+ $Y2=0
r51 19 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r52 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 15 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r54 15 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r55 13 18 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.77 $Y=0 $X2=0.72
+ $Y2=0
r56 13 14 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=0 $X2=0.935
+ $Y2=0
r57 12 14 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=0 $X2=0.935
+ $Y2=0
r58 11 31 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.99
+ $Y2=0
r59 11 12 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.1
+ $Y2=0
r60 7 14 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0
r61 7 9 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0.47
r62 2 36 91 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_NDIFF $count=2 $X=1.68
+ $Y=0.345 $X2=2.16 $Y2=0.58
r63 1 9 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.77
+ $Y=0.345 $X2=0.935 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_1%A_250_69# 1 2 3 12 14 15 20 21 24
r35 22 24 1.85214 $w=2.78e-07 $l=4.5e-08 $layer=LI1_cond $X=3.57 $Y=0.425
+ $X2=3.57 $Y2=0.47
r36 20 22 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.43 $Y=0.34
+ $X2=3.57 $Y2=0.425
r37 20 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.43 $Y=0.34 $X2=2.73
+ $Y2=0.34
r38 17 19 19.6161 $w=2.33e-07 $l=4e-07 $layer=LI1_cond $X=2.612 $Y=0.87
+ $X2=2.612 $Y2=0.47
r39 16 21 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=2.612 $Y=0.425
+ $X2=2.73 $Y2=0.34
r40 16 19 2.20681 $w=2.33e-07 $l=4.5e-08 $layer=LI1_cond $X=2.612 $Y=0.425
+ $X2=2.612 $Y2=0.47
r41 14 17 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.495 $Y=0.955
+ $X2=2.612 $Y2=0.87
r42 14 15 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.495 $Y=0.955
+ $X2=1.485 $Y2=0.955
r43 10 15 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=1.377 $Y=0.87
+ $X2=1.485 $Y2=0.955
r44 10 12 21.4408 $w=2.13e-07 $l=4e-07 $layer=LI1_cond $X=1.377 $Y=0.87
+ $X2=1.377 $Y2=0.47
r45 3 24 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=3.38
+ $Y=0.345 $X2=3.545 $Y2=0.47
r46 2 19 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.45
+ $Y=0.345 $X2=2.59 $Y2=0.47
r47 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.25
+ $Y=0.345 $X2=1.39 $Y2=0.47
.ends

