* File: sky130_fd_sc_lp__dlrbn_2.pxi.spice
* Created: Fri Aug 28 10:25:40 2020
* 
x_PM_SKY130_FD_SC_LP__DLRBN_2%GATE_N N_GATE_N_c_188_n N_GATE_N_M1007_g
+ N_GATE_N_M1026_g N_GATE_N_c_194_n GATE_N GATE_N GATE_N GATE_N N_GATE_N_c_190_n
+ N_GATE_N_c_191_n PM_SKY130_FD_SC_LP__DLRBN_2%GATE_N
x_PM_SKY130_FD_SC_LP__DLRBN_2%A_113_144# N_A_113_144#_M1007_d
+ N_A_113_144#_M1026_d N_A_113_144#_c_219_n N_A_113_144#_M1016_g
+ N_A_113_144#_M1012_g N_A_113_144#_c_229_n N_A_113_144#_M1025_g
+ N_A_113_144#_c_231_n N_A_113_144#_M1024_g N_A_113_144#_c_222_n
+ N_A_113_144#_c_223_n N_A_113_144#_c_233_n N_A_113_144#_c_224_n
+ N_A_113_144#_c_225_n N_A_113_144#_c_235_n N_A_113_144#_c_236_n
+ N_A_113_144#_c_226_n N_A_113_144#_c_227_n N_A_113_144#_c_237_n
+ PM_SKY130_FD_SC_LP__DLRBN_2%A_113_144#
x_PM_SKY130_FD_SC_LP__DLRBN_2%D N_D_c_322_n N_D_M1017_g N_D_M1008_g D D
+ N_D_c_325_n PM_SKY130_FD_SC_LP__DLRBN_2%D
x_PM_SKY130_FD_SC_LP__DLRBN_2%A_162_40# N_A_162_40#_M1016_s N_A_162_40#_M1012_s
+ N_A_162_40#_c_356_n N_A_162_40#_M1019_g N_A_162_40#_c_358_n
+ N_A_162_40#_c_359_n N_A_162_40#_M1015_g N_A_162_40#_c_361_n
+ N_A_162_40#_c_362_n N_A_162_40#_c_367_n N_A_162_40#_c_368_n
+ N_A_162_40#_c_363_n N_A_162_40#_c_364_n N_A_162_40#_c_365_n
+ PM_SKY130_FD_SC_LP__DLRBN_2%A_162_40#
x_PM_SKY130_FD_SC_LP__DLRBN_2%A_392_144# N_A_392_144#_M1017_d
+ N_A_392_144#_M1008_d N_A_392_144#_c_437_n N_A_392_144#_c_438_n
+ N_A_392_144#_c_439_n N_A_392_144#_M1018_g N_A_392_144#_c_441_n
+ N_A_392_144#_M1014_g N_A_392_144#_c_442_n N_A_392_144#_c_450_n
+ N_A_392_144#_c_451_n N_A_392_144#_c_443_n N_A_392_144#_c_444_n
+ N_A_392_144#_c_445_n N_A_392_144#_c_446_n N_A_392_144#_c_447_n
+ N_A_392_144#_c_448_n PM_SKY130_FD_SC_LP__DLRBN_2%A_392_144#
x_PM_SKY130_FD_SC_LP__DLRBN_2%A_942_252# N_A_942_252#_M1027_s
+ N_A_942_252#_M1020_d N_A_942_252#_M1005_g N_A_942_252#_M1004_g
+ N_A_942_252#_M1009_g N_A_942_252#_M1000_g N_A_942_252#_M1022_g
+ N_A_942_252#_M1021_g N_A_942_252#_M1010_g N_A_942_252#_M1011_g
+ N_A_942_252#_c_532_n N_A_942_252#_c_533_n N_A_942_252#_c_534_n
+ N_A_942_252#_c_535_n N_A_942_252#_c_536_n N_A_942_252#_c_537_n
+ N_A_942_252#_c_548_n N_A_942_252#_c_568_p N_A_942_252#_c_558_p
+ N_A_942_252#_c_549_n N_A_942_252#_c_646_p N_A_942_252#_c_550_n
+ N_A_942_252#_c_538_n N_A_942_252#_c_539_n N_A_942_252#_c_540_n
+ N_A_942_252#_c_578_p PM_SKY130_FD_SC_LP__DLRBN_2%A_942_252#
x_PM_SKY130_FD_SC_LP__DLRBN_2%A_591_155# N_A_591_155#_M1025_d
+ N_A_591_155#_M1024_d N_A_591_155#_c_681_n N_A_591_155#_c_682_n
+ N_A_591_155#_c_674_n N_A_591_155#_c_675_n N_A_591_155#_M1027_g
+ N_A_591_155#_c_685_n N_A_591_155#_M1020_g N_A_591_155#_c_677_n
+ N_A_591_155#_c_678_n N_A_591_155#_c_688_n N_A_591_155#_c_689_n
+ N_A_591_155#_c_679_n N_A_591_155#_c_680_n N_A_591_155#_c_690_n
+ N_A_591_155#_c_691_n N_A_591_155#_c_692_n
+ PM_SKY130_FD_SC_LP__DLRBN_2%A_591_155#
x_PM_SKY130_FD_SC_LP__DLRBN_2%RESET_B N_RESET_B_M1002_g N_RESET_B_M1006_g
+ RESET_B RESET_B RESET_B N_RESET_B_c_777_n N_RESET_B_c_778_n
+ PM_SKY130_FD_SC_LP__DLRBN_2%RESET_B
x_PM_SKY130_FD_SC_LP__DLRBN_2%A_1555_367# N_A_1555_367#_M1011_d
+ N_A_1555_367#_M1010_d N_A_1555_367#_M1003_g N_A_1555_367#_M1001_g
+ N_A_1555_367#_c_814_n N_A_1555_367#_M1013_g N_A_1555_367#_M1023_g
+ N_A_1555_367#_c_817_n N_A_1555_367#_c_823_n N_A_1555_367#_c_818_n
+ N_A_1555_367#_c_824_n N_A_1555_367#_c_825_n N_A_1555_367#_c_819_n
+ N_A_1555_367#_c_820_n PM_SKY130_FD_SC_LP__DLRBN_2%A_1555_367#
x_PM_SKY130_FD_SC_LP__DLRBN_2%VPWR N_VPWR_M1026_s N_VPWR_M1012_d N_VPWR_M1018_d
+ N_VPWR_M1020_s N_VPWR_M1006_d N_VPWR_M1021_s N_VPWR_M1001_s N_VPWR_M1023_s
+ N_VPWR_c_878_n N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n N_VPWR_c_882_n
+ N_VPWR_c_883_n N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n N_VPWR_c_887_n
+ N_VPWR_c_888_n N_VPWR_c_889_n N_VPWR_c_890_n N_VPWR_c_891_n VPWR
+ N_VPWR_c_892_n N_VPWR_c_893_n N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n
+ N_VPWR_c_897_n N_VPWR_c_898_n N_VPWR_c_899_n N_VPWR_c_900_n N_VPWR_c_877_n
+ PM_SKY130_FD_SC_LP__DLRBN_2%VPWR
x_PM_SKY130_FD_SC_LP__DLRBN_2%A_606_359# N_A_606_359#_M1024_s
+ N_A_606_359#_M1005_d N_A_606_359#_c_1003_n N_A_606_359#_c_1004_n
+ N_A_606_359#_c_1005_n PM_SKY130_FD_SC_LP__DLRBN_2%A_606_359#
x_PM_SKY130_FD_SC_LP__DLRBN_2%Q N_Q_M1009_d N_Q_M1000_d N_Q_c_1038_n
+ N_Q_c_1040_n N_Q_c_1039_n Q N_Q_c_1057_n PM_SKY130_FD_SC_LP__DLRBN_2%Q
x_PM_SKY130_FD_SC_LP__DLRBN_2%Q_N N_Q_N_M1003_s N_Q_N_M1001_d Q_N Q_N Q_N Q_N
+ Q_N N_Q_N_c_1066_n PM_SKY130_FD_SC_LP__DLRBN_2%Q_N
x_PM_SKY130_FD_SC_LP__DLRBN_2%VGND N_VGND_M1007_s N_VGND_M1016_d N_VGND_M1014_d
+ N_VGND_M1002_d N_VGND_M1022_s N_VGND_M1003_d N_VGND_M1013_d N_VGND_c_1084_n
+ N_VGND_c_1085_n N_VGND_c_1086_n N_VGND_c_1087_n N_VGND_c_1088_n
+ N_VGND_c_1089_n N_VGND_c_1090_n N_VGND_c_1091_n N_VGND_c_1092_n VGND
+ N_VGND_c_1093_n N_VGND_c_1094_n N_VGND_c_1095_n N_VGND_c_1096_n
+ N_VGND_c_1097_n N_VGND_c_1098_n N_VGND_c_1099_n N_VGND_c_1100_n
+ N_VGND_c_1101_n N_VGND_c_1102_n N_VGND_c_1103_n N_VGND_c_1104_n
+ PM_SKY130_FD_SC_LP__DLRBN_2%VGND
x_PM_SKY130_FD_SC_LP__DLRBN_2%A_508_155# N_A_508_155#_M1025_s
+ N_A_508_155#_M1014_s N_A_508_155#_c_1204_n N_A_508_155#_c_1196_n
+ N_A_508_155#_c_1197_n PM_SKY130_FD_SC_LP__DLRBN_2%A_508_155#
x_PM_SKY130_FD_SC_LP__DLRBN_2%A_677_155# N_A_677_155#_M1019_d
+ N_A_677_155#_M1004_d N_A_677_155#_c_1222_n N_A_677_155#_c_1223_n
+ PM_SKY130_FD_SC_LP__DLRBN_2%A_677_155#
cc_1 VNB N_GATE_N_c_188_n 0.0189248f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.733
cc_2 VNB GATE_N 0.0207677f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_GATE_N_c_190_n 0.023095f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.415
cc_4 VNB N_GATE_N_c_191_n 0.0226348f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.25
cc_5 VNB N_A_113_144#_c_219_n 0.0176816f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.685
cc_6 VNB N_A_113_144#_M1012_g 0.00206566f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_113_144#_M1025_g 0.0356758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_113_144#_c_222_n 0.0613417f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.415
cc_9 VNB N_A_113_144#_c_223_n 0.0160057f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.665
cc_10 VNB N_A_113_144#_c_224_n 0.00247161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_113_144#_c_225_n 0.0016003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_113_144#_c_226_n 0.00330095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_113_144#_c_227_n 0.00285794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_D_c_322_n 0.0165959f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.437
cc_15 VNB N_D_M1008_g 0.00211356f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.92
cc_16 VNB D 0.00644055f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.685
cc_17 VNB N_D_c_325_n 0.0388017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_162_40#_c_356_n 0.166769f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.685
cc_19 VNB N_A_162_40#_M1019_g 0.0359906f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_20 VNB N_A_162_40#_c_358_n 0.0344702f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_21 VNB N_A_162_40#_c_359_n 0.00761329f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_22 VNB N_A_162_40#_M1015_g 0.0101787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_162_40#_c_361_n 0.00381661f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.415
cc_24 VNB N_A_162_40#_c_362_n 0.00616386f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.415
cc_25 VNB N_A_162_40#_c_363_n 0.00204064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_162_40#_c_364_n 0.00172415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_162_40#_c_365_n 0.0477742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_392_144#_c_437_n 0.0240126f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.685
cc_29 VNB N_A_392_144#_c_438_n 0.0126173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_392_144#_c_439_n 0.00691914f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.92
cc_31 VNB N_A_392_144#_M1018_g 0.034517f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_32 VNB N_A_392_144#_c_441_n 0.0175105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_392_144#_c_442_n 0.0141882f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.415
cc_34 VNB N_A_392_144#_c_443_n 0.0123222f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.415
cc_35 VNB N_A_392_144#_c_444_n 0.010845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_392_144#_c_445_n 0.0012924f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=2.035
cc_37 VNB N_A_392_144#_c_446_n 0.0178301f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=2.405
cc_38 VNB N_A_392_144#_c_447_n 0.0391115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_392_144#_c_448_n 0.00764162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_942_252#_M1005_g 0.00135402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_942_252#_M1004_g 0.038858f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_42 VNB N_A_942_252#_M1009_g 0.0207568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_942_252#_M1022_g 0.0229139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_942_252#_M1011_g 0.025904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_942_252#_c_532_n 0.0288362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_942_252#_c_533_n 0.0181656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_942_252#_c_534_n 0.00577872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_942_252#_c_535_n 0.0216058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_942_252#_c_536_n 0.0362362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_942_252#_c_537_n 0.0171717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_942_252#_c_538_n 0.00112395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_942_252#_c_539_n 0.0263479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_942_252#_c_540_n 0.00219983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_591_155#_c_674_n 0.0134123f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_55 VNB N_A_591_155#_c_675_n 0.00615187f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_56 VNB N_A_591_155#_M1027_g 0.0344547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_591_155#_c_677_n 0.00232228f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.415
cc_58 VNB N_A_591_155#_c_678_n 4.79822e-19 $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.25
cc_59 VNB N_A_591_155#_c_679_n 0.0112233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_591_155#_c_680_n 7.99442e-19 $X=-0.19 $Y=-0.245 $X2=0.277
+ $Y2=1.665
cc_61 VNB N_RESET_B_M1006_g 0.00327085f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.92
cc_62 VNB RESET_B 0.0149142f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.685
cc_63 VNB N_RESET_B_c_777_n 0.0285578f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.415
cc_64 VNB N_RESET_B_c_778_n 0.0170092f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.295
cc_65 VNB N_A_1555_367#_M1003_g 0.0246435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1555_367#_M1001_g 7.30661e-19 $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_67 VNB N_A_1555_367#_c_814_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1555_367#_M1013_g 0.0285202f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.415
cc_69 VNB N_A_1555_367#_M1023_g 0.0155486f $X=-0.19 $Y=-0.245 $X2=0.277
+ $Y2=1.295
cc_70 VNB N_A_1555_367#_c_817_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1555_367#_c_818_n 0.0147124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1555_367#_c_819_n 0.00297614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1555_367#_c_820_n 0.0366348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VPWR_c_877_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_Q_c_1038_n 0.00156739f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.92
cc_76 VNB N_Q_c_1039_n 0.00158703f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_77 VNB N_Q_N_c_1066_n 0.00827268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1084_n 0.0120573f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.25
cc_79 VNB N_VGND_c_1085_n 0.0437266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1086_n 0.0111135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1087_n 0.0104754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1088_n 0.00703937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1089_n 0.0245608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1090_n 0.0190926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1091_n 0.0111284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1092_n 0.0512481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1093_n 0.0295305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1094_n 0.0670976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1095_n 0.0443289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1096_n 0.0188039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1097_n 0.0218935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1098_n 0.0156559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1099_n 0.00370274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1100_n 0.00423165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1101_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1102_n 0.00596278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1103_n 0.00549216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1104_n 0.528129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_508_155#_c_1196_n 0.00284385f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_100 VNB N_A_508_155#_c_1197_n 0.00873717f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_101 VNB N_A_677_155#_c_1222_n 0.0219093f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=2.685
cc_102 VNB N_A_677_155#_c_1223_n 0.00704237f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_103 VPB N_GATE_N_c_188_n 0.00706052f $X=-0.19 $Y=1.655 $X2=0.407 $Y2=1.733
cc_104 VPB N_GATE_N_M1026_g 0.0435686f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.685
cc_105 VPB N_GATE_N_c_194_n 0.0235691f $X=-0.19 $Y=1.655 $X2=0.407 $Y2=1.92
cc_106 VPB GATE_N 0.0353714f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_107 VPB N_A_113_144#_M1012_g 0.0220005f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_108 VPB N_A_113_144#_c_229_n 0.0932647f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_109 VPB N_A_113_144#_M1025_g 0.0749852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_113_144#_c_231_n 0.0280035f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.415
cc_111 VPB N_A_113_144#_M1024_g 0.0418909f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_113_144#_c_233_n 0.00664245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_113_144#_c_225_n 0.0261092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_113_144#_c_235_n 0.00327581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_113_144#_c_236_n 0.0134787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_113_144#_c_237_n 0.0433305f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_D_M1008_g 0.0233251f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.92
cc_118 VPB D 0.0103536f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.685
cc_119 VPB N_A_162_40#_M1015_g 0.0178934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_162_40#_c_367_n 0.00309226f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.415
cc_121 VPB N_A_162_40#_c_368_n 0.0077371f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.295
cc_122 VPB N_A_162_40#_c_364_n 0.00219428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_392_144#_M1018_g 0.0209667f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_124 VPB N_A_392_144#_c_450_n 0.00622126f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.415
cc_125 VPB N_A_392_144#_c_451_n 0.00723881f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.295
cc_126 VPB N_A_392_144#_c_443_n 0.00320907f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.415
cc_127 VPB N_A_942_252#_M1005_g 0.0237261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_942_252#_M1000_g 0.0194868f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.415
cc_129 VPB N_A_942_252#_M1021_g 0.021358f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=2.035
cc_130 VPB N_A_942_252#_M1010_g 0.0257327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_942_252#_c_532_n 0.00262466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_942_252#_c_533_n 0.00557482f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_942_252#_c_534_n 3.79508e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_942_252#_c_548_n 0.00158822f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_942_252#_c_549_n 0.00107746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_942_252#_c_550_n 0.00145336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_942_252#_c_539_n 0.00850494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_591_155#_c_681_n 0.107634f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.685
cc_139 VPB N_A_591_155#_c_682_n 0.0769051f $X=-0.19 $Y=1.655 $X2=0.407 $Y2=1.92
cc_140 VPB N_A_591_155#_c_674_n 0.00794187f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_141 VPB N_A_591_155#_c_675_n 0.00398463f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_142 VPB N_A_591_155#_c_685_n 0.018472f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_591_155#_c_677_n 0.00204578f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.415
cc_144 VPB N_A_591_155#_c_678_n 0.00563737f $X=-0.19 $Y=1.655 $X2=0.407 $Y2=1.25
cc_145 VPB N_A_591_155#_c_688_n 0.0114342f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.295
cc_146 VPB N_A_591_155#_c_689_n 0.00539956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_591_155#_c_690_n 0.00387404f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=2.405
cc_148 VPB N_A_591_155#_c_691_n 0.0456364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_591_155#_c_692_n 0.00595279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_M1006_g 0.0186363f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.92
cc_151 VPB RESET_B 0.00129868f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.685
cc_152 VPB N_A_1555_367#_M1001_g 0.0235482f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_153 VPB N_A_1555_367#_M1023_g 0.0272177f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.295
cc_154 VPB N_A_1555_367#_c_823_n 0.00511683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_1555_367#_c_824_n 0.0150072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_1555_367#_c_825_n 0.00168299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_1555_367#_c_819_n 0.00144079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_878_n 0.0124576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_879_n 0.0212482f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.665
cc_160 VPB N_VPWR_c_880_n 0.0311624f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=2.405
cc_161 VPB N_VPWR_c_881_n 0.0197049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_882_n 0.00449364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_883_n 3.21238e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_884_n 0.0195267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_885_n 0.0275633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_886_n 0.0111025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_887_n 0.0653578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_888_n 0.0298299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_889_n 0.00477947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_890_n 0.0278421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_891_n 0.00459045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_892_n 0.0682706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_893_n 0.0150561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_894_n 0.0153449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_895_n 0.0238029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_896_n 0.0151073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_897_n 0.00583335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_898_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_899_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_900_n 0.00497525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_877_n 0.103989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_606_359#_c_1003_n 0.0122363f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.685
cc_183 VPB N_A_606_359#_c_1004_n 0.00257609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_606_359#_c_1005_n 0.0075249f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_185 VPB N_Q_c_1040_n 0.00116944f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_186 VPB N_Q_c_1039_n 0.00108064f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_187 VPB N_Q_N_c_1066_n 0.00425363f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 GATE_N N_A_113_144#_c_222_n 2.4546e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_189 N_GATE_N_c_190_n N_A_113_144#_c_222_n 0.0206348f $X=0.385 $Y=1.415 $X2=0
+ $Y2=0
cc_190 GATE_N N_A_113_144#_c_224_n 0.00301646f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_191 N_GATE_N_c_191_n N_A_113_144#_c_224_n 0.00699015f $X=0.407 $Y=1.25 $X2=0
+ $Y2=0
cc_192 N_GATE_N_c_188_n N_A_113_144#_c_225_n 0.0191448f $X=0.407 $Y=1.733 $X2=0
+ $Y2=0
cc_193 GATE_N N_A_113_144#_c_225_n 0.0663458f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_194 N_GATE_N_M1026_g N_A_113_144#_c_235_n 8.33328e-19 $X=0.52 $Y=2.685 $X2=0
+ $Y2=0
cc_195 N_GATE_N_c_191_n N_A_113_144#_c_226_n 4.43964e-19 $X=0.407 $Y=1.25 $X2=0
+ $Y2=0
cc_196 GATE_N N_A_113_144#_c_227_n 0.0268194f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_197 N_GATE_N_c_190_n N_A_113_144#_c_227_n 0.00248201f $X=0.385 $Y=1.415 $X2=0
+ $Y2=0
cc_198 N_GATE_N_M1026_g N_A_113_144#_c_237_n 0.00314792f $X=0.52 $Y=2.685 $X2=0
+ $Y2=0
cc_199 N_GATE_N_c_191_n N_A_162_40#_c_362_n 0.0025442f $X=0.407 $Y=1.25 $X2=0
+ $Y2=0
cc_200 GATE_N N_VPWR_M1026_s 0.00285862f $X=0.155 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_201 N_GATE_N_M1026_g N_VPWR_c_879_n 0.00987068f $X=0.52 $Y=2.685 $X2=0 $Y2=0
cc_202 GATE_N N_VPWR_c_879_n 0.0238082f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_203 N_GATE_N_M1026_g N_VPWR_c_888_n 0.00414769f $X=0.52 $Y=2.685 $X2=0 $Y2=0
cc_204 N_GATE_N_M1026_g N_VPWR_c_877_n 0.00826848f $X=0.52 $Y=2.685 $X2=0 $Y2=0
cc_205 GATE_N N_VPWR_c_877_n 0.00335395f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_206 GATE_N N_VGND_c_1085_n 0.0274351f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_207 N_GATE_N_c_190_n N_VGND_c_1085_n 0.00121027f $X=0.385 $Y=1.415 $X2=0
+ $Y2=0
cc_208 N_GATE_N_c_191_n N_VGND_c_1085_n 0.00952974f $X=0.407 $Y=1.25 $X2=0 $Y2=0
cc_209 N_GATE_N_c_191_n N_VGND_c_1093_n 0.00306407f $X=0.407 $Y=1.25 $X2=0 $Y2=0
cc_210 N_GATE_N_c_191_n N_VGND_c_1104_n 0.00372921f $X=0.407 $Y=1.25 $X2=0 $Y2=0
cc_211 N_A_113_144#_c_219_n N_D_c_322_n 0.0120579f $X=1.455 $Y=1.25 $X2=-0.19
+ $Y2=-0.245
cc_212 N_A_113_144#_M1012_g N_D_M1008_g 0.0194915f $X=1.495 $Y=2.115 $X2=0 $Y2=0
cc_213 N_A_113_144#_c_229_n N_D_M1008_g 0.00936846f $X=2.805 $Y=2.88 $X2=0 $Y2=0
cc_214 N_A_113_144#_c_219_n D 3.0994e-19 $X=1.455 $Y=1.25 $X2=0 $Y2=0
cc_215 N_A_113_144#_c_223_n D 0.00479337f $X=1.475 $Y=1.415 $X2=0 $Y2=0
cc_216 N_A_113_144#_M1025_g N_D_c_325_n 0.0110969f $X=2.88 $Y=0.985 $X2=0 $Y2=0
cc_217 N_A_113_144#_c_223_n N_D_c_325_n 0.021559f $X=1.475 $Y=1.415 $X2=0 $Y2=0
cc_218 N_A_113_144#_c_219_n N_A_162_40#_c_356_n 0.00908082f $X=1.455 $Y=1.25
+ $X2=0 $Y2=0
cc_219 N_A_113_144#_M1025_g N_A_162_40#_c_356_n 0.00636915f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_220 N_A_113_144#_M1025_g N_A_162_40#_M1019_g 0.0222092f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_221 N_A_113_144#_M1024_g N_A_162_40#_c_359_n 0.0111303f $X=3.37 $Y=2.005
+ $X2=0 $Y2=0
cc_222 N_A_113_144#_M1024_g N_A_162_40#_M1015_g 0.0224099f $X=3.37 $Y=2.005
+ $X2=0 $Y2=0
cc_223 N_A_113_144#_c_226_n N_A_162_40#_c_361_n 4.78424e-19 $X=0.705 $Y=0.865
+ $X2=0 $Y2=0
cc_224 N_A_113_144#_c_219_n N_A_162_40#_c_362_n 0.00636363f $X=1.455 $Y=1.25
+ $X2=0 $Y2=0
cc_225 N_A_113_144#_c_226_n N_A_162_40#_c_362_n 0.0112176f $X=0.705 $Y=0.865
+ $X2=0 $Y2=0
cc_226 N_A_113_144#_c_222_n N_A_162_40#_c_367_n 0.0051022f $X=1.38 $Y=1.415
+ $X2=0 $Y2=0
cc_227 N_A_113_144#_c_225_n N_A_162_40#_c_367_n 0.0459993f $X=0.735 $Y=2.52
+ $X2=0 $Y2=0
cc_228 N_A_113_144#_c_236_n N_A_162_40#_c_368_n 0.0150456f $X=1.355 $Y=2.94
+ $X2=0 $Y2=0
cc_229 N_A_113_144#_c_237_n N_A_162_40#_c_368_n 0.00453155f $X=1.52 $Y=2.94
+ $X2=0 $Y2=0
cc_230 N_A_113_144#_c_219_n N_A_162_40#_c_363_n 0.00198593f $X=1.455 $Y=1.25
+ $X2=0 $Y2=0
cc_231 N_A_113_144#_c_222_n N_A_162_40#_c_363_n 0.00621555f $X=1.38 $Y=1.415
+ $X2=0 $Y2=0
cc_232 N_A_113_144#_c_224_n N_A_162_40#_c_363_n 0.0112176f $X=0.73 $Y=1.25 $X2=0
+ $Y2=0
cc_233 N_A_113_144#_c_219_n N_A_162_40#_c_364_n 0.00490768f $X=1.455 $Y=1.25
+ $X2=0 $Y2=0
cc_234 N_A_113_144#_M1012_g N_A_162_40#_c_364_n 0.00620632f $X=1.495 $Y=2.115
+ $X2=0 $Y2=0
cc_235 N_A_113_144#_c_222_n N_A_162_40#_c_364_n 0.0159607f $X=1.38 $Y=1.415
+ $X2=0 $Y2=0
cc_236 N_A_113_144#_c_223_n N_A_162_40#_c_364_n 0.0042497f $X=1.475 $Y=1.415
+ $X2=0 $Y2=0
cc_237 N_A_113_144#_c_224_n N_A_162_40#_c_364_n 0.00486831f $X=0.73 $Y=1.25
+ $X2=0 $Y2=0
cc_238 N_A_113_144#_c_225_n N_A_162_40#_c_364_n 0.00705545f $X=0.735 $Y=2.52
+ $X2=0 $Y2=0
cc_239 N_A_113_144#_c_227_n N_A_162_40#_c_364_n 0.0229044f $X=0.97 $Y=1.415
+ $X2=0 $Y2=0
cc_240 N_A_113_144#_c_222_n N_A_162_40#_c_365_n 0.00677113f $X=1.38 $Y=1.415
+ $X2=0 $Y2=0
cc_241 N_A_113_144#_M1025_g N_A_392_144#_c_450_n 0.00110417f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_242 N_A_113_144#_c_229_n N_A_392_144#_c_451_n 0.010244f $X=2.805 $Y=2.88
+ $X2=0 $Y2=0
cc_243 N_A_113_144#_M1025_g N_A_392_144#_c_451_n 0.00130391f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_244 N_A_113_144#_M1025_g N_A_392_144#_c_443_n 0.00407982f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_245 N_A_113_144#_M1025_g N_A_392_144#_c_444_n 2.20914e-19 $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_246 N_A_113_144#_M1025_g N_A_392_144#_c_446_n 4.49332e-19 $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_247 N_A_113_144#_M1025_g N_A_392_144#_c_448_n 3.91561e-19 $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_248 N_A_113_144#_M1025_g N_A_591_155#_c_678_n 0.0222397f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_249 N_A_113_144#_M1024_g N_A_591_155#_c_678_n 0.00116715f $X=3.37 $Y=2.005
+ $X2=0 $Y2=0
cc_250 N_A_113_144#_M1025_g N_A_591_155#_c_688_n 0.0126682f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_251 N_A_113_144#_c_231_n N_A_591_155#_c_688_n 0.00377811f $X=3.295 $Y=2.88
+ $X2=0 $Y2=0
cc_252 N_A_113_144#_M1024_g N_A_591_155#_c_688_n 0.019692f $X=3.37 $Y=2.005
+ $X2=0 $Y2=0
cc_253 N_A_113_144#_c_229_n N_A_591_155#_c_689_n 0.00262328f $X=2.805 $Y=2.88
+ $X2=0 $Y2=0
cc_254 N_A_113_144#_M1025_g N_A_591_155#_c_689_n 0.00735057f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_255 N_A_113_144#_M1025_g N_A_591_155#_c_679_n 0.0152033f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_256 N_A_113_144#_M1025_g N_A_591_155#_c_680_n 0.0105248f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_257 N_A_113_144#_M1024_g N_A_591_155#_c_690_n 0.0067212f $X=3.37 $Y=2.005
+ $X2=0 $Y2=0
cc_258 N_A_113_144#_M1024_g N_A_591_155#_c_691_n 0.00727191f $X=3.37 $Y=2.005
+ $X2=0 $Y2=0
cc_259 N_A_113_144#_M1024_g N_A_591_155#_c_692_n 0.00254892f $X=3.37 $Y=2.005
+ $X2=0 $Y2=0
cc_260 N_A_113_144#_c_235_n N_VPWR_c_879_n 0.0145269f $X=0.9 $Y=2.925 $X2=0
+ $Y2=0
cc_261 N_A_113_144#_M1012_g N_VPWR_c_880_n 0.00809596f $X=1.495 $Y=2.115 $X2=0
+ $Y2=0
cc_262 N_A_113_144#_c_229_n N_VPWR_c_880_n 0.0239885f $X=2.805 $Y=2.88 $X2=0
+ $Y2=0
cc_263 N_A_113_144#_c_236_n N_VPWR_c_880_n 0.023903f $X=1.355 $Y=2.94 $X2=0
+ $Y2=0
cc_264 N_A_113_144#_c_237_n N_VPWR_c_880_n 0.00208705f $X=1.52 $Y=2.94 $X2=0
+ $Y2=0
cc_265 N_A_113_144#_c_229_n N_VPWR_c_888_n 0.00437818f $X=2.805 $Y=2.88 $X2=0
+ $Y2=0
cc_266 N_A_113_144#_c_235_n N_VPWR_c_888_n 0.0185661f $X=0.9 $Y=2.925 $X2=0
+ $Y2=0
cc_267 N_A_113_144#_c_236_n N_VPWR_c_888_n 0.0404966f $X=1.355 $Y=2.94 $X2=0
+ $Y2=0
cc_268 N_A_113_144#_c_237_n N_VPWR_c_888_n 0.00577541f $X=1.52 $Y=2.94 $X2=0
+ $Y2=0
cc_269 N_A_113_144#_c_229_n N_VPWR_c_892_n 0.0367894f $X=2.805 $Y=2.88 $X2=0
+ $Y2=0
cc_270 N_A_113_144#_c_229_n N_VPWR_c_877_n 0.0480995f $X=2.805 $Y=2.88 $X2=0
+ $Y2=0
cc_271 N_A_113_144#_c_235_n N_VPWR_c_877_n 0.0100976f $X=0.9 $Y=2.925 $X2=0
+ $Y2=0
cc_272 N_A_113_144#_c_236_n N_VPWR_c_877_n 0.0220946f $X=1.355 $Y=2.94 $X2=0
+ $Y2=0
cc_273 N_A_113_144#_c_237_n N_VPWR_c_877_n 0.00800665f $X=1.52 $Y=2.94 $X2=0
+ $Y2=0
cc_274 N_A_113_144#_M1024_g N_A_606_359#_c_1003_n 0.00916504f $X=3.37 $Y=2.005
+ $X2=0 $Y2=0
cc_275 N_A_113_144#_M1025_g N_A_606_359#_c_1004_n 0.00258901f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_276 N_A_113_144#_M1024_g N_A_606_359#_c_1004_n 0.00507882f $X=3.37 $Y=2.005
+ $X2=0 $Y2=0
cc_277 N_A_113_144#_c_224_n N_VGND_c_1085_n 6.21674e-19 $X=0.73 $Y=1.25 $X2=0
+ $Y2=0
cc_278 N_A_113_144#_c_226_n N_VGND_c_1085_n 0.0131206f $X=0.705 $Y=0.865 $X2=0
+ $Y2=0
cc_279 N_A_113_144#_c_219_n N_VGND_c_1086_n 9.47161e-19 $X=1.455 $Y=1.25 $X2=0
+ $Y2=0
cc_280 N_A_113_144#_c_226_n N_VGND_c_1093_n 0.00346289f $X=0.705 $Y=0.865 $X2=0
+ $Y2=0
cc_281 N_A_113_144#_c_219_n N_VGND_c_1104_n 7.07383e-19 $X=1.455 $Y=1.25 $X2=0
+ $Y2=0
cc_282 N_A_113_144#_c_226_n N_VGND_c_1104_n 0.00570654f $X=0.705 $Y=0.865 $X2=0
+ $Y2=0
cc_283 N_A_113_144#_M1025_g N_A_508_155#_c_1197_n 0.011102f $X=2.88 $Y=0.985
+ $X2=0 $Y2=0
cc_284 N_D_c_322_n N_A_162_40#_c_356_n 0.00924127f $X=1.885 $Y=1.25 $X2=0 $Y2=0
cc_285 N_D_c_322_n N_A_162_40#_c_362_n 8.89533e-19 $X=1.885 $Y=1.25 $X2=0 $Y2=0
cc_286 D N_A_162_40#_c_364_n 0.0427051f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_287 N_D_c_325_n N_A_162_40#_c_364_n 2.25016e-19 $X=2.08 $Y=1.415 $X2=0 $Y2=0
cc_288 N_D_M1008_g N_A_392_144#_c_450_n 0.00349749f $X=2.08 $Y=2.115 $X2=0 $Y2=0
cc_289 N_D_M1008_g N_A_392_144#_c_451_n 0.00442198f $X=2.08 $Y=2.115 $X2=0 $Y2=0
cc_290 N_D_c_322_n N_A_392_144#_c_443_n 0.00519907f $X=1.885 $Y=1.25 $X2=0 $Y2=0
cc_291 D N_A_392_144#_c_443_n 0.0419097f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_292 N_D_c_325_n N_A_392_144#_c_443_n 0.0070568f $X=2.08 $Y=1.415 $X2=0 $Y2=0
cc_293 N_D_c_322_n N_A_392_144#_c_444_n 0.00216486f $X=1.885 $Y=1.25 $X2=0 $Y2=0
cc_294 N_D_c_322_n N_A_392_144#_c_448_n 4.53275e-19 $X=1.885 $Y=1.25 $X2=0 $Y2=0
cc_295 D N_A_392_144#_c_448_n 0.00336958f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_296 N_D_c_325_n N_A_392_144#_c_448_n 0.00567191f $X=2.08 $Y=1.415 $X2=0 $Y2=0
cc_297 N_D_M1008_g N_A_591_155#_c_689_n 0.00273699f $X=2.08 $Y=2.115 $X2=0 $Y2=0
cc_298 N_D_M1008_g N_VPWR_c_880_n 0.00814833f $X=2.08 $Y=2.115 $X2=0 $Y2=0
cc_299 D N_VPWR_c_880_n 0.0224027f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_300 N_D_c_325_n N_VPWR_c_880_n 8.34534e-19 $X=2.08 $Y=1.415 $X2=0 $Y2=0
cc_301 N_D_c_322_n N_VGND_c_1086_n 0.00144303f $X=1.885 $Y=1.25 $X2=0 $Y2=0
cc_302 D N_VGND_c_1086_n 0.0173485f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_303 N_D_c_322_n N_VGND_c_1104_n 8.46057e-19 $X=1.885 $Y=1.25 $X2=0 $Y2=0
cc_304 N_D_c_322_n N_A_508_155#_c_1196_n 2.80528e-19 $X=1.885 $Y=1.25 $X2=0
+ $Y2=0
cc_305 N_A_162_40#_M1019_g N_A_392_144#_c_437_n 0.0169613f $X=3.31 $Y=0.985
+ $X2=0 $Y2=0
cc_306 N_A_162_40#_c_358_n N_A_392_144#_c_439_n 0.010157f $X=3.82 $Y=1.38 $X2=0
+ $Y2=0
cc_307 N_A_162_40#_c_358_n N_A_392_144#_M1018_g 0.0803638f $X=3.82 $Y=1.38 $X2=0
+ $Y2=0
cc_308 N_A_162_40#_c_356_n N_A_392_144#_c_445_n 0.00831118f $X=3.235 $Y=0.275
+ $X2=0 $Y2=0
cc_309 N_A_162_40#_c_356_n N_A_392_144#_c_446_n 0.0283225f $X=3.235 $Y=0.275
+ $X2=0 $Y2=0
cc_310 N_A_162_40#_M1019_g N_A_392_144#_c_446_n 0.00656387f $X=3.31 $Y=0.985
+ $X2=0 $Y2=0
cc_311 N_A_162_40#_c_356_n N_A_392_144#_c_447_n 0.0182746f $X=3.235 $Y=0.275
+ $X2=0 $Y2=0
cc_312 N_A_162_40#_c_356_n N_A_392_144#_c_448_n 0.00534942f $X=3.235 $Y=0.275
+ $X2=0 $Y2=0
cc_313 N_A_162_40#_c_359_n N_A_591_155#_c_679_n 0.00239126f $X=3.385 $Y=1.38
+ $X2=0 $Y2=0
cc_314 N_A_162_40#_M1015_g N_A_591_155#_c_679_n 0.00366911f $X=3.895 $Y=2.115
+ $X2=0 $Y2=0
cc_315 N_A_162_40#_M1019_g N_A_591_155#_c_680_n 0.0101054f $X=3.31 $Y=0.985
+ $X2=0 $Y2=0
cc_316 N_A_162_40#_c_359_n N_A_591_155#_c_680_n 0.00751231f $X=3.385 $Y=1.38
+ $X2=0 $Y2=0
cc_317 N_A_162_40#_M1015_g N_A_591_155#_c_691_n 0.00977216f $X=3.895 $Y=2.115
+ $X2=0 $Y2=0
cc_318 N_A_162_40#_M1015_g N_A_591_155#_c_692_n 0.0148953f $X=3.895 $Y=2.115
+ $X2=0 $Y2=0
cc_319 N_A_162_40#_c_368_n N_VPWR_c_880_n 0.0140782f $X=1.28 $Y=1.94 $X2=0 $Y2=0
cc_320 N_A_162_40#_M1015_g N_VPWR_c_881_n 6.75621e-19 $X=3.895 $Y=2.115 $X2=0
+ $Y2=0
cc_321 N_A_162_40#_c_358_n N_A_606_359#_c_1003_n 0.00730971f $X=3.82 $Y=1.38
+ $X2=0 $Y2=0
cc_322 N_A_162_40#_c_359_n N_A_606_359#_c_1003_n 6.94889e-19 $X=3.385 $Y=1.38
+ $X2=0 $Y2=0
cc_323 N_A_162_40#_M1015_g N_A_606_359#_c_1003_n 0.0126513f $X=3.895 $Y=2.115
+ $X2=0 $Y2=0
cc_324 N_A_162_40#_c_359_n N_A_606_359#_c_1004_n 0.00160432f $X=3.385 $Y=1.38
+ $X2=0 $Y2=0
cc_325 N_A_162_40#_M1015_g N_A_606_359#_c_1004_n 6.63216e-19 $X=3.895 $Y=2.115
+ $X2=0 $Y2=0
cc_326 N_A_162_40#_c_361_n N_VGND_c_1085_n 0.00779361f $X=1.24 $Y=0.45 $X2=0
+ $Y2=0
cc_327 N_A_162_40#_c_362_n N_VGND_c_1085_n 0.0075246f $X=1.24 $Y=0.915 $X2=0
+ $Y2=0
cc_328 N_A_162_40#_c_365_n N_VGND_c_1085_n 0.00514483f $X=0.975 $Y=0.275 $X2=0
+ $Y2=0
cc_329 N_A_162_40#_c_356_n N_VGND_c_1086_n 0.0199466f $X=3.235 $Y=0.275 $X2=0
+ $Y2=0
cc_330 N_A_162_40#_c_361_n N_VGND_c_1086_n 0.0137118f $X=1.24 $Y=0.45 $X2=0
+ $Y2=0
cc_331 N_A_162_40#_c_362_n N_VGND_c_1086_n 0.0332053f $X=1.24 $Y=0.915 $X2=0
+ $Y2=0
cc_332 N_A_162_40#_c_365_n N_VGND_c_1086_n 7.11833e-19 $X=0.975 $Y=0.275 $X2=0
+ $Y2=0
cc_333 N_A_162_40#_c_361_n N_VGND_c_1093_n 0.0314699f $X=1.24 $Y=0.45 $X2=0
+ $Y2=0
cc_334 N_A_162_40#_c_365_n N_VGND_c_1093_n 0.0157158f $X=0.975 $Y=0.275 $X2=0
+ $Y2=0
cc_335 N_A_162_40#_c_356_n N_VGND_c_1094_n 0.0303994f $X=3.235 $Y=0.275 $X2=0
+ $Y2=0
cc_336 N_A_162_40#_c_356_n N_VGND_c_1104_n 0.0533292f $X=3.235 $Y=0.275 $X2=0
+ $Y2=0
cc_337 N_A_162_40#_c_361_n N_VGND_c_1104_n 0.0192531f $X=1.24 $Y=0.45 $X2=0
+ $Y2=0
cc_338 N_A_162_40#_c_365_n N_VGND_c_1104_n 0.00853508f $X=0.975 $Y=0.275 $X2=0
+ $Y2=0
cc_339 N_A_162_40#_c_356_n N_A_508_155#_c_1196_n 0.0012902f $X=3.235 $Y=0.275
+ $X2=0 $Y2=0
cc_340 N_A_162_40#_c_356_n N_A_508_155#_c_1197_n 0.00220413f $X=3.235 $Y=0.275
+ $X2=0 $Y2=0
cc_341 N_A_162_40#_M1019_g N_A_508_155#_c_1197_n 0.0155002f $X=3.31 $Y=0.985
+ $X2=0 $Y2=0
cc_342 N_A_162_40#_c_358_n N_A_508_155#_c_1197_n 0.00107033f $X=3.82 $Y=1.38
+ $X2=0 $Y2=0
cc_343 N_A_162_40#_c_358_n N_A_677_155#_c_1222_n 0.0107114f $X=3.82 $Y=1.38
+ $X2=0 $Y2=0
cc_344 N_A_392_144#_M1018_g N_A_942_252#_M1004_g 0.00505872f $X=4.255 $Y=2.115
+ $X2=0 $Y2=0
cc_345 N_A_392_144#_c_441_n N_A_942_252#_M1004_g 0.0179314f $X=4.425 $Y=0.935
+ $X2=0 $Y2=0
cc_346 N_A_392_144#_M1018_g N_A_942_252#_c_535_n 0.00160383f $X=4.255 $Y=2.115
+ $X2=0 $Y2=0
cc_347 N_A_392_144#_M1018_g N_A_942_252#_c_536_n 0.0294976f $X=4.255 $Y=2.115
+ $X2=0 $Y2=0
cc_348 N_A_392_144#_M1018_g N_A_591_155#_c_681_n 0.00548134f $X=4.255 $Y=2.115
+ $X2=0 $Y2=0
cc_349 N_A_392_144#_c_450_n N_A_591_155#_c_678_n 0.0192181f $X=2.295 $Y=2.085
+ $X2=0 $Y2=0
cc_350 N_A_392_144#_c_451_n N_A_591_155#_c_678_n 0.0124027f $X=2.295 $Y=2.28
+ $X2=0 $Y2=0
cc_351 N_A_392_144#_c_443_n N_A_591_155#_c_678_n 0.00875882f $X=2.29 $Y=1.775
+ $X2=0 $Y2=0
cc_352 N_A_392_144#_c_451_n N_A_591_155#_c_689_n 0.011112f $X=2.295 $Y=2.28
+ $X2=0 $Y2=0
cc_353 N_A_392_144#_c_443_n N_A_591_155#_c_679_n 0.00902706f $X=2.29 $Y=1.775
+ $X2=0 $Y2=0
cc_354 N_A_392_144#_c_443_n N_A_591_155#_c_680_n 0.00855184f $X=2.29 $Y=1.775
+ $X2=0 $Y2=0
cc_355 N_A_392_144#_M1018_g N_A_591_155#_c_692_n 0.00191733f $X=4.255 $Y=2.115
+ $X2=0 $Y2=0
cc_356 N_A_392_144#_c_450_n N_VPWR_c_880_n 0.0115604f $X=2.295 $Y=2.085 $X2=0
+ $Y2=0
cc_357 N_A_392_144#_c_451_n N_VPWR_c_880_n 0.0250892f $X=2.295 $Y=2.28 $X2=0
+ $Y2=0
cc_358 N_A_392_144#_M1018_g N_VPWR_c_881_n 0.0085938f $X=4.255 $Y=2.115 $X2=0
+ $Y2=0
cc_359 N_A_392_144#_M1018_g N_VPWR_c_877_n 7.42461e-19 $X=4.255 $Y=2.115 $X2=0
+ $Y2=0
cc_360 N_A_392_144#_c_438_n N_A_606_359#_c_1003_n 9.43288e-19 $X=4.18 $Y=1.01
+ $X2=0 $Y2=0
cc_361 N_A_392_144#_M1018_g N_A_606_359#_c_1003_n 0.0163621f $X=4.255 $Y=2.115
+ $X2=0 $Y2=0
cc_362 N_A_392_144#_c_442_n N_A_606_359#_c_1003_n 7.57803e-19 $X=4.425 $Y=1.01
+ $X2=0 $Y2=0
cc_363 N_A_392_144#_M1018_g N_A_606_359#_c_1005_n 7.18812e-19 $X=4.255 $Y=2.115
+ $X2=0 $Y2=0
cc_364 N_A_392_144#_c_444_n N_VGND_c_1086_n 0.0105305f $X=2.295 $Y=0.7 $X2=0
+ $Y2=0
cc_365 N_A_392_144#_c_445_n N_VGND_c_1086_n 0.00797368f $X=2.38 $Y=0.35 $X2=0
+ $Y2=0
cc_366 N_A_392_144#_c_448_n N_VGND_c_1086_n 0.00148629f $X=2.295 $Y=0.87 $X2=0
+ $Y2=0
cc_367 N_A_392_144#_c_441_n N_VGND_c_1087_n 0.0016771f $X=4.425 $Y=0.935 $X2=0
+ $Y2=0
cc_368 N_A_392_144#_c_446_n N_VGND_c_1087_n 0.00523301f $X=3.79 $Y=0.35 $X2=0
+ $Y2=0
cc_369 N_A_392_144#_c_447_n N_VGND_c_1087_n 0.00126845f $X=3.79 $Y=0.35 $X2=0
+ $Y2=0
cc_370 N_A_392_144#_c_441_n N_VGND_c_1094_n 0.00530499f $X=4.425 $Y=0.935 $X2=0
+ $Y2=0
cc_371 N_A_392_144#_c_445_n N_VGND_c_1094_n 0.0112461f $X=2.38 $Y=0.35 $X2=0
+ $Y2=0
cc_372 N_A_392_144#_c_446_n N_VGND_c_1094_n 0.0982432f $X=3.79 $Y=0.35 $X2=0
+ $Y2=0
cc_373 N_A_392_144#_c_447_n N_VGND_c_1094_n 0.00647615f $X=3.79 $Y=0.35 $X2=0
+ $Y2=0
cc_374 N_A_392_144#_c_448_n N_VGND_c_1094_n 0.00412524f $X=2.295 $Y=0.87 $X2=0
+ $Y2=0
cc_375 N_A_392_144#_c_441_n N_VGND_c_1104_n 0.00534666f $X=4.425 $Y=0.935 $X2=0
+ $Y2=0
cc_376 N_A_392_144#_c_445_n N_VGND_c_1104_n 0.00576194f $X=2.38 $Y=0.35 $X2=0
+ $Y2=0
cc_377 N_A_392_144#_c_446_n N_VGND_c_1104_n 0.053241f $X=3.79 $Y=0.35 $X2=0
+ $Y2=0
cc_378 N_A_392_144#_c_447_n N_VGND_c_1104_n 0.00961399f $X=3.79 $Y=0.35 $X2=0
+ $Y2=0
cc_379 N_A_392_144#_c_448_n N_VGND_c_1104_n 0.00591505f $X=2.295 $Y=0.87 $X2=0
+ $Y2=0
cc_380 N_A_392_144#_c_443_n N_A_508_155#_c_1204_n 0.00830095f $X=2.29 $Y=1.775
+ $X2=0 $Y2=0
cc_381 N_A_392_144#_c_448_n N_A_508_155#_c_1204_n 0.0197174f $X=2.295 $Y=0.87
+ $X2=0 $Y2=0
cc_382 N_A_392_144#_c_444_n N_A_508_155#_c_1196_n 0.00717904f $X=2.295 $Y=0.7
+ $X2=0 $Y2=0
cc_383 N_A_392_144#_c_446_n N_A_508_155#_c_1196_n 0.0164903f $X=3.79 $Y=0.35
+ $X2=0 $Y2=0
cc_384 N_A_392_144#_c_448_n N_A_508_155#_c_1196_n 0.00845692f $X=2.295 $Y=0.87
+ $X2=0 $Y2=0
cc_385 N_A_392_144#_c_437_n N_A_508_155#_c_1197_n 0.012095f $X=3.88 $Y=0.935
+ $X2=0 $Y2=0
cc_386 N_A_392_144#_c_438_n N_A_508_155#_c_1197_n 0.00484381f $X=4.18 $Y=1.01
+ $X2=0 $Y2=0
cc_387 N_A_392_144#_c_441_n N_A_508_155#_c_1197_n 0.00285282f $X=4.425 $Y=0.935
+ $X2=0 $Y2=0
cc_388 N_A_392_144#_c_446_n N_A_508_155#_c_1197_n 0.0832348f $X=3.79 $Y=0.35
+ $X2=0 $Y2=0
cc_389 N_A_392_144#_c_447_n N_A_508_155#_c_1197_n 0.0043898f $X=3.79 $Y=0.35
+ $X2=0 $Y2=0
cc_390 N_A_392_144#_c_438_n N_A_677_155#_c_1222_n 0.00778645f $X=4.18 $Y=1.01
+ $X2=0 $Y2=0
cc_391 N_A_392_144#_c_439_n N_A_677_155#_c_1222_n 0.00598892f $X=3.955 $Y=1.01
+ $X2=0 $Y2=0
cc_392 N_A_392_144#_M1018_g N_A_677_155#_c_1222_n 0.00790699f $X=4.255 $Y=2.115
+ $X2=0 $Y2=0
cc_393 N_A_392_144#_c_442_n N_A_677_155#_c_1222_n 0.0152863f $X=4.425 $Y=1.01
+ $X2=0 $Y2=0
cc_394 N_A_942_252#_M1005_g N_A_591_155#_c_681_n 0.00422034f $X=4.785 $Y=2.005
+ $X2=0 $Y2=0
cc_395 N_A_942_252#_c_548_n N_A_591_155#_c_682_n 0.00820251f $X=5.65 $Y=2.325
+ $X2=0 $Y2=0
cc_396 N_A_942_252#_c_558_p N_A_591_155#_c_682_n 0.00499476f $X=5.735 $Y=2.41
+ $X2=0 $Y2=0
cc_397 N_A_942_252#_c_535_n N_A_591_155#_c_674_n 0.00227287f $X=5.465 $Y=1.465
+ $X2=0 $Y2=0
cc_398 N_A_942_252#_c_548_n N_A_591_155#_c_674_n 0.0109631f $X=5.65 $Y=2.325
+ $X2=0 $Y2=0
cc_399 N_A_942_252#_c_540_n N_A_591_155#_c_674_n 0.0126738f $X=5.6 $Y=1.465
+ $X2=0 $Y2=0
cc_400 N_A_942_252#_M1005_g N_A_591_155#_c_675_n 0.0159925f $X=4.785 $Y=2.005
+ $X2=0 $Y2=0
cc_401 N_A_942_252#_c_535_n N_A_591_155#_c_675_n 0.0107139f $X=5.465 $Y=1.465
+ $X2=0 $Y2=0
cc_402 N_A_942_252#_c_536_n N_A_591_155#_c_675_n 8.27877e-19 $X=4.875 $Y=1.425
+ $X2=0 $Y2=0
cc_403 N_A_942_252#_c_537_n N_A_591_155#_M1027_g 0.0092467f $X=5.63 $Y=0.445
+ $X2=0 $Y2=0
cc_404 N_A_942_252#_c_540_n N_A_591_155#_M1027_g 0.00594255f $X=5.6 $Y=1.465
+ $X2=0 $Y2=0
cc_405 N_A_942_252#_c_548_n N_A_591_155#_c_685_n 0.00344266f $X=5.65 $Y=2.325
+ $X2=0 $Y2=0
cc_406 N_A_942_252#_c_568_p N_A_591_155#_c_685_n 0.0139911f $X=5.935 $Y=2.41
+ $X2=0 $Y2=0
cc_407 N_A_942_252#_c_532_n N_RESET_B_M1006_g 0.0465764f $X=7.25 $Y=1.49 $X2=0
+ $Y2=0
cc_408 N_A_942_252#_c_549_n N_RESET_B_M1006_g 0.0100497f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_409 N_A_942_252#_M1020_d RESET_B 0.001837f $X=5.92 $Y=1.835 $X2=0 $Y2=0
cc_410 N_A_942_252#_M1009_g RESET_B 0.00707132f $X=6.745 $Y=0.72 $X2=0 $Y2=0
cc_411 N_A_942_252#_c_537_n RESET_B 0.00905268f $X=5.63 $Y=0.445 $X2=0 $Y2=0
cc_412 N_A_942_252#_c_548_n RESET_B 0.029912f $X=5.65 $Y=2.325 $X2=0 $Y2=0
cc_413 N_A_942_252#_c_568_p RESET_B 2.7065e-19 $X=5.935 $Y=2.41 $X2=0 $Y2=0
cc_414 N_A_942_252#_c_549_n RESET_B 0.0281521f $X=7.225 $Y=2.41 $X2=0 $Y2=0
cc_415 N_A_942_252#_c_540_n RESET_B 0.0236896f $X=5.6 $Y=1.465 $X2=0 $Y2=0
cc_416 N_A_942_252#_c_578_p RESET_B 0.0149669f $X=6.06 $Y=2.49 $X2=0 $Y2=0
cc_417 N_A_942_252#_M1009_g N_RESET_B_c_777_n 0.021023f $X=6.745 $Y=0.72 $X2=0
+ $Y2=0
cc_418 N_A_942_252#_M1009_g N_RESET_B_c_778_n 0.0180515f $X=6.745 $Y=0.72 $X2=0
+ $Y2=0
cc_419 N_A_942_252#_c_539_n N_A_1555_367#_M1001_g 3.28042e-19 $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_420 N_A_942_252#_M1021_g N_A_1555_367#_c_823_n 3.86425e-19 $X=7.175 $Y=2.465
+ $X2=0 $Y2=0
cc_421 N_A_942_252#_M1010_g N_A_1555_367#_c_823_n 0.00648025f $X=7.7 $Y=2.155
+ $X2=0 $Y2=0
cc_422 N_A_942_252#_c_549_n N_A_1555_367#_c_823_n 0.00626904f $X=7.225 $Y=2.41
+ $X2=0 $Y2=0
cc_423 N_A_942_252#_M1011_g N_A_1555_367#_c_818_n 0.0037909f $X=7.715 $Y=0.93
+ $X2=0 $Y2=0
cc_424 N_A_942_252#_c_538_n N_A_1555_367#_c_818_n 0.0172107f $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_425 N_A_942_252#_c_539_n N_A_1555_367#_c_818_n 0.00813965f $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_426 N_A_942_252#_c_538_n N_A_1555_367#_c_824_n 0.00921278f $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_427 N_A_942_252#_c_539_n N_A_1555_367#_c_824_n 0.00330352f $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_428 N_A_942_252#_M1010_g N_A_1555_367#_c_825_n 0.00403483f $X=7.7 $Y=2.155
+ $X2=0 $Y2=0
cc_429 N_A_942_252#_c_534_n N_A_1555_367#_c_825_n 0.00630225f $X=7.707 $Y=1.49
+ $X2=0 $Y2=0
cc_430 N_A_942_252#_c_550_n N_A_1555_367#_c_825_n 0.0104983f $X=7.402 $Y=2.325
+ $X2=0 $Y2=0
cc_431 N_A_942_252#_c_538_n N_A_1555_367#_c_825_n 0.0207209f $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_432 N_A_942_252#_M1010_g N_A_1555_367#_c_819_n 0.00229383f $X=7.7 $Y=2.155
+ $X2=0 $Y2=0
cc_433 N_A_942_252#_M1011_g N_A_1555_367#_c_819_n 0.00436986f $X=7.715 $Y=0.93
+ $X2=0 $Y2=0
cc_434 N_A_942_252#_c_538_n N_A_1555_367#_c_819_n 0.0110918f $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_435 N_A_942_252#_c_539_n N_A_1555_367#_c_819_n 0.00171921f $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_436 N_A_942_252#_M1011_g N_A_1555_367#_c_820_n 3.61688e-19 $X=7.715 $Y=0.93
+ $X2=0 $Y2=0
cc_437 N_A_942_252#_c_538_n N_A_1555_367#_c_820_n 6.27541e-19 $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_438 N_A_942_252#_c_539_n N_A_1555_367#_c_820_n 0.0218591f $X=7.99 $Y=1.49
+ $X2=0 $Y2=0
cc_439 N_A_942_252#_c_548_n N_VPWR_M1020_s 0.00789799f $X=5.65 $Y=2.325 $X2=0
+ $Y2=0
cc_440 N_A_942_252#_c_558_p N_VPWR_M1020_s 0.00411973f $X=5.735 $Y=2.41 $X2=0
+ $Y2=0
cc_441 N_A_942_252#_c_549_n N_VPWR_M1006_d 0.00434914f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_442 N_A_942_252#_c_549_n N_VPWR_M1021_s 0.0035095f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_443 N_A_942_252#_c_550_n N_VPWR_M1021_s 0.00373515f $X=7.402 $Y=2.325 $X2=0
+ $Y2=0
cc_444 N_A_942_252#_M1005_g N_VPWR_c_881_n 0.00535895f $X=4.785 $Y=2.005 $X2=0
+ $Y2=0
cc_445 N_A_942_252#_c_558_p N_VPWR_c_882_n 0.0129733f $X=5.735 $Y=2.41 $X2=0
+ $Y2=0
cc_446 N_A_942_252#_M1000_g N_VPWR_c_883_n 0.0119622f $X=6.745 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_A_942_252#_M1021_g N_VPWR_c_883_n 0.00164057f $X=7.175 $Y=2.465 $X2=0
+ $Y2=0
cc_448 N_A_942_252#_c_549_n N_VPWR_c_883_n 0.0168972f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_449 N_A_942_252#_M1000_g N_VPWR_c_884_n 0.00171132f $X=6.745 $Y=2.465 $X2=0
+ $Y2=0
cc_450 N_A_942_252#_M1021_g N_VPWR_c_884_n 0.0153692f $X=7.175 $Y=2.465 $X2=0
+ $Y2=0
cc_451 N_A_942_252#_c_549_n N_VPWR_c_884_n 0.0237968f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_452 N_A_942_252#_M1010_g N_VPWR_c_885_n 0.00387011f $X=7.7 $Y=2.155 $X2=0
+ $Y2=0
cc_453 N_A_942_252#_c_578_p N_VPWR_c_893_n 0.0142265f $X=6.06 $Y=2.49 $X2=0
+ $Y2=0
cc_454 N_A_942_252#_M1000_g N_VPWR_c_894_n 0.00564095f $X=6.745 $Y=2.465 $X2=0
+ $Y2=0
cc_455 N_A_942_252#_M1021_g N_VPWR_c_894_n 0.00486043f $X=7.175 $Y=2.465 $X2=0
+ $Y2=0
cc_456 N_A_942_252#_M1010_g N_VPWR_c_895_n 0.00312414f $X=7.7 $Y=2.155 $X2=0
+ $Y2=0
cc_457 N_A_942_252#_M1020_d N_VPWR_c_877_n 0.00246871f $X=5.92 $Y=1.835 $X2=0
+ $Y2=0
cc_458 N_A_942_252#_M1000_g N_VPWR_c_877_n 0.00524988f $X=6.745 $Y=2.465 $X2=0
+ $Y2=0
cc_459 N_A_942_252#_M1021_g N_VPWR_c_877_n 0.00459245f $X=7.175 $Y=2.465 $X2=0
+ $Y2=0
cc_460 N_A_942_252#_M1010_g N_VPWR_c_877_n 0.00410284f $X=7.7 $Y=2.155 $X2=0
+ $Y2=0
cc_461 N_A_942_252#_c_568_p N_VPWR_c_877_n 0.00483499f $X=5.935 $Y=2.41 $X2=0
+ $Y2=0
cc_462 N_A_942_252#_c_558_p N_VPWR_c_877_n 6.19628e-19 $X=5.735 $Y=2.41 $X2=0
+ $Y2=0
cc_463 N_A_942_252#_c_549_n N_VPWR_c_877_n 0.0252579f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_464 N_A_942_252#_c_578_p N_VPWR_c_877_n 0.00925289f $X=6.06 $Y=2.49 $X2=0
+ $Y2=0
cc_465 N_A_942_252#_M1005_g N_A_606_359#_c_1003_n 0.0118015f $X=4.785 $Y=2.005
+ $X2=0 $Y2=0
cc_466 N_A_942_252#_c_535_n N_A_606_359#_c_1003_n 0.00880999f $X=5.465 $Y=1.465
+ $X2=0 $Y2=0
cc_467 N_A_942_252#_M1005_g N_A_606_359#_c_1005_n 0.0066464f $X=4.785 $Y=2.005
+ $X2=0 $Y2=0
cc_468 N_A_942_252#_c_535_n N_A_606_359#_c_1005_n 0.027278f $X=5.465 $Y=1.465
+ $X2=0 $Y2=0
cc_469 N_A_942_252#_c_536_n N_A_606_359#_c_1005_n 0.00129418f $X=4.875 $Y=1.425
+ $X2=0 $Y2=0
cc_470 N_A_942_252#_c_548_n N_A_606_359#_c_1005_n 0.0167758f $X=5.65 $Y=2.325
+ $X2=0 $Y2=0
cc_471 N_A_942_252#_c_549_n N_Q_M1000_d 0.00501287f $X=7.225 $Y=2.41 $X2=0 $Y2=0
cc_472 N_A_942_252#_M1009_g N_Q_c_1038_n 0.00258056f $X=6.745 $Y=0.72 $X2=0
+ $Y2=0
cc_473 N_A_942_252#_M1022_g N_Q_c_1038_n 5.3965e-19 $X=7.175 $Y=0.72 $X2=0 $Y2=0
cc_474 N_A_942_252#_c_532_n N_Q_c_1038_n 0.00135235f $X=7.25 $Y=1.49 $X2=0 $Y2=0
cc_475 N_A_942_252#_M1000_g N_Q_c_1040_n 0.00396943f $X=6.745 $Y=2.465 $X2=0
+ $Y2=0
cc_476 N_A_942_252#_c_532_n N_Q_c_1040_n 0.00129972f $X=7.25 $Y=1.49 $X2=0 $Y2=0
cc_477 N_A_942_252#_c_549_n N_Q_c_1040_n 0.0149496f $X=7.225 $Y=2.41 $X2=0 $Y2=0
cc_478 N_A_942_252#_c_550_n N_Q_c_1040_n 0.0136635f $X=7.402 $Y=2.325 $X2=0
+ $Y2=0
cc_479 N_A_942_252#_M1009_g N_Q_c_1039_n 0.00339022f $X=6.745 $Y=0.72 $X2=0
+ $Y2=0
cc_480 N_A_942_252#_M1000_g N_Q_c_1039_n 0.00277119f $X=6.745 $Y=2.465 $X2=0
+ $Y2=0
cc_481 N_A_942_252#_M1022_g N_Q_c_1039_n 0.00364839f $X=7.175 $Y=0.72 $X2=0
+ $Y2=0
cc_482 N_A_942_252#_M1021_g N_Q_c_1039_n 0.00111912f $X=7.175 $Y=2.465 $X2=0
+ $Y2=0
cc_483 N_A_942_252#_c_532_n N_Q_c_1039_n 0.0176605f $X=7.25 $Y=1.49 $X2=0 $Y2=0
cc_484 N_A_942_252#_c_646_p N_Q_c_1039_n 0.0123662f $X=7.402 $Y=1.575 $X2=0
+ $Y2=0
cc_485 N_A_942_252#_c_550_n N_Q_c_1039_n 0.0128098f $X=7.402 $Y=2.325 $X2=0
+ $Y2=0
cc_486 N_A_942_252#_M1009_g N_Q_c_1057_n 0.00813529f $X=6.745 $Y=0.72 $X2=0
+ $Y2=0
cc_487 N_A_942_252#_M1004_g N_VGND_c_1087_n 0.00340737f $X=4.855 $Y=0.615 $X2=0
+ $Y2=0
cc_488 N_A_942_252#_M1009_g N_VGND_c_1088_n 0.00609025f $X=6.745 $Y=0.72 $X2=0
+ $Y2=0
cc_489 N_A_942_252#_c_537_n N_VGND_c_1088_n 6.71991e-19 $X=5.63 $Y=0.445 $X2=0
+ $Y2=0
cc_490 N_A_942_252#_M1022_g N_VGND_c_1089_n 0.00661079f $X=7.175 $Y=0.72 $X2=0
+ $Y2=0
cc_491 N_A_942_252#_M1011_g N_VGND_c_1089_n 0.00451996f $X=7.715 $Y=0.93 $X2=0
+ $Y2=0
cc_492 N_A_942_252#_c_533_n N_VGND_c_1089_n 0.00521901f $X=7.625 $Y=1.49 $X2=0
+ $Y2=0
cc_493 N_A_942_252#_c_646_p N_VGND_c_1089_n 0.0196061f $X=7.402 $Y=1.575 $X2=0
+ $Y2=0
cc_494 N_A_942_252#_c_538_n N_VGND_c_1089_n 8.23339e-19 $X=7.99 $Y=1.49 $X2=0
+ $Y2=0
cc_495 N_A_942_252#_M1011_g N_VGND_c_1090_n 0.00329734f $X=7.715 $Y=0.93 $X2=0
+ $Y2=0
cc_496 N_A_942_252#_M1004_g N_VGND_c_1095_n 0.00552345f $X=4.855 $Y=0.615 $X2=0
+ $Y2=0
cc_497 N_A_942_252#_c_537_n N_VGND_c_1095_n 0.0165854f $X=5.63 $Y=0.445 $X2=0
+ $Y2=0
cc_498 N_A_942_252#_M1009_g N_VGND_c_1096_n 0.004915f $X=6.745 $Y=0.72 $X2=0
+ $Y2=0
cc_499 N_A_942_252#_M1022_g N_VGND_c_1096_n 0.00522039f $X=7.175 $Y=0.72 $X2=0
+ $Y2=0
cc_500 N_A_942_252#_M1011_g N_VGND_c_1097_n 0.00368595f $X=7.715 $Y=0.93 $X2=0
+ $Y2=0
cc_501 N_A_942_252#_M1004_g N_VGND_c_1104_n 0.00534666f $X=4.855 $Y=0.615 $X2=0
+ $Y2=0
cc_502 N_A_942_252#_M1009_g N_VGND_c_1104_n 0.00938496f $X=6.745 $Y=0.72 $X2=0
+ $Y2=0
cc_503 N_A_942_252#_M1022_g N_VGND_c_1104_n 0.0108352f $X=7.175 $Y=0.72 $X2=0
+ $Y2=0
cc_504 N_A_942_252#_M1011_g N_VGND_c_1104_n 0.00443953f $X=7.715 $Y=0.93 $X2=0
+ $Y2=0
cc_505 N_A_942_252#_c_537_n N_VGND_c_1104_n 0.0102927f $X=5.63 $Y=0.445 $X2=0
+ $Y2=0
cc_506 N_A_942_252#_M1004_g N_A_677_155#_c_1222_n 0.0177511f $X=4.855 $Y=0.615
+ $X2=0 $Y2=0
cc_507 N_A_942_252#_c_535_n N_A_677_155#_c_1222_n 0.0421022f $X=5.465 $Y=1.465
+ $X2=0 $Y2=0
cc_508 N_A_942_252#_c_536_n N_A_677_155#_c_1222_n 0.00475838f $X=4.875 $Y=1.425
+ $X2=0 $Y2=0
cc_509 N_A_942_252#_c_537_n N_A_677_155#_c_1222_n 0.0134002f $X=5.63 $Y=0.445
+ $X2=0 $Y2=0
cc_510 N_A_942_252#_M1004_g N_A_677_155#_c_1223_n 0.00630349f $X=4.855 $Y=0.615
+ $X2=0 $Y2=0
cc_511 N_A_942_252#_c_537_n N_A_677_155#_c_1223_n 0.0335897f $X=5.63 $Y=0.445
+ $X2=0 $Y2=0
cc_512 N_A_591_155#_c_677_n N_RESET_B_M1006_g 0.0399405f $X=5.845 $Y=1.65 $X2=0
+ $Y2=0
cc_513 N_A_591_155#_M1027_g RESET_B 0.00675604f $X=5.845 $Y=0.72 $X2=0 $Y2=0
cc_514 N_A_591_155#_c_685_n RESET_B 0.00893176f $X=5.845 $Y=1.725 $X2=0 $Y2=0
cc_515 N_A_591_155#_c_677_n RESET_B 0.00406703f $X=5.845 $Y=1.65 $X2=0 $Y2=0
cc_516 N_A_591_155#_c_677_n N_RESET_B_c_777_n 0.0427543f $X=5.845 $Y=1.65 $X2=0
+ $Y2=0
cc_517 N_A_591_155#_M1027_g N_RESET_B_c_778_n 0.0427543f $X=5.845 $Y=0.72 $X2=0
+ $Y2=0
cc_518 N_A_591_155#_c_681_n N_VPWR_c_881_n 0.0298801f $X=5.28 $Y=3.03 $X2=0
+ $Y2=0
cc_519 N_A_591_155#_c_682_n N_VPWR_c_881_n 0.0142785f $X=5.355 $Y=2.955 $X2=0
+ $Y2=0
cc_520 N_A_591_155#_c_690_n N_VPWR_c_881_n 0.0330211f $X=3.965 $Y=2.94 $X2=0
+ $Y2=0
cc_521 N_A_591_155#_c_691_n N_VPWR_c_881_n 0.00407707f $X=3.965 $Y=2.94 $X2=0
+ $Y2=0
cc_522 N_A_591_155#_c_692_n N_VPWR_c_881_n 0.0240516f $X=3.68 $Y=2.22 $X2=0
+ $Y2=0
cc_523 N_A_591_155#_c_682_n N_VPWR_c_882_n 0.0111555f $X=5.355 $Y=2.955 $X2=0
+ $Y2=0
cc_524 N_A_591_155#_c_685_n N_VPWR_c_882_n 0.00366673f $X=5.845 $Y=1.725 $X2=0
+ $Y2=0
cc_525 N_A_591_155#_c_685_n N_VPWR_c_883_n 5.57473e-19 $X=5.845 $Y=1.725 $X2=0
+ $Y2=0
cc_526 N_A_591_155#_c_681_n N_VPWR_c_890_n 0.0229955f $X=5.28 $Y=3.03 $X2=0
+ $Y2=0
cc_527 N_A_591_155#_c_688_n N_VPWR_c_892_n 0.00957164f $X=3.515 $Y=2.44 $X2=0
+ $Y2=0
cc_528 N_A_591_155#_c_689_n N_VPWR_c_892_n 0.00266576f $X=2.87 $Y=2.44 $X2=0
+ $Y2=0
cc_529 N_A_591_155#_c_690_n N_VPWR_c_892_n 0.0167839f $X=3.965 $Y=2.94 $X2=0
+ $Y2=0
cc_530 N_A_591_155#_c_691_n N_VPWR_c_892_n 0.0110745f $X=3.965 $Y=2.94 $X2=0
+ $Y2=0
cc_531 N_A_591_155#_c_692_n N_VPWR_c_892_n 0.00461844f $X=3.68 $Y=2.22 $X2=0
+ $Y2=0
cc_532 N_A_591_155#_c_685_n N_VPWR_c_893_n 0.00585385f $X=5.845 $Y=1.725 $X2=0
+ $Y2=0
cc_533 N_A_591_155#_c_681_n N_VPWR_c_877_n 0.0507977f $X=5.28 $Y=3.03 $X2=0
+ $Y2=0
cc_534 N_A_591_155#_c_685_n N_VPWR_c_877_n 0.00743389f $X=5.845 $Y=1.725 $X2=0
+ $Y2=0
cc_535 N_A_591_155#_c_688_n N_VPWR_c_877_n 0.0172056f $X=3.515 $Y=2.44 $X2=0
+ $Y2=0
cc_536 N_A_591_155#_c_689_n N_VPWR_c_877_n 0.00469963f $X=2.87 $Y=2.44 $X2=0
+ $Y2=0
cc_537 N_A_591_155#_c_690_n N_VPWR_c_877_n 0.0108843f $X=3.965 $Y=2.94 $X2=0
+ $Y2=0
cc_538 N_A_591_155#_c_691_n N_VPWR_c_877_n 0.00781325f $X=3.965 $Y=2.94 $X2=0
+ $Y2=0
cc_539 N_A_591_155#_c_692_n N_VPWR_c_877_n 0.00789651f $X=3.68 $Y=2.22 $X2=0
+ $Y2=0
cc_540 N_A_591_155#_M1024_d N_A_606_359#_c_1003_n 0.00295165f $X=3.445 $Y=1.795
+ $X2=0 $Y2=0
cc_541 N_A_591_155#_c_688_n N_A_606_359#_c_1003_n 0.00714148f $X=3.515 $Y=2.44
+ $X2=0 $Y2=0
cc_542 N_A_591_155#_c_692_n N_A_606_359#_c_1003_n 0.0316116f $X=3.68 $Y=2.22
+ $X2=0 $Y2=0
cc_543 N_A_591_155#_c_678_n N_A_606_359#_c_1004_n 0.0248562f $X=2.785 $Y=2.285
+ $X2=0 $Y2=0
cc_544 N_A_591_155#_c_688_n N_A_606_359#_c_1004_n 0.0202655f $X=3.515 $Y=2.44
+ $X2=0 $Y2=0
cc_545 N_A_591_155#_c_679_n N_A_606_359#_c_1004_n 0.0167909f $X=3.095 $Y=1.425
+ $X2=0 $Y2=0
cc_546 N_A_591_155#_c_682_n N_A_606_359#_c_1005_n 0.00449324f $X=5.355 $Y=2.955
+ $X2=0 $Y2=0
cc_547 N_A_591_155#_c_692_n A_794_359# 0.00147842f $X=3.68 $Y=2.22 $X2=-0.19
+ $Y2=-0.245
cc_548 N_A_591_155#_M1027_g N_VGND_c_1095_n 0.00522039f $X=5.845 $Y=0.72 $X2=0
+ $Y2=0
cc_549 N_A_591_155#_M1027_g N_VGND_c_1104_n 0.0109202f $X=5.845 $Y=0.72 $X2=0
+ $Y2=0
cc_550 N_A_591_155#_c_679_n N_A_508_155#_c_1204_n 0.00305114f $X=3.095 $Y=1.425
+ $X2=0 $Y2=0
cc_551 N_A_591_155#_M1025_d N_A_508_155#_c_1197_n 0.00176773f $X=2.955 $Y=0.775
+ $X2=0 $Y2=0
cc_552 N_A_591_155#_c_679_n N_A_508_155#_c_1197_n 0.00356936f $X=3.095 $Y=1.425
+ $X2=0 $Y2=0
cc_553 N_A_591_155#_c_680_n N_A_508_155#_c_1197_n 0.0166128f $X=3.095 $Y=1.07
+ $X2=0 $Y2=0
cc_554 RESET_B N_VPWR_M1006_d 0.00371401f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_555 N_RESET_B_M1006_g N_VPWR_c_883_n 0.00887602f $X=6.275 $Y=2.465 $X2=0
+ $Y2=0
cc_556 N_RESET_B_M1006_g N_VPWR_c_893_n 0.00564095f $X=6.275 $Y=2.465 $X2=0
+ $Y2=0
cc_557 N_RESET_B_M1006_g N_VPWR_c_877_n 0.00519715f $X=6.275 $Y=2.465 $X2=0
+ $Y2=0
cc_558 N_RESET_B_M1006_g N_Q_c_1039_n 4.12412e-19 $X=6.275 $Y=2.465 $X2=0 $Y2=0
cc_559 RESET_B N_Q_c_1039_n 0.0618476f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_560 N_RESET_B_c_777_n N_Q_c_1039_n 2.52588e-19 $X=6.295 $Y=1.415 $X2=0 $Y2=0
cc_561 N_RESET_B_c_778_n N_Q_c_1057_n 6.97664e-19 $X=6.295 $Y=1.25 $X2=0 $Y2=0
cc_562 RESET_B N_VGND_c_1088_n 0.0278086f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_563 N_RESET_B_c_777_n N_VGND_c_1088_n 0.0010452f $X=6.295 $Y=1.415 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_778_n N_VGND_c_1088_n 0.00394727f $X=6.295 $Y=1.25 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_778_n N_VGND_c_1095_n 0.00522039f $X=6.295 $Y=1.25 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_778_n N_VGND_c_1104_n 0.0100951f $X=6.295 $Y=1.25 $X2=0 $Y2=0
cc_567 N_A_1555_367#_c_824_n N_VPWR_M1001_s 0.00275572f $X=8.365 $Y=1.84 $X2=0
+ $Y2=0
cc_568 N_A_1555_367#_M1001_g N_VPWR_c_885_n 0.0144732f $X=8.685 $Y=2.465 $X2=0
+ $Y2=0
cc_569 N_A_1555_367#_M1023_g N_VPWR_c_885_n 7.25278e-19 $X=9.115 $Y=2.465 $X2=0
+ $Y2=0
cc_570 N_A_1555_367#_c_823_n N_VPWR_c_885_n 0.0211306f $X=7.915 $Y=1.98 $X2=0
+ $Y2=0
cc_571 N_A_1555_367#_c_824_n N_VPWR_c_885_n 0.0212472f $X=8.365 $Y=1.84 $X2=0
+ $Y2=0
cc_572 N_A_1555_367#_c_820_n N_VPWR_c_885_n 9.38299e-19 $X=8.562 $Y=1.385 $X2=0
+ $Y2=0
cc_573 N_A_1555_367#_M1023_g N_VPWR_c_887_n 0.00764209f $X=9.115 $Y=2.465 $X2=0
+ $Y2=0
cc_574 N_A_1555_367#_M1001_g N_VPWR_c_896_n 0.00525069f $X=8.685 $Y=2.465 $X2=0
+ $Y2=0
cc_575 N_A_1555_367#_M1023_g N_VPWR_c_896_n 0.00585385f $X=9.115 $Y=2.465 $X2=0
+ $Y2=0
cc_576 N_A_1555_367#_M1001_g N_VPWR_c_877_n 0.00886509f $X=8.685 $Y=2.465 $X2=0
+ $Y2=0
cc_577 N_A_1555_367#_M1023_g N_VPWR_c_877_n 0.011478f $X=9.115 $Y=2.465 $X2=0
+ $Y2=0
cc_578 N_A_1555_367#_c_823_n N_VPWR_c_877_n 0.0104273f $X=7.915 $Y=1.98 $X2=0
+ $Y2=0
cc_579 N_A_1555_367#_M1003_g N_Q_N_c_1066_n 0.0023234f $X=8.685 $Y=0.69 $X2=0
+ $Y2=0
cc_580 N_A_1555_367#_c_814_n N_Q_N_c_1066_n 0.0162773f $X=9.04 $Y=1.385 $X2=0
+ $Y2=0
cc_581 N_A_1555_367#_M1013_g N_Q_N_c_1066_n 0.00588371f $X=9.115 $Y=0.69 $X2=0
+ $Y2=0
cc_582 N_A_1555_367#_M1023_g N_Q_N_c_1066_n 0.0104972f $X=9.115 $Y=2.465 $X2=0
+ $Y2=0
cc_583 N_A_1555_367#_c_818_n N_Q_N_c_1066_n 0.00940486f $X=8.365 $Y=1 $X2=0
+ $Y2=0
cc_584 N_A_1555_367#_c_824_n N_Q_N_c_1066_n 0.00985831f $X=8.365 $Y=1.84 $X2=0
+ $Y2=0
cc_585 N_A_1555_367#_c_819_n N_Q_N_c_1066_n 0.0456233f $X=8.53 $Y=1.475 $X2=0
+ $Y2=0
cc_586 N_A_1555_367#_c_820_n N_Q_N_c_1066_n 0.00372991f $X=8.562 $Y=1.385 $X2=0
+ $Y2=0
cc_587 N_A_1555_367#_c_818_n N_VGND_M1003_d 0.00379195f $X=8.365 $Y=1 $X2=0
+ $Y2=0
cc_588 N_A_1555_367#_M1003_g N_VGND_c_1090_n 0.0108458f $X=8.685 $Y=0.69 $X2=0
+ $Y2=0
cc_589 N_A_1555_367#_M1013_g N_VGND_c_1090_n 5.01913e-19 $X=9.115 $Y=0.69 $X2=0
+ $Y2=0
cc_590 N_A_1555_367#_c_818_n N_VGND_c_1090_n 0.0238937f $X=8.365 $Y=1 $X2=0
+ $Y2=0
cc_591 N_A_1555_367#_c_820_n N_VGND_c_1090_n 7.37395e-19 $X=8.562 $Y=1.385 $X2=0
+ $Y2=0
cc_592 N_A_1555_367#_M1013_g N_VGND_c_1092_n 0.00702119f $X=9.115 $Y=0.69 $X2=0
+ $Y2=0
cc_593 N_A_1555_367#_M1003_g N_VGND_c_1098_n 0.00530359f $X=8.685 $Y=0.69 $X2=0
+ $Y2=0
cc_594 N_A_1555_367#_M1013_g N_VGND_c_1098_n 0.00550375f $X=9.115 $Y=0.69 $X2=0
+ $Y2=0
cc_595 N_A_1555_367#_M1003_g N_VGND_c_1104_n 0.00941735f $X=8.685 $Y=0.69 $X2=0
+ $Y2=0
cc_596 N_A_1555_367#_M1013_g N_VGND_c_1104_n 0.0111259f $X=9.115 $Y=0.69 $X2=0
+ $Y2=0
cc_597 N_VPWR_M1018_d N_A_606_359#_c_1003_n 0.00337793f $X=4.33 $Y=1.795 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_881_n N_A_606_359#_c_1003_n 0.0219076f $X=4.475 $Y=2.245 $X2=0
+ $Y2=0
cc_599 N_VPWR_c_881_n N_A_606_359#_c_1005_n 0.00384115f $X=4.475 $Y=2.245 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_877_n N_Q_M1000_d 0.00408795f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_601 N_VPWR_c_877_n N_Q_N_M1001_d 0.00362709f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_602 N_VPWR_c_887_n N_Q_N_c_1066_n 0.00152843f $X=9.33 $Y=1.98 $X2=0 $Y2=0
cc_603 N_VPWR_c_896_n N_Q_N_c_1066_n 0.0142265f $X=9.205 $Y=3.33 $X2=0 $Y2=0
cc_604 N_VPWR_c_877_n N_Q_N_c_1066_n 0.00925289f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_605 N_A_606_359#_c_1003_n A_794_359# 0.00141317f $X=4.835 $Y=1.86 $X2=-0.19
+ $Y2=1.655
cc_606 N_A_606_359#_c_1003_n N_A_677_155#_c_1222_n 0.0368825f $X=4.835 $Y=1.86
+ $X2=0 $Y2=0
cc_607 N_Q_c_1038_n N_VGND_c_1089_n 9.52992e-19 $X=6.93 $Y=1.155 $X2=0 $Y2=0
cc_608 N_Q_c_1057_n N_VGND_c_1096_n 0.0103941f $X=6.96 $Y=0.505 $X2=0 $Y2=0
cc_609 N_Q_c_1057_n N_VGND_c_1104_n 0.00982997f $X=6.96 $Y=0.505 $X2=0 $Y2=0
cc_610 N_Q_N_c_1066_n N_VGND_c_1090_n 0.0170201f $X=8.9 $Y=0.42 $X2=0 $Y2=0
cc_611 N_Q_N_c_1066_n N_VGND_c_1092_n 0.00265464f $X=8.9 $Y=0.42 $X2=0 $Y2=0
cc_612 N_Q_N_c_1066_n N_VGND_c_1098_n 0.0170614f $X=8.9 $Y=0.42 $X2=0 $Y2=0
cc_613 N_Q_N_c_1066_n N_VGND_c_1104_n 0.00925289f $X=8.9 $Y=0.42 $X2=0 $Y2=0
cc_614 N_VGND_c_1094_n N_A_508_155#_c_1197_n 0.00729258f $X=4.545 $Y=0 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1104_n N_A_508_155#_c_1197_n 0.0145177f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_616 N_VGND_c_1087_n N_A_677_155#_c_1222_n 0.0140743f $X=4.64 $Y=0.6 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1095_n N_A_677_155#_c_1223_n 0.00834666f $X=6.295 $Y=0 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1104_n N_A_677_155#_c_1223_n 0.0102973f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_619 N_A_508_155#_c_1197_n N_A_677_155#_M1019_d 0.00280397f $X=4.21 $Y=0.7
+ $X2=-0.19 $Y2=-0.245
cc_620 N_A_508_155#_c_1197_n N_A_677_155#_c_1222_n 0.0649641f $X=4.21 $Y=0.7
+ $X2=0 $Y2=0
