* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4bb_lp A_N B_N C D VGND VNB VPB VPWR X
X0 a_291_409# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_461_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_896_47# a_461_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_704_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR C a_461_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_272_51# B_N a_291_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_461_47# a_896_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_626_47# C a_704_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_461_47# a_291_409# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VPWR a_27_51# a_461_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_114_51# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_27_51# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_461_47# a_27_51# a_548_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_51# A_N a_114_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND B_N a_272_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VPWR a_461_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_548_47# a_291_409# a_626_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
