* File: sky130_fd_sc_lp__o41a_lp.pex.spice
* Created: Fri Aug 28 11:19:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41A_LP%A1 3 7 11 12 13 16 17
c35 7 0 1.79304e-19 $X=0.515 $Y=0.495
r36 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.52
+ $Y=1.355 $X2=0.52 $Y2=1.355
r37 13 17 4.99854 $w=6.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=1.525
+ $X2=0.52 $Y2=1.525
r38 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.52 $Y=1.695
+ $X2=0.52 $Y2=1.355
r39 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.695
+ $X2=0.52 $Y2=1.86
r40 10 16 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.19
+ $X2=0.52 $Y2=1.355
r41 7 10 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.515 $Y=0.495
+ $X2=0.515 $Y2=1.19
r42 3 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.56 $Y=2.56 $X2=0.56
+ $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_LP%A2 3 7 11 12 13 14 15 16 22 23
r46 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.09
+ $Y=1.395 $X2=1.09 $Y2=1.395
r47 15 16 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.12 $Y=2.405
+ $X2=1.12 $Y2=2.775
r48 14 15 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.12 $Y=2.035
+ $X2=1.12 $Y2=2.405
r49 13 14 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=2.035
r50 13 23 7.97845 $w=3.88e-07 $l=2.7e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.395
r51 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.09 $Y=1.735
+ $X2=1.09 $Y2=1.395
r52 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.735
+ $X2=1.09 $Y2=1.9
r53 10 22 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.23
+ $X2=1.09 $Y2=1.395
r54 7 10 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.105 $Y=0.495
+ $X2=1.105 $Y2=1.23
r55 3 12 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.05 $Y=2.56 $X2=1.05
+ $Y2=1.9
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_LP%A3 3 7 11 12 13 14 15 16 22 23
r42 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.66
+ $Y=1.395 $X2=1.66 $Y2=1.395
r43 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=2.405
+ $X2=1.66 $Y2=2.775
r44 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=2.035
+ $X2=1.66 $Y2=2.405
r45 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=1.665
+ $X2=1.66 $Y2=2.035
r46 13 23 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.66 $Y=1.665
+ $X2=1.66 $Y2=1.395
r47 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.66 $Y=1.735
+ $X2=1.66 $Y2=1.395
r48 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.735
+ $X2=1.66 $Y2=1.9
r49 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.23
+ $X2=1.66 $Y2=1.395
r50 7 12 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.62 $Y=2.56 $X2=1.62
+ $Y2=1.9
r51 3 10 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.57 $Y=0.495
+ $X2=1.57 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_LP%A4 3 8 10 11 13 14 15 16 17 18 19 25 26
c54 11 0 2.55406e-19 $X=2.077 $Y=0.93
r55 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.2
+ $Y=1.395 $X2=2.2 $Y2=1.395
r56 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.2 $Y=2.405 $X2=2.2
+ $Y2=2.775
r57 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.2 $Y=2.035 $X2=2.2
+ $Y2=2.405
r58 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.2 $Y=1.665 $X2=2.2
+ $Y2=2.035
r59 16 26 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.2 $Y=1.665 $X2=2.2
+ $Y2=1.395
r60 14 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.2 $Y=1.735 $X2=2.2
+ $Y2=1.395
r61 14 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.735
+ $X2=2.2 $Y2=1.9
r62 13 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.23 $X2=2.2
+ $Y2=1.395
r63 11 13 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.11 $Y=0.93 $X2=2.11
+ $Y2=1.23
r64 10 11 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=2.077 $Y=0.78
+ $X2=2.077 $Y2=0.93
r65 8 15 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.16 $Y=2.56 $X2=2.16
+ $Y2=1.9
r66 3 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.045 $Y=0.495
+ $X2=2.045 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_LP%B1 1 3 5 6 8 12 14
r55 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.835
+ $Y=1.345 $X2=2.835 $Y2=1.345
r56 14 18 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.12 $Y=1.345
+ $X2=2.835 $Y2=1.345
r57 10 12 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.475 $Y=0.855
+ $X2=2.745 $Y2=0.855
r58 6 17 61.5611 $w=2.86e-07 $l=4.02492e-07 $layer=POLY_cond $X=2.975 $Y=1.705
+ $X2=2.885 $Y2=1.345
r59 6 8 212.428 $w=2.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.975 $Y=1.705
+ $X2=2.975 $Y2=2.56
r60 5 17 38.6549 $w=2.86e-07 $l=2.24332e-07 $layer=POLY_cond $X=2.745 $Y=1.18
+ $X2=2.885 $Y2=1.345
r61 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.745 $Y=0.93
+ $X2=2.745 $Y2=0.855
r62 4 5 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.745 $Y=0.93
+ $X2=2.745 $Y2=1.18
r63 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.475 $Y=0.78
+ $X2=2.475 $Y2=0.855
r64 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.475 $Y=0.78 $X2=2.475
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_LP%A_457_412# 1 2 9 13 17 21 23 26 30 34 35 36
+ 37 41 43 44 45
c84 35 0 7.90676e-20 $X=2.855 $Y=0.915
c85 26 0 3.87244e-20 $X=2.69 $Y=0.495
r86 43 45 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=1.355
+ $X2=3.58 $Y2=1.19
r87 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.58
+ $Y=1.355 $X2=3.58 $Y2=1.355
r88 41 43 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.58 $Y=1.69
+ $X2=3.58 $Y2=1.355
r89 38 45 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.5 $Y=1 $X2=3.5
+ $Y2=1.19
r90 36 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.415 $Y=1.775
+ $X2=3.58 $Y2=1.69
r91 36 37 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.415 $Y=1.775
+ $X2=2.875 $Y2=1.775
r92 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.415 $Y=0.915
+ $X2=3.5 $Y2=1
r93 34 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.415 $Y=0.915
+ $X2=2.855 $Y2=0.915
r94 30 32 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.71 $Y=2.205
+ $X2=2.71 $Y2=2.9
r95 28 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.71 $Y=1.86
+ $X2=2.875 $Y2=1.775
r96 28 30 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.71 $Y=1.86
+ $X2=2.71 $Y2=2.205
r97 24 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.69 $Y=0.83
+ $X2=2.855 $Y2=0.915
r98 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.69 $Y=0.83
+ $X2=2.69 $Y2=0.495
r99 22 44 53.3155 $w=3.55e-07 $l=3.28e-07 $layer=POLY_cond $X=3.567 $Y=1.683
+ $X2=3.567 $Y2=1.355
r100 22 23 33.8903 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=3.567 $Y=1.683
+ $X2=3.567 $Y2=1.86
r101 21 44 2.43821 $w=3.55e-07 $l=1.5e-08 $layer=POLY_cond $X=3.567 $Y=1.34
+ $X2=3.567 $Y2=1.355
r102 13 23 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.62 $Y=2.56 $X2=3.62
+ $Y2=1.86
r103 7 21 25.9344 $w=3.55e-07 $l=1.5e-07 $layer=POLY_cond $X=3.645 $Y=1.19
+ $X2=3.645 $Y2=1.34
r104 7 17 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.825 $Y=1.19
+ $X2=3.825 $Y2=0.445
r105 7 9 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.465 $Y=1.19
+ $X2=3.465 $Y2=0.445
r106 2 32 400 $w=1.7e-07 $l=1.03082e-06 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=2.06 $X2=2.71 $Y2=2.9
r107 2 30 400 $w=1.7e-07 $l=4.92189e-07 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=2.06 $X2=2.71 $Y2=2.205
r108 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.285 $X2=2.69 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_LP%VPWR 1 2 7 9 15 19 21 28 29 35
r41 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 29 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 26 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.24 $Y2=3.33
r46 26 28 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=4.08 $Y2=3.33
r47 25 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 24 25 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 22 32 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=3.33 $X2=0.23
+ $Y2=3.33
r50 22 24 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 21 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=3.33
+ $X2=3.24 $Y2=3.33
r52 21 24 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=3.075 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 19 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 19 25 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.24 $Y=2.205
+ $X2=3.24 $Y2=2.915
r56 13 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=3.245
+ $X2=3.24 $Y2=3.33
r57 13 18 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.24 $Y=3.245
+ $X2=3.24 $Y2=2.915
r58 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.295 $Y=2.205
+ $X2=0.295 $Y2=2.915
r59 7 32 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.23 $Y2=3.33
r60 7 12 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.915
r61 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.1
+ $Y=2.06 $X2=3.24 $Y2=2.915
r62 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.1
+ $Y=2.06 $X2=3.24 $Y2=2.205
r63 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.06 $X2=0.295 $Y2=2.915
r64 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.06 $X2=0.295 $Y2=2.205
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_LP%X 1 2 7 8 9 10 11 12 13 32
r27 33 49 1.89893 $w=4.83e-07 $l=7.7e-08 $layer=LI1_cond $X=3.962 $Y=2.282
+ $X2=3.962 $Y2=2.205
r28 32 47 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=4.085 $Y=2.035
+ $X2=4.085 $Y2=2.04
r29 13 39 3.08268 $w=4.83e-07 $l=1.25e-07 $layer=LI1_cond $X=3.962 $Y=2.775
+ $X2=3.962 $Y2=2.9
r30 12 13 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.962 $Y=2.405
+ $X2=3.962 $Y2=2.775
r31 12 33 3.03335 $w=4.83e-07 $l=1.23e-07 $layer=LI1_cond $X=3.962 $Y=2.405
+ $X2=3.962 $Y2=2.282
r32 11 49 3.08268 $w=4.83e-07 $l=1.25e-07 $layer=LI1_cond $X=3.962 $Y=2.08
+ $X2=3.962 $Y2=2.205
r33 11 47 4.03982 $w=4.83e-07 $l=4e-08 $layer=LI1_cond $X=3.962 $Y=2.08
+ $X2=3.962 $Y2=2.04
r34 11 32 1.92074 $w=2.38e-07 $l=4e-08 $layer=LI1_cond $X=4.085 $Y=1.995
+ $X2=4.085 $Y2=2.035
r35 10 11 15.8461 $w=2.38e-07 $l=3.3e-07 $layer=LI1_cond $X=4.085 $Y=1.665
+ $X2=4.085 $Y2=1.995
r36 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.085 $Y=1.295
+ $X2=4.085 $Y2=1.665
r37 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.085 $Y=0.925
+ $X2=4.085 $Y2=1.295
r38 8 45 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=4.085 $Y=0.925
+ $X2=4.085 $Y2=0.675
r39 7 45 8.03684 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.04 $Y=0.47
+ $X2=4.04 $Y2=0.675
r40 2 49 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=2.06 $X2=3.885 $Y2=2.205
r41 2 39 400 $w=1.7e-07 $l=9.07304e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=2.06 $X2=3.885 $Y2=2.9
r42 1 7 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_LP%A_31_57# 1 2 3 12 14 15 18 20 24 26
c54 26 0 1.79304e-19 $X=1.32 $Y=0.945
r55 22 24 17.7476 $w=2.48e-07 $l=3.85e-07 $layer=LI1_cond $X=2.22 $Y=0.88
+ $X2=2.22 $Y2=0.495
r56 21 26 8.61065 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=1.485 $Y=0.965
+ $X2=1.32 $Y2=0.945
r57 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.095 $Y=0.965
+ $X2=2.22 $Y2=0.88
r58 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.095 $Y=0.965
+ $X2=1.485 $Y2=0.965
r59 16 26 0.89609 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=1.32 $Y=0.84
+ $X2=1.32 $Y2=0.945
r60 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.32 $Y=0.84
+ $X2=1.32 $Y2=0.495
r61 14 26 8.61065 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=1.155 $Y=0.925
+ $X2=1.32 $Y2=0.945
r62 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.155 $Y=0.925
+ $X2=0.465 $Y2=0.925
r63 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.3 $Y=0.84
+ $X2=0.465 $Y2=0.925
r64 10 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.3 $Y=0.84 $X2=0.3
+ $Y2=0.495
r65 3 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.285 $X2=2.26 $Y2=0.495
r66 2 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.18
+ $Y=0.285 $X2=1.32 $Y2=0.495
r67 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.285 $X2=0.3 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_LP%VGND 1 2 3 14 16 20 24 26 28 35 36 39 42 45
c55 28 0 1.37614e-19 $X=3.085 $Y=0
r56 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r58 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r59 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r60 36 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r61 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r62 33 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.25
+ $Y2=0
r63 33 35 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=4.08
+ $Y2=0
r64 29 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=1.79
+ $Y2=0
r65 29 31 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=2.16
+ $Y2=0
r66 28 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.25
+ $Y2=0
r67 28 31 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=2.16
+ $Y2=0
r68 26 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r69 26 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r70 26 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r71 22 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0
r72 22 24 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0.43
r73 18 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=0.085
+ $X2=1.79 $Y2=0
r74 18 20 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=1.79 $Y=0.085
+ $X2=1.79 $Y2=0.48
r75 17 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.81
+ $Y2=0
r76 16 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.665 $Y=0 $X2=1.79
+ $Y2=0
r77 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.665 $Y=0 $X2=0.975
+ $Y2=0
r78 12 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=0.085
+ $X2=0.81 $Y2=0
r79 12 14 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.81 $Y=0.085
+ $X2=0.81 $Y2=0.46
r80 3 24 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=3.105
+ $Y=0.235 $X2=3.25 $Y2=0.43
r81 2 20 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.285 $X2=1.83 $Y2=0.48
r82 1 14 182 $w=1.7e-07 $l=2.94788e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.285 $X2=0.81 $Y2=0.46
.ends

