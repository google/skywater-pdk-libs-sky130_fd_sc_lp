* File: sky130_fd_sc_lp__lsbufiso1p_lp.pex.spice
* Created: Wed Sep  2 09:59:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%VGND 1 2 3 4 29 45 49 53 57 70 71 75
+ 78 82 91 98 105
c172 70 0 1.58517e-19 $X=2.87 $Y=3.33
c173 57 0 5.05501e-20 $X=5.665 $Y=3.715
r174 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.955 $Y=3.33
+ $X2=6.955 $Y2=3.33
r175 94 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r176 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r177 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.32
+ $X2=0.72 $Y2=3.32
r178 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r179 86 98 0.132399 $w=4.9e-07 $l=4.75e-07 $layer=MET1_cond $X=6.48 $Y=3.32
+ $X2=6.955 $Y2=3.32
r180 86 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.32
+ $X2=5.52 $Y2=3.32
r181 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r182 83 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=5.665 $Y2=3.33
r183 83 85 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=6.48 $Y2=3.33
r184 82 97 3.44808 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=6.81 $Y=3.33
+ $X2=7.005 $Y2=3.33
r185 82 85 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.81 $Y=3.33
+ $X2=6.48 $Y2=3.33
r186 81 105 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.12 $Y=3.32
+ $X2=3.36 $Y2=3.32
r187 80 81 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r188 78 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.5 $Y=3.33
+ $X2=5.665 $Y2=3.33
r189 78 80 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=5.5 $Y=3.33
+ $X2=3.12 $Y2=3.33
r190 76 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.32
+ $X2=3.12 $Y2=3.32
r191 76 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.32
+ $X2=0.72 $Y2=3.32
r192 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r193 73 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r194 73 75 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r195 71 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.32
+ $X2=5.52 $Y2=3.32
r196 71 105 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.6 $Y=3.32
+ $X2=3.36 $Y2=3.32
r197 69 80 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.04 $Y=3.33 $X2=3.12
+ $Y2=3.33
r198 69 70 3.86674 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.04 $Y=3.33
+ $X2=2.87 $Y2=3.33
r199 64 97 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=6.96 $Y=3.415
+ $X2=7.005 $Y2=3.33
r200 59 97 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=6.96 $Y=3.245
+ $X2=7.005 $Y2=3.33
r201 55 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.665 $Y=3.415
+ $X2=5.665 $Y2=3.33
r202 55 57 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=5.665 $Y=3.415
+ $X2=5.665 $Y2=3.715
r203 51 70 2.84813 $w=3.35e-07 $l=8.74643e-08 $layer=LI1_cond $X=2.865 $Y=3.415
+ $X2=2.87 $Y2=3.33
r204 51 53 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=2.865 $Y=3.415
+ $X2=2.865 $Y2=4.155
r205 47 70 2.84813 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=3.245
+ $X2=2.87 $Y2=3.33
r206 47 49 24.7436 $w=3.38e-07 $l=7.3e-07 $layer=LI1_cond $X=2.87 $Y=3.245
+ $X2=2.87 $Y2=2.515
r207 43 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=3.33
r208 43 45 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=2.44
r209 42 88 3.44808 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r210 41 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r211 41 42 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.39 $Y2=3.33
r212 36 88 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.24 $Y=3.415
+ $X2=0.195 $Y2=3.33
r213 31 88 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.195 $Y2=3.33
r214 29 64 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=6.96 $Y=3.855
+ $X2=6.96 $Y2=3.415
r215 29 59 32.8446 $w=2.98e-07 $l=8.55e-07 $layer=LI1_cond $X=6.96 $Y=2.39
+ $X2=6.96 $Y2=3.245
r216 29 36 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=0.24 $Y=3.855
+ $X2=0.24 $Y2=3.415
r217 29 31 32.8446 $w=2.98e-07 $l=8.55e-07 $layer=LI1_cond $X=0.24 $Y=2.39
+ $X2=0.24 $Y2=3.245
r218 4 57 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.52
+ $Y=3.59 $X2=5.665 $Y2=3.715
r219 3 53 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.74
+ $Y=4.01 $X2=2.865 $Y2=4.155
r220 2 49 91 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=2 $X=2.735
+ $Y=2.23 $X2=2.875 $Y2=2.515
r221 1 45 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=2.23 $X2=0.74 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%VPB 7 9 10 11 12 13 14
r19 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=6.96 $Y=0.925
+ $X2=6.96 $Y2=1.295
r20 12 13 15.3659 $w=2.98e-07 $l=4e-07 $layer=LI1_cond $X=6.96 $Y=0.525 $X2=6.96
+ $Y2=0.925
r21 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.295
r22 9 10 15.3659 $w=2.98e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=0.525 $X2=0.24
+ $Y2=0.925
r23 7 12 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=6.875 $Y=0.32 $X2=6.96 $Y2=0.525
r24 7 9 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0.155
+ $Y=0.32 $X2=0.24 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%DESTVPB 7 9 10 11 12 13 14
r61 13 14 15.558 $w=2.98e-07 $l=4.05e-07 $layer=LI1_cond $X=6.96 $Y=5.7 $X2=6.96
+ $Y2=6.105
r62 12 13 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.96 $Y=5.365
+ $X2=6.96 $Y2=5.7
r63 10 11 15.558 $w=2.98e-07 $l=4.05e-07 $layer=LI1_cond $X=0.24 $Y=5.7 $X2=0.24
+ $Y2=6.105
r64 9 10 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=5.365
+ $X2=0.24 $Y2=5.7
r65 7 13 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=6.875 $Y=5.495 $X2=6.96 $Y2=5.7
r66 7 10 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=0.155 $Y=5.495 $X2=0.24 $Y2=5.7
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_176_987# 1 2 9 13 15 18 21 24 28 31
+ 35
c77 18 0 1.70849e-20 $X=2.24 $Y=5.355
r78 28 30 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=4.235
+ $X2=2.32 $Y2=4.4
r79 25 35 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.165 $Y=5.1
+ $X2=1.315 $Y2=5.1
r80 25 32 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.165 $Y=5.1
+ $X2=0.955 $Y2=5.1
r81 24 26 16.4603 $w=2.52e-07 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=5.1
+ $X2=1.165 $Y2=5.44
r82 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=5.1 $X2=1.165 $Y2=5.1
r83 19 31 3.70735 $w=2.5e-07 $l=2.38642e-07 $layer=LI1_cond $X=2.32 $Y=5.525
+ $X2=2.155 $Y2=5.355
r84 19 21 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.32 $Y=5.525
+ $X2=2.32 $Y2=5.55
r85 18 31 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=5.355
+ $X2=2.155 $Y2=5.355
r86 18 30 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.24 $Y=5.355
+ $X2=2.24 $Y2=4.4
r87 16 26 3.04159 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.33 $Y=5.44
+ $X2=1.165 $Y2=5.44
r88 15 31 2.76166 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=5.44
+ $X2=2.155 $Y2=5.355
r89 15 16 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.155 $Y=5.44
+ $X2=1.33 $Y2=5.44
r90 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.315 $Y=5.265
+ $X2=1.315 $Y2=5.1
r91 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.315 $Y=5.265
+ $X2=1.315 $Y2=5.925
r92 7 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=5.265
+ $X2=0.955 $Y2=5.1
r93 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=5.265
+ $X2=0.955 $Y2=5.925
r94 2 21 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.18
+ $Y=5.425 $X2=2.32 $Y2=5.55
r95 1 28 182 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_NDIFF $count=1 $X=2.18
+ $Y=3.59 $X2=2.32 $Y2=4.235
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A 3 5 7 10 12 13 16 21 22 24 27 31 34
+ 43 51
c72 27 0 3.44129e-20 $X=1.16 $Y=2.775
r73 42 43 61.0986 $w=3.4e-07 $l=3.6e-07 $layer=POLY_cond $X=0.955 $Y=1.96
+ $X2=1.315 $Y2=1.96
r74 39 42 34.7923 $w=3.4e-07 $l=2.05e-07 $layer=POLY_cond $X=0.75 $Y=1.96
+ $X2=0.955 $Y2=1.96
r75 34 51 8.5999 $w=6.03e-07 $l=4.35e-07 $layer=LI1_cond $X=0.725 $Y=1.832
+ $X2=1.16 $Y2=1.832
r76 34 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.955 $X2=0.75 $Y2=1.955
r77 32 46 22.0523 $w=3.06e-07 $l=1.4e-07 $layer=POLY_cond $X=1.405 $Y=2.925
+ $X2=1.405 $Y2=3.065
r78 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.405
+ $Y=2.925 $X2=1.405 $Y2=2.925
r79 28 31 9.41162 $w=2.98e-07 $l=2.45e-07 $layer=LI1_cond $X=1.16 $Y=2.925
+ $X2=1.405 $Y2=2.925
r80 27 28 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.16 $Y=2.775 $X2=1.16
+ $Y2=2.925
r81 26 51 8.37032 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=1.16 $Y=2.135
+ $X2=1.16 $Y2=1.832
r82 26 27 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.16 $Y=2.135
+ $X2=1.16 $Y2=2.775
r83 22 46 24.3585 $w=3.06e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.315 $Y=3.14
+ $X2=1.405 $Y2=3.065
r84 22 24 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.315 $Y=3.14
+ $X2=1.315 $Y2=4.01
r85 19 32 38.535 $w=3.06e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.315 $Y=2.76
+ $X2=1.405 $Y2=2.925
r86 19 21 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.315 $Y=2.76
+ $X2=1.315 $Y2=2.44
r87 18 43 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.315 $Y=2.13
+ $X2=1.315 $Y2=1.96
r88 18 21 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.315 $Y=2.13
+ $X2=1.315 $Y2=2.44
r89 14 43 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.315 $Y=1.79
+ $X2=1.315 $Y2=1.96
r90 14 16 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=1.315 $Y=1.79
+ $X2=1.315 $Y2=0.735
r91 12 46 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.24 $Y=3.065
+ $X2=1.405 $Y2=3.065
r92 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.24 $Y=3.065
+ $X2=1.03 $Y2=3.065
r93 8 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.955 $Y=3.14
+ $X2=1.03 $Y2=3.065
r94 8 10 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=0.955 $Y=3.14
+ $X2=0.955 $Y2=4.01
r95 5 42 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.955 $Y=2.13
+ $X2=0.955 $Y2=1.96
r96 5 7 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.955 $Y=2.13
+ $X2=0.955 $Y2=2.44
r97 1 42 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.955 $Y=1.79
+ $X2=0.955 $Y2=1.96
r98 1 3 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=0.955 $Y=1.79
+ $X2=0.955 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_278_47# 1 2 7 9 10 11 13 14 16 17 20
+ 26 28 29 31 33
c71 29 0 3.44129e-20 $X=1.98 $Y=2.925
r72 31 33 41.2959 $w=2.98e-07 $l=1.075e-06 $layer=LI1_cond $X=1.565 $Y=1.36
+ $X2=1.565 $Y2=2.435
r73 29 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=2.925
+ $X2=1.98 $Y2=3.09
r74 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.98
+ $Y=2.925 $X2=1.98 $Y2=2.925
r75 26 33 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.98 $Y=2.52
+ $X2=1.53 $Y2=2.52
r76 26 28 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.98 $Y=2.605
+ $X2=1.98 $Y2=2.925
r77 20 23 23.3781 $w=3.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.54 $Y=0.38
+ $X2=1.54 $Y2=1.09
r78 18 31 6.02978 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=1.54 $Y=1.185
+ $X2=1.54 $Y2=1.36
r79 18 23 3.12806 $w=3.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.54 $Y=1.185
+ $X2=1.54 $Y2=1.09
r80 14 17 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=2.105 $Y=3.515
+ $X2=2.087 $Y2=3.44
r81 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.105 $Y=3.515
+ $X2=2.105 $Y2=4.01
r82 13 17 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=2.07 $Y=3.365
+ $X2=2.087 $Y2=3.44
r83 13 39 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=2.07 $Y=3.365
+ $X2=2.07 $Y2=3.09
r84 10 17 5.30422 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=1.995 $Y=3.44
+ $X2=2.087 $Y2=3.44
r85 10 11 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.995 $Y=3.44
+ $X2=1.82 $Y2=3.44
r86 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.745 $Y=3.515
+ $X2=1.82 $Y2=3.44
r87 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.745 $Y=3.515
+ $X2=1.745 $Y2=4.01
r88 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.39
+ $Y=0.235 $X2=1.53 $Y2=1.09
r89 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.39
+ $Y=0.235 $X2=1.53 $Y2=0.38
r90 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.39
+ $Y=2.23 $X2=1.53 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_123_718# 1 2 7 9 10 12 13 14 17 21
+ 25 29 35 37 40 41 44 45 46 48 49 51 54 56 57 61 65 66 79
c157 79 0 5.05501e-20 $X=6.24 $Y=5.03
c158 14 0 1.8723e-19 $X=2.18 $Y=5.275
c159 7 0 1.70849e-20 $X=1.745 $Y=5.35
r160 66 74 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.58 $Y=5.1
+ $X2=2.58 $Y2=5.275
r161 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=5.1 $X2=2.58 $Y2=5.1
r162 62 69 3.32414 $w=2.9e-07 $l=2e-08 $layer=POLY_cond $X=1.765 $Y=5.142
+ $X2=1.745 $Y2=5.142
r163 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=5.1 $X2=1.765 $Y2=5.1
r164 56 57 5.31505 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.75 $Y=5.57
+ $X2=0.75 $Y2=5.435
r165 52 79 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.97 $Y=5.03
+ $X2=6.24 $Y2=5.03
r166 52 76 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.97 $Y=5.03 $X2=5.88
+ $Y2=5.03
r167 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.97
+ $Y=5.03 $X2=5.97 $Y2=5.03
r168 49 51 50.8123 $w=3.28e-07 $l=1.455e-06 $layer=LI1_cond $X=4.515 $Y=5.03
+ $X2=5.97 $Y2=5.03
r169 47 49 7.68689 $w=3.3e-07 $l=2.04316e-07 $layer=LI1_cond $X=4.427 $Y=5.195
+ $X2=4.515 $Y2=5.03
r170 47 48 65.9117 $w=1.73e-07 $l=1.04e-06 $layer=LI1_cond $X=4.427 $Y=5.195
+ $X2=4.427 $Y2=6.235
r171 45 48 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=4.34 $Y=6.32
+ $X2=4.427 $Y2=6.235
r172 45 46 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.34 $Y=6.32
+ $X2=3.8 $Y2=6.32
r173 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.715 $Y=6.235
+ $X2=3.8 $Y2=6.32
r174 43 44 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.715 $Y=5.285
+ $X2=3.715 $Y2=6.235
r175 41 43 6.89401 $w=2.05e-07 $l=1.39155e-07 $layer=LI1_cond $X=3.63 $Y=5.182
+ $X2=3.715 $Y2=5.285
r176 41 65 52.2084 $w=2.03e-07 $l=9.65e-07 $layer=LI1_cond $X=3.63 $Y=5.182
+ $X2=2.665 $Y2=5.182
r177 40 61 10.1403 $w=1.73e-07 $l=1.6e-07 $layer=LI1_cond $X=1.605 $Y=5.097
+ $X2=1.765 $Y2=5.097
r178 39 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.605 $Y=4.82
+ $X2=1.605 $Y2=5.01
r179 38 54 3.01551 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.855 $Y=4.735
+ $X2=0.715 $Y2=4.735
r180 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.52 $Y=4.735
+ $X2=1.605 $Y2=4.82
r181 37 38 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.52 $Y=4.735
+ $X2=0.855 $Y2=4.735
r182 33 56 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.75 $Y=5.61 $X2=0.75
+ $Y2=5.57
r183 33 35 22.0611 $w=3.48e-07 $l=6.7e-07 $layer=LI1_cond $X=0.75 $Y=5.61
+ $X2=0.75 $Y2=6.28
r184 31 54 3.49088 $w=2.67e-07 $l=9.12688e-08 $layer=LI1_cond $X=0.702 $Y=4.82
+ $X2=0.715 $Y2=4.735
r185 31 57 27.7942 $w=2.53e-07 $l=6.15e-07 $layer=LI1_cond $X=0.702 $Y=4.82
+ $X2=0.702 $Y2=5.435
r186 27 54 3.49088 $w=2.67e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=4.65
+ $X2=0.715 $Y2=4.735
r187 27 29 37.0428 $w=2.78e-07 $l=9e-07 $layer=LI1_cond $X=0.715 $Y=4.65
+ $X2=0.715 $Y2=3.75
r188 23 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.24 $Y=5.195
+ $X2=6.24 $Y2=5.03
r189 23 25 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=6.24 $Y=5.195
+ $X2=6.24 $Y2=5.925
r190 19 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.24 $Y=4.865
+ $X2=6.24 $Y2=5.03
r191 19 21 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=6.24 $Y=4.865
+ $X2=6.24 $Y2=4.01
r192 15 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.88 $Y=5.195
+ $X2=5.88 $Y2=5.03
r193 15 17 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=5.88 $Y=5.195
+ $X2=5.88 $Y2=5.925
r194 13 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=5.275
+ $X2=2.58 $Y2=5.275
r195 13 14 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=2.415 $Y=5.275
+ $X2=2.18 $Y2=5.275
r196 10 14 23.6571 $w=2.9e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.105 $Y=5.35
+ $X2=2.18 $Y2=5.275
r197 10 62 56.5103 $w=2.9e-07 $l=4.31648e-07 $layer=POLY_cond $X=2.105 $Y=5.35
+ $X2=1.765 $Y2=5.142
r198 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.105 $Y=5.35
+ $X2=2.105 $Y2=5.925
r199 7 69 18.1727 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.745 $Y=5.35
+ $X2=1.745 $Y2=5.142
r200 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.745 $Y=5.35
+ $X2=1.745 $Y2=5.925
r201 2 56 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=5.425 $X2=0.74 $Y2=5.57
r202 2 35 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=5.425 $X2=0.74 $Y2=6.28
r203 1 29 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=3.59 $X2=0.74 $Y2=3.75
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%SLEEP 1 3 6 8 10 13 15 16 19 21 26
c67 1 0 1.58517e-19 $X=3.08 $Y=4.505
r68 27 28 9.29477 $w=3.63e-07 $l=7e-08 $layer=POLY_cond $X=3.44 $Y=4.687
+ $X2=3.51 $Y2=4.687
r69 25 27 24.5647 $w=3.63e-07 $l=1.85e-07 $layer=POLY_cond $X=3.255 $Y=4.687
+ $X2=3.44 $Y2=4.687
r70 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.255
+ $Y=4.705 $X2=3.255 $Y2=4.705
r71 23 25 23.2369 $w=3.63e-07 $l=1.75e-07 $layer=POLY_cond $X=3.08 $Y=4.687
+ $X2=3.255 $Y2=4.687
r72 21 26 3.84148 $w=4.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.12 $Y=4.707
+ $X2=3.255 $Y2=4.707
r73 17 19 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=3.87 $Y=4.655
+ $X2=3.87 $Y2=5.925
r74 16 28 27.0016 $w=3.63e-07 $l=1.39549e-07 $layer=POLY_cond $X=3.585 $Y=4.58
+ $X2=3.51 $Y2=4.687
r75 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.795 $Y=4.58
+ $X2=3.87 $Y2=4.655
r76 15 16 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.795 $Y=4.58
+ $X2=3.585 $Y2=4.58
r77 11 28 23.5056 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.51 $Y=4.87
+ $X2=3.51 $Y2=4.687
r78 11 13 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=3.51 $Y=4.87
+ $X2=3.51 $Y2=5.925
r79 8 27 23.5056 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=3.44 $Y=4.505
+ $X2=3.44 $Y2=4.687
r80 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.44 $Y=4.505 $X2=3.44
+ $Y2=4.22
r81 4 23 23.5056 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.08 $Y=4.87
+ $X2=3.08 $Y2=4.687
r82 4 6 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=3.08 $Y=4.87
+ $X2=3.08 $Y2=5.925
r83 1 23 23.5056 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=3.08 $Y=4.505
+ $X2=3.08 $Y2=4.687
r84 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.08 $Y=4.505 $X2=3.08
+ $Y2=4.22
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_517_420# 1 2 7 9 10 11 14 17 18 19
+ 22 24 28 30 32 34 35 36 37 38 39 41 45 53
r99 45 54 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.995 $Y=3.75
+ $X2=3.995 $Y2=3.84
r100 45 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=3.75
+ $X2=3.995 $Y2=3.585
r101 44 47 10.7413 $w=4.6e-07 $l=4.05e-07 $layer=LI1_cond $X=3.785 $Y=3.75
+ $X2=3.785 $Y2=4.155
r102 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.995
+ $Y=3.75 $X2=3.995 $Y2=3.75
r103 39 41 35.4909 $w=1.98e-07 $l=6.4e-07 $layer=LI1_cond $X=4.07 $Y=4.91
+ $X2=4.07 $Y2=5.55
r104 38 39 24.0086 $w=1.68e-07 $l=3.68e-07 $layer=LI1_cond $X=3.702 $Y=4.825
+ $X2=4.07 $Y2=4.825
r105 37 47 5.44365 $w=4.6e-07 $l=1.19499e-07 $layer=LI1_cond $X=3.702 $Y=4.24
+ $X2=3.785 $Y2=4.155
r106 37 38 25.6098 $w=2.23e-07 $l=5e-07 $layer=LI1_cond $X=3.702 $Y=4.24
+ $X2=3.702 $Y2=4.74
r107 32 34 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.88 $Y=4.505
+ $X2=5.88 $Y2=4.01
r108 31 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.525 $Y=4.58
+ $X2=5.45 $Y2=4.58
r109 30 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.805 $Y=4.58
+ $X2=5.88 $Y2=4.505
r110 30 31 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.805 $Y=4.58
+ $X2=5.525 $Y2=4.58
r111 26 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.45 $Y=4.655
+ $X2=5.45 $Y2=4.58
r112 26 28 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=5.45 $Y=4.655
+ $X2=5.45 $Y2=5.925
r113 25 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.165 $Y=4.58
+ $X2=5.09 $Y2=4.58
r114 24 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.375 $Y=4.58
+ $X2=5.45 $Y2=4.58
r115 24 25 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.375 $Y=4.58
+ $X2=5.165 $Y2=4.58
r116 20 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.09 $Y=4.655
+ $X2=5.09 $Y2=4.58
r117 20 22 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=5.09 $Y=4.655
+ $X2=5.09 $Y2=5.925
r118 18 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.015 $Y=4.58
+ $X2=5.09 $Y2=4.58
r119 18 19 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=5.015 $Y=4.58
+ $X2=4.67 $Y2=4.58
r120 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.595 $Y=4.505
+ $X2=4.67 $Y2=4.58
r121 16 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.595 $Y=3.915
+ $X2=4.595 $Y2=4.505
r122 15 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.16 $Y=3.84
+ $X2=3.995 $Y2=3.84
r123 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.52 $Y=3.84
+ $X2=4.595 $Y2=3.915
r124 14 15 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.52 $Y=3.84
+ $X2=4.16 $Y2=3.84
r125 12 53 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.905 $Y=3.295
+ $X2=3.905 $Y2=3.585
r126 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.83 $Y=3.22
+ $X2=3.905 $Y2=3.295
r127 10 11 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=3.83 $Y=3.22
+ $X2=2.735 $Y2=3.22
r128 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.66 $Y=3.145
+ $X2=2.735 $Y2=3.22
r129 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.66 $Y=3.145
+ $X2=2.66 $Y2=2.65
r130 2 41 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.945
+ $Y=5.425 $X2=4.085 $Y2=5.55
r131 1 47 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=4.01 $X2=3.655 $Y2=4.155
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%VPWR 1 6 10 12 22 23 26 33
r24 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r25 22 23 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r26 20 33 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.36
+ $Y2=0
r27 20 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r28 19 22 375.786 $w=1.68e-07 $l=5.76e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=6.96
+ $Y2=0
r29 19 20 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r30 17 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.74
+ $Y2=0
r31 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.2
+ $Y2=0
r32 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r33 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r34 12 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.74
+ $Y2=0
r35 12 14 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.24
+ $Y2=0
r36 10 23 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=6.96
+ $Y2=0
r37 10 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.36
+ $Y2=0
r38 6 8 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.74 $Y=0.38 $X2=0.74
+ $Y2=1.09
r39 4 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0
r40 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.38
r41 1 8 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.74 $Y2=1.09
r42 1 6 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.74 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_278_1085# 1 2 9 11 12 13 15
r35 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=6.235
+ $X2=2.865 $Y2=6.32
r36 13 15 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.865 $Y=6.235
+ $X2=2.865 $Y2=5.6
r37 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=6.32
+ $X2=2.865 $Y2=6.32
r38 11 12 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=2.7 $Y=6.32
+ $X2=1.695 $Y2=6.32
r39 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.53 $Y=6.235
+ $X2=1.695 $Y2=6.32
r40 7 9 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.53 $Y=6.235
+ $X2=1.53 $Y2=5.78
r41 2 18 400 $w=1.7e-07 $l=9.17701e-07 $layer=licon1_PDIFF $count=1 $X=2.735
+ $Y=5.425 $X2=2.865 $Y2=6.28
r42 2 15 400 $w=1.7e-07 $l=2.3103e-07 $layer=licon1_PDIFF $count=1 $X=2.735
+ $Y=5.425 $X2=2.865 $Y2=5.6
r43 1 9 300 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=2 $X=1.39
+ $Y=5.425 $X2=1.53 $Y2=5.78
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%DESTPWR 1 2 9 15 18 19 20 29 38 39 42
+ 48
r74 42 43 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=6.66
+ $X2=5.52 $Y2=6.66
r75 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=6.66
+ $X2=6.96 $Y2=6.66
r76 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=6.66 $X2=6.96
+ $Y2=6.66
r77 36 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=6.66 $X2=5.52
+ $Y2=6.66
r78 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=6.66 $X2=6.96
+ $Y2=6.66
r79 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=6.66 $X2=6
+ $Y2=6.66
r80 33 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.83 $Y=6.66
+ $X2=5.665 $Y2=6.66
r81 33 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.83 $Y=6.66 $X2=6
+ $Y2=6.66
r82 29 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.5 $Y=6.66
+ $X2=5.665 $Y2=6.66
r83 29 31 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=5.5 $Y=6.66 $X2=3.6
+ $Y2=6.66
r84 28 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.12 $Y=6.66
+ $X2=3.36 $Y2=6.66
r85 27 28 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=6.66
+ $X2=3.12 $Y2=6.66
r86 24 28 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=0.24 $Y=6.66
+ $X2=3.12 $Y2=6.66
r87 23 27 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=6.66
+ $X2=3.12 $Y2=6.66
r88 23 24 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=6.66
+ $X2=0.24 $Y2=6.66
r89 20 43 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=6.66
+ $X2=5.52 $Y2=6.66
r90 20 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.6 $Y=6.66
+ $X2=3.36 $Y2=6.66
r91 20 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=6.66
+ $X2=3.6 $Y2=6.66
r92 18 27 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.21 $Y=6.66 $X2=3.12
+ $Y2=6.66
r93 18 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=6.66
+ $X2=3.295 $Y2=6.66
r94 17 31 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.38 $Y=6.66 $X2=3.6
+ $Y2=6.66
r95 17 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.38 $Y=6.66
+ $X2=3.295 $Y2=6.66
r96 13 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.665 $Y=6.575
+ $X2=5.665 $Y2=6.66
r97 13 15 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=5.665 $Y=6.575
+ $X2=5.665 $Y2=5.925
r98 9 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.295 $Y=5.62
+ $X2=3.295 $Y2=6.3
r99 7 19 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=6.575
+ $X2=3.295 $Y2=6.66
r100 7 12 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.295 $Y=6.575
+ $X2=3.295 $Y2=6.3
r101 2 15 300 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=2 $X=5.525
+ $Y=5.425 $X2=5.665 $Y2=5.925
r102 1 12 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=5.425 $X2=3.295 $Y2=6.3
r103 1 9 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=5.425 $X2=3.295 $Y2=5.62
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%X 1 2 3 10 12 14 18 19 20 21 22 23 24
+ 35 47
r47 33 47 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=6.455 $Y=5.42
+ $X2=6.455 $Y2=5.365
r48 24 54 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=6.455 $Y=6.105
+ $X2=6.455 $Y2=6.28
r49 23 24 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.455 $Y=5.735
+ $X2=6.455 $Y2=6.105
r50 23 48 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.455 $Y=5.735
+ $X2=6.455 $Y2=5.59
r51 22 33 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=5.505
+ $X2=6.455 $Y2=5.42
r52 22 48 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=5.505
+ $X2=6.455 $Y2=5.59
r53 22 47 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.455 $Y=5.35
+ $X2=6.455 $Y2=5.365
r54 21 22 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=6.455 $Y=4.995
+ $X2=6.455 $Y2=5.35
r55 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.455 $Y=4.625
+ $X2=6.455 $Y2=4.995
r56 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.455 $Y=4.255
+ $X2=6.455 $Y2=4.625
r57 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.455 $Y=3.885
+ $X2=6.455 $Y2=4.255
r58 18 35 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.455 $Y=3.885
+ $X2=6.455 $Y2=3.735
r59 15 17 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.04 $Y=5.505
+ $X2=4.875 $Y2=5.505
r60 14 22 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.29 $Y=5.505
+ $X2=6.455 $Y2=5.505
r61 14 15 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=6.29 $Y=5.505
+ $X2=5.04 $Y2=5.505
r62 10 17 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=5.59
+ $X2=4.875 $Y2=5.505
r63 10 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.875 $Y=5.59
+ $X2=4.875 $Y2=6.3
r64 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.315
+ $Y=5.425 $X2=6.455 $Y2=5.57
r65 3 54 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.315
+ $Y=5.425 $X2=6.455 $Y2=6.28
r66 2 17 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=4.73
+ $Y=5.425 $X2=4.875 $Y2=5.585
r67 2 12 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=4.73
+ $Y=5.425 $X2=4.875 $Y2=6.3
r68 1 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.315
+ $Y=3.59 $X2=6.455 $Y2=3.735
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_278_718# 1 2 9 13 16 18 19
c38 18 0 1.8723e-19 $X=1.53 $Y=3.75
r39 16 19 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.4 $Y=3.585
+ $X2=2.4 $Y2=3.09
r40 11 19 6.27261 $w=2.13e-07 $l=1.07e-07 $layer=LI1_cond $X=2.422 $Y=2.983
+ $X2=2.422 $Y2=3.09
r41 11 13 26.1578 $w=2.13e-07 $l=4.88e-07 $layer=LI1_cond $X=2.422 $Y=2.983
+ $X2=2.422 $Y2=2.495
r42 10 18 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.645 $Y=3.67
+ $X2=1.505 $Y2=3.67
r43 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.315 $Y=3.67
+ $X2=2.4 $Y2=3.585
r44 9 10 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.315 $Y=3.67
+ $X2=1.645 $Y2=3.67
r45 2 13 91 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=2 $X=2.32
+ $Y=2.23 $X2=2.445 $Y2=2.495
r46 1 18 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=1.39
+ $Y=3.59 $X2=1.53 $Y2=3.75
.ends

