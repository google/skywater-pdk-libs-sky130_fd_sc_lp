* File: sky130_fd_sc_lp__einvn_8.pxi.spice
* Created: Fri Aug 28 10:33:04 2020
* 
x_PM_SKY130_FD_SC_LP__EINVN_8%A_110_57# N_A_110_57#_M1023_d N_A_110_57#_M1010_d
+ N_A_110_57#_c_159_n N_A_110_57#_c_160_n N_A_110_57#_c_161_n
+ N_A_110_57#_M1004_g N_A_110_57#_c_162_n N_A_110_57#_c_163_n
+ N_A_110_57#_M1012_g N_A_110_57#_c_164_n N_A_110_57#_c_165_n
+ N_A_110_57#_M1014_g N_A_110_57#_c_166_n N_A_110_57#_c_167_n
+ N_A_110_57#_M1016_g N_A_110_57#_c_168_n N_A_110_57#_c_169_n
+ N_A_110_57#_M1026_g N_A_110_57#_c_170_n N_A_110_57#_c_171_n
+ N_A_110_57#_M1027_g N_A_110_57#_c_172_n N_A_110_57#_c_173_n
+ N_A_110_57#_M1028_g N_A_110_57#_c_174_n N_A_110_57#_c_175_n
+ N_A_110_57#_M1033_g N_A_110_57#_c_176_n N_A_110_57#_c_177_n
+ N_A_110_57#_c_178_n N_A_110_57#_c_179_n N_A_110_57#_c_180_n
+ N_A_110_57#_c_181_n N_A_110_57#_c_182_n N_A_110_57#_c_183_n
+ N_A_110_57#_c_184_n N_A_110_57#_c_185_n N_A_110_57#_c_186_n
+ PM_SKY130_FD_SC_LP__EINVN_8%A_110_57#
x_PM_SKY130_FD_SC_LP__EINVN_8%TE_B N_TE_B_M1023_g N_TE_B_c_319_n N_TE_B_M1010_g
+ N_TE_B_c_302_n N_TE_B_c_303_n N_TE_B_c_322_n N_TE_B_M1001_g N_TE_B_c_304_n
+ N_TE_B_c_324_n N_TE_B_M1006_g N_TE_B_c_305_n N_TE_B_c_326_n N_TE_B_M1011_g
+ N_TE_B_c_306_n N_TE_B_c_328_n N_TE_B_M1018_g N_TE_B_c_307_n N_TE_B_c_330_n
+ N_TE_B_M1022_g N_TE_B_c_308_n N_TE_B_c_332_n N_TE_B_M1024_g N_TE_B_c_309_n
+ N_TE_B_c_334_n N_TE_B_M1025_g N_TE_B_c_310_n N_TE_B_c_336_n N_TE_B_M1030_g
+ N_TE_B_c_311_n N_TE_B_c_312_n N_TE_B_c_313_n N_TE_B_c_314_n N_TE_B_c_315_n
+ N_TE_B_c_316_n N_TE_B_c_317_n TE_B TE_B TE_B TE_B N_TE_B_c_318_n TE_B
+ PM_SKY130_FD_SC_LP__EINVN_8%TE_B
x_PM_SKY130_FD_SC_LP__EINVN_8%A N_A_c_461_n N_A_M1000_g N_A_M1003_g N_A_c_463_n
+ N_A_M1002_g N_A_M1007_g N_A_c_465_n N_A_M1005_g N_A_M1008_g N_A_c_467_n
+ N_A_M1013_g N_A_M1009_g N_A_c_469_n N_A_M1015_g N_A_M1020_g N_A_c_471_n
+ N_A_M1017_g N_A_M1021_g N_A_c_473_n N_A_M1019_g N_A_M1029_g N_A_c_475_n
+ N_A_M1032_g N_A_M1031_g A A N_A_c_477_n PM_SKY130_FD_SC_LP__EINVN_8%A
x_PM_SKY130_FD_SC_LP__EINVN_8%VPWR N_VPWR_M1010_s N_VPWR_M1001_d N_VPWR_M1011_d
+ N_VPWR_M1022_d N_VPWR_M1025_d N_VPWR_c_602_n N_VPWR_c_603_n N_VPWR_c_604_n
+ N_VPWR_c_605_n N_VPWR_c_606_n N_VPWR_c_607_n N_VPWR_c_608_n N_VPWR_c_609_n
+ N_VPWR_c_610_n N_VPWR_c_611_n VPWR N_VPWR_c_612_n N_VPWR_c_613_n
+ N_VPWR_c_614_n N_VPWR_c_601_n N_VPWR_c_616_n N_VPWR_c_617_n N_VPWR_c_618_n
+ PM_SKY130_FD_SC_LP__EINVN_8%VPWR
x_PM_SKY130_FD_SC_LP__EINVN_8%A_305_367# N_A_305_367#_M1001_s
+ N_A_305_367#_M1006_s N_A_305_367#_M1018_s N_A_305_367#_M1024_s
+ N_A_305_367#_M1030_s N_A_305_367#_M1007_d N_A_305_367#_M1009_d
+ N_A_305_367#_M1021_d N_A_305_367#_M1031_d N_A_305_367#_c_729_n
+ N_A_305_367#_c_735_n N_A_305_367#_c_730_n N_A_305_367#_c_797_n
+ N_A_305_367#_c_737_n N_A_305_367#_c_801_n N_A_305_367#_c_738_n
+ N_A_305_367#_c_805_n N_A_305_367#_c_731_n N_A_305_367#_c_809_n
+ N_A_305_367#_c_773_n N_A_305_367#_c_833_p N_A_305_367#_c_775_n
+ N_A_305_367#_c_777_n N_A_305_367#_c_778_n N_A_305_367#_c_780_n
+ N_A_305_367#_c_781_n N_A_305_367#_c_732_n N_A_305_367#_c_733_n
+ N_A_305_367#_c_769_n N_A_305_367#_c_770_n N_A_305_367#_c_771_n
+ N_A_305_367#_c_821_n N_A_305_367#_c_823_n N_A_305_367#_c_825_n
+ PM_SKY130_FD_SC_LP__EINVN_8%A_305_367#
x_PM_SKY130_FD_SC_LP__EINVN_8%Z N_Z_M1000_s N_Z_M1005_s N_Z_M1015_s N_Z_M1019_s
+ N_Z_M1003_s N_Z_M1008_s N_Z_M1020_s N_Z_M1029_s N_Z_c_864_n N_Z_c_861_n
+ N_Z_c_862_n N_Z_c_878_n N_Z_c_882_n N_Z_c_858_n N_Z_c_888_n N_Z_c_859_n Z Z Z
+ Z Z Z N_Z_c_860_n PM_SKY130_FD_SC_LP__EINVN_8%Z
x_PM_SKY130_FD_SC_LP__EINVN_8%VGND N_VGND_M1023_s N_VGND_M1004_d N_VGND_M1014_d
+ N_VGND_M1026_d N_VGND_M1028_d N_VGND_c_943_n N_VGND_c_944_n N_VGND_c_945_n
+ N_VGND_c_946_n N_VGND_c_947_n N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n
+ N_VGND_c_951_n N_VGND_c_952_n N_VGND_c_953_n N_VGND_c_954_n N_VGND_c_955_n
+ VGND N_VGND_c_956_n N_VGND_c_957_n N_VGND_c_958_n
+ PM_SKY130_FD_SC_LP__EINVN_8%VGND
x_PM_SKY130_FD_SC_LP__EINVN_8%A_305_47# N_A_305_47#_M1004_s N_A_305_47#_M1012_s
+ N_A_305_47#_M1016_s N_A_305_47#_M1027_s N_A_305_47#_M1033_s
+ N_A_305_47#_M1002_d N_A_305_47#_M1013_d N_A_305_47#_M1017_d
+ N_A_305_47#_M1032_d N_A_305_47#_c_1060_n N_A_305_47#_c_1061_n
+ N_A_305_47#_c_1062_n N_A_305_47#_c_1063_n N_A_305_47#_c_1064_n
+ N_A_305_47#_c_1065_n N_A_305_47#_c_1066_n N_A_305_47#_c_1067_n
+ N_A_305_47#_c_1068_n N_A_305_47#_c_1200_n N_A_305_47#_c_1069_n
+ N_A_305_47#_c_1125_n N_A_305_47#_c_1130_n N_A_305_47#_c_1070_n
+ N_A_305_47#_c_1071_n N_A_305_47#_c_1072_n N_A_305_47#_c_1073_n
+ N_A_305_47#_c_1074_n N_A_305_47#_c_1135_n N_A_305_47#_c_1140_n
+ PM_SKY130_FD_SC_LP__EINVN_8%A_305_47#
cc_1 VNB N_A_110_57#_c_159_n 0.0239185f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.265
cc_2 VNB N_A_110_57#_c_160_n 0.0125595f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.265
cc_3 VNB N_A_110_57#_c_161_n 0.019504f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.185
cc_4 VNB N_A_110_57#_c_162_n 0.00969604f $X=-0.19 $Y=-0.245 $X2=2.22 $Y2=1.265
cc_5 VNB N_A_110_57#_c_163_n 0.0161528f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.185
cc_6 VNB N_A_110_57#_c_164_n 0.0103904f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.265
cc_7 VNB N_A_110_57#_c_165_n 0.0161528f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.185
cc_8 VNB N_A_110_57#_c_166_n 0.00969604f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.265
cc_9 VNB N_A_110_57#_c_167_n 0.0161528f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=1.185
cc_10 VNB N_A_110_57#_c_168_n 0.0103904f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.265
cc_11 VNB N_A_110_57#_c_169_n 0.0161528f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.185
cc_12 VNB N_A_110_57#_c_170_n 0.00969604f $X=-0.19 $Y=-0.245 $X2=3.94 $Y2=1.265
cc_13 VNB N_A_110_57#_c_171_n 0.0161528f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=1.185
cc_14 VNB N_A_110_57#_c_172_n 0.0103904f $X=-0.19 $Y=-0.245 $X2=4.37 $Y2=1.265
cc_15 VNB N_A_110_57#_c_173_n 0.0161528f $X=-0.19 $Y=-0.245 $X2=4.445 $Y2=1.185
cc_16 VNB N_A_110_57#_c_174_n 0.0164987f $X=-0.19 $Y=-0.245 $X2=4.8 $Y2=1.265
cc_17 VNB N_A_110_57#_c_175_n 0.0163877f $X=-0.19 $Y=-0.245 $X2=4.875 $Y2=1.185
cc_18 VNB N_A_110_57#_c_176_n 0.00406978f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.265
cc_19 VNB N_A_110_57#_c_177_n 0.00406978f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.265
cc_20 VNB N_A_110_57#_c_178_n 0.00406978f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.265
cc_21 VNB N_A_110_57#_c_179_n 0.00406978f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=1.265
cc_22 VNB N_A_110_57#_c_180_n 0.00406978f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.265
cc_23 VNB N_A_110_57#_c_181_n 0.00406978f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=1.265
cc_24 VNB N_A_110_57#_c_182_n 0.00406978f $X=-0.19 $Y=-0.245 $X2=4.445 $Y2=1.265
cc_25 VNB N_A_110_57#_c_183_n 0.00250006f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.43
cc_26 VNB N_A_110_57#_c_184_n 0.004735f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.98
cc_27 VNB N_A_110_57#_c_185_n 0.0074406f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.83
cc_28 VNB N_A_110_57#_c_186_n 0.0509946f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.83
cc_29 VNB N_TE_B_M1023_g 0.0282184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_TE_B_c_302_n 0.0195562f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.265
cc_31 VNB N_TE_B_c_303_n 0.0665148f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.185
cc_32 VNB N_TE_B_c_304_n 0.00757833f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.265
cc_33 VNB N_TE_B_c_305_n 0.00757827f $X=-0.19 $Y=-0.245 $X2=2.37 $Y2=1.265
cc_34 VNB N_TE_B_c_306_n 0.00757833f $X=-0.19 $Y=-0.245 $X2=2.8 $Y2=1.265
cc_35 VNB N_TE_B_c_307_n 0.00757827f $X=-0.19 $Y=-0.245 $X2=3.23 $Y2=1.265
cc_36 VNB N_TE_B_c_308_n 0.00757833f $X=-0.19 $Y=-0.245 $X2=3.66 $Y2=1.265
cc_37 VNB N_TE_B_c_309_n 0.00757827f $X=-0.19 $Y=-0.245 $X2=4.09 $Y2=1.265
cc_38 VNB N_TE_B_c_310_n 0.0137088f $X=-0.19 $Y=-0.245 $X2=4.52 $Y2=1.265
cc_39 VNB N_TE_B_c_311_n 0.00412531f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.265
cc_40 VNB N_TE_B_c_312_n 0.00412531f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.265
cc_41 VNB N_TE_B_c_313_n 0.00412531f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.265
cc_42 VNB N_TE_B_c_314_n 0.00412531f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=1.265
cc_43 VNB N_TE_B_c_315_n 0.00412531f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.265
cc_44 VNB N_TE_B_c_316_n 0.00412531f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=1.265
cc_45 VNB N_TE_B_c_317_n 0.00412531f $X=-0.19 $Y=-0.245 $X2=4.445 $Y2=1.265
cc_46 VNB N_TE_B_c_318_n 0.0268092f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.83
cc_47 VNB N_A_c_461_n 0.0164056f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.285
cc_48 VNB N_A_M1003_g 0.00839416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_c_463_n 0.016196f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.265
cc_50 VNB N_A_M1007_g 0.00706341f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.265
cc_51 VNB N_A_c_465_n 0.0161714f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=0.655
cc_52 VNB N_A_M1008_g 0.00702562f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.655
cc_53 VNB N_A_c_467_n 0.0158137f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.265
cc_54 VNB N_A_M1009_g 0.00590672f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.265
cc_55 VNB N_A_c_469_n 0.0158137f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.185
cc_56 VNB N_A_M1020_g 0.00590672f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=1.185
cc_57 VNB N_A_c_471_n 0.0158138f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=0.655
cc_58 VNB N_A_M1021_g 0.00590672f $X=-0.19 $Y=-0.245 $X2=4.445 $Y2=0.655
cc_59 VNB N_A_c_473_n 0.0158138f $X=-0.19 $Y=-0.245 $X2=4.52 $Y2=1.265
cc_60 VNB N_A_M1029_g 0.00590672f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.265
cc_61 VNB N_A_c_475_n 0.0215271f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.265
cc_62 VNB N_A_M1031_g 0.0111406f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.665
cc_63 VNB N_A_c_477_n 0.174854f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.83
cc_64 VNB N_VPWR_c_601_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_Z_c_858_n 0.00108157f $X=-0.19 $Y=-0.245 $X2=4.875 $Y2=0.655
cc_66 VNB N_Z_c_859_n 0.00106072f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=1.265
cc_67 VNB N_Z_c_860_n 0.0103654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_943_n 0.0109056f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=0.655
cc_69 VNB N_VGND_c_944_n 0.0374186f $X=-0.19 $Y=-0.245 $X2=2.37 $Y2=1.265
cc_70 VNB N_VGND_c_945_n 0.00705838f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.265
cc_71 VNB N_VGND_c_946_n 0.00645267f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=0.655
cc_72 VNB N_VGND_c_947_n 0.00645267f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=0.655
cc_73 VNB N_VGND_c_948_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=3.94 $Y2=1.265
cc_74 VNB N_VGND_c_949_n 0.00706729f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=0.655
cc_75 VNB N_VGND_c_950_n 0.0427099f $X=-0.19 $Y=-0.245 $X2=4.445 $Y2=1.185
cc_76 VNB N_VGND_c_951_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.445 $Y2=0.655
cc_77 VNB N_VGND_c_952_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=4.8 $Y2=1.265
cc_78 VNB N_VGND_c_953_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.52 $Y2=1.265
cc_79 VNB N_VGND_c_954_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=4.875 $Y2=1.185
cc_80 VNB N_VGND_c_955_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.875 $Y2=0.655
cc_81 VNB N_VGND_c_956_n 0.10375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_957_n 0.458514f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.875
cc_83 VNB N_VGND_c_958_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_305_47#_c_1060_n 0.0202326f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=0.655
cc_85 VNB N_A_305_47#_c_1061_n 0.00347392f $X=-0.19 $Y=-0.245 $X2=3.94 $Y2=1.265
cc_86 VNB N_A_305_47#_c_1062_n 0.00324387f $X=-0.19 $Y=-0.245 $X2=3.66 $Y2=1.265
cc_87 VNB N_A_305_47#_c_1063_n 0.00158555f $X=-0.19 $Y=-0.245 $X2=4.015
+ $Y2=0.655
cc_88 VNB N_A_305_47#_c_1064_n 0.00347392f $X=-0.19 $Y=-0.245 $X2=4.09 $Y2=1.265
cc_89 VNB N_A_305_47#_c_1065_n 0.00158555f $X=-0.19 $Y=-0.245 $X2=4.8 $Y2=1.265
cc_90 VNB N_A_305_47#_c_1066_n 0.00347392f $X=-0.19 $Y=-0.245 $X2=4.875
+ $Y2=1.185
cc_91 VNB N_A_305_47#_c_1067_n 0.00158555f $X=-0.19 $Y=-0.245 $X2=1.865
+ $Y2=1.265
cc_92 VNB N_A_305_47#_c_1068_n 0.00759676f $X=-0.19 $Y=-0.245 $X2=2.725
+ $Y2=1.265
cc_93 VNB N_A_305_47#_c_1069_n 0.00372355f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.665
cc_94 VNB N_A_305_47#_c_1070_n 0.00746637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_305_47#_c_1071_n 0.0380389f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.83
cc_96 VNB N_A_305_47#_c_1072_n 0.00153519f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.83
cc_97 VNB N_A_305_47#_c_1073_n 0.00153519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_305_47#_c_1074_n 0.00153519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VPB N_A_110_57#_c_184_n 0.0126369f $X=-0.19 $Y=1.655 $X2=1.13 $Y2=1.98
cc_100 VPB N_TE_B_c_319_n 0.023589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_TE_B_c_302_n 0.0269392f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=1.265
cc_102 VPB N_TE_B_c_303_n 0.0358014f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=1.185
cc_103 VPB N_TE_B_c_322_n 0.019358f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=0.655
cc_104 VPB N_TE_B_c_304_n 0.0049284f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=1.265
cc_105 VPB N_TE_B_c_324_n 0.0150524f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=0.655
cc_106 VPB N_TE_B_c_305_n 0.0049284f $X=-0.19 $Y=1.655 $X2=2.37 $Y2=1.265
cc_107 VPB N_TE_B_c_326_n 0.0150524f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=0.655
cc_108 VPB N_TE_B_c_306_n 0.0049284f $X=-0.19 $Y=1.655 $X2=2.8 $Y2=1.265
cc_109 VPB N_TE_B_c_328_n 0.0150524f $X=-0.19 $Y=1.655 $X2=3.155 $Y2=0.655
cc_110 VPB N_TE_B_c_307_n 0.0049284f $X=-0.19 $Y=1.655 $X2=3.23 $Y2=1.265
cc_111 VPB N_TE_B_c_330_n 0.0150524f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=0.655
cc_112 VPB N_TE_B_c_308_n 0.0049284f $X=-0.19 $Y=1.655 $X2=3.66 $Y2=1.265
cc_113 VPB N_TE_B_c_332_n 0.0150524f $X=-0.19 $Y=1.655 $X2=4.015 $Y2=0.655
cc_114 VPB N_TE_B_c_309_n 0.0049284f $X=-0.19 $Y=1.655 $X2=4.09 $Y2=1.265
cc_115 VPB N_TE_B_c_334_n 0.0150524f $X=-0.19 $Y=1.655 $X2=4.445 $Y2=0.655
cc_116 VPB N_TE_B_c_310_n 0.00711562f $X=-0.19 $Y=1.655 $X2=4.52 $Y2=1.265
cc_117 VPB N_TE_B_c_336_n 0.0151133f $X=-0.19 $Y=1.655 $X2=4.875 $Y2=0.655
cc_118 VPB N_TE_B_c_311_n 0.00111435f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=1.265
cc_119 VPB N_TE_B_c_312_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.265
cc_120 VPB N_TE_B_c_313_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=1.265
cc_121 VPB N_TE_B_c_314_n 0.00111435f $X=-0.19 $Y=1.655 $X2=3.155 $Y2=1.265
cc_122 VPB N_TE_B_c_315_n 0.00111435f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=1.265
cc_123 VPB N_TE_B_c_316_n 0.00111435f $X=-0.19 $Y=1.655 $X2=4.015 $Y2=1.265
cc_124 VPB N_TE_B_c_317_n 0.00111435f $X=-0.19 $Y=1.655 $X2=4.445 $Y2=1.265
cc_125 VPB TE_B 0.0695331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_M1003_g 0.019476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_M1007_g 0.0185045f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=1.265
cc_128 VPB N_A_M1008_g 0.0185143f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=0.655
cc_129 VPB N_A_M1009_g 0.0182686f $X=-0.19 $Y=1.655 $X2=3.51 $Y2=1.265
cc_130 VPB N_A_M1020_g 0.0182686f $X=-0.19 $Y=1.655 $X2=4.015 $Y2=1.185
cc_131 VPB N_A_M1021_g 0.0182686f $X=-0.19 $Y=1.655 $X2=4.445 $Y2=0.655
cc_132 VPB N_A_M1029_g 0.0182686f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=1.265
cc_133 VPB N_A_M1031_g 0.0268065f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.665
cc_134 VPB N_VPWR_c_602_n 0.00672171f $X=-0.19 $Y=1.655 $X2=2.37 $Y2=1.265
cc_135 VPB N_VPWR_c_603_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=3.155 $Y2=1.185
cc_136 VPB N_VPWR_c_604_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=3.585 $Y2=0.655
cc_137 VPB N_VPWR_c_605_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=4.015 $Y2=0.655
cc_138 VPB N_VPWR_c_606_n 0.0129398f $X=-0.19 $Y=1.655 $X2=4.445 $Y2=0.655
cc_139 VPB N_VPWR_c_607_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=4.875 $Y2=1.185
cc_140 VPB N_VPWR_c_608_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.265
cc_141 VPB N_VPWR_c_609_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=1.265
cc_142 VPB N_VPWR_c_610_n 0.0129398f $X=-0.19 $Y=1.655 $X2=3.155 $Y2=1.265
cc_143 VPB N_VPWR_c_611_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=1.265
cc_144 VPB N_VPWR_c_612_n 0.0187638f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.665
cc_145 VPB N_VPWR_c_613_n 0.0285647f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.98
cc_146 VPB N_VPWR_c_614_n 0.101972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_601_n 0.0767562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_616_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_617_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_618_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_305_367#_c_729_n 0.0102152f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=0.655
cc_152 VPB N_A_305_367#_c_730_n 0.00149049f $X=-0.19 $Y=1.655 $X2=4.015
+ $Y2=0.655
cc_153 VPB N_A_305_367#_c_731_n 0.0034393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_305_367#_c_732_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_305_367#_c_733_n 0.0512487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_Z_c_861_n 0.00225871f $X=-0.19 $Y=1.655 $X2=3.66 $Y2=1.265
cc_157 VPB N_Z_c_862_n 0.00230427f $X=-0.19 $Y=1.655 $X2=4.015 $Y2=1.185
cc_158 VPB N_Z_c_860_n 0.00202898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 N_A_110_57#_c_183_n N_TE_B_M1023_g 0.00124045f $X=0.69 $Y=0.43 $X2=0
+ $Y2=0
cc_160 N_A_110_57#_c_184_n N_TE_B_M1023_g 9.42755e-19 $X=1.13 $Y=1.98 $X2=0
+ $Y2=0
cc_161 N_A_110_57#_c_186_n N_TE_B_M1023_g 0.0116695f $X=1.15 $Y=0.83 $X2=0 $Y2=0
cc_162 N_A_110_57#_c_184_n N_TE_B_c_319_n 0.0189977f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_163 N_A_110_57#_c_159_n N_TE_B_c_302_n 0.0158549f $X=1.79 $Y=1.265 $X2=0
+ $Y2=0
cc_164 N_A_110_57#_c_184_n N_TE_B_c_302_n 0.0201767f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_165 N_A_110_57#_c_160_n N_TE_B_c_303_n 0.0192026f $X=1.315 $Y=1.265 $X2=0
+ $Y2=0
cc_166 N_A_110_57#_c_184_n N_TE_B_c_303_n 0.00520013f $X=1.13 $Y=1.98 $X2=0
+ $Y2=0
cc_167 N_A_110_57#_c_185_n N_TE_B_c_303_n 0.0074479f $X=1.15 $Y=0.83 $X2=0 $Y2=0
cc_168 N_A_110_57#_c_184_n N_TE_B_c_322_n 5.51926e-19 $X=1.13 $Y=1.98 $X2=0
+ $Y2=0
cc_169 N_A_110_57#_c_162_n N_TE_B_c_304_n 0.0158549f $X=2.22 $Y=1.265 $X2=0
+ $Y2=0
cc_170 N_A_110_57#_c_164_n N_TE_B_c_305_n 0.0158549f $X=2.65 $Y=1.265 $X2=0
+ $Y2=0
cc_171 N_A_110_57#_c_166_n N_TE_B_c_306_n 0.0158549f $X=3.08 $Y=1.265 $X2=0
+ $Y2=0
cc_172 N_A_110_57#_c_168_n N_TE_B_c_307_n 0.0158549f $X=3.51 $Y=1.265 $X2=0
+ $Y2=0
cc_173 N_A_110_57#_c_170_n N_TE_B_c_308_n 0.0158549f $X=3.94 $Y=1.265 $X2=0
+ $Y2=0
cc_174 N_A_110_57#_c_172_n N_TE_B_c_309_n 0.0158549f $X=4.37 $Y=1.265 $X2=0
+ $Y2=0
cc_175 N_A_110_57#_c_174_n N_TE_B_c_310_n 0.0158549f $X=4.8 $Y=1.265 $X2=0 $Y2=0
cc_176 N_A_110_57#_c_176_n N_TE_B_c_311_n 0.0158549f $X=1.865 $Y=1.265 $X2=0
+ $Y2=0
cc_177 N_A_110_57#_c_177_n N_TE_B_c_312_n 0.0158549f $X=2.295 $Y=1.265 $X2=0
+ $Y2=0
cc_178 N_A_110_57#_c_178_n N_TE_B_c_313_n 0.0158549f $X=2.725 $Y=1.265 $X2=0
+ $Y2=0
cc_179 N_A_110_57#_c_179_n N_TE_B_c_314_n 0.0158549f $X=3.155 $Y=1.265 $X2=0
+ $Y2=0
cc_180 N_A_110_57#_c_180_n N_TE_B_c_315_n 0.0158549f $X=3.585 $Y=1.265 $X2=0
+ $Y2=0
cc_181 N_A_110_57#_c_181_n N_TE_B_c_316_n 0.0158549f $X=4.015 $Y=1.265 $X2=0
+ $Y2=0
cc_182 N_A_110_57#_c_182_n N_TE_B_c_317_n 0.0158549f $X=4.445 $Y=1.265 $X2=0
+ $Y2=0
cc_183 N_A_110_57#_c_160_n N_TE_B_c_318_n 0.001031f $X=1.315 $Y=1.265 $X2=0
+ $Y2=0
cc_184 N_A_110_57#_c_184_n N_TE_B_c_318_n 0.0303969f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_185 N_A_110_57#_c_185_n N_TE_B_c_318_n 0.0151152f $X=1.15 $Y=0.83 $X2=0 $Y2=0
cc_186 N_A_110_57#_c_184_n TE_B 0.00503842f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_187 N_A_110_57#_c_175_n N_A_c_461_n 0.0111703f $X=4.875 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_110_57#_c_174_n N_A_c_477_n 0.0111703f $X=4.8 $Y=1.265 $X2=0 $Y2=0
cc_189 N_A_110_57#_c_184_n N_VPWR_c_602_n 0.045869f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_190 N_A_110_57#_c_184_n N_VPWR_c_613_n 0.021117f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_191 N_A_110_57#_M1010_d N_VPWR_c_601_n 0.00215158f $X=0.99 $Y=1.835 $X2=0
+ $Y2=0
cc_192 N_A_110_57#_c_184_n N_VPWR_c_601_n 0.0126604f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_193 N_A_110_57#_c_184_n N_A_305_367#_c_729_n 0.0940211f $X=1.13 $Y=1.98 $X2=0
+ $Y2=0
cc_194 N_A_110_57#_c_159_n N_A_305_367#_c_735_n 5.15742e-19 $X=1.79 $Y=1.265
+ $X2=0 $Y2=0
cc_195 N_A_110_57#_c_184_n N_A_305_367#_c_730_n 0.0216832f $X=1.13 $Y=1.98 $X2=0
+ $Y2=0
cc_196 N_A_110_57#_c_164_n N_A_305_367#_c_737_n 5.15742e-19 $X=2.65 $Y=1.265
+ $X2=0 $Y2=0
cc_197 N_A_110_57#_c_168_n N_A_305_367#_c_738_n 5.15742e-19 $X=3.51 $Y=1.265
+ $X2=0 $Y2=0
cc_198 N_A_110_57#_c_172_n N_A_305_367#_c_731_n 4.80142e-19 $X=4.37 $Y=1.265
+ $X2=0 $Y2=0
cc_199 N_A_110_57#_c_183_n N_VGND_c_944_n 0.00137572f $X=0.69 $Y=0.43 $X2=0
+ $Y2=0
cc_200 N_A_110_57#_c_161_n N_VGND_c_945_n 0.00424645f $X=1.865 $Y=1.185 $X2=0
+ $Y2=0
cc_201 N_A_110_57#_c_162_n N_VGND_c_945_n 0.00228818f $X=2.22 $Y=1.265 $X2=0
+ $Y2=0
cc_202 N_A_110_57#_c_163_n N_VGND_c_945_n 0.0027833f $X=2.295 $Y=1.185 $X2=0
+ $Y2=0
cc_203 N_A_110_57#_c_165_n N_VGND_c_946_n 0.0027833f $X=2.725 $Y=1.185 $X2=0
+ $Y2=0
cc_204 N_A_110_57#_c_166_n N_VGND_c_946_n 0.00228818f $X=3.08 $Y=1.265 $X2=0
+ $Y2=0
cc_205 N_A_110_57#_c_167_n N_VGND_c_946_n 0.0027833f $X=3.155 $Y=1.185 $X2=0
+ $Y2=0
cc_206 N_A_110_57#_c_169_n N_VGND_c_947_n 0.0027833f $X=3.585 $Y=1.185 $X2=0
+ $Y2=0
cc_207 N_A_110_57#_c_170_n N_VGND_c_947_n 0.00228818f $X=3.94 $Y=1.265 $X2=0
+ $Y2=0
cc_208 N_A_110_57#_c_171_n N_VGND_c_947_n 0.0027833f $X=4.015 $Y=1.185 $X2=0
+ $Y2=0
cc_209 N_A_110_57#_c_171_n N_VGND_c_948_n 0.00585385f $X=4.015 $Y=1.185 $X2=0
+ $Y2=0
cc_210 N_A_110_57#_c_173_n N_VGND_c_948_n 0.00585385f $X=4.445 $Y=1.185 $X2=0
+ $Y2=0
cc_211 N_A_110_57#_c_173_n N_VGND_c_949_n 0.0027833f $X=4.445 $Y=1.185 $X2=0
+ $Y2=0
cc_212 N_A_110_57#_c_174_n N_VGND_c_949_n 0.00228818f $X=4.8 $Y=1.265 $X2=0
+ $Y2=0
cc_213 N_A_110_57#_c_175_n N_VGND_c_949_n 0.00424645f $X=4.875 $Y=1.185 $X2=0
+ $Y2=0
cc_214 N_A_110_57#_c_161_n N_VGND_c_950_n 0.00585385f $X=1.865 $Y=1.185 $X2=0
+ $Y2=0
cc_215 N_A_110_57#_c_183_n N_VGND_c_950_n 0.0134832f $X=0.69 $Y=0.43 $X2=0 $Y2=0
cc_216 N_A_110_57#_c_185_n N_VGND_c_950_n 0.0087537f $X=1.15 $Y=0.83 $X2=0 $Y2=0
cc_217 N_A_110_57#_c_186_n N_VGND_c_950_n 0.00574822f $X=1.15 $Y=0.83 $X2=0
+ $Y2=0
cc_218 N_A_110_57#_c_163_n N_VGND_c_952_n 0.00585385f $X=2.295 $Y=1.185 $X2=0
+ $Y2=0
cc_219 N_A_110_57#_c_165_n N_VGND_c_952_n 0.00585385f $X=2.725 $Y=1.185 $X2=0
+ $Y2=0
cc_220 N_A_110_57#_c_167_n N_VGND_c_954_n 0.00585385f $X=3.155 $Y=1.185 $X2=0
+ $Y2=0
cc_221 N_A_110_57#_c_169_n N_VGND_c_954_n 0.00585385f $X=3.585 $Y=1.185 $X2=0
+ $Y2=0
cc_222 N_A_110_57#_c_175_n N_VGND_c_956_n 0.00585385f $X=4.875 $Y=1.185 $X2=0
+ $Y2=0
cc_223 N_A_110_57#_c_161_n N_VGND_c_957_n 0.0118221f $X=1.865 $Y=1.185 $X2=0
+ $Y2=0
cc_224 N_A_110_57#_c_163_n N_VGND_c_957_n 0.0105224f $X=2.295 $Y=1.185 $X2=0
+ $Y2=0
cc_225 N_A_110_57#_c_165_n N_VGND_c_957_n 0.0105224f $X=2.725 $Y=1.185 $X2=0
+ $Y2=0
cc_226 N_A_110_57#_c_167_n N_VGND_c_957_n 0.0105224f $X=3.155 $Y=1.185 $X2=0
+ $Y2=0
cc_227 N_A_110_57#_c_169_n N_VGND_c_957_n 0.0105224f $X=3.585 $Y=1.185 $X2=0
+ $Y2=0
cc_228 N_A_110_57#_c_171_n N_VGND_c_957_n 0.0105224f $X=4.015 $Y=1.185 $X2=0
+ $Y2=0
cc_229 N_A_110_57#_c_173_n N_VGND_c_957_n 0.0105224f $X=4.445 $Y=1.185 $X2=0
+ $Y2=0
cc_230 N_A_110_57#_c_175_n N_VGND_c_957_n 0.0105477f $X=4.875 $Y=1.185 $X2=0
+ $Y2=0
cc_231 N_A_110_57#_c_183_n N_VGND_c_957_n 0.00793704f $X=0.69 $Y=0.43 $X2=0
+ $Y2=0
cc_232 N_A_110_57#_c_185_n N_VGND_c_957_n 0.014669f $X=1.15 $Y=0.83 $X2=0 $Y2=0
cc_233 N_A_110_57#_c_186_n N_VGND_c_957_n 0.00926103f $X=1.15 $Y=0.83 $X2=0
+ $Y2=0
cc_234 N_A_110_57#_c_159_n N_A_305_47#_c_1060_n 0.0119277f $X=1.79 $Y=1.265
+ $X2=0 $Y2=0
cc_235 N_A_110_57#_c_161_n N_A_305_47#_c_1060_n 0.00313635f $X=1.865 $Y=1.185
+ $X2=0 $Y2=0
cc_236 N_A_110_57#_c_184_n N_A_305_47#_c_1060_n 0.0187399f $X=1.13 $Y=1.98 $X2=0
+ $Y2=0
cc_237 N_A_110_57#_c_185_n N_A_305_47#_c_1060_n 0.0310382f $X=1.15 $Y=0.83 $X2=0
+ $Y2=0
cc_238 N_A_110_57#_c_186_n N_A_305_47#_c_1060_n 0.00278505f $X=1.15 $Y=0.83
+ $X2=0 $Y2=0
cc_239 N_A_110_57#_c_159_n N_A_305_47#_c_1061_n 4.55988e-19 $X=1.79 $Y=1.265
+ $X2=0 $Y2=0
cc_240 N_A_110_57#_c_162_n N_A_305_47#_c_1061_n 0.00704942f $X=2.22 $Y=1.265
+ $X2=0 $Y2=0
cc_241 N_A_110_57#_c_164_n N_A_305_47#_c_1061_n 4.55988e-19 $X=2.65 $Y=1.265
+ $X2=0 $Y2=0
cc_242 N_A_110_57#_c_176_n N_A_305_47#_c_1061_n 0.00854977f $X=1.865 $Y=1.265
+ $X2=0 $Y2=0
cc_243 N_A_110_57#_c_177_n N_A_305_47#_c_1061_n 0.00854977f $X=2.295 $Y=1.265
+ $X2=0 $Y2=0
cc_244 N_A_110_57#_c_159_n N_A_305_47#_c_1062_n 0.00427593f $X=1.79 $Y=1.265
+ $X2=0 $Y2=0
cc_245 N_A_110_57#_c_184_n N_A_305_47#_c_1062_n 0.0189433f $X=1.13 $Y=1.98 $X2=0
+ $Y2=0
cc_246 N_A_110_57#_c_163_n N_A_305_47#_c_1063_n 0.00187564f $X=2.295 $Y=1.185
+ $X2=0 $Y2=0
cc_247 N_A_110_57#_c_164_n N_A_305_47#_c_1063_n 0.0101061f $X=2.65 $Y=1.265
+ $X2=0 $Y2=0
cc_248 N_A_110_57#_c_165_n N_A_305_47#_c_1063_n 0.00187564f $X=2.725 $Y=1.185
+ $X2=0 $Y2=0
cc_249 N_A_110_57#_c_164_n N_A_305_47#_c_1064_n 4.55988e-19 $X=2.65 $Y=1.265
+ $X2=0 $Y2=0
cc_250 N_A_110_57#_c_166_n N_A_305_47#_c_1064_n 0.00704942f $X=3.08 $Y=1.265
+ $X2=0 $Y2=0
cc_251 N_A_110_57#_c_168_n N_A_305_47#_c_1064_n 4.55988e-19 $X=3.51 $Y=1.265
+ $X2=0 $Y2=0
cc_252 N_A_110_57#_c_178_n N_A_305_47#_c_1064_n 0.00854977f $X=2.725 $Y=1.265
+ $X2=0 $Y2=0
cc_253 N_A_110_57#_c_179_n N_A_305_47#_c_1064_n 0.00854977f $X=3.155 $Y=1.265
+ $X2=0 $Y2=0
cc_254 N_A_110_57#_c_167_n N_A_305_47#_c_1065_n 0.00187564f $X=3.155 $Y=1.185
+ $X2=0 $Y2=0
cc_255 N_A_110_57#_c_168_n N_A_305_47#_c_1065_n 0.0101061f $X=3.51 $Y=1.265
+ $X2=0 $Y2=0
cc_256 N_A_110_57#_c_169_n N_A_305_47#_c_1065_n 0.00187564f $X=3.585 $Y=1.185
+ $X2=0 $Y2=0
cc_257 N_A_110_57#_c_168_n N_A_305_47#_c_1066_n 4.55988e-19 $X=3.51 $Y=1.265
+ $X2=0 $Y2=0
cc_258 N_A_110_57#_c_170_n N_A_305_47#_c_1066_n 0.00704942f $X=3.94 $Y=1.265
+ $X2=0 $Y2=0
cc_259 N_A_110_57#_c_172_n N_A_305_47#_c_1066_n 4.55988e-19 $X=4.37 $Y=1.265
+ $X2=0 $Y2=0
cc_260 N_A_110_57#_c_180_n N_A_305_47#_c_1066_n 0.00854977f $X=3.585 $Y=1.265
+ $X2=0 $Y2=0
cc_261 N_A_110_57#_c_181_n N_A_305_47#_c_1066_n 0.00854977f $X=4.015 $Y=1.265
+ $X2=0 $Y2=0
cc_262 N_A_110_57#_c_171_n N_A_305_47#_c_1067_n 0.00187564f $X=4.015 $Y=1.185
+ $X2=0 $Y2=0
cc_263 N_A_110_57#_c_172_n N_A_305_47#_c_1067_n 0.00997154f $X=4.37 $Y=1.265
+ $X2=0 $Y2=0
cc_264 N_A_110_57#_c_173_n N_A_305_47#_c_1067_n 0.00187564f $X=4.445 $Y=1.185
+ $X2=0 $Y2=0
cc_265 N_A_110_57#_c_172_n N_A_305_47#_c_1068_n 4.55988e-19 $X=4.37 $Y=1.265
+ $X2=0 $Y2=0
cc_266 N_A_110_57#_c_174_n N_A_305_47#_c_1068_n 0.016146f $X=4.8 $Y=1.265 $X2=0
+ $Y2=0
cc_267 N_A_110_57#_c_182_n N_A_305_47#_c_1068_n 0.00854977f $X=4.445 $Y=1.265
+ $X2=0 $Y2=0
cc_268 N_A_110_57#_c_175_n N_A_305_47#_c_1069_n 0.00353987f $X=4.875 $Y=1.185
+ $X2=0 $Y2=0
cc_269 N_A_110_57#_c_164_n N_A_305_47#_c_1072_n 0.00300205f $X=2.65 $Y=1.265
+ $X2=0 $Y2=0
cc_270 N_A_110_57#_c_168_n N_A_305_47#_c_1073_n 0.00300205f $X=3.51 $Y=1.265
+ $X2=0 $Y2=0
cc_271 N_A_110_57#_c_172_n N_A_305_47#_c_1074_n 0.00300205f $X=4.37 $Y=1.265
+ $X2=0 $Y2=0
cc_272 N_TE_B_c_310_n N_A_M1003_g 0.0250876f $X=4.8 $Y=1.64 $X2=0 $Y2=0
cc_273 N_TE_B_c_319_n N_VPWR_c_602_n 0.00878211f $X=0.915 $Y=1.725 $X2=0 $Y2=0
cc_274 N_TE_B_c_303_n N_VPWR_c_602_n 0.00615812f $X=0.99 $Y=1.64 $X2=0 $Y2=0
cc_275 N_TE_B_c_318_n N_VPWR_c_602_n 0.0153853f $X=0.61 $Y=1.46 $X2=0 $Y2=0
cc_276 TE_B N_VPWR_c_602_n 0.08652f $X=0.24 $Y=1.665 $X2=0 $Y2=0
cc_277 N_TE_B_c_322_n N_VPWR_c_603_n 0.0164399f $X=1.865 $Y=1.725 $X2=0 $Y2=0
cc_278 N_TE_B_c_304_n N_VPWR_c_603_n 5.05051e-19 $X=2.22 $Y=1.64 $X2=0 $Y2=0
cc_279 N_TE_B_c_324_n N_VPWR_c_603_n 0.0144597f $X=2.295 $Y=1.725 $X2=0 $Y2=0
cc_280 N_TE_B_c_326_n N_VPWR_c_603_n 7.27171e-19 $X=2.725 $Y=1.725 $X2=0 $Y2=0
cc_281 N_TE_B_c_324_n N_VPWR_c_604_n 7.27171e-19 $X=2.295 $Y=1.725 $X2=0 $Y2=0
cc_282 N_TE_B_c_326_n N_VPWR_c_604_n 0.0144597f $X=2.725 $Y=1.725 $X2=0 $Y2=0
cc_283 N_TE_B_c_306_n N_VPWR_c_604_n 5.05051e-19 $X=3.08 $Y=1.64 $X2=0 $Y2=0
cc_284 N_TE_B_c_328_n N_VPWR_c_604_n 0.0144597f $X=3.155 $Y=1.725 $X2=0 $Y2=0
cc_285 N_TE_B_c_330_n N_VPWR_c_604_n 7.27171e-19 $X=3.585 $Y=1.725 $X2=0 $Y2=0
cc_286 N_TE_B_c_328_n N_VPWR_c_605_n 7.27171e-19 $X=3.155 $Y=1.725 $X2=0 $Y2=0
cc_287 N_TE_B_c_330_n N_VPWR_c_605_n 0.0144597f $X=3.585 $Y=1.725 $X2=0 $Y2=0
cc_288 N_TE_B_c_308_n N_VPWR_c_605_n 5.05051e-19 $X=3.94 $Y=1.64 $X2=0 $Y2=0
cc_289 N_TE_B_c_332_n N_VPWR_c_605_n 0.0144597f $X=4.015 $Y=1.725 $X2=0 $Y2=0
cc_290 N_TE_B_c_334_n N_VPWR_c_605_n 7.27171e-19 $X=4.445 $Y=1.725 $X2=0 $Y2=0
cc_291 N_TE_B_c_332_n N_VPWR_c_606_n 0.00486043f $X=4.015 $Y=1.725 $X2=0 $Y2=0
cc_292 N_TE_B_c_334_n N_VPWR_c_606_n 0.00486043f $X=4.445 $Y=1.725 $X2=0 $Y2=0
cc_293 N_TE_B_c_332_n N_VPWR_c_607_n 7.27171e-19 $X=4.015 $Y=1.725 $X2=0 $Y2=0
cc_294 N_TE_B_c_334_n N_VPWR_c_607_n 0.0144597f $X=4.445 $Y=1.725 $X2=0 $Y2=0
cc_295 N_TE_B_c_310_n N_VPWR_c_607_n 5.05051e-19 $X=4.8 $Y=1.64 $X2=0 $Y2=0
cc_296 N_TE_B_c_336_n N_VPWR_c_607_n 0.0156326f $X=4.875 $Y=1.725 $X2=0 $Y2=0
cc_297 N_TE_B_c_324_n N_VPWR_c_608_n 0.00486043f $X=2.295 $Y=1.725 $X2=0 $Y2=0
cc_298 N_TE_B_c_326_n N_VPWR_c_608_n 0.00486043f $X=2.725 $Y=1.725 $X2=0 $Y2=0
cc_299 N_TE_B_c_328_n N_VPWR_c_610_n 0.00486043f $X=3.155 $Y=1.725 $X2=0 $Y2=0
cc_300 N_TE_B_c_330_n N_VPWR_c_610_n 0.00486043f $X=3.585 $Y=1.725 $X2=0 $Y2=0
cc_301 TE_B N_VPWR_c_612_n 0.0127207f $X=0.24 $Y=1.665 $X2=0 $Y2=0
cc_302 N_TE_B_c_319_n N_VPWR_c_613_n 0.00579312f $X=0.915 $Y=1.725 $X2=0 $Y2=0
cc_303 N_TE_B_c_322_n N_VPWR_c_613_n 0.00486043f $X=1.865 $Y=1.725 $X2=0 $Y2=0
cc_304 N_TE_B_c_336_n N_VPWR_c_614_n 0.00486043f $X=4.875 $Y=1.725 $X2=0 $Y2=0
cc_305 N_TE_B_c_319_n N_VPWR_c_601_n 0.0130517f $X=0.915 $Y=1.725 $X2=0 $Y2=0
cc_306 N_TE_B_c_322_n N_VPWR_c_601_n 0.00954696f $X=1.865 $Y=1.725 $X2=0 $Y2=0
cc_307 N_TE_B_c_324_n N_VPWR_c_601_n 0.00824727f $X=2.295 $Y=1.725 $X2=0 $Y2=0
cc_308 N_TE_B_c_326_n N_VPWR_c_601_n 0.00824727f $X=2.725 $Y=1.725 $X2=0 $Y2=0
cc_309 N_TE_B_c_328_n N_VPWR_c_601_n 0.00824727f $X=3.155 $Y=1.725 $X2=0 $Y2=0
cc_310 N_TE_B_c_330_n N_VPWR_c_601_n 0.00824727f $X=3.585 $Y=1.725 $X2=0 $Y2=0
cc_311 N_TE_B_c_332_n N_VPWR_c_601_n 0.00824727f $X=4.015 $Y=1.725 $X2=0 $Y2=0
cc_312 N_TE_B_c_334_n N_VPWR_c_601_n 0.00824727f $X=4.445 $Y=1.725 $X2=0 $Y2=0
cc_313 N_TE_B_c_336_n N_VPWR_c_601_n 0.0082726f $X=4.875 $Y=1.725 $X2=0 $Y2=0
cc_314 TE_B N_VPWR_c_601_n 0.0112374f $X=0.24 $Y=1.665 $X2=0 $Y2=0
cc_315 N_TE_B_c_319_n N_A_305_367#_c_729_n 0.00187619f $X=0.915 $Y=1.725 $X2=0
+ $Y2=0
cc_316 N_TE_B_c_302_n N_A_305_367#_c_735_n 5.27972e-19 $X=1.79 $Y=1.64 $X2=0
+ $Y2=0
cc_317 N_TE_B_c_322_n N_A_305_367#_c_735_n 0.0134493f $X=1.865 $Y=1.725 $X2=0
+ $Y2=0
cc_318 N_TE_B_c_304_n N_A_305_367#_c_735_n 0.00525471f $X=2.22 $Y=1.64 $X2=0
+ $Y2=0
cc_319 N_TE_B_c_324_n N_A_305_367#_c_735_n 0.0125573f $X=2.295 $Y=1.725 $X2=0
+ $Y2=0
cc_320 N_TE_B_c_305_n N_A_305_367#_c_735_n 5.27972e-19 $X=2.65 $Y=1.64 $X2=0
+ $Y2=0
cc_321 N_TE_B_c_311_n N_A_305_367#_c_735_n 0.00184441f $X=1.865 $Y=1.64 $X2=0
+ $Y2=0
cc_322 N_TE_B_c_312_n N_A_305_367#_c_735_n 0.00184441f $X=2.295 $Y=1.64 $X2=0
+ $Y2=0
cc_323 N_TE_B_c_319_n N_A_305_367#_c_730_n 5.9011e-19 $X=0.915 $Y=1.725 $X2=0
+ $Y2=0
cc_324 N_TE_B_c_302_n N_A_305_367#_c_730_n 0.00912496f $X=1.79 $Y=1.64 $X2=0
+ $Y2=0
cc_325 N_TE_B_c_305_n N_A_305_367#_c_737_n 5.27972e-19 $X=2.65 $Y=1.64 $X2=0
+ $Y2=0
cc_326 N_TE_B_c_326_n N_A_305_367#_c_737_n 0.0125573f $X=2.725 $Y=1.725 $X2=0
+ $Y2=0
cc_327 N_TE_B_c_306_n N_A_305_367#_c_737_n 0.00525471f $X=3.08 $Y=1.64 $X2=0
+ $Y2=0
cc_328 N_TE_B_c_328_n N_A_305_367#_c_737_n 0.0125573f $X=3.155 $Y=1.725 $X2=0
+ $Y2=0
cc_329 N_TE_B_c_307_n N_A_305_367#_c_737_n 5.27972e-19 $X=3.51 $Y=1.64 $X2=0
+ $Y2=0
cc_330 N_TE_B_c_313_n N_A_305_367#_c_737_n 0.00184441f $X=2.725 $Y=1.64 $X2=0
+ $Y2=0
cc_331 N_TE_B_c_314_n N_A_305_367#_c_737_n 0.00184441f $X=3.155 $Y=1.64 $X2=0
+ $Y2=0
cc_332 N_TE_B_c_307_n N_A_305_367#_c_738_n 5.27972e-19 $X=3.51 $Y=1.64 $X2=0
+ $Y2=0
cc_333 N_TE_B_c_330_n N_A_305_367#_c_738_n 0.0125573f $X=3.585 $Y=1.725 $X2=0
+ $Y2=0
cc_334 N_TE_B_c_308_n N_A_305_367#_c_738_n 0.00525471f $X=3.94 $Y=1.64 $X2=0
+ $Y2=0
cc_335 N_TE_B_c_332_n N_A_305_367#_c_738_n 0.0125573f $X=4.015 $Y=1.725 $X2=0
+ $Y2=0
cc_336 N_TE_B_c_309_n N_A_305_367#_c_738_n 5.27972e-19 $X=4.37 $Y=1.64 $X2=0
+ $Y2=0
cc_337 N_TE_B_c_315_n N_A_305_367#_c_738_n 0.00184441f $X=3.585 $Y=1.64 $X2=0
+ $Y2=0
cc_338 N_TE_B_c_316_n N_A_305_367#_c_738_n 0.00184441f $X=4.015 $Y=1.64 $X2=0
+ $Y2=0
cc_339 N_TE_B_c_309_n N_A_305_367#_c_731_n 5.27972e-19 $X=4.37 $Y=1.64 $X2=0
+ $Y2=0
cc_340 N_TE_B_c_334_n N_A_305_367#_c_731_n 0.0125024f $X=4.445 $Y=1.725 $X2=0
+ $Y2=0
cc_341 N_TE_B_c_310_n N_A_305_367#_c_731_n 0.00755325f $X=4.8 $Y=1.64 $X2=0
+ $Y2=0
cc_342 N_TE_B_c_336_n N_A_305_367#_c_731_n 0.0122683f $X=4.875 $Y=1.725 $X2=0
+ $Y2=0
cc_343 N_TE_B_c_317_n N_A_305_367#_c_731_n 0.00184441f $X=4.445 $Y=1.64 $X2=0
+ $Y2=0
cc_344 N_TE_B_c_305_n N_A_305_367#_c_769_n 0.00475798f $X=2.65 $Y=1.64 $X2=0
+ $Y2=0
cc_345 N_TE_B_c_307_n N_A_305_367#_c_770_n 0.00475798f $X=3.51 $Y=1.64 $X2=0
+ $Y2=0
cc_346 N_TE_B_c_309_n N_A_305_367#_c_771_n 0.00475798f $X=4.37 $Y=1.64 $X2=0
+ $Y2=0
cc_347 N_TE_B_M1023_g N_VGND_c_944_n 0.0058048f $X=0.475 $Y=0.705 $X2=0 $Y2=0
cc_348 N_TE_B_c_303_n N_VGND_c_944_n 0.00168578f $X=0.99 $Y=1.64 $X2=0 $Y2=0
cc_349 N_TE_B_c_318_n N_VGND_c_944_n 0.0231146f $X=0.61 $Y=1.46 $X2=0 $Y2=0
cc_350 N_TE_B_M1023_g N_VGND_c_950_n 0.0053602f $X=0.475 $Y=0.705 $X2=0 $Y2=0
cc_351 N_TE_B_M1023_g N_VGND_c_957_n 0.01173f $X=0.475 $Y=0.705 $X2=0 $Y2=0
cc_352 N_TE_B_c_302_n N_A_305_47#_c_1061_n 0.00445188f $X=1.79 $Y=1.64 $X2=0
+ $Y2=0
cc_353 N_TE_B_c_302_n N_A_305_47#_c_1062_n 0.00225083f $X=1.79 $Y=1.64 $X2=0
+ $Y2=0
cc_354 N_TE_B_c_305_n N_A_305_47#_c_1064_n 0.00445188f $X=2.65 $Y=1.64 $X2=0
+ $Y2=0
cc_355 N_TE_B_c_307_n N_A_305_47#_c_1066_n 0.00445188f $X=3.51 $Y=1.64 $X2=0
+ $Y2=0
cc_356 N_TE_B_c_309_n N_A_305_47#_c_1068_n 0.00438275f $X=4.37 $Y=1.64 $X2=0
+ $Y2=0
cc_357 N_TE_B_c_305_n N_A_305_47#_c_1072_n 0.00210288f $X=2.65 $Y=1.64 $X2=0
+ $Y2=0
cc_358 N_TE_B_c_307_n N_A_305_47#_c_1073_n 0.00210288f $X=3.51 $Y=1.64 $X2=0
+ $Y2=0
cc_359 N_TE_B_c_309_n N_A_305_47#_c_1074_n 0.00210288f $X=4.37 $Y=1.64 $X2=0
+ $Y2=0
cc_360 N_A_M1003_g N_VPWR_c_607_n 0.00109252f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_361 N_A_M1003_g N_VPWR_c_614_n 0.00357877f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_362 N_A_M1007_g N_VPWR_c_614_n 0.00357877f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A_M1008_g N_VPWR_c_614_n 0.00357877f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_364 N_A_M1009_g N_VPWR_c_614_n 0.00357877f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_365 N_A_M1020_g N_VPWR_c_614_n 0.00357877f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_366 N_A_M1021_g N_VPWR_c_614_n 0.00357877f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_367 N_A_M1029_g N_VPWR_c_614_n 0.00357877f $X=7.885 $Y=2.465 $X2=0 $Y2=0
cc_368 N_A_M1031_g N_VPWR_c_614_n 0.00357877f $X=8.315 $Y=2.465 $X2=0 $Y2=0
cc_369 N_A_M1003_g N_VPWR_c_601_n 0.00537654f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_370 N_A_M1007_g N_VPWR_c_601_n 0.0053512f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_371 N_A_M1008_g N_VPWR_c_601_n 0.0053512f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_372 N_A_M1009_g N_VPWR_c_601_n 0.0053512f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_373 N_A_M1020_g N_VPWR_c_601_n 0.0053512f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A_M1021_g N_VPWR_c_601_n 0.0053512f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_375 N_A_M1029_g N_VPWR_c_601_n 0.0053512f $X=7.885 $Y=2.465 $X2=0 $Y2=0
cc_376 N_A_M1031_g N_VPWR_c_601_n 0.00665089f $X=8.315 $Y=2.465 $X2=0 $Y2=0
cc_377 N_A_M1003_g N_A_305_367#_c_731_n 0.00155056f $X=5.305 $Y=2.465 $X2=0
+ $Y2=0
cc_378 N_A_M1003_g N_A_305_367#_c_773_n 0.0115031f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_379 N_A_M1007_g N_A_305_367#_c_773_n 0.0114565f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A_M1008_g N_A_305_367#_c_775_n 0.0115031f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_381 N_A_M1009_g N_A_305_367#_c_775_n 0.0115031f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_382 N_A_c_477_n N_A_305_367#_c_777_n 3.75556e-19 $X=8.315 $Y=1.35 $X2=0 $Y2=0
cc_383 N_A_M1020_g N_A_305_367#_c_778_n 0.0115031f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_384 N_A_M1021_g N_A_305_367#_c_778_n 0.0115031f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_385 N_A_c_477_n N_A_305_367#_c_780_n 3.75556e-19 $X=8.315 $Y=1.35 $X2=0 $Y2=0
cc_386 N_A_M1029_g N_A_305_367#_c_781_n 0.0115031f $X=7.885 $Y=2.465 $X2=0 $Y2=0
cc_387 N_A_M1031_g N_A_305_367#_c_781_n 0.0115031f $X=8.315 $Y=2.465 $X2=0 $Y2=0
cc_388 N_A_M1031_g N_A_305_367#_c_733_n 0.0029331f $X=8.315 $Y=2.465 $X2=0 $Y2=0
cc_389 N_A_M1003_g N_Z_c_864_n 0.01237f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_390 N_A_M1007_g N_Z_c_864_n 0.0136935f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_391 N_A_M1008_g N_Z_c_864_n 6.56666e-19 $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_392 N_A_c_461_n N_Z_c_861_n 0.00395163f $X=5.305 $Y=1.185 $X2=0 $Y2=0
cc_393 N_A_c_463_n N_Z_c_861_n 0.0124788f $X=5.735 $Y=1.185 $X2=0 $Y2=0
cc_394 N_A_M1007_g N_Z_c_861_n 0.0117018f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_395 N_A_c_465_n N_Z_c_861_n 0.0140602f $X=6.165 $Y=1.185 $X2=0 $Y2=0
cc_396 N_A_M1008_g N_Z_c_861_n 0.0128612f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_397 A N_Z_c_861_n 0.0841442f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_398 N_A_c_477_n N_Z_c_861_n 0.00680243f $X=8.315 $Y=1.35 $X2=0 $Y2=0
cc_399 N_A_M1003_g N_Z_c_862_n 0.0040804f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_400 N_A_M1007_g N_Z_c_862_n 0.00258557f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_401 A N_Z_c_862_n 0.0276081f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_402 N_A_c_477_n N_Z_c_862_n 0.00232957f $X=8.315 $Y=1.35 $X2=0 $Y2=0
cc_403 N_A_M1007_g N_Z_c_878_n 6.56666e-19 $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_404 N_A_M1008_g N_Z_c_878_n 0.0136935f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_405 N_A_M1009_g N_Z_c_878_n 0.0136935f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_406 N_A_M1020_g N_Z_c_878_n 6.56666e-19 $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_407 N_A_M1009_g N_Z_c_882_n 6.56666e-19 $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_408 N_A_M1020_g N_Z_c_882_n 0.0136935f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_409 N_A_M1021_g N_Z_c_882_n 0.0136935f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_410 N_A_M1029_g N_Z_c_882_n 6.56666e-19 $X=7.885 $Y=2.465 $X2=0 $Y2=0
cc_411 N_A_c_469_n N_Z_c_858_n 0.00137536f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_412 N_A_c_471_n N_Z_c_858_n 0.00137599f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_413 N_A_M1021_g N_Z_c_888_n 6.56666e-19 $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_414 N_A_M1029_g N_Z_c_888_n 0.0136935f $X=7.885 $Y=2.465 $X2=0 $Y2=0
cc_415 N_A_M1031_g N_Z_c_888_n 0.0128496f $X=8.315 $Y=2.465 $X2=0 $Y2=0
cc_416 N_A_c_473_n N_Z_c_859_n 0.00139595f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_417 N_A_c_475_n N_Z_c_859_n 0.00186692f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_418 N_A_c_465_n N_Z_c_860_n 0.00421371f $X=6.165 $Y=1.185 $X2=0 $Y2=0
cc_419 N_A_M1008_g N_Z_c_860_n 0.00824293f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_420 N_A_c_467_n N_Z_c_860_n 0.00639949f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_421 N_A_M1009_g N_Z_c_860_n 0.0165798f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_422 N_A_c_469_n N_Z_c_860_n 0.00834088f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_423 N_A_M1020_g N_Z_c_860_n 0.0170518f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_424 N_A_c_471_n N_Z_c_860_n 0.00834088f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_425 N_A_M1021_g N_Z_c_860_n 0.0170573f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_426 N_A_c_473_n N_Z_c_860_n 0.00825947f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_427 N_A_M1029_g N_Z_c_860_n 0.0167817f $X=7.885 $Y=2.465 $X2=0 $Y2=0
cc_428 N_A_c_475_n N_Z_c_860_n 0.00149168f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_429 N_A_M1031_g N_Z_c_860_n 0.0163822f $X=8.315 $Y=2.465 $X2=0 $Y2=0
cc_430 A N_Z_c_860_n 0.0277655f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_431 N_A_c_477_n N_Z_c_860_n 0.100819f $X=8.315 $Y=1.35 $X2=0 $Y2=0
cc_432 N_A_c_461_n N_VGND_c_956_n 0.00357877f $X=5.305 $Y=1.185 $X2=0 $Y2=0
cc_433 N_A_c_463_n N_VGND_c_956_n 0.00357877f $X=5.735 $Y=1.185 $X2=0 $Y2=0
cc_434 N_A_c_465_n N_VGND_c_956_n 0.00357877f $X=6.165 $Y=1.185 $X2=0 $Y2=0
cc_435 N_A_c_467_n N_VGND_c_956_n 0.00357842f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_436 N_A_c_469_n N_VGND_c_956_n 0.00357842f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_437 N_A_c_471_n N_VGND_c_956_n 0.00357842f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_438 N_A_c_473_n N_VGND_c_956_n 0.00357842f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_439 N_A_c_475_n N_VGND_c_956_n 0.00357877f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_440 N_A_c_461_n N_VGND_c_957_n 0.00537654f $X=5.305 $Y=1.185 $X2=0 $Y2=0
cc_441 N_A_c_463_n N_VGND_c_957_n 0.0053512f $X=5.735 $Y=1.185 $X2=0 $Y2=0
cc_442 N_A_c_465_n N_VGND_c_957_n 0.0053512f $X=6.165 $Y=1.185 $X2=0 $Y2=0
cc_443 N_A_c_467_n N_VGND_c_957_n 0.00535118f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_444 N_A_c_469_n N_VGND_c_957_n 0.00535118f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_445 N_A_c_471_n N_VGND_c_957_n 0.00535118f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_446 N_A_c_473_n N_VGND_c_957_n 0.00535118f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_447 N_A_c_475_n N_VGND_c_957_n 0.00665089f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_448 A N_A_305_47#_c_1068_n 0.0196111f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_449 N_A_c_477_n N_A_305_47#_c_1068_n 0.00566904f $X=8.315 $Y=1.35 $X2=0 $Y2=0
cc_450 N_A_c_461_n N_A_305_47#_c_1069_n 0.00431169f $X=5.305 $Y=1.185 $X2=0
+ $Y2=0
cc_451 A N_A_305_47#_c_1069_n 0.0080339f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_452 N_A_c_461_n N_A_305_47#_c_1125_n 0.0142368f $X=5.305 $Y=1.185 $X2=0 $Y2=0
cc_453 N_A_c_463_n N_A_305_47#_c_1125_n 0.0101209f $X=5.735 $Y=1.185 $X2=0 $Y2=0
cc_454 N_A_c_465_n N_A_305_47#_c_1125_n 0.0101938f $X=6.165 $Y=1.185 $X2=0 $Y2=0
cc_455 N_A_c_467_n N_A_305_47#_c_1125_n 0.0108825f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_456 N_A_c_477_n N_A_305_47#_c_1125_n 2.74016e-19 $X=8.315 $Y=1.35 $X2=0 $Y2=0
cc_457 N_A_c_469_n N_A_305_47#_c_1130_n 0.0105205f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_458 N_A_c_471_n N_A_305_47#_c_1130_n 0.0105205f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_459 N_A_c_473_n N_A_305_47#_c_1070_n 0.0105205f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_460 N_A_c_475_n N_A_305_47#_c_1070_n 0.012237f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_461 N_A_c_475_n N_A_305_47#_c_1071_n 0.00269856f $X=8.315 $Y=1.185 $X2=0
+ $Y2=0
cc_462 N_A_c_465_n N_A_305_47#_c_1135_n 7.61713e-19 $X=6.165 $Y=1.185 $X2=0
+ $Y2=0
cc_463 N_A_c_467_n N_A_305_47#_c_1135_n 0.00835573f $X=6.595 $Y=1.185 $X2=0
+ $Y2=0
cc_464 N_A_c_469_n N_A_305_47#_c_1135_n 0.0089814f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_465 N_A_c_471_n N_A_305_47#_c_1135_n 5.39928e-19 $X=7.455 $Y=1.185 $X2=0
+ $Y2=0
cc_466 N_A_c_477_n N_A_305_47#_c_1135_n 7.00643e-19 $X=8.315 $Y=1.35 $X2=0 $Y2=0
cc_467 N_A_c_469_n N_A_305_47#_c_1140_n 5.40824e-19 $X=7.025 $Y=1.185 $X2=0
+ $Y2=0
cc_468 N_A_c_471_n N_A_305_47#_c_1140_n 0.0088546f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_469 N_A_c_473_n N_A_305_47#_c_1140_n 0.00893811f $X=7.885 $Y=1.185 $X2=0
+ $Y2=0
cc_470 N_A_c_475_n N_A_305_47#_c_1140_n 5.47147e-19 $X=8.315 $Y=1.185 $X2=0
+ $Y2=0
cc_471 N_A_c_477_n N_A_305_47#_c_1140_n 7.00643e-19 $X=8.315 $Y=1.35 $X2=0 $Y2=0
cc_472 N_VPWR_c_601_n N_A_305_367#_M1001_s 0.00371702f $X=8.88 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_473 N_VPWR_c_601_n N_A_305_367#_M1006_s 0.00536646f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_601_n N_A_305_367#_M1018_s 0.00536646f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_601_n N_A_305_367#_M1024_s 0.00536646f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_601_n N_A_305_367#_M1030_s 0.00376627f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_601_n N_A_305_367#_M1007_d 0.00223565f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_601_n N_A_305_367#_M1009_d 0.00223565f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_601_n N_A_305_367#_M1021_d 0.00223565f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_601_n N_A_305_367#_M1031_d 0.00215161f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_613_n N_A_305_367#_c_729_n 0.0178111f $X=1.915 $Y=3.33 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_601_n N_A_305_367#_c_729_n 0.0100304f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_483 N_VPWR_M1001_d N_A_305_367#_c_735_n 0.00178571f $X=1.94 $Y=1.835 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_603_n N_A_305_367#_c_735_n 0.0175375f $X=2.08 $Y=2.18 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_608_n N_A_305_367#_c_797_n 0.0124525f $X=2.775 $Y=3.33 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_601_n N_A_305_367#_c_797_n 0.00730901f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_487 N_VPWR_M1011_d N_A_305_367#_c_737_n 0.00178571f $X=2.8 $Y=1.835 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_604_n N_A_305_367#_c_737_n 0.0175375f $X=2.94 $Y=2.18 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_610_n N_A_305_367#_c_801_n 0.0124525f $X=3.635 $Y=3.33 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_601_n N_A_305_367#_c_801_n 0.00730901f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_491 N_VPWR_M1022_d N_A_305_367#_c_738_n 0.00178571f $X=3.66 $Y=1.835 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_605_n N_A_305_367#_c_738_n 0.0175375f $X=3.8 $Y=2.18 $X2=0 $Y2=0
cc_493 N_VPWR_c_606_n N_A_305_367#_c_805_n 0.0124525f $X=4.495 $Y=3.33 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_601_n N_A_305_367#_c_805_n 0.00730901f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_495 N_VPWR_M1025_d N_A_305_367#_c_731_n 0.00178571f $X=4.52 $Y=1.835 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_607_n N_A_305_367#_c_731_n 0.0175375f $X=4.66 $Y=2.18 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_614_n N_A_305_367#_c_809_n 0.0125234f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_601_n N_A_305_367#_c_809_n 0.00738148f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_614_n N_A_305_367#_c_773_n 0.0361172f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_601_n N_A_305_367#_c_773_n 0.023676f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_501 N_VPWR_c_614_n N_A_305_367#_c_775_n 0.0361172f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_601_n N_A_305_367#_c_775_n 0.023676f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_503 N_VPWR_c_614_n N_A_305_367#_c_778_n 0.0361172f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_601_n N_A_305_367#_c_778_n 0.023676f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_505 N_VPWR_c_614_n N_A_305_367#_c_781_n 0.0361172f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_601_n N_A_305_367#_c_781_n 0.023676f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_507 N_VPWR_c_614_n N_A_305_367#_c_732_n 0.0179183f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_601_n N_A_305_367#_c_732_n 0.0101029f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_614_n N_A_305_367#_c_821_n 0.0125234f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_601_n N_A_305_367#_c_821_n 0.00738676f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_614_n N_A_305_367#_c_823_n 0.0125234f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_601_n N_A_305_367#_c_823_n 0.00738676f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_614_n N_A_305_367#_c_825_n 0.0125234f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_514 N_VPWR_c_601_n N_A_305_367#_c_825_n 0.00738676f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_601_n N_Z_M1003_s 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_516 N_VPWR_c_601_n N_Z_M1008_s 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_517 N_VPWR_c_601_n N_Z_M1020_s 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_518 N_VPWR_c_601_n N_Z_M1029_s 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_519 N_A_305_367#_c_773_n N_Z_M1003_s 0.00332344f $X=5.855 $Y=2.99 $X2=0 $Y2=0
cc_520 N_A_305_367#_c_775_n N_Z_M1008_s 0.00332344f $X=6.715 $Y=2.99 $X2=0 $Y2=0
cc_521 N_A_305_367#_c_778_n N_Z_M1020_s 0.00332344f $X=7.575 $Y=2.99 $X2=0 $Y2=0
cc_522 N_A_305_367#_c_781_n N_Z_M1029_s 0.00332344f $X=8.435 $Y=2.99 $X2=0 $Y2=0
cc_523 N_A_305_367#_c_773_n N_Z_c_864_n 0.0159805f $X=5.855 $Y=2.99 $X2=0 $Y2=0
cc_524 N_A_305_367#_M1007_d N_Z_c_861_n 0.00181369f $X=5.81 $Y=1.835 $X2=0 $Y2=0
cc_525 N_A_305_367#_c_833_p N_Z_c_861_n 0.0130379f $X=5.95 $Y=2.22 $X2=0 $Y2=0
cc_526 N_A_305_367#_c_731_n N_Z_c_862_n 0.0150174f $X=4.995 $Y=1.8 $X2=0 $Y2=0
cc_527 N_A_305_367#_c_775_n N_Z_c_878_n 0.0159805f $X=6.715 $Y=2.99 $X2=0 $Y2=0
cc_528 N_A_305_367#_c_778_n N_Z_c_882_n 0.0159805f $X=7.575 $Y=2.99 $X2=0 $Y2=0
cc_529 N_A_305_367#_c_781_n N_Z_c_888_n 0.0159805f $X=8.435 $Y=2.99 $X2=0 $Y2=0
cc_530 N_A_305_367#_M1009_d N_Z_c_860_n 0.00188202f $X=6.67 $Y=1.835 $X2=0 $Y2=0
cc_531 N_A_305_367#_M1021_d N_Z_c_860_n 0.00188202f $X=7.53 $Y=1.835 $X2=0 $Y2=0
cc_532 N_A_305_367#_c_777_n N_Z_c_860_n 0.0143367f $X=6.81 $Y=2.22 $X2=0 $Y2=0
cc_533 N_A_305_367#_c_780_n N_Z_c_860_n 0.0143367f $X=7.67 $Y=2.22 $X2=0 $Y2=0
cc_534 N_A_305_367#_c_733_n N_Z_c_860_n 0.00246889f $X=8.53 $Y=1.99 $X2=0 $Y2=0
cc_535 N_A_305_367#_c_735_n N_A_305_47#_c_1061_n 0.0448297f $X=2.415 $Y=1.8
+ $X2=0 $Y2=0
cc_536 N_A_305_367#_c_735_n N_A_305_47#_c_1062_n 0.00286013f $X=2.415 $Y=1.8
+ $X2=0 $Y2=0
cc_537 N_A_305_367#_c_730_n N_A_305_47#_c_1062_n 0.0231769f $X=1.745 $Y=1.8
+ $X2=0 $Y2=0
cc_538 N_A_305_367#_c_737_n N_A_305_47#_c_1064_n 0.0448297f $X=3.275 $Y=1.8
+ $X2=0 $Y2=0
cc_539 N_A_305_367#_c_738_n N_A_305_47#_c_1066_n 0.0448297f $X=4.135 $Y=1.8
+ $X2=0 $Y2=0
cc_540 N_A_305_367#_c_731_n N_A_305_47#_c_1068_n 0.0657039f $X=4.995 $Y=1.8
+ $X2=0 $Y2=0
cc_541 N_A_305_367#_c_735_n N_A_305_47#_c_1072_n 0.00286013f $X=2.415 $Y=1.8
+ $X2=0 $Y2=0
cc_542 N_A_305_367#_c_737_n N_A_305_47#_c_1072_n 0.00286013f $X=3.275 $Y=1.8
+ $X2=0 $Y2=0
cc_543 N_A_305_367#_c_769_n N_A_305_47#_c_1072_n 0.0169369f $X=2.51 $Y=1.8 $X2=0
+ $Y2=0
cc_544 N_A_305_367#_c_737_n N_A_305_47#_c_1073_n 0.00286013f $X=3.275 $Y=1.8
+ $X2=0 $Y2=0
cc_545 N_A_305_367#_c_738_n N_A_305_47#_c_1073_n 0.00286013f $X=4.135 $Y=1.8
+ $X2=0 $Y2=0
cc_546 N_A_305_367#_c_770_n N_A_305_47#_c_1073_n 0.0169369f $X=3.37 $Y=1.8 $X2=0
+ $Y2=0
cc_547 N_A_305_367#_c_738_n N_A_305_47#_c_1074_n 0.00286013f $X=4.135 $Y=1.8
+ $X2=0 $Y2=0
cc_548 N_A_305_367#_c_731_n N_A_305_47#_c_1074_n 0.00286013f $X=4.995 $Y=1.8
+ $X2=0 $Y2=0
cc_549 N_A_305_367#_c_771_n N_A_305_47#_c_1074_n 0.0169369f $X=4.23 $Y=1.8 $X2=0
+ $Y2=0
cc_550 N_Z_M1000_s N_VGND_c_957_n 0.00225186f $X=5.38 $Y=0.235 $X2=0 $Y2=0
cc_551 N_Z_M1005_s N_VGND_c_957_n 0.00225186f $X=6.24 $Y=0.235 $X2=0 $Y2=0
cc_552 N_Z_M1015_s N_VGND_c_957_n 0.00225186f $X=7.1 $Y=0.235 $X2=0 $Y2=0
cc_553 N_Z_M1019_s N_VGND_c_957_n 0.00225186f $X=7.96 $Y=0.235 $X2=0 $Y2=0
cc_554 N_Z_c_861_n N_A_305_47#_M1002_d 0.003322f $X=6.215 $Y=1.78 $X2=0 $Y2=0
cc_555 N_Z_M1000_s N_A_305_47#_c_1125_n 0.00329623f $X=5.38 $Y=0.235 $X2=0 $Y2=0
cc_556 N_Z_M1005_s N_A_305_47#_c_1125_n 0.00329237f $X=6.24 $Y=0.235 $X2=0 $Y2=0
cc_557 N_Z_c_861_n N_A_305_47#_c_1125_n 0.0483298f $X=6.215 $Y=1.78 $X2=0 $Y2=0
cc_558 N_Z_c_860_n N_A_305_47#_c_1125_n 0.0158479f $X=8.1 $Y=1.282 $X2=0 $Y2=0
cc_559 N_Z_M1015_s N_A_305_47#_c_1130_n 0.00332344f $X=7.1 $Y=0.235 $X2=0 $Y2=0
cc_560 N_Z_c_858_n N_A_305_47#_c_1130_n 0.0126348f $X=7.24 $Y=0.76 $X2=0 $Y2=0
cc_561 N_Z_M1019_s N_A_305_47#_c_1070_n 0.00332344f $X=7.96 $Y=0.235 $X2=0 $Y2=0
cc_562 N_Z_c_859_n N_A_305_47#_c_1070_n 0.0126348f $X=8.1 $Y=0.76 $X2=0 $Y2=0
cc_563 N_Z_c_859_n N_A_305_47#_c_1071_n 0.00152254f $X=8.1 $Y=0.76 $X2=0 $Y2=0
cc_564 N_Z_c_860_n N_A_305_47#_c_1135_n 0.0246504f $X=8.1 $Y=1.282 $X2=0 $Y2=0
cc_565 N_Z_c_860_n N_A_305_47#_c_1140_n 0.0246504f $X=8.1 $Y=1.282 $X2=0 $Y2=0
cc_566 N_VGND_c_957_n N_A_305_47#_M1004_s 0.00249946f $X=8.88 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_567 N_VGND_c_957_n N_A_305_47#_M1012_s 0.00293134f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_568 N_VGND_c_957_n N_A_305_47#_M1016_s 0.00293134f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_569 N_VGND_c_957_n N_A_305_47#_M1027_s 0.00293134f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_570 N_VGND_c_957_n N_A_305_47#_M1033_s 0.00254871f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_c_957_n N_A_305_47#_M1002_d 0.00223577f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_957_n N_A_305_47#_M1013_d 0.00223559f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_c_957_n N_A_305_47#_M1017_d 0.00223559f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_574 N_VGND_c_957_n N_A_305_47#_M1032_d 0.00211942f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_575 N_VGND_c_945_n N_A_305_47#_c_1060_n 0.0031603f $X=2.08 $Y=0.38 $X2=0
+ $Y2=0
cc_576 N_VGND_c_950_n N_A_305_47#_c_1060_n 0.0190529f $X=1.95 $Y=0 $X2=0 $Y2=0
cc_577 N_VGND_c_957_n N_A_305_47#_c_1060_n 0.0113912f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_578 N_VGND_c_945_n N_A_305_47#_c_1061_n 0.0211735f $X=2.08 $Y=0.38 $X2=0
+ $Y2=0
cc_579 N_VGND_c_945_n N_A_305_47#_c_1063_n 0.00313008f $X=2.08 $Y=0.38 $X2=0
+ $Y2=0
cc_580 N_VGND_c_946_n N_A_305_47#_c_1063_n 0.00313008f $X=2.94 $Y=0.38 $X2=0
+ $Y2=0
cc_581 N_VGND_c_952_n N_A_305_47#_c_1063_n 0.0149362f $X=2.81 $Y=0 $X2=0 $Y2=0
cc_582 N_VGND_c_957_n N_A_305_47#_c_1063_n 0.0100304f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_583 N_VGND_c_946_n N_A_305_47#_c_1064_n 0.0211735f $X=2.94 $Y=0.38 $X2=0
+ $Y2=0
cc_584 N_VGND_c_946_n N_A_305_47#_c_1065_n 0.00313008f $X=2.94 $Y=0.38 $X2=0
+ $Y2=0
cc_585 N_VGND_c_947_n N_A_305_47#_c_1065_n 0.00313008f $X=3.8 $Y=0.38 $X2=0
+ $Y2=0
cc_586 N_VGND_c_954_n N_A_305_47#_c_1065_n 0.0149362f $X=3.67 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_957_n N_A_305_47#_c_1065_n 0.0100304f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_947_n N_A_305_47#_c_1066_n 0.0211735f $X=3.8 $Y=0.38 $X2=0 $Y2=0
cc_589 N_VGND_c_947_n N_A_305_47#_c_1067_n 0.00313008f $X=3.8 $Y=0.38 $X2=0
+ $Y2=0
cc_590 N_VGND_c_948_n N_A_305_47#_c_1067_n 0.0149362f $X=4.53 $Y=0 $X2=0 $Y2=0
cc_591 N_VGND_c_949_n N_A_305_47#_c_1067_n 0.00313008f $X=4.66 $Y=0.38 $X2=0
+ $Y2=0
cc_592 N_VGND_c_957_n N_A_305_47#_c_1067_n 0.0100304f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_593 N_VGND_c_949_n N_A_305_47#_c_1068_n 0.0211735f $X=4.66 $Y=0.38 $X2=0
+ $Y2=0
cc_594 N_VGND_c_956_n N_A_305_47#_c_1200_n 0.0137653f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_c_957_n N_A_305_47#_c_1200_n 0.00874748f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_596 N_VGND_c_949_n N_A_305_47#_c_1069_n 0.00309615f $X=4.66 $Y=0.38 $X2=0
+ $Y2=0
cc_597 N_VGND_c_956_n N_A_305_47#_c_1125_n 0.0824976f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_c_957_n N_A_305_47#_c_1125_n 0.0525837f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_599 N_VGND_c_956_n N_A_305_47#_c_1130_n 0.0298674f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_600 N_VGND_c_957_n N_A_305_47#_c_1130_n 0.0187823f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_601 N_VGND_c_956_n N_A_305_47#_c_1070_n 0.0509189f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_c_957_n N_A_305_47#_c_1070_n 0.0313885f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_603 N_VGND_c_956_n N_A_305_47#_c_1135_n 0.0191147f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_957_n N_A_305_47#_c_1135_n 0.0124713f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_605 N_VGND_c_956_n N_A_305_47#_c_1140_n 0.0191147f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_606 N_VGND_c_957_n N_A_305_47#_c_1140_n 0.0124713f $X=8.88 $Y=0 $X2=0 $Y2=0
