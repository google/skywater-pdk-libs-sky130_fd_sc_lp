* File: sky130_fd_sc_lp__a311oi_0.pex.spice
* Created: Fri Aug 28 09:58:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311OI_0%A3 4 7 9 11 13 14 15 18 22 24 25 26 31
r43 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.525
+ $Y=1.245 $X2=0.525 $Y2=1.245
r44 25 26 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r45 25 32 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=0.64 $Y=1.295 $X2=0.64
+ $Y2=1.245
r46 24 32 9.21954 $w=3.98e-07 $l=3.2e-07 $layer=LI1_cond $X=0.64 $Y=0.925
+ $X2=0.64 $Y2=1.245
r47 20 22 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.615 $Y=2.14
+ $X2=0.715 $Y2=2.14
r48 16 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.615 $Y=0.84
+ $X2=0.825 $Y2=0.84
r49 14 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.525 $Y=1.585
+ $X2=0.525 $Y2=1.245
r50 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.585
+ $X2=0.525 $Y2=1.75
r51 13 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.08
+ $X2=0.525 $Y2=1.245
r52 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.825 $Y=0.765
+ $X2=0.825 $Y2=0.84
r53 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.825 $Y=0.765
+ $X2=0.825 $Y2=0.445
r54 5 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.715 $Y=2.215
+ $X2=0.715 $Y2=2.14
r55 5 7 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.715 $Y=2.215 $X2=0.715
+ $Y2=2.685
r56 4 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=2.065
+ $X2=0.615 $Y2=2.14
r57 4 15 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=0.615 $Y=2.065
+ $X2=0.615 $Y2=1.75
r58 1 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=0.915
+ $X2=0.615 $Y2=0.84
r59 1 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=0.915
+ $X2=0.615 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_0%A2 3 7 11 12 13 14 15 16 22
c49 11 0 1.4009e-19 $X=1.095 $Y=1.66
c50 7 0 1.63173e-19 $X=1.185 $Y=0.445
r51 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.095
+ $Y=1.32 $X2=1.095 $Y2=1.32
r52 16 23 13.0358 $w=3.03e-07 $l=3.45e-07 $layer=LI1_cond $X=1.162 $Y=1.665
+ $X2=1.162 $Y2=1.32
r53 15 23 0.944625 $w=3.03e-07 $l=2.5e-08 $layer=LI1_cond $X=1.162 $Y=1.295
+ $X2=1.162 $Y2=1.32
r54 14 15 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=1.162 $Y=0.925
+ $X2=1.162 $Y2=1.295
r55 13 14 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=1.162 $Y=0.555
+ $X2=1.162 $Y2=0.925
r56 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.095 $Y=1.66
+ $X2=1.095 $Y2=1.32
r57 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.66
+ $X2=1.095 $Y2=1.825
r58 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.155
+ $X2=1.095 $Y2=1.32
r59 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.185 $Y=0.445
+ $X2=1.185 $Y2=1.155
r60 3 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.145 $Y=2.685
+ $X2=1.145 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_0%A1 3 7 11 12 13 14 18
c41 11 0 1.4009e-19 $X=1.635 $Y=1.66
r42 13 14 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.652 $Y=1.295
+ $X2=1.652 $Y2=1.665
r43 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.635
+ $Y=1.32 $X2=1.635 $Y2=1.32
r44 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.635 $Y=1.66
+ $X2=1.635 $Y2=1.32
r45 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.66
+ $X2=1.635 $Y2=1.825
r46 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.155
+ $X2=1.635 $Y2=1.32
r47 7 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.575 $Y=2.685
+ $X2=1.575 $Y2=1.825
r48 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.545 $Y=0.445
+ $X2=1.545 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_0%B1 3 7 10 12 13 14 15 16 17 18 25 27 34
c58 15 0 1.21381e-19 $X=2.16 $Y=1.295
r59 28 34 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=2.155 $Y=1.695
+ $X2=2.155 $Y2=1.665
r60 25 27 35.3006 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.24
+ $X2=2.205 $Y2=1.075
r61 17 18 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.192 $Y=2.035
+ $X2=2.192 $Y2=2.405
r62 17 42 7.90892 $w=2.53e-07 $l=1.75e-07 $layer=LI1_cond $X=2.192 $Y=2.035
+ $X2=2.192 $Y2=1.86
r63 16 42 5.44459 $w=3.28e-07 $l=1.38e-07 $layer=LI1_cond $X=2.155 $Y=1.722
+ $X2=2.155 $Y2=1.86
r64 16 28 0.942908 $w=3.28e-07 $l=2.7e-08 $layer=LI1_cond $X=2.155 $Y=1.722
+ $X2=2.155 $Y2=1.695
r65 16 34 0.97783 $w=3.28e-07 $l=2.8e-08 $layer=LI1_cond $X=2.155 $Y=1.637
+ $X2=2.155 $Y2=1.665
r66 15 16 13.8642 $w=3.28e-07 $l=3.97e-07 $layer=LI1_cond $X=2.155 $Y=1.24
+ $X2=2.155 $Y2=1.637
r67 15 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.235
+ $Y=1.24 $X2=2.235 $Y2=1.24
r68 13 27 50.526 $w=2.1e-07 $l=1.6e-07 $layer=POLY_cond $X=2.115 $Y=0.915
+ $X2=2.115 $Y2=1.075
r69 12 13 52.88 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=2.075 $Y=0.765
+ $X2=2.075 $Y2=0.915
r70 10 14 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.085 $Y=2.685 $X2=2.085
+ $Y2=1.745
r71 7 14 49.7341 $w=3.9e-07 $l=1.95e-07 $layer=POLY_cond $X=2.205 $Y=1.55
+ $X2=2.205 $Y2=1.745
r72 6 25 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=2.205 $Y=1.27 $X2=2.205
+ $Y2=1.24
r73 6 7 39.929 $w=3.9e-07 $l=2.8e-07 $layer=POLY_cond $X=2.205 $Y=1.27 $X2=2.205
+ $Y2=1.55
r74 3 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.005 $Y=0.445
+ $X2=2.005 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_0%C1 3 6 9 15 16 17 22
c36 22 0 1.21381e-19 $X=2.775 $Y=1.63
r37 22 24 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.63
+ $X2=2.805 $Y2=1.465
r38 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.775
+ $Y=1.63 $X2=2.775 $Y2=1.63
r39 16 17 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.675 $Y=1.665
+ $X2=2.675 $Y2=2.035
r40 16 23 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=1.665
+ $X2=2.675 $Y2=1.63
r41 15 23 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.675 $Y=1.295
+ $X2=2.675 $Y2=1.63
r42 9 24 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.775 $Y=0.445
+ $X2=2.775 $Y2=1.465
r43 6 11 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.805 $Y=2.06
+ $X2=2.445 $Y2=2.06
r44 5 22 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=2.805 $Y=1.66 $X2=2.805
+ $Y2=1.63
r45 5 6 46.3462 $w=3.9e-07 $l=3.25e-07 $layer=POLY_cond $X=2.805 $Y=1.66
+ $X2=2.805 $Y2=1.985
r46 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.445 $Y=2.135
+ $X2=2.445 $Y2=2.06
r47 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.445 $Y=2.135
+ $X2=2.445 $Y2=2.685
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_0%VPWR 1 2 9 13 16 17 19 20 21 34 35
r37 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 21 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 21 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 19 28 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.23 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 19 20 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.23 $Y=3.33
+ $X2=1.365 $Y2=3.33
r47 18 31 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.5 $Y=3.33 $X2=1.68
+ $Y2=3.33
r48 18 20 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.5 $Y=3.33
+ $X2=1.365 $Y2=3.33
r49 16 24 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.335 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 16 17 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.335 $Y=3.33
+ $X2=0.482 $Y2=3.33
r51 15 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.63 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 15 17 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.63 $Y=3.33
+ $X2=0.482 $Y2=3.33
r53 11 20 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=3.245
+ $X2=1.365 $Y2=3.33
r54 11 13 31.3721 $w=2.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.365 $Y=3.245
+ $X2=1.365 $Y2=2.51
r55 7 17 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.482 $Y=3.245
+ $X2=0.482 $Y2=3.33
r56 7 9 28.3228 $w=2.93e-07 $l=7.25e-07 $layer=LI1_cond $X=0.482 $Y=3.245
+ $X2=0.482 $Y2=2.52
r57 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=2.365 $X2=1.36 $Y2=2.51
r58 1 9 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.375
+ $Y=2.365 $X2=0.5 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_0%A_158_473# 1 2 9 11 12 15
r31 13 15 17.1586 $w=2.23e-07 $l=3.35e-07 $layer=LI1_cond $X=1.782 $Y=2.175
+ $X2=1.782 $Y2=2.51
r32 11 13 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=1.67 $Y=2.09
+ $X2=1.782 $Y2=2.175
r33 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.67 $Y=2.09
+ $X2=1.06 $Y2=2.09
r34 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.93 $Y=2.175
+ $X2=1.06 $Y2=2.09
r35 7 9 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=0.93 $Y=2.175
+ $X2=0.93 $Y2=2.51
r36 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.65
+ $Y=2.365 $X2=1.79 $Y2=2.51
r37 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.79
+ $Y=2.365 $X2=0.93 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_0%Y 1 2 3 12 14 15 16 17 18 19 20 21 34 41 57
c47 15 0 1.63173e-19 $X=1.92 $Y=0.82
r48 39 57 6.80322 $w=2.45e-07 $l=3.4e-07 $layer=LI1_cond $X=3.152 $Y=2.345
+ $X2=3.152 $Y2=2.685
r49 38 41 0.94077 $w=2.43e-07 $l=2e-08 $layer=LI1_cond $X=3.152 $Y=0.905
+ $X2=3.152 $Y2=0.925
r50 21 57 0.56286 $w=6.78e-07 $l=3.2e-08 $layer=LI1_cond $X=3.12 $Y=2.685
+ $X2=3.152 $Y2=2.685
r51 21 52 8.09112 $w=6.78e-07 $l=4.6e-07 $layer=LI1_cond $X=3.12 $Y=2.685
+ $X2=2.66 $Y2=2.685
r52 21 39 0.6115 $w=2.43e-07 $l=1.3e-08 $layer=LI1_cond $X=3.152 $Y=2.332
+ $X2=3.152 $Y2=2.345
r53 20 21 13.9704 $w=2.43e-07 $l=2.97e-07 $layer=LI1_cond $X=3.152 $Y=2.035
+ $X2=3.152 $Y2=2.332
r54 19 20 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.152 $Y=1.665
+ $X2=3.152 $Y2=2.035
r55 18 19 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.152 $Y=1.295
+ $X2=3.152 $Y2=1.665
r56 17 32 2.86771 $w=3.32e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=0.82
+ $X2=3.065 $Y2=0.735
r57 17 38 2.86771 $w=3.32e-07 $l=1.22327e-07 $layer=LI1_cond $X=3.065 $Y=0.82
+ $X2=3.152 $Y2=0.905
r58 17 18 15.899 $w=2.43e-07 $l=3.38e-07 $layer=LI1_cond $X=3.152 $Y=0.957
+ $X2=3.152 $Y2=1.295
r59 17 41 1.50523 $w=2.43e-07 $l=3.2e-08 $layer=LI1_cond $X=3.152 $Y=0.957
+ $X2=3.152 $Y2=0.925
r60 16 32 4.93904 $w=4.18e-07 $l=1.8e-07 $layer=LI1_cond $X=3.065 $Y=0.555
+ $X2=3.065 $Y2=0.735
r61 16 34 3.0183 $w=4.18e-07 $l=1.1e-07 $layer=LI1_cond $X=3.065 $Y=0.555
+ $X2=3.065 $Y2=0.445
r62 14 17 3.83825 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.855 $Y=0.82
+ $X2=3.065 $Y2=0.82
r63 14 15 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.855 $Y=0.82 $X2=1.92
+ $Y2=0.82
r64 10 15 7.72402 $w=1.7e-07 $l=2.01057e-07 $layer=LI1_cond $X=1.757 $Y=0.735
+ $X2=1.92 $Y2=0.82
r65 10 12 10.2833 $w=3.23e-07 $l=2.9e-07 $layer=LI1_cond $X=1.757 $Y=0.735
+ $X2=1.757 $Y2=0.445
r66 3 52 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.52
+ $Y=2.365 $X2=2.66 $Y2=2.51
r67 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.235 $X2=2.99 $Y2=0.445
r68 1 12 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=1.62
+ $Y=0.235 $X2=1.775 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_0%VGND 1 2 8 9 13 14 27 30
r39 29 30 9.74588 $w=6.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.56 $Y=0.24
+ $X2=2.685 $Y2=0.24
r40 25 29 7.36048 $w=6.48e-07 $l=4e-07 $layer=LI1_cond $X=2.16 $Y=0.24 $X2=2.56
+ $Y2=0.24
r41 25 27 8.73382 $w=6.48e-07 $l=7e-08 $layer=LI1_cond $X=2.16 $Y=0.24 $X2=2.09
+ $Y2=0.24
r42 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r43 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 20 22 2.15409 $w=6.23e-07 $l=1.1e-07 $layer=LI1_cond $X=0.61 $Y=0.262
+ $X2=0.72 $Y2=0.262
r45 18 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r46 17 20 7.24559 $w=6.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.262
+ $X2=0.61 $Y2=0.262
r47 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 14 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r49 13 30 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=2.685
+ $Y2=0
r50 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r51 9 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r52 9 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r53 8 22 8.35809 $w=6.23e-07 $l=2.88191e-07 $layer=LI1_cond $X=0.775 $Y=0
+ $X2=0.72 $Y2=0.262
r54 8 27 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=0.775 $Y=0 $X2=2.09
+ $Y2=0
r55 2 29 91 $w=1.7e-07 $l=5.56417e-07 $layer=licon1_NDIFF $count=2 $X=2.08
+ $Y=0.235 $X2=2.56 $Y2=0.4
r56 1 20 91 $w=1.7e-07 $l=5.60245e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.61 $Y2=0.445
.ends

