# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__fa_m
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__fa_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.265000 2.495000 0.465000 ;
        RECT 1.115000 0.465000 2.245000 0.640000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 2.340000 2.305000 2.510000 ;
        RECT 1.085000 2.510000 1.415000 2.875000 ;
        RECT 2.135000 2.510000 2.305000 2.615000 ;
        RECT 2.135000 2.615000 3.690000 2.825000 ;
        RECT 2.135000 2.825000 6.515000 2.995000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 2.690000 1.955000 3.065000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 0.695000 0.520000 1.025000 ;
        RECT 0.155000 1.025000 0.345000 2.860000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.100000 0.735000 7.525000 0.945000 ;
        RECT 7.335000 0.945000 7.525000 2.860000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.525000  1.205000 0.695000 1.365000 ;
      RECT 0.525000  1.365000 5.615000 1.535000 ;
      RECT 0.525000  2.005000 0.855000 3.245000 ;
      RECT 0.740000  0.085000 0.930000 0.935000 ;
      RECT 1.470000  0.835000 1.800000 1.365000 ;
      RECT 1.530000  1.535000 1.740000 2.145000 ;
      RECT 1.960000  1.715000 3.265000 1.885000 ;
      RECT 1.960000  1.885000 2.170000 2.145000 ;
      RECT 1.980000  0.835000 2.310000 1.015000 ;
      RECT 1.980000  1.015000 3.265000 1.185000 ;
      RECT 2.485000  2.065000 2.815000 2.265000 ;
      RECT 2.485000  2.265000 4.040000 2.425000 ;
      RECT 2.485000  2.425000 7.000000 2.435000 ;
      RECT 2.515000  0.645000 2.845000 0.835000 ;
      RECT 2.675000  0.085000 2.845000 0.645000 ;
      RECT 3.055000  0.735000 3.265000 1.015000 ;
      RECT 3.055000  1.885000 3.265000 2.085000 ;
      RECT 3.820000  0.085000 4.030000 0.905000 ;
      RECT 3.820000  2.065000 4.040000 2.265000 ;
      RECT 3.870000  2.435000 7.000000 2.595000 ;
      RECT 4.250000  0.705000 4.440000 1.005000 ;
      RECT 4.250000  1.005000 5.320000 1.175000 ;
      RECT 4.250000  1.715000 5.320000 1.885000 ;
      RECT 4.250000  1.885000 4.460000 2.245000 ;
      RECT 4.620000  0.085000 4.950000 0.825000 ;
      RECT 4.680000  2.065000 4.890000 2.425000 ;
      RECT 5.110000  1.885000 5.320000 2.245000 ;
      RECT 5.130000  0.705000 5.320000 1.005000 ;
      RECT 5.580000  0.705000 5.965000 1.035000 ;
      RECT 5.580000  1.915000 5.965000 2.245000 ;
      RECT 5.795000  1.035000 5.965000 1.125000 ;
      RECT 5.795000  1.125000 7.155000 1.295000 ;
      RECT 5.795000  1.295000 5.965000 1.915000 ;
      RECT 6.670000  2.125000 7.000000 2.425000 ;
      RECT 6.730000  0.085000 6.920000 0.905000 ;
      RECT 6.830000  2.595000 7.000000 3.245000 ;
      RECT 6.985000  1.295000 7.155000 1.795000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__fa_m
END LIBRARY
