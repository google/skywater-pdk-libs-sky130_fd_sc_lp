* File: sky130_fd_sc_lp__and3b_2.spice
* Created: Wed Sep  2 09:32:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and3b_2.pex.spice"
.subckt sky130_fd_sc_lp__and3b_2  VNB VPB A_N C B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_N_M1005_g N_A_27_137#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.127033 AS=0.1113 PD=0.96 PS=1.37 NRD=70.692 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_204_27#_M1009_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.254067 PD=1.12 PS=1.92 NRD=0 NRS=14.28 M=1 R=5.6 SA=75000.5
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1010 N_X_M1009_d N_A_204_27#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.327867 PD=1.12 PS=2.19333 NRD=0 NRS=17.136 M=1 R=5.6 SA=75001
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1003 A_489_137# N_C_M1003_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.163933 PD=0.63 PS=1.09667 NRD=14.28 NRS=95.796 M=1 R=2.8 SA=75002.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 A_561_137# N_B_M1006_g A_489_137# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75002.4 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_204_27#_M1007_d N_A_27_137#_M1007_g A_561_137# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0819 PD=1.41 PS=0.81 NRD=5.712 NRS=39.996 M=1 R=2.8
+ SA=75003 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_N_M1008_g N_A_27_137#_M1008_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.105 AS=0.1113 PD=0.835 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1008_d N_A_204_27#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.315 AS=0.1764 PD=2.505 PS=1.54 NRD=9.8894 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_204_27#_M1011_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.39375 AS=0.1764 PD=2.91 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1000 N_A_204_27#_M1000_d N_C_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.13125 PD=0.7 PS=0.97 NRD=0 NRS=180.57 M=1 R=2.8 SA=75002
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_A_204_27#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.07665 AS=0.0588 PD=0.785 PS=0.7 NRD=28.1316 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_204_27#_M1002_d N_A_27_137#_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.07665 PD=1.37 PS=0.785 NRD=0 NRS=11.7215 M=1 R=2.8
+ SA=75003 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__and3b_2.pxi.spice"
*
.ends
*
*
