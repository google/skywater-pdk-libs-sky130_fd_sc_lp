* File: sky130_fd_sc_lp__dlrtp_lp2.spice
* Created: Fri Aug 28 10:27:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrtp_lp2.pex.spice"
.subckt sky130_fd_sc_lp__dlrtp_lp2  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1016 A_114_122# N_D_M1016_g N_A_27_122#_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_D_M1004_g A_114_122# VNB NSHORT L=0.15 W=0.42
+ AD=0.103162 AS=0.0504 PD=1.095 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.4 A=0.063 P=1.14 MULT=1
MM1017 A_294_185# N_GATE_M1017_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.103162 PD=0.63 PS=1.095 NRD=14.28 NRS=54.456 M=1 R=2.8
+ SA=75000.4 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_256_405#_M1008_d N_GATE_M1008_g A_294_185# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 A_500_47# N_A_256_405#_M1021_g N_A_413_47#_M1021_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_256_405#_M1023_g A_500_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1010 A_658_47# N_A_27_122#_M1010_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1011 N_A_736_47#_M1011_d N_A_413_47#_M1011_g A_658_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1018 A_850_47# N_A_256_405#_M1018_g N_A_736_47#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_898_21#_M1015_g A_850_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.3024 AS=0.0504 PD=2.28 PS=0.66 NRD=124.284 NRS=18.564 M=1 R=2.8
+ SA=75002.3 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 A_1216_57# N_A_736_47#_M1002_g N_A_898_21#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_RESET_B_M1003_g A_1216_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1012 A_1380_57# N_A_898_21#_M1012_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_Q_M1013_d N_A_898_21#_M1013_g A_1380_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1022_d N_D_M1022_g N_A_27_122#_M1022_s VPB PHIGHVT L=0.25 W=1
+ AD=0.186125 AS=0.285 PD=1.43 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1014 N_A_256_405#_M1014_d N_GATE_M1014_g N_VPWR_M1022_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.186125 PD=2.57 PS=1.43 NRD=0 NRS=16.7253 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A_256_405#_M1001_g N_A_413_47#_M1001_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.405 AS=0.285 PD=1.81 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125005 A=0.25 P=2.5 MULT=1
MM1005 A_740_419# N_A_27_122#_M1005_g N_VPWR_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.405 PD=1.24 PS=1.81 NRD=12.7853 NRS=104.39 M=1 R=4 SA=125001
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1019 N_A_736_47#_M1019_d N_A_256_405#_M1019_g A_740_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125002
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1006 A_944_419# N_A_413_47#_M1006_g N_A_736_47#_M1019_d VPB PHIGHVT L=0.25 W=1
+ AD=0.125 AS=0.14 PD=1.25 PS=1.28 NRD=13.7703 NRS=0 M=1 R=4 SA=125002 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A_898_21#_M1009_g A_944_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.2275 AS=0.125 PD=1.455 PS=1.25 NRD=18.715 NRS=13.7703 M=1 R=4 SA=125003
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1020 N_A_898_21#_M1020_d N_A_736_47#_M1020_g N_VPWR_M1009_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.2275 PD=1.28 PS=1.455 NRD=0 NRS=15.7403 M=1 R=4 SA=125003
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_RESET_B_M1007_g N_A_898_21#_M1020_d VPB PHIGHVT L=0.25
+ W=1 AD=0.1625 AS=0.14 PD=1.325 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1000 N_Q_M1000_d N_A_898_21#_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.1625 PD=2.57 PS=1.325 NRD=0 NRS=8.8453 M=1 R=4 SA=125005
+ SB=125000 A=0.25 P=2.5 MULT=1
DX24_noxref VNB VPB NWDIODE A=14.7041 P=20.23
*
.include "sky130_fd_sc_lp__dlrtp_lp2.pxi.spice"
*
.ends
*
*
