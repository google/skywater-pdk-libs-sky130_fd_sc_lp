* File: sky130_fd_sc_lp__a32o_lp.spice
* Created: Fri Aug 28 10:01:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32o_lp.pex.spice"
.subckt sky130_fd_sc_lp__a32o_lp  VNB VPB B2 B1 A1 A2 A3 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1001 A_137_141# N_B2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.4
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_137_419#_M1010_d N_B1_M1010_g A_137_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1008 A_329_141# N_A1_M1008_g N_A_137_419#_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0882 PD=0.84 PS=0.84 NRD=44.28 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1011 A_443_141# N_A2_M1011_g A_329_141# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0882 PD=0.84 PS=0.84 NRD=44.28 NRS=44.28 M=1 R=2.8 SA=75001.7 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A3_M1009_g A_443_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.09975 AS=0.0882 PD=0.895 PS=0.84 NRD=24.276 NRS=44.28 M=1 R=2.8
+ SA=75002.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1005 A_682_141# N_A_137_419#_M1005_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.09975 PD=0.66 PS=0.895 NRD=18.564 NRS=31.428 M=1 R=2.8
+ SA=75002.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_137_419#_M1002_g A_682_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.1575 AS=0.0504 PD=1.59 PS=0.66 NRD=25.704 NRS=18.564 M=1 R=2.8 SA=75003.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1006 N_A_137_419#_M1006_d N_B2_M1006_g N_A_30_419#_M1006_s VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1000 N_A_30_419#_M1000_d N_B1_M1000_g N_A_137_419#_M1006_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_30_419#_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.18 AS=0.14 PD=1.36 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1012 N_A_30_419#_M1012_d N_A2_M1012_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.18 PD=1.28 PS=1.36 NRD=0 NRS=15.7403 M=1 R=4 SA=125002 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_A3_M1003_g N_A_30_419#_M1012_d VPB PHIGHVT L=0.25 W=1
+ AD=0.3825 AS=0.14 PD=1.765 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1004 N_X_M1004_d N_A_137_419#_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.3825 PD=2.57 PS=1.765 NRD=0 NRS=82.7203 M=1 R=4 SA=125003
+ SB=125000 A=0.25 P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__a32o_lp.pxi.spice"
*
.ends
*
*
