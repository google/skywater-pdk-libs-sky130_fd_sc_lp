# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a21boi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a21boi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.415000 5.165000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.030000 1.075000 5.605000 1.210000 ;
        RECT 3.030000 1.210000 6.605000 1.245000 ;
        RECT 3.030000 1.245000 3.315000 1.515000 ;
        RECT 5.335000 1.245000 6.605000 1.515000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.210000 0.805000 1.750000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.646400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275000 0.370000 1.485000 0.700000 ;
        RECT 1.315000 0.700000 1.485000 1.035000 ;
        RECT 1.315000 1.035000 2.860000 1.205000 ;
        RECT 1.505000 1.715000 2.860000 1.750000 ;
        RECT 1.505000 1.750000 2.725000 2.035000 ;
        RECT 1.505000 2.035000 1.765000 2.485000 ;
        RECT 2.135000 0.255000 2.365000 0.695000 ;
        RECT 2.135000 0.695000 4.885000 0.895000 ;
        RECT 2.135000 0.895000 2.860000 1.035000 ;
        RECT 2.435000 2.035000 2.725000 2.665000 ;
        RECT 2.545000 1.205000 2.860000 1.715000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.125000  1.920000 1.195000 2.090000 ;
      RECT 0.125000  2.090000 0.385000 3.075000 ;
      RECT 0.325000  0.255000 0.605000 0.870000 ;
      RECT 0.325000  0.870000 1.145000 1.040000 ;
      RECT 0.555000  2.260000 0.885000 3.245000 ;
      RECT 0.775000  0.085000 1.105000 0.690000 ;
      RECT 0.975000  1.040000 1.145000 1.375000 ;
      RECT 0.975000  1.375000 2.375000 1.545000 ;
      RECT 0.975000  1.545000 1.195000 1.920000 ;
      RECT 1.075000  2.260000 1.335000 2.665000 ;
      RECT 1.075000  2.665000 2.265000 2.835000 ;
      RECT 1.075000  2.835000 3.095000 3.075000 ;
      RECT 1.655000  0.085000 1.965000 0.865000 ;
      RECT 1.935000  2.205000 2.265000 2.665000 ;
      RECT 2.535000  0.085000 3.095000 0.525000 ;
      RECT 2.895000  1.920000 6.605000 1.925000 ;
      RECT 2.895000  1.925000 5.665000 2.090000 ;
      RECT 2.895000  2.090000 3.095000 2.835000 ;
      RECT 3.265000  0.255000 5.315000 0.525000 ;
      RECT 3.265000  2.260000 4.455000 2.495000 ;
      RECT 3.265000  2.495000 3.595000 3.245000 ;
      RECT 3.765000  2.665000 4.815000 3.065000 ;
      RECT 4.625000  2.090000 4.815000 2.665000 ;
      RECT 4.985000  2.260000 5.315000 3.245000 ;
      RECT 5.055000  0.525000 5.315000 0.735000 ;
      RECT 5.055000  0.735000 6.135000 0.905000 ;
      RECT 5.335000  1.685000 6.605000 1.920000 ;
      RECT 5.485000  0.085000 5.715000 0.565000 ;
      RECT 5.485000  2.090000 5.665000 3.075000 ;
      RECT 5.845000  2.105000 6.175000 3.245000 ;
      RECT 5.885000  0.255000 6.135000 0.735000 ;
      RECT 5.905000  0.905000 6.135000 1.040000 ;
      RECT 6.305000  0.085000 6.605000 1.040000 ;
      RECT 6.345000  1.925000 6.605000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__a21boi_4
END LIBRARY
