* File: sky130_fd_sc_lp__buf_2.spice
* Created: Wed Sep  2 09:34:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__buf_2.pex.spice"
.subckt sky130_fd_sc_lp__buf_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_X_M1000_d N_A_90_21#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1003 N_X_M1000_d N_A_90_21#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2786 PD=1.12 PS=2.09333 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1004 N_A_90_21#_M1004_d N_A_M1004_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1393 PD=1.37 PS=1.04667 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_90_21#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_X_M1001_d N_A_90_21#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.430588 PD=1.54 PS=2.58632 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1002 N_A_90_21#_M1002_d N_A_M1002_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.218712 PD=1.81 PS=1.31368 NRD=0 NRS=144.657 M=1 R=4.26667
+ SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__buf_2.pxi.spice"
*
.ends
*
*
