* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__decap_12 VGND VNB VPB VPWR
M1000 VGND VPWR VGND VNB nshort w=1e+06u l=4e+06u
+  ad=5.5e+11p pd=5.1e+06u as=0p ps=0u
M1001 VPWR VGND VPWR VPB phighvt w=1e+06u l=4e+06u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
.ends
