* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__inputiso1p_lp A SLEEP VGND VNB VPB VPWR X
X0 a_493_93# a_161_489# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_245_489# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_177_93# A a_161_489# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_161_489# SLEEP a_335_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_335_93# SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_161_489# a_493_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND A a_177_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_161_489# A a_245_489# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_161_489# a_493_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_493_367# a_161_489# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
