* File: sky130_fd_sc_lp__o32ai_4.pxi.spice
* Created: Wed Sep  2 10:26:57 2020
* 
x_PM_SKY130_FD_SC_LP__O32AI_4%B2 N_B2_M1003_g N_B2_M1006_g N_B2_M1018_g
+ N_B2_M1014_g N_B2_M1020_g N_B2_M1025_g N_B2_M1027_g N_B2_M1028_g B2 B2 B2 B2
+ N_B2_c_145_n N_B2_c_146_n PM_SKY130_FD_SC_LP__O32AI_4%B2
x_PM_SKY130_FD_SC_LP__O32AI_4%B1 N_B1_M1001_g N_B1_M1013_g N_B1_M1015_g
+ N_B1_M1023_g N_B1_M1024_g N_B1_M1029_g N_B1_M1039_g N_B1_M1037_g B1 B1 B1 B1
+ N_B1_c_228_n PM_SKY130_FD_SC_LP__O32AI_4%B1
x_PM_SKY130_FD_SC_LP__O32AI_4%A3 N_A3_M1009_g N_A3_M1021_g N_A3_M1002_g
+ N_A3_M1008_g N_A3_M1031_g N_A3_M1030_g N_A3_M1034_g N_A3_M1033_g A3 A3 A3 A3
+ N_A3_c_317_n PM_SKY130_FD_SC_LP__O32AI_4%A3
x_PM_SKY130_FD_SC_LP__O32AI_4%A2 N_A2_M1005_g N_A2_c_403_n N_A2_M1004_g
+ N_A2_M1016_g N_A2_c_405_n N_A2_M1010_g N_A2_M1022_g N_A2_c_407_n N_A2_M1019_g
+ N_A2_M1038_g N_A2_c_409_n N_A2_c_410_n N_A2_c_411_n N_A2_M1032_g A2 A2 A2 A2
+ N_A2_c_412_n PM_SKY130_FD_SC_LP__O32AI_4%A2
x_PM_SKY130_FD_SC_LP__O32AI_4%A1 N_A1_c_486_n N_A1_M1007_g N_A1_M1000_g
+ N_A1_c_487_n N_A1_M1011_g N_A1_M1012_g N_A1_c_488_n N_A1_M1035_g N_A1_M1017_g
+ N_A1_c_489_n N_A1_M1036_g N_A1_M1026_g A1 A1 A1 A1 N_A1_c_491_n N_A1_c_492_n
+ PM_SKY130_FD_SC_LP__O32AI_4%A1
x_PM_SKY130_FD_SC_LP__O32AI_4%A_30_367# N_A_30_367#_M1006_d N_A_30_367#_M1014_d
+ N_A_30_367#_M1028_d N_A_30_367#_M1023_s N_A_30_367#_M1037_s
+ N_A_30_367#_c_555_n N_A_30_367#_c_556_n N_A_30_367#_c_560_n
+ N_A_30_367#_c_573_p N_A_30_367#_c_562_n N_A_30_367#_c_578_p
+ N_A_30_367#_c_564_n N_A_30_367#_c_565_n N_A_30_367#_c_567_n
+ N_A_30_367#_c_593_p N_A_30_367#_c_581_p N_A_30_367#_c_557_n
+ PM_SKY130_FD_SC_LP__O32AI_4%A_30_367#
x_PM_SKY130_FD_SC_LP__O32AI_4%Y N_Y_M1003_d N_Y_M1020_d N_Y_M1001_d N_Y_M1024_d
+ N_Y_M1006_s N_Y_M1025_s N_Y_M1002_d N_Y_M1030_d N_Y_c_740_p N_Y_c_609_n
+ N_Y_c_610_n N_Y_c_627_n N_Y_c_744_p N_Y_c_611_n N_Y_c_748_p N_Y_c_612_n
+ N_Y_c_752_p N_Y_c_613_n N_Y_c_677_n N_Y_c_681_n N_Y_c_614_n N_Y_c_633_n
+ N_Y_c_615_n N_Y_c_616_n N_Y_c_617_n N_Y_c_619_n N_Y_c_691_n N_Y_c_693_n Y Y
+ PM_SKY130_FD_SC_LP__O32AI_4%Y
x_PM_SKY130_FD_SC_LP__O32AI_4%VPWR N_VPWR_M1013_d N_VPWR_M1029_d N_VPWR_M1000_d
+ N_VPWR_M1012_d N_VPWR_M1026_d N_VPWR_c_770_n N_VPWR_c_771_n N_VPWR_c_772_n
+ N_VPWR_c_773_n N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n N_VPWR_c_777_n
+ N_VPWR_c_778_n N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n
+ N_VPWR_c_783_n N_VPWR_c_784_n VPWR N_VPWR_c_785_n N_VPWR_c_769_n
+ PM_SKY130_FD_SC_LP__O32AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O32AI_4%A_829_349# N_A_829_349#_M1002_s
+ N_A_829_349#_M1008_s N_A_829_349#_M1033_s N_A_829_349#_M1016_d
+ N_A_829_349#_M1038_d N_A_829_349#_c_896_n N_A_829_349#_c_897_n
+ N_A_829_349#_c_898_n N_A_829_349#_c_928_n N_A_829_349#_c_899_n
+ N_A_829_349#_c_931_n N_A_829_349#_c_900_n N_A_829_349#_c_954_p
+ N_A_829_349#_c_901_n N_A_829_349#_c_902_n N_A_829_349#_c_903_n
+ N_A_829_349#_c_904_n N_A_829_349#_c_905_n
+ PM_SKY130_FD_SC_LP__O32AI_4%A_829_349#
x_PM_SKY130_FD_SC_LP__O32AI_4%A_1256_349# N_A_1256_349#_M1005_s
+ N_A_1256_349#_M1022_s N_A_1256_349#_M1000_s N_A_1256_349#_M1017_s
+ N_A_1256_349#_c_996_n N_A_1256_349#_c_958_n N_A_1256_349#_c_959_n
+ N_A_1256_349#_c_999_n N_A_1256_349#_c_960_n N_A_1256_349#_c_988_n
+ N_A_1256_349#_c_961_n N_A_1256_349#_c_992_n N_A_1256_349#_c_962_n
+ N_A_1256_349#_c_982_n PM_SKY130_FD_SC_LP__O32AI_4%A_1256_349#
x_PM_SKY130_FD_SC_LP__O32AI_4%A_30_47# N_A_30_47#_M1003_s N_A_30_47#_M1018_s
+ N_A_30_47#_M1027_s N_A_30_47#_M1015_s N_A_30_47#_M1039_s N_A_30_47#_M1021_s
+ N_A_30_47#_M1034_s N_A_30_47#_M1010_s N_A_30_47#_M1032_s N_A_30_47#_M1011_d
+ N_A_30_47#_M1036_d N_A_30_47#_c_1003_n N_A_30_47#_c_1010_n N_A_30_47#_c_1004_n
+ N_A_30_47#_c_1012_n N_A_30_47#_c_1020_n N_A_30_47#_c_1022_n
+ N_A_30_47#_c_1024_n N_A_30_47#_c_1025_n N_A_30_47#_c_1036_n
+ N_A_30_47#_c_1027_n N_A_30_47#_c_1038_n N_A_30_47#_c_1040_n
+ N_A_30_47#_c_1041_n N_A_30_47#_c_1049_n N_A_30_47#_c_1135_p
+ N_A_30_47#_c_1053_n N_A_30_47#_c_1130_p N_A_30_47#_c_1061_n
+ N_A_30_47#_c_1131_p N_A_30_47#_c_1005_n N_A_30_47#_c_1006_n
+ N_A_30_47#_c_1014_n N_A_30_47#_c_1018_n N_A_30_47#_c_1030_n
+ N_A_30_47#_c_1042_n N_A_30_47#_c_1043_n N_A_30_47#_c_1057_n
+ N_A_30_47#_c_1059_n N_A_30_47#_c_1070_n PM_SKY130_FD_SC_LP__O32AI_4%A_30_47#
x_PM_SKY130_FD_SC_LP__O32AI_4%VGND N_VGND_M1009_d N_VGND_M1031_d N_VGND_M1004_d
+ N_VGND_M1019_d N_VGND_M1007_s N_VGND_M1035_s N_VGND_c_1167_n N_VGND_c_1168_n
+ N_VGND_c_1169_n N_VGND_c_1170_n N_VGND_c_1171_n N_VGND_c_1172_n
+ N_VGND_c_1173_n N_VGND_c_1174_n N_VGND_c_1175_n N_VGND_c_1176_n
+ N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n VGND N_VGND_c_1180_n
+ N_VGND_c_1181_n N_VGND_c_1182_n N_VGND_c_1183_n N_VGND_c_1184_n
+ N_VGND_c_1185_n PM_SKY130_FD_SC_LP__O32AI_4%VGND
cc_1 VNB N_B2_M1003_g 0.0303823f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_2 VNB N_B2_M1006_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_3 VNB N_B2_M1018_g 0.0209293f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.655
cc_4 VNB N_B2_M1014_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_5 VNB N_B2_M1020_g 0.0209293f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_6 VNB N_B2_M1025_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_7 VNB N_B2_M1027_g 0.0211935f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_8 VNB N_B2_M1028_g 0.00114276f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_9 VNB N_B2_c_145_n 0.0135836f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.46
cc_10 VNB N_B2_c_146_n 0.104193f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.46
cc_11 VNB N_B1_M1001_g 0.0238213f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_12 VNB N_B1_M1015_g 0.0234721f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.655
cc_13 VNB N_B1_M1024_g 0.0234721f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_14 VNB N_B1_M1039_g 0.0254637f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_15 VNB B1 0.00317876f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_16 VNB N_B1_c_228_n 0.0775041f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.567
cc_17 VNB N_A3_M1009_g 0.0201802f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_18 VNB N_A3_M1021_g 0.0196169f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_19 VNB N_A3_M1031_g 0.0206533f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_20 VNB N_A3_M1034_g 0.024446f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_21 VNB A3 0.00260128f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_22 VNB N_A3_c_317_n 0.0889009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_M1005_g 0.00256042f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_24 VNB N_A2_c_403_n 0.0193166f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.625
cc_25 VNB N_A2_M1016_g 0.00249068f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.655
cc_26 VNB N_A2_c_405_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A2_M1022_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.295
cc_28 VNB N_A2_c_407_n 0.018931f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_29 VNB N_A2_M1038_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A2_c_409_n 0.0293414f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_31 VNB N_A2_c_410_n 0.0794657f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_32 VNB N_A2_c_411_n 0.0419057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A2_c_412_n 0.00189034f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.46
cc_34 VNB N_A1_c_486_n 0.0166505f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.295
cc_35 VNB N_A1_c_487_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A1_c_488_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_37 VNB N_A1_c_489_n 0.0218823f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_38 VNB A1 0.0134162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A1_c_491_n 0.0760484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A1_c_492_n 0.0984116f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.46
cc_41 VNB N_Y_c_609_n 0.00322376f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_42 VNB N_Y_c_610_n 0.0032169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_611_n 0.0085839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_612_n 0.00351696f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.46
cc_45 VNB N_Y_c_613_n 0.0196465f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.46
cc_46 VNB N_Y_c_614_n 0.0037417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_615_n 0.00150375f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.567
cc_48 VNB N_Y_c_616_n 0.00164567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_Y_c_617_n 0.00206898f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.567
cc_50 VNB N_VPWR_c_769_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_30_47#_c_1003_n 0.0294275f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_52 VNB N_A_30_47#_c_1004_n 0.00746637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_30_47#_c_1005_n 0.00740486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_30_47#_c_1006_n 0.0233935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1167_n 4.2118e-19 $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.625
cc_56 VNB N_VGND_c_1168_n 0.00225941f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.295
cc_57 VNB N_VGND_c_1169_n 4.05289e-19 $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.625
cc_58 VNB N_VGND_c_1170_n 3.22457e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_59 VNB N_VGND_c_1171_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1172_n 0.0937972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1173_n 0.00436274f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.46
cc_62 VNB N_VGND_c_1174_n 0.0155317f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.46
cc_63 VNB N_VGND_c_1175_n 0.00509914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1176_n 0.0158116f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.46
cc_65 VNB N_VGND_c_1177_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.46
cc_66 VNB N_VGND_c_1178_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.46
cc_67 VNB N_VGND_c_1179_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.46
cc_68 VNB N_VGND_c_1180_n 0.0219286f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.567
cc_69 VNB N_VGND_c_1181_n 0.0148029f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.567
cc_70 VNB N_VGND_c_1182_n 0.0247634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1183_n 0.501448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1184_n 0.00449511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1185_n 0.0181368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VPB N_B2_M1006_g 0.0254418f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_75 VPB N_B2_M1014_g 0.0189466f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_76 VPB N_B2_M1025_g 0.0189466f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_77 VPB N_B2_M1028_g 0.0194637f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_78 VPB N_B2_c_145_n 0.0165558f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.46
cc_79 VPB N_B1_M1013_g 0.0184325f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_80 VPB N_B1_M1023_g 0.0178551f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_81 VPB N_B1_M1029_g 0.0178551f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_82 VPB N_B1_M1037_g 0.0240279f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_83 VPB B1 0.0116982f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_84 VPB N_B1_c_228_n 0.0199687f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.567
cc_85 VPB N_A3_M1002_g 0.0217292f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.655
cc_86 VPB N_A3_M1008_g 0.0173999f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_87 VPB N_A3_M1030_g 0.0174041f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_88 VPB N_A3_M1033_g 0.0180953f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_89 VPB A3 0.003845f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_90 VPB N_A3_c_317_n 0.0257471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A2_M1005_g 0.0201136f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.655
cc_92 VPB N_A2_M1016_g 0.0191384f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.655
cc_93 VPB N_A2_M1022_g 0.0191411f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.295
cc_94 VPB N_A2_M1038_g 0.0255214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A1_M1000_g 0.0221774f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_96 VPB N_A1_M1012_g 0.017618f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.625
cc_97 VPB N_A1_M1017_g 0.017618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A1_M1026_g 0.026336f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=0.655
cc_99 VPB N_A1_c_492_n 0.0107279f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.46
cc_100 VPB N_A_30_367#_c_555_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_30_367#_c_556_n 0.0378712f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=0.655
cc_102 VPB N_A_30_367#_c_557_n 0.00782378f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.46
cc_103 VPB N_Y_c_614_n 0.00148593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_Y_c_619_n 0.0132426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_770_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.35 $Y2=0.655
cc_106 VPB N_VPWR_c_771_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_107 VPB N_VPWR_c_772_n 0.0138448f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=0.655
cc_108 VPB N_VPWR_c_773_n 3.16049e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_774_n 0.0559723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_775_n 0.0546648f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.46
cc_111 VPB N_VPWR_c_776_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_777_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.46
cc_113 VPB N_VPWR_c_778_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.46
cc_114 VPB N_VPWR_c_779_n 0.10748f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.46
cc_115 VPB N_VPWR_c_780_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.46
cc_116 VPB N_VPWR_c_781_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.46
cc_117 VPB N_VPWR_c_782_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.46
cc_118 VPB N_VPWR_c_783_n 0.0148832f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.46
cc_119 VPB N_VPWR_c_784_n 0.00555219f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=1.46
cc_120 VPB N_VPWR_c_785_n 0.0145539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_769_n 0.0948618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_829_349#_c_896_n 0.00593693f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=0.655
cc_123 VPB N_A_829_349#_c_897_n 0.00223571f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_829_349#_c_898_n 0.0037234f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.625
cc_125 VPB N_A_829_349#_c_899_n 0.00216451f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=0.655
cc_126 VPB N_A_829_349#_c_900_n 0.00205771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_829_349#_c_901_n 0.00621886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_829_349#_c_902_n 0.00910797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_829_349#_c_903_n 0.00185632f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.46
cc_130 VPB N_A_829_349#_c_904_n 0.00196551f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.46
cc_131 VPB N_A_829_349#_c_905_n 0.00189272f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.46
cc_132 VPB N_A_1256_349#_c_958_n 0.00237782f $X=-0.19 $Y=1.655 $X2=1.35
+ $Y2=0.655
cc_133 VPB N_A_1256_349#_c_959_n 0.00285182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_1256_349#_c_960_n 0.0235224f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=0.655
cc_135 VPB N_A_1256_349#_c_961_n 0.0109075f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_136 VPB N_A_1256_349#_c_962_n 0.00215817f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.46
cc_137 N_B2_M1027_g N_B1_M1001_g 0.0264707f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_138 N_B2_M1028_g N_B1_M1013_g 0.0314921f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_139 N_B2_M1028_g B1 3.64523e-19 $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_140 N_B2_c_145_n B1 0.0241139f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_141 N_B2_c_146_n B1 3.09501e-19 $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_142 N_B2_c_145_n N_B1_c_228_n 6.89561e-19 $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_143 N_B2_c_146_n N_B1_c_228_n 0.0221693f $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_144 N_B2_c_145_n N_A_30_367#_c_556_n 0.0175239f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_145 N_B2_c_146_n N_A_30_367#_c_556_n 0.00113953f $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_146 N_B2_M1006_g N_A_30_367#_c_560_n 0.0115031f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B2_M1014_g N_A_30_367#_c_560_n 0.0115031f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_148 N_B2_M1025_g N_A_30_367#_c_562_n 0.0114565f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_149 N_B2_M1028_g N_A_30_367#_c_562_n 0.0104327f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_150 N_B2_M1028_g N_A_30_367#_c_564_n 0.00446092f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_151 N_B2_M1018_g N_Y_c_609_n 0.0119717f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_152 N_B2_M1020_g N_Y_c_609_n 0.0122536f $X=1.35 $Y=0.655 $X2=0 $Y2=0
cc_153 N_B2_c_145_n N_Y_c_609_n 0.043886f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_154 N_B2_c_146_n N_Y_c_609_n 0.00241702f $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_155 N_B2_M1003_g N_Y_c_610_n 0.0031967f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_156 N_B2_c_145_n N_Y_c_610_n 0.0171288f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_157 N_B2_c_146_n N_Y_c_610_n 0.00251039f $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_158 N_B2_M1014_g N_Y_c_627_n 0.01115f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B2_M1025_g N_Y_c_627_n 0.01115f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_160 N_B2_c_145_n N_Y_c_627_n 0.0359705f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_161 N_B2_c_146_n N_Y_c_627_n 5.04482e-19 $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_162 N_B2_M1027_g N_Y_c_611_n 0.0122536f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_163 N_B2_c_145_n N_Y_c_611_n 0.0125191f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_164 N_B2_M1006_g N_Y_c_633_n 0.0110566f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_165 N_B2_M1014_g N_Y_c_633_n 0.0101524f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_166 N_B2_M1025_g N_Y_c_633_n 5.66402e-19 $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_167 N_B2_c_145_n N_Y_c_633_n 0.0233849f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_168 N_B2_c_146_n N_Y_c_633_n 5.70981e-19 $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_169 N_B2_c_145_n N_Y_c_615_n 0.0141497f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_170 N_B2_c_146_n N_Y_c_615_n 0.00251039f $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_171 N_B2_M1028_g N_Y_c_619_n 0.00872087f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_172 N_B2_c_145_n N_Y_c_619_n 0.00647385f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_173 N_B2_M1014_g Y 5.65733e-19 $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_174 N_B2_M1025_g Y 0.0101524f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_175 N_B2_M1028_g Y 0.0135252f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_176 N_B2_c_145_n Y 0.0262103f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_177 N_B2_c_146_n Y 5.70981e-19 $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_178 N_B2_M1028_g N_VPWR_c_770_n 0.00104138f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_179 N_B2_M1006_g N_VPWR_c_775_n 0.00357877f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_180 N_B2_M1014_g N_VPWR_c_775_n 0.00357877f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B2_M1025_g N_VPWR_c_775_n 0.00357877f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B2_M1028_g N_VPWR_c_775_n 0.00357877f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B2_M1006_g N_VPWR_c_769_n 0.00629771f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_184 N_B2_M1014_g N_VPWR_c_769_n 0.0053512f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_185 N_B2_M1025_g N_VPWR_c_769_n 0.0053512f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B2_M1028_g N_VPWR_c_769_n 0.0054589f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_187 N_B2_M1003_g N_A_30_47#_c_1003_n 0.00246707f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_188 N_B2_c_145_n N_A_30_47#_c_1003_n 0.0143788f $X=1.69 $Y=1.46 $X2=0 $Y2=0
cc_189 N_B2_c_146_n N_A_30_47#_c_1003_n 0.00564732f $X=1.78 $Y=1.46 $X2=0 $Y2=0
cc_190 N_B2_M1003_g N_A_30_47#_c_1010_n 0.012237f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_191 N_B2_M1018_g N_A_30_47#_c_1010_n 0.00836084f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_192 N_B2_M1020_g N_A_30_47#_c_1012_n 0.00836084f $X=1.35 $Y=0.655 $X2=0 $Y2=0
cc_193 N_B2_M1027_g N_A_30_47#_c_1012_n 0.00836084f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_194 N_B2_M1003_g N_A_30_47#_c_1014_n 5.10997e-19 $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_195 N_B2_M1018_g N_A_30_47#_c_1014_n 0.00639472f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_196 N_B2_M1020_g N_A_30_47#_c_1014_n 0.0062862f $X=1.35 $Y=0.655 $X2=0 $Y2=0
cc_197 N_B2_M1027_g N_A_30_47#_c_1014_n 5.02748e-19 $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_198 N_B2_M1020_g N_A_30_47#_c_1018_n 5.02748e-19 $X=1.35 $Y=0.655 $X2=0 $Y2=0
cc_199 N_B2_M1027_g N_A_30_47#_c_1018_n 0.0062862f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_200 N_B2_M1003_g N_VGND_c_1172_n 0.00357877f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_201 N_B2_M1018_g N_VGND_c_1172_n 0.00357842f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_202 N_B2_M1020_g N_VGND_c_1172_n 0.00357842f $X=1.35 $Y=0.655 $X2=0 $Y2=0
cc_203 N_B2_M1027_g N_VGND_c_1172_n 0.00357842f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_204 N_B2_M1003_g N_VGND_c_1183_n 0.00643216f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_205 N_B2_M1018_g N_VGND_c_1183_n 0.00535118f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_206 N_B2_M1020_g N_VGND_c_1183_n 0.00535118f $X=1.35 $Y=0.655 $X2=0 $Y2=0
cc_207 N_B2_M1027_g N_VGND_c_1183_n 0.00537652f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_208 N_B1_M1039_g N_A3_M1009_g 0.0272252f $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_209 B1 N_A3_M1002_g 3.46383e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_210 N_B1_c_228_n N_A3_M1002_g 0.0010129f $X=3.59 $Y=1.51 $X2=0 $Y2=0
cc_211 N_B1_M1037_g A3 4.72957e-19 $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_212 B1 A3 0.0249591f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_213 N_B1_c_228_n A3 0.00127015f $X=3.59 $Y=1.51 $X2=0 $Y2=0
cc_214 N_B1_c_228_n N_A3_c_317_n 0.0158253f $X=3.59 $Y=1.51 $X2=0 $Y2=0
cc_215 N_B1_M1013_g N_A_30_367#_c_565_n 0.0125619f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_216 N_B1_M1023_g N_A_30_367#_c_565_n 0.0125125f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_217 N_B1_M1029_g N_A_30_367#_c_567_n 0.0125619f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B1_M1037_g N_A_30_367#_c_567_n 0.0125619f $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_219 N_B1_M1001_g N_Y_c_611_n 0.0125413f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_220 B1 N_Y_c_611_n 0.0143378f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_221 N_B1_c_228_n N_Y_c_611_n 0.00163409f $X=3.59 $Y=1.51 $X2=0 $Y2=0
cc_222 N_B1_M1015_g N_Y_c_612_n 0.0125854f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_223 N_B1_M1024_g N_Y_c_612_n 0.0125072f $X=3.07 $Y=0.655 $X2=0 $Y2=0
cc_224 B1 N_Y_c_612_n 0.0365751f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B1_c_228_n N_Y_c_612_n 0.00247231f $X=3.59 $Y=1.51 $X2=0 $Y2=0
cc_226 N_B1_M1039_g N_Y_c_613_n 0.0130599f $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_227 B1 N_Y_c_613_n 0.0182894f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B1_c_228_n N_Y_c_613_n 0.00430806f $X=3.59 $Y=1.51 $X2=0 $Y2=0
cc_229 B1 N_Y_c_616_n 0.0118717f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_230 N_B1_c_228_n N_Y_c_616_n 0.0025758f $X=3.59 $Y=1.51 $X2=0 $Y2=0
cc_231 N_B1_M1039_g N_Y_c_617_n 3.32503e-19 $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_232 B1 N_Y_c_617_n 0.0135439f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B1_c_228_n N_Y_c_617_n 0.00257251f $X=3.59 $Y=1.51 $X2=0 $Y2=0
cc_234 N_B1_M1013_g N_Y_c_619_n 0.0106442f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_235 N_B1_M1023_g N_Y_c_619_n 0.0104926f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_236 N_B1_M1029_g N_Y_c_619_n 0.0104926f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B1_M1037_g N_Y_c_619_n 0.0125331f $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_238 B1 N_Y_c_619_n 0.111409f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_239 N_B1_c_228_n N_Y_c_619_n 0.00288353f $X=3.59 $Y=1.51 $X2=0 $Y2=0
cc_240 N_B1_M1013_g Y 7.94691e-19 $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B1_M1013_g N_VPWR_c_770_n 0.0118761f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B1_M1023_g N_VPWR_c_770_n 0.0106714f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B1_M1029_g N_VPWR_c_770_n 5.78645e-19 $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B1_M1023_g N_VPWR_c_771_n 5.78645e-19 $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B1_M1029_g N_VPWR_c_771_n 0.0106714f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B1_M1037_g N_VPWR_c_771_n 0.012364f $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B1_M1013_g N_VPWR_c_775_n 0.00486043f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B1_M1023_g N_VPWR_c_777_n 0.00486043f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_249 N_B1_M1029_g N_VPWR_c_777_n 0.00486043f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_250 N_B1_M1037_g N_VPWR_c_779_n 0.00486043f $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_251 N_B1_M1013_g N_VPWR_c_769_n 0.00835496f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_252 N_B1_M1023_g N_VPWR_c_769_n 0.00824727f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_253 N_B1_M1029_g N_VPWR_c_769_n 0.00824727f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_254 N_B1_M1037_g N_VPWR_c_769_n 0.00954696f $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_255 N_B1_M1001_g N_A_30_47#_c_1020_n 0.00836084f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_256 N_B1_M1015_g N_A_30_47#_c_1020_n 0.00836084f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_257 N_B1_M1024_g N_A_30_47#_c_1022_n 0.008789f $X=3.07 $Y=0.655 $X2=0 $Y2=0
cc_258 N_B1_M1039_g N_A_30_47#_c_1022_n 0.00875768f $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_259 N_B1_M1039_g N_A_30_47#_c_1024_n 6.34972e-19 $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_260 N_B1_M1024_g N_A_30_47#_c_1025_n 4.45884e-19 $X=3.07 $Y=0.655 $X2=0 $Y2=0
cc_261 N_B1_M1039_g N_A_30_47#_c_1025_n 0.0033428f $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_262 N_B1_M1039_g N_A_30_47#_c_1027_n 0.00207083f $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_263 N_B1_M1001_g N_A_30_47#_c_1018_n 0.00628588f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_264 N_B1_M1015_g N_A_30_47#_c_1018_n 5.02725e-19 $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_265 N_B1_M1001_g N_A_30_47#_c_1030_n 4.43872e-19 $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_266 N_B1_M1015_g N_A_30_47#_c_1030_n 0.00628722f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_267 N_B1_M1024_g N_A_30_47#_c_1030_n 0.0061293f $X=3.07 $Y=0.655 $X2=0 $Y2=0
cc_268 N_B1_M1039_g N_A_30_47#_c_1030_n 4.9709e-19 $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_269 N_B1_M1039_g N_VGND_c_1167_n 9.37539e-19 $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_270 N_B1_M1001_g N_VGND_c_1172_n 0.00357842f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_271 N_B1_M1015_g N_VGND_c_1172_n 0.00357842f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_272 N_B1_M1024_g N_VGND_c_1172_n 0.00357842f $X=3.07 $Y=0.655 $X2=0 $Y2=0
cc_273 N_B1_M1039_g N_VGND_c_1172_n 0.00357842f $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_274 N_B1_M1001_g N_VGND_c_1183_n 0.00537652f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_275 N_B1_M1015_g N_VGND_c_1183_n 0.00535118f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_276 N_B1_M1024_g N_VGND_c_1183_n 0.00535118f $X=3.07 $Y=0.655 $X2=0 $Y2=0
cc_277 N_B1_M1039_g N_VGND_c_1183_n 0.00561868f $X=3.5 $Y=0.655 $X2=0 $Y2=0
cc_278 N_A3_M1033_g N_A2_M1005_g 0.0242688f $X=5.775 $Y=2.375 $X2=0 $Y2=0
cc_279 N_A3_M1034_g N_A2_c_410_n 9.35895e-19 $X=5.47 $Y=0.655 $X2=0 $Y2=0
cc_280 N_A3_c_317_n N_A2_c_410_n 0.0242688f $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_281 N_A3_c_317_n N_A2_c_412_n 2.12391e-19 $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_282 N_A3_M1002_g N_A_30_367#_c_557_n 4.07938e-19 $X=4.485 $Y=2.375 $X2=0
+ $Y2=0
cc_283 A3 N_Y_M1002_d 0.00181504f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_284 A3 N_Y_M1030_d 0.00181948f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_285 N_A3_M1009_g N_Y_c_613_n 0.0110126f $X=4.04 $Y=0.655 $X2=0 $Y2=0
cc_286 N_A3_M1021_g N_Y_c_613_n 0.0108858f $X=4.47 $Y=0.655 $X2=0 $Y2=0
cc_287 N_A3_M1031_g N_Y_c_613_n 0.011278f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_288 N_A3_M1034_g N_Y_c_613_n 0.0125998f $X=5.47 $Y=0.655 $X2=0 $Y2=0
cc_289 A3 N_Y_c_613_n 0.127275f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_290 N_A3_c_317_n N_Y_c_613_n 0.0227189f $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_291 N_A3_M1008_g N_Y_c_677_n 0.0129934f $X=4.915 $Y=2.375 $X2=0 $Y2=0
cc_292 N_A3_M1030_g N_Y_c_677_n 0.0126248f $X=5.345 $Y=2.375 $X2=0 $Y2=0
cc_293 A3 N_Y_c_677_n 0.0476503f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_294 N_A3_c_317_n N_Y_c_677_n 4.6067e-19 $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_295 N_A3_M1008_g N_Y_c_681_n 5.57395e-19 $X=4.915 $Y=2.375 $X2=0 $Y2=0
cc_296 N_A3_M1030_g N_Y_c_681_n 0.00779921f $X=5.345 $Y=2.375 $X2=0 $Y2=0
cc_297 N_A3_M1030_g N_Y_c_614_n 8.89824e-19 $X=5.345 $Y=2.375 $X2=0 $Y2=0
cc_298 N_A3_M1034_g N_Y_c_614_n 0.00200076f $X=5.47 $Y=0.655 $X2=0 $Y2=0
cc_299 N_A3_M1033_g N_Y_c_614_n 0.007117f $X=5.775 $Y=2.375 $X2=0 $Y2=0
cc_300 A3 N_Y_c_614_n 0.0308557f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_301 N_A3_c_317_n N_Y_c_614_n 0.0102717f $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_302 N_A3_M1002_g N_Y_c_619_n 0.015034f $X=4.485 $Y=2.375 $X2=0 $Y2=0
cc_303 A3 N_Y_c_619_n 0.0416794f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_304 N_A3_c_317_n N_Y_c_619_n 0.00195452f $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_305 A3 N_Y_c_691_n 0.0143942f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_306 N_A3_c_317_n N_Y_c_691_n 5.25617e-19 $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_307 N_A3_M1033_g N_Y_c_693_n 0.0160527f $X=5.775 $Y=2.375 $X2=0 $Y2=0
cc_308 N_A3_c_317_n N_Y_c_693_n 4.61857e-19 $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_309 N_A3_M1002_g N_VPWR_c_779_n 0.00302501f $X=4.485 $Y=2.375 $X2=0 $Y2=0
cc_310 N_A3_M1008_g N_VPWR_c_779_n 0.00302501f $X=4.915 $Y=2.375 $X2=0 $Y2=0
cc_311 N_A3_M1030_g N_VPWR_c_779_n 0.00302501f $X=5.345 $Y=2.375 $X2=0 $Y2=0
cc_312 N_A3_M1033_g N_VPWR_c_779_n 0.00302501f $X=5.775 $Y=2.375 $X2=0 $Y2=0
cc_313 N_A3_M1002_g N_VPWR_c_769_n 0.0048466f $X=4.485 $Y=2.375 $X2=0 $Y2=0
cc_314 N_A3_M1008_g N_VPWR_c_769_n 0.00434671f $X=4.915 $Y=2.375 $X2=0 $Y2=0
cc_315 N_A3_M1030_g N_VPWR_c_769_n 0.00431035f $X=5.345 $Y=2.375 $X2=0 $Y2=0
cc_316 N_A3_M1033_g N_VPWR_c_769_n 0.00435646f $X=5.775 $Y=2.375 $X2=0 $Y2=0
cc_317 A3 N_A_829_349#_M1002_s 0.00227983f $X=5.435 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_318 A3 N_A_829_349#_M1008_s 0.00181948f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_319 N_A3_M1002_g N_A_829_349#_c_897_n 0.0132832f $X=4.485 $Y=2.375 $X2=0
+ $Y2=0
cc_320 N_A3_M1008_g N_A_829_349#_c_897_n 0.0118965f $X=4.915 $Y=2.375 $X2=0
+ $Y2=0
cc_321 N_A3_M1030_g N_A_829_349#_c_899_n 0.0125383f $X=5.345 $Y=2.375 $X2=0
+ $Y2=0
cc_322 N_A3_M1033_g N_A_829_349#_c_899_n 0.0118965f $X=5.775 $Y=2.375 $X2=0
+ $Y2=0
cc_323 N_A3_M1008_g N_A_829_349#_c_903_n 8.24137e-19 $X=4.915 $Y=2.375 $X2=0
+ $Y2=0
cc_324 N_A3_M1033_g N_A_829_349#_c_904_n 8.05012e-19 $X=5.775 $Y=2.375 $X2=0
+ $Y2=0
cc_325 N_A3_M1009_g N_A_30_47#_c_1024_n 0.00183873f $X=4.04 $Y=0.655 $X2=0 $Y2=0
cc_326 N_A3_M1009_g N_A_30_47#_c_1025_n 0.00499461f $X=4.04 $Y=0.655 $X2=0 $Y2=0
cc_327 N_A3_M1009_g N_A_30_47#_c_1036_n 0.0122131f $X=4.04 $Y=0.655 $X2=0 $Y2=0
cc_328 N_A3_M1021_g N_A_30_47#_c_1036_n 0.00963355f $X=4.47 $Y=0.655 $X2=0 $Y2=0
cc_329 N_A3_M1031_g N_A_30_47#_c_1038_n 0.00692874f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_330 N_A3_M1034_g N_A_30_47#_c_1038_n 3.68824e-19 $X=5.47 $Y=0.655 $X2=0 $Y2=0
cc_331 N_A3_M1034_g N_A_30_47#_c_1040_n 0.00314833f $X=5.47 $Y=0.655 $X2=0 $Y2=0
cc_332 N_A3_c_317_n N_A_30_47#_c_1041_n 4.94962e-19 $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_333 N_A3_M1031_g N_A_30_47#_c_1042_n 0.00317387f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_334 N_A3_M1031_g N_A_30_47#_c_1043_n 0.00896496f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_335 N_A3_M1034_g N_A_30_47#_c_1043_n 0.0100268f $X=5.47 $Y=0.655 $X2=0 $Y2=0
cc_336 N_A3_M1009_g N_VGND_c_1167_n 0.00810046f $X=4.04 $Y=0.655 $X2=0 $Y2=0
cc_337 N_A3_M1021_g N_VGND_c_1167_n 0.00697246f $X=4.47 $Y=0.655 $X2=0 $Y2=0
cc_338 N_A3_M1031_g N_VGND_c_1167_n 4.61686e-19 $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_339 N_A3_M1031_g N_VGND_c_1168_n 0.00300641f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_340 N_A3_M1034_g N_VGND_c_1168_n 0.00824166f $X=5.47 $Y=0.655 $X2=0 $Y2=0
cc_341 N_A3_M1009_g N_VGND_c_1172_n 0.00355956f $X=4.04 $Y=0.655 $X2=0 $Y2=0
cc_342 N_A3_M1021_g N_VGND_c_1174_n 0.00355956f $X=4.47 $Y=0.655 $X2=0 $Y2=0
cc_343 N_A3_M1031_g N_VGND_c_1174_n 0.00417814f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_344 N_A3_M1034_g N_VGND_c_1180_n 0.00355956f $X=5.47 $Y=0.655 $X2=0 $Y2=0
cc_345 N_A3_M1009_g N_VGND_c_1183_n 0.00452069f $X=4.04 $Y=0.655 $X2=0 $Y2=0
cc_346 N_A3_M1021_g N_VGND_c_1183_n 0.0044169f $X=4.47 $Y=0.655 $X2=0 $Y2=0
cc_347 N_A3_M1031_g N_VGND_c_1183_n 0.00609256f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_348 N_A3_M1034_g N_VGND_c_1183_n 0.00563228f $X=5.47 $Y=0.655 $X2=0 $Y2=0
cc_349 N_A2_c_411_n N_A1_c_486_n 0.0124275f $X=8.025 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_350 N_A2_c_411_n A1 3.51084e-19 $X=8.025 $Y=1.185 $X2=0 $Y2=0
cc_351 N_A2_c_412_n A1 0.0201927f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_352 N_A2_c_411_n N_A1_c_492_n 0.0224405f $X=8.025 $Y=1.185 $X2=0 $Y2=0
cc_353 N_A2_c_412_n N_A1_c_492_n 3.51084e-19 $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_354 N_A2_c_403_n N_Y_c_613_n 0.0048144f $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_355 N_A2_c_403_n N_Y_c_614_n 5.75192e-19 $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_356 N_A2_c_410_n N_Y_c_614_n 0.00885933f $X=7.57 $Y=1.35 $X2=0 $Y2=0
cc_357 N_A2_c_412_n N_Y_c_614_n 0.0216521f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_358 N_A2_M1005_g N_Y_c_693_n 0.00151f $X=6.205 $Y=2.375 $X2=0 $Y2=0
cc_359 N_A2_M1038_g N_VPWR_c_772_n 0.00143393f $X=7.495 $Y=2.375 $X2=0 $Y2=0
cc_360 N_A2_M1005_g N_VPWR_c_779_n 0.00302501f $X=6.205 $Y=2.375 $X2=0 $Y2=0
cc_361 N_A2_M1016_g N_VPWR_c_779_n 0.00302501f $X=6.635 $Y=2.375 $X2=0 $Y2=0
cc_362 N_A2_M1022_g N_VPWR_c_779_n 0.00302501f $X=7.065 $Y=2.375 $X2=0 $Y2=0
cc_363 N_A2_M1038_g N_VPWR_c_779_n 0.00302501f $X=7.495 $Y=2.375 $X2=0 $Y2=0
cc_364 N_A2_M1005_g N_VPWR_c_769_n 0.00435646f $X=6.205 $Y=2.375 $X2=0 $Y2=0
cc_365 N_A2_M1016_g N_VPWR_c_769_n 0.00434671f $X=6.635 $Y=2.375 $X2=0 $Y2=0
cc_366 N_A2_M1022_g N_VPWR_c_769_n 0.00434671f $X=7.065 $Y=2.375 $X2=0 $Y2=0
cc_367 N_A2_M1038_g N_VPWR_c_769_n 0.0048466f $X=7.495 $Y=2.375 $X2=0 $Y2=0
cc_368 N_A2_M1005_g N_A_829_349#_c_900_n 0.0127027f $X=6.205 $Y=2.375 $X2=0
+ $Y2=0
cc_369 N_A2_M1016_g N_A_829_349#_c_900_n 0.0127216f $X=6.635 $Y=2.375 $X2=0
+ $Y2=0
cc_370 N_A2_M1022_g N_A_829_349#_c_901_n 0.0127216f $X=7.065 $Y=2.375 $X2=0
+ $Y2=0
cc_371 N_A2_M1038_g N_A_829_349#_c_901_n 0.0132832f $X=7.495 $Y=2.375 $X2=0
+ $Y2=0
cc_372 N_A2_M1016_g N_A_1256_349#_c_958_n 0.013787f $X=6.635 $Y=2.375 $X2=0
+ $Y2=0
cc_373 N_A2_M1022_g N_A_1256_349#_c_958_n 0.0138996f $X=7.065 $Y=2.375 $X2=0
+ $Y2=0
cc_374 N_A2_c_410_n N_A_1256_349#_c_958_n 0.0026979f $X=7.57 $Y=1.35 $X2=0 $Y2=0
cc_375 N_A2_c_412_n N_A_1256_349#_c_958_n 0.0433986f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_376 N_A2_M1005_g N_A_1256_349#_c_959_n 9.04234e-19 $X=6.205 $Y=2.375 $X2=0
+ $Y2=0
cc_377 N_A2_c_410_n N_A_1256_349#_c_959_n 0.0027894f $X=7.57 $Y=1.35 $X2=0 $Y2=0
cc_378 N_A2_c_412_n N_A_1256_349#_c_959_n 0.0212944f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_379 N_A2_M1038_g N_A_1256_349#_c_960_n 0.0159867f $X=7.495 $Y=2.375 $X2=0
+ $Y2=0
cc_380 N_A2_c_409_n N_A_1256_349#_c_960_n 0.0157255f $X=7.95 $Y=1.35 $X2=0 $Y2=0
cc_381 N_A2_c_412_n N_A_1256_349#_c_960_n 0.0591566f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_382 N_A2_c_410_n N_A_1256_349#_c_962_n 0.0027894f $X=7.57 $Y=1.35 $X2=0 $Y2=0
cc_383 N_A2_c_412_n N_A_1256_349#_c_962_n 0.0221295f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_384 N_A2_c_403_n N_A_30_47#_c_1040_n 0.0129479f $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_385 N_A2_c_405_n N_A_30_47#_c_1040_n 7.14109e-19 $X=6.795 $Y=1.185 $X2=0
+ $Y2=0
cc_386 N_A2_c_410_n N_A_30_47#_c_1040_n 0.00497272f $X=7.57 $Y=1.35 $X2=0 $Y2=0
cc_387 N_A2_c_412_n N_A_30_47#_c_1040_n 0.0101854f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_388 N_A2_c_403_n N_A_30_47#_c_1049_n 0.00817198f $X=6.365 $Y=1.185 $X2=0
+ $Y2=0
cc_389 N_A2_c_405_n N_A_30_47#_c_1049_n 0.0124062f $X=6.795 $Y=1.185 $X2=0 $Y2=0
cc_390 N_A2_c_410_n N_A_30_47#_c_1049_n 0.00271364f $X=7.57 $Y=1.35 $X2=0 $Y2=0
cc_391 N_A2_c_412_n N_A_30_47#_c_1049_n 0.0351765f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_392 N_A2_c_407_n N_A_30_47#_c_1053_n 0.0144386f $X=7.225 $Y=1.185 $X2=0 $Y2=0
cc_393 N_A2_c_410_n N_A_30_47#_c_1053_n 0.0115594f $X=7.57 $Y=1.35 $X2=0 $Y2=0
cc_394 N_A2_c_411_n N_A_30_47#_c_1053_n 0.0144386f $X=8.025 $Y=1.185 $X2=0 $Y2=0
cc_395 N_A2_c_412_n N_A_30_47#_c_1053_n 0.0650792f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_396 N_A2_c_410_n N_A_30_47#_c_1057_n 0.00280606f $X=7.57 $Y=1.35 $X2=0 $Y2=0
cc_397 N_A2_c_412_n N_A_30_47#_c_1057_n 0.0157444f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_398 N_A2_c_411_n N_A_30_47#_c_1059_n 0.00237027f $X=8.025 $Y=1.185 $X2=0
+ $Y2=0
cc_399 N_A2_c_412_n N_A_30_47#_c_1059_n 0.00647368f $X=8.05 $Y=1.35 $X2=0 $Y2=0
cc_400 N_A2_c_403_n N_VGND_c_1169_n 0.00896863f $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_401 N_A2_c_405_n N_VGND_c_1169_n 0.00681318f $X=6.795 $Y=1.185 $X2=0 $Y2=0
cc_402 N_A2_c_407_n N_VGND_c_1169_n 5.27055e-19 $X=7.225 $Y=1.185 $X2=0 $Y2=0
cc_403 N_A2_c_411_n N_VGND_c_1170_n 5.68058e-19 $X=8.025 $Y=1.185 $X2=0 $Y2=0
cc_404 N_A2_c_411_n N_VGND_c_1176_n 0.00585385f $X=8.025 $Y=1.185 $X2=0 $Y2=0
cc_405 N_A2_c_403_n N_VGND_c_1180_n 0.0038873f $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_406 N_A2_c_405_n N_VGND_c_1181_n 0.00486043f $X=6.795 $Y=1.185 $X2=0 $Y2=0
cc_407 N_A2_c_407_n N_VGND_c_1181_n 0.00585385f $X=7.225 $Y=1.185 $X2=0 $Y2=0
cc_408 N_A2_c_403_n N_VGND_c_1183_n 0.00732762f $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_409 N_A2_c_405_n N_VGND_c_1183_n 0.00824727f $X=6.795 $Y=1.185 $X2=0 $Y2=0
cc_410 N_A2_c_407_n N_VGND_c_1183_n 0.0113749f $X=7.225 $Y=1.185 $X2=0 $Y2=0
cc_411 N_A2_c_411_n N_VGND_c_1183_n 0.0115052f $X=8.025 $Y=1.185 $X2=0 $Y2=0
cc_412 N_A2_c_407_n N_VGND_c_1185_n 0.00317857f $X=7.225 $Y=1.185 $X2=0 $Y2=0
cc_413 N_A2_c_411_n N_VGND_c_1185_n 0.00324785f $X=8.025 $Y=1.185 $X2=0 $Y2=0
cc_414 N_A1_M1000_g N_VPWR_c_772_n 0.0178144f $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_415 N_A1_M1012_g N_VPWR_c_772_n 7.52633e-19 $X=8.93 $Y=2.465 $X2=0 $Y2=0
cc_416 N_A1_M1000_g N_VPWR_c_773_n 7.52633e-19 $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_417 N_A1_M1012_g N_VPWR_c_773_n 0.0160914f $X=8.93 $Y=2.465 $X2=0 $Y2=0
cc_418 N_A1_M1017_g N_VPWR_c_773_n 0.0161833f $X=9.36 $Y=2.465 $X2=0 $Y2=0
cc_419 N_A1_M1026_g N_VPWR_c_773_n 7.68857e-19 $X=9.79 $Y=2.465 $X2=0 $Y2=0
cc_420 N_A1_M1026_g N_VPWR_c_774_n 0.00762775f $X=9.79 $Y=2.465 $X2=0 $Y2=0
cc_421 A1 N_VPWR_c_774_n 0.0150295f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_422 N_A1_c_491_n N_VPWR_c_774_n 0.00629308f $X=10.29 $Y=1.35 $X2=0 $Y2=0
cc_423 N_A1_M1000_g N_VPWR_c_781_n 0.00486043f $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_424 N_A1_M1012_g N_VPWR_c_781_n 0.00486043f $X=8.93 $Y=2.465 $X2=0 $Y2=0
cc_425 N_A1_M1017_g N_VPWR_c_783_n 0.00486043f $X=9.36 $Y=2.465 $X2=0 $Y2=0
cc_426 N_A1_M1026_g N_VPWR_c_783_n 0.00585385f $X=9.79 $Y=2.465 $X2=0 $Y2=0
cc_427 N_A1_M1000_g N_VPWR_c_769_n 0.00824727f $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_428 N_A1_M1012_g N_VPWR_c_769_n 0.00824727f $X=8.93 $Y=2.465 $X2=0 $Y2=0
cc_429 N_A1_M1017_g N_VPWR_c_769_n 0.00824727f $X=9.36 $Y=2.465 $X2=0 $Y2=0
cc_430 N_A1_M1026_g N_VPWR_c_769_n 0.0116533f $X=9.79 $Y=2.465 $X2=0 $Y2=0
cc_431 N_A1_M1000_g N_A_829_349#_c_902_n 0.0017431f $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_432 N_A1_M1000_g N_A_1256_349#_c_960_n 0.0163803f $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_433 A1 N_A_1256_349#_c_960_n 0.0138945f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_434 N_A1_M1012_g N_A_1256_349#_c_961_n 0.0142932f $X=8.93 $Y=2.465 $X2=0
+ $Y2=0
cc_435 N_A1_M1017_g N_A_1256_349#_c_961_n 0.0140113f $X=9.36 $Y=2.465 $X2=0
+ $Y2=0
cc_436 N_A1_M1026_g N_A_1256_349#_c_961_n 0.00522089f $X=9.79 $Y=2.465 $X2=0
+ $Y2=0
cc_437 A1 N_A_1256_349#_c_961_n 0.0667685f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_438 N_A1_c_492_n N_A_1256_349#_c_961_n 0.00878722f $X=9.865 $Y=1.425 $X2=0
+ $Y2=0
cc_439 A1 N_A_1256_349#_c_982_n 0.0150076f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_440 N_A1_c_492_n N_A_1256_349#_c_982_n 0.00524049f $X=9.865 $Y=1.425 $X2=0
+ $Y2=0
cc_441 N_A1_c_486_n N_A_30_47#_c_1061_n 0.0122595f $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_442 N_A1_c_487_n N_A_30_47#_c_1061_n 0.0122595f $X=8.93 $Y=1.185 $X2=0 $Y2=0
cc_443 A1 N_A_30_47#_c_1061_n 0.0390584f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_444 N_A1_c_492_n N_A_30_47#_c_1061_n 0.00249428f $X=9.865 $Y=1.425 $X2=0
+ $Y2=0
cc_445 N_A1_c_488_n N_A_30_47#_c_1005_n 0.0122595f $X=9.36 $Y=1.185 $X2=0 $Y2=0
cc_446 N_A1_c_489_n N_A_30_47#_c_1005_n 0.0122595f $X=9.79 $Y=1.185 $X2=0 $Y2=0
cc_447 A1 N_A_30_47#_c_1005_n 0.0614573f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_448 N_A1_c_491_n N_A_30_47#_c_1005_n 0.00620367f $X=10.29 $Y=1.35 $X2=0 $Y2=0
cc_449 N_A1_c_492_n N_A_30_47#_c_1005_n 0.00249428f $X=9.865 $Y=1.425 $X2=0
+ $Y2=0
cc_450 A1 N_A_30_47#_c_1070_n 0.0144542f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_451 N_A1_c_492_n N_A_30_47#_c_1070_n 0.00258646f $X=9.865 $Y=1.425 $X2=0
+ $Y2=0
cc_452 N_A1_c_486_n N_VGND_c_1170_n 0.0103045f $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_453 N_A1_c_487_n N_VGND_c_1170_n 0.0100888f $X=8.93 $Y=1.185 $X2=0 $Y2=0
cc_454 N_A1_c_488_n N_VGND_c_1170_n 5.75816e-19 $X=9.36 $Y=1.185 $X2=0 $Y2=0
cc_455 N_A1_c_487_n N_VGND_c_1171_n 5.75816e-19 $X=8.93 $Y=1.185 $X2=0 $Y2=0
cc_456 N_A1_c_488_n N_VGND_c_1171_n 0.0100888f $X=9.36 $Y=1.185 $X2=0 $Y2=0
cc_457 N_A1_c_489_n N_VGND_c_1171_n 0.011776f $X=9.79 $Y=1.185 $X2=0 $Y2=0
cc_458 N_A1_c_486_n N_VGND_c_1176_n 0.00486043f $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_459 N_A1_c_487_n N_VGND_c_1178_n 0.00486043f $X=8.93 $Y=1.185 $X2=0 $Y2=0
cc_460 N_A1_c_488_n N_VGND_c_1178_n 0.00486043f $X=9.36 $Y=1.185 $X2=0 $Y2=0
cc_461 N_A1_c_489_n N_VGND_c_1182_n 0.00486043f $X=9.79 $Y=1.185 $X2=0 $Y2=0
cc_462 N_A1_c_486_n N_VGND_c_1183_n 0.00837755f $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_463 N_A1_c_487_n N_VGND_c_1183_n 0.00824727f $X=8.93 $Y=1.185 $X2=0 $Y2=0
cc_464 N_A1_c_488_n N_VGND_c_1183_n 0.00824727f $X=9.36 $Y=1.185 $X2=0 $Y2=0
cc_465 N_A1_c_489_n N_VGND_c_1183_n 0.00936453f $X=9.79 $Y=1.185 $X2=0 $Y2=0
cc_466 N_A_30_367#_c_560_n N_Y_M1006_s 0.00332344f $X=1.04 $Y=2.99 $X2=0 $Y2=0
cc_467 N_A_30_367#_c_562_n N_Y_M1025_s 0.00332344f $X=1.935 $Y=2.99 $X2=0 $Y2=0
cc_468 N_A_30_367#_M1014_d N_Y_c_627_n 0.00334931f $X=0.995 $Y=1.835 $X2=0 $Y2=0
cc_469 N_A_30_367#_c_573_p N_Y_c_627_n 0.0135055f $X=1.135 $Y=2.435 $X2=0 $Y2=0
cc_470 N_A_30_367#_c_560_n N_Y_c_633_n 0.0159805f $X=1.04 $Y=2.99 $X2=0 $Y2=0
cc_471 N_A_30_367#_M1028_d N_Y_c_619_n 0.0090222f $X=1.855 $Y=1.835 $X2=0 $Y2=0
cc_472 N_A_30_367#_M1023_s N_Y_c_619_n 0.00333177f $X=2.75 $Y=1.835 $X2=0 $Y2=0
cc_473 N_A_30_367#_M1037_s N_Y_c_619_n 0.00834034f $X=3.61 $Y=1.835 $X2=0 $Y2=0
cc_474 N_A_30_367#_c_578_p N_Y_c_619_n 0.0144818f $X=2.03 $Y=2.45 $X2=0 $Y2=0
cc_475 N_A_30_367#_c_565_n N_Y_c_619_n 0.0324646f $X=2.795 $Y=2.36 $X2=0 $Y2=0
cc_476 N_A_30_367#_c_567_n N_Y_c_619_n 0.0324646f $X=3.655 $Y=2.36 $X2=0 $Y2=0
cc_477 N_A_30_367#_c_581_p N_Y_c_619_n 0.0135055f $X=2.89 $Y=2.435 $X2=0 $Y2=0
cc_478 N_A_30_367#_c_557_n N_Y_c_619_n 0.020301f $X=3.75 $Y=2.435 $X2=0 $Y2=0
cc_479 N_A_30_367#_c_562_n Y 0.0184743f $X=1.935 $Y=2.99 $X2=0 $Y2=0
cc_480 N_A_30_367#_c_578_p Y 0.0149698f $X=2.03 $Y=2.45 $X2=0 $Y2=0
cc_481 N_A_30_367#_c_564_n Y 0.0213468f $X=2.03 $Y=2.905 $X2=0 $Y2=0
cc_482 N_A_30_367#_c_565_n N_VPWR_M1013_d 0.00344712f $X=2.795 $Y=2.36 $X2=-0.19
+ $Y2=1.655
cc_483 N_A_30_367#_c_567_n N_VPWR_M1029_d 0.00344712f $X=3.655 $Y=2.36 $X2=0
+ $Y2=0
cc_484 N_A_30_367#_c_565_n N_VPWR_c_770_n 0.0171443f $X=2.795 $Y=2.36 $X2=0
+ $Y2=0
cc_485 N_A_30_367#_c_567_n N_VPWR_c_771_n 0.0171443f $X=3.655 $Y=2.36 $X2=0
+ $Y2=0
cc_486 N_A_30_367#_c_555_n N_VPWR_c_775_n 0.0179183f $X=0.24 $Y=2.905 $X2=0
+ $Y2=0
cc_487 N_A_30_367#_c_560_n N_VPWR_c_775_n 0.0361172f $X=1.04 $Y=2.99 $X2=0 $Y2=0
cc_488 N_A_30_367#_c_562_n N_VPWR_c_775_n 0.0509116f $X=1.935 $Y=2.99 $X2=0
+ $Y2=0
cc_489 N_A_30_367#_c_593_p N_VPWR_c_775_n 0.0125234f $X=1.135 $Y=2.99 $X2=0
+ $Y2=0
cc_490 N_A_30_367#_c_581_p N_VPWR_c_777_n 0.0124525f $X=2.89 $Y=2.435 $X2=0
+ $Y2=0
cc_491 N_A_30_367#_c_557_n N_VPWR_c_779_n 0.0178111f $X=3.75 $Y=2.435 $X2=0
+ $Y2=0
cc_492 N_A_30_367#_M1006_d N_VPWR_c_769_n 0.00215161f $X=0.15 $Y=1.835 $X2=0
+ $Y2=0
cc_493 N_A_30_367#_M1014_d N_VPWR_c_769_n 0.00223565f $X=0.995 $Y=1.835 $X2=0
+ $Y2=0
cc_494 N_A_30_367#_M1028_d N_VPWR_c_769_n 0.00404775f $X=1.855 $Y=1.835 $X2=0
+ $Y2=0
cc_495 N_A_30_367#_M1023_s N_VPWR_c_769_n 0.00536646f $X=2.75 $Y=1.835 $X2=0
+ $Y2=0
cc_496 N_A_30_367#_M1037_s N_VPWR_c_769_n 0.00371702f $X=3.61 $Y=1.835 $X2=0
+ $Y2=0
cc_497 N_A_30_367#_c_555_n N_VPWR_c_769_n 0.0101082f $X=0.24 $Y=2.905 $X2=0
+ $Y2=0
cc_498 N_A_30_367#_c_560_n N_VPWR_c_769_n 0.023676f $X=1.04 $Y=2.99 $X2=0 $Y2=0
cc_499 N_A_30_367#_c_562_n N_VPWR_c_769_n 0.0323787f $X=1.935 $Y=2.99 $X2=0
+ $Y2=0
cc_500 N_A_30_367#_c_593_p N_VPWR_c_769_n 0.00738676f $X=1.135 $Y=2.99 $X2=0
+ $Y2=0
cc_501 N_A_30_367#_c_581_p N_VPWR_c_769_n 0.00730901f $X=2.89 $Y=2.435 $X2=0
+ $Y2=0
cc_502 N_A_30_367#_c_557_n N_VPWR_c_769_n 0.0100304f $X=3.75 $Y=2.435 $X2=0
+ $Y2=0
cc_503 N_A_30_367#_c_557_n N_A_829_349#_c_896_n 0.048326f $X=3.75 $Y=2.435 $X2=0
+ $Y2=0
cc_504 N_A_30_367#_c_557_n N_A_829_349#_c_898_n 0.0136671f $X=3.75 $Y=2.435
+ $X2=0 $Y2=0
cc_505 N_Y_c_619_n N_VPWR_M1013_d 0.00333608f $X=4.57 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_506 N_Y_c_619_n N_VPWR_M1029_d 0.00333608f $X=4.57 $Y=2.015 $X2=0 $Y2=0
cc_507 N_Y_M1006_s N_VPWR_c_769_n 0.00225186f $X=0.565 $Y=1.835 $X2=0 $Y2=0
cc_508 N_Y_M1025_s N_VPWR_c_769_n 0.00225186f $X=1.425 $Y=1.835 $X2=0 $Y2=0
cc_509 N_Y_c_619_n N_A_829_349#_M1002_s 0.00486436f $X=4.57 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_510 N_Y_c_677_n N_A_829_349#_M1008_s 0.00336353f $X=5.415 $Y=2.015 $X2=0
+ $Y2=0
cc_511 N_Y_c_614_n N_A_829_349#_M1033_s 0.00215545f $X=5.92 $Y=1.93 $X2=0 $Y2=0
cc_512 N_Y_c_693_n N_A_829_349#_M1033_s 0.00309954f $X=5.92 $Y=2.015 $X2=0 $Y2=0
cc_513 N_Y_c_619_n N_A_829_349#_c_896_n 0.0202165f $X=4.57 $Y=2.015 $X2=0 $Y2=0
cc_514 N_Y_M1002_d N_A_829_349#_c_897_n 0.00176461f $X=4.56 $Y=1.745 $X2=0 $Y2=0
cc_515 N_Y_c_691_n N_A_829_349#_c_897_n 0.0126348f $X=4.7 $Y=2.095 $X2=0 $Y2=0
cc_516 N_Y_c_677_n N_A_829_349#_c_928_n 0.0135055f $X=5.415 $Y=2.015 $X2=0 $Y2=0
cc_517 N_Y_M1030_d N_A_829_349#_c_899_n 0.00176461f $X=5.42 $Y=1.745 $X2=0 $Y2=0
cc_518 N_Y_c_681_n N_A_829_349#_c_899_n 0.0127809f $X=5.547 $Y=2.1 $X2=0 $Y2=0
cc_519 N_Y_c_693_n N_A_829_349#_c_931_n 0.00793666f $X=5.92 $Y=2.015 $X2=0 $Y2=0
cc_520 N_Y_c_614_n N_A_1256_349#_c_959_n 0.00690884f $X=5.92 $Y=1.93 $X2=0 $Y2=0
cc_521 N_Y_c_609_n N_A_30_47#_M1018_s 0.00176461f $X=1.47 $Y=1.09 $X2=0 $Y2=0
cc_522 N_Y_c_611_n N_A_30_47#_M1027_s 0.00176461f $X=2.33 $Y=1.09 $X2=0 $Y2=0
cc_523 N_Y_c_612_n N_A_30_47#_M1015_s 0.00176461f $X=3.19 $Y=1.09 $X2=0 $Y2=0
cc_524 N_Y_c_613_n N_A_30_47#_M1039_s 0.00306584f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_525 N_Y_c_613_n N_A_30_47#_M1021_s 0.00250873f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_526 N_Y_c_613_n N_A_30_47#_M1034_s 0.00652081f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_527 N_Y_c_610_n N_A_30_47#_c_1003_n 0.00166417f $X=0.8 $Y=1.09 $X2=0 $Y2=0
cc_528 N_Y_M1003_d N_A_30_47#_c_1010_n 0.00332344f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_529 N_Y_c_740_p N_A_30_47#_c_1010_n 0.0124813f $X=0.705 $Y=0.76 $X2=0 $Y2=0
cc_530 N_Y_c_609_n N_A_30_47#_c_1010_n 0.00306745f $X=1.47 $Y=1.09 $X2=0 $Y2=0
cc_531 N_Y_M1020_d N_A_30_47#_c_1012_n 0.00332344f $X=1.425 $Y=0.235 $X2=0 $Y2=0
cc_532 N_Y_c_609_n N_A_30_47#_c_1012_n 0.00306745f $X=1.47 $Y=1.09 $X2=0 $Y2=0
cc_533 N_Y_c_744_p N_A_30_47#_c_1012_n 0.0124813f $X=1.565 $Y=0.76 $X2=0 $Y2=0
cc_534 N_Y_c_611_n N_A_30_47#_c_1012_n 0.00306745f $X=2.33 $Y=1.09 $X2=0 $Y2=0
cc_535 N_Y_M1001_d N_A_30_47#_c_1020_n 0.00332344f $X=2.285 $Y=0.235 $X2=0 $Y2=0
cc_536 N_Y_c_611_n N_A_30_47#_c_1020_n 0.00306745f $X=2.33 $Y=1.09 $X2=0 $Y2=0
cc_537 N_Y_c_748_p N_A_30_47#_c_1020_n 0.0124813f $X=2.425 $Y=0.76 $X2=0 $Y2=0
cc_538 N_Y_c_612_n N_A_30_47#_c_1020_n 0.00306745f $X=3.19 $Y=1.09 $X2=0 $Y2=0
cc_539 N_Y_M1024_d N_A_30_47#_c_1022_n 0.00333487f $X=3.145 $Y=0.235 $X2=0 $Y2=0
cc_540 N_Y_c_612_n N_A_30_47#_c_1022_n 0.00319377f $X=3.19 $Y=1.09 $X2=0 $Y2=0
cc_541 N_Y_c_752_p N_A_30_47#_c_1022_n 0.0126023f $X=3.285 $Y=0.78 $X2=0 $Y2=0
cc_542 N_Y_c_613_n N_A_30_47#_c_1022_n 0.00324593f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_543 N_Y_c_613_n N_A_30_47#_c_1036_n 0.0343548f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_544 N_Y_c_613_n N_A_30_47#_c_1027_n 0.0217249f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_545 N_Y_c_613_n N_A_30_47#_c_1040_n 0.00405725f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_546 N_Y_c_613_n N_A_30_47#_c_1041_n 0.0150152f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_547 N_Y_c_609_n N_A_30_47#_c_1014_n 0.0168576f $X=1.47 $Y=1.09 $X2=0 $Y2=0
cc_548 N_Y_c_611_n N_A_30_47#_c_1018_n 0.0168576f $X=2.33 $Y=1.09 $X2=0 $Y2=0
cc_549 N_Y_c_612_n N_A_30_47#_c_1030_n 0.0168576f $X=3.19 $Y=1.09 $X2=0 $Y2=0
cc_550 N_Y_c_613_n N_A_30_47#_c_1042_n 0.0208046f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_551 N_Y_c_613_n N_A_30_47#_c_1043_n 0.0542761f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_552 N_Y_c_613_n N_VGND_M1009_d 0.00176891f $X=5.835 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_553 N_Y_c_613_n N_VGND_M1031_d 0.00251484f $X=5.835 $Y=1.08 $X2=0 $Y2=0
cc_554 N_Y_M1003_d N_VGND_c_1183_n 0.00225186f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_555 N_Y_M1020_d N_VGND_c_1183_n 0.00225186f $X=1.425 $Y=0.235 $X2=0 $Y2=0
cc_556 N_Y_M1001_d N_VGND_c_1183_n 0.00225186f $X=2.285 $Y=0.235 $X2=0 $Y2=0
cc_557 N_Y_M1024_d N_VGND_c_1183_n 0.00225186f $X=3.145 $Y=0.235 $X2=0 $Y2=0
cc_558 N_VPWR_c_779_n N_A_829_349#_c_897_n 0.0386886f $X=8.12 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_769_n N_A_829_349#_c_897_n 0.02175f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_560 N_VPWR_c_779_n N_A_829_349#_c_898_n 0.0193554f $X=8.12 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_769_n N_A_829_349#_c_898_n 0.010497f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_779_n N_A_829_349#_c_899_n 0.0380182f $X=8.12 $Y=3.33 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_769_n N_A_829_349#_c_899_n 0.0213705f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_779_n N_A_829_349#_c_900_n 0.0373973f $X=8.12 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_769_n N_A_829_349#_c_900_n 0.0209975f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_772_n N_A_829_349#_c_901_n 0.0116404f $X=8.285 $Y=2.09 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_779_n N_A_829_349#_c_901_n 0.0591891f $X=8.12 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_769_n N_A_829_349#_c_901_n 0.0328424f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_772_n N_A_829_349#_c_902_n 0.0575668f $X=8.285 $Y=2.09 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_779_n N_A_829_349#_c_903_n 0.0182801f $X=8.12 $Y=3.33 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_769_n N_A_829_349#_c_903_n 0.00991381f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_572 N_VPWR_c_779_n N_A_829_349#_c_904_n 0.0193554f $X=8.12 $Y=3.33 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_769_n N_A_829_349#_c_904_n 0.010497f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_779_n N_A_829_349#_c_905_n 0.0186386f $X=8.12 $Y=3.33 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_769_n N_A_829_349#_c_905_n 0.0101082f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_769_n N_A_1256_349#_M1000_s 0.00536646f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_769_n N_A_1256_349#_M1017_s 0.00397496f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_772_n N_A_1256_349#_c_960_n 0.0244345f $X=8.285 $Y=2.09 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_781_n N_A_1256_349#_c_988_n 0.0124525f $X=8.98 $Y=3.33 $X2=0
+ $Y2=0
cc_580 N_VPWR_c_769_n N_A_1256_349#_c_988_n 0.00730901f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_581 N_VPWR_c_773_n N_A_1256_349#_c_961_n 0.0216087f $X=9.145 $Y=2.09 $X2=0
+ $Y2=0
cc_582 N_VPWR_c_774_n N_A_1256_349#_c_961_n 0.00166417f $X=10.005 $Y=1.98 $X2=0
+ $Y2=0
cc_583 N_VPWR_c_783_n N_A_1256_349#_c_992_n 0.0138717f $X=9.88 $Y=3.33 $X2=0
+ $Y2=0
cc_584 N_VPWR_c_769_n N_A_1256_349#_c_992_n 0.00886411f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_585 N_A_829_349#_c_900_n N_A_1256_349#_M1005_s 0.00176461f $X=6.715 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_586 N_A_829_349#_c_901_n N_A_1256_349#_M1022_s 0.00176461f $X=7.58 $Y=2.99
+ $X2=0 $Y2=0
cc_587 N_A_829_349#_c_900_n N_A_1256_349#_c_996_n 0.0126348f $X=6.715 $Y=2.99
+ $X2=0 $Y2=0
cc_588 N_A_829_349#_M1016_d N_A_1256_349#_c_958_n 0.00176461f $X=6.71 $Y=1.745
+ $X2=0 $Y2=0
cc_589 N_A_829_349#_c_954_p N_A_1256_349#_c_958_n 0.0135055f $X=6.85 $Y=2.17
+ $X2=0 $Y2=0
cc_590 N_A_829_349#_c_901_n N_A_1256_349#_c_999_n 0.0126348f $X=7.58 $Y=2.99
+ $X2=0 $Y2=0
cc_591 N_A_829_349#_M1038_d N_A_1256_349#_c_960_n 0.00262981f $X=7.57 $Y=1.745
+ $X2=0 $Y2=0
cc_592 N_A_829_349#_c_902_n N_A_1256_349#_c_960_n 0.0202165f $X=7.71 $Y=2.17
+ $X2=0 $Y2=0
cc_593 N_A_1256_349#_c_960_n N_A_30_47#_c_1059_n 0.00509225f $X=8.62 $Y=1.75
+ $X2=0 $Y2=0
cc_594 N_A_30_47#_c_1036_n N_VGND_M1009_d 0.00333053f $X=4.59 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_595 N_A_30_47#_c_1043_n N_VGND_M1031_d 0.00469582f $X=5.59 $Y=0.54 $X2=0
+ $Y2=0
cc_596 N_A_30_47#_c_1049_n N_VGND_M1004_d 0.00417571f $X=6.915 $Y=0.955 $X2=0
+ $Y2=0
cc_597 N_A_30_47#_c_1053_n N_VGND_M1019_d 0.0128715f $X=8.11 $Y=0.955 $X2=0
+ $Y2=0
cc_598 N_A_30_47#_c_1061_n N_VGND_M1007_s 0.00329816f $X=9.05 $Y=0.955 $X2=0
+ $Y2=0
cc_599 N_A_30_47#_c_1005_n N_VGND_M1035_s 0.00329816f $X=9.91 $Y=0.955 $X2=0
+ $Y2=0
cc_600 N_A_30_47#_c_1024_n N_VGND_c_1167_n 0.0133291f $X=3.715 $Y=0.445 $X2=0
+ $Y2=0
cc_601 N_A_30_47#_c_1025_n N_VGND_c_1167_n 0.00260495f $X=3.715 $Y=0.655 $X2=0
+ $Y2=0
cc_602 N_A_30_47#_c_1036_n N_VGND_c_1167_n 0.016098f $X=4.59 $Y=0.74 $X2=0 $Y2=0
cc_603 N_A_30_47#_c_1043_n N_VGND_c_1168_n 0.0197854f $X=5.59 $Y=0.54 $X2=0
+ $Y2=0
cc_604 N_A_30_47#_c_1049_n N_VGND_c_1169_n 0.00928814f $X=6.915 $Y=0.955 $X2=0
+ $Y2=0
cc_605 N_A_30_47#_c_1061_n N_VGND_c_1170_n 0.0170777f $X=9.05 $Y=0.955 $X2=0
+ $Y2=0
cc_606 N_A_30_47#_c_1005_n N_VGND_c_1171_n 0.0170777f $X=9.91 $Y=0.955 $X2=0
+ $Y2=0
cc_607 N_A_30_47#_c_1010_n N_VGND_c_1172_n 0.0319341f $X=0.97 $Y=0.34 $X2=0
+ $Y2=0
cc_608 N_A_30_47#_c_1004_n N_VGND_c_1172_n 0.0189827f $X=0.4 $Y=0.34 $X2=0 $Y2=0
cc_609 N_A_30_47#_c_1012_n N_VGND_c_1172_n 0.0298674f $X=1.83 $Y=0.34 $X2=0
+ $Y2=0
cc_610 N_A_30_47#_c_1020_n N_VGND_c_1172_n 0.0298674f $X=2.69 $Y=0.34 $X2=0
+ $Y2=0
cc_611 N_A_30_47#_c_1022_n N_VGND_c_1172_n 0.0300582f $X=3.55 $Y=0.35 $X2=0
+ $Y2=0
cc_612 N_A_30_47#_c_1024_n N_VGND_c_1172_n 0.0208876f $X=3.715 $Y=0.445 $X2=0
+ $Y2=0
cc_613 N_A_30_47#_c_1036_n N_VGND_c_1172_n 0.00293018f $X=4.59 $Y=0.74 $X2=0
+ $Y2=0
cc_614 N_A_30_47#_c_1014_n N_VGND_c_1172_n 0.0188892f $X=1.135 $Y=0.38 $X2=0
+ $Y2=0
cc_615 N_A_30_47#_c_1018_n N_VGND_c_1172_n 0.0188892f $X=1.995 $Y=0.38 $X2=0
+ $Y2=0
cc_616 N_A_30_47#_c_1030_n N_VGND_c_1172_n 0.0188892f $X=2.855 $Y=0.38 $X2=0
+ $Y2=0
cc_617 N_A_30_47#_c_1036_n N_VGND_c_1174_n 0.00235176f $X=4.59 $Y=0.74 $X2=0
+ $Y2=0
cc_618 N_A_30_47#_c_1038_n N_VGND_c_1174_n 0.0203777f $X=4.755 $Y=0.375 $X2=0
+ $Y2=0
cc_619 N_A_30_47#_c_1043_n N_VGND_c_1174_n 0.00235176f $X=5.59 $Y=0.54 $X2=0
+ $Y2=0
cc_620 N_A_30_47#_c_1130_p N_VGND_c_1176_n 0.0168584f $X=8.24 $Y=0.42 $X2=0
+ $Y2=0
cc_621 N_A_30_47#_c_1131_p N_VGND_c_1178_n 0.0124525f $X=9.145 $Y=0.42 $X2=0
+ $Y2=0
cc_622 N_A_30_47#_c_1040_n N_VGND_c_1180_n 0.00559624f $X=6.175 $Y=0.54 $X2=0
+ $Y2=0
cc_623 N_A_30_47#_c_1041_n N_VGND_c_1180_n 0.0398659f $X=5.875 $Y=0.54 $X2=0
+ $Y2=0
cc_624 N_A_30_47#_c_1043_n N_VGND_c_1180_n 0.00235176f $X=5.59 $Y=0.54 $X2=0
+ $Y2=0
cc_625 N_A_30_47#_c_1135_p N_VGND_c_1181_n 0.0136943f $X=7.01 $Y=0.42 $X2=0
+ $Y2=0
cc_626 N_A_30_47#_c_1006_n N_VGND_c_1182_n 0.0178111f $X=10.005 $Y=0.42 $X2=0
+ $Y2=0
cc_627 N_A_30_47#_M1003_s N_VGND_c_1183_n 0.00215159f $X=0.15 $Y=0.235 $X2=0
+ $Y2=0
cc_628 N_A_30_47#_M1018_s N_VGND_c_1183_n 0.00223559f $X=0.995 $Y=0.235 $X2=0
+ $Y2=0
cc_629 N_A_30_47#_M1027_s N_VGND_c_1183_n 0.00223559f $X=1.855 $Y=0.235 $X2=0
+ $Y2=0
cc_630 N_A_30_47#_M1015_s N_VGND_c_1183_n 0.00223559f $X=2.715 $Y=0.235 $X2=0
+ $Y2=0
cc_631 N_A_30_47#_M1039_s N_VGND_c_1183_n 0.00346783f $X=3.575 $Y=0.235 $X2=0
+ $Y2=0
cc_632 N_A_30_47#_M1021_s N_VGND_c_1183_n 0.00297296f $X=4.545 $Y=0.235 $X2=0
+ $Y2=0
cc_633 N_A_30_47#_M1034_s N_VGND_c_1183_n 0.00649977f $X=5.545 $Y=0.235 $X2=0
+ $Y2=0
cc_634 N_A_30_47#_M1010_s N_VGND_c_1183_n 0.0041489f $X=6.87 $Y=0.235 $X2=0
+ $Y2=0
cc_635 N_A_30_47#_M1032_s N_VGND_c_1183_n 0.00451078f $X=8.1 $Y=0.235 $X2=0
+ $Y2=0
cc_636 N_A_30_47#_M1011_d N_VGND_c_1183_n 0.00536646f $X=9.005 $Y=0.235 $X2=0
+ $Y2=0
cc_637 N_A_30_47#_M1036_d N_VGND_c_1183_n 0.00371702f $X=9.865 $Y=0.235 $X2=0
+ $Y2=0
cc_638 N_A_30_47#_c_1010_n N_VGND_c_1183_n 0.0201012f $X=0.97 $Y=0.34 $X2=0
+ $Y2=0
cc_639 N_A_30_47#_c_1004_n N_VGND_c_1183_n 0.0112745f $X=0.4 $Y=0.34 $X2=0 $Y2=0
cc_640 N_A_30_47#_c_1012_n N_VGND_c_1183_n 0.0187823f $X=1.83 $Y=0.34 $X2=0
+ $Y2=0
cc_641 N_A_30_47#_c_1020_n N_VGND_c_1183_n 0.0187823f $X=2.69 $Y=0.34 $X2=0
+ $Y2=0
cc_642 N_A_30_47#_c_1022_n N_VGND_c_1183_n 0.0188286f $X=3.55 $Y=0.35 $X2=0
+ $Y2=0
cc_643 N_A_30_47#_c_1024_n N_VGND_c_1183_n 0.0125837f $X=3.715 $Y=0.445 $X2=0
+ $Y2=0
cc_644 N_A_30_47#_c_1036_n N_VGND_c_1183_n 0.0108837f $X=4.59 $Y=0.74 $X2=0
+ $Y2=0
cc_645 N_A_30_47#_c_1038_n N_VGND_c_1183_n 0.0125108f $X=4.755 $Y=0.375 $X2=0
+ $Y2=0
cc_646 N_A_30_47#_c_1040_n N_VGND_c_1183_n 0.00526241f $X=6.175 $Y=0.54 $X2=0
+ $Y2=0
cc_647 N_A_30_47#_c_1041_n N_VGND_c_1183_n 0.022616f $X=5.875 $Y=0.54 $X2=0
+ $Y2=0
cc_648 N_A_30_47#_c_1135_p N_VGND_c_1183_n 0.00866972f $X=7.01 $Y=0.42 $X2=0
+ $Y2=0
cc_649 N_A_30_47#_c_1130_p N_VGND_c_1183_n 0.0104192f $X=8.24 $Y=0.42 $X2=0
+ $Y2=0
cc_650 N_A_30_47#_c_1131_p N_VGND_c_1183_n 0.00730901f $X=9.145 $Y=0.42 $X2=0
+ $Y2=0
cc_651 N_A_30_47#_c_1006_n N_VGND_c_1183_n 0.0100304f $X=10.005 $Y=0.42 $X2=0
+ $Y2=0
cc_652 N_A_30_47#_c_1014_n N_VGND_c_1183_n 0.0124024f $X=1.135 $Y=0.38 $X2=0
+ $Y2=0
cc_653 N_A_30_47#_c_1018_n N_VGND_c_1183_n 0.0124024f $X=1.995 $Y=0.38 $X2=0
+ $Y2=0
cc_654 N_A_30_47#_c_1030_n N_VGND_c_1183_n 0.0124024f $X=2.855 $Y=0.38 $X2=0
+ $Y2=0
cc_655 N_A_30_47#_c_1043_n N_VGND_c_1183_n 0.00973063f $X=5.59 $Y=0.54 $X2=0
+ $Y2=0
cc_656 N_A_30_47#_c_1053_n N_VGND_c_1185_n 0.0436082f $X=8.11 $Y=0.955 $X2=0
+ $Y2=0
