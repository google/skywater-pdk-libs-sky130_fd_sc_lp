* File: sky130_fd_sc_lp__and3_1.pxi.spice
* Created: Fri Aug 28 10:05:51 2020
* 
x_PM_SKY130_FD_SC_LP__AND3_1%A N_A_M1005_g N_A_M1002_g A N_A_c_56_n
+ PM_SKY130_FD_SC_LP__AND3_1%A
x_PM_SKY130_FD_SC_LP__AND3_1%B N_B_M1006_g N_B_M1007_g B N_B_c_85_n
+ PM_SKY130_FD_SC_LP__AND3_1%B
x_PM_SKY130_FD_SC_LP__AND3_1%C N_C_M1004_g N_C_M1000_g C C C C C N_C_c_116_n
+ N_C_c_117_n C PM_SKY130_FD_SC_LP__AND3_1%C
x_PM_SKY130_FD_SC_LP__AND3_1%A_61_367# N_A_61_367#_M1002_s N_A_61_367#_M1005_s
+ N_A_61_367#_M1007_d N_A_61_367#_M1001_g N_A_61_367#_M1003_g
+ N_A_61_367#_c_165_n N_A_61_367#_c_174_n N_A_61_367#_c_166_n
+ N_A_61_367#_c_167_n N_A_61_367#_c_176_n N_A_61_367#_c_168_n
+ N_A_61_367#_c_169_n N_A_61_367#_c_170_n N_A_61_367#_c_171_n
+ N_A_61_367#_c_172_n PM_SKY130_FD_SC_LP__AND3_1%A_61_367#
x_PM_SKY130_FD_SC_LP__AND3_1%VPWR N_VPWR_M1005_d N_VPWR_M1000_d N_VPWR_c_247_n
+ N_VPWR_c_248_n N_VPWR_c_249_n N_VPWR_c_250_n VPWR N_VPWR_c_251_n
+ N_VPWR_c_252_n N_VPWR_c_246_n N_VPWR_c_254_n PM_SKY130_FD_SC_LP__AND3_1%VPWR
x_PM_SKY130_FD_SC_LP__AND3_1%X N_X_M1001_d N_X_M1003_d X X X X X X X N_X_c_275_n
+ X PM_SKY130_FD_SC_LP__AND3_1%X
x_PM_SKY130_FD_SC_LP__AND3_1%VGND N_VGND_M1004_d N_VGND_c_293_n N_VGND_c_294_n
+ N_VGND_c_295_n VGND N_VGND_c_296_n N_VGND_c_297_n
+ PM_SKY130_FD_SC_LP__AND3_1%VGND
cc_1 VNB N_A_M1005_g 0.0141755f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.045
cc_2 VNB N_A_M1002_g 0.038899f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.475
cc_3 VNB A 0.00328655f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_c_56_n 0.0318699f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.27
cc_5 VNB N_B_M1006_g 0.0330128f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.045
cc_6 VNB N_B_M1007_g 0.012058f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.475
cc_7 VNB B 0.00451813f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_B_c_85_n 0.0275276f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.27
cc_9 VNB N_C_M1004_g 0.0418281f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.045
cc_10 VNB N_C_M1000_g 0.00607467f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.475
cc_11 VNB C 8.35218e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C_c_116_n 0.0336645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C_c_117_n 0.00460633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_61_367#_M1001_g 0.0251019f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.27
cc_15 VNB N_A_61_367#_M1003_g 0.00126934f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.27
cc_16 VNB N_A_61_367#_c_165_n 0.0319038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_61_367#_c_166_n 0.00630523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_61_367#_c_167_n 0.0227102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_61_367#_c_168_n 0.0015531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_61_367#_c_169_n 0.033649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_61_367#_c_170_n 0.00508882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_61_367#_c_171_n 0.00343242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_61_367#_c_172_n 0.0389438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_246_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB X 0.0287167f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_26 VNB N_X_c_275_n 0.0339723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0156323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_293_n 0.00661825f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.475
cc_29 VNB N_VGND_c_294_n 0.0535174f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_30 VNB N_VGND_c_295_n 0.00632158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_296_n 0.0232341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_297_n 0.186847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A_M1005_g 0.0294376f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.045
cc_34 VPB N_B_M1007_g 0.0246705f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=0.475
cc_35 VPB N_C_M1000_g 0.0227263f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=0.475
cc_36 VPB C 0.00297052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB C 0.0159178f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.27
cc_38 VPB C 0.00307308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_61_367#_M1003_g 0.0269763f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.27
cc_40 VPB N_A_61_367#_c_174_n 0.0263498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_61_367#_c_166_n 0.00476118f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_61_367#_c_176_n 9.68691e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_61_367#_c_170_n 0.0059747f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_247_n 0.0556395f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_45 VPB N_VPWR_c_248_n 0.0208376f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.27
cc_46 VPB N_VPWR_c_249_n 0.0255325f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.27
cc_47 VPB N_VPWR_c_250_n 0.00535984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_251_n 0.0276675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_252_n 0.0159542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_246_n 0.100555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_254_n 0.00612933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB X 0.0595412f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_53 N_A_M1002_g N_B_M1006_g 0.0358509f $X=0.67 $Y=0.475 $X2=0 $Y2=0
cc_54 N_A_M1005_g N_B_M1007_g 0.0244879f $X=0.645 $Y=2.045 $X2=0 $Y2=0
cc_55 A B 0.0263531f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A_c_56_n B 3.62375e-19 $X=0.58 $Y=1.27 $X2=0 $Y2=0
cc_57 A N_B_c_85_n 0.00110775f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_58 N_A_c_56_n N_B_c_85_n 0.0358509f $X=0.58 $Y=1.27 $X2=0 $Y2=0
cc_59 N_A_M1005_g N_A_61_367#_c_165_n 0.00373495f $X=0.645 $Y=2.045 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_A_61_367#_c_165_n 0.00363706f $X=0.67 $Y=0.475 $X2=0 $Y2=0
cc_61 A N_A_61_367#_c_165_n 0.0247707f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A_c_56_n N_A_61_367#_c_165_n 0.00806477f $X=0.58 $Y=1.27 $X2=0 $Y2=0
cc_63 N_A_M1005_g N_A_61_367#_c_174_n 0.0021737f $X=0.645 $Y=2.045 $X2=0 $Y2=0
cc_64 N_A_M1005_g N_A_61_367#_c_166_n 0.016526f $X=0.645 $Y=2.045 $X2=0 $Y2=0
cc_65 A N_A_61_367#_c_166_n 0.0184789f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A_c_56_n N_A_61_367#_c_166_n 7.68921e-19 $X=0.58 $Y=1.27 $X2=0 $Y2=0
cc_67 N_A_M1002_g N_A_61_367#_c_167_n 0.0086436f $X=0.67 $Y=0.475 $X2=0 $Y2=0
cc_68 A N_A_61_367#_c_167_n 0.0144766f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_M1002_g N_A_61_367#_c_169_n 0.0156998f $X=0.67 $Y=0.475 $X2=0 $Y2=0
cc_70 A N_A_61_367#_c_169_n 0.0111149f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_c_56_n N_A_61_367#_c_169_n 0.00473998f $X=0.58 $Y=1.27 $X2=0 $Y2=0
cc_72 A N_A_61_367#_c_170_n 0.0066825f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A_c_56_n N_A_61_367#_c_170_n 0.00393882f $X=0.58 $Y=1.27 $X2=0 $Y2=0
cc_74 N_A_M1005_g N_VPWR_c_247_n 0.00360463f $X=0.645 $Y=2.045 $X2=0 $Y2=0
cc_75 N_A_M1002_g N_VGND_c_294_n 0.00522167f $X=0.67 $Y=0.475 $X2=0 $Y2=0
cc_76 N_A_M1002_g N_VGND_c_297_n 0.00669905f $X=0.67 $Y=0.475 $X2=0 $Y2=0
cc_77 N_B_M1006_g N_C_M1004_g 0.0330787f $X=1.06 $Y=0.475 $X2=0 $Y2=0
cc_78 B N_C_M1004_g 0.00105098f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B_c_85_n N_C_M1004_g 0.0213609f $X=1.15 $Y=1.27 $X2=0 $Y2=0
cc_80 N_B_M1007_g C 0.00111381f $X=1.095 $Y=2.045 $X2=0 $Y2=0
cc_81 N_B_M1007_g N_C_c_116_n 0.017264f $X=1.095 $Y=2.045 $X2=0 $Y2=0
cc_82 N_B_M1007_g N_C_c_117_n 7.31916e-19 $X=1.095 $Y=2.045 $X2=0 $Y2=0
cc_83 B N_C_c_117_n 0.027262f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_84 N_B_c_85_n N_C_c_117_n 9.73062e-19 $X=1.15 $Y=1.27 $X2=0 $Y2=0
cc_85 N_B_M1007_g C 2.25551e-19 $X=1.095 $Y=2.045 $X2=0 $Y2=0
cc_86 N_B_M1007_g N_A_61_367#_c_166_n 0.0147748f $X=1.095 $Y=2.045 $X2=0 $Y2=0
cc_87 B N_A_61_367#_c_166_n 0.0274819f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B_c_85_n N_A_61_367#_c_166_n 0.00426987f $X=1.15 $Y=1.27 $X2=0 $Y2=0
cc_89 N_B_M1006_g N_A_61_367#_c_167_n 0.0119214f $X=1.06 $Y=0.475 $X2=0 $Y2=0
cc_90 B N_A_61_367#_c_167_n 0.0262222f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B_c_85_n N_A_61_367#_c_167_n 0.0041736f $X=1.15 $Y=1.27 $X2=0 $Y2=0
cc_92 N_B_M1007_g N_A_61_367#_c_176_n 9.86245e-19 $X=1.095 $Y=2.045 $X2=0 $Y2=0
cc_93 N_B_M1006_g N_A_61_367#_c_169_n 0.00232236f $X=1.06 $Y=0.475 $X2=0 $Y2=0
cc_94 N_B_M1007_g N_VPWR_c_247_n 0.00187795f $X=1.095 $Y=2.045 $X2=0 $Y2=0
cc_95 N_B_M1006_g N_VGND_c_294_n 0.00555245f $X=1.06 $Y=0.475 $X2=0 $Y2=0
cc_96 N_B_M1006_g N_VGND_c_297_n 0.00617788f $X=1.06 $Y=0.475 $X2=0 $Y2=0
cc_97 N_C_M1004_g N_A_61_367#_M1001_g 0.0243514f $X=1.6 $Y=0.475 $X2=0 $Y2=0
cc_98 N_C_c_116_n N_A_61_367#_M1001_g 0.00407639f $X=1.69 $Y=1.38 $X2=0 $Y2=0
cc_99 N_C_c_117_n N_A_61_367#_M1001_g 3.55941e-19 $X=1.685 $Y=1.52 $X2=0 $Y2=0
cc_100 N_C_M1000_g N_A_61_367#_M1003_g 0.00821703f $X=1.6 $Y=2.045 $X2=0 $Y2=0
cc_101 C N_A_61_367#_M1003_g 0.00463219f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_102 N_C_M1000_g N_A_61_367#_c_166_n 0.00140141f $X=1.6 $Y=2.045 $X2=0 $Y2=0
cc_103 C N_A_61_367#_c_166_n 0.013766f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_104 N_C_M1004_g N_A_61_367#_c_167_n 0.0129595f $X=1.6 $Y=0.475 $X2=0 $Y2=0
cc_105 N_C_c_116_n N_A_61_367#_c_167_n 0.00320359f $X=1.69 $Y=1.38 $X2=0 $Y2=0
cc_106 N_C_c_117_n N_A_61_367#_c_167_n 0.0208086f $X=1.685 $Y=1.52 $X2=0 $Y2=0
cc_107 N_C_M1000_g N_A_61_367#_c_176_n 0.00154238f $X=1.6 $Y=2.045 $X2=0 $Y2=0
cc_108 C N_A_61_367#_c_176_n 0.0315517f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_109 N_C_M1004_g N_A_61_367#_c_168_n 0.00368307f $X=1.6 $Y=0.475 $X2=0 $Y2=0
cc_110 N_C_c_116_n N_A_61_367#_c_168_n 6.36029e-19 $X=1.69 $Y=1.38 $X2=0 $Y2=0
cc_111 N_C_c_117_n N_A_61_367#_c_168_n 0.0153627f $X=1.685 $Y=1.52 $X2=0 $Y2=0
cc_112 N_C_M1000_g N_A_61_367#_c_171_n 2.73006e-19 $X=1.6 $Y=2.045 $X2=0 $Y2=0
cc_113 C N_A_61_367#_c_171_n 0.00908958f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_114 N_C_c_116_n N_A_61_367#_c_171_n 0.00160409f $X=1.69 $Y=1.38 $X2=0 $Y2=0
cc_115 N_C_c_117_n N_A_61_367#_c_171_n 0.0169277f $X=1.685 $Y=1.52 $X2=0 $Y2=0
cc_116 N_C_M1000_g N_A_61_367#_c_172_n 0.00259092f $X=1.6 $Y=2.045 $X2=0 $Y2=0
cc_117 C N_A_61_367#_c_172_n 2.51352e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_118 N_C_c_116_n N_A_61_367#_c_172_n 0.0148798f $X=1.69 $Y=1.38 $X2=0 $Y2=0
cc_119 C N_VPWR_M1000_d 0.00402737f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_120 C N_VPWR_c_247_n 0.00347656f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_121 C N_VPWR_c_247_n 0.0223741f $X=1.68 $Y=2.405 $X2=0 $Y2=0
cc_122 N_C_M1000_g N_VPWR_c_248_n 0.00203551f $X=1.6 $Y=2.045 $X2=0 $Y2=0
cc_123 C N_VPWR_c_248_n 0.0909454f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_124 C N_VPWR_c_251_n 0.00988231f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_125 C N_VPWR_c_246_n 0.00927996f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_126 N_C_M1004_g N_VGND_c_293_n 0.0126039f $X=1.6 $Y=0.475 $X2=0 $Y2=0
cc_127 N_C_M1004_g N_VGND_c_294_n 0.00555245f $X=1.6 $Y=0.475 $X2=0 $Y2=0
cc_128 N_C_M1004_g N_VGND_c_297_n 0.00646315f $X=1.6 $Y=0.475 $X2=0 $Y2=0
cc_129 N_A_61_367#_c_166_n N_VPWR_c_247_n 0.0188586f $X=1.185 $Y=1.69 $X2=0
+ $Y2=0
cc_130 N_A_61_367#_M1003_g N_VPWR_c_248_n 0.0291959f $X=2.385 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_A_61_367#_c_171_n N_VPWR_c_248_n 0.0316193f $X=2.23 $Y=1.47 $X2=0 $Y2=0
cc_132 N_A_61_367#_c_172_n N_VPWR_c_248_n 0.00628191f $X=2.385 $Y=1.47 $X2=0
+ $Y2=0
cc_133 N_A_61_367#_M1003_g N_VPWR_c_252_n 0.00525069f $X=2.385 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_61_367#_M1003_g N_VPWR_c_246_n 0.00981609f $X=2.385 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_61_367#_M1001_g X 0.00365917f $X=2.195 $Y=0.685 $X2=0 $Y2=0
cc_136 N_A_61_367#_c_168_n X 0.00755745f $X=2.035 $Y=1.305 $X2=0 $Y2=0
cc_137 N_A_61_367#_c_171_n X 0.0261531f $X=2.23 $Y=1.47 $X2=0 $Y2=0
cc_138 N_A_61_367#_c_172_n X 0.0201044f $X=2.385 $Y=1.47 $X2=0 $Y2=0
cc_139 N_A_61_367#_M1001_g N_X_c_275_n 0.00368004f $X=2.195 $Y=0.685 $X2=0 $Y2=0
cc_140 N_A_61_367#_c_168_n X 0.00730356f $X=2.035 $Y=1.305 $X2=0 $Y2=0
cc_141 N_A_61_367#_c_171_n X 0.00234263f $X=2.23 $Y=1.47 $X2=0 $Y2=0
cc_142 N_A_61_367#_c_172_n X 0.00719266f $X=2.385 $Y=1.47 $X2=0 $Y2=0
cc_143 N_A_61_367#_c_167_n N_VGND_M1004_d 0.00637277f $X=1.945 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A_61_367#_c_168_n N_VGND_M1004_d 0.00213205f $X=2.035 $Y=1.305
+ $X2=-0.19 $Y2=-0.245
cc_145 N_A_61_367#_M1001_g N_VGND_c_293_n 0.00508647f $X=2.195 $Y=0.685 $X2=0
+ $Y2=0
cc_146 N_A_61_367#_c_167_n N_VGND_c_293_n 0.0263558f $X=1.945 $Y=0.85 $X2=0
+ $Y2=0
cc_147 N_A_61_367#_c_169_n N_VGND_c_294_n 0.0231875f $X=0.455 $Y=0.475 $X2=0
+ $Y2=0
cc_148 N_A_61_367#_M1001_g N_VGND_c_296_n 0.00555245f $X=2.195 $Y=0.685 $X2=0
+ $Y2=0
cc_149 N_A_61_367#_M1001_g N_VGND_c_297_n 0.0115897f $X=2.195 $Y=0.685 $X2=0
+ $Y2=0
cc_150 N_A_61_367#_c_167_n N_VGND_c_297_n 0.0417954f $X=1.945 $Y=0.85 $X2=0
+ $Y2=0
cc_151 N_A_61_367#_c_169_n N_VGND_c_297_n 0.0177232f $X=0.455 $Y=0.475 $X2=0
+ $Y2=0
cc_152 N_VPWR_c_246_n N_X_M1003_d 0.00336915f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_153 N_VPWR_c_248_n X 0.049486f $X=2.03 $Y=1.975 $X2=0 $Y2=0
cc_154 N_VPWR_c_252_n X 0.0203165f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_155 N_VPWR_c_246_n X 0.0115856f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_156 N_X_c_275_n N_VGND_c_293_n 6.35167e-19 $X=2.41 $Y=0.42 $X2=0 $Y2=0
cc_157 N_X_c_275_n N_VGND_c_296_n 0.0357f $X=2.41 $Y=0.42 $X2=0 $Y2=0
cc_158 N_X_c_275_n N_VGND_c_297_n 0.0193611f $X=2.41 $Y=0.42 $X2=0 $Y2=0
