# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__mux2i_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935000 1.425000 4.715000 1.750000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.885000 1.425000 5.670000 1.750000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.945000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.345000 0.790000 1.855000 ;
        RECT 0.610000 1.855000 1.850000 2.120000 ;
        RECT 1.680000 1.405000 2.275000 1.670000 ;
        RECT 1.680000 1.670000 1.850000 1.855000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  1.785000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.870000 1.580000 3.710000 1.920000 ;
        RECT 2.870000 1.920000 5.430000 2.090000 ;
        RECT 3.380000 0.965000 4.650000 1.075000 ;
        RECT 3.380000 1.075000 5.590000 1.245000 ;
        RECT 3.380000 1.245000 3.710000 1.580000 ;
        RECT 4.240000 2.090000 5.430000 2.100000 ;
        RECT 4.240000 2.100000 4.570000 2.735000 ;
        RECT 4.320000 0.605000 4.650000 0.965000 ;
        RECT 5.135000 2.100000 5.430000 3.075000 ;
        RECT 5.330000 0.330000 5.590000 1.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.180000  0.255000 0.630000 0.985000 ;
      RECT 0.180000  0.985000 1.130000 1.155000 ;
      RECT 0.180000  1.155000 0.440000 3.075000 ;
      RECT 0.710000  2.290000 1.040000 3.245000 ;
      RECT 0.800000  0.085000 1.130000 0.815000 ;
      RECT 0.960000  1.155000 1.130000 1.415000 ;
      RECT 0.960000  1.415000 1.435000 1.585000 ;
      RECT 1.230000  2.290000 1.560000 2.600000 ;
      RECT 1.230000  2.600000 3.475000 2.770000 ;
      RECT 1.230000  2.770000 1.560000 2.970000 ;
      RECT 1.300000  0.255000 1.530000 1.065000 ;
      RECT 1.300000  1.065000 3.210000 1.235000 ;
      RECT 1.700000  0.085000 1.920000 0.675000 ;
      RECT 1.700000  0.675000 2.850000 0.895000 ;
      RECT 1.740000  2.940000 2.070000 3.245000 ;
      RECT 2.090000  0.255000 5.160000 0.435000 ;
      RECT 2.090000  0.435000 2.420000 0.505000 ;
      RECT 2.250000  1.840000 2.580000 2.260000 ;
      RECT 2.250000  2.260000 4.070000 2.430000 ;
      RECT 2.795000  2.940000 3.125000 3.245000 ;
      RECT 3.020000  0.605000 4.140000 0.795000 ;
      RECT 3.020000  0.795000 3.210000 1.065000 ;
      RECT 3.305000  2.770000 3.475000 2.905000 ;
      RECT 3.305000  2.905000 4.965000 3.075000 ;
      RECT 3.810000  2.430000 4.070000 2.735000 ;
      RECT 4.740000  2.270000 4.965000 2.905000 ;
      RECT 4.830000  0.435000 5.160000 0.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__mux2i_2
