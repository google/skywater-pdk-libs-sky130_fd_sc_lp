* File: sky130_fd_sc_lp__bufinv_8.spice
* Created: Wed Sep  2 09:35:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__bufinv_8.pex.spice"
.subckt sky130_fd_sc_lp__bufinv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_82_23#_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A_82_23#_M1005_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1005_d N_A_82_23#_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_82_23#_M1013_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1013_d N_A_82_23#_M1014_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1016_d N_A_82_23#_M1016_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1016_d N_A_82_23#_M1022_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1023 N_VGND_M1023_d N_A_82_23#_M1023_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_A_82_23#_M1002_d N_A_876_23#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.231 AS=0.1176 PD=2.23 PS=1.12 NRD=1.428 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1008 N_A_82_23#_M1008_d N_A_876_23#_M1008_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1015 N_A_82_23#_M1008_d N_A_876_23#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1018 N_A_876_23#_M1018_d N_A_M1018_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_A_82_23#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1000_d N_A_82_23#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_A_82_23#_M1006_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1009 N_Y_M1006_d N_A_82_23#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1011_d N_A_82_23#_M1011_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1017 N_Y_M1011_d N_A_82_23#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1019 N_Y_M1019_d N_A_82_23#_M1019_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1020 N_Y_M1019_d N_A_82_23#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A_876_23#_M1001_g N_A_82_23#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1001_d N_A_876_23#_M1010_g N_A_82_23#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1021_d N_A_876_23#_M1021_g N_A_82_23#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1012 N_A_876_23#_M1012_d N_A_M1012_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=12.3463 P=16.97
*
.include "sky130_fd_sc_lp__bufinv_8.pxi.spice"
*
.ends
*
*
