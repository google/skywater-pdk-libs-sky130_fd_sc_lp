* File: sky130_fd_sc_lp__invkapwr_1.pxi.spice
* Created: Wed Sep  2 09:56:26 2020
* 
x_PM_SKY130_FD_SC_LP__INVKAPWR_1%A N_A_M1000_g N_A_M1001_g N_A_c_26_n
+ N_A_M1002_g A A A PM_SKY130_FD_SC_LP__INVKAPWR_1%A
x_PM_SKY130_FD_SC_LP__INVKAPWR_1%KAPWR N_KAPWR_M1000_d N_KAPWR_M1002_d KAPWR
+ N_KAPWR_c_57_n N_KAPWR_c_58_n N_KAPWR_c_59_n KAPWR
+ PM_SKY130_FD_SC_LP__INVKAPWR_1%KAPWR
x_PM_SKY130_FD_SC_LP__INVKAPWR_1%Y N_Y_M1001_s N_Y_M1000_s N_Y_c_78_n N_Y_c_82_n
+ Y Y Y PM_SKY130_FD_SC_LP__INVKAPWR_1%Y
x_PM_SKY130_FD_SC_LP__INVKAPWR_1%VGND N_VGND_M1001_d N_VGND_c_104_n
+ N_VGND_c_105_n VGND N_VGND_c_106_n N_VGND_c_107_n
+ PM_SKY130_FD_SC_LP__INVKAPWR_1%VGND
x_PM_SKY130_FD_SC_LP__INVKAPWR_1%VPWR VPWR N_VPWR_c_118_n VPWR
+ PM_SKY130_FD_SC_LP__INVKAPWR_1%VPWR
cc_1 VNB N_A_M1001_g 0.0417082f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.56
cc_2 VNB N_A_c_26_n 0.102616f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.6
cc_3 VNB N_A_M1002_g 0.00312369f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.53
cc_4 VNB A 0.0438986f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_Y_c_78_n 0.00194427f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.6
cc_6 VNB Y 0.019474f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB Y 0.0178819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB Y 0.00353325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_VGND_c_104_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_105_n 0.0228715f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.56
cc_11 VNB N_VGND_c_106_n 0.0327369f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.53
cc_12 VNB N_VGND_c_107_n 0.122328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB VPWR 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.775
cc_14 VPB N_A_M1000_g 0.0407045f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.53
cc_15 VPB N_A_c_26_n 0.0173042f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.6
cc_16 VPB N_A_M1002_g 0.0453799f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.53
cc_17 VPB A 0.0114762f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_18 VPB N_KAPWR_c_57_n 0.0240449f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.53
cc_19 VPB N_KAPWR_c_58_n 0.0249745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_20 VPB N_KAPWR_c_59_n 0.0256445f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.27
cc_21 VPB N_Y_c_82_n 0.00451878f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_22 VPB Y 0.0162053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_23 VPB VPWR 0.0491993f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.775
cc_24 VPB N_VPWR_c_118_n 0.0442176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 N_A_M1000_g N_KAPWR_c_57_n 0.00793401f $X=0.535 $Y=2.53 $X2=0 $Y2=0
cc_26 N_A_c_26_n N_KAPWR_c_57_n 0.00138689f $X=0.965 $Y=1.6 $X2=0 $Y2=0
cc_27 N_A_M1002_g N_KAPWR_c_57_n 4.31856e-19 $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_28 A N_KAPWR_c_57_n 0.0149329f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_29 N_A_M1002_g N_KAPWR_c_58_n 0.00117107f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_30 N_A_M1000_g N_KAPWR_c_59_n 0.00657544f $X=0.535 $Y=2.53 $X2=0 $Y2=0
cc_31 N_A_M1002_g N_KAPWR_c_59_n 0.00758551f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_32 N_A_M1001_g N_Y_c_78_n 0.00304928f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_33 A N_Y_c_78_n 0.0835948f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_34 N_A_M1000_g N_Y_c_82_n 0.00541707f $X=0.535 $Y=2.53 $X2=0 $Y2=0
cc_35 N_A_M1002_g N_Y_c_82_n 0.00598611f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_36 N_A_M1001_g Y 0.0176135f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_37 N_A_c_26_n Y 0.009494f $X=0.965 $Y=1.6 $X2=0 $Y2=0
cc_38 N_A_c_26_n Y 0.0295942f $X=0.965 $Y=1.6 $X2=0 $Y2=0
cc_39 N_A_c_26_n Y 0.00932139f $X=0.965 $Y=1.6 $X2=0 $Y2=0
cc_40 N_A_M1002_g Y 0.0205729f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_41 N_A_M1001_g N_VGND_c_105_n 0.013725f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_42 N_A_M1001_g N_VGND_c_106_n 0.00396895f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_43 N_A_M1001_g N_VGND_c_107_n 0.00422451f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_44 A N_VGND_c_107_n 0.0151652f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_45 N_A_M1000_g VPWR 0.00318874f $X=0.535 $Y=2.53 $X2=-0.19 $Y2=-0.245
cc_46 N_A_M1002_g VPWR 0.00318874f $X=0.965 $Y=2.53 $X2=-0.19 $Y2=-0.245
cc_47 N_A_M1000_g N_VPWR_c_118_n 0.00555753f $X=0.535 $Y=2.53 $X2=0 $Y2=0
cc_48 N_A_M1002_g N_VPWR_c_118_n 0.00570944f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_49 N_KAPWR_c_59_n N_Y_M1000_s 0.00322372f $X=1.175 $Y=2.81 $X2=0 $Y2=0
cc_50 N_KAPWR_c_57_n N_Y_c_82_n 0.0286267f $X=0.32 $Y=2.345 $X2=0 $Y2=0
cc_51 N_KAPWR_c_58_n N_Y_c_82_n 0.00679416f $X=1.18 $Y=2.345 $X2=0 $Y2=0
cc_52 N_KAPWR_c_59_n N_Y_c_82_n 0.0232419f $X=1.175 $Y=2.81 $X2=0 $Y2=0
cc_53 N_KAPWR_c_58_n Y 0.0136765f $X=1.18 $Y=2.345 $X2=0 $Y2=0
cc_54 N_KAPWR_c_57_n VPWR 0.00138124f $X=0.32 $Y=2.345 $X2=-0.19 $Y2=1.655
cc_55 N_KAPWR_c_58_n VPWR 0.00126281f $X=1.18 $Y=2.345 $X2=-0.19 $Y2=1.655
cc_56 N_KAPWR_c_59_n VPWR 0.138365f $X=1.175 $Y=2.81 $X2=-0.19 $Y2=1.655
cc_57 N_KAPWR_c_57_n N_VPWR_c_118_n 0.0121699f $X=0.32 $Y=2.345 $X2=0 $Y2=0
cc_58 N_KAPWR_c_58_n N_VPWR_c_118_n 0.0114619f $X=1.18 $Y=2.345 $X2=0 $Y2=0
cc_59 N_KAPWR_c_59_n N_VPWR_c_118_n 0.003541f $X=1.175 $Y=2.81 $X2=0 $Y2=0
cc_60 Y N_VGND_c_105_n 0.0212507f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_61 N_Y_c_78_n N_VGND_c_106_n 0.00706712f $X=0.75 $Y=0.56 $X2=0 $Y2=0
cc_62 N_Y_c_78_n N_VGND_c_107_n 0.00711097f $X=0.75 $Y=0.56 $X2=0 $Y2=0
cc_63 Y N_VGND_c_107_n 0.00673873f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_64 N_Y_c_82_n VPWR 8.5012e-19 $X=0.75 $Y=2.345 $X2=-0.19 $Y2=-0.245
cc_65 N_Y_c_82_n N_VPWR_c_118_n 0.0068611f $X=0.75 $Y=2.345 $X2=0 $Y2=0
