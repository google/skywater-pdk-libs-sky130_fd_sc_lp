* File: sky130_fd_sc_lp__o211ai_2.pxi.spice
* Created: Fri Aug 28 11:02:56 2020
* 
x_PM_SKY130_FD_SC_LP__O211AI_2%C1 N_C1_c_82_n N_C1_M1009_g N_C1_M1008_g
+ N_C1_c_84_n N_C1_M1010_g N_C1_M1015_g C1 C1 N_C1_c_87_n
+ PM_SKY130_FD_SC_LP__O211AI_2%C1
x_PM_SKY130_FD_SC_LP__O211AI_2%B1 N_B1_c_126_n N_B1_M1002_g N_B1_M1003_g
+ N_B1_c_128_n N_B1_M1006_g N_B1_M1011_g B1 B1 N_B1_c_130_n N_B1_c_131_n
+ PM_SKY130_FD_SC_LP__O211AI_2%B1
x_PM_SKY130_FD_SC_LP__O211AI_2%A2 N_A2_c_178_n N_A2_M1005_g N_A2_M1007_g
+ N_A2_c_179_n N_A2_M1014_g N_A2_M1013_g N_A2_c_180_n A2 A2 N_A2_c_181_n
+ N_A2_c_182_n N_A2_c_183_n PM_SKY130_FD_SC_LP__O211AI_2%A2
x_PM_SKY130_FD_SC_LP__O211AI_2%A1 N_A1_c_237_n N_A1_M1000_g N_A1_M1001_g
+ N_A1_c_238_n N_A1_M1012_g N_A1_M1004_g N_A1_c_239_n N_A1_c_240_n A1
+ N_A1_c_242_n PM_SKY130_FD_SC_LP__O211AI_2%A1
x_PM_SKY130_FD_SC_LP__O211AI_2%VPWR N_VPWR_M1008_s N_VPWR_M1015_s N_VPWR_M1011_d
+ N_VPWR_M1001_d N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n
+ N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n VPWR N_VPWR_c_288_n
+ N_VPWR_c_289_n N_VPWR_c_290_n N_VPWR_c_280_n N_VPWR_c_292_n N_VPWR_c_293_n
+ PM_SKY130_FD_SC_LP__O211AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O211AI_2%Y N_Y_M1009_d N_Y_M1008_d N_Y_M1003_s N_Y_M1007_s
+ N_Y_c_351_n N_Y_c_393_n N_Y_c_352_n N_Y_c_386_n N_Y_c_353_n N_Y_c_354_n Y Y Y
+ Y Y Y N_Y_c_367_n Y PM_SKY130_FD_SC_LP__O211AI_2%Y
x_PM_SKY130_FD_SC_LP__O211AI_2%A_487_367# N_A_487_367#_M1007_d
+ N_A_487_367#_M1013_d N_A_487_367#_M1004_s N_A_487_367#_c_406_n
+ N_A_487_367#_c_412_n N_A_487_367#_c_407_n N_A_487_367#_c_429_n
+ N_A_487_367#_c_408_n N_A_487_367#_c_409_n N_A_487_367#_c_410_n
+ PM_SKY130_FD_SC_LP__O211AI_2%A_487_367#
x_PM_SKY130_FD_SC_LP__O211AI_2%A_31_65# N_A_31_65#_M1009_s N_A_31_65#_M1010_s
+ N_A_31_65#_M1006_s N_A_31_65#_c_442_n N_A_31_65#_c_443_n N_A_31_65#_c_444_n
+ N_A_31_65#_c_451_n N_A_31_65#_c_445_n N_A_31_65#_c_446_n
+ PM_SKY130_FD_SC_LP__O211AI_2%A_31_65#
x_PM_SKY130_FD_SC_LP__O211AI_2%A_286_65# N_A_286_65#_M1002_d N_A_286_65#_M1005_s
+ N_A_286_65#_M1000_s N_A_286_65#_c_470_n N_A_286_65#_c_471_n
+ N_A_286_65#_c_472_n N_A_286_65#_c_473_n N_A_286_65#_c_474_n
+ PM_SKY130_FD_SC_LP__O211AI_2%A_286_65#
x_PM_SKY130_FD_SC_LP__O211AI_2%VGND N_VGND_M1005_d N_VGND_M1014_d N_VGND_M1012_d
+ N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n
+ N_VGND_c_522_n N_VGND_c_523_n VGND N_VGND_c_524_n N_VGND_c_525_n
+ N_VGND_c_526_n N_VGND_c_527_n PM_SKY130_FD_SC_LP__O211AI_2%VGND
cc_1 VNB N_C1_c_82_n 0.0201579f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.275
cc_2 VNB N_C1_M1008_g 0.00302368f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_3 VNB N_C1_c_84_n 0.0159689f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.275
cc_4 VNB N_C1_M1015_g 0.00237041f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_5 VNB C1 0.0205877f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_C1_c_87_n 0.0702627f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.44
cc_7 VNB N_B1_c_126_n 0.0158295f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.275
cc_8 VNB N_B1_M1003_g 0.00257133f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_9 VNB N_B1_c_128_n 0.0194524f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.275
cc_10 VNB N_B1_M1011_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_11 VNB N_B1_c_130_n 0.0117483f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.44
cc_12 VNB N_B1_c_131_n 0.0457306f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.44
cc_13 VNB N_A2_c_178_n 0.0209132f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.275
cc_14 VNB N_A2_c_179_n 0.0150745f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.275
cc_15 VNB N_A2_c_180_n 0.00129035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_181_n 0.0705886f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.665
cc_17 VNB N_A2_c_182_n 0.0145063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_183_n 0.00302006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_237_n 0.0150745f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.275
cc_20 VNB N_A1_c_238_n 0.0212386f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.275
cc_21 VNB N_A1_c_239_n 0.00153477f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.44
cc_22 VNB N_A1_c_240_n 0.00129035f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.44
cc_23 VNB A1 0.0401833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_242_n 0.0718416f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.665
cc_25 VNB N_VPWR_c_280_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB Y 0.0011264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_31_65#_c_442_n 0.0241979f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_28 VNB N_A_31_65#_c_443_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_31_65#_c_444_n 0.00955931f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_A_31_65#_c_445_n 0.00890199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_31_65#_c_446_n 0.00138314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_286_65#_c_470_n 0.00992764f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.745
cc_33 VNB N_A_286_65#_c_471_n 0.00140017f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_34 VNB N_A_286_65#_c_472_n 0.00615342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_286_65#_c_473_n 0.00140017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_286_65#_c_474_n 0.00110528f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.295
cc_37 VNB N_VGND_c_517_n 0.00743735f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_38 VNB N_VGND_c_518_n 7.15834e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_39 VNB N_VGND_c_519_n 0.0343095f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.44
cc_40 VNB N_VGND_c_520_n 0.013269f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.44
cc_41 VNB N_VGND_c_521_n 0.00469972f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.44
cc_42 VNB N_VGND_c_522_n 0.013269f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.295
cc_43 VNB N_VGND_c_523_n 0.00532387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_524_n 0.0583799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_525_n 0.0134401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_526_n 0.280627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_527_n 0.00532387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_C1_M1008_g 0.0251188f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_49 VPB N_C1_M1015_g 0.0186943f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_50 VPB C1 0.00764551f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_51 VPB N_B1_M1003_g 0.0191231f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_52 VPB N_B1_M1011_g 0.0251964f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_53 VPB N_A2_M1007_g 0.024771f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_54 VPB N_A2_M1013_g 0.0189785f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_55 VPB N_A2_c_181_n 0.00444146f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=1.665
cc_56 VPB N_A1_M1001_g 0.0183535f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_57 VPB N_A1_M1004_g 0.0245761f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_58 VPB N_A1_c_242_n 0.00444228f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=1.665
cc_59 VPB N_VPWR_c_281_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_60 VPB N_VPWR_c_282_n 0.0482554f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_61 VPB N_VPWR_c_283_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.44
cc_62 VPB N_VPWR_c_284_n 0.0127521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_285_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_286_n 0.0364572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_287_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_288_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_289_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_290_n 0.0236496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_280_n 0.0658237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_292_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_293_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_Y_c_351_n 0.00426037f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_73 VPB N_Y_c_352_n 0.0250152f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.44
cc_74 VPB N_Y_c_353_n 8.77875e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_Y_c_354_n 0.00162876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB Y 6.3801e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_487_367#_c_406_n 0.00804601f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_78 VPB N_A_487_367#_c_407_n 0.00194261f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_79 VPB N_A_487_367#_c_408_n 0.0124462f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.44
cc_80 VPB N_A_487_367#_c_409_n 0.00340953f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.44
cc_81 VPB N_A_487_367#_c_410_n 0.0433415f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.44
cc_82 N_C1_c_84_n N_B1_c_126_n 0.0156538f $X=0.925 $Y=1.275 $X2=-0.19 $Y2=-0.245
cc_83 N_C1_M1015_g N_B1_M1003_g 0.0232709f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_84 N_C1_c_84_n N_B1_c_130_n 0.00281761f $X=0.925 $Y=1.275 $X2=0 $Y2=0
cc_85 N_C1_c_87_n N_B1_c_131_n 0.0197002f $X=0.925 $Y=1.44 $X2=0 $Y2=0
cc_86 N_C1_M1008_g N_VPWR_c_282_n 0.0203882f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_87 N_C1_M1015_g N_VPWR_c_282_n 7.73851e-19 $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_88 C1 N_VPWR_c_282_n 0.0268575f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_89 N_C1_c_87_n N_VPWR_c_282_n 0.00156499f $X=0.925 $Y=1.44 $X2=0 $Y2=0
cc_90 N_C1_M1008_g N_VPWR_c_283_n 7.25756e-19 $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_91 N_C1_M1015_g N_VPWR_c_283_n 0.0141914f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_92 N_C1_M1008_g N_VPWR_c_288_n 0.00486043f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_93 N_C1_M1015_g N_VPWR_c_288_n 0.00486043f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_94 N_C1_M1008_g N_VPWR_c_280_n 0.00824727f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_95 N_C1_M1015_g N_VPWR_c_280_n 0.00824727f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_96 N_C1_M1015_g N_Y_c_351_n 0.0141566f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_97 N_C1_M1008_g N_Y_c_353_n 0.00237496f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_98 N_C1_M1015_g N_Y_c_353_n 0.00227113f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_99 N_C1_c_82_n Y 0.00635526f $X=0.495 $Y=1.275 $X2=0 $Y2=0
cc_100 N_C1_c_84_n Y 0.00252456f $X=0.925 $Y=1.275 $X2=0 $Y2=0
cc_101 N_C1_c_82_n Y 0.00169907f $X=0.495 $Y=1.275 $X2=0 $Y2=0
cc_102 N_C1_M1008_g Y 0.00131041f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_103 N_C1_c_84_n Y 0.00280302f $X=0.925 $Y=1.275 $X2=0 $Y2=0
cc_104 N_C1_M1015_g Y 0.00415694f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_105 C1 Y 0.0400764f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_106 N_C1_c_87_n Y 0.0206299f $X=0.925 $Y=1.44 $X2=0 $Y2=0
cc_107 N_C1_c_82_n N_Y_c_367_n 0.00441594f $X=0.495 $Y=1.275 $X2=0 $Y2=0
cc_108 N_C1_c_84_n N_Y_c_367_n 0.0041995f $X=0.925 $Y=1.275 $X2=0 $Y2=0
cc_109 C1 N_A_31_65#_c_442_n 0.0247205f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_110 N_C1_c_87_n N_A_31_65#_c_442_n 0.00169895f $X=0.925 $Y=1.44 $X2=0 $Y2=0
cc_111 N_C1_c_82_n N_A_31_65#_c_443_n 0.0125695f $X=0.495 $Y=1.275 $X2=0 $Y2=0
cc_112 N_C1_c_84_n N_A_31_65#_c_443_n 0.0119687f $X=0.925 $Y=1.275 $X2=0 $Y2=0
cc_113 N_C1_c_82_n N_VGND_c_524_n 0.00302501f $X=0.495 $Y=1.275 $X2=0 $Y2=0
cc_114 N_C1_c_84_n N_VGND_c_524_n 0.00302501f $X=0.925 $Y=1.275 $X2=0 $Y2=0
cc_115 N_C1_c_82_n N_VGND_c_526_n 0.00471248f $X=0.495 $Y=1.275 $X2=0 $Y2=0
cc_116 N_C1_c_84_n N_VGND_c_526_n 0.00435646f $X=0.925 $Y=1.275 $X2=0 $Y2=0
cc_117 N_B1_c_128_n N_A2_c_181_n 8.36064e-19 $X=1.785 $Y=1.275 $X2=0 $Y2=0
cc_118 N_B1_c_130_n N_A2_c_181_n 3.12906e-19 $X=1.74 $Y=1.44 $X2=0 $Y2=0
cc_119 N_B1_c_131_n N_A2_c_181_n 0.00404661f $X=1.785 $Y=1.44 $X2=0 $Y2=0
cc_120 N_B1_c_128_n N_A2_c_182_n 8.45562e-19 $X=1.785 $Y=1.275 $X2=0 $Y2=0
cc_121 N_B1_c_130_n N_A2_c_182_n 0.0281513f $X=1.74 $Y=1.44 $X2=0 $Y2=0
cc_122 N_B1_c_131_n N_A2_c_182_n 0.00405429f $X=1.785 $Y=1.44 $X2=0 $Y2=0
cc_123 N_B1_M1003_g N_VPWR_c_283_n 0.0141914f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B1_M1011_g N_VPWR_c_283_n 7.25756e-19 $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B1_M1003_g N_VPWR_c_284_n 7.25756e-19 $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B1_M1011_g N_VPWR_c_284_n 0.0159418f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B1_M1003_g N_VPWR_c_289_n 0.00486043f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_128 N_B1_M1011_g N_VPWR_c_289_n 0.00486043f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_129 N_B1_M1003_g N_VPWR_c_280_n 0.00824727f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_130 N_B1_M1011_g N_VPWR_c_280_n 0.00824727f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_131 N_B1_M1003_g N_Y_c_351_n 0.0134905f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_132 N_B1_c_130_n N_Y_c_351_n 0.0254721f $X=1.74 $Y=1.44 $X2=0 $Y2=0
cc_133 N_B1_c_131_n N_Y_c_351_n 0.00106178f $X=1.785 $Y=1.44 $X2=0 $Y2=0
cc_134 N_B1_M1011_g N_Y_c_352_n 0.0155776f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_135 N_B1_c_130_n N_Y_c_352_n 0.0134993f $X=1.74 $Y=1.44 $X2=0 $Y2=0
cc_136 N_B1_c_131_n N_Y_c_352_n 0.00106178f $X=1.785 $Y=1.44 $X2=0 $Y2=0
cc_137 N_B1_c_130_n N_Y_c_354_n 0.012542f $X=1.74 $Y=1.44 $X2=0 $Y2=0
cc_138 N_B1_c_131_n N_Y_c_354_n 0.00248053f $X=1.785 $Y=1.44 $X2=0 $Y2=0
cc_139 N_B1_M1003_g Y 7.50734e-19 $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_140 N_B1_c_130_n Y 0.0259326f $X=1.74 $Y=1.44 $X2=0 $Y2=0
cc_141 N_B1_c_131_n Y 6.54318e-19 $X=1.785 $Y=1.44 $X2=0 $Y2=0
cc_142 N_B1_c_126_n N_Y_c_367_n 8.79119e-19 $X=1.355 $Y=1.275 $X2=0 $Y2=0
cc_143 N_B1_M1011_g N_A_487_367#_c_406_n 0.00139782f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_B1_c_130_n N_A_31_65#_c_451_n 0.0152553f $X=1.74 $Y=1.44 $X2=0 $Y2=0
cc_145 N_B1_c_126_n N_A_31_65#_c_445_n 0.0155889f $X=1.355 $Y=1.275 $X2=0 $Y2=0
cc_146 N_B1_c_128_n N_A_31_65#_c_445_n 0.0144613f $X=1.785 $Y=1.275 $X2=0 $Y2=0
cc_147 N_B1_c_130_n N_A_31_65#_c_445_n 0.00431892f $X=1.74 $Y=1.44 $X2=0 $Y2=0
cc_148 N_B1_c_126_n N_A_286_65#_c_470_n 0.00278809f $X=1.355 $Y=1.275 $X2=0
+ $Y2=0
cc_149 N_B1_c_128_n N_A_286_65#_c_470_n 0.012131f $X=1.785 $Y=1.275 $X2=0 $Y2=0
cc_150 N_B1_c_130_n N_A_286_65#_c_470_n 0.030256f $X=1.74 $Y=1.44 $X2=0 $Y2=0
cc_151 N_B1_c_131_n N_A_286_65#_c_470_n 5.96813e-19 $X=1.785 $Y=1.44 $X2=0 $Y2=0
cc_152 N_B1_c_128_n N_VGND_c_517_n 0.00184346f $X=1.785 $Y=1.275 $X2=0 $Y2=0
cc_153 N_B1_c_126_n N_VGND_c_524_n 0.00302501f $X=1.355 $Y=1.275 $X2=0 $Y2=0
cc_154 N_B1_c_128_n N_VGND_c_524_n 0.00302501f $X=1.785 $Y=1.275 $X2=0 $Y2=0
cc_155 N_B1_c_126_n N_VGND_c_526_n 0.00435646f $X=1.355 $Y=1.275 $X2=0 $Y2=0
cc_156 N_B1_c_128_n N_VGND_c_526_n 0.0048466f $X=1.785 $Y=1.275 $X2=0 $Y2=0
cc_157 N_A2_c_179_n N_A1_c_237_n 0.0201362f $X=3.205 $Y=1.21 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A2_M1013_g N_A1_M1001_g 0.0201362f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A2_c_180_n N_A1_c_240_n 0.00950855f $X=3.115 $Y=1.505 $X2=0 $Y2=0
cc_160 N_A2_c_181_n N_A1_c_240_n 2.12265e-19 $X=3.205 $Y=1.44 $X2=0 $Y2=0
cc_161 N_A2_c_180_n N_A1_c_242_n 2.12265e-19 $X=3.115 $Y=1.505 $X2=0 $Y2=0
cc_162 N_A2_c_181_n N_A1_c_242_n 0.0201362f $X=3.205 $Y=1.44 $X2=0 $Y2=0
cc_163 N_A2_M1007_g N_VPWR_c_284_n 0.00214936f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A2_M1013_g N_VPWR_c_285_n 0.00109252f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A2_M1007_g N_VPWR_c_286_n 0.00357877f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A2_M1013_g N_VPWR_c_286_n 0.00357877f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A2_M1007_g N_VPWR_c_280_n 0.00665089f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A2_M1013_g N_VPWR_c_280_n 0.00537654f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A2_M1007_g N_Y_c_352_n 0.0148281f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A2_M1013_g N_Y_c_352_n 0.00295925f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A2_c_180_n N_Y_c_352_n 0.0264029f $X=3.115 $Y=1.505 $X2=0 $Y2=0
cc_172 N_A2_c_181_n N_Y_c_352_n 0.00414098f $X=3.205 $Y=1.44 $X2=0 $Y2=0
cc_173 N_A2_c_182_n N_Y_c_352_n 0.0587936f $X=2.538 $Y=1.392 $X2=0 $Y2=0
cc_174 N_A2_M1007_g N_Y_c_386_n 0.0144173f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A2_M1013_g N_Y_c_386_n 0.00845257f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A2_M1007_g N_A_487_367#_c_412_n 0.0114565f $X=2.775 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A2_M1013_g N_A_487_367#_c_412_n 0.0115031f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A2_M1013_g N_A_487_367#_c_409_n 6.13138e-19 $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A2_c_178_n N_A_31_65#_c_445_n 9.55167e-19 $X=2.775 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A2_c_178_n N_A_286_65#_c_470_n 0.0142607f $X=2.775 $Y=1.21 $X2=0 $Y2=0
cc_181 N_A2_c_180_n N_A_286_65#_c_470_n 0.00475695f $X=3.115 $Y=1.505 $X2=0
+ $Y2=0
cc_182 N_A2_c_181_n N_A_286_65#_c_470_n 0.00143281f $X=3.205 $Y=1.44 $X2=0 $Y2=0
cc_183 N_A2_c_182_n N_A_286_65#_c_470_n 0.0509949f $X=2.538 $Y=1.392 $X2=0 $Y2=0
cc_184 N_A2_c_178_n N_A_286_65#_c_471_n 6.56187e-19 $X=2.775 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A2_c_179_n N_A_286_65#_c_471_n 6.56187e-19 $X=3.205 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A2_c_179_n N_A_286_65#_c_472_n 0.0101357f $X=3.205 $Y=1.21 $X2=0 $Y2=0
cc_187 N_A2_c_180_n N_A_286_65#_c_472_n 0.0131833f $X=3.115 $Y=1.505 $X2=0 $Y2=0
cc_188 N_A2_c_181_n N_A_286_65#_c_472_n 0.00383431f $X=3.205 $Y=1.44 $X2=0 $Y2=0
cc_189 N_A2_c_178_n N_A_286_65#_c_474_n 0.00311892f $X=2.775 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A2_c_180_n N_A_286_65#_c_474_n 0.0137115f $X=3.115 $Y=1.505 $X2=0 $Y2=0
cc_191 N_A2_c_181_n N_A_286_65#_c_474_n 0.00634873f $X=3.205 $Y=1.44 $X2=0 $Y2=0
cc_192 N_A2_c_183_n N_A_286_65#_c_474_n 0.00458153f $X=2.735 $Y=1.392 $X2=0
+ $Y2=0
cc_193 N_A2_c_178_n N_VGND_c_517_n 0.0102853f $X=2.775 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A2_c_179_n N_VGND_c_517_n 5.14896e-19 $X=3.205 $Y=1.21 $X2=0 $Y2=0
cc_195 N_A2_c_178_n N_VGND_c_518_n 5.63271e-19 $X=2.775 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A2_c_179_n N_VGND_c_518_n 0.010882f $X=3.205 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A2_c_178_n N_VGND_c_520_n 0.00465098f $X=2.775 $Y=1.21 $X2=0 $Y2=0
cc_198 N_A2_c_179_n N_VGND_c_520_n 0.00465098f $X=3.205 $Y=1.21 $X2=0 $Y2=0
cc_199 N_A2_c_178_n N_VGND_c_526_n 0.00443946f $X=2.775 $Y=1.21 $X2=0 $Y2=0
cc_200 N_A2_c_179_n N_VGND_c_526_n 0.00822759f $X=3.205 $Y=1.21 $X2=0 $Y2=0
cc_201 N_A1_M1001_g N_VPWR_c_285_n 0.0153413f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A1_M1004_g N_VPWR_c_285_n 0.0161459f $X=4.065 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A1_M1001_g N_VPWR_c_286_n 0.00486043f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A1_M1004_g N_VPWR_c_290_n 0.00486043f $X=4.065 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A1_M1001_g N_VPWR_c_280_n 0.0082726f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A1_M1004_g N_VPWR_c_280_n 0.00935029f $X=4.065 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A1_M1001_g N_A_487_367#_c_408_n 0.0129567f $X=3.635 $Y=2.465 $X2=0
+ $Y2=0
cc_208 N_A1_M1004_g N_A_487_367#_c_408_n 0.0137084f $X=4.065 $Y=2.465 $X2=0
+ $Y2=0
cc_209 N_A1_c_239_n N_A_487_367#_c_408_n 0.0231891f $X=4.305 $Y=1.4 $X2=0 $Y2=0
cc_210 N_A1_c_240_n N_A_487_367#_c_408_n 0.0440106f $X=4.115 $Y=1.4 $X2=0 $Y2=0
cc_211 N_A1_c_242_n N_A_487_367#_c_408_n 0.00417724f $X=4.065 $Y=1.44 $X2=0
+ $Y2=0
cc_212 N_A1_c_237_n N_A_286_65#_c_472_n 0.0101567f $X=3.635 $Y=1.21 $X2=0 $Y2=0
cc_213 N_A1_c_238_n N_A_286_65#_c_472_n 0.00349191f $X=4.065 $Y=1.21 $X2=0 $Y2=0
cc_214 N_A1_c_239_n N_A_286_65#_c_472_n 0.00327024f $X=4.305 $Y=1.4 $X2=0 $Y2=0
cc_215 N_A1_c_240_n N_A_286_65#_c_472_n 0.0276566f $X=4.115 $Y=1.4 $X2=0 $Y2=0
cc_216 N_A1_c_242_n N_A_286_65#_c_472_n 0.0103512f $X=4.065 $Y=1.44 $X2=0 $Y2=0
cc_217 N_A1_c_237_n N_A_286_65#_c_473_n 6.56187e-19 $X=3.635 $Y=1.21 $X2=0 $Y2=0
cc_218 N_A1_c_238_n N_A_286_65#_c_473_n 6.56187e-19 $X=4.065 $Y=1.21 $X2=0 $Y2=0
cc_219 N_A1_c_237_n N_VGND_c_518_n 0.0108921f $X=3.635 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A1_c_238_n N_VGND_c_518_n 5.89866e-19 $X=4.065 $Y=1.21 $X2=0 $Y2=0
cc_221 N_A1_c_237_n N_VGND_c_519_n 6.26644e-19 $X=3.635 $Y=1.21 $X2=0 $Y2=0
cc_222 N_A1_c_238_n N_VGND_c_519_n 0.0162439f $X=4.065 $Y=1.21 $X2=0 $Y2=0
cc_223 N_A1_c_239_n N_VGND_c_519_n 0.0250514f $X=4.305 $Y=1.4 $X2=0 $Y2=0
cc_224 N_A1_c_242_n N_VGND_c_519_n 0.00506784f $X=4.065 $Y=1.44 $X2=0 $Y2=0
cc_225 N_A1_c_237_n N_VGND_c_522_n 0.00465098f $X=3.635 $Y=1.21 $X2=0 $Y2=0
cc_226 N_A1_c_238_n N_VGND_c_522_n 0.00465098f $X=4.065 $Y=1.21 $X2=0 $Y2=0
cc_227 N_A1_c_237_n N_VGND_c_526_n 0.00822759f $X=3.635 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A1_c_238_n N_VGND_c_526_n 0.00822759f $X=4.065 $Y=1.21 $X2=0 $Y2=0
cc_229 N_VPWR_c_280_n N_Y_M1008_d 0.00536646f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_230 N_VPWR_c_280_n N_Y_M1003_s 0.00536646f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_231 N_VPWR_c_280_n N_Y_M1007_s 0.00225186f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_232 N_VPWR_M1015_s N_Y_c_351_n 0.00176461f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_233 N_VPWR_c_283_n N_Y_c_351_n 0.0170777f $X=1.14 $Y=2.185 $X2=0 $Y2=0
cc_234 N_VPWR_c_289_n N_Y_c_393_n 0.0124525f $X=1.835 $Y=3.33 $X2=0 $Y2=0
cc_235 N_VPWR_c_280_n N_Y_c_393_n 0.00730901f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_236 N_VPWR_M1011_d N_Y_c_352_n 0.00265333f $X=1.86 $Y=1.835 $X2=0 $Y2=0
cc_237 N_VPWR_c_284_n N_Y_c_352_n 0.0220026f $X=2 $Y=2.185 $X2=0 $Y2=0
cc_238 N_VPWR_c_288_n Y 0.0124525f $X=0.975 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_c_280_n Y 0.00730901f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_240 N_VPWR_c_280_n N_A_487_367#_M1007_d 0.00215161f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_241 N_VPWR_c_280_n N_A_487_367#_M1013_d 0.00376627f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_280_n N_A_487_367#_M1004_s 0.00371702f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_284_n N_A_487_367#_c_406_n 0.0532774f $X=2 $Y=2.185 $X2=0 $Y2=0
cc_244 N_VPWR_c_286_n N_A_487_367#_c_412_n 0.0361172f $X=3.685 $Y=3.33 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_280_n N_A_487_367#_c_412_n 0.023676f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_246 N_VPWR_c_284_n N_A_487_367#_c_407_n 0.0121616f $X=2 $Y=2.185 $X2=0 $Y2=0
cc_247 N_VPWR_c_286_n N_A_487_367#_c_407_n 0.0179183f $X=3.685 $Y=3.33 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_280_n N_A_487_367#_c_407_n 0.0101082f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_286_n N_A_487_367#_c_429_n 0.0125234f $X=3.685 $Y=3.33 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_280_n N_A_487_367#_c_429_n 0.00738676f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_251 N_VPWR_M1001_d N_A_487_367#_c_408_n 0.00176461f $X=3.71 $Y=1.835 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_285_n N_A_487_367#_c_408_n 0.0170777f $X=3.85 $Y=2.185 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_290_n N_A_487_367#_c_410_n 0.0178111f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_280_n N_A_487_367#_c_410_n 0.0100304f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_255 N_Y_c_352_n N_A_487_367#_M1007_d 0.00265333f $X=2.825 $Y=1.845 $X2=-0.19
+ $Y2=-0.245
cc_256 N_Y_c_352_n N_A_487_367#_c_406_n 0.0202165f $X=2.825 $Y=1.845 $X2=0 $Y2=0
cc_257 N_Y_M1007_s N_A_487_367#_c_412_n 0.00332344f $X=2.85 $Y=1.835 $X2=0 $Y2=0
cc_258 N_Y_c_386_n N_A_487_367#_c_412_n 0.0159805f $X=2.99 $Y=1.97 $X2=0 $Y2=0
cc_259 N_Y_c_352_n N_A_487_367#_c_409_n 0.0106597f $X=2.825 $Y=1.845 $X2=0 $Y2=0
cc_260 N_Y_M1009_d N_A_31_65#_c_443_n 0.00176461f $X=0.57 $Y=0.325 $X2=0 $Y2=0
cc_261 N_Y_c_367_n N_A_31_65#_c_443_n 0.0159533f $X=0.71 $Y=0.68 $X2=0 $Y2=0
cc_262 N_A_487_367#_c_408_n N_A_286_65#_c_472_n 0.00156656f $X=4.185 $Y=1.845
+ $X2=0 $Y2=0
cc_263 N_A_487_367#_c_409_n N_A_286_65#_c_472_n 0.00748144f $X=3.515 $Y=1.845
+ $X2=0 $Y2=0
cc_264 N_A_31_65#_c_445_n N_A_286_65#_M1002_d 0.00172844f $X=2 $Y=0.48 $X2=-0.19
+ $Y2=-0.245
cc_265 N_A_31_65#_M1006_s N_A_286_65#_c_470_n 0.00989588f $X=1.86 $Y=0.325 $X2=0
+ $Y2=0
cc_266 N_A_31_65#_c_445_n N_A_286_65#_c_470_n 0.0442327f $X=2 $Y=0.48 $X2=0
+ $Y2=0
cc_267 N_A_31_65#_c_445_n N_VGND_c_517_n 0.0277572f $X=2 $Y=0.48 $X2=0 $Y2=0
cc_268 N_A_31_65#_c_443_n N_VGND_c_524_n 0.0422287f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_269 N_A_31_65#_c_444_n N_VGND_c_524_n 0.0200723f $X=0.375 $Y=0.34 $X2=0 $Y2=0
cc_270 N_A_31_65#_c_445_n N_VGND_c_524_n 0.0625346f $X=2 $Y=0.48 $X2=0 $Y2=0
cc_271 N_A_31_65#_c_446_n N_VGND_c_524_n 0.0136205f $X=1.14 $Y=0.47 $X2=0 $Y2=0
cc_272 N_A_31_65#_c_443_n N_VGND_c_526_n 0.0238173f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_273 N_A_31_65#_c_444_n N_VGND_c_526_n 0.0108858f $X=0.375 $Y=0.34 $X2=0 $Y2=0
cc_274 N_A_31_65#_c_445_n N_VGND_c_526_n 0.0342537f $X=2 $Y=0.48 $X2=0 $Y2=0
cc_275 N_A_31_65#_c_446_n N_VGND_c_526_n 0.00738676f $X=1.14 $Y=0.47 $X2=0 $Y2=0
cc_276 N_A_286_65#_c_470_n N_VGND_M1005_d 0.00502116f $X=2.895 $Y=0.92 $X2=-0.19
+ $Y2=-0.245
cc_277 N_A_286_65#_c_472_n N_VGND_M1014_d 0.00176461f $X=3.755 $Y=1.165 $X2=0
+ $Y2=0
cc_278 N_A_286_65#_c_470_n N_VGND_c_517_n 0.0217739f $X=2.895 $Y=0.92 $X2=0
+ $Y2=0
cc_279 N_A_286_65#_c_471_n N_VGND_c_517_n 0.0147868f $X=2.99 $Y=0.42 $X2=0 $Y2=0
cc_280 N_A_286_65#_c_471_n N_VGND_c_518_n 0.0211656f $X=2.99 $Y=0.42 $X2=0 $Y2=0
cc_281 N_A_286_65#_c_472_n N_VGND_c_518_n 0.0170777f $X=3.755 $Y=1.165 $X2=0
+ $Y2=0
cc_282 N_A_286_65#_c_473_n N_VGND_c_518_n 0.0247302f $X=3.85 $Y=0.42 $X2=0 $Y2=0
cc_283 N_A_286_65#_c_473_n N_VGND_c_519_n 0.0296081f $X=3.85 $Y=0.42 $X2=0 $Y2=0
cc_284 N_A_286_65#_c_471_n N_VGND_c_520_n 0.0134771f $X=2.99 $Y=0.42 $X2=0 $Y2=0
cc_285 N_A_286_65#_c_473_n N_VGND_c_522_n 0.0134771f $X=3.85 $Y=0.42 $X2=0 $Y2=0
cc_286 N_A_286_65#_c_470_n N_VGND_c_526_n 0.0157096f $X=2.895 $Y=0.92 $X2=0
+ $Y2=0
cc_287 N_A_286_65#_c_471_n N_VGND_c_526_n 0.00730901f $X=2.99 $Y=0.42 $X2=0
+ $Y2=0
cc_288 N_A_286_65#_c_473_n N_VGND_c_526_n 0.00730901f $X=3.85 $Y=0.42 $X2=0
+ $Y2=0
