* File: sky130_fd_sc_lp__decapkapwr_4.pex.spice
* Created: Wed Sep  2 09:42:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_4%VGND 1 7 9 11 14 17 19 26 29 32 42
r31 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r32 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 36 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r34 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 33 38 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.25
+ $Y2=0
r36 33 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=1.2 $Y2=0
r37 32 41 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.685
+ $Y2=0
r38 32 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.2
+ $Y2=0
r39 29 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r40 29 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r41 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.77 $X2=0.575 $Y2=1.77
r42 23 26 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.335 $Y=1.77
+ $X2=0.575 $Y2=1.77
r43 19 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.615 $Y=0.36
+ $X2=1.615 $Y2=1.04
r44 17 41 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.685 $Y2=0
r45 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0.36
r46 14 16 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.335 $Y=0.38
+ $X2=0.335 $Y2=1.06
r47 12 23 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.335 $Y=1.605
+ $X2=0.335 $Y2=1.77
r48 12 16 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.335 $Y=1.605
+ $X2=0.335 $Y2=1.06
r49 11 38 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.25 $Y2=0
r50 11 14 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.38
r51 7 27 22.6591 $w=1e-06 $l=4.09268e-07 $layer=POLY_cond $X=0.91 $Y=1.935
+ $X2=0.575 $Y2=1.77
r52 7 9 33.9353 $w=1e-06 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.935 $X2=0.91
+ $Y2=2.595
r53 1 21 121.333 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=1.615 $Y2=1.04
r54 1 19 121.333 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=1.615 $Y2=0.36
r55 1 16 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=0.335 $Y2=1.06
r56 1 14 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=0.335 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_4%KAPWR 1 7 9 11 13 14 16 23 26 34
r36 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.705 $Y=2.81
+ $X2=1.705 $Y2=2.81
r37 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.215 $Y=2.81
+ $X2=0.215 $Y2=2.81
r38 23 34 0.407181 $w=2.7e-07 $l=7.45e-07 $layer=MET1_cond $X=0.96 $Y=2.81
+ $X2=1.705 $Y2=2.81
r39 23 30 0.407181 $w=2.7e-07 $l=7.45e-07 $layer=MET1_cond $X=0.96 $Y=2.81
+ $X2=0.215 $Y2=2.81
r40 19 26 44.365 $w=8.68e-07 $l=9.34987e-07 $layer=POLY_cond $X=1.345 $Y=1.51
+ $X2=0.992 $Y2=0.735
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.345
+ $Y=1.51 $X2=1.345 $Y2=1.51
r42 14 33 3.07376 $w=4.05e-07 $l=2e-07 $layer=LI1_cond $X=1.587 $Y=2.675
+ $X2=1.587 $Y2=2.875
r43 14 16 10.9553 $w=4.03e-07 $l=3.85e-07 $layer=LI1_cond $X=1.587 $Y=2.675
+ $X2=1.587 $Y2=2.29
r44 13 18 8.32511 $w=3.33e-07 $l=2.42e-07 $layer=LI1_cond $X=1.587 $Y=1.507
+ $X2=1.345 $Y2=1.507
r45 13 16 17.5001 $w=4.03e-07 $l=6.15e-07 $layer=LI1_cond $X=1.587 $Y=1.675
+ $X2=1.587 $Y2=2.29
r46 12 29 3.69365 $w=2.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.425 $Y=2.81
+ $X2=0.26 $Y2=2.875
r47 11 33 4.10347 $w=2.7e-07 $l=2.32237e-07 $layer=LI1_cond $X=1.385 $Y=2.81
+ $X2=1.587 $Y2=2.875
r48 11 12 40.9757 $w=2.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.385 $Y=2.81
+ $X2=0.425 $Y2=2.81
r49 7 29 3.21187 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=0.26 $Y=2.675 $X2=0.26
+ $Y2=2.875
r50 7 9 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.26 $Y=2.675
+ $X2=0.26 $Y2=2.27
r51 1 33 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.095 $X2=1.55 $Y2=2.97
r52 1 29 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.095 $X2=0.26 $Y2=2.95
r53 1 16 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.095 $X2=1.55 $Y2=2.29
r54 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.095 $X2=0.26 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_4%VPWR 1 8 14
r14 5 14 0.0081048 $w=1.92e-06 $l=1.22e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.96 $Y2=3.208
r15 5 8 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33 $X2=1.68
+ $Y2=3.33
r16 4 8 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.68
+ $Y2=3.33
r17 4 5 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33 $X2=0.24
+ $Y2=3.33
r18 1 14 6.64328e-05 $w=1.92e-06 $l=1e-09 $layer=MET1_cond $X=0.96 $Y=3.207
+ $X2=0.96 $Y2=3.208
.ends

