* File: sky130_fd_sc_lp__sdfxtp_4.spice
* Created: Wed Sep  2 10:36:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfxtp_4.pex.spice"
.subckt sky130_fd_sc_lp__sdfxtp_4  VNB VPB D SCE SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* SCE	SCE
* D	D
* VPB	VPB
* VNB	VNB
MM1035 N_VGND_M1035_d N_SCE_M1035_g N_A_91_123#_M1035_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1037 A_260_123# N_A_91_123#_M1037_g N_VGND_M1035_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07245 AS=0.0588 PD=0.765 PS=0.7 NRD=33.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1030 N_A_359_123#_M1030_d N_D_M1030_g A_260_123# VNB NSHORT L=0.15 W=0.42
+ AD=0.0987 AS=0.07245 PD=0.89 PS=0.765 NRD=27.132 NRS=33.564 M=1 R=2.8
+ SA=75001.1 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1000 A_483_123# N_SCE_M1000_g N_A_359_123#_M1030_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0987 PD=0.63 PS=0.89 NRD=14.28 NRS=27.132 M=1 R=2.8 SA=75001.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_SCD_M1026_g A_483_123# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1028 N_A_641_123#_M1028_d N_CLK_M1028_g N_VGND_M1026_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1512 AS=0.0588 PD=1.56 PS=0.7 NRD=27.132 NRS=0 M=1 R=2.8
+ SA=75002.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1006 N_A_850_51#_M1006_d N_A_641_123#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_1053_125#_M1009_d N_A_641_123#_M1009_g N_A_359_123#_M1009_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.063 AS=0.1113 PD=0.72 PS=1.37 NRD=5.712 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1010 A_1143_125# N_A_850_51#_M1010_g N_A_1053_125#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.063 PD=0.72 PS=0.72 NRD=27.132 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_1203_99#_M1012_g A_1143_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.227196 AS=0.063 PD=1.35113 PS=0.72 NRD=138.84 NRS=27.132 M=1 R=2.8
+ SA=75001.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1019 N_A_1203_99#_M1019_d N_A_1053_125#_M1019_g N_VGND_M1012_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.138023 AS=0.346204 PD=1.24981 PS=2.05887 NRD=0 NRS=81.552
+ M=1 R=4.26667 SA=75001.4 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1033 N_A_1475_449#_M1033_d N_A_850_51#_M1033_g N_A_1203_99#_M1019_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.10815 AS=0.0905774 PD=0.935 PS=0.820189 NRD=67.14
+ NRS=34.284 M=1 R=2.8 SA=75001.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1034 A_1670_61# N_A_641_123#_M1034_g N_A_1475_449#_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.05775 AS=0.10815 PD=0.695 PS=0.935 NRD=23.568 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1673_409#_M1029_g A_1670_61# VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.05775 PD=0.81 PS=0.695 NRD=28.56 NRS=23.568 M=1 R=2.8
+ SA=75002.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_A_1673_409#_M1013_d N_A_1475_449#_M1013_g N_VGND_M1029_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A_1673_409#_M1005_g N_Q_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1014_d N_A_1673_409#_M1014_g N_Q_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1014_d N_A_1673_409#_M1017_g N_Q_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1025 N_VGND_M1025_d N_A_1673_409#_M1025_g N_Q_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1027 N_VPWR_M1027_d N_SCE_M1027_g N_A_91_123#_M1027_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1016 A_296_491# N_SCE_M1016_g N_VPWR_M1027_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1020 N_A_359_123#_M1020_d N_D_M1020_g A_296_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 A_454_491# N_A_91_123#_M1007_g N_A_359_123#_M1020_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=32.308 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_SCD_M1001_g A_454_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1008 AS=0.1024 PD=0.955 PS=0.96 NRD=10.7562 NRS=32.308 M=1 R=4.26667
+ SA=75001.9 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1031 N_A_641_123#_M1031_d N_CLK_M1031_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1008 PD=1.81 PS=0.955 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_A_850_51#_M1003_d N_A_641_123#_M1003_g N_VPWR_M1003_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.3424 PD=1.81 PS=2.35 NRD=0 NRS=83.0946 M=1
+ R=4.26667 SA=75000.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_1053_125#_M1008_d N_A_850_51#_M1008_g N_A_359_123#_M1008_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.10745 AS=0.1113 PD=0.96 PS=1.37 NRD=44.5417 NRS=0
+ M=1 R=2.8 SA=75000.2 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1022 A_1199_449# N_A_641_123#_M1022_g N_A_1053_125#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.10745 PD=0.63 PS=0.96 NRD=23.443 NRS=44.5417 M=1 R=2.8
+ SA=75000.7 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_1203_99#_M1021_g A_1199_449# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.123333 AS=0.0441 PD=0.926667 PS=0.63 NRD=111.935 NRS=23.443 M=1 R=2.8
+ SA=75001.1 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1002 N_A_1203_99#_M1002_d N_A_1053_125#_M1002_g N_VPWR_M1021_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.246667 PD=1.12 PS=1.85333 NRD=0 NRS=19.9167 M=1
+ R=5.6 SA=75001 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1023 N_A_1475_449#_M1023_d N_A_641_123#_M1023_g N_A_1203_99#_M1002_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2464 AS=0.1176 PD=1.96 PS=1.12 NRD=82.0702 NRS=0
+ M=1 R=5.6 SA=75001.4 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1032 A_1631_507# N_A_850_51#_M1032_g N_A_1475_449#_M1023_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1232 PD=0.63 PS=0.98 NRD=23.443 NRS=0 M=1 R=2.8 SA=75002
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_1673_409#_M1018_g A_1631_507# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.131775 AS=0.0441 PD=0.9725 PS=0.63 NRD=192.292 NRS=23.443 M=1
+ R=2.8 SA=75002.3 SB=75001 A=0.063 P=1.14 MULT=1
MM1015 N_A_1673_409#_M1015_d N_A_1475_449#_M1015_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.395325 PD=3.05 PS=2.9175 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A_1673_409#_M1004_g N_Q_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_1673_409#_M1011_g N_Q_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1024 N_VPWR_M1011_d N_A_1673_409#_M1024_g N_Q_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1036 N_VPWR_M1036_d N_A_1673_409#_M1036_g N_Q_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX38_noxref VNB VPB NWDIODE A=23.2371 P=28.77
c_132 VNB 0 3.22859e-19 $X=0 $Y=0
c_243 VPB 0 1.42881e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfxtp_4.pxi.spice"
*
.ends
*
*
