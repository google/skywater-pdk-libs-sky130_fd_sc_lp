* File: sky130_fd_sc_lp__clkinv_2.pxi.spice
* Created: Fri Aug 28 10:17:54 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINV_2%A N_A_M1001_g N_A_M1002_g N_A_M1000_g N_A_M1004_g
+ N_A_M1003_g A A N_A_c_36_n N_A_c_37_n PM_SKY130_FD_SC_LP__CLKINV_2%A
x_PM_SKY130_FD_SC_LP__CLKINV_2%Y N_Y_M1000_d N_Y_M1001_s N_Y_M1002_s N_Y_c_112_p
+ N_Y_c_84_n N_Y_c_85_n N_Y_c_113_p N_Y_c_79_n N_Y_c_86_n N_Y_c_87_n N_Y_c_80_n
+ Y Y N_Y_c_83_n PM_SKY130_FD_SC_LP__CLKINV_2%Y
x_PM_SKY130_FD_SC_LP__CLKINV_2%VPWR N_VPWR_M1001_d N_VPWR_M1004_d N_VPWR_c_125_n
+ N_VPWR_c_126_n N_VPWR_c_127_n VPWR N_VPWR_c_128_n N_VPWR_c_129_n
+ N_VPWR_c_130_n N_VPWR_c_124_n PM_SKY130_FD_SC_LP__CLKINV_2%VPWR
x_PM_SKY130_FD_SC_LP__CLKINV_2%VGND N_VGND_M1000_s N_VGND_M1003_s N_VGND_c_151_n
+ N_VGND_c_152_n N_VGND_c_153_n VGND N_VGND_c_154_n N_VGND_c_155_n
+ N_VGND_c_156_n N_VGND_c_157_n PM_SKY130_FD_SC_LP__CLKINV_2%VGND
cc_1 VNB N_A_M1000_g 0.0525956f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.56
cc_2 VNB N_A_M1003_g 0.0435876f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=0.56
cc_3 VNB N_A_c_36_n 0.0293436f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.46
cc_4 VNB N_A_c_37_n 0.084547f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.485
cc_5 VNB N_Y_c_79_n 0.00149799f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.485
cc_6 VNB N_Y_c_80_n 0.00456845f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.485
cc_7 VNB Y 0.00295631f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.46
cc_8 VNB Y 0.0291489f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.485
cc_9 VNB N_Y_c_83_n 0.0103855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VPWR_c_124_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.377
cc_11 VNB N_VGND_c_151_n 0.0256902f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.295
cc_12 VNB N_VGND_c_152_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.56
cc_13 VNB N_VGND_c_153_n 0.0222797f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.675
cc_14 VNB N_VGND_c_154_n 0.0223503f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=1.295
cc_15 VNB N_VGND_c_155_n 0.0160313f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_16 VNB N_VGND_c_156_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.46
cc_17 VNB N_VGND_c_157_n 0.152942f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.46
cc_18 VPB N_A_M1001_g 0.0233545f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_19 VPB N_A_M1002_g 0.0176925f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_20 VPB N_A_M1004_g 0.0223382f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_21 VPB N_A_c_37_n 0.00870531f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.485
cc_22 VPB N_Y_c_84_n 0.00234264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_23 VPB N_Y_c_85_n 0.0176848f $X=-0.19 $Y=1.655 $X2=1.445 $Y2=1.295
cc_24 VPB N_Y_c_86_n 0.0132482f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.46
cc_25 VPB N_Y_c_87_n 0.00209286f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.485
cc_26 VPB Y 0.00298715f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.485
cc_27 VPB N_VPWR_c_125_n 0.00461568f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.295
cc_28 VPB N_VPWR_c_126_n 0.0142571f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.675
cc_29 VPB N_VPWR_c_127_n 0.00460237f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_30 VPB N_VPWR_c_128_n 0.0183554f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_31 VPB N_VPWR_c_129_n 0.0167406f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.485
cc_32 VPB N_VPWR_c_130_n 0.00497514f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=1.46
cc_33 VPB N_VPWR_c_124_n 0.051331f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.377
cc_34 N_A_M1001_g N_Y_c_84_n 0.0153265f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_35 N_A_M1002_g N_Y_c_84_n 0.0143812f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_36 N_A_c_36_n N_Y_c_84_n 0.0436107f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_37 N_A_c_37_n N_Y_c_84_n 0.002829f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_38 N_A_M1000_g N_Y_c_79_n 0.00189162f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_39 N_A_M1003_g N_Y_c_79_n 0.00180689f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_40 N_A_M1004_g N_Y_c_86_n 0.0159989f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_41 N_A_c_36_n N_Y_c_86_n 0.0110823f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_42 N_A_c_37_n N_Y_c_86_n 0.00322171f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_43 N_A_c_36_n N_Y_c_87_n 0.0219511f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_44 N_A_c_37_n N_Y_c_87_n 0.00314903f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_45 N_A_M1000_g N_Y_c_80_n 0.006617f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_46 N_A_c_36_n N_Y_c_80_n 0.0198419f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_47 N_A_c_37_n N_Y_c_80_n 6.24756e-19 $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_48 N_A_M1003_g Y 0.0152312f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_49 N_A_c_36_n Y 0.00755553f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_50 N_A_M1003_g Y 0.0205853f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_51 N_A_c_36_n Y 0.0267298f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_52 N_A_c_37_n Y 0.00240773f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_53 N_A_M1001_g N_VPWR_c_125_n 0.00309734f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_54 N_A_M1002_g N_VPWR_c_125_n 0.0016342f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_55 N_A_M1004_g N_VPWR_c_127_n 0.00341773f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_56 N_A_M1001_g N_VPWR_c_128_n 0.00585385f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_57 N_A_M1002_g N_VPWR_c_129_n 0.00585385f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_58 N_A_M1004_g N_VPWR_c_129_n 0.00585385f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VPWR_c_124_n 0.0116543f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_VPWR_c_124_n 0.0106302f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_61 N_A_M1004_g N_VPWR_c_124_n 0.0116375f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_VGND_c_151_n 0.00406185f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_63 N_A_c_36_n N_VGND_c_151_n 0.0110952f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_64 N_A_c_37_n N_VGND_c_151_n 0.00153298f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_65 N_A_M1000_g N_VGND_c_153_n 5.44985e-19 $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_66 N_A_M1003_g N_VGND_c_153_n 0.00957799f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_67 N_A_M1000_g N_VGND_c_155_n 0.00478016f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_68 N_A_M1003_g N_VGND_c_155_n 0.00396895f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_69 N_A_M1000_g N_VGND_c_157_n 0.0096052f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_70 N_A_M1003_g N_VGND_c_157_n 0.00397666f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_71 N_Y_c_84_n N_VPWR_M1001_d 0.00176461f $X=1.01 $Y=1.8 $X2=-0.19 $Y2=-0.245
cc_72 N_Y_c_86_n N_VPWR_M1004_d 0.00246823f $X=1.595 $Y=1.8 $X2=0 $Y2=0
cc_73 N_Y_c_84_n N_VPWR_c_125_n 0.0135055f $X=1.01 $Y=1.8 $X2=0 $Y2=0
cc_74 N_Y_c_86_n N_VPWR_c_127_n 0.0176763f $X=1.595 $Y=1.8 $X2=0 $Y2=0
cc_75 N_Y_c_112_p N_VPWR_c_128_n 0.0135826f $X=0.28 $Y=2 $X2=0 $Y2=0
cc_76 N_Y_c_113_p N_VPWR_c_129_n 0.012556f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_77 N_Y_M1001_s N_VPWR_c_124_n 0.00254606f $X=0.155 $Y=1.835 $X2=0 $Y2=0
cc_78 N_Y_M1002_s N_VPWR_c_124_n 0.00302905f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_79 N_Y_c_112_p N_VPWR_c_124_n 0.00969167f $X=0.28 $Y=2 $X2=0 $Y2=0
cc_80 N_Y_c_113_p N_VPWR_c_124_n 0.00988321f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_81 Y N_VGND_c_153_n 0.00530131f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_82 N_Y_c_83_n N_VGND_c_153_n 0.0165893f $X=1.687 $Y=1.04 $X2=0 $Y2=0
cc_83 N_Y_c_79_n N_VGND_c_155_n 0.00717541f $X=1.23 $Y=0.56 $X2=0 $Y2=0
cc_84 N_Y_c_79_n N_VGND_c_157_n 0.00799322f $X=1.23 $Y=0.56 $X2=0 $Y2=0
cc_85 Y N_VGND_c_157_n 0.00538134f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_86 N_Y_c_83_n N_VGND_c_157_n 6.73317e-19 $X=1.687 $Y=1.04 $X2=0 $Y2=0
