* File: sky130_fd_sc_lp__nand3b_1.pxi.spice
* Created: Fri Aug 28 10:49:44 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3B_1%A_N N_A_N_M1005_g N_A_N_M1004_g A_N N_A_N_c_47_n
+ N_A_N_c_48_n PM_SKY130_FD_SC_LP__NAND3B_1%A_N
x_PM_SKY130_FD_SC_LP__NAND3B_1%C N_C_M1002_g N_C_M1007_g C N_C_c_75_n N_C_c_78_n
+ PM_SKY130_FD_SC_LP__NAND3B_1%C
x_PM_SKY130_FD_SC_LP__NAND3B_1%B N_B_M1003_g N_B_M1000_g B N_B_c_107_n
+ N_B_c_108_n PM_SKY130_FD_SC_LP__NAND3B_1%B
x_PM_SKY130_FD_SC_LP__NAND3B_1%A_84_131# N_A_84_131#_M1005_s N_A_84_131#_M1004_s
+ N_A_84_131#_M1006_g N_A_84_131#_M1001_g N_A_84_131#_c_142_n
+ N_A_84_131#_c_143_n N_A_84_131#_c_144_n N_A_84_131#_c_150_n
+ N_A_84_131#_c_145_n N_A_84_131#_c_146_n N_A_84_131#_c_147_n
+ PM_SKY130_FD_SC_LP__NAND3B_1%A_84_131#
x_PM_SKY130_FD_SC_LP__NAND3B_1%VPWR N_VPWR_M1004_d N_VPWR_M1003_d N_VPWR_c_198_n
+ N_VPWR_c_199_n N_VPWR_c_200_n N_VPWR_c_201_n N_VPWR_c_202_n N_VPWR_c_203_n
+ VPWR N_VPWR_c_204_n N_VPWR_c_197_n PM_SKY130_FD_SC_LP__NAND3B_1%VPWR
x_PM_SKY130_FD_SC_LP__NAND3B_1%Y N_Y_M1006_d N_Y_M1007_d N_Y_M1001_d N_Y_c_231_n
+ N_Y_c_233_n N_Y_c_236_n Y Y Y Y Y Y Y Y N_Y_c_228_n
+ PM_SKY130_FD_SC_LP__NAND3B_1%Y
x_PM_SKY130_FD_SC_LP__NAND3B_1%VGND N_VGND_M1005_d N_VGND_c_265_n N_VGND_c_266_n
+ N_VGND_c_267_n VGND N_VGND_c_268_n N_VGND_c_269_n
+ PM_SKY130_FD_SC_LP__NAND3B_1%VGND
cc_1 VNB N_A_N_M1005_g 0.0319121f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.865
cc_2 VNB N_A_N_c_47_n 0.0262629f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.51
cc_3 VNB N_A_N_c_48_n 0.00176211f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.51
cc_4 VNB N_C_M1002_g 0.0274268f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.865
cc_5 VNB N_C_c_75_n 0.0253514f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.51
cc_6 VNB N_B_M1000_g 0.0240206f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.045
cc_7 VNB N_B_c_107_n 0.0239395f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.51
cc_8 VNB N_B_c_108_n 0.00176211f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.51
cc_9 VNB N_A_84_131#_M1001_g 0.00777961f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.51
cc_10 VNB N_A_84_131#_c_142_n 0.0199061f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.675
cc_11 VNB N_A_84_131#_c_143_n 0.0387922f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.51
cc_12 VNB N_A_84_131#_c_144_n 0.0336875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_84_131#_c_145_n 0.00316314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_84_131#_c_146_n 0.0349348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_84_131#_c_147_n 0.0198338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_197_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB Y 0.0387571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_228_n 0.0337381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_265_n 0.0171306f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.045
cc_20 VNB N_VGND_c_266_n 0.0282373f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.51
cc_21 VNB N_VGND_c_267_n 0.00711686f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.51
cc_22 VNB N_VGND_c_268_n 0.0506028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_269_n 0.182284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VPB N_A_N_M1004_g 0.0294525f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.045
cc_25 VPB N_A_N_c_47_n 0.0065075f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.51
cc_26 VPB N_A_N_c_48_n 0.0044482f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.51
cc_27 VPB N_C_M1007_g 0.022164f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.045
cc_28 VPB N_C_c_75_n 0.00648093f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.51
cc_29 VPB N_C_c_78_n 0.00340787f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.51
cc_30 VPB N_B_M1003_g 0.0189618f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.865
cc_31 VPB N_B_c_107_n 0.00632607f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.51
cc_32 VPB N_B_c_108_n 0.00334344f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.51
cc_33 VPB N_A_84_131#_M1001_g 0.0241647f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.51
cc_34 VPB N_A_84_131#_c_142_n 0.0137762f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.675
cc_35 VPB N_A_84_131#_c_150_n 0.0258825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_198_n 0.034417f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_37 VPB N_VPWR_c_199_n 0.00233412f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.675
cc_38 VPB N_VPWR_c_200_n 0.0301467f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.665
cc_39 VPB N_VPWR_c_201_n 0.00574121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_202_n 0.0170386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_203_n 0.00519718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_204_n 0.02026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_197_n 0.0780881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB Y 0.0582653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB Y 0.0144375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 N_A_N_M1005_g N_C_M1002_g 0.0172594f $X=0.76 $Y=0.865 $X2=0 $Y2=0
cc_47 N_A_N_M1004_g N_C_M1007_g 0.0136549f $X=0.76 $Y=2.045 $X2=0 $Y2=0
cc_48 N_A_N_c_47_n N_C_c_75_n 0.0215729f $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_49 N_A_N_c_48_n N_C_c_75_n 0.00142573f $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_50 N_A_N_M1004_g N_C_c_78_n 2.59842e-19 $X=0.76 $Y=2.045 $X2=0 $Y2=0
cc_51 N_A_N_c_47_n N_C_c_78_n 2.88395e-19 $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_52 N_A_N_c_48_n N_C_c_78_n 0.0262648f $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_53 N_A_N_M1005_g N_A_84_131#_c_142_n 0.00250416f $X=0.76 $Y=0.865 $X2=0 $Y2=0
cc_54 N_A_N_M1004_g N_A_84_131#_c_142_n 0.00413488f $X=0.76 $Y=2.045 $X2=0 $Y2=0
cc_55 N_A_N_c_47_n N_A_84_131#_c_142_n 0.00854217f $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_56 N_A_N_c_48_n N_A_84_131#_c_142_n 0.0239191f $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_57 N_A_N_M1005_g N_A_84_131#_c_143_n 0.0167027f $X=0.76 $Y=0.865 $X2=0 $Y2=0
cc_58 N_A_N_M1005_g N_A_84_131#_c_144_n 4.27702e-19 $X=0.76 $Y=0.865 $X2=0 $Y2=0
cc_59 N_A_N_c_47_n N_A_84_131#_c_144_n 0.00454115f $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_60 N_A_N_c_48_n N_A_84_131#_c_144_n 0.0282684f $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_61 N_A_N_M1004_g N_A_84_131#_c_150_n 0.00429565f $X=0.76 $Y=2.045 $X2=0 $Y2=0
cc_62 N_A_N_c_47_n N_A_84_131#_c_150_n 9.55994e-19 $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_63 N_A_N_c_48_n N_A_84_131#_c_150_n 0.0141221f $X=0.67 $Y=1.51 $X2=0 $Y2=0
cc_64 N_A_N_M1004_g N_VPWR_c_198_n 0.00366436f $X=0.76 $Y=2.045 $X2=0 $Y2=0
cc_65 N_A_N_M1005_g N_VGND_c_265_n 0.0141352f $X=0.76 $Y=0.865 $X2=0 $Y2=0
cc_66 N_A_N_M1005_g N_VGND_c_266_n 0.00359024f $X=0.76 $Y=0.865 $X2=0 $Y2=0
cc_67 N_A_N_M1005_g N_VGND_c_269_n 0.00418172f $X=0.76 $Y=0.865 $X2=0 $Y2=0
cc_68 N_C_M1007_g N_B_M1003_g 0.0188528f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_69 N_C_M1002_g N_B_M1000_g 0.0538164f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_70 N_C_c_75_n N_B_c_107_n 0.0215729f $X=1.21 $Y=1.51 $X2=0 $Y2=0
cc_71 N_C_c_78_n N_B_c_107_n 2.88395e-19 $X=1.21 $Y=1.51 $X2=0 $Y2=0
cc_72 N_C_c_75_n N_B_c_108_n 0.00186964f $X=1.21 $Y=1.51 $X2=0 $Y2=0
cc_73 N_C_c_78_n N_B_c_108_n 0.0259188f $X=1.21 $Y=1.51 $X2=0 $Y2=0
cc_74 N_C_M1002_g N_A_84_131#_c_143_n 0.0156709f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_75 N_C_c_75_n N_A_84_131#_c_143_n 0.00443962f $X=1.21 $Y=1.51 $X2=0 $Y2=0
cc_76 N_C_c_78_n N_A_84_131#_c_143_n 0.0241855f $X=1.21 $Y=1.51 $X2=0 $Y2=0
cc_77 N_C_M1007_g N_VPWR_c_198_n 0.00632283f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_78 N_C_c_75_n N_VPWR_c_198_n 8.37776e-19 $X=1.21 $Y=1.51 $X2=0 $Y2=0
cc_79 N_C_c_78_n N_VPWR_c_198_n 0.011076f $X=1.21 $Y=1.51 $X2=0 $Y2=0
cc_80 N_C_M1007_g N_VPWR_c_202_n 0.0054895f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_81 N_C_M1007_g N_VPWR_c_197_n 0.0110907f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_82 N_C_M1007_g N_Y_c_231_n 0.00209314f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_83 N_C_c_78_n N_Y_c_231_n 0.00192368f $X=1.21 $Y=1.51 $X2=0 $Y2=0
cc_84 N_C_M1007_g N_Y_c_233_n 0.0117938f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_85 N_C_M1002_g N_VGND_c_265_n 0.00676437f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_86 N_C_M1002_g N_VGND_c_268_n 0.00585385f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_87 N_C_M1002_g N_VGND_c_269_n 0.0120894f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_88 N_B_M1003_g N_A_84_131#_M1001_g 0.0319177f $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_89 N_B_c_108_n N_A_84_131#_M1001_g 8.27458e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_90 N_B_M1000_g N_A_84_131#_c_143_n 0.0152051f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_91 N_B_c_107_n N_A_84_131#_c_143_n 0.00454708f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_92 N_B_c_108_n N_A_84_131#_c_143_n 0.02736f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_93 N_B_M1000_g N_A_84_131#_c_145_n 6.73426e-19 $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_94 N_B_c_107_n N_A_84_131#_c_145_n 8.87114e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_95 N_B_c_108_n N_A_84_131#_c_145_n 0.0056352f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_96 N_B_c_107_n N_A_84_131#_c_146_n 0.0207536f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_97 N_B_c_108_n N_A_84_131#_c_146_n 9.51592e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_98 N_B_M1000_g N_A_84_131#_c_147_n 0.0549488f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_99 N_B_M1003_g N_VPWR_c_199_n 0.00291503f $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_100 N_B_M1003_g N_VPWR_c_202_n 0.00583607f $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_101 N_B_M1003_g N_VPWR_c_197_n 0.0106324f $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_102 N_B_c_107_n N_Y_c_231_n 2.28961e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_103 N_B_c_108_n N_Y_c_231_n 0.00607567f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_104 N_B_M1003_g N_Y_c_236_n 0.0131658f $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_105 N_B_c_107_n N_Y_c_236_n 5.1995e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_106 N_B_c_108_n N_Y_c_236_n 0.0180034f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_107 N_B_c_108_n Y 0.00704184f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_108 N_B_M1000_g N_Y_c_228_n 0.00334754f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_109 N_B_M1000_g N_VGND_c_268_n 0.00585385f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_110 N_B_M1000_g N_VGND_c_269_n 0.011138f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_111 N_A_84_131#_c_143_n N_VPWR_c_198_n 0.00486676f $X=2.125 $Y=1.17 $X2=0
+ $Y2=0
cc_112 N_A_84_131#_M1001_g N_VPWR_c_199_n 0.0155086f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_84_131#_M1001_g N_VPWR_c_204_n 0.00544582f $X=2.2 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_84_131#_M1001_g N_VPWR_c_197_n 0.0102513f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_84_131#_c_143_n N_Y_c_231_n 0.00432421f $X=2.125 $Y=1.17 $X2=0 $Y2=0
cc_116 N_A_84_131#_M1001_g N_Y_c_236_n 0.0141146f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_84_131#_c_143_n N_Y_c_236_n 0.00506761f $X=2.125 $Y=1.17 $X2=0 $Y2=0
cc_118 N_A_84_131#_c_145_n N_Y_c_236_n 0.00607732f $X=2.25 $Y=1.17 $X2=0 $Y2=0
cc_119 N_A_84_131#_c_145_n Y 0.00224207f $X=2.25 $Y=1.17 $X2=0 $Y2=0
cc_120 N_A_84_131#_c_146_n Y 0.00316214f $X=2.29 $Y=1.35 $X2=0 $Y2=0
cc_121 N_A_84_131#_M1001_g Y 0.00834263f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_84_131#_c_145_n Y 0.0330156f $X=2.25 $Y=1.17 $X2=0 $Y2=0
cc_123 N_A_84_131#_c_146_n Y 0.00821274f $X=2.29 $Y=1.35 $X2=0 $Y2=0
cc_124 N_A_84_131#_c_147_n Y 0.00351952f $X=2.29 $Y=1.185 $X2=0 $Y2=0
cc_125 N_A_84_131#_c_145_n N_Y_c_228_n 0.011781f $X=2.25 $Y=1.17 $X2=0 $Y2=0
cc_126 N_A_84_131#_c_146_n N_Y_c_228_n 0.00365125f $X=2.29 $Y=1.35 $X2=0 $Y2=0
cc_127 N_A_84_131#_c_147_n N_Y_c_228_n 0.0176737f $X=2.29 $Y=1.185 $X2=0 $Y2=0
cc_128 N_A_84_131#_c_143_n N_VGND_c_265_n 0.0267957f $X=2.125 $Y=1.17 $X2=0
+ $Y2=0
cc_129 N_A_84_131#_c_147_n N_VGND_c_268_n 0.00482548f $X=2.29 $Y=1.185 $X2=0
+ $Y2=0
cc_130 N_A_84_131#_c_144_n N_VGND_c_269_n 0.0201697f $X=0.65 $Y=1.01 $X2=0 $Y2=0
cc_131 N_A_84_131#_c_147_n N_VGND_c_269_n 0.00949816f $X=2.29 $Y=1.185 $X2=0
+ $Y2=0
cc_132 N_VPWR_c_197_n N_Y_M1007_d 0.00293134f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_133 N_VPWR_c_197_n N_Y_M1001_d 0.00336915f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_134 N_VPWR_c_202_n N_Y_c_233_n 0.0165751f $X=1.805 $Y=3.33 $X2=0 $Y2=0
cc_135 N_VPWR_c_197_n N_Y_c_233_n 0.0108194f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_136 N_VPWR_M1003_d N_Y_c_236_n 0.00587357f $X=1.805 $Y=1.835 $X2=0 $Y2=0
cc_137 N_VPWR_c_199_n N_Y_c_236_n 0.0174033f $X=1.97 $Y=2.365 $X2=0 $Y2=0
cc_138 N_VPWR_c_204_n Y 0.0335785f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_139 N_VPWR_c_197_n Y 0.0187779f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_140 N_Y_c_228_n N_VGND_c_268_n 0.0349786f $X=2.415 $Y=0.38 $X2=0 $Y2=0
cc_141 N_Y_M1006_d N_VGND_c_269_n 0.00215817f $X=2.275 $Y=0.235 $X2=0 $Y2=0
cc_142 N_Y_c_228_n N_VGND_c_269_n 0.0222253f $X=2.415 $Y=0.38 $X2=0 $Y2=0
cc_143 N_VGND_c_269_n A_275_47# 0.0130629f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_144 N_VGND_c_269_n A_366_47# 0.0126346f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
