* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_27_519# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_27_519# a_254_55# a_284_81# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_710_117# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR S1 a_1245_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_284_81# S0 a_196_519# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_793_117# a_254_55# a_968_501# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_799_501# S0 a_793_117# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_968_501# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_212_81# a_254_55# a_284_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_284_81# S0 a_33_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_1635_149# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_1635_149# a_1245_21# a_793_117# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_793_117# a_254_55# a_879_117# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_33_81# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR A2 a_799_501# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_284_81# S1 a_1635_149# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VGND A0 a_212_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND S1 a_1245_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_710_117# S0 a_793_117# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1635_149# a_1245_21# a_284_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_1635_149# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 VPWR A0 a_196_519# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_254_55# S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_254_55# S0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_793_117# S1 a_1635_149# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND A2 a_879_117# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
