* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a22o_m A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_85_317# B2 a_265_501# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND A2 a_265_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_85_317# B1 a_445_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_445_125# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR A2 a_265_501# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 X a_85_317# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_265_501# B1 a_85_317# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_265_125# A1 a_85_317# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_85_317# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_265_501# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
