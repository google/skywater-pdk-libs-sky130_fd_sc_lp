* File: sky130_fd_sc_lp__iso1n_lp2.spice
* Created: Wed Sep  2 09:58:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__iso1n_lp2.pex.spice"
.subckt sky130_fd_sc_lp__iso1n_lp2  VNB VPB SLEEP_B A VPWR X KAGND VGND
* 
* KAGND	KAGND
* X	X
* VPWR	VPWR
* A	A
* SLEEP_B	SLEEP_B
* VPB	VPB
* VNB	VNB
MM1001 A_114_109# N_SLEEP_B_M1001_g N_A_27_109#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1006 N_KAGND_M1006_d N_SLEEP_B_M1006_g A_114_109# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1008 A_272_109# N_A_27_109#_M1008_g N_KAGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1004 N_A_350_109#_M1004_d N_A_27_109#_M1004_g A_272_109# VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 A_452_109# N_A_M1011_g N_A_350_109#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0756 PD=0.63 PS=0.78 NRD=14.28 NRS=22.848 M=1 R=2.8 SA=75001.9
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 N_KAGND_M1009_d N_A_M1009_g A_452_109# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.3 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1010 A_610_109# N_A_350_109#_M1010_g N_KAGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_350_109#_M1005_g A_610_109# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_SLEEP_B_M1000_g N_A_27_109#_M1000_s VPB PHIGHVT L=0.25
+ W=1 AD=0.16 AS=0.285 PD=1.32 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1007 A_300_409# N_A_27_109#_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.16 PD=1.24 PS=1.32 NRD=12.7853 NRS=7.8603 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1002 N_A_350_109#_M1002_d N_A_M1002_g A_300_409# VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.12 PD=2.57 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1003 N_X_M1003_d N_A_350_109#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_62 VPB 0 1.20445e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__iso1n_lp2.pxi.spice"
*
.ends
*
*
