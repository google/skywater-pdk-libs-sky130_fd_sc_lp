* File: sky130_fd_sc_lp__o221a_1.pex.spice
* Created: Fri Aug 28 11:07:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221A_1%C1 3 7 9 10 11 12 14 15 25 33
r41 27 33 2.40092 $w=2.38e-07 $l=5e-08 $layer=LI1_cond $X=0.205 $Y=1.345
+ $X2=0.205 $Y2=1.295
r42 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.42
+ $Y=1.51 $X2=0.42 $Y2=1.51
r43 14 15 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.205 $Y=2.035
+ $X2=0.205 $Y2=2.405
r44 12 25 5.12197 $w=4.03e-07 $l=1.8e-07 $layer=LI1_cond $X=0.24 $Y=1.547
+ $X2=0.42 $Y2=1.547
r45 12 27 0.995938 $w=4.03e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.547
+ $X2=0.205 $Y2=1.547
r46 12 27 3.79848 $w=2.4e-07 $l=2.03e-07 $layer=LI1_cond $X=0.205 $Y=1.75
+ $X2=0.205 $Y2=1.547
r47 12 14 9.97569 $w=4.08e-07 $l=2.85e-07 $layer=LI1_cond $X=0.205 $Y=1.75
+ $X2=0.205 $Y2=2.035
r48 12 33 0.864332 $w=2.38e-07 $l=1.8e-08 $layer=LI1_cond $X=0.205 $Y=1.277
+ $X2=0.205 $Y2=1.295
r49 11 12 16.9025 $w=2.38e-07 $l=3.52e-07 $layer=LI1_cond $X=0.205 $Y=0.925
+ $X2=0.205 $Y2=1.277
r50 9 24 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=0.745 $Y=1.51
+ $X2=0.42 $Y2=1.51
r51 9 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.745 $Y=1.51
+ $X2=0.82 $Y2=1.51
r52 5 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.82 $Y=1.675
+ $X2=0.82 $Y2=1.51
r53 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.82 $Y=1.675 $X2=0.82
+ $Y2=2.465
r54 1 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.82 $Y=1.345
+ $X2=0.82 $Y2=1.51
r55 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.82 $Y=1.345 $X2=0.82
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%B1 3 6 8 9 13 15
c40 15 0 1.46826e-19 $X=1.27 $Y=1.21
r41 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.27 $Y=1.375
+ $X2=1.27 $Y2=1.54
r42 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.27 $Y=1.375
+ $X2=1.27 $Y2=1.21
r43 8 9 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.245 $Y=1.295
+ $X2=1.245 $Y2=1.665
r44 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.375 $X2=1.27 $Y2=1.375
r45 6 16 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.36 $Y=2.465
+ $X2=1.36 $Y2=1.54
r46 3 15 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.29 $Y=0.665
+ $X2=1.29 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%B2 3 6 8 11 12 13
c37 13 0 1.78828e-19 $X=1.815 $Y=1.195
c38 12 0 1.83534e-19 $X=1.82 $Y=1.36
r39 11 14 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.36
+ $X2=1.815 $Y2=1.525
r40 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.36
+ $X2=1.815 $Y2=1.195
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.36 $X2=1.82 $Y2=1.36
r42 8 12 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.68 $Y=1.36 $X2=1.82
+ $Y2=1.36
r43 6 14 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.75 $Y=2.465 $X2=1.75
+ $Y2=1.525
r44 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.72 $Y=0.665
+ $X2=1.72 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%A2 3 6 8 9 13 15
c33 13 0 1.78828e-19 $X=2.515 $Y=1.35
c34 6 0 3.67072e-20 $X=2.67 $Y=2.465
r35 13 16 46.6684 $w=4.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.525 $Y=1.35
+ $X2=2.525 $Y2=1.515
r36 13 15 46.6684 $w=4.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.525 $Y=1.35
+ $X2=2.525 $Y2=1.185
r37 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.515
+ $Y=1.35 $X2=2.515 $Y2=1.35
r38 9 14 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.35
+ $X2=2.515 $Y2=1.35
r39 8 14 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.16 $Y=1.35
+ $X2=2.515 $Y2=1.35
r40 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.67 $Y=2.465
+ $X2=2.67 $Y2=1.515
r41 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.67 $Y=0.655
+ $X2=2.67 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%A1 3 7 8 11 13
c32 11 0 1.51321e-19 $X=3.12 $Y=1.35
c33 3 0 1.03873e-19 $X=3.03 $Y=2.465
r34 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.35
+ $X2=3.12 $Y2=1.515
r35 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.35
+ $X2=3.12 $Y2=1.185
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.35 $X2=3.12 $Y2=1.35
r37 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.1 $Y=0.655 $X2=3.1
+ $Y2=1.185
r38 3 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.03 $Y=2.465
+ $X2=3.03 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%A_96_49# 1 2 3 12 15 19 23 26 27 28 31 33 36
+ 39 45 53 54 57
r98 54 58 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=3.692 $Y=1.35
+ $X2=3.692 $Y2=1.515
r99 54 57 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=3.692 $Y=1.35
+ $X2=3.692 $Y2=1.185
r100 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.67
+ $Y=1.35 $X2=3.67 $Y2=1.35
r101 50 53 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.48 $Y=1.35
+ $X2=3.67 $Y2=1.35
r102 48 49 0.50437 $w=8.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.215 $Y=1.98
+ $X2=2.215 $Y2=2.015
r103 45 48 2.88212 $w=8.28e-07 $l=2e-07 $layer=LI1_cond $X=2.215 $Y=1.78
+ $X2=2.215 $Y2=1.98
r104 42 44 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.605 $Y=2.015
+ $X2=0.85 $Y2=2.015
r105 35 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.48 $Y=1.515
+ $X2=3.48 $Y2=1.35
r106 35 36 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.48 $Y=1.515
+ $X2=3.48 $Y2=1.695
r107 34 45 10.4562 $w=1.7e-07 $l=4.15e-07 $layer=LI1_cond $X=2.63 $Y=1.78
+ $X2=2.215 $Y2=1.78
r108 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.395 $Y=1.78
+ $X2=3.48 $Y2=1.695
r109 33 34 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.395 $Y=1.78
+ $X2=2.63 $Y2=1.78
r110 29 49 1.2249 $w=8.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=2.1
+ $X2=2.215 $Y2=2.015
r111 29 31 11.6726 $w=8.28e-07 $l=8.1e-07 $layer=LI1_cond $X=2.215 $Y=2.1
+ $X2=2.215 $Y2=2.91
r112 28 44 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=2.015
+ $X2=0.85 $Y2=2.015
r113 27 49 10.4562 $w=1.7e-07 $l=4.15e-07 $layer=LI1_cond $X=1.8 $Y=2.015
+ $X2=2.215 $Y2=2.015
r114 27 28 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.8 $Y=2.015
+ $X2=0.935 $Y2=2.015
r115 26 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=1.93
+ $X2=0.85 $Y2=2.015
r116 25 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=1.175
+ $X2=0.85 $Y2=1.09
r117 25 26 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.85 $Y=1.175
+ $X2=0.85 $Y2=1.93
r118 23 42 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=0.625 $Y=2.91
+ $X2=0.625 $Y2=2.1
r119 17 39 15.5273 $w=1.68e-07 $l=2.38e-07 $layer=LI1_cond $X=0.612 $Y=1.09
+ $X2=0.85 $Y2=1.09
r120 17 19 28.6885 $w=2.33e-07 $l=5.85e-07 $layer=LI1_cond $X=0.612 $Y=1.005
+ $X2=0.612 $Y2=0.42
r121 15 58 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.605 $Y=2.465
+ $X2=3.605 $Y2=1.515
r122 12 57 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.57 $Y=0.655
+ $X2=3.57 $Y2=1.185
r123 3 48 200 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=3 $X=1.825
+ $Y=1.835 $X2=1.965 $Y2=1.98
r124 3 31 200 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=3 $X=1.825
+ $Y=1.835 $X2=1.965 $Y2=2.91
r125 2 42 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.48
+ $Y=1.835 $X2=0.605 $Y2=2.095
r126 2 23 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.48
+ $Y=1.835 $X2=0.605 $Y2=2.91
r127 1 19 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=0.48
+ $Y=0.245 $X2=0.605 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%VPWR 1 2 9 13 18 19 20 22 32 33 36
r44 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r47 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=1.09 $Y2=3.33
r49 27 29 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 25 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.09 $Y2=3.33
r53 22 24 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 20 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 20 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 18 29 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.14 $Y=3.33 $X2=3.12
+ $Y2=3.33
r57 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=3.33
+ $X2=3.305 $Y2=3.33
r58 17 32 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.47 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.47 $Y=3.33
+ $X2=3.305 $Y2=3.33
r60 13 16 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.305 $Y=2.12
+ $X2=3.305 $Y2=2.95
r61 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=3.245
+ $X2=3.305 $Y2=3.33
r62 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=3.245
+ $X2=3.305 $Y2=2.95
r63 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=3.245 $X2=1.09
+ $Y2=3.33
r64 7 9 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=1.09 $Y=3.245 $X2=1.09
+ $Y2=2.375
r65 2 16 400 $w=1.7e-07 $l=1.21088e-06 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=1.835 $X2=3.305 $Y2=2.95
r66 2 13 400 $w=1.7e-07 $l=3.71786e-07 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=1.835 $X2=3.305 $Y2=2.12
r67 1 9 300 $w=1.7e-07 $l=6.3e-07 $layer=licon1_PDIFF $count=2 $X=0.895 $Y=1.835
+ $X2=1.09 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%X 1 2 7 8 9 10 11 12 13 28 29 38
c25 29 0 1.03873e-19 $X=3.945 $Y=2.315
r26 23 28 1.11527 $w=3.08e-07 $l=3e-08 $layer=LI1_cond $X=4.08 $Y=1.695 $X2=4.08
+ $Y2=1.665
r27 13 33 7.01149 $w=5.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.945 $Y=2.775
+ $X2=3.945 $Y2=2.435
r28 12 33 0.618661 $w=5.78e-07 $l=3e-08 $layer=LI1_cond $X=3.945 $Y=2.405
+ $X2=3.945 $Y2=2.435
r29 12 29 1.85598 $w=5.78e-07 $l=9e-08 $layer=LI1_cond $X=3.945 $Y=2.405
+ $X2=3.945 $Y2=2.315
r30 11 29 5.97626 $w=5.8e-07 $l=2.8e-07 $layer=LI1_cond $X=3.945 $Y=2.035
+ $X2=3.945 $Y2=2.315
r31 11 47 1.24953 $w=5.37e-07 $l=5.5e-08 $layer=LI1_cond $X=3.945 $Y=2.035
+ $X2=3.945 $Y2=1.98
r32 10 47 5.86145 $w=5.37e-07 $l=2.58e-07 $layer=LI1_cond $X=3.945 $Y=1.722
+ $X2=3.945 $Y2=1.98
r33 10 23 2.77513 $w=5.37e-07 $l=1.47885e-07 $layer=LI1_cond $X=3.945 $Y=1.722
+ $X2=4.08 $Y2=1.695
r34 10 28 1.04092 $w=3.08e-07 $l=2.8e-08 $layer=LI1_cond $X=4.08 $Y=1.637
+ $X2=4.08 $Y2=1.665
r35 9 10 12.714 $w=3.08e-07 $l=3.42e-07 $layer=LI1_cond $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.637
r36 9 44 10.4092 $w=3.08e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.015
r37 8 44 4.46876 $w=5.83e-07 $l=9e-08 $layer=LI1_cond $X=3.942 $Y=0.925
+ $X2=3.942 $Y2=1.015
r38 7 8 7.56494 $w=5.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.942 $Y=0.555
+ $X2=3.942 $Y2=0.925
r39 7 38 2.76018 $w=5.83e-07 $l=1.35e-07 $layer=LI1_cond $X=3.942 $Y=0.555
+ $X2=3.942 $Y2=0.42
r40 2 47 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.68
+ $Y=1.835 $X2=3.82 $Y2=1.98
r41 2 33 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=3.68
+ $Y=1.835 $X2=3.82 $Y2=2.435
r42 1 38 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.645
+ $Y=0.235 $X2=3.785 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%A_179_49# 1 2 9 12 13
r24 13 16 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.935 $Y=0.34
+ $X2=1.935 $Y2=0.55
r25 10 12 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=0.34
+ $X2=1.065 $Y2=0.34
r26 9 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=0.34
+ $X2=1.935 $Y2=0.34
r27 9 10 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.77 $Y=0.34 $X2=1.23
+ $Y2=0.34
r28 2 16 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.795
+ $Y=0.245 $X2=1.935 $Y2=0.55
r29 1 12 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=0.895
+ $Y=0.245 $X2=1.065 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%A_273_49# 1 2 7 11 14
c22 7 0 1.51321e-19 $X=2.79 $Y=0.93
r23 14 16 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.5 $Y=0.76 $X2=1.5
+ $Y2=0.93
r24 9 11 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=2.885 $Y=0.845
+ $X2=2.885 $Y2=0.42
r25 8 16 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.6 $Y=0.93 $X2=1.5
+ $Y2=0.93
r26 7 9 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.79 $Y=0.93
+ $X2=2.885 $Y2=0.845
r27 7 8 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.79 $Y=0.93 $X2=1.6
+ $Y2=0.93
r28 2 11 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.745
+ $Y=0.235 $X2=2.885 $Y2=0.42
r29 1 14 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=1.365
+ $Y=0.245 $X2=1.505 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r53 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r54 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r55 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r56 24 28 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r57 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 21 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r59 21 25 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=0.24
+ $Y2=0
r60 21 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r61 19 31 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.15 $Y=0 $X2=3.12
+ $Y2=0
r62 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=0 $X2=3.315
+ $Y2=0
r63 18 34 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.48 $Y=0 $X2=4.08
+ $Y2=0
r64 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.48 $Y=0 $X2=3.315
+ $Y2=0
r65 16 28 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.29 $Y=0 $X2=2.16
+ $Y2=0
r66 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=0 $X2=2.455
+ $Y2=0
r67 15 31 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.62 $Y=0 $X2=3.12
+ $Y2=0
r68 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=0 $X2=2.455
+ $Y2=0
r69 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0
r70 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0.38
r71 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=0.085
+ $X2=2.455 $Y2=0
r72 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.455 $Y=0.085
+ $X2=2.455 $Y2=0.55
r73 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.175
+ $Y=0.235 $X2=3.315 $Y2=0.38
r74 1 9 182 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_NDIFF $count=1 $X=2.33
+ $Y=0.235 $X2=2.455 $Y2=0.55
.ends

