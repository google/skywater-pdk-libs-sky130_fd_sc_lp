* File: sky130_fd_sc_lp__dlxtp_lp.pex.spice
* Created: Fri Aug 28 10:29:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%GATE 3 7 11 15 17 18 22
r39 17 18 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.74 $Y=1.645
+ $X2=0.74 $Y2=2.035
r40 17 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.74
+ $Y=1.645 $X2=0.74 $Y2=1.645
r41 13 22 92.2311 $w=2.7e-07 $l=5.94559e-07 $layer=POLY_cond $X=0.885 $Y=2.15
+ $X2=0.69 $Y2=1.645
r42 13 15 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.885 $Y=2.15
+ $X2=0.885 $Y2=2.67
r43 9 22 31.5348 $w=2.7e-07 $l=2.33345e-07 $layer=POLY_cond $X=0.855 $Y=1.48
+ $X2=0.69 $Y2=1.645
r44 9 11 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.855 $Y=1.48
+ $X2=0.855 $Y2=0.72
r45 5 22 92.2311 $w=2.7e-07 $l=5.94559e-07 $layer=POLY_cond $X=0.495 $Y=2.15
+ $X2=0.69 $Y2=1.645
r46 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.495 $Y=2.15
+ $X2=0.495 $Y2=2.67
r47 1 22 31.5348 $w=2.7e-07 $l=1.95e-07 $layer=POLY_cond $X=0.495 $Y=1.645
+ $X2=0.69 $Y2=1.645
r48 1 3 389.702 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.495 $Y=1.645
+ $X2=0.495 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%D 3 7 11 15 17 23 24
c46 3 0 1.39673e-19 $X=1.315 $Y=0.72
r47 22 24 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.435 $Y=1.985
+ $X2=1.675 $Y2=1.985
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.435
+ $Y=1.985 $X2=1.435 $Y2=1.985
r49 19 22 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.315 $Y=1.985
+ $X2=1.435 $Y2=1.985
r50 17 23 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.435 $Y2=1.985
r51 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=2.15
+ $X2=1.675 $Y2=1.985
r52 13 15 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.675 $Y=2.15
+ $X2=1.675 $Y2=2.67
r53 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.82
+ $X2=1.675 $Y2=1.985
r54 9 11 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=1.675 $Y=1.82
+ $X2=1.675 $Y2=0.72
r55 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.315 $Y=2.15
+ $X2=1.315 $Y2=1.985
r56 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.315 $Y=2.15
+ $X2=1.315 $Y2=2.67
r57 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.315 $Y=1.82
+ $X2=1.315 $Y2=1.985
r58 1 3 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=1.315 $Y=1.82
+ $X2=1.315 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%A_27_102# 1 2 8 11 13 17 21 25 29 31 35 39
+ 41 44 48 50 52 54 56 57 61 68 74 78
c154 78 0 3.48291e-20 $X=4.105 $Y=1.72
c155 68 0 3.48291e-20 $X=4.105 $Y=1.67
c156 52 0 1.39673e-19 $X=2.98 $Y=1.51
c157 29 0 1.30072e-19 $X=4.045 $Y=2.775
c158 21 0 1.98648e-19 $X=3.065 $Y=2.775
r159 74 75 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.145 $Y=1.5
+ $X2=3.145 $Y2=1.425
r160 72 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.81
+ $X2=4.105 $Y2=1.975
r161 72 78 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.105 $Y=1.81
+ $X2=4.105 $Y2=1.72
r162 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=1.81 $X2=4.105 $Y2=1.81
r163 68 71 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=4.105 $Y=1.67
+ $X2=4.105 $Y2=1.81
r164 65 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.59
+ $X2=3.145 $Y2=1.755
r165 65 74 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.145 $Y=1.59
+ $X2=3.145 $Y2=1.5
r166 64 66 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.145 $Y=1.59
+ $X2=3.145 $Y2=1.67
r167 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.145
+ $Y=1.59 $X2=3.145 $Y2=1.59
r168 61 64 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.145 $Y=1.51
+ $X2=3.145 $Y2=1.59
r169 57 59 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.46 $Y=1.215
+ $X2=1.46 $Y2=1.51
r170 55 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=1.67
+ $X2=3.145 $Y2=1.67
r171 54 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.94 $Y=1.67
+ $X2=4.105 $Y2=1.67
r172 54 55 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.94 $Y=1.67
+ $X2=3.31 $Y2=1.67
r173 53 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=1.51
+ $X2=1.46 $Y2=1.51
r174 52 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.98 $Y=1.51
+ $X2=3.145 $Y2=1.51
r175 52 53 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=2.98 $Y=1.51
+ $X2=1.545 $Y2=1.51
r176 51 56 3.3199 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.215
+ $X2=0.28 $Y2=1.215
r177 50 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=1.215
+ $X2=1.46 $Y2=1.215
r178 50 51 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.375 $Y=1.215
+ $X2=0.445 $Y2=1.215
r179 46 56 3.24686 $w=2.9e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.24 $Y=1.3
+ $X2=0.28 $Y2=1.215
r180 46 48 55.0868 $w=2.48e-07 $l=1.195e-06 $layer=LI1_cond $X=0.24 $Y=1.3
+ $X2=0.24 $Y2=2.495
r181 42 56 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=1.13
+ $X2=0.28 $Y2=1.215
r182 42 44 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=1.13
+ $X2=0.28 $Y2=0.72
r183 37 39 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.675 $Y=1.11
+ $X2=2.845 $Y2=1.11
r184 33 35 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=4.835 $Y=1.645
+ $X2=4.835 $Y2=0.445
r185 32 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=1.72
+ $X2=4.105 $Y2=1.72
r186 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.76 $Y=1.72
+ $X2=4.835 $Y2=1.645
r187 31 32 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=4.76 $Y=1.72
+ $X2=4.27 $Y2=1.72
r188 29 81 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.045 $Y=2.775
+ $X2=4.045 $Y2=1.975
r189 25 75 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.235 $Y=0.445
+ $X2=3.235 $Y2=1.425
r190 21 77 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.065 $Y=2.775
+ $X2=3.065 $Y2=1.755
r191 15 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.845 $Y=1.035
+ $X2=2.845 $Y2=1.11
r192 15 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.845 $Y=1.035
+ $X2=2.845 $Y2=0.445
r193 14 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.75 $Y=1.5
+ $X2=2.675 $Y2=1.5
r194 13 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.98 $Y=1.5
+ $X2=3.145 $Y2=1.5
r195 13 14 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.98 $Y=1.5
+ $X2=2.75 $Y2=1.5
r196 9 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.675 $Y=1.575
+ $X2=2.675 $Y2=1.5
r197 9 11 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=2.675 $Y=1.575
+ $X2=2.675 $Y2=2.775
r198 8 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.675 $Y=1.425
+ $X2=2.675 $Y2=1.5
r199 7 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.675 $Y=1.185
+ $X2=2.675 $Y2=1.11
r200 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.675 $Y=1.185
+ $X2=2.675 $Y2=1.425
r201 2 48 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.35 $X2=0.28 $Y2=2.495
r202 1 44 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.51 $X2=0.28 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%A_350_102# 1 2 11 15 19 23 27 28 29 30 31
+ 32 36 38 45 50
c101 38 0 1.08596e-19 $X=3.715 $Y=1.16
c102 36 0 3.48291e-20 $X=3.565 $Y=2.13
c103 32 0 3.48291e-20 $X=3.565 $Y=2.05
r104 42 50 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.715 $Y=1.24
+ $X2=3.875 $Y2=1.24
r105 42 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.715 $Y=1.24
+ $X2=3.625 $Y2=1.24
r106 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.715
+ $Y=1.24 $X2=3.715 $Y2=1.24
r107 38 41 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.715 $Y=1.16
+ $X2=3.715 $Y2=1.24
r108 36 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=2.13
+ $X2=3.565 $Y2=2.295
r109 36 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=2.13
+ $X2=3.565 $Y2=1.965
r110 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.565
+ $Y=2.13 $X2=3.565 $Y2=2.13
r111 32 35 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.565 $Y=2.05
+ $X2=3.565 $Y2=2.13
r112 29 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=2.05
+ $X2=3.565 $Y2=2.05
r113 29 30 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=3.4 $Y=2.05
+ $X2=2.055 $Y2=2.05
r114 27 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=1.16
+ $X2=3.715 $Y2=1.16
r115 27 28 97.5348 $w=1.68e-07 $l=1.495e-06 $layer=LI1_cond $X=3.55 $Y=1.16
+ $X2=2.055 $Y2=1.16
r116 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=2.135
+ $X2=2.055 $Y2=2.05
r117 25 31 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.97 $Y=2.135
+ $X2=1.97 $Y2=2.33
r118 23 31 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=2.495
+ $X2=1.89 $Y2=2.33
r119 17 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.89 $Y=1.075
+ $X2=2.055 $Y2=1.16
r120 17 19 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.89 $Y=1.075
+ $X2=1.89 $Y2=0.72
r121 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.875 $Y=1.075
+ $X2=3.875 $Y2=1.24
r122 13 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.875 $Y=1.075
+ $X2=3.875 $Y2=0.445
r123 11 46 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.655 $Y=2.775
+ $X2=3.655 $Y2=2.295
r124 7 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.625 $Y=1.405
+ $X2=3.625 $Y2=1.24
r125 7 45 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.625 $Y=1.405
+ $X2=3.625 $Y2=1.965
r126 2 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.75
+ $Y=2.35 $X2=1.89 $Y2=2.495
r127 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.51 $X2=1.89 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%A_463_491# 1 2 9 13 15 20 22 23 24 25 29 30
+ 33 34 35
c112 34 0 8.98036e-20 $X=4.73 $Y=2.35
c113 33 0 1.30072e-19 $X=4.73 $Y=2.35
c114 30 0 1.08596e-19 $X=4.355 $Y=1.02
c115 23 0 1.98648e-19 $X=2.625 $Y=2.56
r116 34 41 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.73 $Y=2.35
+ $X2=4.59 $Y2=2.35
r117 33 35 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=4.672 $Y=2.35
+ $X2=4.672 $Y2=2.185
r118 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.73
+ $Y=2.35 $X2=4.73 $Y2=2.35
r119 30 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.02
+ $X2=4.355 $Y2=0.855
r120 29 31 5.90323 $w=3.72e-07 $l=1.8e-07 $layer=LI1_cond $X=4.355 $Y=0.955
+ $X2=4.535 $Y2=0.955
r121 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.355
+ $Y=1.02 $X2=4.355 $Y2=1.02
r122 26 31 5.3395 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.535 $Y=1.185
+ $X2=4.535 $Y2=0.955
r123 26 35 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=4.535 $Y=1.185
+ $X2=4.535 $Y2=2.185
r124 24 29 11.8335 $w=3.72e-07 $l=3.14245e-07 $layer=LI1_cond $X=4.105 $Y=0.81
+ $X2=4.355 $Y2=0.955
r125 24 25 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=4.105 $Y=0.81
+ $X2=2.795 $Y2=0.81
r126 22 33 5.4385 $w=4.43e-07 $l=2.1e-07 $layer=LI1_cond $X=4.672 $Y=2.56
+ $X2=4.672 $Y2=2.35
r127 22 23 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=4.45 $Y=2.56
+ $X2=2.625 $Y2=2.56
r128 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.63 $Y=0.725
+ $X2=2.795 $Y2=0.81
r129 18 20 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.63 $Y=0.725
+ $X2=2.63 $Y2=0.47
r130 15 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.46 $Y=2.645
+ $X2=2.625 $Y2=2.56
r131 15 17 3.88182 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=2.46 $Y=2.645
+ $X2=2.46 $Y2=2.75
r132 11 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=2.515
+ $X2=4.59 $Y2=2.35
r133 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.59 $Y=2.515
+ $X2=4.59 $Y2=2.885
r134 9 39 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.265 $Y=0.445
+ $X2=4.265 $Y2=0.855
r135 2 17 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=2.455 $X2=2.46 $Y2=2.75
r136 1 20 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.63 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%A_1027_407# 1 2 9 13 19 23 27 31 33 34 35
+ 39 42 45 51 54 58 60 61 68
c110 61 0 1.43975e-19 $X=6.52 $Y=1.47
c111 34 0 3.8192e-20 $X=5.217 $Y=2.185
r112 58 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.315 $Y=1.09
+ $X2=5.315 $Y2=1.255
r113 58 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.315 $Y=1.09
+ $X2=5.315 $Y2=0.925
r114 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.315
+ $Y=1.09 $X2=5.315 $Y2=1.09
r115 54 57 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.315 $Y=1.01
+ $X2=5.315 $Y2=1.09
r116 52 68 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=7.36 $Y=1.47
+ $X2=7.655 $Y2=1.47
r117 52 65 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.36 $Y=1.47
+ $X2=7.295 $Y2=1.47
r118 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.36
+ $Y=1.47 $X2=7.36 $Y2=1.47
r119 49 61 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.685 $Y=1.47
+ $X2=6.52 $Y2=1.47
r120 49 51 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.685 $Y=1.47
+ $X2=7.36 $Y2=1.47
r121 45 47 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=6.52 $Y=1.98
+ $X2=6.52 $Y2=2.9
r122 43 61 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=1.635
+ $X2=6.52 $Y2=1.47
r123 43 45 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.52 $Y=1.635
+ $X2=6.52 $Y2=1.98
r124 42 61 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=1.305
+ $X2=6.52 $Y2=1.47
r125 41 60 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.095
+ $X2=6.52 $Y2=1.01
r126 41 42 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.52 $Y=1.095
+ $X2=6.52 $Y2=1.305
r127 37 60 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.925
+ $X2=6.52 $Y2=1.01
r128 37 39 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.52 $Y=0.925
+ $X2=6.52 $Y2=0.43
r129 36 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.48 $Y=1.01
+ $X2=5.315 $Y2=1.01
r130 35 60 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.355 $Y=1.01
+ $X2=6.52 $Y2=1.01
r131 35 36 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=6.355 $Y=1.01
+ $X2=5.48 $Y2=1.01
r132 33 34 65.3429 $w=1.65e-07 $l=1.5e-07 $layer=POLY_cond $X=5.217 $Y=2.035
+ $X2=5.217 $Y2=2.185
r133 33 64 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.225 $Y=2.035
+ $X2=5.225 $Y2=1.255
r134 29 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.635
+ $X2=7.655 $Y2=1.47
r135 29 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.655 $Y=1.635
+ $X2=7.655 $Y2=2.465
r136 25 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.305
+ $X2=7.655 $Y2=1.47
r137 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.655 $Y=1.305
+ $X2=7.655 $Y2=0.685
r138 21 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.295 $Y=1.635
+ $X2=7.295 $Y2=1.47
r139 21 23 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.295 $Y=1.635
+ $X2=7.295 $Y2=2.465
r140 17 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.295 $Y=1.305
+ $X2=7.295 $Y2=1.47
r141 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.295 $Y=1.305
+ $X2=7.295 $Y2=0.685
r142 13 63 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.225 $Y=0.445
+ $X2=5.225 $Y2=0.925
r143 9 34 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=5.21 $Y=2.885 $X2=5.21
+ $Y2=2.185
r144 2 47 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=1.835 $X2=6.52 $Y2=2.9
r145 2 45 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=1.835 $X2=6.52 $Y2=1.98
r146 1 39 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=6.38
+ $Y=0.235 $X2=6.52 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%A_824_491# 1 2 9 13 17 21 23 28 30 31 32 34
+ 40 49
c101 32 0 1.27996e-19 $X=5.245 $Y=1.52
c102 13 0 1.43975e-19 $X=5.945 $Y=2.465
r103 45 47 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.915 $Y=1.44
+ $X2=5.945 $Y2=1.44
r104 41 49 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=6.005 $Y=1.44
+ $X2=6.305 $Y2=1.44
r105 41 47 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.005 $Y=1.44
+ $X2=5.945 $Y2=1.44
r106 40 43 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.005 $Y=1.44
+ $X2=6.005 $Y2=1.52
r107 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.005
+ $Y=1.44 $X2=6.005 $Y2=1.44
r108 36 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.885 $Y=1.52
+ $X2=5.16 $Y2=1.52
r109 32 38 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.245 $Y=1.52
+ $X2=5.16 $Y2=1.52
r110 31 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.84 $Y=1.52
+ $X2=6.005 $Y2=1.52
r111 31 32 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.84 $Y=1.52
+ $X2=5.245 $Y2=1.52
r112 29 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=1.605
+ $X2=5.16 $Y2=1.52
r113 29 30 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=5.16 $Y=1.605
+ $X2=5.16 $Y2=2.825
r114 28 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=1.435
+ $X2=4.885 $Y2=1.52
r115 27 34 10.0093 $w=3.23e-07 $l=3.52916e-07 $layer=LI1_cond $X=4.885 $Y=0.675
+ $X2=4.62 $Y2=0.47
r116 27 28 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.885 $Y=0.675
+ $X2=4.885 $Y2=1.435
r117 23 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.075 $Y=2.93
+ $X2=5.16 $Y2=2.825
r118 23 25 43.0433 $w=2.08e-07 $l=8.15e-07 $layer=LI1_cond $X=5.075 $Y=2.93
+ $X2=4.26 $Y2=2.93
r119 19 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.605
+ $X2=6.305 $Y2=1.44
r120 19 21 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.305 $Y=1.605
+ $X2=6.305 $Y2=2.465
r121 15 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.275
+ $X2=6.305 $Y2=1.44
r122 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.305 $Y=1.275
+ $X2=6.305 $Y2=0.655
r123 11 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.945 $Y=1.605
+ $X2=5.945 $Y2=1.44
r124 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.945 $Y=1.605
+ $X2=5.945 $Y2=2.465
r125 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.275
+ $X2=5.915 $Y2=1.44
r126 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.915 $Y=1.275
+ $X2=5.915 $Y2=0.655
r127 2 25 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=2.455 $X2=4.26 $Y2=2.93
r128 1 34 182 $w=1.7e-07 $l=3.79737e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=0.235 $X2=4.62 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%VPWR 1 2 3 4 15 19 23 29 34 35 37 38 39 41
+ 56 62 63 66 69
r95 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r96 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r97 63 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=6.96 $Y2=3.33
r98 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r99 60 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=3.33
+ $X2=7.08 $Y2=3.33
r100 60 62 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.245 $Y=3.33
+ $X2=7.92 $Y2=3.33
r101 59 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r102 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r103 56 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=3.33
+ $X2=7.08 $Y2=3.33
r104 56 58 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=6.915 $Y=3.33
+ $X2=6 $Y2=3.33
r105 55 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r106 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r107 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r109 49 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r110 49 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 48 49 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.1 $Y2=3.33
r113 46 48 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 44 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=1.1 $Y2=3.33
r117 41 43 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 39 55 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 39 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r120 37 54 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.565 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=3.33
+ $X2=5.73 $Y2=3.33
r122 36 58 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.895 $Y=3.33
+ $X2=6 $Y2=3.33
r123 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.895 $Y=3.33
+ $X2=5.73 $Y2=3.33
r124 34 48 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.36 $Y2=3.33
r126 33 51 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=3.6 $Y2=3.33
r127 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=3.36 $Y2=3.33
r128 29 32 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=7.08 $Y=1.98
+ $X2=7.08 $Y2=2.95
r129 27 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=3.245
+ $X2=7.08 $Y2=3.33
r130 27 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.08 $Y=3.245
+ $X2=7.08 $Y2=2.95
r131 23 26 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=5.73 $Y=1.98
+ $X2=5.73 $Y2=2.95
r132 21 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.73 $Y=3.245
+ $X2=5.73 $Y2=3.33
r133 21 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.73 $Y=3.245
+ $X2=5.73 $Y2=2.95
r134 17 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=3.245
+ $X2=3.36 $Y2=3.33
r135 17 19 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.36 $Y=3.245
+ $X2=3.36 $Y2=2.99
r136 13 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=3.245 $X2=1.1
+ $Y2=3.33
r137 13 15 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=1.1 $Y=3.245
+ $X2=1.1 $Y2=2.495
r138 4 32 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=6.935
+ $Y=1.835 $X2=7.08 $Y2=2.95
r139 4 29 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.935
+ $Y=1.835 $X2=7.08 $Y2=1.98
r140 3 26 600 $w=1.7e-07 $l=5.66039e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=2.675 $X2=5.73 $Y2=2.95
r141 3 23 300 $w=1.7e-07 $l=8.90112e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=2.675 $X2=5.73 $Y2=1.98
r142 2 19 600 $w=1.7e-07 $l=6.35551e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=2.455 $X2=3.36 $Y2=2.99
r143 1 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.96
+ $Y=2.35 $X2=1.1 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%Q 1 2 7 8 9 10 11 12 13 22
r15 13 40 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=7.87 $Y=2.775
+ $X2=7.87 $Y2=2.9
r16 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.87 $Y=2.405
+ $X2=7.87 $Y2=2.775
r17 11 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.87 $Y=1.98
+ $X2=7.87 $Y2=2.405
r18 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=7.87 $Y=1.665
+ $X2=7.87 $Y2=1.98
r19 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.87 $Y=1.295
+ $X2=7.87 $Y2=1.665
r20 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.87 $Y=0.925 $X2=7.87
+ $Y2=1.295
r21 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.87 $Y=0.555 $X2=7.87
+ $Y2=0.925
r22 7 22 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=7.87 $Y=0.555
+ $X2=7.87 $Y2=0.43
r23 2 40 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.835 $X2=7.87 $Y2=2.9
r24 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.835 $X2=7.87 $Y2=1.98
r25 1 22 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=7.73
+ $Y=0.265 $X2=7.87 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP%VGND 1 2 3 4 15 19 23 27 29 31 36 41 46 53
+ 54 57 60 63 66
r94 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r95 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r96 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r97 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r98 54 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=6.96
+ $Y2=0
r99 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r100 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=0 $X2=7.08
+ $Y2=0
r101 51 53 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.245 $Y=0
+ $X2=7.92 $Y2=0
r102 50 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r103 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r104 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r105 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.445
+ $Y2=0
r106 47 49 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=6
+ $Y2=0
r107 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=7.08
+ $Y2=0
r108 46 49 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6
+ $Y2=0
r109 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r110 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r111 42 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.45
+ $Y2=0
r112 42 44 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=3.615 $Y=0
+ $X2=5.04 $Y2=0
r113 41 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.28 $Y=0 $X2=5.445
+ $Y2=0
r114 41 44 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.28 $Y=0 $X2=5.04
+ $Y2=0
r115 40 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r116 40 58 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=1.2
+ $Y2=0
r117 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r118 37 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r119 37 39 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=3.12 $Y2=0
r120 36 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=0 $X2=3.45
+ $Y2=0
r121 36 39 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=0
+ $X2=3.12 $Y2=0
r122 34 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r123 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r124 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r125 31 33 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r126 29 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r127 29 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r128 25 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0
r129 25 27 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0.41
r130 21 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=0.085
+ $X2=5.445 $Y2=0
r131 21 23 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.445 $Y=0.085
+ $X2=5.445 $Y2=0.445
r132 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=0.085
+ $X2=3.45 $Y2=0
r133 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.45 $Y=0.085
+ $X2=3.45 $Y2=0.38
r134 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r135 13 15 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.72
r136 4 27 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.935
+ $Y=0.265 $X2=7.08 $Y2=0.41
r137 3 23 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.3
+ $Y=0.235 $X2=5.445 $Y2=0.445
r138 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.31
+ $Y=0.235 $X2=3.45 $Y2=0.38
r139 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.51 $X2=1.07 $Y2=0.72
.ends

