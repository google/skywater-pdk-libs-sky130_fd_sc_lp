* NGSPICE file created from sky130_fd_sc_lp__dfsbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
M1000 a_129_179# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=2.6113e+12p ps=2.327e+07u
M1001 VPWR a_2227_367# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1002 a_129_179# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.9105e+12p ps=1.806e+07u
M1003 a_1173_125# a_593_125# VGND VNB nshort w=640000u l=150000u
+  ad=4.875e+11p pd=4.51e+06u as=0p ps=0u
M1004 VPWR a_1360_451# Q_N VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1005 a_1360_451# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=3.906e+11p pd=3.83e+06u as=0p ps=0u
M1006 VPWR a_129_179# a_191_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1007 VGND a_1360_451# a_1533_258# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 a_507_125# D VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1009 a_1360_451# a_129_179# a_1288_451# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1010 a_1288_451# a_593_125# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1677_91# a_1533_258# a_1280_159# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.226e+11p ps=2.74e+06u
M1012 Q a_2227_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1013 VPWR a_1533_258# a_1468_451# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.365e+11p ps=1.49e+06u
M1014 VGND SET_B a_1677_91# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q_N a_1360_451# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 Q a_2227_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR SET_B a_721_99# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=4.053e+11p ps=2.77e+06u
M1018 a_2227_367# a_1360_451# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1019 a_721_99# a_593_125# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1360_451# a_129_179# a_1280_159# VNB nshort w=420000u l=150000u
+  ad=2.158e+11p pd=2.03e+06u as=0p ps=0u
M1021 a_679_125# a_191_21# a_593_125# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1022 VGND SET_B a_996_169# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1023 a_996_169# a_593_125# a_721_99# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1024 VPWR a_1360_451# a_1533_258# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1025 VGND a_721_99# a_679_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1173_125# a_191_21# a_1360_451# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_2227_367# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_701_535# a_129_179# a_593_125# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.344e+11p ps=1.48e+06u
M1029 a_1468_451# a_191_21# a_1360_451# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_1360_451# Q_N VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_721_99# a_701_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_507_125# D VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1033 a_593_125# a_129_179# a_507_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2227_367# a_1360_451# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1035 Q_N a_1360_451# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_129_179# a_191_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1037 a_593_125# a_191_21# a_507_125# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

