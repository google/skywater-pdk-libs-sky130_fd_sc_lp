* NGSPICE file created from sky130_fd_sc_lp__nor4bb_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor4bb_lp A B C_N D_N VGND VNB VPB VPWR Y
M1000 a_245_409# a_430_21# Y VPB phighvt w=1e+06u l=250000u
+  ad=5.7e+11p pd=5.14e+06u as=2.85e+11p ps=2.57e+06u
M1001 VGND C_N a_144_47# VNB nshort w=420000u l=150000u
+  ad=4.242e+11p pd=4.54e+06u as=8.82e+10p ps=1.26e+06u
M1002 a_624_47# B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1003 a_788_409# B a_352_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=5.7e+11p ps=5.14e+06u
M1004 Y B a_624_47# VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=0p ps=0u
M1005 VPWR C_N a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=6.05e+11p pd=5.21e+06u as=2.85e+11p ps=2.57e+06u
M1006 a_430_21# D_N VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1007 a_144_47# C_N a_27_409# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1008 a_302_47# a_27_409# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 Y a_27_409# a_302_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_782_47# A Y VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1011 VPWR A a_788_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A a_782_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_460_47# a_430_21# Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1014 VGND a_430_21# a_460_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_980_47# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1016 a_352_409# a_27_409# a_245_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_430_21# D_N a_980_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends

