# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdlclkp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdlclkp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.035000 0.555000 1.705000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.075000 0.265000 8.515000 0.595000 ;
        RECT 8.115000 2.060000 8.515000 3.065000 ;
        RECT 8.285000 0.595000 8.515000 2.060000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.390000 1.570000 2.150000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.580000 5.655000 2.150000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.855000 ;
      RECT 0.445000  1.885000 0.905000 2.615000 ;
      RECT 0.445000  2.615000 2.225000 2.785000 ;
      RECT 0.445000  2.785000 0.775000 2.900000 ;
      RECT 0.735000  0.485000 1.265000 1.040000 ;
      RECT 0.735000  1.040000 2.405000 1.210000 ;
      RECT 0.735000  1.210000 0.905000 1.885000 ;
      RECT 1.545000  2.965000 1.875000 3.245000 ;
      RECT 1.725000  0.085000 2.055000 0.860000 ;
      RECT 1.780000  1.390000 2.110000 2.265000 ;
      RECT 1.780000  2.265000 2.575000 2.435000 ;
      RECT 2.055000  2.785000 3.265000 3.045000 ;
      RECT 2.235000  0.265000 3.505000 0.435000 ;
      RECT 2.235000  0.435000 2.405000 1.040000 ;
      RECT 2.290000  1.390000 3.200000 1.720000 ;
      RECT 2.290000  1.720000 2.620000 2.085000 ;
      RECT 2.405000  2.435000 4.145000 2.605000 ;
      RECT 2.595000  0.615000 2.970000 0.945000 ;
      RECT 2.800000  0.945000 2.970000 1.390000 ;
      RECT 3.175000  0.435000 3.505000 0.675000 ;
      RECT 3.380000  0.880000 5.265000 1.050000 ;
      RECT 3.380000  1.050000 3.550000 2.005000 ;
      RECT 3.380000  2.005000 3.795000 2.255000 ;
      RECT 3.685000  0.265000 3.935000 0.880000 ;
      RECT 3.730000  1.495000 4.145000 1.825000 ;
      RECT 3.975000  1.230000 6.045000 1.400000 ;
      RECT 3.975000  1.400000 4.145000 1.495000 ;
      RECT 3.975000  1.825000 4.145000 2.435000 ;
      RECT 4.325000  1.580000 4.655000 2.330000 ;
      RECT 4.325000  2.330000 5.420000 2.490000 ;
      RECT 4.325000  2.490000 7.925000 2.500000 ;
      RECT 4.425000  0.085000 4.755000 0.675000 ;
      RECT 4.525000  2.680000 4.855000 3.245000 ;
      RECT 4.935000  0.765000 5.265000 0.880000 ;
      RECT 5.090000  2.500000 7.925000 2.660000 ;
      RECT 5.090000  2.660000 5.420000 3.045000 ;
      RECT 5.445000  0.265000 5.775000 0.505000 ;
      RECT 5.445000  0.505000 6.395000 0.675000 ;
      RECT 5.715000  0.940000 6.045000 1.230000 ;
      RECT 5.835000  1.400000 6.045000 2.060000 ;
      RECT 5.835000  2.060000 6.165000 2.310000 ;
      RECT 6.225000  0.675000 6.395000 1.580000 ;
      RECT 6.225000  1.580000 6.515000 1.750000 ;
      RECT 6.345000  1.750000 6.515000 2.490000 ;
      RECT 6.365000  2.840000 6.695000 3.245000 ;
      RECT 6.585000  0.085000 6.835000 1.400000 ;
      RECT 6.895000  2.060000 7.575000 2.230000 ;
      RECT 6.895000  2.230000 7.225000 2.310000 ;
      RECT 7.265000  0.085000 7.595000 0.680000 ;
      RECT 7.325000  0.935000 8.105000 1.105000 ;
      RECT 7.325000  1.105000 7.575000 2.060000 ;
      RECT 7.505000  2.840000 7.835000 3.245000 ;
      RECT 7.755000  1.315000 8.085000 1.645000 ;
      RECT 7.755000  1.645000 7.925000 2.490000 ;
      RECT 7.775000  0.775000 8.105000 0.935000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_lp__sdlclkp_lp
