* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 X a_36_67# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_36_67# C1 a_119_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_235_367# B2 a_36_67# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_36_67# A2 a_461_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_461_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_119_67# B1 a_205_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_36_67# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_205_67# B2 a_119_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND A2 a_205_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR a_36_67# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR B1 a_235_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 X a_36_67# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_205_67# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VGND a_36_67# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
