* File: sky130_fd_sc_lp__o21ba_1.pex.spice
* Created: Wed Sep  2 10:16:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BA_1%A_84_28# 1 2 7 9 12 15 16 17 19 20 21 25 26
+ 27 28 30 36 43
r83 34 43 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=0.65 $Y=1.385
+ $X2=0.695 $Y2=1.385
r84 34 40 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.65 $Y=1.385
+ $X2=0.495 $Y2=1.385
r85 33 36 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.65 $Y=1.385 $X2=0.85
+ $Y2=1.385
r86 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.65
+ $Y=1.385 $X2=0.65 $Y2=1.385
r87 28 39 2.8525 $w=2.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.66 $Y=2.1 $X2=2.66
+ $Y2=2.012
r88 28 30 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.66 $Y=2.1
+ $X2=2.66 $Y2=2.435
r89 26 39 4.376 $w=1.75e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=2.012
+ $X2=2.66 $Y2=2.012
r90 26 27 13.626 $w=1.73e-07 $l=2.15e-07 $layer=LI1_cond $X=2.525 $Y=2.012
+ $X2=2.31 $Y2=2.012
r91 23 27 7.00809 $w=1.75e-07 $l=1.55531e-07 $layer=LI1_cond $X=2.192 $Y=1.925
+ $X2=2.31 $Y2=2.012
r92 23 25 73.315 $w=2.33e-07 $l=1.495e-06 $layer=LI1_cond $X=2.192 $Y=1.925
+ $X2=2.192 $Y2=0.43
r93 22 25 0.245201 $w=2.33e-07 $l=5e-09 $layer=LI1_cond $X=2.192 $Y=0.425
+ $X2=2.192 $Y2=0.43
r94 20 22 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.075 $Y=0.34
+ $X2=2.192 $Y2=0.425
r95 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.075 $Y=0.34
+ $X2=1.305 $Y2=0.34
r96 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.305 $Y2=0.34
r97 18 19 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.22 $Y2=0.87
r98 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.135 $Y=0.955
+ $X2=1.22 $Y2=0.87
r99 16 17 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.135 $Y=0.955
+ $X2=0.935 $Y2=0.955
r100 15 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=1.22
+ $X2=0.85 $Y2=1.385
r101 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.85 $Y=1.04
+ $X2=0.935 $Y2=0.955
r102 14 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.85 $Y=1.04
+ $X2=0.85 $Y2=1.22
r103 10 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.695 $Y=1.55
+ $X2=0.695 $Y2=1.385
r104 10 12 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=0.695 $Y=1.55
+ $X2=0.695 $Y2=2.465
r105 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=1.385
r106 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=0.69
r107 2 39 600 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.835 $X2=2.63 $Y2=2.01
r108 2 30 300 $w=1.7e-07 $l=6.75278e-07 $layer=licon1_PDIFF $count=2 $X=2.47
+ $Y=1.835 $X2=2.63 $Y2=2.435
r109 1 25 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=2.055
+ $Y=0.255 $X2=2.18 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_1%B1_N 3 6 8 9 13 15
r33 13 16 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=1.385
+ $X2=1.23 $Y2=1.55
r34 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=1.385
+ $X2=1.23 $Y2=1.22
r35 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.385 $X2=1.22 $Y2=1.385
r36 9 14 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=1.205 $Y=1.665
+ $X2=1.205 $Y2=1.385
r37 8 14 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=1.205 $Y=1.295
+ $X2=1.205 $Y2=1.385
r38 6 16 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.33 $Y=2.045
+ $X2=1.33 $Y2=1.55
r39 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.33 $Y=0.9 $X2=1.33
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_1%A_281_138# 1 2 7 9 12 14 15 18 23 24 27
r37 27 29 5.82291 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.69 $Y=1.385
+ $X2=1.69 $Y2=1.55
r38 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.385 $X2=1.81 $Y2=1.385
r39 24 29 15.4345 $w=2.78e-07 $l=3.75e-07 $layer=LI1_cond $X=1.615 $Y=1.925
+ $X2=1.615 $Y2=1.55
r40 23 24 4.48843 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.59 $Y=2.045
+ $X2=1.59 $Y2=1.925
r41 16 27 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=1.69 $Y=1.335 $X2=1.69
+ $Y2=1.385
r42 16 18 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=1.335
+ $X2=1.69 $Y2=0.965
r43 14 28 89.1793 $w=3.3e-07 $l=5.1e-07 $layer=POLY_cond $X=2.32 $Y=1.385
+ $X2=1.81 $Y2=1.385
r44 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.32 $Y=1.385
+ $X2=2.395 $Y2=1.385
r45 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.55
+ $X2=2.395 $Y2=1.385
r46 10 12 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=2.395 $Y=1.55
+ $X2=2.395 $Y2=2.465
r47 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.22
+ $X2=2.395 $Y2=1.385
r48 7 9 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.395 $Y=1.22
+ $X2=2.395 $Y2=0.675
r49 2 23 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=1.835 $X2=1.59 $Y2=2.045
r50 1 18 182 $w=1.7e-07 $l=3.78153e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.69 $X2=1.65 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_1%A2 3 7 9 10 14
c35 14 0 1.25093e-19 $X=2.875 $Y=1.51
c36 7 0 5.33748e-20 $X=2.845 $Y=2.465
r37 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.51
+ $X2=2.875 $Y2=1.675
r38 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.51
+ $X2=2.875 $Y2=1.345
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.875
+ $Y=1.51 $X2=2.875 $Y2=1.51
r40 10 15 8.68765 $w=3.23e-07 $l=2.45e-07 $layer=LI1_cond $X=3.12 $Y=1.587
+ $X2=2.875 $Y2=1.587
r41 9 15 8.33305 $w=3.23e-07 $l=2.35e-07 $layer=LI1_cond $X=2.64 $Y=1.587
+ $X2=2.875 $Y2=1.587
r42 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.845 $Y=2.465
+ $X2=2.845 $Y2=1.675
r43 3 16 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.825 $Y=0.675
+ $X2=2.825 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_1%A1 3 7 9 14 15
c26 15 0 5.33748e-20 $X=3.55 $Y=1.46
r27 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.46 $X2=3.55 $Y2=1.46
r28 11 14 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=3.355 $Y=1.46
+ $X2=3.55 $Y2=1.46
r29 9 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.46
r30 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.625
+ $X2=3.355 $Y2=1.46
r31 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.355 $Y=1.625
+ $X2=3.355 $Y2=2.465
r32 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.295
+ $X2=3.355 $Y2=1.46
r33 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.355 $Y=1.295
+ $X2=3.355 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_1%X 1 2 7 8 9 10 11 12 13 24 44 48
r17 44 45 5.81366 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.33 $Y=1.98
+ $X2=0.33 $Y2=1.815
r18 34 48 0.610244 $w=4.88e-07 $l=2.5e-08 $layer=LI1_cond $X=0.33 $Y=2.06
+ $X2=0.33 $Y2=2.035
r19 13 41 3.29532 $w=4.88e-07 $l=1.35e-07 $layer=LI1_cond $X=0.33 $Y=2.775
+ $X2=0.33 $Y2=2.91
r20 12 13 9.03161 $w=4.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.33 $Y=2.405
+ $X2=0.33 $Y2=2.775
r21 11 48 0.732293 $w=4.88e-07 $l=3e-08 $layer=LI1_cond $X=0.33 $Y=2.005
+ $X2=0.33 $Y2=2.035
r22 11 44 0.610244 $w=4.88e-07 $l=2.5e-08 $layer=LI1_cond $X=0.33 $Y=2.005
+ $X2=0.33 $Y2=1.98
r23 11 12 7.68908 $w=4.88e-07 $l=3.15e-07 $layer=LI1_cond $X=0.33 $Y=2.09
+ $X2=0.33 $Y2=2.405
r24 11 34 0.732293 $w=4.88e-07 $l=3e-08 $layer=LI1_cond $X=0.33 $Y=2.09 $X2=0.33
+ $Y2=2.06
r25 10 45 5.76222 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=0.235 $Y=1.665
+ $X2=0.235 $Y2=1.815
r26 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.665
r27 8 9 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=0.925
+ $X2=0.235 $Y2=1.295
r28 7 8 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=0.555
+ $X2=0.235 $Y2=0.925
r29 7 24 5.18599 $w=2.98e-07 $l=1.35e-07 $layer=LI1_cond $X=0.235 $Y=0.555
+ $X2=0.235 $Y2=0.42
r30 2 44 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.835 $X2=0.48 $Y2=1.98
r31 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.835 $X2=0.48 $Y2=2.91
r32 1 24 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.27 $X2=0.28 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_1%VPWR 1 2 3 12 18 20 22 27 28 29 35 39 45 49
r44 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 43 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 40 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.18 $Y2=3.33
r50 40 42 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 39 48 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.622 $Y2=3.33
r52 39 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 35 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.18 $Y2=3.33
r55 35 37 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 33 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 29 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 29 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 27 32 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 27 28 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.745 $Y=3.33 $X2=1
+ $Y2=3.33
r62 26 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 26 28 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.255 $Y=3.33 $X2=1
+ $Y2=3.33
r64 22 25 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=3.57 $Y=2.005
+ $X2=3.57 $Y2=2.95
r65 20 48 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.622 $Y2=3.33
r66 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.57 $Y2=2.95
r67 16 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=3.33
r68 16 18 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=2.38
r69 12 15 11.4917 $w=5.08e-07 $l=4.9e-07 $layer=LI1_cond $X=1 $Y=2.01 $X2=1
+ $Y2=2.5
r70 10 28 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=3.33
r71 10 15 17.4721 $w=5.08e-07 $l=7.45e-07 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=2.5
r72 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.835 $X2=3.57 $Y2=2.95
r73 3 22 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.835 $X2=3.57 $Y2=2.005
r74 2 18 300 $w=1.7e-07 $l=6.04276e-07 $layer=licon1_PDIFF $count=2 $X=2.055
+ $Y=1.835 $X2=2.18 $Y2=2.38
r75 1 15 300 $w=1.7e-07 $l=7.31659e-07 $layer=licon1_PDIFF $count=2 $X=0.77
+ $Y=1.835 $X2=0.91 $Y2=2.5
r76 1 12 600 $w=1.7e-07 $l=3.2078e-07 $layer=licon1_PDIFF $count=1 $X=0.77
+ $Y=1.835 $X2=1.015 $Y2=2.01
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r43 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r46 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r47 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.07
+ $Y2=0
r48 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.6
+ $Y2=0
r49 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r50 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r51 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r53 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 23 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.735
+ $Y2=0
r55 23 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.2
+ $Y2=0
r56 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.07
+ $Y2=0
r57 22 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.64
+ $Y2=0
r58 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r59 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r60 17 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.735
+ $Y2=0
r61 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.24
+ $Y2=0
r62 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r63 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r64 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0
r65 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0.4
r66 7 36 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0
r67 7 9 15.526 $w=3.58e-07 $l=4.85e-07 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0.57
r68 2 13 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=2.9
+ $Y=0.255 $X2=3.07 $Y2=0.4
r69 1 9 182 $w=1.7e-07 $l=3.69459e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.27 $X2=0.725 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_1%A_494_51# 1 2 9 11 12 15
c21 12 0 1.25093e-19 $X=2.715 $Y=1.12
r22 13 15 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.57 $Y=1.035
+ $X2=3.57 $Y2=0.4
r23 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.405 $Y=1.12
+ $X2=3.57 $Y2=1.035
r24 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.405 $Y=1.12
+ $X2=2.715 $Y2=1.12
r25 7 12 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=2.597 $Y=1.035
+ $X2=2.715 $Y2=1.12
r26 7 9 29.6693 $w=2.33e-07 $l=6.05e-07 $layer=LI1_cond $X=2.597 $Y=1.035
+ $X2=2.597 $Y2=0.43
r27 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.43
+ $Y=0.255 $X2=3.57 $Y2=0.4
r28 1 9 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.47
+ $Y=0.255 $X2=2.61 $Y2=0.43
.ends

