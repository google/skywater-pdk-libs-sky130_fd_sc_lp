* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2a_lp A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_674_416# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VPWR A1_N a_298_416# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_604_142# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_86_22# B2 a_674_416# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_298_416# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VPWR a_298_416# a_86_22# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VGND B1 a_604_142# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_274_48# A2_N a_298_416# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_86_22# a_298_416# a_604_142# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_86_22# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_116_48# a_86_22# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_86_22# a_116_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND A1_N a_274_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
