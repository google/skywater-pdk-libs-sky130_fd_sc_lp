* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_281_138# B1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.0941e+12p ps=9.59e+06u
M1001 a_84_28# a_281_138# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.78e+11p pd=3.12e+06u as=0p ps=0u
M1002 a_494_51# a_281_138# a_84_28# VNB nshort w=840000u l=150000u
+  ad=4.578e+11p pd=4.45e+06u as=2.226e+11p ps=2.21e+06u
M1003 a_584_367# A2 a_84_28# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.536e+11p pd=3.24e+06u as=0p ps=0u
M1004 VPWR A1 a_584_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_84_28# X VNB nshort w=840000u l=150000u
+  ad=7.35e+11p pd=5.49e+06u as=2.394e+11p ps=2.25e+06u
M1006 a_281_138# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1007 VGND A2 a_494_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_84_28# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1009 a_494_51# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
