# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__bushold0_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__bushold0_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN RESET
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.525000 1.355000 2.195000 ;
    END
  END RESET
  PIN X
    ANTENNADIFFAREA  0.228900 ;
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485000 1.525000 0.815000 2.365000 ;
        RECT 0.485000 2.365000 2.315000 2.535000 ;
        RECT 1.225000 0.255000 1.525000 0.840000 ;
        RECT 1.225000 0.840000 2.315000 1.015000 ;
        RECT 2.025000 1.015000 2.315000 2.365000 ;
        RECT 2.025000 2.535000 2.315000 3.050000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.085000  1.055000 0.625000 1.185000 ;
      RECT 0.085000  1.185000 1.855000 1.355000 ;
      RECT 0.085000  1.355000 0.315000 2.720000 ;
      RECT 0.085000  2.720000 0.425000 3.050000 ;
      RECT 0.335000  0.255000 0.625000 1.055000 ;
      RECT 0.795000  0.085000 1.055000 0.610000 ;
      RECT 0.835000  2.720000 1.165000 3.245000 ;
      RECT 1.605000  1.355000 1.855000 2.195000 ;
      RECT 1.975000  0.085000 2.305000 0.610000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_lp__bushold0_1
END LIBRARY
