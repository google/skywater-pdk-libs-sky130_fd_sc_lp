* File: sky130_fd_sc_lp__a311o_2.pxi.spice
* Created: Wed Sep  2 09:25:08 2020
* 
x_PM_SKY130_FD_SC_LP__A311O_2%A_85_21# N_A_85_21#_M1000_d N_A_85_21#_M1008_d
+ N_A_85_21#_M1002_d N_A_85_21#_c_67_n N_A_85_21#_M1012_g N_A_85_21#_M1001_g
+ N_A_85_21#_c_69_n N_A_85_21#_c_70_n N_A_85_21#_M1013_g N_A_85_21#_c_71_n
+ N_A_85_21#_M1004_g N_A_85_21#_c_73_n N_A_85_21#_c_74_n N_A_85_21#_c_75_n
+ N_A_85_21#_c_89_p N_A_85_21#_c_171_p N_A_85_21#_c_82_n N_A_85_21#_c_129_p
+ N_A_85_21#_c_175_p N_A_85_21#_c_76_n N_A_85_21#_c_83_n N_A_85_21#_c_77_n
+ N_A_85_21#_c_78_n N_A_85_21#_c_107_p PM_SKY130_FD_SC_LP__A311O_2%A_85_21#
x_PM_SKY130_FD_SC_LP__A311O_2%A3 N_A3_M1005_g N_A3_M1010_g A3 N_A3_c_197_n
+ N_A3_c_198_n PM_SKY130_FD_SC_LP__A311O_2%A3
x_PM_SKY130_FD_SC_LP__A311O_2%A2 N_A2_M1006_g N_A2_M1009_g A2 N_A2_c_230_n
+ N_A2_c_231_n PM_SKY130_FD_SC_LP__A311O_2%A2
x_PM_SKY130_FD_SC_LP__A311O_2%A1 N_A1_M1000_g N_A1_M1011_g A1 N_A1_c_263_n
+ N_A1_c_264_n PM_SKY130_FD_SC_LP__A311O_2%A1
x_PM_SKY130_FD_SC_LP__A311O_2%B1 N_B1_M1003_g N_B1_M1007_g B1 B1 N_B1_c_296_n
+ N_B1_c_297_n PM_SKY130_FD_SC_LP__A311O_2%B1
x_PM_SKY130_FD_SC_LP__A311O_2%C1 N_C1_c_327_n N_C1_M1008_g N_C1_M1002_g C1
+ N_C1_c_330_n PM_SKY130_FD_SC_LP__A311O_2%C1
x_PM_SKY130_FD_SC_LP__A311O_2%VPWR N_VPWR_M1001_s N_VPWR_M1004_s N_VPWR_M1009_d
+ N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_358_n
+ N_VPWR_c_359_n N_VPWR_c_360_n VPWR N_VPWR_c_361_n N_VPWR_c_353_n
+ N_VPWR_c_363_n PM_SKY130_FD_SC_LP__A311O_2%VPWR
x_PM_SKY130_FD_SC_LP__A311O_2%X N_X_M1012_s N_X_M1001_d N_X_c_410_n X X X X X X
+ X N_X_c_412_n X PM_SKY130_FD_SC_LP__A311O_2%X
x_PM_SKY130_FD_SC_LP__A311O_2%A_341_367# N_A_341_367#_M1005_d
+ N_A_341_367#_M1011_d N_A_341_367#_c_441_n N_A_341_367#_c_447_n
+ N_A_341_367#_c_442_n N_A_341_367#_c_443_n N_A_341_367#_c_445_n
+ PM_SKY130_FD_SC_LP__A311O_2%A_341_367#
x_PM_SKY130_FD_SC_LP__A311O_2%VGND N_VGND_M1012_d N_VGND_M1013_d N_VGND_M1003_d
+ N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n
+ VGND N_VGND_c_479_n N_VGND_c_480_n N_VGND_c_481_n N_VGND_c_482_n
+ PM_SKY130_FD_SC_LP__A311O_2%VGND
cc_1 VNB N_A_85_21#_c_67_n 0.0215272f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_2 VNB N_A_85_21#_M1001_g 0.0237353f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.465
cc_3 VNB N_A_85_21#_c_69_n 0.0120874f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.26
cc_4 VNB N_A_85_21#_c_70_n 0.0177049f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.185
cc_5 VNB N_A_85_21#_c_71_n 0.0330087f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.515
cc_6 VNB N_A_85_21#_M1004_g 0.00733047f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.465
cc_7 VNB N_A_85_21#_c_73_n 0.0151359f $X=-0.19 $Y=-0.245 $X2=0.537 $Y2=1.26
cc_8 VNB N_A_85_21#_c_74_n 0.00260664f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.35
cc_9 VNB N_A_85_21#_c_75_n 0.00146397f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.695
cc_10 VNB N_A_85_21#_c_76_n 0.00742189f $X=-0.19 $Y=-0.245 $X2=3.75 $Y2=0.93
cc_11 VNB N_A_85_21#_c_77_n 0.0229172f $X=-0.19 $Y=-0.245 $X2=3.895 $Y2=0.42
cc_12 VNB N_A_85_21#_c_78_n 8.37735e-19 $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.515
cc_13 VNB N_A3_M1005_g 0.0082987f $X=-0.19 $Y=-0.245 $X2=3.755 $Y2=1.835
cc_14 VNB A3 0.00685705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_c_197_n 0.0278854f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_16 VNB N_A3_c_198_n 0.0180061f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.335
cc_17 VNB N_A2_M1009_g 0.00819075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A2 0.00576765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_230_n 0.0306735f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_20 VNB N_A2_c_231_n 0.0174287f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.335
cc_21 VNB N_A1_M1011_g 0.00819075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A1 0.00564417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_263_n 0.0306098f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_24 VNB N_A1_c_264_n 0.019046f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.335
cc_25 VNB N_B1_M1007_g 0.00765658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB B1 0.00875679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B1_c_296_n 0.0279491f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.335
cc_28 VNB N_B1_c_297_n 0.0185641f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.465
cc_29 VNB N_C1_c_327_n 0.0237919f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=0.235
cc_30 VNB N_C1_M1002_g 0.0107928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB C1 0.0256801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_C1_c_330_n 0.0506368f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.335
cc_33 VNB N_VPWR_c_353_n 0.183584f $X=-0.19 $Y=-0.245 $X2=3.75 $Y2=0.93
cc_34 VNB N_X_c_410_n 6.93921e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB X 8.10132e-19 $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.335
cc_36 VNB N_X_c_412_n 0.00208358f $X=-0.19 $Y=-0.245 $X2=0.537 $Y2=1.26
cc_37 VNB N_VGND_c_474_n 0.0116069f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_38 VNB N_VGND_c_475_n 0.0487051f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_39 VNB N_VGND_c_476_n 0.0055721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_477_n 0.046745f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.185
cc_41 VNB N_VGND_c_478_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.655
cc_42 VNB N_VGND_c_479_n 0.0149091f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.465
cc_43 VNB N_VGND_c_480_n 0.0226629f $X=-0.19 $Y=-0.245 $X2=3.73 $Y2=1.785
cc_44 VNB N_VGND_c_481_n 0.235761f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.785
cc_45 VNB N_VGND_c_482_n 0.0123187f $X=-0.19 $Y=-0.245 $X2=3.895 $Y2=1.875
cc_46 VPB N_A_85_21#_M1001_g 0.0265098f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.465
cc_47 VPB N_A_85_21#_M1004_g 0.0210093f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.465
cc_48 VPB N_A_85_21#_c_75_n 4.19665e-19 $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.695
cc_49 VPB N_A_85_21#_c_82_n 0.0429727f $X=-0.19 $Y=1.655 $X2=3.73 $Y2=1.785
cc_50 VPB N_A_85_21#_c_83_n 0.0466985f $X=-0.19 $Y=1.655 $X2=3.895 $Y2=1.98
cc_51 VPB N_A3_M1005_g 0.0208086f $X=-0.19 $Y=1.655 $X2=3.755 $Y2=1.835
cc_52 VPB N_A2_M1009_g 0.0215545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A1_M1011_g 0.0215545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B1_M1007_g 0.0193532f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_C1_M1002_g 0.0251825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_354_n 0.0135853f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.185
cc_57 VPB N_VPWR_c_355_n 0.0635876f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.655
cc_58 VPB N_VPWR_c_356_n 0.0190923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_357_n 0.00564356f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.655
cc_60 VPB N_VPWR_c_358_n 0.00564356f $X=-0.19 $Y=1.655 $X2=0.537 $Y2=1.26
cc_61 VPB N_VPWR_c_359_n 0.0217315f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.35
cc_62 VPB N_VPWR_c_360_n 0.00632158f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.35
cc_63 VPB N_VPWR_c_361_n 0.0509561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_353_n 0.0552252f $X=-0.19 $Y=1.655 $X2=3.75 $Y2=0.93
cc_65 VPB N_VPWR_c_363_n 0.00632158f $X=-0.19 $Y=1.655 $X2=3.895 $Y2=2.95
cc_66 VPB X 0.00122414f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.335
cc_67 N_A_85_21#_M1004_g N_A3_M1005_g 0.031914f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A_85_21#_c_75_n N_A3_M1005_g 0.00325856f $X=1.16 $Y=1.695 $X2=0 $Y2=0
cc_69 N_A_85_21#_c_82_n N_A3_M1005_g 0.0155928f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_70 N_A_85_21#_c_71_n A3 4.0736e-19 $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_71 N_A_85_21#_c_74_n A3 0.0235285f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_72 N_A_85_21#_c_89_p A3 0.0240806f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_73 N_A_85_21#_c_82_n A3 0.0291344f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_74 N_A_85_21#_c_71_n N_A3_c_197_n 0.0214627f $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_75 N_A_85_21#_c_74_n N_A3_c_197_n 0.00108002f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_76 N_A_85_21#_c_89_p N_A3_c_197_n 0.00418644f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_77 N_A_85_21#_c_82_n N_A3_c_197_n 0.00123311f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_78 N_A_85_21#_c_70_n N_A3_c_198_n 0.00987982f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_79 N_A_85_21#_c_74_n N_A3_c_198_n 0.00334685f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_80 N_A_85_21#_c_89_p N_A3_c_198_n 0.0125968f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_81 N_A_85_21#_c_82_n N_A2_M1009_g 0.012393f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_82 N_A_85_21#_c_89_p A2 0.0235468f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_83 N_A_85_21#_c_82_n A2 0.0252525f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_84 N_A_85_21#_c_89_p N_A2_c_230_n 0.00111032f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_85 N_A_85_21#_c_82_n N_A2_c_230_n 0.00127412f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_86 N_A_85_21#_c_89_p N_A2_c_231_n 0.0124119f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_87 N_A_85_21#_c_82_n N_A1_M1011_g 0.0126492f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_88 N_A_85_21#_c_89_p A1 0.0128194f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_89 N_A_85_21#_c_82_n A1 0.02453f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_90 N_A_85_21#_c_107_p A1 0.0100434f $X=2.87 $Y=0.93 $X2=0 $Y2=0
cc_91 N_A_85_21#_c_82_n N_A1_c_263_n 0.00126f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_92 N_A_85_21#_c_107_p N_A1_c_263_n 0.0019056f $X=2.87 $Y=0.93 $X2=0 $Y2=0
cc_93 N_A_85_21#_c_89_p N_A1_c_264_n 0.010517f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_94 N_A_85_21#_c_82_n N_B1_M1007_g 0.0148719f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_95 N_A_85_21#_c_83_n N_B1_M1007_g 0.00394678f $X=3.895 $Y=1.98 $X2=0 $Y2=0
cc_96 N_A_85_21#_c_82_n B1 0.0531606f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_97 N_A_85_21#_c_76_n B1 0.0439922f $X=3.75 $Y=0.93 $X2=0 $Y2=0
cc_98 N_A_85_21#_c_107_p B1 0.00139459f $X=2.87 $Y=0.93 $X2=0 $Y2=0
cc_99 N_A_85_21#_c_82_n N_B1_c_296_n 0.00123311f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_100 N_A_85_21#_c_76_n N_B1_c_296_n 0.00418644f $X=3.75 $Y=0.93 $X2=0 $Y2=0
cc_101 N_A_85_21#_c_76_n N_B1_c_297_n 0.0105231f $X=3.75 $Y=0.93 $X2=0 $Y2=0
cc_102 N_A_85_21#_c_77_n N_B1_c_297_n 8.45867e-19 $X=3.895 $Y=0.42 $X2=0 $Y2=0
cc_103 N_A_85_21#_c_76_n N_C1_c_327_n 0.011968f $X=3.75 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_104 N_A_85_21#_c_77_n N_C1_c_327_n 0.00926328f $X=3.895 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_105 N_A_85_21#_c_82_n N_C1_M1002_g 0.017073f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_106 N_A_85_21#_c_83_n N_C1_M1002_g 0.0260918f $X=3.895 $Y=1.98 $X2=0 $Y2=0
cc_107 N_A_85_21#_c_82_n C1 0.0164787f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_108 N_A_85_21#_c_76_n C1 0.0170114f $X=3.75 $Y=0.93 $X2=0 $Y2=0
cc_109 N_A_85_21#_c_82_n N_C1_c_330_n 0.00787312f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_110 N_A_85_21#_c_76_n N_C1_c_330_n 0.00422869f $X=3.75 $Y=0.93 $X2=0 $Y2=0
cc_111 N_A_85_21#_c_82_n N_VPWR_M1004_s 0.00345945f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_112 N_A_85_21#_c_129_p N_VPWR_M1004_s 0.00167177f $X=1.245 $Y=1.785 $X2=0
+ $Y2=0
cc_113 N_A_85_21#_c_82_n N_VPWR_M1009_d 0.00532109f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_114 N_A_85_21#_M1001_g N_VPWR_c_355_n 0.00885808f $X=0.575 $Y=2.465 $X2=0
+ $Y2=0
cc_115 N_A_85_21#_c_73_n N_VPWR_c_355_n 0.00136241f $X=0.537 $Y=1.26 $X2=0 $Y2=0
cc_116 N_A_85_21#_M1001_g N_VPWR_c_356_n 0.00564131f $X=0.575 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_85_21#_M1004_g N_VPWR_c_356_n 0.00585385f $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_85_21#_c_71_n N_VPWR_c_357_n 3.13519e-19 $X=1.005 $Y=1.515 $X2=0
+ $Y2=0
cc_119 N_A_85_21#_M1004_g N_VPWR_c_357_n 0.0145975f $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_85_21#_c_82_n N_VPWR_c_357_n 0.0190746f $X=3.73 $Y=1.785 $X2=0 $Y2=0
cc_121 N_A_85_21#_c_129_p N_VPWR_c_357_n 0.0084752f $X=1.245 $Y=1.785 $X2=0
+ $Y2=0
cc_122 N_A_85_21#_c_83_n N_VPWR_c_361_n 0.0210467f $X=3.895 $Y=1.98 $X2=0 $Y2=0
cc_123 N_A_85_21#_M1002_d N_VPWR_c_353_n 0.00215158f $X=3.755 $Y=1.835 $X2=0
+ $Y2=0
cc_124 N_A_85_21#_M1001_g N_VPWR_c_353_n 0.0111233f $X=0.575 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_85_21#_M1004_g N_VPWR_c_353_n 0.0112505f $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_126 N_A_85_21#_c_83_n N_VPWR_c_353_n 0.0125689f $X=3.895 $Y=1.98 $X2=0 $Y2=0
cc_127 N_A_85_21#_M1001_g N_X_c_410_n 0.00873334f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_85_21#_M1004_g N_X_c_410_n 0.00239475f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A_85_21#_c_75_n N_X_c_410_n 0.00921753f $X=1.16 $Y=1.695 $X2=0 $Y2=0
cc_130 N_A_85_21#_c_78_n N_X_c_410_n 0.0169419f $X=1.115 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A_85_21#_M1001_g X 0.0136863f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A_85_21#_c_129_p X 0.00883267f $X=1.245 $Y=1.785 $X2=0 $Y2=0
cc_133 N_A_85_21#_M1001_g X 0.00134506f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A_85_21#_c_69_n X 0.00166885f $X=0.855 $Y=1.26 $X2=0 $Y2=0
cc_135 N_A_85_21#_c_71_n X 0.00115671f $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_85_21#_c_67_n N_X_c_412_n 0.00313789f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_137 N_A_85_21#_M1001_g N_X_c_412_n 0.00425435f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A_85_21#_c_69_n N_X_c_412_n 0.0105447f $X=0.855 $Y=1.26 $X2=0 $Y2=0
cc_139 N_A_85_21#_c_70_n N_X_c_412_n 0.00132459f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_140 N_A_85_21#_c_71_n N_X_c_412_n 0.00128254f $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A_85_21#_c_73_n N_X_c_412_n 0.00695144f $X=0.537 $Y=1.26 $X2=0 $Y2=0
cc_142 N_A_85_21#_c_74_n N_X_c_412_n 0.0169419f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_143 N_A_85_21#_M1001_g X 0.0120787f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_85_21#_c_82_n N_A_341_367#_M1005_d 0.00176773f $X=3.73 $Y=1.785
+ $X2=-0.19 $Y2=-0.245
cc_145 N_A_85_21#_c_82_n N_A_341_367#_M1011_d 0.00176773f $X=3.73 $Y=1.785 $X2=0
+ $Y2=0
cc_146 N_A_85_21#_c_82_n N_A_341_367#_c_441_n 0.0172972f $X=3.73 $Y=1.785 $X2=0
+ $Y2=0
cc_147 N_A_85_21#_c_82_n N_A_341_367#_c_442_n 0.0502156f $X=3.73 $Y=1.785 $X2=0
+ $Y2=0
cc_148 N_A_85_21#_c_82_n N_A_341_367#_c_443_n 0.0172972f $X=3.73 $Y=1.785 $X2=0
+ $Y2=0
cc_149 N_A_85_21#_c_83_n N_A_341_367#_c_443_n 0.00499344f $X=3.895 $Y=1.98 $X2=0
+ $Y2=0
cc_150 N_A_85_21#_c_83_n N_A_341_367#_c_445_n 0.0235322f $X=3.895 $Y=1.98 $X2=0
+ $Y2=0
cc_151 N_A_85_21#_c_82_n A_657_367# 0.00791466f $X=3.73 $Y=1.785 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_85_21#_c_74_n N_VGND_M1013_d 8.58642e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_153 N_A_85_21#_c_89_p N_VGND_M1013_d 0.0137531f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_154 N_A_85_21#_c_171_p N_VGND_M1013_d 0.00252966f $X=1.245 $Y=0.93 $X2=0
+ $Y2=0
cc_155 N_A_85_21#_c_76_n N_VGND_M1003_d 0.0058207f $X=3.75 $Y=0.93 $X2=0 $Y2=0
cc_156 N_A_85_21#_c_67_n N_VGND_c_475_n 0.00702751f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_157 N_A_85_21#_c_76_n N_VGND_c_476_n 0.0219723f $X=3.75 $Y=0.93 $X2=0 $Y2=0
cc_158 N_A_85_21#_c_175_p N_VGND_c_477_n 0.0212513f $X=2.87 $Y=0.38 $X2=0 $Y2=0
cc_159 N_A_85_21#_c_67_n N_VGND_c_479_n 0.00585385f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_160 N_A_85_21#_c_70_n N_VGND_c_479_n 0.00487821f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_161 N_A_85_21#_c_77_n N_VGND_c_480_n 0.0196832f $X=3.895 $Y=0.42 $X2=0 $Y2=0
cc_162 N_A_85_21#_M1000_d N_VGND_c_481_n 0.00350322f $X=2.675 $Y=0.235 $X2=0
+ $Y2=0
cc_163 N_A_85_21#_M1008_d N_VGND_c_481_n 0.00215158f $X=3.755 $Y=0.235 $X2=0
+ $Y2=0
cc_164 N_A_85_21#_c_67_n N_VGND_c_481_n 0.0114915f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_165 N_A_85_21#_c_70_n N_VGND_c_481_n 0.00824731f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A_85_21#_c_89_p N_VGND_c_481_n 0.0344835f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_167 N_A_85_21#_c_171_p N_VGND_c_481_n 9.31834e-19 $X=1.245 $Y=0.93 $X2=0
+ $Y2=0
cc_168 N_A_85_21#_c_175_p N_VGND_c_481_n 0.0127519f $X=2.87 $Y=0.38 $X2=0 $Y2=0
cc_169 N_A_85_21#_c_76_n N_VGND_c_481_n 0.0120825f $X=3.75 $Y=0.93 $X2=0 $Y2=0
cc_170 N_A_85_21#_c_77_n N_VGND_c_481_n 0.0118828f $X=3.895 $Y=0.42 $X2=0 $Y2=0
cc_171 N_A_85_21#_c_67_n N_VGND_c_482_n 6.00882e-19 $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_172 N_A_85_21#_c_70_n N_VGND_c_482_n 0.0119671f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_173 N_A_85_21#_c_71_n N_VGND_c_482_n 7.9281e-19 $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A_85_21#_c_89_p N_VGND_c_482_n 0.0274261f $X=2.705 $Y=0.93 $X2=0 $Y2=0
cc_175 N_A_85_21#_c_171_p N_VGND_c_482_n 0.0177173f $X=1.245 $Y=0.93 $X2=0 $Y2=0
cc_176 N_A_85_21#_c_89_p A_355_47# 0.0056012f $X=2.705 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_177 N_A_85_21#_c_89_p A_427_47# 0.012197f $X=2.705 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_178 A3 A2 0.0272043f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A3_c_197_n A2 3.63963e-19 $X=1.61 $Y=1.35 $X2=0 $Y2=0
cc_180 N_A3_M1005_g N_A2_c_230_n 0.0285329f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A3_c_197_n N_A2_c_230_n 0.0449631f $X=1.61 $Y=1.35 $X2=0 $Y2=0
cc_182 A3 N_A2_c_231_n 0.00197313f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A3_c_198_n N_A2_c_231_n 0.0449631f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_184 N_A3_M1005_g N_VPWR_c_357_n 0.0138976f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A3_M1005_g N_VPWR_c_359_n 0.00549284f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A3_M1005_g N_VPWR_c_353_n 0.0104373f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A3_M1005_g N_A_341_367#_c_441_n 0.0022433f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A3_M1005_g N_A_341_367#_c_447_n 0.0101065f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A3_c_198_n N_VGND_c_477_n 0.00487821f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_190 N_A3_c_198_n N_VGND_c_481_n 0.00446189f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_191 N_A3_c_198_n N_VGND_c_482_n 0.0166995f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_192 N_A2_M1009_g N_A1_M1011_g 0.0284258f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_193 A2 A1 0.0283653f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A2_c_230_n A1 0.00103548f $X=2.15 $Y=1.36 $X2=0 $Y2=0
cc_195 N_A2_c_230_n N_A1_c_263_n 0.0214125f $X=2.15 $Y=1.36 $X2=0 $Y2=0
cc_196 A2 N_A1_c_264_n 0.00107665f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A2_c_231_n N_A1_c_264_n 0.036177f $X=2.15 $Y=1.195 $X2=0 $Y2=0
cc_198 N_A2_M1009_g N_VPWR_c_358_n 0.0107817f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A2_M1009_g N_VPWR_c_359_n 0.00549284f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A2_M1009_g N_VPWR_c_353_n 0.010663f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_201 N_A2_M1009_g N_A_341_367#_c_441_n 7.32094e-19 $X=2.06 $Y=2.465 $X2=0
+ $Y2=0
cc_202 N_A2_M1009_g N_A_341_367#_c_447_n 0.0129587f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A2_M1009_g N_A_341_367#_c_442_n 0.0123084f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A2_M1009_g N_A_341_367#_c_445_n 8.44338e-19 $X=2.06 $Y=2.465 $X2=0
+ $Y2=0
cc_205 N_A2_c_231_n N_VGND_c_477_n 0.00585385f $X=2.15 $Y=1.195 $X2=0 $Y2=0
cc_206 N_A2_c_231_n N_VGND_c_481_n 0.00666612f $X=2.15 $Y=1.195 $X2=0 $Y2=0
cc_207 N_A2_c_231_n N_VGND_c_482_n 0.00338156f $X=2.15 $Y=1.195 $X2=0 $Y2=0
cc_208 N_A1_c_263_n N_B1_M1007_g 0.0285322f $X=2.69 $Y=1.36 $X2=0 $Y2=0
cc_209 A1 B1 0.0285755f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_210 N_A1_c_263_n B1 0.00209836f $X=2.69 $Y=1.36 $X2=0 $Y2=0
cc_211 A1 N_B1_c_296_n 3.71332e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_212 N_A1_c_263_n N_B1_c_296_n 0.0199439f $X=2.69 $Y=1.36 $X2=0 $Y2=0
cc_213 N_A1_c_264_n N_B1_c_297_n 0.0122901f $X=2.69 $Y=1.195 $X2=0 $Y2=0
cc_214 N_A1_M1011_g N_VPWR_c_358_n 0.0108912f $X=2.78 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A1_M1011_g N_VPWR_c_361_n 0.00549284f $X=2.78 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A1_M1011_g N_VPWR_c_353_n 0.010663f $X=2.78 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A1_M1011_g N_A_341_367#_c_447_n 8.49511e-19 $X=2.78 $Y=2.465 $X2=0
+ $Y2=0
cc_218 N_A1_M1011_g N_A_341_367#_c_442_n 0.0123084f $X=2.78 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A1_M1011_g N_A_341_367#_c_443_n 7.32094e-19 $X=2.78 $Y=2.465 $X2=0
+ $Y2=0
cc_220 N_A1_M1011_g N_A_341_367#_c_445_n 0.0127916f $X=2.78 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A1_c_264_n N_VGND_c_477_n 0.00585385f $X=2.69 $Y=1.195 $X2=0 $Y2=0
cc_222 N_A1_c_264_n N_VGND_c_481_n 0.00702334f $X=2.69 $Y=1.195 $X2=0 $Y2=0
cc_223 B1 N_C1_c_327_n 0.00146201f $X=3.515 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_224 N_B1_c_296_n N_C1_c_327_n 0.0214298f $X=3.23 $Y=1.35 $X2=-0.19 $Y2=-0.245
cc_225 N_B1_c_297_n N_C1_c_327_n 0.0256101f $X=3.23 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_226 B1 C1 0.0273733f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_227 N_B1_M1007_g N_C1_c_330_n 0.0637441f $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_228 B1 N_C1_c_330_n 0.0118564f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_229 N_B1_M1007_g N_VPWR_c_361_n 0.00549284f $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_230 N_B1_M1007_g N_VPWR_c_353_n 0.0101744f $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_231 N_B1_M1007_g N_A_341_367#_c_443_n 0.00346817f $X=3.21 $Y=2.465 $X2=0
+ $Y2=0
cc_232 N_B1_M1007_g N_A_341_367#_c_445_n 0.016217f $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_233 N_B1_c_297_n N_VGND_c_476_n 0.00574528f $X=3.23 $Y=1.185 $X2=0 $Y2=0
cc_234 N_B1_c_297_n N_VGND_c_477_n 0.00585385f $X=3.23 $Y=1.185 $X2=0 $Y2=0
cc_235 N_B1_c_297_n N_VGND_c_481_n 0.00684837f $X=3.23 $Y=1.185 $X2=0 $Y2=0
cc_236 N_C1_M1002_g N_VPWR_c_361_n 0.0054895f $X=3.68 $Y=2.465 $X2=0 $Y2=0
cc_237 N_C1_M1002_g N_VPWR_c_353_n 0.0112045f $X=3.68 $Y=2.465 $X2=0 $Y2=0
cc_238 N_C1_M1002_g N_A_341_367#_c_443_n 5.12803e-19 $X=3.68 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_C1_M1002_g N_A_341_367#_c_445_n 0.00257172f $X=3.68 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_C1_c_327_n N_VGND_c_476_n 0.00395775f $X=3.68 $Y=1.195 $X2=0 $Y2=0
cc_241 N_C1_c_327_n N_VGND_c_480_n 0.00579312f $X=3.68 $Y=1.195 $X2=0 $Y2=0
cc_242 N_C1_c_327_n N_VGND_c_481_n 0.00754289f $X=3.68 $Y=1.195 $X2=0 $Y2=0
cc_243 N_VPWR_c_353_n N_X_M1001_d 0.00310528f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_355_n X 0.0464612f $X=0.36 $Y=1.98 $X2=0 $Y2=0
cc_245 N_VPWR_c_356_n X 0.0157159f $X=1.15 $Y=3.33 $X2=0 $Y2=0
cc_246 N_VPWR_c_353_n X 0.010282f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_247 N_VPWR_c_353_n N_A_341_367#_M1005_d 0.00223819f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_248 N_VPWR_c_353_n N_A_341_367#_M1011_d 0.00223819f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_357_n N_A_341_367#_c_441_n 0.0123489f $X=1.315 $Y=2.13 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_357_n N_A_341_367#_c_447_n 0.058188f $X=1.315 $Y=2.13 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_358_n N_A_341_367#_c_447_n 0.0392681f $X=2.425 $Y=2.495 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_359_n N_A_341_367#_c_447_n 0.0177952f $X=2.26 $Y=3.33 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_353_n N_A_341_367#_c_447_n 0.0123247f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_254 N_VPWR_M1009_d N_A_341_367#_c_442_n 0.0149054f $X=2.135 $Y=1.835 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_358_n N_A_341_367#_c_442_n 0.0266856f $X=2.425 $Y=2.495 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_358_n N_A_341_367#_c_445_n 0.040512f $X=2.425 $Y=2.495 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_361_n N_A_341_367#_c_445_n 0.0177952f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_353_n N_A_341_367#_c_445_n 0.0123247f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_353_n A_657_367# 0.0137053f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_260 N_X_c_412_n N_VGND_c_475_n 0.00152359f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_261 N_X_c_412_n N_VGND_c_479_n 0.0138717f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_262 N_X_M1012_s N_VGND_c_481_n 0.00397496f $X=0.575 $Y=0.235 $X2=0 $Y2=0
cc_263 N_X_c_412_n N_VGND_c_481_n 0.00886411f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_264 N_VGND_c_481_n A_355_47# 0.00309736f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_265 N_VGND_c_481_n A_427_47# 0.00576233f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
