* File: sky130_fd_sc_lp__or2_4.pex.spice
* Created: Fri Aug 28 11:21:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2_4%B 3 6 8 9 12 13 14 18
c31 13 0 3.10066e-20 $X=0.24 $Y=1.295
c32 9 0 1.17514e-19 $X=0.37 $Y=1.335
r33 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.355
+ $Y=1.375 $X2=0.355 $Y2=1.375
r34 14 19 9.41432 $w=3.53e-07 $l=2.9e-07 $layer=LI1_cond $X=0.262 $Y=1.665
+ $X2=0.262 $Y2=1.375
r35 13 19 2.59705 $w=3.53e-07 $l=8e-08 $layer=LI1_cond $X=0.262 $Y=1.295
+ $X2=0.262 $Y2=1.375
r36 11 18 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.355 $Y=1.575
+ $X2=0.355 $Y2=1.375
r37 11 12 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.37 $Y=1.575
+ $X2=0.37 $Y2=1.725
r38 9 18 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.355 $Y=1.335
+ $X2=0.355 $Y2=1.375
r39 8 9 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.37 $Y=1.185 $X2=0.37
+ $Y2=1.335
r40 6 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.725
r41 3 8 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.655
+ $X2=0.475 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_4%A 3 7 9 12 13
c45 3 0 3.10066e-20 $X=0.835 $Y=2.465
r46 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.675
r47 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.345
r48 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.51 $X2=0.925 $Y2=1.51
r49 9 13 5.76222 $w=4.08e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=1.55
+ $X2=0.925 $Y2=1.55
r50 7 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.92 $Y=0.655
+ $X2=0.92 $Y2=1.345
r51 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.835 $Y=2.465
+ $X2=0.835 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_4%A_27_367# 1 2 9 13 17 21 25 29 33 37 39 41 43
+ 47 49 50 52 54 60 65 72
c118 43 0 1.17514e-19 $X=1.19 $Y=2.015
r119 69 70 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.84 $Y=1.5
+ $X2=2.27 $Y2=1.5
r120 61 72 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.52 $Y=1.5 $X2=2.7
+ $Y2=1.5
r121 61 70 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.52 $Y=1.5
+ $X2=2.27 $Y2=1.5
r122 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.5 $X2=2.52 $Y2=1.5
r123 58 69 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.5 $Y=1.5 $X2=1.84
+ $Y2=1.5
r124 58 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.5 $Y=1.5 $X2=1.41
+ $Y2=1.5
r125 57 60 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.5 $Y=1.5
+ $X2=2.52 $Y2=1.5
r126 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.5 $Y=1.5
+ $X2=1.5 $Y2=1.5
r127 55 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=1.5
+ $X2=1.275 $Y2=1.5
r128 55 57 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.36 $Y=1.5 $X2=1.5
+ $Y2=1.5
r129 53 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=1.585
+ $X2=1.275 $Y2=1.5
r130 53 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.275 $Y=1.585
+ $X2=1.275 $Y2=1.93
r131 52 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=1.415
+ $X2=1.275 $Y2=1.5
r132 51 52 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.275 $Y=1.175
+ $X2=1.275 $Y2=1.415
r133 49 51 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.19 $Y=1.08
+ $X2=1.275 $Y2=1.175
r134 49 50 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=1.19 $Y=1.08
+ $X2=0.83 $Y2=1.08
r135 45 50 6.86407 $w=1.9e-07 $l=1.50167e-07 $layer=LI1_cond $X=0.72 $Y=0.985
+ $X2=0.83 $Y2=1.08
r136 45 47 29.5968 $w=2.18e-07 $l=5.65e-07 $layer=LI1_cond $X=0.72 $Y=0.985
+ $X2=0.72 $Y2=0.42
r137 44 64 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=2.015
+ $X2=0.26 $Y2=2.015
r138 43 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.19 $Y=2.015
+ $X2=1.275 $Y2=1.93
r139 43 44 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.19 $Y=2.015
+ $X2=0.425 $Y2=2.015
r140 39 64 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.1 $X2=0.26
+ $Y2=2.015
r141 39 41 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.26 $Y=2.1
+ $X2=0.26 $Y2=2.95
r142 35 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.665
+ $X2=2.7 $Y2=1.5
r143 35 37 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.7 $Y=1.665 $X2=2.7
+ $Y2=2.465
r144 31 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.335
+ $X2=2.7 $Y2=1.5
r145 31 33 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.7 $Y=1.335
+ $X2=2.7 $Y2=0.655
r146 27 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.665
+ $X2=2.27 $Y2=1.5
r147 27 29 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.27 $Y=1.665
+ $X2=2.27 $Y2=2.465
r148 23 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.335
+ $X2=2.27 $Y2=1.5
r149 23 25 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.27 $Y=1.335
+ $X2=2.27 $Y2=0.655
r150 19 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=1.665
+ $X2=1.84 $Y2=1.5
r151 19 21 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.84 $Y=1.665
+ $X2=1.84 $Y2=2.465
r152 15 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=1.335
+ $X2=1.84 $Y2=1.5
r153 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.84 $Y=1.335
+ $X2=1.84 $Y2=0.655
r154 11 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.665
+ $X2=1.41 $Y2=1.5
r155 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.41 $Y=1.665
+ $X2=1.41 $Y2=2.465
r156 7 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.335
+ $X2=1.41 $Y2=1.5
r157 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.41 $Y=1.335
+ $X2=1.41 $Y2=0.655
r158 2 64 400 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.03
r159 2 41 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r160 1 47 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.705 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_4%VPWR 1 2 3 12 16 22 27 28 29 30 31 32 34 48 50
r49 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 45 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 39 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.125 $Y2=3.33
r54 39 41 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 34 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=1.125 $Y2=3.33
r58 34 36 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 32 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 32 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 32 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 30 44 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.915 $Y2=3.33
r64 29 47 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=3.08 $Y=3.33 $X2=3.12
+ $Y2=3.33
r65 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=2.915 $Y2=3.33
r66 27 41 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=2.055 $Y2=3.33
r68 26 44 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.22 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=3.33
+ $X2=2.055 $Y2=3.33
r70 22 25 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.915 $Y=2.2
+ $X2=2.915 $Y2=2.95
r71 20 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=3.33
r72 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=2.95
r73 16 19 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.2
+ $X2=2.055 $Y2=2.97
r74 14 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=3.33
r75 14 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=2.97
r76 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=3.245
+ $X2=1.125 $Y2=3.33
r77 10 12 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=1.125 $Y=3.245
+ $X2=1.125 $Y2=2.38
r78 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.915 $Y2=2.95
r79 3 22 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.915 $Y2=2.2
r80 2 19 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.97
r81 2 16 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.2
r82 1 12 300 $w=1.7e-07 $l=6.43584e-07 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=1.835 $X2=1.125 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41 42
+ 44 45 49 51
r60 49 51 1.37196 $w=4.18e-07 $l=5e-08 $layer=LI1_cond $X=3.065 $Y=1.245
+ $X2=3.065 $Y2=1.295
r61 44 49 2.50256 $w=4.2e-07 $l=9e-08 $layer=LI1_cond $X=3.065 $Y=1.155
+ $X2=3.065 $Y2=1.245
r62 44 45 9.68601 $w=4.18e-07 $l=3.53e-07 $layer=LI1_cond $X=3.065 $Y=1.312
+ $X2=3.065 $Y2=1.665
r63 44 51 0.466465 $w=4.18e-07 $l=1.7e-08 $layer=LI1_cond $X=3.065 $Y=1.312
+ $X2=3.065 $Y2=1.295
r64 43 45 2.46952 $w=4.18e-07 $l=9e-08 $layer=LI1_cond $X=3.065 $Y=1.755
+ $X2=3.065 $Y2=1.665
r65 40 42 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.58 $Y=1.85
+ $X2=2.485 $Y2=1.85
r66 39 43 8.16006 $w=1.9e-07 $l=2.53081e-07 $layer=LI1_cond $X=2.855 $Y=1.85
+ $X2=3.065 $Y2=1.755
r67 39 40 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=2.855 $Y=1.85
+ $X2=2.58 $Y2=1.85
r68 38 41 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.58 $Y=1.155
+ $X2=2.485 $Y2=1.155
r69 37 44 5.83931 $w=1.8e-07 $l=2.1e-07 $layer=LI1_cond $X=2.855 $Y=1.155
+ $X2=3.065 $Y2=1.155
r70 37 38 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=2.855 $Y=1.155
+ $X2=2.58 $Y2=1.155
r71 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.485 $Y=1.98
+ $X2=2.485 $Y2=2.91
r72 31 42 1.34256 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.485 $Y=1.945
+ $X2=2.485 $Y2=1.85
r73 31 33 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=2.485 $Y=1.945
+ $X2=2.485 $Y2=1.98
r74 27 41 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=2.485 $Y=1.065
+ $X2=2.485 $Y2=1.155
r75 27 29 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=2.485 $Y=1.065
+ $X2=2.485 $Y2=0.42
r76 25 42 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.39 $Y=1.85
+ $X2=2.485 $Y2=1.85
r77 25 26 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=2.39 $Y=1.85 $X2=1.72
+ $Y2=1.85
r78 23 41 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.39 $Y=1.155
+ $X2=2.485 $Y2=1.155
r79 23 24 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.39 $Y=1.155
+ $X2=1.72 $Y2=1.155
r80 19 21 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=1.63 $Y=1.98 $X2=1.63
+ $Y2=2.91
r81 17 26 6.82297 $w=1.9e-07 $l=1.32571e-07 $layer=LI1_cond $X=1.63 $Y=1.945
+ $X2=1.72 $Y2=1.85
r82 17 19 2.15657 $w=1.78e-07 $l=3.5e-08 $layer=LI1_cond $X=1.63 $Y=1.945
+ $X2=1.63 $Y2=1.98
r83 13 24 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=1.625 $Y=1.065
+ $X2=1.72 $Y2=1.155
r84 13 15 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=1.625 $Y=1.065
+ $X2=1.625 $Y2=0.42
r85 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.835 $X2=2.485 $Y2=2.91
r86 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.835 $X2=2.485 $Y2=1.98
r87 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=2.91
r88 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=1.98
r89 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.345
+ $Y=0.235 $X2=2.485 $Y2=0.42
r90 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.235 $X2=1.625 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_4%VGND 1 2 3 4 13 15 19 23 27 30 31 32 33 34 35
+ 37 51 56
r56 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r57 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r59 48 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r60 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r61 42 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.33 $Y=0 $X2=1.165
+ $Y2=0
r62 42 44 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.33 $Y=0 $X2=1.68
+ $Y2=0
r63 41 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r64 41 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r65 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 38 53 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r67 38 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r68 37 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1 $Y=0 $X2=1.165
+ $Y2=0
r69 37 40 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.72
+ $Y2=0
r70 35 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r71 35 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r72 35 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r73 33 47 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.64
+ $Y2=0
r74 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.915
+ $Y2=0
r75 32 50 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.12
+ $Y2=0
r76 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.915
+ $Y2=0
r77 30 44 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.68
+ $Y2=0
r78 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.055
+ $Y2=0
r79 29 47 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.64
+ $Y2=0
r80 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.055
+ $Y2=0
r81 25 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0
r82 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.38
r83 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0
r84 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0.38
r85 17 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0
r86 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0.36
r87 13 53 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r88 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r89 4 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.775
+ $Y=0.235 $X2=2.915 $Y2=0.38
r90 3 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.915
+ $Y=0.235 $X2=2.055 $Y2=0.38
r91 2 19 91 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=2 $X=0.995
+ $Y=0.235 $X2=1.165 $Y2=0.36
r92 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

