* File: sky130_fd_sc_lp__or4_0.spice
* Created: Wed Sep  2 10:31:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4_0.pex.spice"
.subckt sky130_fd_sc_lp__or4_0  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1000 N_A_54_482#_M1000_d N_D_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_C_M1009_g N_A_54_482#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0588 PD=1.04 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_54_482#_M1007_d N_B_M1007_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1302 PD=0.7 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_54_482#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=12.852 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_54_482#_M1001_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0735 PD=1.46 PS=0.77 NRD=0 NRS=7.14 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_137_482# N_D_M1005_g N_A_54_482#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.1113 PD=0.72 PS=1.37 NRD=44.5417 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1003 A_227_482# N_C_M1003_g A_137_482# VPB PHIGHVT L=0.15 W=0.42 AD=0.063
+ AS=0.063 PD=0.72 PS=0.72 NRD=44.5417 NRS=44.5417 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 A_317_482# N_B_M1006_g A_227_482# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.063 PD=0.63 PS=0.72 NRD=23.443 NRS=44.5417 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g A_317_482# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.140581 AS=0.0441 PD=1.05 PS=0.63 NRD=131.182 NRS=23.443 M=1 R=2.8
+ SA=75001.4 SB=75001 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_54_482#_M1004_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.214219 PD=1.81 PS=1.6 NRD=0 NRS=6.1464 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__or4_0.pxi.spice"
*
.ends
*
*
