* File: sky130_fd_sc_lp__sdfxtp_1.pex.spice
* Created: Wed Sep  2 10:36:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%A_78_123# 1 2 7 11 15 19 22 24 25 28 29 34
+ 40 42
c90 40 0 1.36701e-19 $X=1.07 $Y=1.82
c91 28 0 5.78633e-20 $X=2.15 $Y=2.13
r92 40 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.82
+ $X2=1.07 $Y2=1.655
r93 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.82 $X2=1.07 $Y2=1.82
r94 37 39 8.37255 $w=6.63e-07 $l=4.55e-07 $layer=LI1_cond $X=0.615 $Y=2.062
+ $X2=1.07 $Y2=2.062
r95 31 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.18 $Y=0.8
+ $X2=0.515 $Y2=0.8
r96 29 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=2.13
+ $X2=2.15 $Y2=2.295
r97 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=2.13 $X2=2.15 $Y2=2.13
r98 26 28 8.16314 $w=2.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.115 $Y=2.3
+ $X2=2.115 $Y2=2.13
r99 25 39 10.7777 $w=6.63e-07 $l=3.97019e-07 $layer=LI1_cond $X=1.235 $Y=2.385
+ $X2=1.07 $Y2=2.062
r100 24 26 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.995 $Y=2.385
+ $X2=2.115 $Y2=2.3
r101 24 25 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.995 $Y=2.385
+ $X2=1.235 $Y2=2.385
r102 20 37 4.82816 $w=3.3e-07 $l=4.08e-07 $layer=LI1_cond $X=0.615 $Y=2.47
+ $X2=0.615 $Y2=2.062
r103 20 22 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.615 $Y=2.47
+ $X2=0.615 $Y2=2.6
r104 19 37 8.00453 $w=6.63e-07 $l=6.05202e-07 $layer=LI1_cond $X=0.18 $Y=1.655
+ $X2=0.615 $Y2=2.062
r105 18 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.18 $Y=0.965
+ $X2=0.18 $Y2=0.8
r106 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.18 $Y=0.965
+ $X2=0.18 $Y2=1.655
r107 15 46 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.13 $Y=2.775
+ $X2=2.13 $Y2=2.295
r108 11 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.16 $Y=0.825
+ $X2=1.16 $Y2=1.415
r109 7 17 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.145 $Y=1.505
+ $X2=1.145 $Y2=1.415
r110 7 42 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.145 $Y=1.505
+ $X2=1.145 $Y2=1.655
r111 2 22 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.49
+ $Y=2.455 $X2=0.615 $Y2=2.6
r112 1 34 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.39
+ $Y=0.615 $X2=0.515 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%D 3 7 11 12 13 14 15 16 17 24
c50 3 0 6.71236e-20 $X=1.52 $Y=0.825
r51 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.61
+ $Y=1.45 $X2=1.61 $Y2=1.45
r52 16 17 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.615 $Y=1.665
+ $X2=1.615 $Y2=2.035
r53 16 25 7.74298 $w=3.18e-07 $l=2.15e-07 $layer=LI1_cond $X=1.615 $Y=1.665
+ $X2=1.615 $Y2=1.45
r54 15 25 5.58215 $w=3.18e-07 $l=1.55e-07 $layer=LI1_cond $X=1.615 $Y=1.295
+ $X2=1.615 $Y2=1.45
r55 14 15 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.615 $Y=0.925
+ $X2=1.615 $Y2=1.295
r56 13 14 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.615 $Y=0.555
+ $X2=1.615 $Y2=0.925
r57 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.61 $Y=1.79
+ $X2=1.61 $Y2=1.45
r58 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.79
+ $X2=1.61 $Y2=1.955
r59 10 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.285
+ $X2=1.61 $Y2=1.45
r60 7 12 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.7 $Y=2.775 $X2=1.7
+ $Y2=1.955
r61 3 10 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.52 $Y=0.825
+ $X2=1.52 $Y2=1.285
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%SCE 2 6 7 9 10 11 12 13 14 16 19 24 25 31
r68 29 31 10.1474 $w=2.85e-07 $l=6e-08 $layer=POLY_cond $X=0.53 $Y=1.31 $X2=0.59
+ $Y2=1.31
r69 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.31 $X2=0.53 $Y2=1.31
r70 24 25 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.31 $X2=1.2
+ $Y2=1.31
r71 24 30 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.72 $Y=1.31
+ $X2=0.53 $Y2=1.31
r72 21 23 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.59 $Y=2.27
+ $X2=0.83 $Y2=2.27
r73 17 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.245 $Y=0.275
+ $X2=2.245 $Y2=0.825
r74 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.34 $Y=2.345
+ $X2=1.34 $Y2=2.775
r75 13 23 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.27
+ $X2=0.83 $Y2=2.27
r76 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.265 $Y=2.27
+ $X2=1.34 $Y2=2.345
r77 12 13 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.265 $Y=2.27
+ $X2=0.905 $Y2=2.27
r78 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.17 $Y=0.2
+ $X2=2.245 $Y2=0.275
r79 10 11 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=2.17 $Y=0.2
+ $X2=0.805 $Y2=0.2
r80 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.345
+ $X2=0.83 $Y2=2.27
r81 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.83 $Y=2.345 $X2=0.83
+ $Y2=2.775
r82 4 31 23.6772 $w=2.85e-07 $l=2.24332e-07 $layer=POLY_cond $X=0.73 $Y=1.145
+ $X2=0.59 $Y2=1.31
r83 4 6 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.73 $Y=1.145 $X2=0.73
+ $Y2=0.825
r84 3 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.73 $Y=0.275
+ $X2=0.805 $Y2=0.2
r85 3 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.73 $Y=0.275 $X2=0.73
+ $Y2=0.825
r86 2 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.59 $Y=2.195
+ $X2=0.59 $Y2=2.27
r87 1 31 17.7656 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.475
+ $X2=0.59 $Y2=1.31
r88 1 2 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.59 $Y=1.475 $X2=0.59
+ $Y2=2.195
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%SCD 3 7 9 10 14
c49 7 0 2.6087e-19 $X=2.605 $Y=0.825
r50 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.59
+ $X2=2.515 $Y2=1.755
r51 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.59
+ $X2=2.515 $Y2=1.425
r52 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.515
+ $Y=1.59 $X2=2.515 $Y2=1.59
r53 10 15 4.80185 $w=2.98e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.645
+ $X2=2.515 $Y2=1.645
r54 9 15 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=2.16 $Y=1.645
+ $X2=2.515 $Y2=1.645
r55 7 16 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.605 $Y=0.825 $X2=2.605
+ $Y2=1.425
r56 3 17 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.6 $Y=2.775 $X2=2.6
+ $Y2=1.755
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%CLK 3 7 9 10 11 16
c48 16 0 1.76152e-19 $X=3.34 $Y=1.375
c49 9 0 9.46395e-20 $X=3.6 $Y=1.295
r50 16 19 82.2934 $w=5.15e-07 $l=5.05e-07 $layer=POLY_cond $X=3.247 $Y=1.375
+ $X2=3.247 $Y2=1.88
r51 16 18 46.971 $w=5.15e-07 $l=1.65e-07 $layer=POLY_cond $X=3.247 $Y=1.375
+ $X2=3.247 $Y2=1.21
r52 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.34
+ $Y=1.375 $X2=3.34 $Y2=1.375
r53 10 11 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.475 $Y=1.665
+ $X2=3.475 $Y2=2.035
r54 10 17 7.59565 $w=4.38e-07 $l=2.9e-07 $layer=LI1_cond $X=3.475 $Y=1.665
+ $X2=3.475 $Y2=1.375
r55 9 17 2.09535 $w=4.38e-07 $l=8e-08 $layer=LI1_cond $X=3.475 $Y=1.295
+ $X2=3.475 $Y2=1.375
r56 7 19 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=3.065 $Y=2.775
+ $X2=3.065 $Y2=1.88
r57 3 18 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.065 $Y=0.825
+ $X2=3.065 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%A_628_123# 1 2 9 12 16 20 24 28 30 32 33 34
+ 35 36 42 44 45 46 47 49 50 51 52 58 59 62 65 66 69 70 74 75 76 80 81 82 91
c227 81 0 5.86445e-20 $X=7.435 $Y=1.92
c228 76 0 6.8524e-20 $X=5.845 $Y=2.72
c229 75 0 6.83332e-20 $X=4.05 $Y=2.47
c230 74 0 1.44144e-19 $X=3.95 $Y=0.93
c231 69 0 9.01006e-21 $X=8.155 $Y=1.02
c232 44 0 1.76152e-19 $X=3.865 $Y=2.47
c233 36 0 1.6623e-19 $X=3.865 $Y=0.85
c234 35 0 7.51337e-20 $X=5.635 $Y=1.61
c235 34 0 1.76508e-19 $X=5.255 $Y=1.61
c236 20 0 3.05678e-20 $X=5.71 $Y=2.455
r237 81 86 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.435 $Y=1.92
+ $X2=7.22 $Y2=1.92
r238 80 83 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=7.477 $Y=1.92
+ $X2=7.477 $Y2=2.085
r239 80 82 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=7.477 $Y=1.92
+ $X2=7.477 $Y2=1.755
r240 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.435
+ $Y=1.92 $X2=7.435 $Y2=1.92
r241 76 77 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.845 $Y=2.72
+ $X2=5.845 $Y2=2.98
r242 73 74 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.95
+ $Y=0.93 $X2=3.95 $Y2=0.93
r243 70 91 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.155 $Y=1.02
+ $X2=8.155 $Y2=0.855
r244 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.155
+ $Y=1.02 $X2=8.155 $Y2=1.02
r245 67 69 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=8.12 $Y=1.295
+ $X2=8.12 $Y2=1.02
r246 65 67 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.99 $Y=1.38
+ $X2=8.12 $Y2=1.295
r247 65 66 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.99 $Y=1.38
+ $X2=7.605 $Y2=1.38
r248 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.52 $Y=1.465
+ $X2=7.605 $Y2=1.38
r249 63 82 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.52 $Y=1.465
+ $X2=7.52 $Y2=1.755
r250 62 83 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.435 $Y=2.635
+ $X2=7.435 $Y2=2.085
r251 60 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=2.72
+ $X2=5.845 $Y2=2.72
r252 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.35 $Y=2.72
+ $X2=7.435 $Y2=2.635
r253 59 60 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=7.35 $Y=2.72
+ $X2=5.93 $Y2=2.72
r254 58 76 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.635
+ $X2=5.845 $Y2=2.72
r255 57 58 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=5.845 $Y=1.705
+ $X2=5.845 $Y2=2.635
r256 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.63
+ $Y=1.61 $X2=5.63 $Y2=1.61
r257 52 57 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.76 $Y=1.61
+ $X2=5.845 $Y2=1.705
r258 52 54 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=5.76 $Y=1.61
+ $X2=5.63 $Y2=1.61
r259 50 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2.98
+ $X2=5.845 $Y2=2.98
r260 50 51 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=5.76 $Y=2.98
+ $X2=4.235 $Y2=2.98
r261 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.15 $Y=2.895
+ $X2=4.235 $Y2=2.98
r262 48 75 3.46198 $w=2.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.15 $Y=2.555
+ $X2=4.05 $Y2=2.47
r263 48 49 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.15 $Y=2.555
+ $X2=4.15 $Y2=2.895
r264 47 75 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=2.385
+ $X2=4.05 $Y2=2.47
r265 46 73 2.96797 $w=3.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.05 $Y=0.985
+ $X2=4.05 $Y2=0.85
r266 46 47 43.606 $w=3.68e-07 $l=1.4e-06 $layer=LI1_cond $X=4.05 $Y=0.985
+ $X2=4.05 $Y2=2.385
r267 44 75 3.05049 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.865 $Y=2.47
+ $X2=4.05 $Y2=2.47
r268 44 45 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.865 $Y=2.47
+ $X2=3.445 $Y2=2.47
r269 40 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.28 $Y=2.555
+ $X2=3.445 $Y2=2.47
r270 40 42 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.28 $Y=2.555
+ $X2=3.28 $Y2=2.6
r271 36 73 4.06722 $w=2.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.865 $Y=0.85
+ $X2=4.05 $Y2=0.85
r272 36 38 24.9696 $w=2.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.865 $Y=0.85
+ $X2=3.28 $Y2=0.85
r273 35 55 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=5.635 $Y=1.61
+ $X2=5.63 $Y2=1.61
r274 34 55 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=5.255 $Y=1.61
+ $X2=5.63 $Y2=1.61
r275 32 74 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=3.95 $Y=1.285
+ $X2=3.95 $Y2=0.93
r276 32 33 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.955 $Y=1.285
+ $X2=3.955 $Y2=1.435
r277 30 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=0.765
+ $X2=3.95 $Y2=0.93
r278 28 91 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.245 $Y=0.535
+ $X2=8.245 $Y2=0.855
r279 22 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.22 $Y=2.085
+ $X2=7.22 $Y2=1.92
r280 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.22 $Y=2.085
+ $X2=7.22 $Y2=2.665
r281 18 35 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.71 $Y=1.775
+ $X2=5.635 $Y2=1.61
r282 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.71 $Y=1.775
+ $X2=5.71 $Y2=2.455
r283 14 34 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.18 $Y=1.445
+ $X2=5.255 $Y2=1.61
r284 14 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.18 $Y=1.445
+ $X2=5.18 $Y2=0.835
r285 12 33 661.468 $w=1.5e-07 $l=1.29e-06 $layer=POLY_cond $X=4.05 $Y=2.725
+ $X2=4.05 $Y2=1.435
r286 9 30 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.04 $Y=0.445
+ $X2=4.04 $Y2=0.765
r287 2 42 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.14
+ $Y=2.455 $X2=3.28 $Y2=2.6
r288 1 38 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.14
+ $Y=0.615 $X2=3.28 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%A_823_47# 1 2 7 8 9 11 14 17 19 20 21 24 27
+ 33 34 38 42 44 45 46 48 49 50 53 54 56 61 63
c164 63 0 9.01006e-21 $X=7.585 $Y=0.865
c165 53 0 5.86445e-20 $X=7.6 $Y=1.03
c166 19 0 1.38024e-19 $X=7.585 $Y=1.395
c167 7 0 1.71289e-19 $X=5.205 $Y=2.06
r168 54 63 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.585 $Y=1.03
+ $X2=7.585 $Y2=0.865
r169 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.6
+ $Y=1.03 $X2=7.6 $Y2=1.03
r170 51 53 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=7.6 $Y=0.555
+ $X2=7.6 $Y2=1.03
r171 49 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.435 $Y=0.47
+ $X2=7.6 $Y2=0.555
r172 49 50 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.435 $Y=0.47
+ $X2=6.905 $Y2=0.47
r173 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.82 $Y=0.555
+ $X2=6.905 $Y2=0.47
r174 47 48 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.82 $Y=0.555
+ $X2=6.82 $Y2=0.815
r175 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.735 $Y=0.9
+ $X2=6.82 $Y2=0.815
r176 45 46 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=6.735 $Y=0.9
+ $X2=5.85 $Y2=0.9
r177 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.765 $Y=0.815
+ $X2=5.85 $Y2=0.9
r178 43 44 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.765 $Y=0.485
+ $X2=5.765 $Y2=0.815
r179 42 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=0.35
+ $X2=5.63 $Y2=0.515
r180 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.63
+ $Y=0.35 $X2=5.63 $Y2=0.35
r181 39 56 4.56504 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=4.595 $Y=0.375
+ $X2=4.5 $Y2=0.375
r182 39 41 54.2172 $w=2.18e-07 $l=1.035e-06 $layer=LI1_cond $X=4.595 $Y=0.375
+ $X2=5.63 $Y2=0.375
r183 38 43 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.68 $Y=0.375
+ $X2=5.765 $Y2=0.485
r184 38 41 2.61919 $w=2.18e-07 $l=5e-08 $layer=LI1_cond $X=5.68 $Y=0.375
+ $X2=5.63 $Y2=0.375
r185 33 36 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=4.5 $Y=1.63 $X2=4.5
+ $Y2=2.56
r186 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.5
+ $Y=1.63 $X2=4.5 $Y2=1.63
r187 31 56 1.87542 $w=1.9e-07 $l=1.1e-07 $layer=LI1_cond $X=4.5 $Y=0.485 $X2=4.5
+ $Y2=0.375
r188 31 33 66.8373 $w=1.88e-07 $l=1.145e-06 $layer=LI1_cond $X=4.5 $Y=0.485
+ $X2=4.5 $Y2=1.63
r189 27 56 4.56504 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=4.405 $Y=0.375
+ $X2=4.5 $Y2=0.375
r190 27 29 7.85757 $w=2.18e-07 $l=1.5e-07 $layer=LI1_cond $X=4.405 $Y=0.375
+ $X2=4.255 $Y2=0.375
r191 26 34 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.5 $Y=1.985
+ $X2=4.5 $Y2=1.63
r192 22 24 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=8 $Y=1.545 $X2=8
+ $Y2=2.685
r193 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.925 $Y=1.47
+ $X2=8 $Y2=1.545
r194 20 21 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=7.925 $Y=1.47
+ $X2=7.765 $Y2=1.47
r195 19 21 33.3473 $w=1.5e-07 $l=2.14243e-07 $layer=POLY_cond $X=7.585 $Y=1.395
+ $X2=7.765 $Y2=1.47
r196 18 54 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=7.585 $Y=1.045
+ $X2=7.585 $Y2=1.03
r197 18 19 56.1013 $w=3.6e-07 $l=3.5e-07 $layer=POLY_cond $X=7.585 $Y=1.045
+ $X2=7.585 $Y2=1.395
r198 17 63 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=7.48 $Y=0.535
+ $X2=7.48 $Y2=0.865
r199 14 61 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.61 $Y=0.835
+ $X2=5.61 $Y2=0.515
r200 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.28 $Y=2.135
+ $X2=5.28 $Y2=2.455
r201 8 26 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.665 $Y=2.06
+ $X2=4.5 $Y2=1.985
r202 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.205 $Y=2.06
+ $X2=5.28 $Y2=2.135
r203 7 8 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.205 $Y=2.06
+ $X2=4.665 $Y2=2.06
r204 2 36 600 $w=1.7e-07 $l=4.45814e-07 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=2.405 $X2=4.5 $Y2=2.56
r205 1 29 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.115
+ $Y=0.235 $X2=4.255 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%A_1201_99# 1 2 9 13 15 18 21 24 27
c65 15 0 7.51337e-20 $X=7 $Y=2.075
r66 26 27 10.0716 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=7.132 $Y=1.165
+ $X2=7.132 $Y2=1.335
r67 24 26 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=7.17 $Y=0.9
+ $X2=7.17 $Y2=1.165
r68 21 29 9.3345 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=7.085 $Y=1.685
+ $X2=7.085 $Y2=2.075
r69 21 27 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.085 $Y=1.685
+ $X2=7.085 $Y2=1.335
r70 18 32 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=6.182 $Y=1.85
+ $X2=6.182 $Y2=2.015
r71 18 31 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=6.182 $Y=1.85
+ $X2=6.182 $Y2=1.685
r72 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.195
+ $Y=1.85 $X2=6.195 $Y2=1.85
r73 15 29 2.03444 $w=7.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=2.075 $X2=7.085
+ $Y2=2.075
r74 15 17 12.3441 $w=7.78e-07 $l=8.05e-07 $layer=LI1_cond $X=7 $Y=2.075
+ $X2=6.195 $Y2=2.075
r75 13 32 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6.08 $Y=2.455
+ $X2=6.08 $Y2=2.015
r76 9 31 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=6.08 $Y=0.835
+ $X2=6.08 $Y2=1.685
r77 2 29 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=6.865
+ $Y=2.245 $X2=7.005 $Y2=2.38
r78 1 24 182 $w=1.7e-07 $l=5.96992e-07 $layer=licon1_NDIFF $count=1 $X=6.935
+ $Y=0.405 $X2=7.16 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%A_1051_125# 1 2 9 13 16 19 21 23 25 27 34
+ 35
c87 21 0 1.76508e-19 $X=5.465 $Y=2.045
c88 16 0 1.71289e-19 $X=5.2 $Y=1.875
r89 35 39 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=6.752 $Y=1.34
+ $X2=6.752 $Y2=1.505
r90 35 38 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=6.752 $Y=1.34
+ $X2=6.752 $Y2=1.175
r91 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.735
+ $Y=1.34 $X2=6.735 $Y2=1.34
r92 26 27 2.06925 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=5.51 $Y=1.26
+ $X2=5.312 $Y2=1.26
r93 25 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.65 $Y=1.26
+ $X2=6.735 $Y2=1.26
r94 25 26 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=6.65 $Y=1.26
+ $X2=5.51 $Y2=1.26
r95 21 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.465 $Y=1.96
+ $X2=5.2 $Y2=1.96
r96 21 23 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=5.465 $Y=2.045
+ $X2=5.465 $Y2=2.45
r97 17 27 4.36305 $w=2.07e-07 $l=1.16619e-07 $layer=LI1_cond $X=5.387 $Y=1.175
+ $X2=5.312 $Y2=1.26
r98 17 19 16.6987 $w=2.43e-07 $l=3.55e-07 $layer=LI1_cond $X=5.387 $Y=1.175
+ $X2=5.387 $Y2=0.82
r99 16 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.2 $Y=1.875 $X2=5.2
+ $Y2=1.96
r100 15 27 4.36305 $w=2.07e-07 $l=1.4854e-07 $layer=LI1_cond $X=5.2 $Y=1.345
+ $X2=5.312 $Y2=1.26
r101 15 16 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.2 $Y=1.345
+ $X2=5.2 $Y2=1.875
r102 13 38 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.86 $Y=0.725
+ $X2=6.86 $Y2=1.175
r103 9 39 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=6.79 $Y=2.665
+ $X2=6.79 $Y2=1.505
r104 2 23 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=2.245 $X2=5.495 $Y2=2.45
r105 1 19 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=5.255
+ $Y=0.625 $X2=5.395 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%A_1657_383# 1 2 9 13 15 17 19 22 24 25 28
+ 32 36 39 41 42 43 47 53
r94 48 53 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.615 $Y=1.5 $X2=9.615
+ $Y2=1.41
r95 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.615
+ $Y=1.5 $X2=9.615 $Y2=1.5
r96 44 47 6.51381 $w=2.28e-07 $l=1.3e-07 $layer=LI1_cond $X=9.485 $Y=1.53
+ $X2=9.615 $Y2=1.53
r97 41 43 4.27425 $w=2.37e-07 $l=1.24439e-07 $layer=LI1_cond $X=9.485 $Y=1.985
+ $X2=9.417 $Y2=2.08
r98 40 44 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.485 $Y=1.645
+ $X2=9.485 $Y2=1.53
r99 40 41 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.485 $Y=1.645
+ $X2=9.485 $Y2=1.985
r100 39 44 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.485 $Y=1.415
+ $X2=9.485 $Y2=1.53
r101 39 42 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.485 $Y=1.415
+ $X2=9.485 $Y2=0.985
r102 34 43 4.27425 $w=2.37e-07 $l=9.5e-08 $layer=LI1_cond $X=9.417 $Y=2.175
+ $X2=9.417 $Y2=2.08
r103 34 36 0.944625 $w=3.03e-07 $l=2.5e-08 $layer=LI1_cond $X=9.417 $Y=2.175
+ $X2=9.417 $Y2=2.2
r104 30 42 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.405 $Y=0.82
+ $X2=9.405 $Y2=0.985
r105 30 32 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=9.405 $Y=0.82
+ $X2=9.405 $Y2=0.48
r106 28 52 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=8.482 $Y=2.08
+ $X2=8.482 $Y2=2.245
r107 28 51 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=8.482 $Y=2.08
+ $X2=8.482 $Y2=1.915
r108 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.45
+ $Y=2.08 $X2=8.45 $Y2=2.08
r109 25 43 2.15711 $w=1.9e-07 $l=1.52e-07 $layer=LI1_cond $X=9.265 $Y=2.08
+ $X2=9.417 $Y2=2.08
r110 25 27 47.5742 $w=1.88e-07 $l=8.15e-07 $layer=LI1_cond $X=9.265 $Y=2.08
+ $X2=8.45 $Y2=2.08
r111 20 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.085 $Y=1.485
+ $X2=10.085 $Y2=1.41
r112 20 22 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=10.085 $Y=1.485
+ $X2=10.085 $Y2=2.465
r113 17 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.085 $Y=1.335
+ $X2=10.085 $Y2=1.41
r114 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.085 $Y=1.335
+ $X2=10.085 $Y2=0.805
r115 16 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.78 $Y=1.41
+ $X2=9.615 $Y2=1.41
r116 15 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.01 $Y=1.41
+ $X2=10.085 $Y2=1.41
r117 15 16 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=10.01 $Y=1.41
+ $X2=9.78 $Y2=1.41
r118 13 51 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=8.605 $Y=0.535
+ $X2=8.605 $Y2=1.915
r119 9 52 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.51 $Y=2.685
+ $X2=8.51 $Y2=2.245
r120 2 36 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.21
+ $Y=2.055 $X2=9.35 $Y2=2.2
r121 1 32 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=9.205
+ $Y=0.325 $X2=9.345 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%A_1459_449# 1 2 9 13 17 18 20 21 25 26 28
+ 31 32 37 39
c103 28 0 1.38024e-19 $X=8.505 $Y=1.305
r104 35 37 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=7.775 $Y=2.68
+ $X2=7.87 $Y2=2.68
r105 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.055
+ $Y=1.39 $X2=9.055 $Y2=1.39
r106 29 39 2.80976 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.59 $Y=1.56
+ $X2=8.505 $Y2=1.56
r107 29 31 10.9054 $w=5.08e-07 $l=4.65e-07 $layer=LI1_cond $X=8.59 $Y=1.56
+ $X2=9.055 $Y2=1.56
r108 28 39 3.9231 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=8.505 $Y=1.305
+ $X2=8.505 $Y2=1.56
r109 27 28 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=8.505 $Y=0.675
+ $X2=8.505 $Y2=1.305
r110 25 39 2.80976 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=8.42 $Y=1.73
+ $X2=8.505 $Y2=1.56
r111 25 26 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.42 $Y=1.73
+ $X2=7.955 $Y2=1.73
r112 21 27 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.42 $Y=0.51
+ $X2=8.505 $Y2=0.675
r113 21 23 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=8.42 $Y=0.51
+ $X2=8.03 $Y2=0.51
r114 20 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.87 $Y=2.515
+ $X2=7.87 $Y2=2.68
r115 19 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.87 $Y=1.815
+ $X2=7.955 $Y2=1.73
r116 19 20 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.87 $Y=1.815
+ $X2=7.87 $Y2=2.515
r117 17 32 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.055 $Y=1.73
+ $X2=9.055 $Y2=1.39
r118 17 18 44.4756 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.055 $Y=1.73
+ $X2=9.055 $Y2=1.895
r119 16 32 43.7316 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.055 $Y=1.225
+ $X2=9.055 $Y2=1.39
r120 13 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.135 $Y=2.475
+ $X2=9.135 $Y2=1.895
r121 9 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.13 $Y=0.645
+ $X2=9.13 $Y2=1.225
r122 2 35 600 $w=1.7e-07 $l=6.62722e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=2.245 $X2=7.775 $Y2=2.68
r123 1 23 182 $w=1.7e-07 $l=5.59911e-07 $layer=licon1_NDIFF $count=1 $X=7.555
+ $Y=0.325 $X2=8.03 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%VPWR 1 2 3 4 5 6 21 25 29 33 37 42 43 45 46
+ 47 49 61 68 76 83 84 87 90 97 100
c125 84 0 3.05678e-20 $X=10.32 $Y=3.33
c126 21 0 1.36701e-19 $X=1.08 $Y=2.805
r127 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r128 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r129 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r130 90 93 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.495 $Y=3.06
+ $X2=6.495 $Y2=3.33
r131 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 84 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r133 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r134 81 100 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=9.975 $Y=3.33
+ $X2=9.857 $Y2=3.33
r135 81 83 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.975 $Y=3.33
+ $X2=10.32 $Y2=3.33
r136 80 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r137 80 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r138 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r139 77 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.085 $Y=3.33
+ $X2=8.92 $Y2=3.33
r140 77 79 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.085 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 76 100 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=9.74 $Y=3.33
+ $X2=9.857 $Y2=3.33
r142 76 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.74 $Y=3.33
+ $X2=9.36 $Y2=3.33
r143 75 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r144 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r145 72 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r146 72 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r147 71 74 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r148 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r149 69 93 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.66 $Y=3.33
+ $X2=6.495 $Y2=3.33
r150 69 71 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.66 $Y=3.33 $X2=6.96
+ $Y2=3.33
r151 68 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.92 $Y2=3.33
r152 68 74 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.4 $Y2=3.33
r153 67 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r154 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r155 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r156 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r157 61 93 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.33 $Y=3.33
+ $X2=6.495 $Y2=3.33
r158 61 66 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.33 $Y=3.33 $X2=6
+ $Y2=3.33
r159 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r160 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r161 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r162 57 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r163 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r164 54 87 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=1.097 $Y2=3.33
r165 54 56 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=2.64 $Y2=3.33
r166 52 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r167 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r168 49 87 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=1.097 $Y2=3.33
r169 49 51 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.72 $Y2=3.33
r170 47 67 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33 $X2=6
+ $Y2=3.33
r171 47 64 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.08 $Y2=3.33
r172 45 59 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.635 $Y=3.33
+ $X2=3.6 $Y2=3.33
r173 45 46 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.635 $Y=3.33
+ $X2=3.765 $Y2=3.33
r174 44 63 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.895 $Y=3.33
+ $X2=4.08 $Y2=3.33
r175 44 46 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.895 $Y=3.33
+ $X2=3.765 $Y2=3.33
r176 42 56 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.64 $Y2=3.33
r177 42 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.85 $Y2=3.33
r178 41 59 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.6 $Y2=3.33
r179 41 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.85 $Y2=3.33
r180 37 40 47.5689 $w=2.33e-07 $l=9.7e-07 $layer=LI1_cond $X=9.857 $Y=1.98
+ $X2=9.857 $Y2=2.95
r181 35 100 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=9.857 $Y=3.245
+ $X2=9.857 $Y2=3.33
r182 35 40 14.4668 $w=2.33e-07 $l=2.95e-07 $layer=LI1_cond $X=9.857 $Y=3.245
+ $X2=9.857 $Y2=2.95
r183 31 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.92 $Y=3.245
+ $X2=8.92 $Y2=3.33
r184 31 33 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=8.92 $Y=3.245
+ $X2=8.92 $Y2=2.43
r185 27 46 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=3.245
+ $X2=3.765 $Y2=3.33
r186 27 29 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=3.765 $Y=3.245
+ $X2=3.765 $Y2=2.89
r187 23 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=3.33
r188 23 25 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=2.825
r189 19 87 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.097 $Y=3.245
+ $X2=1.097 $Y2=3.33
r190 19 21 17.189 $w=2.93e-07 $l=4.4e-07 $layer=LI1_cond $X=1.097 $Y=3.245
+ $X2=1.097 $Y2=2.805
r191 6 40 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=9.745
+ $Y=1.835 $X2=9.87 $Y2=2.95
r192 6 37 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.745
+ $Y=1.835 $X2=9.87 $Y2=1.98
r193 5 33 300 $w=1.7e-07 $l=3.56791e-07 $layer=licon1_PDIFF $count=2 $X=8.585
+ $Y=2.475 $X2=8.92 $Y2=2.43
r194 4 90 600 $w=1.7e-07 $l=9.70219e-07 $layer=licon1_PDIFF $count=1 $X=6.155
+ $Y=2.245 $X2=6.495 $Y2=3.06
r195 3 29 600 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=2.405 $X2=3.8 $Y2=2.89
r196 2 25 600 $w=1.7e-07 $l=4.44916e-07 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=2.455 $X2=2.84 $Y2=2.825
r197 1 21 600 $w=1.7e-07 $l=4.28661e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=2.455 $X2=1.08 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%A_319_123# 1 2 3 4 13 19 21 22 24 25 28 30
+ 34 36 37 43 44 46
c122 37 0 5.78633e-20 $X=2.785 $Y=2.405
r123 44 50 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.04 $Y=2.39
+ $X2=4.85 $Y2=2.39
r124 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.405
+ $X2=5.04 $Y2=2.405
r125 40 49 5.49324 $w=3.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=2.405
+ $X2=2.57 $Y2=2.49
r126 40 46 10.595 $w=3.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.57 $Y=2.405
+ $X2=2.57 $Y2=2.12
r127 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=2.405
+ $X2=2.64 $Y2=2.405
r128 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=2.405
+ $X2=2.64 $Y2=2.405
r129 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.405
+ $X2=5.04 $Y2=2.405
r130 36 37 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=4.895 $Y=2.405
+ $X2=2.785 $Y2=2.405
r131 31 34 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.85 $Y=0.83
+ $X2=4.965 $Y2=0.83
r132 30 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.85 $Y=2.225
+ $X2=4.85 $Y2=2.39
r133 29 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.85 $Y=0.995
+ $X2=4.85 $Y2=0.83
r134 29 30 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=4.85 $Y=0.995
+ $X2=4.85 $Y2=2.225
r135 27 28 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=2.035
r136 26 46 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.725 $Y=2.12
+ $X2=2.57 $Y2=2.12
r137 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=2.12
+ $X2=2.99 $Y2=2.035
r138 25 26 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.905 $Y=2.12
+ $X2=2.725 $Y2=2.12
r139 24 49 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.5 $Y=2.64 $X2=2.5
+ $Y2=2.49
r140 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=1.24
+ $X2=2.99 $Y2=1.325
r141 21 22 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.905 $Y=1.24
+ $X2=2.195 $Y2=1.24
r142 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.07 $Y=1.155
+ $X2=2.195 $Y2=1.24
r143 17 19 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=2.07 $Y=1.155
+ $X2=2.07 $Y2=0.85
r144 13 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=2.805
+ $X2=2.5 $Y2=2.64
r145 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.415 $Y=2.805
+ $X2=1.915 $Y2=2.805
r146 4 44 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.94
+ $Y=2.245 $X2=5.065 $Y2=2.39
r147 3 15 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.775
+ $Y=2.455 $X2=1.915 $Y2=2.805
r148 2 34 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.625 $X2=4.965 $Y2=0.83
r149 1 19 182 $w=1.7e-07 $l=5.39861e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.615 $X2=2.03 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%Q 1 2 7 8 9 10 11 12 13
r13 13 39 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=10.33 $Y=2.775
+ $X2=10.33 $Y2=2.91
r14 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.33 $Y=2.405
+ $X2=10.33 $Y2=2.775
r15 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.33 $Y=1.98
+ $X2=10.33 $Y2=2.405
r16 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.33 $Y=1.665
+ $X2=10.33 $Y2=1.98
r17 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.33 $Y=1.295
+ $X2=10.33 $Y2=1.665
r18 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.33 $Y=0.925
+ $X2=10.33 $Y2=1.295
r19 7 8 16.8598 $w=2.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.33 $Y=0.53
+ $X2=10.33 $Y2=0.925
r20 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.835 $X2=10.3 $Y2=2.91
r21 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.835 $X2=10.3 $Y2=1.98
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.16
+ $Y=0.385 $X2=10.3 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_1%VGND 1 2 3 4 5 6 21 25 29 33 35 39 43 46 47
+ 49 50 52 53 54 69 76 83 84 87 90 93
c113 84 0 6.71236e-20 $X=10.32 $Y=0
c114 69 0 1.44144e-19 $X=6.225 $Y=0
r115 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r116 90 91 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r117 88 91 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.88
+ $Y2=0
r118 87 88 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r119 84 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r120 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r121 81 93 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=10.025 $Y=0
+ $X2=9.882 $Y2=0
r122 81 83 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.025 $Y=0
+ $X2=10.32 $Y2=0
r123 80 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r124 80 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r125 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r126 77 90 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=9.02 $Y=0 $X2=8.915
+ $Y2=0
r127 77 79 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.02 $Y=0 $X2=9.36
+ $Y2=0
r128 76 93 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=9.74 $Y=0 $X2=9.882
+ $Y2=0
r129 76 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.74 $Y=0 $X2=9.36
+ $Y2=0
r130 75 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r131 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r132 71 74 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r133 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r134 69 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.39
+ $Y2=0
r135 69 74 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6
+ $Y2=0
r136 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r137 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r138 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r139 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r140 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r141 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r142 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r143 58 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r144 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r145 54 75 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=6
+ $Y2=0
r146 54 72 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=4.08
+ $Y2=0
r147 52 67 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.66 $Y=0 $X2=3.6
+ $Y2=0
r148 52 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.66 $Y=0 $X2=3.79
+ $Y2=0
r149 51 71 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.92 $Y=0 $X2=4.08
+ $Y2=0
r150 51 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.92 $Y=0 $X2=3.79
+ $Y2=0
r151 49 64 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.655 $Y=0 $X2=2.64
+ $Y2=0
r152 49 50 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.655 $Y=0 $X2=2.8
+ $Y2=0
r153 48 67 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=3.6
+ $Y2=0
r154 48 50 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.8
+ $Y2=0
r155 46 57 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.84 $Y=0 $X2=0.72
+ $Y2=0
r156 46 47 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.84 $Y=0 $X2=0.945
+ $Y2=0
r157 45 61 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=1.2
+ $Y2=0
r158 45 47 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=0.945
+ $Y2=0
r159 41 93 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=9.882 $Y=0.085
+ $X2=9.882 $Y2=0
r160 41 43 17.9943 $w=2.83e-07 $l=4.45e-07 $layer=LI1_cond $X=9.882 $Y=0.085
+ $X2=9.882 $Y2=0.53
r161 37 90 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.915 $Y=0.085
+ $X2=8.915 $Y2=0
r162 37 39 20.3333 $w=2.08e-07 $l=3.85e-07 $layer=LI1_cond $X=8.915 $Y=0.085
+ $X2=8.915 $Y2=0.47
r163 36 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.39
+ $Y2=0
r164 35 90 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.81 $Y=0 $X2=8.915
+ $Y2=0
r165 35 36 147.118 $w=1.68e-07 $l=2.255e-06 $layer=LI1_cond $X=8.81 $Y=0
+ $X2=6.555 $Y2=0
r166 31 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.39 $Y2=0
r167 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.39 $Y2=0.55
r168 27 53 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0
r169 27 29 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0.38
r170 23 50 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0
r171 23 25 27.2215 $w=2.88e-07 $l=6.85e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.77
r172 19 47 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.945 $Y=0.085
+ $X2=0.945 $Y2=0
r173 19 21 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=0.945 $Y=0.085
+ $X2=0.945 $Y2=0.76
r174 6 43 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=9.745
+ $Y=0.385 $X2=9.87 $Y2=0.53
r175 5 39 91 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=2 $X=8.68
+ $Y=0.325 $X2=8.915 $Y2=0.47
r176 4 33 182 $w=1.7e-07 $l=2.69907e-07 $layer=licon1_NDIFF $count=1 $X=6.155
+ $Y=0.625 $X2=6.39 $Y2=0.55
r177 3 29 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.7
+ $Y=0.235 $X2=3.825 $Y2=0.38
r178 2 25 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.68
+ $Y=0.615 $X2=2.82 $Y2=0.77
r179 1 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.805
+ $Y=0.615 $X2=0.945 $Y2=0.76
.ends

