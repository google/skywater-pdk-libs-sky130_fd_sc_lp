* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VGND S a_266_132# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_518_434# a_488_106# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_105_22# A0 a_446_132# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_105_22# A1 a_518_434# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_266_132# A1 a_105_22# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_105_22# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VPWR S a_288_434# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND S a_488_106# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_446_132# a_488_106# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR S a_488_106# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 X a_105_22# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_288_434# A0 a_105_22# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
