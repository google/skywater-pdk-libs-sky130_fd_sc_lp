* File: sky130_fd_sc_lp__inv_lp.pxi.spice
* Created: Fri Aug 28 10:38:42 2020
* 
x_PM_SKY130_FD_SC_LP__INV_LP%A N_A_M1000_g N_A_M1001_g N_A_M1002_g A A
+ N_A_c_27_n PM_SKY130_FD_SC_LP__INV_LP%A
x_PM_SKY130_FD_SC_LP__INV_LP%VPWR N_VPWR_M1001_s N_VPWR_c_49_n N_VPWR_c_50_n
+ N_VPWR_c_51_n VPWR N_VPWR_c_52_n N_VPWR_c_48_n PM_SKY130_FD_SC_LP__INV_LP%VPWR
x_PM_SKY130_FD_SC_LP__INV_LP%Y N_Y_M1002_d N_Y_M1001_d Y Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__INV_LP%Y
x_PM_SKY130_FD_SC_LP__INV_LP%VGND N_VGND_M1000_s N_VGND_c_79_n N_VGND_c_80_n
+ VGND N_VGND_c_81_n N_VGND_c_82_n PM_SKY130_FD_SC_LP__INV_LP%VGND
cc_1 VNB N_A_M1000_g 0.0278525f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.545
cc_2 VNB N_A_M1001_g 0.00225235f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.48
cc_3 VNB N_A_M1002_g 0.0249157f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.545
cc_4 VNB A 0.0374652f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_A_c_27_n 0.0854047f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.12
cc_6 VNB N_VPWR_c_48_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.12
cc_7 VNB Y 0.0229869f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.48
cc_8 VNB Y 0.044379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_VGND_c_79_n 0.0133568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_80_n 0.0277707f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.48
cc_11 VNB N_VGND_c_81_n 0.0290825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_82_n 0.123637f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_13 VPB N_A_M1001_g 0.0501821f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=2.48
cc_14 VPB A 0.0222253f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_15 VPB N_VPWR_c_49_n 0.0498161f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=2.48
cc_16 VPB N_VPWR_c_50_n 0.0166223f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.545
cc_17 VPB N_VPWR_c_51_n 0.00598038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_18 VPB N_VPWR_c_52_n 0.0200323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_19 VPB N_VPWR_c_48_n 0.0619474f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.12
cc_20 VPB Y 0.0152399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_21 VPB Y 0.0357849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB Y 0.0093975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_23 N_A_M1001_g N_VPWR_c_49_n 0.0264097f $X=0.885 $Y=2.48 $X2=0 $Y2=0
cc_24 A N_VPWR_c_49_n 0.0291672f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_25 N_A_c_27_n N_VPWR_c_49_n 0.00157358f $X=0.635 $Y=1.12 $X2=0 $Y2=0
cc_26 N_A_M1001_g N_VPWR_c_52_n 0.00687065f $X=0.885 $Y=2.48 $X2=0 $Y2=0
cc_27 N_A_M1001_g N_VPWR_c_48_n 0.0131127f $X=0.885 $Y=2.48 $X2=0 $Y2=0
cc_28 N_A_M1000_g Y 0.00130204f $X=0.545 $Y=0.545 $X2=0 $Y2=0
cc_29 N_A_M1002_g Y 0.0104538f $X=0.935 $Y=0.545 $X2=0 $Y2=0
cc_30 N_A_M1002_g Y 0.0379424f $X=0.935 $Y=0.545 $X2=0 $Y2=0
cc_31 A Y 0.0503992f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_32 N_A_M1001_g Y 0.0159088f $X=0.885 $Y=2.48 $X2=0 $Y2=0
cc_33 N_A_M1001_g Y 0.00451956f $X=0.885 $Y=2.48 $X2=0 $Y2=0
cc_34 N_A_M1000_g N_VGND_c_80_n 0.0142118f $X=0.545 $Y=0.545 $X2=0 $Y2=0
cc_35 N_A_M1002_g N_VGND_c_80_n 0.00197399f $X=0.935 $Y=0.545 $X2=0 $Y2=0
cc_36 A N_VGND_c_80_n 0.0291689f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_37 N_A_M1000_g N_VGND_c_81_n 0.00407525f $X=0.545 $Y=0.545 $X2=0 $Y2=0
cc_38 N_A_M1002_g N_VGND_c_81_n 0.00461273f $X=0.935 $Y=0.545 $X2=0 $Y2=0
cc_39 N_A_M1000_g N_VGND_c_82_n 0.00777674f $X=0.545 $Y=0.545 $X2=0 $Y2=0
cc_40 N_A_M1002_g N_VGND_c_82_n 0.00910201f $X=0.935 $Y=0.545 $X2=0 $Y2=0
cc_41 N_VPWR_c_52_n Y 0.0158357f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_42 N_VPWR_c_48_n Y 0.0121432f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_43 N_VPWR_c_49_n Y 0.0684934f $X=0.62 $Y=2.125 $X2=0 $Y2=0
cc_44 Y N_VGND_c_80_n 0.0145731f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_45 Y N_VGND_c_81_n 0.016801f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_46 Y N_VGND_c_82_n 0.0122049f $X=1.115 $Y=0.47 $X2=0 $Y2=0
