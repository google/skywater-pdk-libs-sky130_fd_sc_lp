* File: sky130_fd_sc_lp__ha_4.spice
* Created: Fri Aug 28 10:36:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ha_4.pex.spice"
.subckt sky130_fd_sc_lp__ha_4  VNB VPB A B VPWR SUM COUT VGND
* 
* VGND	VGND
* COUT	COUT
* SUM	SUM
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1009 N_SUM_M1009_d N_A_110_263#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75005 A=0.126 P=1.98 MULT=1
MM1021 N_SUM_M1009_d N_A_110_263#_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.6 A=0.126 P=1.98 MULT=1
MM1022 N_SUM_M1022_d N_A_110_263#_M1022_g N_VGND_M1021_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.2 A=0.126 P=1.98 MULT=1
MM1034 N_SUM_M1022_d N_A_110_263#_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75003.8 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1034_s N_A_454_263#_M1016_g N_COUT_M1016_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1019_d N_A_454_263#_M1019_g N_COUT_M1016_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1030 N_VGND_M1019_d N_A_454_263#_M1030_g N_COUT_M1030_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1033 N_VGND_M1033_d N_A_454_263#_M1033_g N_COUT_M1030_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=1.428 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1020 N_A_851_47#_M1020_d N_A_M1020_g N_VGND_M1033_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=9.996 M=1 R=5.6 SA=75003.7
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1001 N_A_454_263#_M1001_d N_B_M1001_g N_A_851_47#_M1020_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1002 N_A_454_263#_M1001_d N_B_M1002_g N_A_851_47#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.136 M=1 R=5.6
+ SA=75004.6 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1031 N_A_851_47#_M1002_s N_A_M1031_g N_VGND_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.2226 PD=1.16 PS=2.21 NRD=3.564 NRS=0 M=1 R=5.6 SA=75005.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_B_M1010_g N_A_1284_65#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1848 AS=0.2226 PD=1.28 PS=2.21 NRD=11.424 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1011 N_A_1284_65#_M1011_d N_A_M1011_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1848 PD=1.12 PS=1.28 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.8
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1024 N_A_1284_65#_M1011_d N_A_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2625 PD=1.12 PS=1.465 NRD=0 NRS=36.78 M=1 R=5.6 SA=75001.2
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1029 N_VGND_M1024_s N_B_M1029_g N_A_1284_65#_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2625 AS=0.1176 PD=1.465 PS=1.12 NRD=36.78 NRS=0 M=1 R=5.6 SA=75002
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_110_263#_M1005_d N_A_454_263#_M1005_g N_A_1284_65#_M1029_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75002.4 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1026 N_A_110_263#_M1005_d N_A_454_263#_M1026_g N_A_1284_65#_M1026_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.3528 PD=1.12 PS=2.52 NRD=0 NRS=19.284 M=1 R=5.6
+ SA=75002.8 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1003 N_SUM_M1003_d N_A_110_263#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.1 A=0.189 P=2.82 MULT=1
MM1014 N_SUM_M1003_d N_A_110_263#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.6 A=0.189 P=2.82 MULT=1
MM1025 N_SUM_M1025_d N_A_110_263#_M1025_g N_VPWR_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.2 A=0.189 P=2.82 MULT=1
MM1035 N_SUM_M1025_d N_A_110_263#_M1035_g N_VPWR_M1035_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.8 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1035_s N_A_454_263#_M1006_g N_COUT_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A_454_263#_M1012_g N_COUT_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1023 N_VPWR_M1012_d N_A_454_263#_M1023_g N_COUT_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1032 N_VPWR_M1032_d N_A_454_263#_M1032_g N_COUT_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.24885 AS=0.1764 PD=1.655 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1032_d N_A_M1000_g N_A_454_263#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.24885 AS=0.1764 PD=1.655 PS=1.54 NRD=17.9664 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_B_M1007_g N_A_454_263#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1027 N_VPWR_M1007_d N_B_M1027_g N_A_454_263#_M1027_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_A_M1017_g N_A_454_263#_M1027_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1008 N_A_110_263#_M1008_d N_B_M1008_g N_A_1367_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_A_1367_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.360275 AS=0.1764 PD=1.905 PS=1.54 NRD=18.7544 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75002.6 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1013_d N_A_M1018_g N_A_1367_367#_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.360275 AS=0.1764 PD=1.905 PS=1.54 NRD=24.9993 NRS=0 M=1 R=8.4
+ SA=75001.3 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1028 N_A_110_263#_M1028_d N_B_M1028_g N_A_1367_367#_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.28035 AS=0.1764 PD=1.705 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75001.8 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1004 N_A_110_263#_M1028_d N_A_454_263#_M1004_g N_VPWR_M1004_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.28035 AS=0.3402 PD=1.705 PS=1.8 NRD=13.2778 NRS=28.9196 M=1
+ R=8.4 SA=75002.3 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1015 N_A_110_263#_M1015_d N_A_454_263#_M1015_g N_VPWR_M1004_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3402 PD=3.05 PS=1.8 NRD=0 NRS=11.7215 M=1 R=8.4
+ SA=75003 SB=75000.2 A=0.189 P=2.82 MULT=1
DX36_noxref VNB VPB NWDIODE A=19.5079 P=24.65
c_109 VNB 0 5.91746e-20 $X=0 $Y=0
c_188 VPB 0 2.95893e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__ha_4.pxi.spice"
*
.ends
*
*
