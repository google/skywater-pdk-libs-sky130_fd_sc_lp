* File: sky130_fd_sc_lp__sdlclkp_2.pxi.spice
* Created: Fri Aug 28 11:31:30 2020
* 
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%SCE N_SCE_c_168_n N_SCE_M1005_g N_SCE_M1021_g
+ N_SCE_c_170_n SCE SCE SCE SCE N_SCE_c_172_n N_SCE_c_173_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%SCE
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%GATE N_GATE_M1017_g N_GATE_M1010_g
+ N_GATE_c_196_n N_GATE_c_201_n GATE N_GATE_c_198_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%GATE
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%A_282_70# N_A_282_70#_M1020_d
+ N_A_282_70#_M1007_d N_A_282_70#_c_240_n N_A_282_70#_c_250_n
+ N_A_282_70#_M1002_g N_A_282_70#_M1015_g N_A_282_70#_c_242_n
+ N_A_282_70#_c_243_n N_A_282_70#_c_244_n N_A_282_70#_c_245_n
+ N_A_282_70#_c_246_n N_A_282_70#_c_255_n N_A_282_70#_c_247_n
+ N_A_282_70#_c_256_n N_A_282_70#_c_248_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%A_282_70#
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%A_250_443# N_A_250_443#_M1023_s
+ N_A_250_443#_M1003_s N_A_250_443#_c_327_n N_A_250_443#_c_317_n
+ N_A_250_443#_M1020_g N_A_250_443#_c_328_n N_A_250_443#_c_329_n
+ N_A_250_443#_c_318_n N_A_250_443#_M1007_g N_A_250_443#_c_320_n
+ N_A_250_443#_c_321_n N_A_250_443#_c_322_n N_A_250_443#_M1014_g
+ N_A_250_443#_M1018_g N_A_250_443#_c_333_n N_A_250_443#_c_323_n
+ N_A_250_443#_c_324_n N_A_250_443#_c_363_n N_A_250_443#_c_325_n
+ N_A_250_443#_c_326_n N_A_250_443#_c_335_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%A_250_443#
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%A_742_107# N_A_742_107#_M1016_d
+ N_A_742_107#_M1019_d N_A_742_107#_M1013_g N_A_742_107#_M1011_g
+ N_A_742_107#_M1008_g N_A_742_107#_c_449_n N_A_742_107#_c_450_n
+ N_A_742_107#_M1000_g N_A_742_107#_c_458_n N_A_742_107#_c_459_n
+ N_A_742_107#_c_451_n N_A_742_107#_c_460_n N_A_742_107#_c_461_n
+ N_A_742_107#_c_452_n N_A_742_107#_c_463_n N_A_742_107#_c_464_n
+ N_A_742_107#_c_465_n N_A_742_107#_c_466_n N_A_742_107#_c_516_p
+ N_A_742_107#_c_453_n N_A_742_107#_c_454_n N_A_742_107#_c_469_n
+ N_A_742_107#_c_470_n N_A_742_107#_c_455_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%A_742_107#
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%A_614_133# N_A_614_133#_M1014_d
+ N_A_614_133#_M1002_d N_A_614_133#_M1016_g N_A_614_133#_M1019_g
+ N_A_614_133#_c_588_n N_A_614_133#_c_589_n N_A_614_133#_c_590_n
+ N_A_614_133#_c_591_n N_A_614_133#_c_592_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%A_614_133#
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%CLK N_CLK_c_649_n N_CLK_M1023_g N_CLK_c_650_n
+ N_CLK_M1003_g N_CLK_c_651_n N_CLK_M1006_g N_CLK_c_656_n N_CLK_M1022_g CLK CLK
+ CLK CLK PM_SKY130_FD_SC_LP__SDLCLKP_2%CLK
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%A_1235_429# N_A_1235_429#_M1008_d
+ N_A_1235_429#_M1022_d N_A_1235_429#_M1001_g N_A_1235_429#_M1004_g
+ N_A_1235_429#_M1012_g N_A_1235_429#_M1009_g N_A_1235_429#_c_719_n
+ N_A_1235_429#_c_720_n N_A_1235_429#_c_729_n N_A_1235_429#_c_721_n
+ N_A_1235_429#_c_722_n N_A_1235_429#_c_723_n N_A_1235_429#_c_731_n
+ N_A_1235_429#_c_724_n N_A_1235_429#_c_725_n N_A_1235_429#_c_733_n
+ N_A_1235_429#_c_767_p N_A_1235_429#_c_726_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%A_1235_429#
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%VPWR N_VPWR_M1021_s N_VPWR_M1007_s
+ N_VPWR_M1011_d N_VPWR_M1003_d N_VPWR_M1000_d N_VPWR_M1009_d N_VPWR_c_814_n
+ N_VPWR_c_815_n N_VPWR_c_816_n N_VPWR_c_817_n N_VPWR_c_818_n N_VPWR_c_819_n
+ N_VPWR_c_820_n N_VPWR_c_821_n N_VPWR_c_822_n N_VPWR_c_823_n VPWR
+ N_VPWR_c_824_n N_VPWR_c_825_n N_VPWR_c_826_n N_VPWR_c_827_n N_VPWR_c_828_n
+ N_VPWR_c_829_n N_VPWR_c_830_n N_VPWR_c_813_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%VPWR
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%A_110_70# N_A_110_70#_M1005_d
+ N_A_110_70#_M1014_s N_A_110_70#_M1017_d N_A_110_70#_M1002_s
+ N_A_110_70#_c_913_n N_A_110_70#_c_918_n N_A_110_70#_c_992_p
+ N_A_110_70#_c_919_n N_A_110_70#_c_920_n N_A_110_70#_c_921_n
+ N_A_110_70#_c_922_n N_A_110_70#_c_923_n N_A_110_70#_c_914_n
+ N_A_110_70#_c_924_n N_A_110_70#_c_915_n N_A_110_70#_c_925_n
+ N_A_110_70#_c_916_n PM_SKY130_FD_SC_LP__SDLCLKP_2%A_110_70#
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%GCLK N_GCLK_M1001_s N_GCLK_M1004_s
+ N_GCLK_c_998_n GCLK GCLK GCLK GCLK N_GCLK_c_995_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%GCLK
x_PM_SKY130_FD_SC_LP__SDLCLKP_2%VGND N_VGND_M1005_s N_VGND_M1010_d
+ N_VGND_M1013_d N_VGND_M1023_d N_VGND_M1001_d N_VGND_M1012_d N_VGND_c_1015_n
+ N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n
+ N_VGND_c_1020_n N_VGND_c_1021_n VGND N_VGND_c_1022_n N_VGND_c_1023_n
+ N_VGND_c_1024_n N_VGND_c_1025_n N_VGND_c_1026_n N_VGND_c_1027_n
+ N_VGND_c_1028_n N_VGND_c_1029_n N_VGND_c_1030_n N_VGND_c_1031_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_2%VGND
cc_1 VNB N_SCE_c_168_n 0.0246172f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.353
cc_2 VNB N_SCE_M1021_g 0.00659088f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_3 VNB N_SCE_c_170_n 0.0246924f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.55
cc_4 VNB SCE 0.0332865f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_SCE_c_172_n 0.0246924f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_6 VNB N_SCE_c_173_n 0.0212493f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_7 VNB N_GATE_M1010_g 0.0421666f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_8 VNB N_GATE_c_196_n 0.0118339f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_9 VNB GATE 0.00422564f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_GATE_c_198_n 0.0195022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_282_70#_c_240_n 0.0173511f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_12 VNB N_A_282_70#_M1015_g 0.0326363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_282_70#_c_242_n 0.00333718f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.045
cc_14 VNB N_A_282_70#_c_243_n 0.0082903f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_15 VNB N_A_282_70#_c_244_n 0.00497581f $X=-0.19 $Y=-0.245 $X2=0.25 $Y2=1.295
cc_16 VNB N_A_282_70#_c_245_n 0.0024144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_282_70#_c_246_n 0.00674704f $X=-0.19 $Y=-0.245 $X2=0.25 $Y2=2.035
cc_18 VNB N_A_282_70#_c_247_n 0.00263764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_282_70#_c_248_n 0.00148566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_250_443#_c_317_n 0.0190861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_250_443#_c_318_n 0.014984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_250_443#_M1007_g 0.0185894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_250_443#_c_320_n 0.0423928f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_24 VNB N_A_250_443#_c_321_n 0.0886184f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_25 VNB N_A_250_443#_c_322_n 0.0173683f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_26 VNB N_A_250_443#_c_323_n 0.0356084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_250_443#_c_324_n 0.0172136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_250_443#_c_325_n 0.0788146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_250_443#_c_326_n 0.00686595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_742_107#_M1013_g 0.0365089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_742_107#_M1008_g 0.0453384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_742_107#_c_449_n 0.0267338f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.045
cc_33 VNB N_A_742_107#_c_450_n 0.00820386f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_34 VNB N_A_742_107#_c_451_n 0.00392934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_742_107#_c_452_n 0.0115728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_742_107#_c_453_n 0.0164939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_742_107#_c_454_n 0.00172515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_742_107#_c_455_n 0.0117672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_614_133#_M1016_g 0.0249367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_614_133#_M1019_g 0.00564691f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_41 VNB N_A_614_133#_c_588_n 0.0049002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_614_133#_c_589_n 0.0195891f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.045
cc_43 VNB N_A_614_133#_c_590_n 0.00522796f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_44 VNB N_A_614_133#_c_591_n 0.00259157f $X=-0.19 $Y=-0.245 $X2=0.25 $Y2=1.045
cc_45 VNB N_A_614_133#_c_592_n 0.0384935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_CLK_c_649_n 0.0203505f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.077
cc_47 VNB N_CLK_c_650_n 0.0883915f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.56
cc_48 VNB N_CLK_c_651_n 0.0159318f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_49 VNB CLK 0.00249465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB CLK 7.81659e-19 $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.045
cc_51 VNB N_A_1235_429#_M1001_g 0.0223327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1235_429#_M1004_g 0.0119199f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_53 VNB N_A_1235_429#_M1012_g 0.026336f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.045
cc_54 VNB N_A_1235_429#_M1009_g 0.00146273f $X=-0.19 $Y=-0.245 $X2=0.25
+ $Y2=0.925
cc_55 VNB N_A_1235_429#_c_719_n 0.00615236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1235_429#_c_720_n 0.00870159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1235_429#_c_721_n 0.021736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1235_429#_c_722_n 0.00302211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1235_429#_c_723_n 0.010215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1235_429#_c_724_n 0.00367846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1235_429#_c_725_n 0.0546734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1235_429#_c_726_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VPWR_c_813_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_110_70#_c_913_n 0.0138121f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_65 VNB N_A_110_70#_c_914_n 0.00645625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_110_70#_c_915_n 0.00504204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_110_70#_c_916_n 0.00700864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_GCLK_c_995_n 0.00448819f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_69 VNB N_VGND_c_1015_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.045
cc_70 VNB N_VGND_c_1016_n 0.0210568f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_71 VNB N_VGND_c_1017_n 0.0077039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1018_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.25 $Y2=1.665
cc_73 VNB N_VGND_c_1019_n 0.0119025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1020_n 0.010867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1021_n 0.0400851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1022_n 0.015986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1023_n 0.0700555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1024_n 0.0309833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1025_n 0.0326772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1026_n 0.0159186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1027_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1028_n 0.0155415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1029_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1030_n 0.00548198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1031_n 0.453021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VPB N_SCE_M1021_g 0.0578891f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_87 VPB SCE 0.0242081f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_88 VPB N_GATE_M1017_g 0.0302261f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.88
cc_89 VPB N_GATE_c_196_n 0.0116275f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_90 VPB N_GATE_c_201_n 0.0221293f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_91 VPB GATE 0.00320904f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_92 VPB N_A_282_70#_c_240_n 0.0207148f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_93 VPB N_A_282_70#_c_250_n 0.0302548f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_282_70#_M1002_g 0.0196876f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_95 VPB N_A_282_70#_c_242_n 0.0213147f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.045
cc_96 VPB N_A_282_70#_c_243_n 0.0255264f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=0.88
cc_97 VPB N_A_282_70#_c_246_n 0.00772548f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=2.035
cc_98 VPB N_A_282_70#_c_255_n 0.00146324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_282_70#_c_256_n 0.00407786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_250_443#_c_327_n 0.0428344f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_101 VPB N_A_250_443#_c_328_n 0.166173f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_102 VPB N_A_250_443#_c_329_n 0.0120281f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_103 VPB N_A_250_443#_c_318_n 0.0300935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_250_443#_M1007_g 0.0320996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_250_443#_M1018_g 0.0372066f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=1.295
cc_106 VPB N_A_250_443#_c_333_n 0.0218936f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=2.035
cc_107 VPB N_A_250_443#_c_324_n 0.0102978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_250_443#_c_335_n 0.0074123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_742_107#_M1011_g 0.032868f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_110 VPB N_A_742_107#_M1000_g 0.0206674f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=0.925
cc_111 VPB N_A_742_107#_c_458_n 0.0160555f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=1.295
cc_112 VPB N_A_742_107#_c_459_n 0.0057895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_742_107#_c_460_n 0.00605531f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_742_107#_c_461_n 0.00946291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_742_107#_c_452_n 0.00202204f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_742_107#_c_463_n 0.0101736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_742_107#_c_464_n 0.00459832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_742_107#_c_465_n 0.00752036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_742_107#_c_466_n 4.76509e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_742_107#_c_453_n 0.0120403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_742_107#_c_454_n 0.0079859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_742_107#_c_469_n 0.00449408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_742_107#_c_470_n 0.00100392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_742_107#_c_455_n 0.0276974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_614_133#_M1019_g 0.0259215f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_126 VPB N_A_614_133#_c_588_n 0.0142377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_CLK_c_650_n 0.0227859f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.56
cc_128 VPB N_CLK_M1003_g 0.0310168f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.55
cc_129 VPB N_CLK_c_656_n 0.0210942f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_130 VPB N_CLK_M1022_g 0.0270945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB CLK 0.00183829f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.045
cc_132 VPB N_A_1235_429#_M1004_g 0.0227093f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_133 VPB N_A_1235_429#_M1009_g 0.0215064f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=0.925
cc_134 VPB N_A_1235_429#_c_729_n 0.00702341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_1235_429#_c_723_n 0.00365619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_1235_429#_c_731_n 0.00754068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_1235_429#_c_724_n 0.0220992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_1235_429#_c_733_n 0.00464331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_814_n 0.011036f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.045
cc_140 VPB N_VPWR_c_815_n 0.0368315f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.045
cc_141 VPB N_VPWR_c_816_n 0.00978075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_817_n 0.00830399f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=1.665
cc_143 VPB N_VPWR_c_818_n 0.0158333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_819_n 0.00722481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_820_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_821_n 0.0237814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_822_n 0.0298521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_823_n 0.00631381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_824_n 0.02701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_825_n 0.0587231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_826_n 0.0178619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_827_n 0.0147084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_828_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_829_n 0.00739624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_830_n 0.010398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_813_n 0.0810883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_110_70#_c_913_n 0.00831407f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_158 VPB N_A_110_70#_c_918_n 0.00984158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_110_70#_c_919_n 0.00754362f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=0.925
cc_160 VPB N_A_110_70#_c_920_n 0.00257876f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=1.045
cc_161 VPB N_A_110_70#_c_921_n 0.02643f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=1.295
cc_162 VPB N_A_110_70#_c_922_n 0.00225021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_110_70#_c_923_n 0.00958824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_110_70#_c_924_n 0.00413504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_110_70#_c_925_n 0.00347489f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_110_70#_c_916_n 0.00668545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_GCLK_c_995_n 0.0011933f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.045
cc_168 N_SCE_c_173_n N_GATE_M1010_g 0.0155073f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_169 N_SCE_c_170_n N_GATE_c_196_n 0.0155073f $X=0.352 $Y=1.55 $X2=0 $Y2=0
cc_170 N_SCE_M1021_g N_GATE_c_201_n 0.0737804f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_171 N_SCE_c_172_n N_GATE_c_198_n 0.0155073f $X=0.32 $Y=1.045 $X2=0 $Y2=0
cc_172 N_SCE_M1021_g N_VPWR_c_815_n 0.0114952f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_173 SCE N_VPWR_c_815_n 0.0296692f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_174 N_SCE_M1021_g N_VPWR_c_824_n 0.00428763f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_175 N_SCE_M1021_g N_VPWR_c_813_n 0.00829233f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_176 N_SCE_c_168_n N_A_110_70#_c_913_n 0.00598712f $X=0.352 $Y=1.353 $X2=0
+ $Y2=0
cc_177 N_SCE_M1021_g N_A_110_70#_c_918_n 0.00226923f $X=0.475 $Y=2.66 $X2=0
+ $Y2=0
cc_178 SCE N_A_110_70#_c_914_n 0.099175f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_179 N_SCE_c_173_n N_A_110_70#_c_914_n 0.00598712f $X=0.352 $Y=0.88 $X2=0
+ $Y2=0
cc_180 N_SCE_M1021_g N_A_110_70#_c_924_n 0.00522433f $X=0.475 $Y=2.66 $X2=0
+ $Y2=0
cc_181 SCE N_VGND_c_1016_n 0.0258736f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_182 N_SCE_c_172_n N_VGND_c_1016_n 0.00156152f $X=0.32 $Y=1.045 $X2=0 $Y2=0
cc_183 N_SCE_c_173_n N_VGND_c_1016_n 0.00962719f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_184 N_SCE_c_173_n N_VGND_c_1022_n 0.00396895f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_185 SCE N_VGND_c_1031_n 0.00154673f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_186 N_SCE_c_173_n N_VGND_c_1031_n 0.00771726f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_187 N_GATE_M1010_g N_A_282_70#_c_244_n 4.30318e-19 $X=0.905 $Y=0.56 $X2=0
+ $Y2=0
cc_188 N_GATE_M1010_g N_A_282_70#_c_245_n 9.0643e-19 $X=0.905 $Y=0.56 $X2=0
+ $Y2=0
cc_189 GATE N_A_282_70#_c_245_n 0.0218463f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_190 N_GATE_c_198_n N_A_282_70#_c_245_n 2.5466e-19 $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_191 N_GATE_c_196_n N_A_282_70#_c_255_n 2.98651e-19 $X=0.972 $Y=1.825 $X2=0
+ $Y2=0
cc_192 GATE N_A_282_70#_c_255_n 0.0281797f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_193 N_GATE_M1010_g N_A_282_70#_c_248_n 7.72756e-19 $X=0.905 $Y=0.56 $X2=0
+ $Y2=0
cc_194 N_GATE_M1010_g N_A_250_443#_c_317_n 0.0176135f $X=0.905 $Y=0.56 $X2=0
+ $Y2=0
cc_195 N_GATE_M1017_g N_A_250_443#_c_318_n 0.00550254f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_196 N_GATE_c_196_n N_A_250_443#_c_318_n 0.016234f $X=0.972 $Y=1.825 $X2=0
+ $Y2=0
cc_197 N_GATE_M1010_g N_A_250_443#_c_321_n 0.00687969f $X=0.905 $Y=0.56 $X2=0
+ $Y2=0
cc_198 GATE N_A_250_443#_c_321_n 0.00773516f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_199 N_GATE_c_198_n N_A_250_443#_c_321_n 0.016234f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_200 N_GATE_M1017_g N_A_250_443#_c_333_n 0.0177954f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_201 GATE N_A_250_443#_c_333_n 4.39988e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_202 N_GATE_M1017_g N_VPWR_c_815_n 0.00116793f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_203 N_GATE_M1017_g N_VPWR_c_824_n 0.0030129f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_204 N_GATE_M1017_g N_VPWR_c_813_n 0.00394334f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_205 N_GATE_M1010_g N_A_110_70#_c_913_n 0.0105507f $X=0.905 $Y=0.56 $X2=0
+ $Y2=0
cc_206 N_GATE_c_201_n N_A_110_70#_c_913_n 0.00577749f $X=0.972 $Y=1.975 $X2=0
+ $Y2=0
cc_207 GATE N_A_110_70#_c_913_n 0.0510174f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_208 N_GATE_M1017_g N_A_110_70#_c_918_n 0.0148115f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_209 GATE N_A_110_70#_c_919_n 0.00773076f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_210 N_GATE_M1010_g N_A_110_70#_c_914_n 0.00232933f $X=0.905 $Y=0.56 $X2=0
+ $Y2=0
cc_211 N_GATE_M1017_g N_A_110_70#_c_924_n 0.0134646f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_212 N_GATE_c_201_n N_A_110_70#_c_924_n 0.00763117f $X=0.972 $Y=1.975 $X2=0
+ $Y2=0
cc_213 GATE N_A_110_70#_c_924_n 0.0237764f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_214 N_GATE_M1010_g N_VGND_c_1016_n 5.44985e-19 $X=0.905 $Y=0.56 $X2=0 $Y2=0
cc_215 N_GATE_M1010_g N_VGND_c_1017_n 0.0018259f $X=0.905 $Y=0.56 $X2=0 $Y2=0
cc_216 GATE N_VGND_c_1017_n 0.00719213f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_217 N_GATE_c_198_n N_VGND_c_1017_n 0.00366473f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_218 N_GATE_M1010_g N_VGND_c_1022_n 0.00478016f $X=0.905 $Y=0.56 $X2=0 $Y2=0
cc_219 N_GATE_M1010_g N_VGND_c_1031_n 0.009365f $X=0.905 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A_282_70#_c_244_n N_A_250_443#_c_317_n 0.00202061f $X=1.55 $Y=0.56
+ $X2=0 $Y2=0
cc_221 N_A_282_70#_M1002_g N_A_250_443#_c_328_n 0.00907339f $X=3.225 $Y=2.495
+ $X2=0 $Y2=0
cc_222 N_A_282_70#_c_245_n N_A_250_443#_c_318_n 0.00543061f $X=1.6 $Y=1.585
+ $X2=0 $Y2=0
cc_223 N_A_282_70#_c_255_n N_A_250_443#_c_318_n 0.0110276f $X=1.715 $Y=1.75
+ $X2=0 $Y2=0
cc_224 N_A_282_70#_c_242_n N_A_250_443#_M1007_g 0.00292589f $X=2.695 $Y=1.66
+ $X2=0 $Y2=0
cc_225 N_A_282_70#_c_243_n N_A_250_443#_M1007_g 0.0214229f $X=2.62 $Y=1.75 $X2=0
+ $Y2=0
cc_226 N_A_282_70#_c_245_n N_A_250_443#_M1007_g 0.00522472f $X=1.6 $Y=1.585
+ $X2=0 $Y2=0
cc_227 N_A_282_70#_c_246_n N_A_250_443#_M1007_g 0.0217557f $X=2.305 $Y=1.75
+ $X2=0 $Y2=0
cc_228 N_A_282_70#_c_256_n N_A_250_443#_M1007_g 0.00924201f $X=2.39 $Y=2.21
+ $X2=0 $Y2=0
cc_229 N_A_282_70#_c_243_n N_A_250_443#_c_320_n 0.0461415f $X=2.62 $Y=1.75 $X2=0
+ $Y2=0
cc_230 N_A_282_70#_c_246_n N_A_250_443#_c_320_n 2.98923e-19 $X=2.305 $Y=1.75
+ $X2=0 $Y2=0
cc_231 N_A_282_70#_c_247_n N_A_250_443#_c_320_n 0.00143385f $X=2.415 $Y=1.915
+ $X2=0 $Y2=0
cc_232 N_A_282_70#_c_244_n N_A_250_443#_c_321_n 0.0135109f $X=1.55 $Y=0.56 $X2=0
+ $Y2=0
cc_233 N_A_282_70#_c_245_n N_A_250_443#_c_321_n 0.0187578f $X=1.6 $Y=1.585 $X2=0
+ $Y2=0
cc_234 N_A_282_70#_c_246_n N_A_250_443#_c_321_n 0.0125032f $X=2.305 $Y=1.75
+ $X2=0 $Y2=0
cc_235 N_A_282_70#_c_248_n N_A_250_443#_c_321_n 0.0150946f $X=1.567 $Y=1.125
+ $X2=0 $Y2=0
cc_236 N_A_282_70#_M1015_g N_A_250_443#_c_322_n 0.0219938f $X=3.425 $Y=0.875
+ $X2=0 $Y2=0
cc_237 N_A_282_70#_M1002_g N_A_250_443#_M1018_g 0.0117752f $X=3.225 $Y=2.495
+ $X2=0 $Y2=0
cc_238 N_A_282_70#_M1015_g N_A_250_443#_c_323_n 0.00966652f $X=3.425 $Y=0.875
+ $X2=0 $Y2=0
cc_239 N_A_282_70#_c_244_n N_A_250_443#_c_363_n 0.0331933f $X=1.55 $Y=0.56 $X2=0
+ $Y2=0
cc_240 N_A_282_70#_c_244_n N_A_250_443#_c_325_n 0.00474252f $X=1.55 $Y=0.56
+ $X2=0 $Y2=0
cc_241 N_A_282_70#_M1015_g N_A_742_107#_M1013_g 0.0371238f $X=3.425 $Y=0.875
+ $X2=0 $Y2=0
cc_242 N_A_282_70#_c_250_n N_A_742_107#_M1011_g 0.0020815f $X=3.15 $Y=2.05 $X2=0
+ $Y2=0
cc_243 N_A_282_70#_c_240_n N_A_742_107#_c_455_n 0.0371238f $X=3.35 $Y=1.66 $X2=0
+ $Y2=0
cc_244 N_A_282_70#_c_240_n N_A_614_133#_c_588_n 0.0124791f $X=3.35 $Y=1.66 $X2=0
+ $Y2=0
cc_245 N_A_282_70#_c_250_n N_A_614_133#_c_588_n 0.00521158f $X=3.15 $Y=2.05
+ $X2=0 $Y2=0
cc_246 N_A_282_70#_M1015_g N_A_614_133#_c_588_n 0.00594538f $X=3.425 $Y=0.875
+ $X2=0 $Y2=0
cc_247 N_A_282_70#_c_242_n N_A_614_133#_c_588_n 3.01255e-19 $X=2.695 $Y=1.66
+ $X2=0 $Y2=0
cc_248 N_A_282_70#_M1015_g N_A_614_133#_c_589_n 2.90519e-19 $X=3.425 $Y=0.875
+ $X2=0 $Y2=0
cc_249 N_A_282_70#_c_240_n N_A_614_133#_c_590_n 0.00967568f $X=3.35 $Y=1.66
+ $X2=0 $Y2=0
cc_250 N_A_282_70#_M1015_g N_A_614_133#_c_590_n 0.0150397f $X=3.425 $Y=0.875
+ $X2=0 $Y2=0
cc_251 N_A_282_70#_M1002_g N_VPWR_c_813_n 9.49986e-19 $X=3.225 $Y=2.495 $X2=0
+ $Y2=0
cc_252 N_A_282_70#_c_244_n N_A_110_70#_c_913_n 0.00542138f $X=1.55 $Y=0.56 $X2=0
+ $Y2=0
cc_253 N_A_282_70#_M1007_d N_A_110_70#_c_919_n 0.00218945f $X=2.055 $Y=2.085
+ $X2=0 $Y2=0
cc_254 N_A_282_70#_c_246_n N_A_110_70#_c_919_n 0.0213737f $X=2.305 $Y=1.75 $X2=0
+ $Y2=0
cc_255 N_A_282_70#_c_255_n N_A_110_70#_c_919_n 0.0138953f $X=1.715 $Y=1.75 $X2=0
+ $Y2=0
cc_256 N_A_282_70#_c_256_n N_A_110_70#_c_919_n 0.0140751f $X=2.39 $Y=2.21 $X2=0
+ $Y2=0
cc_257 N_A_282_70#_M1007_d N_A_110_70#_c_920_n 0.00414523f $X=2.055 $Y=2.085
+ $X2=0 $Y2=0
cc_258 N_A_282_70#_c_256_n N_A_110_70#_c_920_n 0.0288484f $X=2.39 $Y=2.21 $X2=0
+ $Y2=0
cc_259 N_A_282_70#_c_256_n N_A_110_70#_c_921_n 0.0169185f $X=2.39 $Y=2.21 $X2=0
+ $Y2=0
cc_260 N_A_282_70#_M1002_g N_A_110_70#_c_923_n 0.00630067f $X=3.225 $Y=2.495
+ $X2=0 $Y2=0
cc_261 N_A_282_70#_c_244_n N_A_110_70#_c_914_n 0.005047f $X=1.55 $Y=0.56 $X2=0
+ $Y2=0
cc_262 N_A_282_70#_c_250_n N_A_110_70#_c_925_n 0.00974585f $X=3.15 $Y=2.05 $X2=0
+ $Y2=0
cc_263 N_A_282_70#_c_240_n N_A_110_70#_c_916_n 0.00668939f $X=3.35 $Y=1.66 $X2=0
+ $Y2=0
cc_264 N_A_282_70#_c_250_n N_A_110_70#_c_916_n 0.00762016f $X=3.15 $Y=2.05 $X2=0
+ $Y2=0
cc_265 N_A_282_70#_M1002_g N_A_110_70#_c_916_n 0.00334391f $X=3.225 $Y=2.495
+ $X2=0 $Y2=0
cc_266 N_A_282_70#_M1015_g N_A_110_70#_c_916_n 0.00128961f $X=3.425 $Y=0.875
+ $X2=0 $Y2=0
cc_267 N_A_282_70#_c_242_n N_A_110_70#_c_916_n 0.0131499f $X=2.695 $Y=1.66 $X2=0
+ $Y2=0
cc_268 N_A_282_70#_c_247_n N_A_110_70#_c_916_n 0.0251378f $X=2.415 $Y=1.915
+ $X2=0 $Y2=0
cc_269 N_A_282_70#_c_256_n N_A_110_70#_c_916_n 0.0627312f $X=2.39 $Y=2.21 $X2=0
+ $Y2=0
cc_270 N_A_282_70#_M1015_g N_VGND_c_1023_n 6.65218e-19 $X=3.425 $Y=0.875 $X2=0
+ $Y2=0
cc_271 N_A_282_70#_c_244_n N_VGND_c_1023_n 0.00999441f $X=1.55 $Y=0.56 $X2=0
+ $Y2=0
cc_272 N_A_282_70#_c_244_n N_VGND_c_1031_n 0.0105228f $X=1.55 $Y=0.56 $X2=0
+ $Y2=0
cc_273 N_A_250_443#_c_323_n N_A_742_107#_M1016_d 0.00666521f $X=4.985 $Y=0.61
+ $X2=-0.19 $Y2=-0.245
cc_274 N_A_250_443#_c_323_n N_A_742_107#_M1013_g 0.0121865f $X=4.985 $Y=0.61
+ $X2=0 $Y2=0
cc_275 N_A_250_443#_M1018_g N_A_742_107#_M1011_g 0.0395013f $X=3.655 $Y=2.495
+ $X2=0 $Y2=0
cc_276 N_A_250_443#_c_323_n N_A_742_107#_c_451_n 0.0319609f $X=4.985 $Y=0.61
+ $X2=0 $Y2=0
cc_277 N_A_250_443#_c_324_n N_A_742_107#_c_451_n 0.0156181f $X=5.157 $Y=2.115
+ $X2=0 $Y2=0
cc_278 N_A_250_443#_c_324_n N_A_742_107#_c_460_n 0.0154584f $X=5.157 $Y=2.115
+ $X2=0 $Y2=0
cc_279 N_A_250_443#_c_335_n N_A_742_107#_c_460_n 0.0205221f $X=5.295 $Y=2.28
+ $X2=0 $Y2=0
cc_280 N_A_250_443#_c_324_n N_A_742_107#_c_452_n 0.0519953f $X=5.157 $Y=2.115
+ $X2=0 $Y2=0
cc_281 N_A_250_443#_M1003_s N_A_742_107#_c_463_n 0.0073298f $X=5.15 $Y=2.145
+ $X2=0 $Y2=0
cc_282 N_A_250_443#_c_335_n N_A_742_107#_c_463_n 0.0249289f $X=5.295 $Y=2.28
+ $X2=0 $Y2=0
cc_283 N_A_250_443#_c_324_n N_A_742_107#_c_464_n 0.0070373f $X=5.157 $Y=2.115
+ $X2=0 $Y2=0
cc_284 N_A_250_443#_c_335_n N_A_742_107#_c_464_n 0.0113465f $X=5.295 $Y=2.28
+ $X2=0 $Y2=0
cc_285 N_A_250_443#_c_324_n N_A_742_107#_c_466_n 0.00270645f $X=5.157 $Y=2.115
+ $X2=0 $Y2=0
cc_286 N_A_250_443#_c_324_n N_A_742_107#_c_469_n 0.0143864f $X=5.157 $Y=2.115
+ $X2=0 $Y2=0
cc_287 N_A_250_443#_M1018_g N_A_742_107#_c_455_n 0.00123997f $X=3.655 $Y=2.495
+ $X2=0 $Y2=0
cc_288 N_A_250_443#_c_323_n N_A_614_133#_M1014_d 0.00176461f $X=4.985 $Y=0.61
+ $X2=-0.19 $Y2=-0.245
cc_289 N_A_250_443#_c_323_n N_A_614_133#_M1016_g 0.015407f $X=4.985 $Y=0.61
+ $X2=0 $Y2=0
cc_290 N_A_250_443#_c_324_n N_A_614_133#_M1016_g 0.00248798f $X=5.157 $Y=2.115
+ $X2=0 $Y2=0
cc_291 N_A_250_443#_c_326_n N_A_614_133#_M1016_g 0.00432922f $X=5.15 $Y=0.53
+ $X2=0 $Y2=0
cc_292 N_A_250_443#_c_324_n N_A_614_133#_M1019_g 6.76381e-19 $X=5.157 $Y=2.115
+ $X2=0 $Y2=0
cc_293 N_A_250_443#_c_328_n N_A_614_133#_c_588_n 0.00316032f $X=3.58 $Y=3.15
+ $X2=0 $Y2=0
cc_294 N_A_250_443#_M1018_g N_A_614_133#_c_588_n 0.00163989f $X=3.655 $Y=2.495
+ $X2=0 $Y2=0
cc_295 N_A_250_443#_c_323_n N_A_614_133#_c_589_n 0.0209585f $X=4.985 $Y=0.61
+ $X2=0 $Y2=0
cc_296 N_A_250_443#_c_320_n N_A_614_133#_c_590_n 0.00443547f $X=2.92 $Y=1.27
+ $X2=0 $Y2=0
cc_297 N_A_250_443#_c_322_n N_A_614_133#_c_590_n 0.00518912f $X=2.995 $Y=1.195
+ $X2=0 $Y2=0
cc_298 N_A_250_443#_c_323_n N_A_614_133#_c_590_n 0.0257281f $X=4.985 $Y=0.61
+ $X2=0 $Y2=0
cc_299 N_A_250_443#_c_323_n N_A_614_133#_c_591_n 0.00349812f $X=4.985 $Y=0.61
+ $X2=0 $Y2=0
cc_300 N_A_250_443#_c_326_n N_CLK_c_649_n 0.00958755f $X=5.15 $Y=0.53 $X2=-0.19
+ $Y2=-0.245
cc_301 N_A_250_443#_c_324_n N_CLK_c_650_n 0.0178434f $X=5.157 $Y=2.115 $X2=0
+ $Y2=0
cc_302 N_A_250_443#_c_335_n N_CLK_c_650_n 0.00372409f $X=5.295 $Y=2.28 $X2=0
+ $Y2=0
cc_303 N_A_250_443#_c_335_n N_CLK_M1003_g 0.00486941f $X=5.295 $Y=2.28 $X2=0
+ $Y2=0
cc_304 N_A_250_443#_c_324_n CLK 0.0408403f $X=5.157 $Y=2.115 $X2=0 $Y2=0
cc_305 N_A_250_443#_c_324_n CLK 0.0346169f $X=5.157 $Y=2.115 $X2=0 $Y2=0
cc_306 N_A_250_443#_c_335_n CLK 0.00250181f $X=5.295 $Y=2.28 $X2=0 $Y2=0
cc_307 N_A_250_443#_c_327_n N_VPWR_c_816_n 0.0106222f $X=1.325 $Y=3.075 $X2=0
+ $Y2=0
cc_308 N_A_250_443#_c_328_n N_VPWR_c_816_n 0.0242353f $X=3.58 $Y=3.15 $X2=0
+ $Y2=0
cc_309 N_A_250_443#_M1007_g N_VPWR_c_816_n 0.00318265f $X=1.98 $Y=2.405 $X2=0
+ $Y2=0
cc_310 N_A_250_443#_c_333_n N_VPWR_c_816_n 0.00195343f $X=1.505 $Y=2.29 $X2=0
+ $Y2=0
cc_311 N_A_250_443#_M1018_g N_VPWR_c_817_n 0.0141228f $X=3.655 $Y=2.495 $X2=0
+ $Y2=0
cc_312 N_A_250_443#_c_329_n N_VPWR_c_824_n 0.00835149f $X=1.4 $Y=3.15 $X2=0
+ $Y2=0
cc_313 N_A_250_443#_c_328_n N_VPWR_c_825_n 0.0491138f $X=3.58 $Y=3.15 $X2=0
+ $Y2=0
cc_314 N_A_250_443#_c_328_n N_VPWR_c_813_n 0.0652721f $X=3.58 $Y=3.15 $X2=0
+ $Y2=0
cc_315 N_A_250_443#_c_329_n N_VPWR_c_813_n 0.0112815f $X=1.4 $Y=3.15 $X2=0 $Y2=0
cc_316 N_A_250_443#_M1007_g N_VPWR_c_813_n 3.79764e-19 $X=1.98 $Y=2.405 $X2=0
+ $Y2=0
cc_317 N_A_250_443#_c_323_n N_A_110_70#_M1014_s 0.00324619f $X=4.985 $Y=0.61
+ $X2=0 $Y2=0
cc_318 N_A_250_443#_c_333_n N_A_110_70#_c_918_n 0.0107012f $X=1.505 $Y=2.29
+ $X2=0 $Y2=0
cc_319 N_A_250_443#_c_318_n N_A_110_70#_c_919_n 0.00618176f $X=1.505 $Y=2.215
+ $X2=0 $Y2=0
cc_320 N_A_250_443#_M1007_g N_A_110_70#_c_919_n 0.0123933f $X=1.98 $Y=2.405
+ $X2=0 $Y2=0
cc_321 N_A_250_443#_c_333_n N_A_110_70#_c_919_n 0.0193473f $X=1.505 $Y=2.29
+ $X2=0 $Y2=0
cc_322 N_A_250_443#_c_327_n N_A_110_70#_c_920_n 7.45924e-19 $X=1.325 $Y=3.075
+ $X2=0 $Y2=0
cc_323 N_A_250_443#_M1007_g N_A_110_70#_c_920_n 0.0181643f $X=1.98 $Y=2.405
+ $X2=0 $Y2=0
cc_324 N_A_250_443#_c_328_n N_A_110_70#_c_921_n 0.0239109f $X=3.58 $Y=3.15 $X2=0
+ $Y2=0
cc_325 N_A_250_443#_M1018_g N_A_110_70#_c_921_n 0.00522941f $X=3.655 $Y=2.495
+ $X2=0 $Y2=0
cc_326 N_A_250_443#_c_328_n N_A_110_70#_c_922_n 0.00271057f $X=3.58 $Y=3.15
+ $X2=0 $Y2=0
cc_327 N_A_250_443#_M1018_g N_A_110_70#_c_923_n 0.00201355f $X=3.655 $Y=2.495
+ $X2=0 $Y2=0
cc_328 N_A_250_443#_c_320_n N_A_110_70#_c_915_n 0.00639922f $X=2.92 $Y=1.27
+ $X2=0 $Y2=0
cc_329 N_A_250_443#_c_322_n N_A_110_70#_c_915_n 0.00320233f $X=2.995 $Y=1.195
+ $X2=0 $Y2=0
cc_330 N_A_250_443#_c_323_n N_A_110_70#_c_915_n 0.0250958f $X=4.985 $Y=0.61
+ $X2=0 $Y2=0
cc_331 N_A_250_443#_c_325_n N_A_110_70#_c_915_n 0.00662232f $X=2.07 $Y=0.35
+ $X2=0 $Y2=0
cc_332 N_A_250_443#_M1007_g N_A_110_70#_c_916_n 0.00650766f $X=1.98 $Y=2.405
+ $X2=0 $Y2=0
cc_333 N_A_250_443#_c_320_n N_A_110_70#_c_916_n 0.0154906f $X=2.92 $Y=1.27 $X2=0
+ $Y2=0
cc_334 N_A_250_443#_c_321_n N_A_110_70#_c_916_n 0.00130903f $X=2.235 $Y=1.27
+ $X2=0 $Y2=0
cc_335 N_A_250_443#_c_323_n N_VGND_M1013_d 0.00988631f $X=4.985 $Y=0.61 $X2=0
+ $Y2=0
cc_336 N_A_250_443#_c_317_n N_VGND_c_1017_n 0.00234275f $X=1.335 $Y=0.88 $X2=0
+ $Y2=0
cc_337 N_A_250_443#_c_363_n N_VGND_c_1017_n 0.00314643f $X=2.07 $Y=0.35 $X2=0
+ $Y2=0
cc_338 N_A_250_443#_c_325_n N_VGND_c_1017_n 8.98479e-19 $X=2.07 $Y=0.35 $X2=0
+ $Y2=0
cc_339 N_A_250_443#_c_326_n N_VGND_c_1018_n 0.0116048f $X=5.15 $Y=0.53 $X2=0
+ $Y2=0
cc_340 N_A_250_443#_c_317_n N_VGND_c_1023_n 0.00478016f $X=1.335 $Y=0.88 $X2=0
+ $Y2=0
cc_341 N_A_250_443#_c_322_n N_VGND_c_1023_n 6.65218e-19 $X=2.995 $Y=1.195 $X2=0
+ $Y2=0
cc_342 N_A_250_443#_c_323_n N_VGND_c_1023_n 0.0394473f $X=4.985 $Y=0.61 $X2=0
+ $Y2=0
cc_343 N_A_250_443#_c_363_n N_VGND_c_1023_n 0.0221582f $X=2.07 $Y=0.35 $X2=0
+ $Y2=0
cc_344 N_A_250_443#_c_325_n N_VGND_c_1023_n 0.00680296f $X=2.07 $Y=0.35 $X2=0
+ $Y2=0
cc_345 N_A_250_443#_c_323_n N_VGND_c_1024_n 0.0157373f $X=4.985 $Y=0.61 $X2=0
+ $Y2=0
cc_346 N_A_250_443#_c_326_n N_VGND_c_1024_n 0.0106815f $X=5.15 $Y=0.53 $X2=0
+ $Y2=0
cc_347 N_A_250_443#_c_323_n N_VGND_c_1028_n 0.0240258f $X=4.985 $Y=0.61 $X2=0
+ $Y2=0
cc_348 N_A_250_443#_c_317_n N_VGND_c_1031_n 0.00944862f $X=1.335 $Y=0.88 $X2=0
+ $Y2=0
cc_349 N_A_250_443#_c_321_n N_VGND_c_1031_n 0.00235618f $X=2.235 $Y=1.27 $X2=0
+ $Y2=0
cc_350 N_A_250_443#_c_323_n N_VGND_c_1031_n 0.0763924f $X=4.985 $Y=0.61 $X2=0
+ $Y2=0
cc_351 N_A_250_443#_c_363_n N_VGND_c_1031_n 0.0112098f $X=2.07 $Y=0.35 $X2=0
+ $Y2=0
cc_352 N_A_250_443#_c_325_n N_VGND_c_1031_n 0.010124f $X=2.07 $Y=0.35 $X2=0
+ $Y2=0
cc_353 N_A_250_443#_c_326_n N_VGND_c_1031_n 0.00936924f $X=5.15 $Y=0.53 $X2=0
+ $Y2=0
cc_354 N_A_250_443#_c_323_n A_700_133# 0.00178881f $X=4.985 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_355 N_A_742_107#_M1013_g N_A_614_133#_M1016_g 0.029616f $X=3.785 $Y=0.875
+ $X2=0 $Y2=0
cc_356 N_A_742_107#_c_451_n N_A_614_133#_M1016_g 0.00471008f $X=4.73 $Y=0.96
+ $X2=0 $Y2=0
cc_357 N_A_742_107#_c_452_n N_A_614_133#_M1016_g 0.00469274f $X=4.815 $Y=1.745
+ $X2=0 $Y2=0
cc_358 N_A_742_107#_M1013_g N_A_614_133#_M1019_g 7.25336e-19 $X=3.785 $Y=0.875
+ $X2=0 $Y2=0
cc_359 N_A_742_107#_c_459_n N_A_614_133#_M1019_g 0.0159376f $X=4.66 $Y=1.83
+ $X2=0 $Y2=0
cc_360 N_A_742_107#_c_452_n N_A_614_133#_M1019_g 0.0067255f $X=4.815 $Y=1.745
+ $X2=0 $Y2=0
cc_361 N_A_742_107#_c_454_n N_A_614_133#_M1019_g 9.52288e-19 $X=3.875 $Y=1.75
+ $X2=0 $Y2=0
cc_362 N_A_742_107#_c_455_n N_A_614_133#_M1019_g 0.0259297f $X=4.015 $Y=1.75
+ $X2=0 $Y2=0
cc_363 N_A_742_107#_M1011_g N_A_614_133#_c_588_n 0.0052398f $X=4.015 $Y=2.495
+ $X2=0 $Y2=0
cc_364 N_A_742_107#_c_454_n N_A_614_133#_c_588_n 0.0254403f $X=3.875 $Y=1.75
+ $X2=0 $Y2=0
cc_365 N_A_742_107#_c_455_n N_A_614_133#_c_588_n 0.00456856f $X=4.015 $Y=1.75
+ $X2=0 $Y2=0
cc_366 N_A_742_107#_M1013_g N_A_614_133#_c_589_n 0.0122856f $X=3.785 $Y=0.875
+ $X2=0 $Y2=0
cc_367 N_A_742_107#_c_459_n N_A_614_133#_c_589_n 0.0116866f $X=4.66 $Y=1.83
+ $X2=0 $Y2=0
cc_368 N_A_742_107#_c_454_n N_A_614_133#_c_589_n 0.0218791f $X=3.875 $Y=1.75
+ $X2=0 $Y2=0
cc_369 N_A_742_107#_c_455_n N_A_614_133#_c_589_n 0.00264811f $X=4.015 $Y=1.75
+ $X2=0 $Y2=0
cc_370 N_A_742_107#_M1013_g N_A_614_133#_c_590_n 0.0087665f $X=3.785 $Y=0.875
+ $X2=0 $Y2=0
cc_371 N_A_742_107#_M1013_g N_A_614_133#_c_591_n 0.00100606f $X=3.785 $Y=0.875
+ $X2=0 $Y2=0
cc_372 N_A_742_107#_c_459_n N_A_614_133#_c_591_n 0.017556f $X=4.66 $Y=1.83 $X2=0
+ $Y2=0
cc_373 N_A_742_107#_c_451_n N_A_614_133#_c_591_n 0.0078165f $X=4.73 $Y=0.96
+ $X2=0 $Y2=0
cc_374 N_A_742_107#_c_452_n N_A_614_133#_c_591_n 0.0243553f $X=4.815 $Y=1.745
+ $X2=0 $Y2=0
cc_375 N_A_742_107#_c_459_n N_A_614_133#_c_592_n 0.00166702f $X=4.66 $Y=1.83
+ $X2=0 $Y2=0
cc_376 N_A_742_107#_c_451_n N_A_614_133#_c_592_n 0.00355796f $X=4.73 $Y=0.96
+ $X2=0 $Y2=0
cc_377 N_A_742_107#_c_452_n N_A_614_133#_c_592_n 0.00391125f $X=4.815 $Y=1.745
+ $X2=0 $Y2=0
cc_378 N_A_742_107#_c_450_n N_CLK_c_650_n 0.0383023f $X=6.23 $Y=1.39 $X2=0 $Y2=0
cc_379 N_A_742_107#_c_463_n N_CLK_c_650_n 0.00269068f $X=5.785 $Y=2.62 $X2=0
+ $Y2=0
cc_380 N_A_742_107#_c_466_n N_CLK_c_650_n 0.00916573f $X=5.955 $Y=1.82 $X2=0
+ $Y2=0
cc_381 N_A_742_107#_c_516_p N_CLK_c_650_n 0.00154689f $X=6.55 $Y=1.48 $X2=0
+ $Y2=0
cc_382 N_A_742_107#_c_453_n N_CLK_c_650_n 0.00598369f $X=6.55 $Y=1.48 $X2=0
+ $Y2=0
cc_383 N_A_742_107#_c_460_n N_CLK_M1003_g 0.00350187f $X=4.755 $Y=1.97 $X2=0
+ $Y2=0
cc_384 N_A_742_107#_c_461_n N_CLK_M1003_g 0.00525755f $X=4.755 $Y=2.91 $X2=0
+ $Y2=0
cc_385 N_A_742_107#_c_463_n N_CLK_M1003_g 0.0175236f $X=5.785 $Y=2.62 $X2=0
+ $Y2=0
cc_386 N_A_742_107#_c_464_n N_CLK_M1003_g 0.00792112f $X=5.87 $Y=2.535 $X2=0
+ $Y2=0
cc_387 N_A_742_107#_c_466_n N_CLK_M1003_g 6.26132e-19 $X=5.955 $Y=1.82 $X2=0
+ $Y2=0
cc_388 N_A_742_107#_M1008_g N_CLK_c_651_n 0.0383023f $X=6.155 $Y=0.58 $X2=0
+ $Y2=0
cc_389 N_A_742_107#_c_450_n N_CLK_c_656_n 0.00631921f $X=6.23 $Y=1.39 $X2=0
+ $Y2=0
cc_390 N_A_742_107#_c_465_n N_CLK_c_656_n 0.00928371f $X=6.385 $Y=1.82 $X2=0
+ $Y2=0
cc_391 N_A_742_107#_c_466_n N_CLK_c_656_n 0.00613803f $X=5.955 $Y=1.82 $X2=0
+ $Y2=0
cc_392 N_A_742_107#_c_516_p N_CLK_c_656_n 2.26415e-19 $X=6.55 $Y=1.48 $X2=0
+ $Y2=0
cc_393 N_A_742_107#_c_453_n N_CLK_c_656_n 0.00920603f $X=6.55 $Y=1.48 $X2=0
+ $Y2=0
cc_394 N_A_742_107#_M1000_g N_CLK_M1022_g 0.012839f $X=6.53 $Y=2.465 $X2=0 $Y2=0
cc_395 N_A_742_107#_c_458_n N_CLK_M1022_g 0.00920603f $X=6.55 $Y=1.985 $X2=0
+ $Y2=0
cc_396 N_A_742_107#_c_463_n N_CLK_M1022_g 0.00174334f $X=5.785 $Y=2.62 $X2=0
+ $Y2=0
cc_397 N_A_742_107#_c_464_n N_CLK_M1022_g 0.00844482f $X=5.87 $Y=2.535 $X2=0
+ $Y2=0
cc_398 N_A_742_107#_c_465_n N_CLK_M1022_g 0.00758011f $X=6.385 $Y=1.82 $X2=0
+ $Y2=0
cc_399 N_A_742_107#_M1008_g CLK 0.00203706f $X=6.155 $Y=0.58 $X2=0 $Y2=0
cc_400 N_A_742_107#_c_450_n CLK 3.66915e-19 $X=6.23 $Y=1.39 $X2=0 $Y2=0
cc_401 N_A_742_107#_c_466_n CLK 0.00773955f $X=5.955 $Y=1.82 $X2=0 $Y2=0
cc_402 N_A_742_107#_c_516_p CLK 0.00483746f $X=6.55 $Y=1.48 $X2=0 $Y2=0
cc_403 N_A_742_107#_c_453_n CLK 3.75757e-19 $X=6.55 $Y=1.48 $X2=0 $Y2=0
cc_404 N_A_742_107#_M1000_g N_A_1235_429#_M1004_g 0.0115558f $X=6.53 $Y=2.465
+ $X2=0 $Y2=0
cc_405 N_A_742_107#_c_453_n N_A_1235_429#_M1004_g 0.00667877f $X=6.55 $Y=1.48
+ $X2=0 $Y2=0
cc_406 N_A_742_107#_c_449_n N_A_1235_429#_c_719_n 0.00667877f $X=6.385 $Y=1.39
+ $X2=0 $Y2=0
cc_407 N_A_742_107#_M1008_g N_A_1235_429#_c_720_n 0.0158193f $X=6.155 $Y=0.58
+ $X2=0 $Y2=0
cc_408 N_A_742_107#_M1000_g N_A_1235_429#_c_729_n 0.0187878f $X=6.53 $Y=2.465
+ $X2=0 $Y2=0
cc_409 N_A_742_107#_c_458_n N_A_1235_429#_c_729_n 0.00447389f $X=6.55 $Y=1.985
+ $X2=0 $Y2=0
cc_410 N_A_742_107#_c_465_n N_A_1235_429#_c_729_n 0.0243108f $X=6.385 $Y=1.82
+ $X2=0 $Y2=0
cc_411 N_A_742_107#_c_449_n N_A_1235_429#_c_721_n 0.00511351f $X=6.385 $Y=1.39
+ $X2=0 $Y2=0
cc_412 N_A_742_107#_c_516_p N_A_1235_429#_c_721_n 0.0139643f $X=6.55 $Y=1.48
+ $X2=0 $Y2=0
cc_413 N_A_742_107#_M1008_g N_A_1235_429#_c_722_n 0.00718079f $X=6.155 $Y=0.58
+ $X2=0 $Y2=0
cc_414 N_A_742_107#_c_449_n N_A_1235_429#_c_722_n 0.00866645f $X=6.385 $Y=1.39
+ $X2=0 $Y2=0
cc_415 N_A_742_107#_c_465_n N_A_1235_429#_c_722_n 0.00680672f $X=6.385 $Y=1.82
+ $X2=0 $Y2=0
cc_416 N_A_742_107#_c_516_p N_A_1235_429#_c_722_n 0.0130305f $X=6.55 $Y=1.48
+ $X2=0 $Y2=0
cc_417 N_A_742_107#_M1008_g N_A_1235_429#_c_723_n 0.00209774f $X=6.155 $Y=0.58
+ $X2=0 $Y2=0
cc_418 N_A_742_107#_c_449_n N_A_1235_429#_c_723_n 0.00471364f $X=6.385 $Y=1.39
+ $X2=0 $Y2=0
cc_419 N_A_742_107#_M1000_g N_A_1235_429#_c_723_n 0.00186826f $X=6.53 $Y=2.465
+ $X2=0 $Y2=0
cc_420 N_A_742_107#_c_458_n N_A_1235_429#_c_723_n 0.00192518f $X=6.55 $Y=1.985
+ $X2=0 $Y2=0
cc_421 N_A_742_107#_c_465_n N_A_1235_429#_c_723_n 0.0131148f $X=6.385 $Y=1.82
+ $X2=0 $Y2=0
cc_422 N_A_742_107#_c_516_p N_A_1235_429#_c_723_n 0.0256297f $X=6.55 $Y=1.48
+ $X2=0 $Y2=0
cc_423 N_A_742_107#_c_453_n N_A_1235_429#_c_723_n 6.39904e-19 $X=6.55 $Y=1.48
+ $X2=0 $Y2=0
cc_424 N_A_742_107#_M1000_g N_A_1235_429#_c_733_n 2.93951e-19 $X=6.53 $Y=2.465
+ $X2=0 $Y2=0
cc_425 N_A_742_107#_c_458_n N_A_1235_429#_c_733_n 7.38236e-19 $X=6.55 $Y=1.985
+ $X2=0 $Y2=0
cc_426 N_A_742_107#_c_463_n N_A_1235_429#_c_733_n 0.0124196f $X=5.785 $Y=2.62
+ $X2=0 $Y2=0
cc_427 N_A_742_107#_c_464_n N_A_1235_429#_c_733_n 0.0317105f $X=5.87 $Y=2.535
+ $X2=0 $Y2=0
cc_428 N_A_742_107#_c_465_n N_A_1235_429#_c_733_n 0.0217912f $X=6.385 $Y=1.82
+ $X2=0 $Y2=0
cc_429 N_A_742_107#_c_459_n N_VPWR_M1011_d 0.00228497f $X=4.66 $Y=1.83 $X2=0
+ $Y2=0
cc_430 N_A_742_107#_c_463_n N_VPWR_M1003_d 0.00969135f $X=5.785 $Y=2.62 $X2=0
+ $Y2=0
cc_431 N_A_742_107#_c_464_n N_VPWR_M1003_d 0.0113743f $X=5.87 $Y=2.535 $X2=0
+ $Y2=0
cc_432 N_A_742_107#_M1011_g N_VPWR_c_817_n 0.0215505f $X=4.015 $Y=2.495 $X2=0
+ $Y2=0
cc_433 N_A_742_107#_c_459_n N_VPWR_c_817_n 0.031351f $X=4.66 $Y=1.83 $X2=0 $Y2=0
cc_434 N_A_742_107#_c_463_n N_VPWR_c_818_n 0.0251047f $X=5.785 $Y=2.62 $X2=0
+ $Y2=0
cc_435 N_A_742_107#_M1000_g N_VPWR_c_819_n 0.00773264f $X=6.53 $Y=2.465 $X2=0
+ $Y2=0
cc_436 N_A_742_107#_c_461_n N_VPWR_c_822_n 0.0177877f $X=4.755 $Y=2.91 $X2=0
+ $Y2=0
cc_437 N_A_742_107#_c_463_n N_VPWR_c_822_n 0.01197f $X=5.785 $Y=2.62 $X2=0 $Y2=0
cc_438 N_A_742_107#_M1011_g N_VPWR_c_825_n 0.00289833f $X=4.015 $Y=2.495 $X2=0
+ $Y2=0
cc_439 N_A_742_107#_M1000_g N_VPWR_c_826_n 0.00382362f $X=6.53 $Y=2.465 $X2=0
+ $Y2=0
cc_440 N_A_742_107#_M1019_d N_VPWR_c_813_n 0.00368844f $X=4.615 $Y=1.825 $X2=0
+ $Y2=0
cc_441 N_A_742_107#_M1011_g N_VPWR_c_813_n 0.00331732f $X=4.015 $Y=2.495 $X2=0
+ $Y2=0
cc_442 N_A_742_107#_M1000_g N_VPWR_c_813_n 0.00413371f $X=6.53 $Y=2.465 $X2=0
+ $Y2=0
cc_443 N_A_742_107#_c_461_n N_VPWR_c_813_n 0.010026f $X=4.755 $Y=2.91 $X2=0
+ $Y2=0
cc_444 N_A_742_107#_c_463_n N_VPWR_c_813_n 0.022139f $X=5.785 $Y=2.62 $X2=0
+ $Y2=0
cc_445 N_A_742_107#_M1008_g N_VGND_c_1018_n 0.00166921f $X=6.155 $Y=0.58 $X2=0
+ $Y2=0
cc_446 N_A_742_107#_M1008_g N_VGND_c_1019_n 0.00509788f $X=6.155 $Y=0.58 $X2=0
+ $Y2=0
cc_447 N_A_742_107#_M1013_g N_VGND_c_1023_n 6.65218e-19 $X=3.785 $Y=0.875 $X2=0
+ $Y2=0
cc_448 N_A_742_107#_M1008_g N_VGND_c_1025_n 0.00436358f $X=6.155 $Y=0.58 $X2=0
+ $Y2=0
cc_449 N_A_742_107#_M1016_d N_VGND_c_1031_n 0.00288526f $X=4.45 $Y=0.245 $X2=0
+ $Y2=0
cc_450 N_A_742_107#_M1008_g N_VGND_c_1031_n 0.00827976f $X=6.155 $Y=0.58 $X2=0
+ $Y2=0
cc_451 N_A_614_133#_c_592_n N_CLK_c_650_n 0.00350077f $X=4.465 $Y=1.39 $X2=0
+ $Y2=0
cc_452 N_A_614_133#_M1019_g N_VPWR_c_817_n 0.0229556f $X=4.54 $Y=2.455 $X2=0
+ $Y2=0
cc_453 N_A_614_133#_c_588_n N_VPWR_c_817_n 0.0129994f $X=3.44 $Y=2.49 $X2=0
+ $Y2=0
cc_454 N_A_614_133#_M1019_g N_VPWR_c_822_n 0.00477554f $X=4.54 $Y=2.455 $X2=0
+ $Y2=0
cc_455 N_A_614_133#_c_588_n N_VPWR_c_825_n 0.00357547f $X=3.44 $Y=2.49 $X2=0
+ $Y2=0
cc_456 N_A_614_133#_M1019_g N_VPWR_c_813_n 0.00955784f $X=4.54 $Y=2.455 $X2=0
+ $Y2=0
cc_457 N_A_614_133#_c_588_n N_VPWR_c_813_n 0.00608178f $X=3.44 $Y=2.49 $X2=0
+ $Y2=0
cc_458 N_A_614_133#_c_590_n N_A_110_70#_c_915_n 0.0311391f $X=3.21 $Y=0.95 $X2=0
+ $Y2=0
cc_459 N_A_614_133#_c_588_n N_A_110_70#_c_916_n 0.034585f $X=3.44 $Y=2.49 $X2=0
+ $Y2=0
cc_460 N_A_614_133#_M1016_g N_VGND_c_1024_n 0.00400062f $X=4.375 $Y=0.665 $X2=0
+ $Y2=0
cc_461 N_A_614_133#_M1016_g N_VGND_c_1028_n 0.00659856f $X=4.375 $Y=0.665 $X2=0
+ $Y2=0
cc_462 N_A_614_133#_M1016_g N_VGND_c_1031_n 0.00814141f $X=4.375 $Y=0.665 $X2=0
+ $Y2=0
cc_463 N_CLK_c_651_n N_A_1235_429#_c_720_n 0.0020907f $X=5.795 $Y=0.9 $X2=0
+ $Y2=0
cc_464 CLK N_A_1235_429#_c_720_n 0.00752209f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_465 N_CLK_c_650_n N_A_1235_429#_c_722_n 5.64437e-19 $X=5.51 $Y=1.855 $X2=0
+ $Y2=0
cc_466 CLK N_A_1235_429#_c_722_n 0.00664603f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_467 N_CLK_M1003_g N_A_1235_429#_c_733_n 6.94601e-19 $X=5.51 $Y=2.465 $X2=0
+ $Y2=0
cc_468 N_CLK_M1022_g N_A_1235_429#_c_733_n 0.0111327f $X=6.1 $Y=2.465 $X2=0
+ $Y2=0
cc_469 N_CLK_M1003_g N_VPWR_c_818_n 0.00116328f $X=5.51 $Y=2.465 $X2=0 $Y2=0
cc_470 N_CLK_M1022_g N_VPWR_c_818_n 6.30742e-19 $X=6.1 $Y=2.465 $X2=0 $Y2=0
cc_471 N_CLK_M1022_g N_VPWR_c_819_n 4.56228e-19 $X=6.1 $Y=2.465 $X2=0 $Y2=0
cc_472 N_CLK_M1003_g N_VPWR_c_822_n 0.00353281f $X=5.51 $Y=2.465 $X2=0 $Y2=0
cc_473 N_CLK_M1022_g N_VPWR_c_826_n 0.00441517f $X=6.1 $Y=2.465 $X2=0 $Y2=0
cc_474 N_CLK_M1003_g N_VPWR_c_813_n 0.00492109f $X=5.51 $Y=2.465 $X2=0 $Y2=0
cc_475 N_CLK_M1022_g N_VPWR_c_813_n 0.00492109f $X=6.1 $Y=2.465 $X2=0 $Y2=0
cc_476 N_CLK_c_649_n N_VGND_c_1018_n 0.0109346f $X=5.365 $Y=0.9 $X2=0 $Y2=0
cc_477 N_CLK_c_650_n N_VGND_c_1018_n 6.67588e-19 $X=5.51 $Y=1.855 $X2=0 $Y2=0
cc_478 N_CLK_c_651_n N_VGND_c_1018_n 0.00948355f $X=5.795 $Y=0.9 $X2=0 $Y2=0
cc_479 CLK N_VGND_c_1018_n 0.0238495f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_480 N_CLK_c_649_n N_VGND_c_1024_n 0.00383152f $X=5.365 $Y=0.9 $X2=0 $Y2=0
cc_481 N_CLK_c_651_n N_VGND_c_1025_n 0.00383152f $X=5.795 $Y=0.9 $X2=0 $Y2=0
cc_482 N_CLK_c_649_n N_VGND_c_1031_n 0.00762539f $X=5.365 $Y=0.9 $X2=0 $Y2=0
cc_483 N_CLK_c_651_n N_VGND_c_1031_n 0.00623447f $X=5.795 $Y=0.9 $X2=0 $Y2=0
cc_484 CLK N_VGND_c_1031_n 0.00260448f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_485 N_A_1235_429#_c_729_n N_VPWR_M1000_d 0.00479681f $X=6.895 $Y=2.23 $X2=0
+ $Y2=0
cc_486 N_A_1235_429#_c_723_n N_VPWR_M1000_d 0.00521807f $X=7.005 $Y=2.075 $X2=0
+ $Y2=0
cc_487 N_A_1235_429#_c_767_p N_VPWR_M1000_d 0.00374919f $X=7.005 $Y=2.23 $X2=0
+ $Y2=0
cc_488 N_A_1235_429#_c_731_n N_VPWR_M1009_d 0.00310159f $X=7.785 $Y=2.3 $X2=0
+ $Y2=0
cc_489 N_A_1235_429#_c_724_n N_VPWR_M1009_d 0.00315154f $X=7.88 $Y=1.46 $X2=0
+ $Y2=0
cc_490 N_A_1235_429#_M1004_g N_VPWR_c_819_n 0.0185831f $X=7.235 $Y=2.465 $X2=0
+ $Y2=0
cc_491 N_A_1235_429#_M1009_g N_VPWR_c_819_n 0.00202515f $X=7.665 $Y=2.465 $X2=0
+ $Y2=0
cc_492 N_A_1235_429#_c_729_n N_VPWR_c_819_n 0.0215811f $X=6.895 $Y=2.23 $X2=0
+ $Y2=0
cc_493 N_A_1235_429#_c_731_n N_VPWR_c_819_n 0.00182821f $X=7.785 $Y=2.3 $X2=0
+ $Y2=0
cc_494 N_A_1235_429#_c_733_n N_VPWR_c_819_n 0.0126797f $X=6.315 $Y=2.32 $X2=0
+ $Y2=0
cc_495 N_A_1235_429#_c_767_p N_VPWR_c_819_n 0.0187086f $X=7.005 $Y=2.23 $X2=0
+ $Y2=0
cc_496 N_A_1235_429#_M1004_g N_VPWR_c_821_n 0.0020169f $X=7.235 $Y=2.465 $X2=0
+ $Y2=0
cc_497 N_A_1235_429#_M1009_g N_VPWR_c_821_n 0.0181237f $X=7.665 $Y=2.465 $X2=0
+ $Y2=0
cc_498 N_A_1235_429#_c_731_n N_VPWR_c_821_n 0.0241939f $X=7.785 $Y=2.3 $X2=0
+ $Y2=0
cc_499 N_A_1235_429#_c_733_n N_VPWR_c_826_n 0.00698343f $X=6.315 $Y=2.32 $X2=0
+ $Y2=0
cc_500 N_A_1235_429#_M1004_g N_VPWR_c_827_n 0.00486043f $X=7.235 $Y=2.465 $X2=0
+ $Y2=0
cc_501 N_A_1235_429#_M1009_g N_VPWR_c_827_n 0.00486043f $X=7.665 $Y=2.465 $X2=0
+ $Y2=0
cc_502 N_A_1235_429#_M1004_g N_VPWR_c_813_n 0.00835506f $X=7.235 $Y=2.465 $X2=0
+ $Y2=0
cc_503 N_A_1235_429#_M1009_g N_VPWR_c_813_n 0.00835506f $X=7.665 $Y=2.465 $X2=0
+ $Y2=0
cc_504 N_A_1235_429#_c_733_n N_VPWR_c_813_n 0.00857557f $X=6.315 $Y=2.32 $X2=0
+ $Y2=0
cc_505 N_A_1235_429#_c_731_n N_GCLK_M1004_s 0.00809843f $X=7.785 $Y=2.3 $X2=0
+ $Y2=0
cc_506 N_A_1235_429#_M1004_g N_GCLK_c_998_n 0.00331889f $X=7.235 $Y=2.465 $X2=0
+ $Y2=0
cc_507 N_A_1235_429#_M1009_g N_GCLK_c_998_n 0.00235741f $X=7.665 $Y=2.465 $X2=0
+ $Y2=0
cc_508 N_A_1235_429#_c_731_n N_GCLK_c_998_n 0.0169068f $X=7.785 $Y=2.3 $X2=0
+ $Y2=0
cc_509 N_A_1235_429#_M1001_g N_GCLK_c_995_n 0.00241527f $X=7.235 $Y=0.695 $X2=0
+ $Y2=0
cc_510 N_A_1235_429#_M1004_g N_GCLK_c_995_n 0.00335521f $X=7.235 $Y=2.465 $X2=0
+ $Y2=0
cc_511 N_A_1235_429#_M1012_g N_GCLK_c_995_n 0.0200643f $X=7.665 $Y=0.695 $X2=0
+ $Y2=0
cc_512 N_A_1235_429#_M1009_g N_GCLK_c_995_n 0.00441153f $X=7.665 $Y=2.465 $X2=0
+ $Y2=0
cc_513 N_A_1235_429#_c_721_n N_GCLK_c_995_n 0.00697241f $X=6.895 $Y=1.13 $X2=0
+ $Y2=0
cc_514 N_A_1235_429#_c_723_n N_GCLK_c_995_n 0.0391649f $X=7.005 $Y=2.075 $X2=0
+ $Y2=0
cc_515 N_A_1235_429#_c_724_n N_GCLK_c_995_n 0.0477583f $X=7.88 $Y=1.46 $X2=0
+ $Y2=0
cc_516 N_A_1235_429#_c_725_n N_GCLK_c_995_n 0.00705365f $X=7.88 $Y=1.46 $X2=0
+ $Y2=0
cc_517 N_A_1235_429#_c_726_n N_GCLK_c_995_n 0.00983897f $X=7.59 $Y=1.46 $X2=0
+ $Y2=0
cc_518 N_A_1235_429#_c_721_n N_VGND_M1001_d 0.0031702f $X=6.895 $Y=1.13 $X2=0
+ $Y2=0
cc_519 N_A_1235_429#_c_720_n N_VGND_c_1018_n 0.00736062f $X=6.37 $Y=0.555 $X2=0
+ $Y2=0
cc_520 N_A_1235_429#_M1001_g N_VGND_c_1019_n 0.0109411f $X=7.235 $Y=0.695 $X2=0
+ $Y2=0
cc_521 N_A_1235_429#_M1012_g N_VGND_c_1019_n 6.22262e-19 $X=7.665 $Y=0.695 $X2=0
+ $Y2=0
cc_522 N_A_1235_429#_c_720_n N_VGND_c_1019_n 0.0233393f $X=6.37 $Y=0.555 $X2=0
+ $Y2=0
cc_523 N_A_1235_429#_c_721_n N_VGND_c_1019_n 0.0228247f $X=6.895 $Y=1.13 $X2=0
+ $Y2=0
cc_524 N_A_1235_429#_M1012_g N_VGND_c_1021_n 0.00629369f $X=7.665 $Y=0.695 $X2=0
+ $Y2=0
cc_525 N_A_1235_429#_c_724_n N_VGND_c_1021_n 0.0230019f $X=7.88 $Y=1.46 $X2=0
+ $Y2=0
cc_526 N_A_1235_429#_c_725_n N_VGND_c_1021_n 0.002042f $X=7.88 $Y=1.46 $X2=0
+ $Y2=0
cc_527 N_A_1235_429#_c_720_n N_VGND_c_1025_n 0.00924118f $X=6.37 $Y=0.555 $X2=0
+ $Y2=0
cc_528 N_A_1235_429#_M1001_g N_VGND_c_1026_n 0.00489337f $X=7.235 $Y=0.695 $X2=0
+ $Y2=0
cc_529 N_A_1235_429#_M1012_g N_VGND_c_1026_n 0.00511358f $X=7.665 $Y=0.695 $X2=0
+ $Y2=0
cc_530 N_A_1235_429#_M1001_g N_VGND_c_1031_n 0.00877123f $X=7.235 $Y=0.695 $X2=0
+ $Y2=0
cc_531 N_A_1235_429#_M1012_g N_VGND_c_1031_n 0.0102336f $X=7.665 $Y=0.695 $X2=0
+ $Y2=0
cc_532 N_A_1235_429#_c_720_n N_VGND_c_1031_n 0.0112261f $X=6.37 $Y=0.555 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_815_n N_A_110_70#_c_918_n 0.0250121f $X=0.26 $Y=2.495 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_816_n N_A_110_70#_c_918_n 0.0323977f $X=1.63 $Y=2.6 $X2=0 $Y2=0
cc_535 N_VPWR_c_824_n N_A_110_70#_c_918_n 0.0287361f $X=1.465 $Y=3.33 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_813_n N_A_110_70#_c_918_n 0.0226124f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_537 N_VPWR_M1007_s N_A_110_70#_c_919_n 0.00597923f $X=1.475 $Y=2.44 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_816_n N_A_110_70#_c_919_n 0.0265244f $X=1.63 $Y=2.6 $X2=0 $Y2=0
cc_539 N_VPWR_c_816_n N_A_110_70#_c_920_n 0.0292273f $X=1.63 $Y=2.6 $X2=0 $Y2=0
cc_540 N_VPWR_c_825_n N_A_110_70#_c_921_n 0.0635422f $X=4.045 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_813_n N_A_110_70#_c_921_n 0.0339568f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_542 N_VPWR_c_816_n N_A_110_70#_c_922_n 0.0150384f $X=1.63 $Y=2.6 $X2=0 $Y2=0
cc_543 N_VPWR_c_825_n N_A_110_70#_c_922_n 0.0114574f $X=4.045 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_813_n N_A_110_70#_c_922_n 0.00589978f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_815_n N_A_110_70#_c_924_n 4.20713e-19 $X=0.26 $Y=2.495 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_813_n N_GCLK_M1004_s 0.0119922f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_547 N_A_110_70#_c_992_p N_VGND_c_1022_n 0.0071868f $X=0.69 $Y=0.56 $X2=0
+ $Y2=0
cc_548 N_A_110_70#_c_992_p N_VGND_c_1031_n 0.00798886f $X=0.69 $Y=0.56 $X2=0
+ $Y2=0
cc_549 N_A_110_70#_c_914_n N_VGND_c_1031_n 2.45469e-19 $X=0.702 $Y=0.93 $X2=0
+ $Y2=0
cc_550 N_GCLK_c_995_n N_VGND_c_1019_n 0.0240307f $X=7.45 $Y=0.42 $X2=0 $Y2=0
cc_551 N_GCLK_c_995_n N_VGND_c_1021_n 0.0327798f $X=7.45 $Y=0.42 $X2=0 $Y2=0
cc_552 N_GCLK_c_995_n N_VGND_c_1026_n 0.0191277f $X=7.45 $Y=0.42 $X2=0 $Y2=0
cc_553 N_GCLK_c_995_n N_VGND_c_1031_n 0.0103094f $X=7.45 $Y=0.42 $X2=0 $Y2=0
