* File: sky130_fd_sc_lp__nor2_0.pex.spice
* Created: Wed Sep  2 10:07:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2_0%A 2 5 8 10 11 12 13 14 20 22
c25 11 0 2.72248e-20 $X=0.24 $Y=0.925
r26 20 22 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.045
+ $X2=0.402 $Y2=0.88
r27 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.37
+ $Y=1.045 $X2=0.37 $Y2=1.045
r28 13 14 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=2.035
r29 12 13 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.665
r30 12 21 7.78678 $w=3.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.045
r31 11 21 3.73765 $w=3.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.27 $Y=0.925
+ $X2=0.27 $Y2=1.045
r32 8 10 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.525 $Y=2.735
+ $X2=0.525 $Y2=1.55
r33 5 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.525 $Y=0.56
+ $X2=0.525 $Y2=0.88
r34 2 10 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.402 $Y=1.353
+ $X2=0.402 $Y2=1.55
r35 1 20 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.402 $Y=1.077
+ $X2=0.402 $Y2=1.045
r36 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.402 $Y=1.077
+ $X2=0.402 $Y2=1.353
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_0%B 3 7 8 9 10 11 17 19
c27 19 0 2.72248e-20 $X=1.087 $Y=0.88
r28 17 20 83.1449 $w=4.95e-07 $l=5.05e-07 $layer=POLY_cond $X=1.087 $Y=1.045
+ $X2=1.087 $Y2=1.55
r29 17 19 46.3954 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.087 $Y=1.045
+ $X2=1.087 $Y2=0.88
r30 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.045 $X2=1.17 $Y2=1.045
r31 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=1.665
+ $X2=1.205 $Y2=2.035
r32 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=1.295
+ $X2=1.205 $Y2=1.665
r33 9 18 9.60369 $w=2.98e-07 $l=2.5e-07 $layer=LI1_cond $X=1.205 $Y=1.295
+ $X2=1.205 $Y2=1.045
r34 8 18 4.60977 $w=2.98e-07 $l=1.2e-07 $layer=LI1_cond $X=1.205 $Y=0.925
+ $X2=1.205 $Y2=1.045
r35 7 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.955 $Y=0.56
+ $X2=0.955 $Y2=0.88
r36 3 20 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.915 $Y=2.735
+ $X2=0.915 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_0%VPWR 1 4 6 8 12 13
r15 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r16 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r17 10 16 4.48864 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r18 10 12 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=1.2 $Y2=3.33
r19 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33 $X2=1.2
+ $Y2=3.33
r20 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r21 4 16 3.11055 $w=3.1e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.227 $Y2=3.33
r22 4 6 25.4653 $w=3.08e-07 $l=6.85e-07 $layer=LI1_cond $X=0.3 $Y=3.245 $X2=0.3
+ $Y2=2.56
r23 1 6 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=2.415 $X2=0.31 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_0%Y 1 2 7 8 9 10 11 12 22 34
c17 34 0 1.06273e-19 $X=0.72 $Y=2.405
r18 34 35 4.83316 $w=6.68e-07 $l=1e-08 $layer=LI1_cond $X=0.96 $Y=2.405 $X2=0.96
+ $Y2=2.395
r19 12 38 3.83816 $w=6.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.96 $Y=2.775
+ $X2=0.96 $Y2=2.56
r20 11 38 2.10653 $w=6.68e-07 $l=1.18e-07 $layer=LI1_cond $X=0.96 $Y=2.442
+ $X2=0.96 $Y2=2.56
r21 11 34 0.660521 $w=6.68e-07 $l=3.7e-08 $layer=LI1_cond $X=0.96 $Y=2.442
+ $X2=0.96 $Y2=2.405
r22 11 35 1.68434 $w=2.58e-07 $l=3.8e-08 $layer=LI1_cond $X=0.755 $Y=2.357
+ $X2=0.755 $Y2=2.395
r23 10 11 14.2726 $w=2.58e-07 $l=3.22e-07 $layer=LI1_cond $X=0.755 $Y=2.035
+ $X2=0.755 $Y2=2.357
r24 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.755 $Y=1.665
+ $X2=0.755 $Y2=2.035
r25 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.755 $Y=1.295
+ $X2=0.755 $Y2=1.665
r26 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.755 $Y=0.925
+ $X2=0.755 $Y2=1.295
r27 7 22 16.6218 $w=2.58e-07 $l=3.75e-07 $layer=LI1_cond $X=0.755 $Y=0.925
+ $X2=0.755 $Y2=0.55
r28 2 38 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.99
+ $Y=2.415 $X2=1.13 $Y2=2.56
r29 1 22 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.35 $X2=0.74 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_0%VGND 1 2 7 9 11 13 15 17 27
r22 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r23 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r24 18 23 4.48864 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r25 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r26 17 26 4.29523 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.247
+ $Y2=0
r27 17 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.72
+ $Y2=0
r28 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r29 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r30 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r31 11 26 3.06482 $w=2.8e-07 $l=1.07912e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.247 $Y2=0
r32 11 13 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0.505
r33 7 23 3.11055 $w=3.1e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.227 $Y2=0
r34 7 9 15.6137 $w=3.08e-07 $l=4.2e-07 $layer=LI1_cond $X=0.3 $Y=0.085 $X2=0.3
+ $Y2=0.505
r35 2 13 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.35 $X2=1.17 $Y2=0.505
r36 1 9 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.35 $X2=0.31 $Y2=0.505
.ends

