* NGSPICE file created from sky130_fd_sc_lp__and3_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and3_2 A B C VGND VNB VPB VPWR X
M1000 VPWR A a_27_385# VPB phighvt w=420000u l=150000u
+  ad=8.505e+11p pd=7.75e+06u as=2.604e+11p ps=2.92e+06u
M1001 X a_27_385# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1002 X a_27_385# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=5.649e+11p ps=4.96e+06u
M1003 a_27_385# B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_196_47# B a_124_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1005 VGND C a_196_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C a_27_385# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_27_385# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_124_47# A a_27_385# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 VGND a_27_385# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

