* File: sky130_fd_sc_lp__nand4b_1.spice
* Created: Wed Sep  2 10:06:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4b_1.pex.spice"
.subckt sky130_fd_sc_lp__nand4b_1  VNB VPB A_N D C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* D	D
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_N_M1003_g N_A_71_131#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0938 AS=0.1113 PD=0.82 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 A_262_47# N_D_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.1876 PD=1.05 PS=1.64 NRD=7.14 NRS=5.352 M=1 R=5.6 SA=75000.5 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1005 A_334_47# N_C_M1005_g A_262_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75000.8 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1007 A_442_47# N_B_M1007_g A_334_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.1638 PD=1.23 PS=1.23 NRD=19.992 NRS=19.992 M=1 R=5.6 SA=75001.4
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_A_71_131#_M1000_g A_442_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_A_N_M1006_g N_A_71_131#_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0966 AS=0.1113 PD=0.825 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_D_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2898 PD=1.54 PS=2.475 NRD=0 NRS=5.7327 M=1 R=8.4 SA=75000.4
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_C_M1008_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2709 AS=0.1764 PD=1.69 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2709 PD=1.54 PS=1.69 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75001.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_71_131#_M1009_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_53 VPB 0 2.00567e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__nand4b_1.pxi.spice"
*
.ends
*
*
