* File: sky130_fd_sc_lp__mux4_2.pxi.spice
* Created: Fri Aug 28 10:46:12 2020
* 
x_PM_SKY130_FD_SC_LP__MUX4_2%A_80_293# N_A_80_293#_M1023_s N_A_80_293#_M1025_s
+ N_A_80_293#_M1005_g N_A_80_293#_c_163_n N_A_80_293#_c_164_n
+ N_A_80_293#_c_165_n N_A_80_293#_M1003_g N_A_80_293#_c_166_n
+ N_A_80_293#_c_167_n N_A_80_293#_c_171_n N_A_80_293#_c_168_n
+ N_A_80_293#_c_169_n PM_SKY130_FD_SC_LP__MUX4_2%A_80_293#
x_PM_SKY130_FD_SC_LP__MUX4_2%S1 N_S1_M1013_g N_S1_c_224_n N_S1_c_225_n
+ N_S1_c_229_n N_S1_M1017_g N_S1_c_230_n N_S1_c_231_n N_S1_M1025_g N_S1_M1023_g
+ S1 S1 N_S1_c_227_n N_S1_c_228_n PM_SKY130_FD_SC_LP__MUX4_2%S1
x_PM_SKY130_FD_SC_LP__MUX4_2%A_110_125# N_A_110_125#_M1013_d
+ N_A_110_125#_M1005_d N_A_110_125#_M1002_g N_A_110_125#_c_302_n
+ N_A_110_125#_M1015_g N_A_110_125#_M1019_g N_A_110_125#_c_304_n
+ N_A_110_125#_M1024_g N_A_110_125#_c_305_n N_A_110_125#_c_306_n
+ N_A_110_125#_c_307_n N_A_110_125#_c_308_n N_A_110_125#_c_309_n
+ N_A_110_125#_c_310_n N_A_110_125#_c_311_n
+ PM_SKY130_FD_SC_LP__MUX4_2%A_110_125#
x_PM_SKY130_FD_SC_LP__MUX4_2%A3 N_A3_M1021_g N_A3_M1018_g A3 A3 A3 N_A3_c_396_n
+ PM_SKY130_FD_SC_LP__MUX4_2%A3
x_PM_SKY130_FD_SC_LP__MUX4_2%A_859_351# N_A_859_351#_M1006_d
+ N_A_859_351#_M1008_d N_A_859_351#_M1026_g N_A_859_351#_c_433_n
+ N_A_859_351#_c_434_n N_A_859_351#_M1011_g N_A_859_351#_M1027_g
+ N_A_859_351#_c_437_n N_A_859_351#_c_438_n N_A_859_351#_M1001_g
+ N_A_859_351#_c_440_n N_A_859_351#_c_457_n N_A_859_351#_c_441_n
+ N_A_859_351#_c_442_n N_A_859_351#_c_443_n N_A_859_351#_c_444_n
+ N_A_859_351#_c_445_n N_A_859_351#_c_584_p N_A_859_351#_c_446_n
+ N_A_859_351#_c_447_n N_A_859_351#_c_448_n N_A_859_351#_c_449_n
+ N_A_859_351#_c_450_n N_A_859_351#_c_451_n N_A_859_351#_c_452_n
+ N_A_859_351#_c_458_n N_A_859_351#_c_453_n
+ PM_SKY130_FD_SC_LP__MUX4_2%A_859_351#
x_PM_SKY130_FD_SC_LP__MUX4_2%A2 N_A2_c_593_n N_A2_M1010_g N_A2_M1020_g A2 A2
+ PM_SKY130_FD_SC_LP__MUX4_2%A2
x_PM_SKY130_FD_SC_LP__MUX4_2%A1 N_A1_M1007_g N_A1_M1022_g N_A1_c_640_n
+ N_A1_c_645_n A1 A1 N_A1_c_641_n N_A1_c_642_n PM_SKY130_FD_SC_LP__MUX4_2%A1
x_PM_SKY130_FD_SC_LP__MUX4_2%A0 N_A0_M1004_g N_A0_M1016_g A0 A0 N_A0_c_686_n
+ PM_SKY130_FD_SC_LP__MUX4_2%A0
x_PM_SKY130_FD_SC_LP__MUX4_2%S0 N_S0_M1009_g N_S0_c_721_n N_S0_c_722_n
+ N_S0_M1012_g N_S0_c_730_n N_S0_c_731_n N_S0_M1000_g N_S0_c_724_n N_S0_M1014_g
+ N_S0_c_733_n N_S0_M1006_g N_S0_M1008_g N_S0_c_726_n N_S0_c_735_n N_S0_c_727_n
+ N_S0_c_736_n S0 N_S0_c_728_n N_S0_c_769_n PM_SKY130_FD_SC_LP__MUX4_2%S0
x_PM_SKY130_FD_SC_LP__MUX4_2%A_27_125# N_A_27_125#_M1013_s N_A_27_125#_M1009_d
+ N_A_27_125#_M1005_s N_A_27_125#_M1026_d N_A_27_125#_c_833_n
+ N_A_27_125#_c_837_n N_A_27_125#_c_838_n N_A_27_125#_c_839_n
+ N_A_27_125#_c_840_n N_A_27_125#_c_841_n N_A_27_125#_c_834_n
+ N_A_27_125#_c_835_n N_A_27_125#_c_843_n PM_SKY130_FD_SC_LP__MUX4_2%A_27_125#
x_PM_SKY130_FD_SC_LP__MUX4_2%A_196_125# N_A_196_125#_M1003_d
+ N_A_196_125#_M1000_d N_A_196_125#_M1017_d N_A_196_125#_M1027_d
+ N_A_196_125#_c_931_n N_A_196_125#_c_934_n N_A_196_125#_c_932_n
+ N_A_196_125#_c_975_n N_A_196_125#_c_936_n N_A_196_125#_c_937_n
+ N_A_196_125#_c_938_n N_A_196_125#_c_982_n N_A_196_125#_c_939_n
+ N_A_196_125#_c_933_n PM_SKY130_FD_SC_LP__MUX4_2%A_196_125#
x_PM_SKY130_FD_SC_LP__MUX4_2%VPWR N_VPWR_M1025_d N_VPWR_M1019_s N_VPWR_M1010_d
+ N_VPWR_M1016_d N_VPWR_c_1037_n N_VPWR_c_1038_n N_VPWR_c_1039_n N_VPWR_c_1040_n
+ N_VPWR_c_1041_n N_VPWR_c_1042_n N_VPWR_c_1043_n VPWR N_VPWR_c_1044_n
+ N_VPWR_c_1045_n N_VPWR_c_1046_n N_VPWR_c_1047_n N_VPWR_c_1036_n
+ N_VPWR_c_1049_n N_VPWR_c_1050_n N_VPWR_c_1051_n
+ PM_SKY130_FD_SC_LP__MUX4_2%VPWR
x_PM_SKY130_FD_SC_LP__MUX4_2%X N_X_M1015_d N_X_M1002_d X X X X X N_X_c_1133_n
+ PM_SKY130_FD_SC_LP__MUX4_2%X
x_PM_SKY130_FD_SC_LP__MUX4_2%VGND N_VGND_M1023_d N_VGND_M1024_s N_VGND_M1020_d
+ N_VGND_M1004_d N_VGND_c_1155_n N_VGND_c_1156_n N_VGND_c_1157_n VGND
+ N_VGND_c_1158_n N_VGND_c_1159_n N_VGND_c_1160_n N_VGND_c_1161_n
+ N_VGND_c_1162_n N_VGND_c_1163_n N_VGND_c_1164_n N_VGND_c_1165_n
+ N_VGND_c_1166_n N_VGND_c_1167_n PM_SKY130_FD_SC_LP__MUX4_2%VGND
cc_1 VNB N_A_80_293#_M1005_g 0.00254372f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.305
cc_2 VNB N_A_80_293#_c_163_n 0.019954f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.54
cc_3 VNB N_A_80_293#_c_164_n 0.00918052f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.54
cc_4 VNB N_A_80_293#_c_165_n 0.017743f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.155
cc_5 VNB N_A_80_293#_c_166_n 0.0161274f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.115
cc_6 VNB N_A_80_293#_c_167_n 0.00859308f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.32
cc_7 VNB N_A_80_293#_c_168_n 8.06243e-19 $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.825
cc_8 VNB N_A_80_293#_c_169_n 0.0770737f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.49
cc_9 VNB N_S1_M1013_g 0.0428709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_S1_c_224_n 0.127752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_S1_c_225_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_S1_M1023_g 0.0358021f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.32
cc_13 VNB N_S1_c_227_n 0.00229553f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.49
cc_14 VNB N_S1_c_228_n 0.0351338f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.49
cc_15 VNB N_A_110_125#_M1002_g 0.00425265f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=2.305
cc_16 VNB N_A_110_125#_c_302_n 0.0178561f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.54
cc_17 VNB N_A_110_125#_M1019_g 0.00436585f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=1.115
cc_18 VNB N_A_110_125#_c_304_n 0.0187617f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.32
cc_19 VNB N_A_110_125#_c_305_n 0.0117803f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.17
cc_20 VNB N_A_110_125#_c_306_n 0.0157679f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.825
cc_21 VNB N_A_110_125#_c_307_n 0.00458975f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.49
cc_22 VNB N_A_110_125#_c_308_n 0.0108873f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.49
cc_23 VNB N_A_110_125#_c_309_n 0.0108293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_110_125#_c_310_n 0.0114866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_110_125#_c_311_n 0.0632412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A3_M1021_g 0.00669677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A3_M1018_g 0.0213207f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.615
cc_28 VNB A3 0.0120895f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.305
cc_29 VNB N_A3_c_396_n 0.0329453f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.17
cc_30 VNB N_A_859_351#_c_433_n 0.0153313f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.155
cc_31 VNB N_A_859_351#_c_434_n 0.00677107f $X=-0.19 $Y=-0.245 $X2=0.905
+ $Y2=0.835
cc_32 VNB N_A_859_351#_M1011_g 0.015441f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.525
cc_33 VNB N_A_859_351#_M1027_g 0.00723117f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.825
cc_34 VNB N_A_859_351#_c_437_n 0.0154231f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.17
cc_35 VNB N_A_859_351#_c_438_n 0.00673671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_859_351#_M1001_g 0.0155442f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.825
cc_37 VNB N_A_859_351#_c_440_n 0.00741911f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.49
cc_38 VNB N_A_859_351#_c_441_n 0.0143752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_859_351#_c_442_n 0.00178286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_859_351#_c_443_n 0.018688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_859_351#_c_444_n 0.00249631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_859_351#_c_445_n 0.00558082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_859_351#_c_446_n 0.0258772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_859_351#_c_447_n 0.00112393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_859_351#_c_448_n 0.0394835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_859_351#_c_449_n 0.00468383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_859_351#_c_450_n 0.00357846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_859_351#_c_451_n 0.038011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_859_351#_c_452_n 0.00211907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_859_351#_c_453_n 0.0240857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A2_c_593_n 0.0229775f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=0.655
cc_52 VNB N_A2_M1020_g 0.0313379f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.615
cc_53 VNB A2 0.00916735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A1_M1007_g 0.0231167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A1_c_640_n 0.0148947f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.54
cc_56 VNB N_A1_c_641_n 0.0177789f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.32
cc_57 VNB N_A1_c_642_n 0.00267987f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.32
cc_58 VNB N_A0_M1004_g 0.0403475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB A0 0.00953123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A0_c_686_n 0.00888828f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.835
cc_61 VNB N_S0_M1009_g 0.0325318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_S0_c_721_n 0.140507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_S0_c_722_n 0.0125433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_S0_M1000_g 0.0295718f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.835
cc_65 VNB N_S0_c_724_n 0.0930353f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.525
cc_66 VNB N_S0_M1006_g 0.0407678f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.49
cc_67 VNB N_S0_c_726_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_S0_c_727_n 0.0294724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_S0_c_728_n 0.0238526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_27_125#_c_833_n 0.0474944f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.835
cc_71 VNB N_A_27_125#_c_834_n 0.00580522f $X=-0.19 $Y=-0.245 $X2=1.99 $Y2=0.96
cc_72 VNB N_A_27_125#_c_835_n 0.00255394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_196_125#_c_931_n 0.00801867f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.32
cc_74 VNB N_A_196_125#_c_932_n 0.00165487f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=0.96
cc_75 VNB N_A_196_125#_c_933_n 0.00641672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VPWR_c_1036_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_X_c_1133_n 0.00265194f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.32
cc_78 VNB N_VGND_c_1155_n 0.0085932f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.835
cc_79 VNB N_VGND_c_1156_n 0.0138741f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.825
cc_80 VNB N_VGND_c_1157_n 0.0028967f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=0.96
cc_81 VNB N_VGND_c_1158_n 0.0665019f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.49
cc_82 VNB N_VGND_c_1159_n 0.0159664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1160_n 0.0433962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1161_n 0.0361371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1162_n 0.0305084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1163_n 0.444971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1164_n 0.011782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1165_n 0.0101353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1166_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1167_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VPB N_A_80_293#_M1005_g 0.0311578f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.305
cc_92 VPB N_A_80_293#_c_171_n 0.00496829f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.17
cc_93 VPB N_A_80_293#_c_168_n 0.00667952f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.825
cc_94 VPB N_A_80_293#_c_169_n 0.024881f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.49
cc_95 VPB N_S1_c_229_n 0.0176643f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.615
cc_96 VPB N_S1_c_230_n 0.0757269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_S1_c_231_n 0.0109492f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=1.54
cc_98 VPB N_S1_M1025_g 0.0324976f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.835
cc_99 VPB N_S1_c_227_n 0.00217245f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.49
cc_100 VPB N_S1_c_228_n 0.0117883f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=1.49
cc_101 VPB N_A_110_125#_M1002_g 0.0240905f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.305
cc_102 VPB N_A_110_125#_M1019_g 0.0232617f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.115
cc_103 VPB N_A_110_125#_c_305_n 0.00781737f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.17
cc_104 VPB N_A3_M1021_g 0.0329915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB A3 0.00636292f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.305
cc_106 VPB N_A_859_351#_M1026_g 0.0202868f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.305
cc_107 VPB N_A_859_351#_M1027_g 0.0347447f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.825
cc_108 VPB N_A_859_351#_c_440_n 0.0061722f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=1.49
cc_109 VPB N_A_859_351#_c_457_n 0.0122637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_859_351#_c_458_n 0.0471449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_859_351#_c_453_n 0.020405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A2_c_593_n 0.0343664f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=0.655
cc_113 VPB N_A2_M1010_g 0.0211243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB A2 0.009932f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A1_M1022_g 0.0189144f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.615
cc_116 VPB N_A1_c_640_n 0.00708926f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=1.54
cc_117 VPB N_A1_c_645_n 0.0154894f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.54
cc_118 VPB N_A1_c_642_n 0.00490289f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=1.32
cc_119 VPB N_A0_M1016_g 0.0187727f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.615
cc_120 VPB A0 0.0177149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A0_c_686_n 0.0318622f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.835
cc_122 VPB N_S0_M1012_g 0.0352332f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.305
cc_123 VPB N_S0_c_730_n 0.141029f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=1.54
cc_124 VPB N_S0_c_731_n 0.012806f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.54
cc_125 VPB N_S0_M1014_g 0.0384145f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.825
cc_126 VPB N_S0_c_733_n 0.0706895f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.17
cc_127 VPB N_S0_M1008_g 0.0388657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_S0_c_735_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_S0_c_736_n 0.0187076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_S0_c_728_n 0.00800036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_27_125#_c_833_n 0.0528133f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.835
cc_132 VPB N_A_27_125#_c_837_n 0.0221189f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=1.32
cc_133 VPB N_A_27_125#_c_838_n 0.0111967f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=1.32
cc_134 VPB N_A_27_125#_c_839_n 0.00304642f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.17
cc_135 VPB N_A_27_125#_c_840_n 0.0178588f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.17
cc_136 VPB N_A_27_125#_c_841_n 0.00312531f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_27_125#_c_834_n 0.00396293f $X=-0.19 $Y=1.655 $X2=1.99 $Y2=0.96
cc_138 VPB N_A_27_125#_c_843_n 0.00642762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_196_125#_c_934_n 0.00239379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_196_125#_c_932_n 0.00456108f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=0.96
cc_141 VPB N_A_196_125#_c_936_n 0.00352366f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_196_125#_c_937_n 0.00202421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_196_125#_c_938_n 0.00493586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_196_125#_c_939_n 0.00750699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_196_125#_c_933_n 0.00687515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_1037_n 0.0130661f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.835
cc_147 VPB N_VPWR_c_1038_n 0.0133947f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=1.32
cc_148 VPB N_VPWR_c_1039_n 0.0020646f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.825
cc_149 VPB N_VPWR_c_1040_n 0.0139755f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.17
cc_150 VPB N_VPWR_c_1041_n 0.0112794f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=0.96
cc_151 VPB N_VPWR_c_1042_n 0.0429929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_1043_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_1044_n 0.0670509f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_1045_n 0.013538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_1046_n 0.0422265f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_1047_n 0.024975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_1036_n 0.0948006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_1049_n 0.00556078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_1050_n 0.00556078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_1051_n 0.0103613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_X_c_1133_n 0.00334993f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.32
cc_162 N_A_80_293#_c_164_n N_S1_M1013_g 0.00935869f $X=0.55 $Y=1.54 $X2=0 $Y2=0
cc_163 N_A_80_293#_c_165_n N_S1_M1013_g 0.01019f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_164 N_A_80_293#_c_165_n N_S1_c_224_n 0.00737308f $X=0.905 $Y=1.155 $X2=0
+ $Y2=0
cc_165 N_A_80_293#_M1005_g N_S1_c_229_n 0.0104914f $X=0.475 $Y=2.305 $X2=0 $Y2=0
cc_166 N_A_80_293#_c_171_n N_S1_c_229_n 0.0011645f $X=1.73 $Y=2.17 $X2=0 $Y2=0
cc_167 N_A_80_293#_c_169_n N_S1_c_229_n 0.0106605f $X=0.905 $Y=1.49 $X2=0 $Y2=0
cc_168 N_A_80_293#_c_171_n N_S1_c_230_n 7.17636e-19 $X=1.73 $Y=2.17 $X2=0 $Y2=0
cc_169 N_A_80_293#_c_168_n N_S1_M1025_g 0.00898787f $X=1.595 $Y=1.825 $X2=0
+ $Y2=0
cc_170 N_A_80_293#_c_166_n N_S1_M1023_g 0.00653541f $X=1.595 $Y=1.115 $X2=0
+ $Y2=0
cc_171 N_A_80_293#_c_167_n N_S1_M1023_g 0.00227557f $X=1.39 $Y=1.32 $X2=0 $Y2=0
cc_172 N_A_80_293#_c_169_n N_S1_M1023_g 4.02364e-19 $X=0.905 $Y=1.49 $X2=0 $Y2=0
cc_173 N_A_80_293#_c_166_n N_S1_c_227_n 0.0073526f $X=1.595 $Y=1.115 $X2=0 $Y2=0
cc_174 N_A_80_293#_c_167_n N_S1_c_227_n 0.0664216f $X=1.39 $Y=1.32 $X2=0 $Y2=0
cc_175 N_A_80_293#_c_169_n N_S1_c_227_n 3.77347e-19 $X=0.905 $Y=1.49 $X2=0 $Y2=0
cc_176 N_A_80_293#_c_166_n N_S1_c_228_n 0.00500502f $X=1.595 $Y=1.115 $X2=0
+ $Y2=0
cc_177 N_A_80_293#_c_167_n N_S1_c_228_n 0.00898787f $X=1.39 $Y=1.32 $X2=0 $Y2=0
cc_178 N_A_80_293#_c_169_n N_S1_c_228_n 0.0131883f $X=0.905 $Y=1.49 $X2=0 $Y2=0
cc_179 N_A_80_293#_M1005_g N_A_110_125#_c_305_n 0.00448692f $X=0.475 $Y=2.305
+ $X2=0 $Y2=0
cc_180 N_A_80_293#_c_163_n N_A_110_125#_c_305_n 0.0151693f $X=0.83 $Y=1.54 $X2=0
+ $Y2=0
cc_181 N_A_80_293#_c_165_n N_A_110_125#_c_305_n 0.0131692f $X=0.905 $Y=1.155
+ $X2=0 $Y2=0
cc_182 N_A_80_293#_c_165_n N_A_110_125#_c_306_n 0.00357386f $X=0.905 $Y=1.155
+ $X2=0 $Y2=0
cc_183 N_A_80_293#_c_166_n N_A_110_125#_c_306_n 0.00618156f $X=1.595 $Y=1.115
+ $X2=0 $Y2=0
cc_184 N_A_80_293#_c_169_n N_A_110_125#_c_306_n 0.00116654f $X=0.905 $Y=1.49
+ $X2=0 $Y2=0
cc_185 N_A_80_293#_M1023_s N_A_110_125#_c_308_n 0.00415272f $X=1.845 $Y=0.655
+ $X2=0 $Y2=0
cc_186 N_A_80_293#_c_166_n N_A_110_125#_c_308_n 0.0373798f $X=1.595 $Y=1.115
+ $X2=0 $Y2=0
cc_187 N_A_80_293#_c_166_n N_A_110_125#_c_309_n 0.00997749f $X=1.595 $Y=1.115
+ $X2=0 $Y2=0
cc_188 N_A_80_293#_c_165_n N_A_110_125#_c_310_n 0.00370797f $X=0.905 $Y=1.155
+ $X2=0 $Y2=0
cc_189 N_A_80_293#_c_166_n N_A_110_125#_c_310_n 0.00875278f $X=1.595 $Y=1.115
+ $X2=0 $Y2=0
cc_190 N_A_80_293#_c_169_n N_A_110_125#_c_310_n 4.91122e-19 $X=0.905 $Y=1.49
+ $X2=0 $Y2=0
cc_191 N_A_80_293#_c_164_n N_A_27_125#_c_833_n 0.0188802f $X=0.55 $Y=1.54 $X2=0
+ $Y2=0
cc_192 N_A_80_293#_M1005_g N_A_27_125#_c_837_n 0.00701919f $X=0.475 $Y=2.305
+ $X2=0 $Y2=0
cc_193 N_A_80_293#_c_171_n N_A_27_125#_c_840_n 0.0182542f $X=1.73 $Y=2.17 $X2=0
+ $Y2=0
cc_194 N_A_80_293#_c_171_n N_A_27_125#_c_841_n 0.00505094f $X=1.73 $Y=2.17 $X2=0
+ $Y2=0
cc_195 N_A_80_293#_c_168_n N_A_27_125#_c_841_n 0.00167165f $X=1.595 $Y=1.825
+ $X2=0 $Y2=0
cc_196 N_A_80_293#_c_169_n N_A_27_125#_c_841_n 3.54966e-19 $X=0.905 $Y=1.49
+ $X2=0 $Y2=0
cc_197 N_A_80_293#_c_165_n N_A_196_125#_c_931_n 0.00261979f $X=0.905 $Y=1.155
+ $X2=0 $Y2=0
cc_198 N_A_80_293#_c_166_n N_A_196_125#_c_931_n 0.0012825f $X=1.595 $Y=1.115
+ $X2=0 $Y2=0
cc_199 N_A_80_293#_c_169_n N_A_196_125#_c_931_n 0.00674091f $X=0.905 $Y=1.49
+ $X2=0 $Y2=0
cc_200 N_A_80_293#_c_171_n N_A_196_125#_c_934_n 0.0163065f $X=1.73 $Y=2.17 $X2=0
+ $Y2=0
cc_201 N_A_80_293#_c_169_n N_A_196_125#_c_934_n 0.00359017f $X=0.905 $Y=1.49
+ $X2=0 $Y2=0
cc_202 N_A_80_293#_c_165_n N_A_196_125#_c_932_n 0.00583143f $X=0.905 $Y=1.155
+ $X2=0 $Y2=0
cc_203 N_A_80_293#_c_166_n N_A_196_125#_c_932_n 0.00973294f $X=1.595 $Y=1.115
+ $X2=0 $Y2=0
cc_204 N_A_80_293#_c_167_n N_A_196_125#_c_932_n 0.054279f $X=1.39 $Y=1.32 $X2=0
+ $Y2=0
cc_205 N_A_80_293#_c_171_n N_A_196_125#_c_932_n 0.00693188f $X=1.73 $Y=2.17
+ $X2=0 $Y2=0
cc_206 N_A_80_293#_c_169_n N_A_196_125#_c_932_n 0.0275407f $X=0.905 $Y=1.49
+ $X2=0 $Y2=0
cc_207 N_A_80_293#_M1025_s N_A_196_125#_c_936_n 0.00480242f $X=1.605 $Y=2.025
+ $X2=0 $Y2=0
cc_208 N_A_80_293#_c_171_n N_A_196_125#_c_936_n 0.00963864f $X=1.73 $Y=2.17
+ $X2=0 $Y2=0
cc_209 N_A_80_293#_c_168_n N_A_196_125#_c_936_n 0.00624462f $X=1.595 $Y=1.825
+ $X2=0 $Y2=0
cc_210 N_A_80_293#_c_168_n N_A_196_125#_c_937_n 0.0018309f $X=1.595 $Y=1.825
+ $X2=0 $Y2=0
cc_211 N_S1_M1025_g N_A_110_125#_M1002_g 0.0162065f $X=2.04 $Y=2.095 $X2=0 $Y2=0
cc_212 N_S1_c_227_n N_A_110_125#_M1002_g 0.00887191f $X=2.16 $Y=1.45 $X2=0 $Y2=0
cc_213 N_S1_c_224_n N_A_110_125#_c_302_n 0.0213243f $X=2.245 $Y=0.18 $X2=0 $Y2=0
cc_214 N_S1_M1013_g N_A_110_125#_c_305_n 0.00460087f $X=0.475 $Y=0.835 $X2=0
+ $Y2=0
cc_215 N_S1_c_229_n N_A_110_125#_c_305_n 0.00117772f $X=0.905 $Y=2.735 $X2=0
+ $Y2=0
cc_216 N_S1_c_224_n N_A_110_125#_c_306_n 0.0132416f $X=2.245 $Y=0.18 $X2=0 $Y2=0
cc_217 N_S1_M1013_g N_A_110_125#_c_307_n 0.00837236f $X=0.475 $Y=0.835 $X2=0
+ $Y2=0
cc_218 N_S1_c_224_n N_A_110_125#_c_307_n 0.00323716f $X=2.245 $Y=0.18 $X2=0
+ $Y2=0
cc_219 N_S1_c_224_n N_A_110_125#_c_308_n 0.0100927f $X=2.245 $Y=0.18 $X2=0 $Y2=0
cc_220 N_S1_M1023_g N_A_110_125#_c_308_n 0.0171986f $X=2.32 $Y=0.865 $X2=0 $Y2=0
cc_221 N_S1_c_227_n N_A_110_125#_c_308_n 0.00397292f $X=2.16 $Y=1.45 $X2=0 $Y2=0
cc_222 N_S1_c_228_n N_A_110_125#_c_308_n 3.70877e-19 $X=2.32 $Y=1.45 $X2=0 $Y2=0
cc_223 N_S1_M1023_g N_A_110_125#_c_309_n 0.00969043f $X=2.32 $Y=0.865 $X2=0
+ $Y2=0
cc_224 N_S1_c_227_n N_A_110_125#_c_309_n 0.0111347f $X=2.16 $Y=1.45 $X2=0 $Y2=0
cc_225 N_S1_c_224_n N_A_110_125#_c_310_n 0.00390735f $X=2.245 $Y=0.18 $X2=0
+ $Y2=0
cc_226 N_S1_M1023_g N_A_110_125#_c_310_n 0.00425273f $X=2.32 $Y=0.865 $X2=0
+ $Y2=0
cc_227 N_S1_M1023_g N_A_110_125#_c_311_n 0.0228845f $X=2.32 $Y=0.865 $X2=0 $Y2=0
cc_228 N_S1_c_227_n N_A_110_125#_c_311_n 0.0013337f $X=2.16 $Y=1.45 $X2=0 $Y2=0
cc_229 N_S1_c_228_n N_A_110_125#_c_311_n 0.00262851f $X=2.32 $Y=1.45 $X2=0 $Y2=0
cc_230 N_S1_M1013_g N_A_27_125#_c_833_n 0.0033445f $X=0.475 $Y=0.835 $X2=0 $Y2=0
cc_231 N_S1_c_229_n N_A_27_125#_c_833_n 0.00220794f $X=0.905 $Y=2.735 $X2=0
+ $Y2=0
cc_232 N_S1_c_230_n N_A_27_125#_c_837_n 0.0243525f $X=1.965 $Y=2.81 $X2=0 $Y2=0
cc_233 N_S1_c_231_n N_A_27_125#_c_837_n 0.0111087f $X=0.98 $Y=2.81 $X2=0 $Y2=0
cc_234 N_S1_c_229_n N_A_27_125#_c_839_n 0.00292991f $X=0.905 $Y=2.735 $X2=0
+ $Y2=0
cc_235 N_S1_c_230_n N_A_27_125#_c_839_n 0.011291f $X=1.965 $Y=2.81 $X2=0 $Y2=0
cc_236 N_S1_M1025_g N_A_27_125#_c_839_n 0.00372426f $X=2.04 $Y=2.095 $X2=0 $Y2=0
cc_237 N_S1_c_230_n N_A_27_125#_c_840_n 0.00600387f $X=1.965 $Y=2.81 $X2=0 $Y2=0
cc_238 N_S1_M1025_g N_A_27_125#_c_840_n 0.0160019f $X=2.04 $Y=2.095 $X2=0 $Y2=0
cc_239 N_S1_c_227_n N_A_27_125#_c_840_n 0.00824163f $X=2.16 $Y=1.45 $X2=0 $Y2=0
cc_240 N_S1_c_229_n N_A_196_125#_c_934_n 0.00175687f $X=0.905 $Y=2.735 $X2=0
+ $Y2=0
cc_241 N_S1_M1025_g N_A_196_125#_c_934_n 0.00290482f $X=2.04 $Y=2.095 $X2=0
+ $Y2=0
cc_242 N_S1_c_229_n N_A_196_125#_c_932_n 0.00392226f $X=0.905 $Y=2.735 $X2=0
+ $Y2=0
cc_243 N_S1_c_230_n N_A_196_125#_c_936_n 0.00242118f $X=1.965 $Y=2.81 $X2=0
+ $Y2=0
cc_244 N_S1_M1025_g N_A_196_125#_c_936_n 0.00744254f $X=2.04 $Y=2.095 $X2=0
+ $Y2=0
cc_245 N_S1_c_227_n N_A_196_125#_c_936_n 0.0068727f $X=2.16 $Y=1.45 $X2=0 $Y2=0
cc_246 N_S1_c_230_n N_A_196_125#_c_937_n 0.00113835f $X=1.965 $Y=2.81 $X2=0
+ $Y2=0
cc_247 N_S1_M1025_g N_A_196_125#_c_937_n 8.24231e-19 $X=2.04 $Y=2.095 $X2=0
+ $Y2=0
cc_248 N_S1_c_229_n N_A_196_125#_c_938_n 0.00462484f $X=0.905 $Y=2.735 $X2=0
+ $Y2=0
cc_249 N_S1_c_230_n N_A_196_125#_c_938_n 0.00475074f $X=1.965 $Y=2.81 $X2=0
+ $Y2=0
cc_250 N_S1_M1025_g N_A_196_125#_c_938_n 3.47381e-19 $X=2.04 $Y=2.095 $X2=0
+ $Y2=0
cc_251 N_S1_c_227_n N_VPWR_M1025_d 0.00815547f $X=2.16 $Y=1.45 $X2=-0.19
+ $Y2=-0.245
cc_252 N_S1_c_230_n N_VPWR_c_1037_n 0.002253f $X=1.965 $Y=2.81 $X2=0 $Y2=0
cc_253 N_S1_c_230_n N_VPWR_c_1044_n 0.00965885f $X=1.965 $Y=2.81 $X2=0 $Y2=0
cc_254 N_S1_c_231_n N_VPWR_c_1044_n 0.00367387f $X=0.98 $Y=2.81 $X2=0 $Y2=0
cc_255 N_S1_c_230_n N_VPWR_c_1036_n 0.0138913f $X=1.965 $Y=2.81 $X2=0 $Y2=0
cc_256 N_S1_c_225_n N_VGND_c_1158_n 0.0478457f $X=0.55 $Y=0.18 $X2=0 $Y2=0
cc_257 N_S1_c_224_n N_VGND_c_1163_n 0.0464595f $X=2.245 $Y=0.18 $X2=0 $Y2=0
cc_258 N_S1_c_225_n N_VGND_c_1163_n 0.0111284f $X=0.55 $Y=0.18 $X2=0 $Y2=0
cc_259 N_S1_c_224_n N_VGND_c_1164_n 0.00661919f $X=2.245 $Y=0.18 $X2=0 $Y2=0
cc_260 N_A_110_125#_c_311_n N_A3_M1021_g 0.0233209f $X=3.335 $Y=1.352 $X2=0
+ $Y2=0
cc_261 N_A_110_125#_c_304_n N_A3_M1018_g 0.00995961f $X=3.375 $Y=1.185 $X2=0
+ $Y2=0
cc_262 N_A_110_125#_c_304_n A3 0.00144855f $X=3.375 $Y=1.185 $X2=0 $Y2=0
cc_263 N_A_110_125#_c_311_n A3 0.0144322f $X=3.335 $Y=1.352 $X2=0 $Y2=0
cc_264 N_A_110_125#_c_311_n N_A3_c_396_n 0.0103208f $X=3.335 $Y=1.352 $X2=0
+ $Y2=0
cc_265 N_A_110_125#_c_305_n N_A_27_125#_c_833_n 0.0751251f $X=0.69 $Y=0.835
+ $X2=0 $Y2=0
cc_266 N_A_110_125#_c_305_n N_A_27_125#_c_837_n 0.0167441f $X=0.69 $Y=0.835
+ $X2=0 $Y2=0
cc_267 N_A_110_125#_M1002_g N_A_27_125#_c_840_n 0.0149374f $X=2.905 $Y=2.405
+ $X2=0 $Y2=0
cc_268 N_A_110_125#_M1019_g N_A_27_125#_c_840_n 0.01447f $X=3.335 $Y=2.405 $X2=0
+ $Y2=0
cc_269 N_A_110_125#_c_306_n N_A_196_125#_c_931_n 0.0217876f $X=1.465 $Y=0.41
+ $X2=0 $Y2=0
cc_270 N_A_110_125#_c_310_n N_A_196_125#_c_931_n 0.0022182f $X=1.55 $Y=0.41
+ $X2=0 $Y2=0
cc_271 N_A_110_125#_c_305_n N_A_196_125#_c_932_n 0.0919721f $X=0.69 $Y=0.835
+ $X2=0 $Y2=0
cc_272 N_A_110_125#_M1002_g N_A_196_125#_c_936_n 0.00794997f $X=2.905 $Y=2.405
+ $X2=0 $Y2=0
cc_273 N_A_110_125#_M1019_g N_A_196_125#_c_936_n 0.00775984f $X=3.335 $Y=2.405
+ $X2=0 $Y2=0
cc_274 N_A_110_125#_c_305_n N_A_196_125#_c_937_n 0.00134725f $X=0.69 $Y=0.835
+ $X2=0 $Y2=0
cc_275 N_A_110_125#_M1002_g N_VPWR_c_1037_n 0.00968892f $X=2.905 $Y=2.405 $X2=0
+ $Y2=0
cc_276 N_A_110_125#_M1019_g N_VPWR_c_1037_n 0.0011441f $X=3.335 $Y=2.405 $X2=0
+ $Y2=0
cc_277 N_A_110_125#_M1002_g N_VPWR_c_1038_n 0.0011441f $X=2.905 $Y=2.405 $X2=0
+ $Y2=0
cc_278 N_A_110_125#_M1019_g N_VPWR_c_1038_n 0.00968892f $X=3.335 $Y=2.405 $X2=0
+ $Y2=0
cc_279 N_A_110_125#_M1002_g N_VPWR_c_1045_n 0.00323304f $X=2.905 $Y=2.405 $X2=0
+ $Y2=0
cc_280 N_A_110_125#_M1019_g N_VPWR_c_1045_n 0.00323304f $X=3.335 $Y=2.405 $X2=0
+ $Y2=0
cc_281 N_A_110_125#_M1002_g N_VPWR_c_1036_n 0.00406886f $X=2.905 $Y=2.405 $X2=0
+ $Y2=0
cc_282 N_A_110_125#_M1019_g N_VPWR_c_1036_n 0.00406886f $X=3.335 $Y=2.405 $X2=0
+ $Y2=0
cc_283 N_A_110_125#_M1002_g N_X_c_1133_n 0.00706232f $X=2.905 $Y=2.405 $X2=0
+ $Y2=0
cc_284 N_A_110_125#_c_302_n N_X_c_1133_n 0.00143199f $X=2.945 $Y=1.185 $X2=0
+ $Y2=0
cc_285 N_A_110_125#_M1019_g N_X_c_1133_n 0.00263751f $X=3.335 $Y=2.405 $X2=0
+ $Y2=0
cc_286 N_A_110_125#_c_304_n N_X_c_1133_n 0.00257599f $X=3.375 $Y=1.185 $X2=0
+ $Y2=0
cc_287 N_A_110_125#_c_309_n N_X_c_1133_n 0.0322241f $X=2.77 $Y=1.35 $X2=0 $Y2=0
cc_288 N_A_110_125#_c_311_n N_X_c_1133_n 0.0203312f $X=3.335 $Y=1.352 $X2=0
+ $Y2=0
cc_289 N_A_110_125#_c_308_n N_VGND_M1023_d 0.0111692f $X=2.605 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_290 N_A_110_125#_c_309_n N_VGND_M1023_d 0.0083679f $X=2.77 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_291 N_A_110_125#_c_302_n N_VGND_c_1155_n 6.98192e-19 $X=2.945 $Y=1.185 $X2=0
+ $Y2=0
cc_292 N_A_110_125#_c_304_n N_VGND_c_1155_n 0.0204725f $X=3.375 $Y=1.185 $X2=0
+ $Y2=0
cc_293 N_A_110_125#_c_306_n N_VGND_c_1158_n 0.0308545f $X=1.465 $Y=0.41 $X2=0
+ $Y2=0
cc_294 N_A_110_125#_c_307_n N_VGND_c_1158_n 0.0109032f $X=0.775 $Y=0.41 $X2=0
+ $Y2=0
cc_295 N_A_110_125#_c_308_n N_VGND_c_1158_n 0.0196388f $X=2.605 $Y=0.61 $X2=0
+ $Y2=0
cc_296 N_A_110_125#_c_310_n N_VGND_c_1158_n 0.00796697f $X=1.55 $Y=0.41 $X2=0
+ $Y2=0
cc_297 N_A_110_125#_c_302_n N_VGND_c_1159_n 0.00585385f $X=2.945 $Y=1.185 $X2=0
+ $Y2=0
cc_298 N_A_110_125#_c_304_n N_VGND_c_1159_n 0.00486043f $X=3.375 $Y=1.185 $X2=0
+ $Y2=0
cc_299 N_A_110_125#_c_302_n N_VGND_c_1163_n 0.0112095f $X=2.945 $Y=1.185 $X2=0
+ $Y2=0
cc_300 N_A_110_125#_c_304_n N_VGND_c_1163_n 0.00824727f $X=3.375 $Y=1.185 $X2=0
+ $Y2=0
cc_301 N_A_110_125#_c_306_n N_VGND_c_1163_n 0.022048f $X=1.465 $Y=0.41 $X2=0
+ $Y2=0
cc_302 N_A_110_125#_c_307_n N_VGND_c_1163_n 0.00736409f $X=0.775 $Y=0.41 $X2=0
+ $Y2=0
cc_303 N_A_110_125#_c_308_n N_VGND_c_1163_n 0.0265842f $X=2.605 $Y=0.61 $X2=0
+ $Y2=0
cc_304 N_A_110_125#_c_310_n N_VGND_c_1163_n 0.00550625f $X=1.55 $Y=0.41 $X2=0
+ $Y2=0
cc_305 N_A_110_125#_c_302_n N_VGND_c_1164_n 0.00253767f $X=2.945 $Y=1.185 $X2=0
+ $Y2=0
cc_306 N_A_110_125#_c_308_n N_VGND_c_1164_n 0.0255775f $X=2.605 $Y=0.61 $X2=0
+ $Y2=0
cc_307 N_A3_M1021_g N_A_859_351#_c_434_n 0.0113421f $X=4.01 $Y=2.415 $X2=0 $Y2=0
cc_308 A3 N_A_859_351#_c_434_n 0.00240913f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_309 N_A3_c_396_n N_A_859_351#_c_434_n 0.008588f $X=3.96 $Y=1.35 $X2=0 $Y2=0
cc_310 N_A3_M1021_g N_A_859_351#_c_457_n 0.0683863f $X=4.01 $Y=2.415 $X2=0 $Y2=0
cc_311 A3 N_A_859_351#_c_457_n 0.00321951f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_312 N_A3_M1018_g N_A_859_351#_c_448_n 0.00338251f $X=4.05 $Y=0.805 $X2=0
+ $Y2=0
cc_313 N_A3_M1018_g N_S0_M1009_g 0.0390122f $X=4.05 $Y=0.805 $X2=0 $Y2=0
cc_314 N_A3_M1021_g N_A_27_125#_c_840_n 0.0112617f $X=4.01 $Y=2.415 $X2=0 $Y2=0
cc_315 A3 N_A_27_125#_c_840_n 0.0428181f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_316 N_A3_M1021_g N_A_27_125#_c_834_n 5.83359e-19 $X=4.01 $Y=2.415 $X2=0 $Y2=0
cc_317 N_A3_M1018_g N_A_27_125#_c_834_n 0.00245784f $X=4.05 $Y=0.805 $X2=0 $Y2=0
cc_318 A3 N_A_27_125#_c_834_n 0.0723668f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_319 N_A3_M1018_g N_A_27_125#_c_835_n 8.38341e-19 $X=4.05 $Y=0.805 $X2=0 $Y2=0
cc_320 N_A3_M1021_g N_A_27_125#_c_843_n 0.00230415f $X=4.01 $Y=2.415 $X2=0 $Y2=0
cc_321 A3 N_A_27_125#_c_843_n 0.0152689f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_322 N_A3_M1021_g N_A_196_125#_c_936_n 0.00271399f $X=4.01 $Y=2.415 $X2=0
+ $Y2=0
cc_323 A3 N_A_196_125#_c_936_n 0.0210442f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_324 A3 N_VPWR_M1019_s 0.0103747f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_325 N_A3_M1021_g N_VPWR_c_1038_n 0.00194811f $X=4.01 $Y=2.415 $X2=0 $Y2=0
cc_326 N_A3_M1021_g N_VPWR_c_1046_n 0.00338502f $X=4.01 $Y=2.415 $X2=0 $Y2=0
cc_327 N_A3_M1021_g N_VPWR_c_1036_n 0.00477801f $X=4.01 $Y=2.415 $X2=0 $Y2=0
cc_328 A3 N_X_c_1133_n 0.0517781f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_329 N_A3_c_396_n N_X_c_1133_n 2.01051e-19 $X=3.96 $Y=1.35 $X2=0 $Y2=0
cc_330 A3 A_817_419# 0.00171177f $X=3.515 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_331 N_A3_M1018_g N_VGND_c_1155_n 0.0120367f $X=4.05 $Y=0.805 $X2=0 $Y2=0
cc_332 A3 N_VGND_c_1155_n 0.0484144f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_333 N_A3_c_396_n N_VGND_c_1155_n 0.00111517f $X=3.96 $Y=1.35 $X2=0 $Y2=0
cc_334 N_A3_M1018_g N_VGND_c_1160_n 0.00315482f $X=4.05 $Y=0.805 $X2=0 $Y2=0
cc_335 N_A3_M1018_g N_VGND_c_1163_n 0.00353573f $X=4.05 $Y=0.805 $X2=0 $Y2=0
cc_336 N_A_859_351#_M1026_g N_A2_c_593_n 7.71601e-19 $X=4.37 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_337 N_A_859_351#_c_457_n N_A2_c_593_n 0.0017767f $X=4.39 $Y=1.905 $X2=-0.19
+ $Y2=-0.245
cc_338 N_A_859_351#_c_441_n N_A2_c_593_n 0.00221614f $X=5.985 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_339 N_A_859_351#_M1011_g N_A2_M1020_g 0.0268535f $X=4.84 $Y=0.805 $X2=0 $Y2=0
cc_340 N_A_859_351#_c_441_n N_A2_M1020_g 0.0167849f $X=5.985 $Y=1.08 $X2=0 $Y2=0
cc_341 N_A_859_351#_c_442_n N_A2_M1020_g 9.00501e-19 $X=6.07 $Y=0.995 $X2=0
+ $Y2=0
cc_342 N_A_859_351#_c_447_n N_A2_M1020_g 0.00172867f $X=4.86 $Y=1.08 $X2=0 $Y2=0
cc_343 N_A_859_351#_c_448_n N_A2_M1020_g 0.0262896f $X=4.86 $Y=1.315 $X2=0 $Y2=0
cc_344 N_A_859_351#_c_433_n A2 0.00739066f $X=4.695 $Y=1.46 $X2=0 $Y2=0
cc_345 N_A_859_351#_c_440_n A2 0.00208652f $X=4.39 $Y=1.755 $X2=0 $Y2=0
cc_346 N_A_859_351#_c_441_n A2 0.0243706f $X=5.985 $Y=1.08 $X2=0 $Y2=0
cc_347 N_A_859_351#_c_447_n A2 0.0265037f $X=4.86 $Y=1.08 $X2=0 $Y2=0
cc_348 N_A_859_351#_c_441_n N_A1_M1007_g 0.00912571f $X=5.985 $Y=1.08 $X2=0
+ $Y2=0
cc_349 N_A_859_351#_c_442_n N_A1_M1007_g 0.0133592f $X=6.07 $Y=0.995 $X2=0 $Y2=0
cc_350 N_A_859_351#_c_451_n N_A1_M1007_g 0.00319853f $X=6.85 $Y=1.315 $X2=0
+ $Y2=0
cc_351 N_A_859_351#_M1027_g N_A1_c_645_n 0.0444976f $X=6.4 $Y=2.415 $X2=0 $Y2=0
cc_352 N_A_859_351#_c_438_n N_A1_c_641_n 0.0444976f $X=6.475 $Y=1.46 $X2=0 $Y2=0
cc_353 N_A_859_351#_c_441_n N_A1_c_641_n 0.00511067f $X=5.985 $Y=1.08 $X2=0
+ $Y2=0
cc_354 N_A_859_351#_c_438_n N_A1_c_642_n 0.00399921f $X=6.475 $Y=1.46 $X2=0
+ $Y2=0
cc_355 N_A_859_351#_c_441_n N_A1_c_642_n 0.0291805f $X=5.985 $Y=1.08 $X2=0 $Y2=0
cc_356 N_A_859_351#_M1001_g N_A0_M1004_g 0.0212588f $X=6.83 $Y=0.805 $X2=0 $Y2=0
cc_357 N_A_859_351#_c_445_n N_A0_M1004_g 0.0144177f $X=7.85 $Y=1.07 $X2=0 $Y2=0
cc_358 N_A_859_351#_c_449_n N_A0_M1004_g 0.00578001f $X=6.907 $Y=1.07 $X2=0
+ $Y2=0
cc_359 N_A_859_351#_c_450_n N_A0_M1004_g 0.00660503f $X=6.907 $Y=0.985 $X2=0
+ $Y2=0
cc_360 N_A_859_351#_c_451_n N_A0_M1004_g 0.0247407f $X=6.85 $Y=1.315 $X2=0 $Y2=0
cc_361 N_A_859_351#_M1027_g A0 0.00203811f $X=6.4 $Y=2.415 $X2=0 $Y2=0
cc_362 N_A_859_351#_c_445_n A0 0.0195344f $X=7.85 $Y=1.07 $X2=0 $Y2=0
cc_363 N_A_859_351#_c_449_n A0 0.036447f $X=6.907 $Y=1.07 $X2=0 $Y2=0
cc_364 N_A_859_351#_c_451_n A0 0.00705699f $X=6.85 $Y=1.315 $X2=0 $Y2=0
cc_365 N_A_859_351#_c_445_n N_A0_c_686_n 9.69765e-19 $X=7.85 $Y=1.07 $X2=0 $Y2=0
cc_366 N_A_859_351#_c_434_n N_S0_M1009_g 0.00851793f $X=4.485 $Y=1.46 $X2=0
+ $Y2=0
cc_367 N_A_859_351#_M1011_g N_S0_M1009_g 0.0160762f $X=4.84 $Y=0.805 $X2=0 $Y2=0
cc_368 N_A_859_351#_c_447_n N_S0_M1009_g 4.98735e-19 $X=4.86 $Y=1.08 $X2=0 $Y2=0
cc_369 N_A_859_351#_M1011_g N_S0_c_721_n 0.0102931f $X=4.84 $Y=0.805 $X2=0 $Y2=0
cc_370 N_A_859_351#_c_443_n N_S0_c_721_n 0.00186516f $X=6.96 $Y=0.35 $X2=0 $Y2=0
cc_371 N_A_859_351#_c_444_n N_S0_c_721_n 0.00203407f $X=6.155 $Y=0.35 $X2=0
+ $Y2=0
cc_372 N_A_859_351#_M1026_g N_S0_M1012_g 0.0119481f $X=4.37 $Y=2.415 $X2=0 $Y2=0
cc_373 N_A_859_351#_c_448_n N_S0_M1012_g 0.00343455f $X=4.86 $Y=1.315 $X2=0
+ $Y2=0
cc_374 N_A_859_351#_M1027_g N_S0_c_730_n 0.00975027f $X=6.4 $Y=2.415 $X2=0 $Y2=0
cc_375 N_A_859_351#_c_438_n N_S0_M1000_g 0.00852163f $X=6.475 $Y=1.46 $X2=0
+ $Y2=0
cc_376 N_A_859_351#_M1001_g N_S0_M1000_g 0.0156566f $X=6.83 $Y=0.805 $X2=0 $Y2=0
cc_377 N_A_859_351#_c_441_n N_S0_M1000_g 8.01099e-19 $X=5.985 $Y=1.08 $X2=0
+ $Y2=0
cc_378 N_A_859_351#_c_442_n N_S0_M1000_g 0.00460997f $X=6.07 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_859_351#_c_443_n N_S0_M1000_g 0.01352f $X=6.96 $Y=0.35 $X2=0 $Y2=0
cc_380 N_A_859_351#_c_449_n N_S0_M1000_g 5.38308e-19 $X=6.907 $Y=1.07 $X2=0
+ $Y2=0
cc_381 N_A_859_351#_c_450_n N_S0_M1000_g 9.69912e-19 $X=6.907 $Y=0.985 $X2=0
+ $Y2=0
cc_382 N_A_859_351#_M1001_g N_S0_c_724_n 0.00881852f $X=6.83 $Y=0.805 $X2=0
+ $Y2=0
cc_383 N_A_859_351#_c_443_n N_S0_c_724_n 0.0109268f $X=6.96 $Y=0.35 $X2=0 $Y2=0
cc_384 N_A_859_351#_M1027_g N_S0_M1014_g 0.0085797f $X=6.4 $Y=2.415 $X2=0 $Y2=0
cc_385 N_A_859_351#_c_451_n N_S0_M1014_g 0.00340313f $X=6.85 $Y=1.315 $X2=0
+ $Y2=0
cc_386 N_A_859_351#_c_443_n N_S0_M1006_g 7.22755e-19 $X=6.96 $Y=0.35 $X2=0 $Y2=0
cc_387 N_A_859_351#_c_445_n N_S0_M1006_g 0.0192505f $X=7.85 $Y=1.07 $X2=0 $Y2=0
cc_388 N_A_859_351#_c_453_n N_S0_M1006_g 0.00143639f $X=8.227 $Y=2.075 $X2=0
+ $Y2=0
cc_389 N_A_859_351#_c_458_n N_S0_M1008_g 8.98903e-19 $X=8.08 $Y=2.24 $X2=0 $Y2=0
cc_390 N_A_859_351#_c_453_n N_S0_M1008_g 0.00416864f $X=8.227 $Y=2.075 $X2=0
+ $Y2=0
cc_391 N_A_859_351#_c_445_n N_S0_c_727_n 0.00134638f $X=7.85 $Y=1.07 $X2=0 $Y2=0
cc_392 N_A_859_351#_c_446_n N_S0_c_727_n 3.13014e-19 $X=8.3 $Y=1.07 $X2=0 $Y2=0
cc_393 N_A_859_351#_c_452_n N_S0_c_727_n 0.00799241f $X=7.98 $Y=1.07 $X2=0 $Y2=0
cc_394 N_A_859_351#_c_453_n N_S0_c_727_n 0.0179558f $X=8.227 $Y=2.075 $X2=0
+ $Y2=0
cc_395 N_A_859_351#_c_458_n N_S0_c_736_n 0.00373925f $X=8.08 $Y=2.24 $X2=0 $Y2=0
cc_396 N_A_859_351#_c_445_n N_S0_c_769_n 0.00456501f $X=7.85 $Y=1.07 $X2=0 $Y2=0
cc_397 N_A_859_351#_c_446_n N_S0_c_769_n 6.72306e-19 $X=8.3 $Y=1.07 $X2=0 $Y2=0
cc_398 N_A_859_351#_c_449_n N_S0_c_769_n 0.0021367f $X=6.907 $Y=1.07 $X2=0 $Y2=0
cc_399 N_A_859_351#_c_452_n N_S0_c_769_n 0.0224195f $X=7.98 $Y=1.07 $X2=0 $Y2=0
cc_400 N_A_859_351#_c_458_n N_S0_c_769_n 0.0117087f $X=8.08 $Y=2.24 $X2=0 $Y2=0
cc_401 N_A_859_351#_c_453_n N_S0_c_769_n 0.0416816f $X=8.227 $Y=2.075 $X2=0
+ $Y2=0
cc_402 N_A_859_351#_c_447_n N_A_27_125#_M1009_d 3.08127e-19 $X=4.86 $Y=1.08
+ $X2=0 $Y2=0
cc_403 N_A_859_351#_M1026_g N_A_27_125#_c_840_n 0.00451192f $X=4.37 $Y=2.415
+ $X2=0 $Y2=0
cc_404 N_A_859_351#_M1026_g N_A_27_125#_c_834_n 0.0037981f $X=4.37 $Y=2.415
+ $X2=0 $Y2=0
cc_405 N_A_859_351#_c_433_n N_A_27_125#_c_834_n 0.00757469f $X=4.695 $Y=1.46
+ $X2=0 $Y2=0
cc_406 N_A_859_351#_c_434_n N_A_27_125#_c_834_n 0.00412987f $X=4.485 $Y=1.46
+ $X2=0 $Y2=0
cc_407 N_A_859_351#_M1011_g N_A_27_125#_c_834_n 3.7941e-19 $X=4.84 $Y=0.805
+ $X2=0 $Y2=0
cc_408 N_A_859_351#_c_440_n N_A_27_125#_c_834_n 0.00706586f $X=4.39 $Y=1.755
+ $X2=0 $Y2=0
cc_409 N_A_859_351#_c_457_n N_A_27_125#_c_834_n 0.00536489f $X=4.39 $Y=1.905
+ $X2=0 $Y2=0
cc_410 N_A_859_351#_c_447_n N_A_27_125#_c_834_n 0.0289506f $X=4.86 $Y=1.08 $X2=0
+ $Y2=0
cc_411 N_A_859_351#_c_448_n N_A_27_125#_c_834_n 0.00221854f $X=4.86 $Y=1.315
+ $X2=0 $Y2=0
cc_412 N_A_859_351#_c_433_n N_A_27_125#_c_835_n 0.00397405f $X=4.695 $Y=1.46
+ $X2=0 $Y2=0
cc_413 N_A_859_351#_M1011_g N_A_27_125#_c_835_n 0.00602075f $X=4.84 $Y=0.805
+ $X2=0 $Y2=0
cc_414 N_A_859_351#_c_447_n N_A_27_125#_c_835_n 0.00281082f $X=4.86 $Y=1.08
+ $X2=0 $Y2=0
cc_415 N_A_859_351#_c_448_n N_A_27_125#_c_835_n 2.41782e-19 $X=4.86 $Y=1.315
+ $X2=0 $Y2=0
cc_416 N_A_859_351#_M1026_g N_A_27_125#_c_843_n 0.0135794f $X=4.37 $Y=2.415
+ $X2=0 $Y2=0
cc_417 N_A_859_351#_c_433_n N_A_27_125#_c_843_n 0.00476349f $X=4.695 $Y=1.46
+ $X2=0 $Y2=0
cc_418 N_A_859_351#_c_449_n N_A_196_125#_M1000_d 3.9346e-19 $X=6.907 $Y=1.07
+ $X2=0 $Y2=0
cc_419 N_A_859_351#_c_437_n N_A_196_125#_c_975_n 0.00373058f $X=6.685 $Y=1.46
+ $X2=0 $Y2=0
cc_420 N_A_859_351#_M1001_g N_A_196_125#_c_975_n 0.00269774f $X=6.83 $Y=0.805
+ $X2=0 $Y2=0
cc_421 N_A_859_351#_c_443_n N_A_196_125#_c_975_n 0.026793f $X=6.96 $Y=0.35 $X2=0
+ $Y2=0
cc_422 N_A_859_351#_c_449_n N_A_196_125#_c_975_n 0.00277344f $X=6.907 $Y=1.07
+ $X2=0 $Y2=0
cc_423 N_A_859_351#_c_451_n N_A_196_125#_c_975_n 2.35593e-19 $X=6.85 $Y=1.315
+ $X2=0 $Y2=0
cc_424 N_A_859_351#_M1026_g N_A_196_125#_c_936_n 0.00254147f $X=4.37 $Y=2.415
+ $X2=0 $Y2=0
cc_425 N_A_859_351#_M1027_g N_A_196_125#_c_936_n 0.00122262f $X=6.4 $Y=2.415
+ $X2=0 $Y2=0
cc_426 N_A_859_351#_M1027_g N_A_196_125#_c_982_n 9.02358e-19 $X=6.4 $Y=2.415
+ $X2=0 $Y2=0
cc_427 N_A_859_351#_M1027_g N_A_196_125#_c_939_n 0.0163379f $X=6.4 $Y=2.415
+ $X2=0 $Y2=0
cc_428 N_A_859_351#_c_437_n N_A_196_125#_c_939_n 0.00497036f $X=6.685 $Y=1.46
+ $X2=0 $Y2=0
cc_429 N_A_859_351#_M1027_g N_A_196_125#_c_933_n 0.0165019f $X=6.4 $Y=2.415
+ $X2=0 $Y2=0
cc_430 N_A_859_351#_c_437_n N_A_196_125#_c_933_n 0.00820996f $X=6.685 $Y=1.46
+ $X2=0 $Y2=0
cc_431 N_A_859_351#_c_438_n N_A_196_125#_c_933_n 0.00409786f $X=6.475 $Y=1.46
+ $X2=0 $Y2=0
cc_432 N_A_859_351#_M1001_g N_A_196_125#_c_933_n 3.85539e-19 $X=6.83 $Y=0.805
+ $X2=0 $Y2=0
cc_433 N_A_859_351#_c_441_n N_A_196_125#_c_933_n 0.0123251f $X=5.985 $Y=1.08
+ $X2=0 $Y2=0
cc_434 N_A_859_351#_c_449_n N_A_196_125#_c_933_n 0.0314783f $X=6.907 $Y=1.07
+ $X2=0 $Y2=0
cc_435 N_A_859_351#_c_451_n N_A_196_125#_c_933_n 0.00223968f $X=6.85 $Y=1.315
+ $X2=0 $Y2=0
cc_436 N_A_859_351#_M1027_g N_VPWR_c_1039_n 0.00104291f $X=6.4 $Y=2.415 $X2=0
+ $Y2=0
cc_437 N_A_859_351#_M1027_g N_VPWR_c_1040_n 7.57905e-19 $X=6.4 $Y=2.415 $X2=0
+ $Y2=0
cc_438 N_A_859_351#_c_458_n N_VPWR_c_1041_n 0.0255585f $X=8.08 $Y=2.24 $X2=0
+ $Y2=0
cc_439 N_A_859_351#_M1026_g N_VPWR_c_1046_n 0.00336978f $X=4.37 $Y=2.415 $X2=0
+ $Y2=0
cc_440 N_A_859_351#_c_458_n N_VPWR_c_1047_n 0.0108825f $X=8.08 $Y=2.24 $X2=0
+ $Y2=0
cc_441 N_A_859_351#_M1026_g N_VPWR_c_1036_n 0.00477801f $X=4.37 $Y=2.415 $X2=0
+ $Y2=0
cc_442 N_A_859_351#_M1027_g N_VPWR_c_1036_n 9.39239e-19 $X=6.4 $Y=2.415 $X2=0
+ $Y2=0
cc_443 N_A_859_351#_c_458_n N_VPWR_c_1036_n 0.0151975f $X=8.08 $Y=2.24 $X2=0
+ $Y2=0
cc_444 N_A_859_351#_c_441_n N_VGND_M1020_d 0.00898353f $X=5.985 $Y=1.08 $X2=0
+ $Y2=0
cc_445 N_A_859_351#_c_445_n N_VGND_M1004_d 0.00176461f $X=7.85 $Y=1.07 $X2=0
+ $Y2=0
cc_446 N_A_859_351#_c_441_n N_VGND_c_1156_n 0.0266856f $X=5.985 $Y=1.08 $X2=0
+ $Y2=0
cc_447 N_A_859_351#_c_442_n N_VGND_c_1156_n 0.029175f $X=6.07 $Y=0.995 $X2=0
+ $Y2=0
cc_448 N_A_859_351#_c_444_n N_VGND_c_1156_n 0.0150384f $X=6.155 $Y=0.35 $X2=0
+ $Y2=0
cc_449 N_A_859_351#_c_443_n N_VGND_c_1157_n 0.0125438f $X=6.96 $Y=0.35 $X2=0
+ $Y2=0
cc_450 N_A_859_351#_c_445_n N_VGND_c_1157_n 0.0170777f $X=7.85 $Y=1.07 $X2=0
+ $Y2=0
cc_451 N_A_859_351#_c_450_n N_VGND_c_1157_n 0.0233254f $X=6.907 $Y=0.985 $X2=0
+ $Y2=0
cc_452 N_A_859_351#_c_443_n N_VGND_c_1161_n 0.059773f $X=6.96 $Y=0.35 $X2=0
+ $Y2=0
cc_453 N_A_859_351#_c_444_n N_VGND_c_1161_n 0.0114574f $X=6.155 $Y=0.35 $X2=0
+ $Y2=0
cc_454 N_A_859_351#_c_584_p N_VGND_c_1162_n 0.00472305f $X=7.945 $Y=0.805 $X2=0
+ $Y2=0
cc_455 N_A_859_351#_M1011_g N_VGND_c_1163_n 9.39239e-19 $X=4.84 $Y=0.805 $X2=0
+ $Y2=0
cc_456 N_A_859_351#_c_443_n N_VGND_c_1163_n 0.0326189f $X=6.96 $Y=0.35 $X2=0
+ $Y2=0
cc_457 N_A_859_351#_c_444_n N_VGND_c_1163_n 0.00589978f $X=6.155 $Y=0.35 $X2=0
+ $Y2=0
cc_458 N_A_859_351#_c_584_p N_VGND_c_1163_n 0.00770078f $X=7.945 $Y=0.805 $X2=0
+ $Y2=0
cc_459 N_A_859_351#_c_441_n A_983_119# 0.00588299f $X=5.985 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_460 N_A_859_351#_c_447_n A_983_119# 0.00225111f $X=4.86 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_461 N_A_859_351#_c_445_n A_1381_119# 0.00152126f $X=7.85 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_462 N_A_859_351#_c_450_n A_1381_119# 0.00581753f $X=6.907 $Y=0.985 $X2=-0.19
+ $Y2=-0.245
cc_463 N_A2_M1020_g N_A1_M1007_g 0.0127972f $X=5.31 $Y=0.805 $X2=0 $Y2=0
cc_464 N_A2_c_593_n N_A1_c_640_n 0.0195762f $X=5.16 $Y=1.925 $X2=0 $Y2=0
cc_465 A2 N_A1_c_640_n 0.00212926f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_466 N_A2_M1010_g N_A1_c_645_n 2.30152e-19 $X=5.16 $Y=2.415 $X2=0 $Y2=0
cc_467 N_A2_c_593_n N_A1_c_641_n 0.00739747f $X=5.16 $Y=1.925 $X2=0 $Y2=0
cc_468 N_A2_M1020_g N_A1_c_641_n 0.00443729f $X=5.31 $Y=0.805 $X2=0 $Y2=0
cc_469 N_A2_c_593_n N_A1_c_642_n 0.00163484f $X=5.16 $Y=1.925 $X2=0 $Y2=0
cc_470 N_A2_M1010_g N_A1_c_642_n 0.00373044f $X=5.16 $Y=2.415 $X2=0 $Y2=0
cc_471 N_A2_M1020_g N_A1_c_642_n 2.26322e-19 $X=5.31 $Y=0.805 $X2=0 $Y2=0
cc_472 A2 N_A1_c_642_n 0.0283184f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_473 N_A2_M1020_g N_S0_c_721_n 0.0104164f $X=5.31 $Y=0.805 $X2=0 $Y2=0
cc_474 N_A2_M1010_g N_S0_M1012_g 0.0540146f $X=5.16 $Y=2.415 $X2=0 $Y2=0
cc_475 A2 N_S0_M1012_g 0.00422526f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_476 N_A2_M1010_g N_S0_c_730_n 0.0102164f $X=5.16 $Y=2.415 $X2=0 $Y2=0
cc_477 N_A2_c_593_n N_A_27_125#_c_834_n 0.00126931f $X=5.16 $Y=1.925 $X2=0 $Y2=0
cc_478 A2 N_A_27_125#_c_834_n 0.0281199f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_479 N_A2_M1020_g N_A_27_125#_c_835_n 0.00123354f $X=5.31 $Y=0.805 $X2=0 $Y2=0
cc_480 N_A2_M1010_g N_A_27_125#_c_843_n 0.00190446f $X=5.16 $Y=2.415 $X2=0 $Y2=0
cc_481 A2 N_A_27_125#_c_843_n 0.00539238f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_482 N_A2_M1010_g N_A_196_125#_c_936_n 0.00465507f $X=5.16 $Y=2.415 $X2=0
+ $Y2=0
cc_483 A2 N_A_196_125#_c_936_n 0.0182915f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_484 N_A2_c_593_n N_VPWR_c_1039_n 0.00847898f $X=5.16 $Y=1.925 $X2=0 $Y2=0
cc_485 N_A2_M1010_g N_VPWR_c_1039_n 0.0098321f $X=5.16 $Y=2.415 $X2=0 $Y2=0
cc_486 A2 N_VPWR_c_1039_n 0.0295724f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_487 N_A2_M1010_g N_VPWR_c_1040_n 0.00659371f $X=5.16 $Y=2.415 $X2=0 $Y2=0
cc_488 N_A2_M1010_g N_VPWR_c_1036_n 7.88961e-19 $X=5.16 $Y=2.415 $X2=0 $Y2=0
cc_489 N_A2_M1020_g N_VGND_c_1156_n 0.0103875f $X=5.31 $Y=0.805 $X2=0 $Y2=0
cc_490 N_A2_M1020_g N_VGND_c_1163_n 9.39239e-19 $X=5.31 $Y=0.805 $X2=0 $Y2=0
cc_491 N_A1_M1007_g N_S0_c_721_n 0.0090126f $X=6.04 $Y=0.805 $X2=0 $Y2=0
cc_492 N_A1_M1022_g N_S0_c_730_n 0.0102164f $X=6.04 $Y=2.415 $X2=0 $Y2=0
cc_493 N_A1_M1007_g N_S0_M1000_g 0.0400266f $X=6.04 $Y=0.805 $X2=0 $Y2=0
cc_494 N_A1_M1007_g N_A_196_125#_c_975_n 2.3876e-19 $X=6.04 $Y=0.805 $X2=0 $Y2=0
cc_495 N_A1_M1022_g N_A_196_125#_c_936_n 0.00429743f $X=6.04 $Y=2.415 $X2=0
+ $Y2=0
cc_496 N_A1_c_642_n N_A_196_125#_c_936_n 0.00935871f $X=5.95 $Y=1.43 $X2=0 $Y2=0
cc_497 N_A1_M1022_g N_A_196_125#_c_982_n 4.68315e-19 $X=6.04 $Y=2.415 $X2=0
+ $Y2=0
cc_498 N_A1_M1022_g N_A_196_125#_c_939_n 0.00277909f $X=6.04 $Y=2.415 $X2=0
+ $Y2=0
cc_499 N_A1_c_645_n N_A_196_125#_c_939_n 4.1052e-19 $X=5.95 $Y=1.935 $X2=0 $Y2=0
cc_500 N_A1_M1007_g N_A_196_125#_c_933_n 0.00453772f $X=6.04 $Y=0.805 $X2=0
+ $Y2=0
cc_501 N_A1_c_641_n N_A_196_125#_c_933_n 5.49051e-19 $X=5.95 $Y=1.43 $X2=0 $Y2=0
cc_502 N_A1_c_642_n N_A_196_125#_c_933_n 0.0586809f $X=5.95 $Y=1.43 $X2=0 $Y2=0
cc_503 N_A1_c_642_n N_VPWR_M1010_d 0.00152826f $X=5.95 $Y=1.43 $X2=0 $Y2=0
cc_504 N_A1_M1022_g N_VPWR_c_1039_n 0.0105419f $X=6.04 $Y=2.415 $X2=0 $Y2=0
cc_505 N_A1_c_645_n N_VPWR_c_1039_n 7.89247e-19 $X=5.95 $Y=1.935 $X2=0 $Y2=0
cc_506 N_A1_c_642_n N_VPWR_c_1039_n 0.01483f $X=5.95 $Y=1.43 $X2=0 $Y2=0
cc_507 N_A1_M1022_g N_VPWR_c_1040_n 0.00778676f $X=6.04 $Y=2.415 $X2=0 $Y2=0
cc_508 N_A1_M1022_g N_VPWR_c_1036_n 7.88961e-19 $X=6.04 $Y=2.415 $X2=0 $Y2=0
cc_509 N_A1_M1007_g N_VGND_c_1156_n 0.00327014f $X=6.04 $Y=0.805 $X2=0 $Y2=0
cc_510 N_A0_M1004_g N_S0_c_724_n 0.0103107f $X=7.3 $Y=0.805 $X2=0 $Y2=0
cc_511 N_A0_M1016_g N_S0_M1014_g 0.0291078f $X=7.435 $Y=2.415 $X2=0 $Y2=0
cc_512 A0 N_S0_M1014_g 0.00429439f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_513 N_A0_M1016_g N_S0_c_733_n 0.0103107f $X=7.435 $Y=2.415 $X2=0 $Y2=0
cc_514 N_A0_M1004_g N_S0_M1006_g 0.026641f $X=7.3 $Y=0.805 $X2=0 $Y2=0
cc_515 N_A0_M1016_g N_S0_M1008_g 0.0138521f $X=7.435 $Y=2.415 $X2=0 $Y2=0
cc_516 N_A0_M1004_g N_S0_c_728_n 0.00718654f $X=7.3 $Y=0.805 $X2=0 $Y2=0
cc_517 A0 N_S0_c_728_n 0.00190235f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_518 N_A0_c_686_n N_S0_c_728_n 0.018462f $X=7.39 $Y=1.77 $X2=0 $Y2=0
cc_519 N_A0_M1004_g N_S0_c_769_n 0.00126003f $X=7.3 $Y=0.805 $X2=0 $Y2=0
cc_520 A0 N_S0_c_769_n 0.0238286f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_521 N_A0_c_686_n N_S0_c_769_n 6.3357e-19 $X=7.39 $Y=1.77 $X2=0 $Y2=0
cc_522 A0 N_A_196_125#_c_939_n 0.0105027f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_523 A0 N_A_196_125#_c_933_n 0.0239914f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_524 N_A0_M1016_g N_VPWR_c_1041_n 0.0176657f $X=7.435 $Y=2.415 $X2=0 $Y2=0
cc_525 A0 N_VPWR_c_1041_n 0.00908623f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_526 N_A0_c_686_n N_VPWR_c_1041_n 0.00111947f $X=7.39 $Y=1.77 $X2=0 $Y2=0
cc_527 N_A0_M1016_g N_VPWR_c_1036_n 7.88961e-19 $X=7.435 $Y=2.415 $X2=0 $Y2=0
cc_528 N_A0_M1004_g N_VGND_c_1157_n 0.00602979f $X=7.3 $Y=0.805 $X2=0 $Y2=0
cc_529 N_A0_M1004_g N_VGND_c_1163_n 7.88961e-19 $X=7.3 $Y=0.805 $X2=0 $Y2=0
cc_530 N_S0_M1009_g N_A_27_125#_c_834_n 0.0101861f $X=4.41 $Y=0.805 $X2=0 $Y2=0
cc_531 N_S0_M1012_g N_A_27_125#_c_834_n 0.00215034f $X=4.8 $Y=2.415 $X2=0 $Y2=0
cc_532 N_S0_M1009_g N_A_27_125#_c_835_n 0.0090867f $X=4.41 $Y=0.805 $X2=0 $Y2=0
cc_533 N_S0_c_721_n N_A_27_125#_c_835_n 0.00372486f $X=6.325 $Y=0.18 $X2=0 $Y2=0
cc_534 N_S0_M1012_g N_A_27_125#_c_843_n 0.0111771f $X=4.8 $Y=2.415 $X2=0 $Y2=0
cc_535 N_S0_M1000_g N_A_196_125#_c_975_n 0.00602476f $X=6.4 $Y=0.805 $X2=0 $Y2=0
cc_536 N_S0_M1012_g N_A_196_125#_c_936_n 0.00735328f $X=4.8 $Y=2.415 $X2=0 $Y2=0
cc_537 N_S0_c_730_n N_A_196_125#_c_936_n 0.00629547f $X=6.85 $Y=3.15 $X2=0 $Y2=0
cc_538 N_S0_c_730_n N_A_196_125#_c_939_n 0.00611088f $X=6.85 $Y=3.15 $X2=0 $Y2=0
cc_539 N_S0_M1014_g N_A_196_125#_c_939_n 6.49221e-19 $X=6.925 $Y=2.415 $X2=0
+ $Y2=0
cc_540 N_S0_M1000_g N_A_196_125#_c_933_n 0.00873301f $X=6.4 $Y=0.805 $X2=0 $Y2=0
cc_541 N_S0_M1014_g N_A_196_125#_c_933_n 0.00195617f $X=6.925 $Y=2.415 $X2=0
+ $Y2=0
cc_542 N_S0_M1012_g N_VPWR_c_1039_n 0.00173701f $X=4.8 $Y=2.415 $X2=0 $Y2=0
cc_543 N_S0_M1012_g N_VPWR_c_1040_n 0.00798893f $X=4.8 $Y=2.415 $X2=0 $Y2=0
cc_544 N_S0_c_730_n N_VPWR_c_1040_n 0.0506993f $X=6.85 $Y=3.15 $X2=0 $Y2=0
cc_545 N_S0_M1014_g N_VPWR_c_1041_n 0.00821197f $X=6.925 $Y=2.415 $X2=0 $Y2=0
cc_546 N_S0_c_733_n N_VPWR_c_1041_n 0.0222995f $X=7.79 $Y=3.15 $X2=0 $Y2=0
cc_547 N_S0_M1008_g N_VPWR_c_1041_n 0.0274944f $X=7.865 $Y=2.415 $X2=0 $Y2=0
cc_548 N_S0_c_769_n N_VPWR_c_1041_n 0.00183649f $X=7.955 $Y=1.42 $X2=0 $Y2=0
cc_549 N_S0_c_730_n N_VPWR_c_1042_n 0.0484017f $X=6.85 $Y=3.15 $X2=0 $Y2=0
cc_550 N_S0_c_731_n N_VPWR_c_1046_n 0.0176953f $X=4.875 $Y=3.15 $X2=0 $Y2=0
cc_551 N_S0_c_733_n N_VPWR_c_1047_n 0.00486043f $X=7.79 $Y=3.15 $X2=0 $Y2=0
cc_552 N_S0_c_730_n N_VPWR_c_1036_n 0.0457369f $X=6.85 $Y=3.15 $X2=0 $Y2=0
cc_553 N_S0_c_731_n N_VPWR_c_1036_n 0.0107579f $X=4.875 $Y=3.15 $X2=0 $Y2=0
cc_554 N_S0_c_733_n N_VPWR_c_1036_n 0.0336313f $X=7.79 $Y=3.15 $X2=0 $Y2=0
cc_555 N_S0_c_735_n N_VPWR_c_1036_n 0.00926736f $X=6.925 $Y=3.15 $X2=0 $Y2=0
cc_556 N_S0_M1009_g N_VGND_c_1155_n 0.00157608f $X=4.41 $Y=0.805 $X2=0 $Y2=0
cc_557 N_S0_c_722_n N_VGND_c_1155_n 0.011006f $X=4.485 $Y=0.18 $X2=0 $Y2=0
cc_558 N_S0_c_721_n N_VGND_c_1156_n 0.025825f $X=6.325 $Y=0.18 $X2=0 $Y2=0
cc_559 N_S0_M1000_g N_VGND_c_1156_n 9.2728e-19 $X=6.4 $Y=0.805 $X2=0 $Y2=0
cc_560 N_S0_c_724_n N_VGND_c_1157_n 0.0220925f $X=7.655 $Y=0.18 $X2=0 $Y2=0
cc_561 N_S0_M1006_g N_VGND_c_1157_n 0.0245966f $X=7.73 $Y=0.805 $X2=0 $Y2=0
cc_562 N_S0_c_722_n N_VGND_c_1160_n 0.0363768f $X=4.485 $Y=0.18 $X2=0 $Y2=0
cc_563 N_S0_c_721_n N_VGND_c_1161_n 0.0381236f $X=6.325 $Y=0.18 $X2=0 $Y2=0
cc_564 N_S0_c_724_n N_VGND_c_1162_n 0.00486043f $X=7.655 $Y=0.18 $X2=0 $Y2=0
cc_565 N_S0_c_721_n N_VGND_c_1163_n 0.0563285f $X=6.325 $Y=0.18 $X2=0 $Y2=0
cc_566 N_S0_c_722_n N_VGND_c_1163_n 0.00681298f $X=4.485 $Y=0.18 $X2=0 $Y2=0
cc_567 N_S0_c_724_n N_VGND_c_1163_n 0.0342301f $X=7.655 $Y=0.18 $X2=0 $Y2=0
cc_568 N_S0_c_726_n N_VGND_c_1163_n 0.00370104f $X=6.4 $Y=0.18 $X2=0 $Y2=0
cc_569 N_A_27_125#_c_837_n N_A_196_125#_c_936_n 0.00414374f $X=1.465 $Y=2.9
+ $X2=0 $Y2=0
cc_570 N_A_27_125#_c_840_n N_A_196_125#_c_936_n 0.139246f $X=4.345 $Y=2.52 $X2=0
+ $Y2=0
cc_571 N_A_27_125#_c_841_n N_A_196_125#_c_936_n 0.00707712f $X=1.635 $Y=2.52
+ $X2=0 $Y2=0
cc_572 N_A_27_125#_c_843_n N_A_196_125#_c_936_n 0.0474282f $X=4.585 $Y=2.24
+ $X2=0 $Y2=0
cc_573 N_A_27_125#_c_837_n N_A_196_125#_c_937_n 0.00336616f $X=1.465 $Y=2.9
+ $X2=0 $Y2=0
cc_574 N_A_27_125#_c_841_n N_A_196_125#_c_937_n 0.00140753f $X=1.635 $Y=2.52
+ $X2=0 $Y2=0
cc_575 N_A_27_125#_c_837_n N_A_196_125#_c_938_n 0.0153855f $X=1.465 $Y=2.9 $X2=0
+ $Y2=0
cc_576 N_A_27_125#_c_841_n N_A_196_125#_c_938_n 0.0111103f $X=1.635 $Y=2.52
+ $X2=0 $Y2=0
cc_577 N_A_27_125#_c_840_n N_VPWR_M1025_d 0.00654096f $X=4.345 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_578 N_A_27_125#_c_840_n N_VPWR_M1019_s 0.0092167f $X=4.345 $Y=2.52 $X2=0
+ $Y2=0
cc_579 N_A_27_125#_c_840_n N_VPWR_c_1037_n 0.0184364f $X=4.345 $Y=2.52 $X2=0
+ $Y2=0
cc_580 N_A_27_125#_c_840_n N_VPWR_c_1038_n 0.0183881f $X=4.345 $Y=2.52 $X2=0
+ $Y2=0
cc_581 N_A_27_125#_c_843_n N_VPWR_c_1039_n 0.0190693f $X=4.585 $Y=2.24 $X2=0
+ $Y2=0
cc_582 N_A_27_125#_c_843_n N_VPWR_c_1040_n 0.0022889f $X=4.585 $Y=2.24 $X2=0
+ $Y2=0
cc_583 N_A_27_125#_c_837_n N_VPWR_c_1044_n 0.0520412f $X=1.465 $Y=2.9 $X2=0
+ $Y2=0
cc_584 N_A_27_125#_c_838_n N_VPWR_c_1044_n 0.0131604f $X=0.385 $Y=2.9 $X2=0
+ $Y2=0
cc_585 N_A_27_125#_c_840_n N_VPWR_c_1044_n 0.0132112f $X=4.345 $Y=2.52 $X2=0
+ $Y2=0
cc_586 N_A_27_125#_c_840_n N_VPWR_c_1045_n 0.00660734f $X=4.345 $Y=2.52 $X2=0
+ $Y2=0
cc_587 N_A_27_125#_c_840_n N_VPWR_c_1046_n 0.00772706f $X=4.345 $Y=2.52 $X2=0
+ $Y2=0
cc_588 N_A_27_125#_c_843_n N_VPWR_c_1046_n 0.00841306f $X=4.585 $Y=2.24 $X2=0
+ $Y2=0
cc_589 N_A_27_125#_c_837_n N_VPWR_c_1036_n 0.044565f $X=1.465 $Y=2.9 $X2=0 $Y2=0
cc_590 N_A_27_125#_c_838_n N_VPWR_c_1036_n 0.0107298f $X=0.385 $Y=2.9 $X2=0
+ $Y2=0
cc_591 N_A_27_125#_c_840_n N_VPWR_c_1036_n 0.0556694f $X=4.345 $Y=2.52 $X2=0
+ $Y2=0
cc_592 N_A_27_125#_c_843_n N_VPWR_c_1036_n 0.012253f $X=4.585 $Y=2.24 $X2=0
+ $Y2=0
cc_593 N_A_27_125#_c_840_n N_X_M1002_d 0.00396493f $X=4.345 $Y=2.52 $X2=0 $Y2=0
cc_594 N_A_27_125#_c_840_n N_X_c_1133_n 0.0126864f $X=4.345 $Y=2.52 $X2=0 $Y2=0
cc_595 N_A_27_125#_c_840_n A_817_419# 0.00320505f $X=4.345 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_596 N_A_27_125#_c_834_n N_VGND_c_1155_n 0.00660378f $X=4.43 $Y=2.075 $X2=0
+ $Y2=0
cc_597 N_A_27_125#_c_835_n N_VGND_c_1155_n 0.0122097f $X=4.625 $Y=0.73 $X2=0
+ $Y2=0
cc_598 N_A_27_125#_c_833_n N_VGND_c_1158_n 0.00482586f $X=0.26 $Y=0.835 $X2=0
+ $Y2=0
cc_599 N_A_27_125#_c_835_n N_VGND_c_1160_n 0.0094145f $X=4.625 $Y=0.73 $X2=0
+ $Y2=0
cc_600 N_A_27_125#_c_833_n N_VGND_c_1163_n 0.00851678f $X=0.26 $Y=0.835 $X2=0
+ $Y2=0
cc_601 N_A_27_125#_c_835_n N_VGND_c_1163_n 0.0116781f $X=4.625 $Y=0.73 $X2=0
+ $Y2=0
cc_602 N_A_196_125#_c_936_n N_VPWR_M1025_d 0.0209789f $X=6.335 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_603 N_A_196_125#_c_936_n N_VPWR_M1019_s 0.00431059f $X=6.335 $Y=2.405 $X2=0
+ $Y2=0
cc_604 N_A_196_125#_c_936_n N_VPWR_c_1037_n 0.00206261f $X=6.335 $Y=2.405 $X2=0
+ $Y2=0
cc_605 N_A_196_125#_c_936_n N_VPWR_c_1038_n 0.00206261f $X=6.335 $Y=2.405 $X2=0
+ $Y2=0
cc_606 N_A_196_125#_c_936_n N_VPWR_c_1039_n 0.0562588f $X=6.335 $Y=2.405 $X2=0
+ $Y2=0
cc_607 N_A_196_125#_c_982_n N_VPWR_c_1039_n 0.00201059f $X=6.48 $Y=2.405 $X2=0
+ $Y2=0
cc_608 N_A_196_125#_c_939_n N_VPWR_c_1039_n 0.014095f $X=6.665 $Y=2.24 $X2=0
+ $Y2=0
cc_609 N_A_196_125#_c_939_n N_VPWR_c_1040_n 0.00299218f $X=6.665 $Y=2.24 $X2=0
+ $Y2=0
cc_610 N_A_196_125#_c_939_n N_VPWR_c_1041_n 0.00833954f $X=6.665 $Y=2.24 $X2=0
+ $Y2=0
cc_611 N_A_196_125#_c_939_n N_VPWR_c_1042_n 0.0107659f $X=6.665 $Y=2.24 $X2=0
+ $Y2=0
cc_612 N_A_196_125#_c_939_n N_VPWR_c_1036_n 0.0133987f $X=6.665 $Y=2.24 $X2=0
+ $Y2=0
cc_613 N_A_196_125#_c_936_n N_X_M1002_d 0.00363609f $X=6.335 $Y=2.405 $X2=0
+ $Y2=0
cc_614 N_A_196_125#_c_936_n N_X_c_1133_n 0.00670125f $X=6.335 $Y=2.405 $X2=0
+ $Y2=0
cc_615 N_A_196_125#_c_936_n A_817_419# 0.00555716f $X=6.335 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_616 N_A_196_125#_c_936_n A_975_419# 0.00787256f $X=6.335 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_617 N_A_196_125#_c_936_n A_1223_419# 0.0103312f $X=6.335 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_618 N_X_c_1133_n N_VGND_c_1159_n 0.0138717f $X=3.16 $Y=0.42 $X2=0 $Y2=0
cc_619 N_X_M1015_d N_VGND_c_1163_n 0.00397496f $X=3.02 $Y=0.235 $X2=0 $Y2=0
cc_620 N_X_c_1133_n N_VGND_c_1163_n 0.00886411f $X=3.16 $Y=0.42 $X2=0 $Y2=0
