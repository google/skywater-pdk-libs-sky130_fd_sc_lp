* File: sky130_fd_sc_lp__o21ba_m.pex.spice
* Created: Wed Sep  2 10:17:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BA_M%A_88_41# 1 2 9 11 16 19 22 23 28
c60 23 0 1.8319e-19 $X=2.29 $Y=0.39
r61 25 28 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=2.29 $Y=2.82 $X2=2.37
+ $Y2=2.82
r62 21 23 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=2.21 $Y=0.39 $X2=2.29
+ $Y2=0.39
r63 21 22 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0.39
+ $X2=2.045 $Y2=0.39
r64 19 25 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.29 $Y=2.715
+ $X2=2.29 $Y2=2.82
r65 18 23 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.29 $Y=0.495
+ $X2=2.29 $Y2=0.39
r66 18 19 144.834 $w=1.68e-07 $l=2.22e-06 $layer=LI1_cond $X=2.29 $Y=0.495
+ $X2=2.29 $Y2=2.715
r67 16 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=0.37
+ $X2=0.605 $Y2=0.535
r68 15 22 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.605 $Y=0.37
+ $X2=2.045 $Y2=0.37
r69 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=0.37 $X2=0.605 $Y2=0.37
r70 9 11 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=0.68 $Y=1.025
+ $X2=0.68 $Y2=2.045
r71 9 32 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.68 $Y=1.025
+ $X2=0.68 $Y2=0.535
r72 2 28 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.23
+ $Y=2.675 $X2=2.37 $Y2=2.82
r73 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.245 $X2=2.21 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_M%B1_N 3 6 8 9 13 15
c36 9 0 1.49404e-20 $X=1.2 $Y=1.665
r37 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.51
+ $X2=1.13 $Y2=1.675
r38 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.51
+ $X2=1.13 $Y2=1.345
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.51 $X2=1.13 $Y2=1.51
r40 9 14 2.48218 $w=3.23e-07 $l=7e-08 $layer=LI1_cond $X=1.2 $Y=1.587 $X2=1.13
+ $Y2=1.587
r41 8 14 14.5385 $w=3.23e-07 $l=4.1e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=1.13 $Y2=1.587
r42 6 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.205 $Y=2.465
+ $X2=1.205 $Y2=1.675
r43 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.205 $Y=0.815
+ $X2=1.205 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_M%A_256_79# 1 2 9 11 13 17 20 21 23 27 29 33
+ 34 39
c59 20 0 1.49404e-20 $X=2.002 $Y=1.445
r60 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.94
+ $Y=0.94 $X2=1.94 $Y2=0.94
r61 31 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.94 $Y=1.275
+ $X2=1.94 $Y2=0.94
r62 30 37 23.1838 $w=3.21e-07 $l=7.0075e-07 $layer=LI1_cond $X=1.645 $Y=1.36
+ $X2=1.45 $Y2=0.75
r63 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.855 $Y=1.36
+ $X2=1.94 $Y2=1.275
r64 29 30 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.855 $Y=1.36
+ $X2=1.645 $Y2=1.36
r65 27 30 5.9155 $w=3.21e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.56 $Y=1.445
+ $X2=1.645 $Y2=1.36
r66 27 39 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.56 $Y=1.445
+ $X2=1.56 $Y2=1.93
r67 23 25 25.2794 $w=3.08e-07 $l=6.8e-07 $layer=LI1_cond $X=1.49 $Y=2.095
+ $X2=1.49 $Y2=2.775
r68 21 39 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.49 $Y=2.085
+ $X2=1.49 $Y2=1.93
r69 21 23 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=1.49 $Y=2.085
+ $X2=1.49 $Y2=2.095
r70 19 34 33.9804 $w=4.55e-07 $l=2.78e-07 $layer=POLY_cond $X=2.002 $Y=1.218
+ $X2=2.002 $Y2=0.94
r71 19 20 54.6551 $w=4.55e-07 $l=2.27e-07 $layer=POLY_cond $X=2.002 $Y=1.218
+ $X2=2.002 $Y2=1.445
r72 15 34 1.83347 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=2.002 $Y=0.925
+ $X2=2.002 $Y2=0.94
r73 15 17 216.9 $w=1.5e-07 $l=4.23e-07 $layer=POLY_cond $X=2.002 $Y=0.85
+ $X2=2.425 $Y2=0.85
r74 11 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.425 $Y=0.775
+ $X2=2.425 $Y2=0.85
r75 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.425 $Y=0.775
+ $X2=2.425 $Y2=0.455
r76 9 20 738.383 $w=1.5e-07 $l=1.44e-06 $layer=POLY_cond $X=2.155 $Y=2.885
+ $X2=2.155 $Y2=1.445
r77 2 25 400 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=1.28
+ $Y=1.835 $X2=1.42 $Y2=2.775
r78 2 23 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=1.28
+ $Y=1.835 $X2=1.42 $Y2=2.095
r79 1 37 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=1.28
+ $Y=0.395 $X2=1.42 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_M%A2 2 5 9 11 12 13 14 15 21
c41 9 0 1.8319e-19 $X=2.855 $Y=0.455
r42 21 23 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.72 $Y=1.375
+ $X2=2.72 $Y2=1.21
r43 14 15 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.657 $Y=2.035
+ $X2=2.657 $Y2=2.405
r44 13 14 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.657 $Y=1.665
+ $X2=2.657 $Y2=2.035
r45 12 13 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.657 $Y=1.295
+ $X2=2.657 $Y2=1.665
r46 12 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.675
+ $Y=1.375 $X2=2.675 $Y2=1.375
r47 9 23 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.855 $Y=0.455
+ $X2=2.855 $Y2=1.21
r48 5 11 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=2.585 $Y=2.885
+ $X2=2.585 $Y2=1.88
r49 2 11 52.1105 $w=4.2e-07 $l=2.1e-07 $layer=POLY_cond $X=2.72 $Y=1.67 $X2=2.72
+ $Y2=1.88
r50 1 21 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=2.72 $Y=1.42 $X2=2.72
+ $Y2=1.375
r51 1 2 33.1044 $w=4.2e-07 $l=2.5e-07 $layer=POLY_cond $X=2.72 $Y=1.42 $X2=2.72
+ $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_M%A1 3 7 12 16 17 18 19 25
r31 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.335
+ $Y=1.765 $X2=3.335 $Y2=1.765
r32 18 19 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.227 $Y=2.035
+ $X2=3.227 $Y2=2.405
r33 18 26 8.08207 $w=3.83e-07 $l=2.7e-07 $layer=LI1_cond $X=3.227 $Y=2.035
+ $X2=3.227 $Y2=1.765
r34 17 26 2.99336 $w=3.83e-07 $l=1e-07 $layer=LI1_cond $X=3.227 $Y=1.665
+ $X2=3.227 $Y2=1.765
r35 16 17 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.227 $Y=1.295
+ $X2=3.227 $Y2=1.665
r36 15 25 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.335 $Y=1.6
+ $X2=3.335 $Y2=1.765
r37 12 25 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=3.335 $Y=2.12
+ $X2=3.335 $Y2=1.765
r38 9 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.945 $Y=2.195
+ $X2=3.335 $Y2=2.195
r39 7 15 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=3.285 $Y=0.455
+ $X2=3.285 $Y2=1.6
r40 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.945 $Y=2.27
+ $X2=2.945 $Y2=2.195
r41 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.945 $Y=2.27
+ $X2=2.945 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_M%X 1 2 7 9 12 13 14 15 32
r20 32 33 5.96742 $w=4.73e-07 $l=3e-08 $layer=LI1_cond $X=0.392 $Y=2.035
+ $X2=0.392 $Y2=2.005
r21 25 36 3.32384 $w=4.73e-07 $l=1.32e-07 $layer=LI1_cond $X=0.392 $Y=2.242
+ $X2=0.392 $Y2=2.11
r22 14 15 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.392 $Y=2.405
+ $X2=0.392 $Y2=2.775
r23 14 25 4.10444 $w=4.73e-07 $l=1.63e-07 $layer=LI1_cond $X=0.392 $Y=2.405
+ $X2=0.392 $Y2=2.242
r24 13 36 1.20867 $w=4.73e-07 $l=4.8e-08 $layer=LI1_cond $X=0.392 $Y=2.062
+ $X2=0.392 $Y2=2.11
r25 13 32 0.679876 $w=4.73e-07 $l=2.7e-08 $layer=LI1_cond $X=0.392 $Y=2.062
+ $X2=0.392 $Y2=2.035
r26 13 33 1.82674 $w=1.68e-07 $l=2.8e-08 $layer=LI1_cond $X=0.24 $Y=1.977
+ $X2=0.24 $Y2=2.005
r27 12 13 20.3551 $w=1.68e-07 $l=3.12e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.977
r28 11 12 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=0.24 $Y=1.195
+ $X2=0.24 $Y2=1.665
r29 7 11 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.325 $Y=1.09
+ $X2=0.24 $Y2=1.195
r30 7 9 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=0.325 $Y=1.09
+ $X2=0.465 $Y2=1.09
r31 2 36 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.34
+ $Y=1.835 $X2=0.465 $Y2=2.11
r32 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.34
+ $Y=0.815 $X2=0.465 $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_M%VPWR 1 2 3 12 18 22 25 26 28 29 30 39 45 46
+ 49
r44 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 46 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r47 43 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.16 $Y2=3.33
r48 43 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 42 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 39 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.16 $Y2=3.33
r52 39 41 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 34 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 30 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 30 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 28 37 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 28 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.93 $Y2=3.33
r60 27 41 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 27 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.93 $Y2=3.33
r62 25 33 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 25 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.99 $Y2=3.33
r64 24 37 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 24 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.99 $Y2=3.33
r66 20 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=3.245
+ $X2=3.16 $Y2=3.33
r67 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.16 $Y=3.245
+ $X2=3.16 $Y2=2.95
r68 16 29 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r69 16 18 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.95
r70 12 15 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=0.99 $Y=2.27
+ $X2=0.99 $Y2=2.95
r71 10 26 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=3.245
+ $X2=0.99 $Y2=3.33
r72 10 15 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.99 $Y=3.245
+ $X2=0.99 $Y2=2.95
r73 3 22 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=2.675 $X2=3.16 $Y2=2.95
r74 2 18 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.815
+ $Y=2.675 $X2=1.94 $Y2=2.95
r75 1 15 400 $w=1.7e-07 $l=1.22689e-06 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=1.835 $X2=0.99 $Y2=2.95
r76 1 12 400 $w=1.7e-07 $l=5.39861e-07 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=1.835 $X2=0.99 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_M%VGND 1 2 7 8 9 10 13 17 20 21 22 29 30
c52 13 0 7.45681e-20 $X=0.915 $Y=0.96
r53 33 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r54 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 27 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r56 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r57 24 33 3.40825 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=0 $X2=0.13
+ $Y2=0
r58 24 26 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=0 $X2=2.64
+ $Y2=0
r59 22 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r60 22 34 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.24
+ $Y2=0
r61 20 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.64
+ $Y2=0
r62 20 21 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=3.07
+ $Y2=0
r63 19 29 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.6
+ $Y2=0
r64 19 21 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.07
+ $Y2=0
r65 15 21 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0
r66 15 17 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0.39
r67 11 13 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=0.915 $Y=0.805
+ $X2=0.915 $Y2=0.96
r68 9 11 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.81 $Y=0.72
+ $X2=0.915 $Y2=0.805
r69 9 10 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.81 $Y=0.72 $X2=0.26
+ $Y2=0.72
r70 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.175 $Y=0.635
+ $X2=0.26 $Y2=0.72
r71 7 33 3.40825 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.175 $Y=0.085
+ $X2=0.13 $Y2=0
r72 7 8 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.175 $Y=0.085
+ $X2=0.175 $Y2=0.635
r73 2 17 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.245 $X2=3.07 $Y2=0.39
r74 1 13 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.755
+ $Y=0.815 $X2=0.915 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_M%A_500_49# 1 2 9 11 12 15
r28 13 15 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=3.5 $Y=0.735 $X2=3.5
+ $Y2=0.52
r29 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.395 $Y=0.82
+ $X2=3.5 $Y2=0.735
r30 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.395 $Y=0.82
+ $X2=2.745 $Y2=0.82
r31 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.65 $Y=0.735
+ $X2=2.745 $Y2=0.82
r32 7 9 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=2.65 $Y=0.735
+ $X2=2.65 $Y2=0.52
r33 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.36
+ $Y=0.245 $X2=3.5 $Y2=0.52
r34 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.245 $X2=2.64 $Y2=0.52
.ends

