* File: sky130_fd_sc_lp__o221a_4.pex.spice
* Created: Wed Sep  2 10:18:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221A_4%C1 1 3 6 8 10 13 15 16 24
r43 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.485 $Y=1.44
+ $X2=0.915 $Y2=1.44
r44 20 23 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.27 $Y=1.44
+ $X2=0.485 $Y2=1.44
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.44 $X2=0.27 $Y2=1.44
r46 16 21 8.34346 $w=3.29e-07 $l=2.25e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=1.44
r47 15 21 5.3769 $w=3.29e-07 $l=1.45e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.44
r48 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.605
+ $X2=0.915 $Y2=1.44
r49 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.915 $Y=1.605
+ $X2=0.915 $Y2=2.465
r50 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.275
+ $X2=0.915 $Y2=1.44
r51 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.915 $Y=1.275
+ $X2=0.915 $Y2=0.745
r52 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.605
+ $X2=0.485 $Y2=1.44
r53 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.485 $Y=1.605
+ $X2=0.485 $Y2=2.465
r54 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.275
+ $X2=0.485 $Y2=1.44
r55 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.485 $Y=1.275
+ $X2=0.485 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%B1 3 6 8 10 13 15 19 20 22 23 28 30 45
c88 30 0 4.64396e-20 $X=1.365 $Y=1.275
c89 28 0 9.51233e-20 $X=1.365 $Y=1.44
c90 19 0 8.30442e-20 $X=2.99 $Y=1.44
r91 28 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.44
+ $X2=1.365 $Y2=1.605
r92 28 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.44
+ $X2=1.365 $Y2=1.275
r93 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.365
+ $Y=1.44 $X2=1.365 $Y2=1.44
r94 23 45 9.14018 $w=5.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.68 $Y=1.34
+ $X2=1.82 $Y2=1.34
r95 23 29 5.96507 $w=5.63e-07 $l=2.3e-07 $layer=LI1_cond $X=1.595 $Y=1.407
+ $X2=1.365 $Y2=1.407
r96 22 29 4.814 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=1.407
+ $X2=1.365 $Y2=1.407
r97 20 32 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=2.99 $Y=1.44
+ $X2=2.675 $Y2=1.44
r98 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.44 $X2=2.99 $Y2=1.44
r99 17 19 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=3.03 $Y=1.245
+ $X2=3.03 $Y2=1.44
r100 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.905 $Y=1.16
+ $X2=3.03 $Y2=1.245
r101 15 45 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=2.905 $Y=1.16
+ $X2=1.82 $Y2=1.16
r102 11 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.605
+ $X2=2.675 $Y2=1.44
r103 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.675 $Y=1.605
+ $X2=2.675 $Y2=2.465
r104 8 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.275
+ $X2=2.675 $Y2=1.44
r105 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.675 $Y=1.275
+ $X2=2.675 $Y2=0.745
r106 6 31 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.385 $Y=2.465
+ $X2=1.385 $Y2=1.605
r107 3 30 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.345 $Y=0.745
+ $X2=1.345 $Y2=1.275
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%B2 3 7 11 15 17 18 26
c50 26 0 8.30442e-20 $X=2.245 $Y=1.51
c51 18 0 9.51233e-20 $X=2.64 $Y=1.665
c52 11 0 6.83896e-20 $X=2.245 $Y=0.745
r53 24 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.155 $Y=1.51
+ $X2=2.245 $Y2=1.51
r54 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.155
+ $Y=1.51 $X2=2.155 $Y2=1.51
r55 21 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.815 $Y=1.51
+ $X2=2.155 $Y2=1.51
r56 17 18 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=2.64 $Y2=1.592
r57 17 25 0.172006 $w=3.33e-07 $l=5e-09 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=2.155 $Y2=1.592
r58 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.245 $Y=1.675
+ $X2=2.245 $Y2=1.51
r59 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.245 $Y=1.675
+ $X2=2.245 $Y2=2.465
r60 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.245 $Y=1.345
+ $X2=2.245 $Y2=1.51
r61 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.245 $Y=1.345 $X2=2.245
+ $Y2=0.745
r62 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.675
+ $X2=1.815 $Y2=1.51
r63 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.815 $Y=1.675
+ $X2=1.815 $Y2=2.465
r64 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.345
+ $X2=1.815 $Y2=1.51
r65 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.815 $Y=1.345 $X2=1.815
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%A1 3 7 10 14 17 21 23 26 29 30 31 34
c85 30 0 1.13212e-19 $X=4.935 $Y=1.35
r86 29 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.35
+ $X2=4.935 $Y2=1.515
r87 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.35
+ $X2=4.935 $Y2=1.185
r88 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.35 $X2=4.935 $Y2=1.35
r89 23 30 9.82196 $w=4.38e-07 $l=3.75e-07 $layer=LI1_cond $X=4.56 $Y=1.295
+ $X2=4.935 $Y2=1.295
r90 23 34 7.00188 $w=4.38e-07 $l=9.5e-08 $layer=LI1_cond $X=4.56 $Y=1.295
+ $X2=4.465 $Y2=1.295
r91 21 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.35
+ $X2=3.535 $Y2=1.515
r92 21 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.35
+ $X2=3.535 $Y2=1.185
r93 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.535
+ $Y=1.35 $X2=3.535 $Y2=1.35
r94 17 20 6.84263 $w=3.18e-07 $l=1.9e-07 $layer=LI1_cond $X=3.53 $Y=1.16
+ $X2=3.53 $Y2=1.35
r95 16 17 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.69 $Y=1.16 $X2=3.53
+ $Y2=1.16
r96 16 34 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.69 $Y=1.16
+ $X2=4.465 $Y2=1.16
r97 14 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.915 $Y=0.655
+ $X2=4.915 $Y2=1.185
r98 10 32 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.845 $Y=2.465
+ $X2=4.845 $Y2=1.515
r99 7 26 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.625 $Y=0.655
+ $X2=3.625 $Y2=1.185
r100 3 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.555 $Y=2.465
+ $X2=3.555 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%A2 3 7 11 15 17 23 24
r53 24 25 11.4373 $w=2.95e-07 $l=7e-08 $layer=POLY_cond $X=4.415 $Y=1.51
+ $X2=4.485 $Y2=1.51
r54 22 24 46.5661 $w=2.95e-07 $l=2.85e-07 $layer=POLY_cond $X=4.13 $Y=1.51
+ $X2=4.415 $Y2=1.51
r55 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.13
+ $Y=1.51 $X2=4.13 $Y2=1.51
r56 20 22 12.2542 $w=2.95e-07 $l=7.5e-08 $layer=POLY_cond $X=4.055 $Y=1.51
+ $X2=4.13 $Y2=1.51
r57 19 20 11.4373 $w=2.95e-07 $l=7e-08 $layer=POLY_cond $X=3.985 $Y=1.51
+ $X2=4.055 $Y2=1.51
r58 17 23 4.10641 $w=4.33e-07 $l=1.55e-07 $layer=LI1_cond $X=4.077 $Y=1.665
+ $X2=4.077 $Y2=1.51
r59 13 25 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.485 $Y=1.345
+ $X2=4.485 $Y2=1.51
r60 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.485 $Y=1.345
+ $X2=4.485 $Y2=0.655
r61 9 24 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.675
+ $X2=4.415 $Y2=1.51
r62 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.415 $Y=1.675
+ $X2=4.415 $Y2=2.465
r63 5 20 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.055 $Y=1.345
+ $X2=4.055 $Y2=1.51
r64 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.055 $Y=1.345
+ $X2=4.055 $Y2=0.655
r65 1 19 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.675
+ $X2=3.985 $Y2=1.51
r66 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.985 $Y=1.675
+ $X2=3.985 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%A_112_65# 1 2 3 4 15 19 23 27 31 35 39 43 47
+ 50 53 55 59 63 66 67 72 75 77 79 81 90
c155 90 0 1.13212e-19 $X=6.675 $Y=1.49
c156 50 0 4.64396e-20 $X=0.735 $Y=1.93
r157 90 91 5.19077 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=6.675 $Y=1.49
+ $X2=6.71 $Y2=1.49
r158 87 88 5.19077 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=6.245 $Y=1.49
+ $X2=6.28 $Y2=1.49
r159 86 87 58.5815 $w=3.25e-07 $l=3.95e-07 $layer=POLY_cond $X=5.85 $Y=1.49
+ $X2=6.245 $Y2=1.49
r160 85 86 5.19077 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=5.815 $Y=1.49
+ $X2=5.85 $Y2=1.49
r161 82 83 5.19077 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=5.385 $Y=1.49
+ $X2=5.42 $Y2=1.49
r162 73 90 21.5046 $w=3.25e-07 $l=1.45e-07 $layer=POLY_cond $X=6.53 $Y=1.49
+ $X2=6.675 $Y2=1.49
r163 73 88 37.0769 $w=3.25e-07 $l=2.5e-07 $layer=POLY_cond $X=6.53 $Y=1.49
+ $X2=6.28 $Y2=1.49
r164 72 73 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.53
+ $Y=1.49 $X2=6.53 $Y2=1.49
r165 70 85 45.2338 $w=3.25e-07 $l=3.05e-07 $layer=POLY_cond $X=5.51 $Y=1.49
+ $X2=5.815 $Y2=1.49
r166 70 83 13.3477 $w=3.25e-07 $l=9e-08 $layer=POLY_cond $X=5.51 $Y=1.49
+ $X2=5.42 $Y2=1.49
r167 69 72 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=5.51 $Y=1.485
+ $X2=6.53 $Y2=1.485
r168 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.51
+ $Y=1.49 $X2=5.51 $Y2=1.49
r169 67 69 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=5.37 $Y=1.485
+ $X2=5.51 $Y2=1.485
r170 65 67 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.285 $Y=1.585
+ $X2=5.37 $Y2=1.485
r171 65 66 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.285 $Y=1.585
+ $X2=5.285 $Y2=1.93
r172 64 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=2.015
+ $X2=4.2 $Y2=2.015
r173 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.2 $Y=2.015
+ $X2=5.285 $Y2=1.93
r174 63 64 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=5.2 $Y=2.015
+ $X2=4.365 $Y2=2.015
r175 60 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.015
+ $X2=2.03 $Y2=2.015
r176 59 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=2.015
+ $X2=4.2 $Y2=2.015
r177 59 60 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.035 $Y=2.015
+ $X2=2.195 $Y2=2.015
r178 56 77 2.53056 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.865 $Y=2.015
+ $X2=0.735 $Y2=2.015
r179 55 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=2.015
+ $X2=2.03 $Y2=2.015
r180 55 56 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=1.865 $Y=2.015
+ $X2=0.865 $Y2=2.015
r181 51 77 3.91525 $w=2.35e-07 $l=9.66954e-08 $layer=LI1_cond $X=0.71 $Y=2.1
+ $X2=0.735 $Y2=2.015
r182 51 53 19.8052 $w=2.08e-07 $l=3.75e-07 $layer=LI1_cond $X=0.71 $Y=2.1
+ $X2=0.71 $Y2=2.475
r183 50 77 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=1.93
+ $X2=0.735 $Y2=2.015
r184 50 75 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=0.735 $Y=1.93
+ $X2=0.735 $Y2=1.145
r185 45 75 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.7 $Y=0.98
+ $X2=0.7 $Y2=1.145
r186 45 47 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.7 $Y=0.98 $X2=0.7
+ $Y2=0.68
r187 41 91 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.71 $Y=1.655
+ $X2=6.71 $Y2=1.49
r188 41 43 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.71 $Y=1.655
+ $X2=6.71 $Y2=2.465
r189 37 90 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.675 $Y=1.325
+ $X2=6.675 $Y2=1.49
r190 37 39 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.675 $Y=1.325
+ $X2=6.675 $Y2=0.655
r191 33 88 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.28 $Y=1.655
+ $X2=6.28 $Y2=1.49
r192 33 35 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.28 $Y=1.655
+ $X2=6.28 $Y2=2.465
r193 29 87 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.325
+ $X2=6.245 $Y2=1.49
r194 29 31 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.245 $Y=1.325
+ $X2=6.245 $Y2=0.655
r195 25 86 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.85 $Y=1.655
+ $X2=5.85 $Y2=1.49
r196 25 27 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.85 $Y=1.655
+ $X2=5.85 $Y2=2.465
r197 21 85 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.325
+ $X2=5.815 $Y2=1.49
r198 21 23 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.815 $Y=1.325
+ $X2=5.815 $Y2=0.655
r199 17 83 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.42 $Y=1.655
+ $X2=5.42 $Y2=1.49
r200 17 19 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.42 $Y=1.655
+ $X2=5.42 $Y2=2.465
r201 13 82 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.325
+ $X2=5.385 $Y2=1.49
r202 13 15 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.385 $Y=1.325
+ $X2=5.385 $Y2=0.655
r203 4 81 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=4.06
+ $Y=1.835 $X2=4.2 $Y2=2.095
r204 3 79 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=1.89
+ $Y=1.835 $X2=2.03 $Y2=2.095
r205 2 77 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=1.98
r206 2 53 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=2.475
r207 1 47 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.325 $X2=0.7 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 39 43 45 49
+ 51 56 64 69 74 83 86 89 92 96
r101 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r102 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r103 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r104 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r105 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r106 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r107 78 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r108 78 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r109 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 75 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=3.33
+ $X2=6.065 $Y2=3.33
r111 75 77 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.23 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 74 95 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=6.76 $Y=3.33 $X2=6.98
+ $Y2=3.33
r113 74 77 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.76 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 73 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r115 73 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r116 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r117 70 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.135 $Y2=3.33
r118 70 72 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 69 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.9 $Y=3.33
+ $X2=6.065 $Y2=3.33
r120 69 72 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.9 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 65 86 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=3.505 $Y=3.33
+ $X2=3.115 $Y2=3.33
r122 65 67 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.505 $Y=3.33
+ $X2=3.6 $Y2=3.33
r123 64 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.97 $Y=3.33
+ $X2=5.135 $Y2=3.33
r124 64 67 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=4.97 $Y=3.33
+ $X2=3.6 $Y2=3.33
r125 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r127 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 60 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r130 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r131 57 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.15 $Y2=3.33
r132 57 59 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.68 $Y2=3.33
r133 56 86 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=3.115 $Y2=3.33
r134 56 62 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.64 $Y2=3.33
r135 55 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 55 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r137 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 52 80 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r139 52 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 51 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.15 $Y2=3.33
r141 51 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.72 $Y2=3.33
r142 49 90 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r143 49 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r144 49 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r145 45 48 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=6.925 $Y=2.19
+ $X2=6.925 $Y2=2.95
r146 43 95 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=6.925 $Y=3.245
+ $X2=6.98 $Y2=3.33
r147 43 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.925 $Y=3.245
+ $X2=6.925 $Y2=2.95
r148 39 42 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=6.065 $Y=2.19
+ $X2=6.065 $Y2=2.95
r149 37 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.065 $Y=3.245
+ $X2=6.065 $Y2=3.33
r150 37 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.065 $Y=3.245
+ $X2=6.065 $Y2=2.95
r151 33 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.135 $Y=3.245
+ $X2=5.135 $Y2=3.33
r152 33 35 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=5.135 $Y=3.245
+ $X2=5.135 $Y2=2.39
r153 29 86 3.08259 $w=7.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=3.245
+ $X2=3.115 $Y2=3.33
r154 29 31 13.1875 $w=7.78e-07 $l=8.6e-07 $layer=LI1_cond $X=3.115 $Y=3.245
+ $X2=3.115 $Y2=2.385
r155 25 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=3.33
r156 25 27 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=2.385
r157 21 24 31.7795 $w=3.28e-07 $l=9.1e-07 $layer=LI1_cond $X=0.27 $Y=2.04
+ $X2=0.27 $Y2=2.95
r158 19 80 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r159 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.95
r160 6 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.835 $X2=6.925 $Y2=2.95
r161 6 45 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.835 $X2=6.925 $Y2=2.19
r162 5 42 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.925
+ $Y=1.835 $X2=6.065 $Y2=2.95
r163 5 39 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=5.925
+ $Y=1.835 $X2=6.065 $Y2=2.19
r164 4 35 300 $w=1.7e-07 $l=6.5372e-07 $layer=licon1_PDIFF $count=2 $X=4.92
+ $Y=1.835 $X2=5.135 $Y2=2.39
r165 3 31 150 $w=1.7e-07 $l=8.20122e-07 $layer=licon1_PDIFF $count=4 $X=2.75
+ $Y=1.835 $X2=3.34 $Y2=2.385
r166 2 27 300 $w=1.7e-07 $l=6.249e-07 $layer=licon1_PDIFF $count=2 $X=0.99
+ $Y=1.835 $X2=1.15 $Y2=2.385
r167 1 24 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.95
r168 1 21 400 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%A_292_367# 1 2 9 11 12 15
r14 13 15 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=2.46 $Y=2.905
+ $X2=2.46 $Y2=2.435
r15 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.365 $Y=2.99
+ $X2=2.46 $Y2=2.905
r16 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.365 $Y=2.99
+ $X2=1.695 $Y2=2.99
r17 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.59 $Y=2.905
+ $X2=1.695 $Y2=2.99
r18 7 9 24.8225 $w=2.08e-07 $l=4.7e-07 $layer=LI1_cond $X=1.59 $Y=2.905 $X2=1.59
+ $Y2=2.435
r19 2 15 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=2.32
+ $Y=1.835 $X2=2.46 $Y2=2.435
r20 1 9 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%A_726_367# 1 2 9 11 12 15
r16 13 15 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=4.665 $Y=2.905
+ $X2=4.665 $Y2=2.445
r17 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.535 $Y=2.99
+ $X2=4.665 $Y2=2.905
r18 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.535 $Y=2.99
+ $X2=3.865 $Y2=2.99
r19 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.77 $Y=2.905
+ $X2=3.865 $Y2=2.99
r20 7 9 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=3.77 $Y=2.905 $X2=3.77
+ $Y2=2.435
r21 2 15 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=4.49
+ $Y=1.835 $X2=4.63 $Y2=2.445
r22 1 9 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=1.835 $X2=3.77 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41
+ 42 44 45 49 51
r61 49 51 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=6.99 $Y=1.215 $X2=6.99
+ $Y2=1.295
r62 44 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=1.13 $X2=6.99
+ $Y2=1.215
r63 44 45 16.964 $w=2.48e-07 $l=3.68e-07 $layer=LI1_cond $X=6.99 $Y=1.297
+ $X2=6.99 $Y2=1.665
r64 44 51 0.0921954 $w=2.48e-07 $l=2e-09 $layer=LI1_cond $X=6.99 $Y=1.297
+ $X2=6.99 $Y2=1.295
r65 43 45 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=6.99 $Y=1.755 $X2=6.99
+ $Y2=1.665
r66 40 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.59 $Y=1.84
+ $X2=6.495 $Y2=1.84
r67 39 43 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.865 $Y=1.84
+ $X2=6.99 $Y2=1.755
r68 39 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.865 $Y=1.84
+ $X2=6.59 $Y2=1.84
r69 38 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.555 $Y=1.13
+ $X2=6.46 $Y2=1.13
r70 37 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.865 $Y=1.13
+ $X2=6.99 $Y2=1.13
r71 37 38 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.865 $Y=1.13
+ $X2=6.555 $Y2=1.13
r72 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.495 $Y=1.98
+ $X2=6.495 $Y2=2.91
r73 31 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.495 $Y=1.925
+ $X2=6.495 $Y2=1.84
r74 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.495 $Y=1.925
+ $X2=6.495 $Y2=1.98
r75 27 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=1.045
+ $X2=6.46 $Y2=1.13
r76 27 29 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=6.46 $Y=1.045
+ $X2=6.46 $Y2=0.42
r77 25 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.4 $Y=1.84 $X2=6.495
+ $Y2=1.84
r78 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.4 $Y=1.84 $X2=5.73
+ $Y2=1.84
r79 23 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.365 $Y=1.13
+ $X2=6.46 $Y2=1.13
r80 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.365 $Y=1.13
+ $X2=5.695 $Y2=1.13
r81 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=5.635 $Y=1.98
+ $X2=5.635 $Y2=2.91
r82 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.635 $Y=1.925
+ $X2=5.73 $Y2=1.84
r83 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=5.635 $Y=1.925
+ $X2=5.635 $Y2=1.98
r84 13 24 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.58 $Y=1.045
+ $X2=5.695 $Y2=1.13
r85 13 15 31.3164 $w=2.28e-07 $l=6.25e-07 $layer=LI1_cond $X=5.58 $Y=1.045
+ $X2=5.58 $Y2=0.42
r86 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.355
+ $Y=1.835 $X2=6.495 $Y2=2.91
r87 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.355
+ $Y=1.835 $X2=6.495 $Y2=1.98
r88 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.495
+ $Y=1.835 $X2=5.635 $Y2=2.91
r89 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.495
+ $Y=1.835 $X2=5.635 $Y2=1.98
r90 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.32
+ $Y=0.235 $X2=6.46 $Y2=0.42
r91 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.46
+ $Y=0.235 $X2=5.6 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%A_29_65# 1 2 3 4 15 17 18 26 28 29
c38 28 0 6.83896e-20 $X=2.89 $Y=0.47
r39 28 29 6.37863 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=0.405
+ $X2=2.725 $Y2=0.405
r40 24 29 28.1034 $w=2.83e-07 $l=6.95e-07 $layer=LI1_cond $X=2.03 $Y=0.397
+ $X2=2.725 $Y2=0.397
r41 22 26 5.21318 $w=2.27e-07 $l=1.15e-07 $layer=LI1_cond $X=1.265 $Y=0.397
+ $X2=1.15 $Y2=0.397
r42 22 24 30.934 $w=2.83e-07 $l=7.65e-07 $layer=LI1_cond $X=1.265 $Y=0.397
+ $X2=2.03 $Y2=0.397
r43 17 26 5.21318 $w=2.27e-07 $l=1.40641e-07 $layer=LI1_cond $X=1.035 $Y=0.34
+ $X2=1.15 $Y2=0.397
r44 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.035 $Y=0.34
+ $X2=0.365 $Y2=0.34
r45 13 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.235 $Y=0.425
+ $X2=0.365 $Y2=0.34
r46 13 15 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=0.235 $Y=0.425
+ $X2=0.235 $Y2=0.47
r47 4 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.75
+ $Y=0.325 $X2=2.89 $Y2=0.47
r48 3 24 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.325 $X2=2.03 $Y2=0.45
r49 2 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.99
+ $Y=0.325 $X2=1.13 $Y2=0.47
r50 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.325 $X2=0.27 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%A_284_65# 1 2 3 4 13 21 25 27 28
r44 27 28 30.1919 $w=1.78e-07 $l=4.9e-07 $layer=LI1_cond $X=2.645 $Y=0.815
+ $X2=3.135 $Y2=0.815
r45 23 25 48.9138 $w=1.93e-07 $l=8.6e-07 $layer=LI1_cond $X=3.84 $Y=0.807
+ $X2=4.7 $Y2=0.807
r46 21 28 5.60117 $w=1.93e-07 $l=9.7e-08 $layer=LI1_cond $X=3.232 $Y=0.807
+ $X2=3.135 $Y2=0.807
r47 21 23 34.5809 $w=1.93e-07 $l=6.08e-07 $layer=LI1_cond $X=3.232 $Y=0.807
+ $X2=3.84 $Y2=0.807
r48 15 18 48.9138 $w=1.93e-07 $l=8.6e-07 $layer=LI1_cond $X=1.6 $Y=0.807
+ $X2=2.46 $Y2=0.807
r49 13 27 5.60117 $w=1.93e-07 $l=9.7e-08 $layer=LI1_cond $X=2.548 $Y=0.807
+ $X2=2.645 $Y2=0.807
r50 13 18 5.00513 $w=1.93e-07 $l=8.8e-08 $layer=LI1_cond $X=2.548 $Y=0.807
+ $X2=2.46 $Y2=0.807
r51 4 25 182 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_NDIFF $count=1 $X=4.56
+ $Y=0.235 $X2=4.7 $Y2=0.805
r52 3 23 182 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_NDIFF $count=1 $X=3.7
+ $Y=0.235 $X2=3.84 $Y2=0.805
r53 2 18 182 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_NDIFF $count=1 $X=2.32
+ $Y=0.325 $X2=2.46 $Y2=0.805
r54 1 15 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=1.42
+ $Y=0.325 $X2=1.6 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_4%VGND 1 2 3 4 5 18 22 24 28 32 34 36 39 40 41
+ 42 43 55 60 66 69 73
r96 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r97 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r98 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r99 64 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r100 64 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r101 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r102 61 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6.03
+ $Y2=0
r103 61 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.195 $Y=0
+ $X2=6.48 $Y2=0
r104 60 72 4.67153 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=6.725 $Y=0
+ $X2=6.962 $Y2=0
r105 60 63 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.725 $Y=0 $X2=6.48
+ $Y2=0
r106 59 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r107 59 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r108 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r109 56 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.165
+ $Y2=0
r110 56 58 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.295 $Y=0
+ $X2=5.52 $Y2=0
r111 55 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=6.03
+ $Y2=0
r112 55 58 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=5.52
+ $Y2=0
r113 54 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r114 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r115 50 51 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r116 47 51 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=3.12 $Y2=0
r117 46 50 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.12
+ $Y2=0
r118 46 47 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r119 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r120 43 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r121 41 53 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.08
+ $Y2=0
r122 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.27
+ $Y2=0
r123 39 50 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.245 $Y=0
+ $X2=3.12 $Y2=0
r124 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.41
+ $Y2=0
r125 38 53 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.575 $Y=0
+ $X2=4.08 $Y2=0
r126 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=0 $X2=3.41
+ $Y2=0
r127 34 72 3.09464 $w=3.3e-07 $l=1.15521e-07 $layer=LI1_cond $X=6.89 $Y=0.085
+ $X2=6.962 $Y2=0
r128 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.89 $Y=0.085
+ $X2=6.89 $Y2=0.36
r129 30 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0
r130 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0.36
r131 26 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.085
+ $X2=5.165 $Y2=0
r132 26 28 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=5.165 $Y=0.085
+ $X2=5.165 $Y2=0.4
r133 25 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.27
+ $Y2=0
r134 24 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.165
+ $Y2=0
r135 24 25 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=4.435
+ $Y2=0
r136 20 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0
r137 20 22 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0.415
r138 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=0.085
+ $X2=3.41 $Y2=0
r139 16 18 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.41 $Y=0.085
+ $X2=3.41 $Y2=0.415
r140 5 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.75
+ $Y=0.235 $X2=6.89 $Y2=0.36
r141 4 32 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.89
+ $Y=0.235 $X2=6.03 $Y2=0.36
r142 3 28 91 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=2 $X=4.99
+ $Y=0.235 $X2=5.15 $Y2=0.4
r143 2 22 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.13
+ $Y=0.235 $X2=4.27 $Y2=0.415
r144 1 18 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.41 $Y2=0.415
.ends

