# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrtp_lp2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrtp_lp2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.195000 0.805000 1.865000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.005000 2.075000 7.565000 3.065000 ;
        RECT 7.315000 0.265000 7.565000 2.075000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.250000 1.225000 6.595000 1.895000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.495000 1.285000 1.825000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.680000 0.085000 ;
        RECT 0.935000  0.085000 1.265000 1.015000 ;
        RECT 2.835000  0.085000 3.165000 0.545000 ;
        RECT 5.050000  0.085000 5.380000 0.675000 ;
        RECT 6.445000  0.085000 6.775000 0.695000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.680000 3.415000 ;
        RECT 0.645000 2.785000 0.975000 3.245000 ;
        RECT 2.615000 2.665000 2.945000 3.245000 ;
        RECT 5.290000 2.075000 5.620000 3.245000 ;
        RECT 6.430000 2.075000 6.760000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.590000 0.445000 1.015000 ;
      RECT 0.090000 1.015000 0.260000 2.075000 ;
      RECT 0.090000 2.075000 0.445000 2.435000 ;
      RECT 0.090000 2.435000 1.985000 2.605000 ;
      RECT 0.090000 2.605000 0.445000 3.065000 ;
      RECT 1.255000 2.005000 1.635000 2.255000 ;
      RECT 1.465000 1.455000 2.540000 1.785000 ;
      RECT 1.465000 1.785000 1.635000 2.005000 ;
      RECT 1.805000 0.905000 2.135000 1.455000 ;
      RECT 1.815000 1.965000 3.040000 2.135000 ;
      RECT 1.815000 2.135000 1.985000 2.435000 ;
      RECT 2.045000 0.265000 2.485000 0.675000 ;
      RECT 2.165000 2.315000 3.985000 2.485000 ;
      RECT 2.165000 2.485000 2.415000 3.065000 ;
      RECT 2.315000 0.675000 2.485000 0.725000 ;
      RECT 2.315000 0.725000 3.860000 0.895000 ;
      RECT 2.370000 1.075000 3.390000 1.245000 ;
      RECT 2.370000 1.245000 2.540000 1.455000 ;
      RECT 2.750000 1.425000 3.040000 1.965000 ;
      RECT 3.220000 1.245000 3.390000 1.335000 ;
      RECT 3.220000 1.335000 4.170000 1.665000 ;
      RECT 3.570000 0.895000 3.860000 0.925000 ;
      RECT 3.570000 0.925000 4.520000 1.095000 ;
      RECT 3.795000 0.295000 4.870000 0.545000 ;
      RECT 3.815000 1.845000 4.760000 2.015000 ;
      RECT 3.815000 2.015000 3.985000 2.315000 ;
      RECT 4.165000 2.195000 5.110000 2.365000 ;
      RECT 4.165000 2.365000 4.495000 3.065000 ;
      RECT 4.350000 1.095000 4.520000 1.265000 ;
      RECT 4.350000 1.265000 4.760000 1.845000 ;
      RECT 4.700000 0.545000 4.870000 0.855000 ;
      RECT 4.700000 0.855000 5.110000 1.025000 ;
      RECT 4.940000 1.025000 5.110000 1.425000 ;
      RECT 4.940000 1.425000 5.720000 1.755000 ;
      RECT 4.940000 1.755000 5.110000 2.195000 ;
      RECT 5.290000 0.855000 6.070000 0.875000 ;
      RECT 5.290000 0.875000 7.105000 1.025000 ;
      RECT 5.290000 1.025000 5.620000 1.185000 ;
      RECT 5.625000 0.265000 6.070000 0.855000 ;
      RECT 5.900000 1.025000 7.105000 1.045000 ;
      RECT 5.900000 1.045000 6.070000 2.075000 ;
      RECT 5.900000 2.075000 6.230000 3.065000 ;
      RECT 6.775000 1.045000 7.105000 1.545000 ;
  END
END sky130_fd_sc_lp__dlrtp_lp2
