* NGSPICE file created from sky130_fd_sc_lp__a221o_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a221o_m A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_233_535# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.352e+11p ps=2.8e+06u
M1001 a_337_397# B2 a_233_535# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1002 VPWR a_33_153# X VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 VGND B2 a_399_47# VNB nshort w=420000u l=150000u
+  ad=3.003e+11p pd=3.11e+06u as=8.82e+10p ps=1.26e+06u
M1004 VGND a_33_153# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 a_399_47# B1 a_33_153# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.234e+11p ps=3.22e+06u
M1006 a_233_535# B1 a_337_397# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_196_47# A2 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 a_33_153# A1 a_196_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_33_153# C1 a_337_397# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1010 a_233_535# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_33_153# C1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

