* File: sky130_fd_sc_lp__and2b_1.pex.spice
* Created: Fri Aug 28 10:05:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2B_1%A_N 1 3 6 8 14
c32 14 0 2.84594e-19 $X=0.69 $Y=0.93
r33 12 14 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.635 $Y=0.93
+ $X2=0.69 $Y2=0.93
r34 10 12 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.475 $Y=0.93
+ $X2=0.635 $Y2=0.93
r35 8 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=0.93 $X2=0.69 $Y2=0.93
r36 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=1.095
+ $X2=0.635 $Y2=0.93
r37 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.635 $Y=1.095
+ $X2=0.635 $Y2=2.045
r38 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.765
+ $X2=0.475 $Y2=0.93
r39 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.765
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_1%A_27_47# 1 2 7 9 11 13 16 20 24 27
c48 24 0 1.68193e-19 $X=1.14 $Y=1.5
r49 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.5 $X2=1.14 $Y2=1.5
r50 22 27 1.73286 $w=3.3e-07 $l=2.23e-07 $layer=LI1_cond $X=0.54 $Y=1.5
+ $X2=0.317 $Y2=1.5
r51 22 24 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=0.54 $Y=1.5 $X2=1.14
+ $Y2=1.5
r52 18 27 4.71911 $w=3.67e-07 $l=1.65e-07 $layer=LI1_cond $X=0.317 $Y=1.665
+ $X2=0.317 $Y2=1.5
r53 18 20 9.84109 $w=4.43e-07 $l=3.8e-07 $layer=LI1_cond $X=0.317 $Y=1.665
+ $X2=0.317 $Y2=2.045
r54 14 27 4.71911 $w=3.67e-07 $l=1.99825e-07 $layer=LI1_cond $X=0.24 $Y=1.335
+ $X2=0.317 $Y2=1.5
r55 14 16 35.3681 $w=2.88e-07 $l=8.9e-07 $layer=LI1_cond $X=0.24 $Y=1.335
+ $X2=0.24 $Y2=0.445
r56 11 25 60.2754 $w=3.34e-07 $l=3.98052e-07 $layer=POLY_cond $X=1.425 $Y=1.185
+ $X2=1.237 $Y2=1.5
r57 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.425 $Y=1.185
+ $X2=1.425 $Y2=0.865
r58 7 25 38.6287 $w=3.34e-07 $l=1.68464e-07 $layer=POLY_cond $X=1.23 $Y=1.665
+ $X2=1.237 $Y2=1.5
r59 7 9 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.23 $Y=1.665 $X2=1.23
+ $Y2=2.045
r60 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.295
+ $Y=1.835 $X2=0.42 $Y2=2.045
r61 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_1%B 5 8 9 11 18
c32 5 0 1.68193e-19 $X=1.785 $Y=0.865
r33 18 20 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.687 $Y=2.58
+ $X2=1.687 $Y2=2.415
r34 11 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=2.58 $X2=1.68 $Y2=2.58
r35 9 11 7.60421 $w=7.53e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.697 $X2=1.68
+ $Y2=2.697
r36 8 20 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.785 $Y=2.045
+ $X2=1.785 $Y2=2.415
r37 5 8 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.785 $Y=0.865
+ $X2=1.785 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_1%A_217_131# 1 2 9 13 14 19 22 26 27 29 31
c57 19 0 7.4402e-20 $X=1.485 $Y=1.185
r58 27 32 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.257 $Y=1.35
+ $X2=2.257 $Y2=1.515
r59 27 31 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.257 $Y=1.35
+ $X2=2.257 $Y2=1.185
r60 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.35 $X2=2.235 $Y2=1.35
r61 24 29 0.225187 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.695 $Y=1.35
+ $X2=1.545 $Y2=1.35
r62 24 26 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=1.695 $Y=1.35
+ $X2=2.235 $Y2=1.35
r63 20 29 6.67463 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.515
+ $X2=1.545 $Y2=1.35
r64 20 22 18.0549 $w=2.98e-07 $l=4.7e-07 $layer=LI1_cond $X=1.545 $Y=1.515
+ $X2=1.545 $Y2=1.985
r65 19 29 6.67463 $w=2.4e-07 $l=1.92678e-07 $layer=LI1_cond $X=1.485 $Y=1.185
+ $X2=1.545 $Y2=1.35
r66 18 19 9.85859 $w=1.78e-07 $l=1.6e-07 $layer=LI1_cond $X=1.485 $Y=1.025
+ $X2=1.485 $Y2=1.185
r67 14 18 7.61292 $w=3.3e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.395 $Y=0.86
+ $X2=1.485 $Y2=1.025
r68 14 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.395 $Y=0.86
+ $X2=1.21 $Y2=0.86
r69 13 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.37 $Y=0.655
+ $X2=2.37 $Y2=1.185
r70 9 32 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.345 $Y=2.465
+ $X2=2.345 $Y2=1.515
r71 2 22 600 $w=1.7e-07 $l=2.90474e-07 $layer=licon1_PDIFF $count=1 $X=1.305
+ $Y=1.835 $X2=1.53 $Y2=1.985
r72 1 16 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.655 $X2=1.21 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_1%VPWR 1 2 10 14 18 23 25 27 34 35 38 41
r37 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 35 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 32 41 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.15 $Y2=3.33
r42 32 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 28 38 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.797 $Y2=3.33
r46 28 30 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 27 41 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.15 $Y2=3.33
r48 27 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 25 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 25 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 21 23 4.49004 $w=3.83e-07 $l=1.5e-07 $layer=LI1_cond $X=2 $Y=1.957 $X2=2.15
+ $Y2=1.957
r52 15 18 5.4741 $w=2.78e-07 $l=1.33e-07 $layer=LI1_cond $X=0.797 $Y=2.01
+ $X2=0.93 $Y2=2.01
r53 12 41 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r54 12 14 34.7867 $w=2.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.43
r55 11 23 2.81547 $w=2.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.15 $Y=2.15
+ $X2=2.15 $Y2=1.957
r56 11 14 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.15 $Y=2.15
+ $X2=2.15 $Y2=2.43
r57 10 38 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.797 $Y=3.245
+ $X2=0.797 $Y2=3.33
r58 9 15 3.50883 $w=1.75e-07 $l=1.4e-07 $layer=LI1_cond $X=0.797 $Y=2.15
+ $X2=0.797 $Y2=2.01
r59 9 10 69.3974 $w=1.73e-07 $l=1.095e-06 $layer=LI1_cond $X=0.797 $Y=2.15
+ $X2=0.797 $Y2=3.245
r60 2 21 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.835 $X2=2 $Y2=1.985
r61 2 14 300 $w=1.7e-07 $l=7.17409e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.835 $X2=2.13 $Y2=2.43
r62 1 18 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=1.835 $X2=0.93 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_1%X 1 2 7 8 9 10 11 12 13 24 34
r15 34 47 1.13355 $w=3.03e-07 $l=3e-08 $layer=LI1_cond $X=2.642 $Y=1.665
+ $X2=2.642 $Y2=1.695
r16 13 44 4.57588 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=2.625 $Y=2.775
+ $X2=2.625 $Y2=2.91
r17 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.625 $Y=2.405
+ $X2=2.625 $Y2=2.775
r18 11 12 14.4055 $w=3.38e-07 $l=4.25e-07 $layer=LI1_cond $X=2.625 $Y=1.98
+ $X2=2.625 $Y2=2.405
r19 11 35 3.89797 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=2.625 $Y=1.98
+ $X2=2.625 $Y2=1.865
r20 10 35 4.84704 $w=3.38e-07 $l=1.43e-07 $layer=LI1_cond $X=2.625 $Y=1.722
+ $X2=2.625 $Y2=1.865
r21 10 47 1.06308 $w=3.38e-07 $l=2.7e-08 $layer=LI1_cond $X=2.625 $Y=1.722
+ $X2=2.625 $Y2=1.695
r22 10 34 1.05798 $w=3.03e-07 $l=2.8e-08 $layer=LI1_cond $X=2.642 $Y=1.637
+ $X2=2.642 $Y2=1.665
r23 9 10 12.9225 $w=3.03e-07 $l=3.42e-07 $layer=LI1_cond $X=2.642 $Y=1.295
+ $X2=2.642 $Y2=1.637
r24 8 9 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.642 $Y=0.925
+ $X2=2.642 $Y2=1.295
r25 7 8 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.642 $Y=0.555
+ $X2=2.642 $Y2=0.925
r26 7 24 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.642 $Y=0.555
+ $X2=2.642 $Y2=0.42
r27 2 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.835 $X2=2.56 $Y2=2.91
r28 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.835 $X2=2.56 $Y2=1.98
r29 1 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.235 $X2=2.585 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_1%VGND 1 2 9 13 17 19 24 31 32 35 38
c35 32 0 1.28143e-19 $X=2.64 $Y=0
c36 19 0 8.20489e-20 $X=0.555 $Y=0
r37 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 29 38 11.0851 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.077
+ $Y2=0
r42 29 31 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.64
+ $Y2=0
r43 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r44 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 25 35 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.705
+ $Y2=0
r46 25 27 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.68
+ $Y2=0
r47 24 38 11.0851 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2.077
+ $Y2=0
r48 24 27 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.68
+ $Y2=0
r49 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r50 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 19 35 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.705
+ $Y2=0
r52 19 21 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.24
+ $Y2=0
r53 17 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r54 17 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r55 13 15 11.5909 $w=4.83e-07 $l=4.7e-07 $layer=LI1_cond $X=2.077 $Y=0.38
+ $X2=2.077 $Y2=0.85
r56 11 38 1.99554 $w=4.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.077 $Y=0.085
+ $X2=2.077 $Y2=0
r57 11 13 7.27512 $w=4.83e-07 $l=2.95e-07 $layer=LI1_cond $X=2.077 $Y=0.085
+ $X2=2.077 $Y2=0.38
r58 7 35 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r59 7 9 13.2531 $w=2.98e-07 $l=3.45e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.43
r60 2 15 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.655 $X2=2 $Y2=0.85
r61 2 13 182 $w=1.7e-07 $l=4.10061e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.655 $X2=2.155 $Y2=0.38
r62 1 9 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.43
.ends

