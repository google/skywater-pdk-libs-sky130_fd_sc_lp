* File: sky130_fd_sc_lp__or3b_4.spice
* Created: Fri Aug 28 11:24:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or3b_4.pex.spice"
.subckt sky130_fd_sc_lp__or3b_4  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_C_N_M1015_g N_A_49_133#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1218 AS=0.1113 PD=0.963333 PS=1.37 NRD=94.284 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.7 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1015_d N_A_253_23#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2436 AS=0.1176 PD=1.92667 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_253_23#_M1009_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001 SB=75002.5
+ A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1009_d N_A_253_23#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A_253_23#_M1012_g N_X_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1004 N_A_253_23#_M1004_d N_A_M1004_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=5.712 M=1 R=5.6 SA=75002.4
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_B_M1007_g N_A_253_23#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1617 AS=0.1176 PD=1.225 PS=1.12 NRD=7.848 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1006 N_A_253_23#_M1006_d N_A_49_133#_M1006_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1617 PD=2.21 PS=1.225 NRD=0 NRS=7.14 M=1 R=5.6
+ SA=75003.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1014 N_VPWR_M1014_d N_C_N_M1014_g N_A_49_133#_M1014_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.12285 AS=0.1113 PD=0.95 PS=1.37 NRD=111.384 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_253_23#_M1001_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.36855 PD=1.54 PS=2.85 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5 SB=75003
+ A=0.189 P=2.82 MULT=1
MM1002 N_X_M1001_d N_A_253_23#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1008 N_X_M1008_d N_A_253_23#_M1008_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.3
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1013 N_X_M1008_d N_A_253_23#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2457 PD=1.54 PS=1.65 NRD=0 NRS=8.5892 M=1 R=8.4 SA=75001.7
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1010 A_656_367# N_A_M1010_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.2457 PD=1.47 PS=1.65 NRD=7.8012 NRS=8.5892 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 A_728_367# N_B_M1005_g A_656_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75002.6
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1000 N_A_253_23#_M1000_d N_A_49_133#_M1000_g A_728_367# VPB PHIGHVT L=0.15
+ W=1.26 AD=0.378 AS=0.2457 PD=3.12 PS=1.65 NRD=2.6004 NRS=21.8867 M=1 R=8.4
+ SA=75003.2 SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__or3b_4.pxi.spice"
*
.ends
*
*
