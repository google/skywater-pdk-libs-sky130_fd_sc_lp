* File: sky130_fd_sc_lp__a31oi_4.pxi.spice
* Created: Fri Aug 28 10:00:13 2020
* 
x_PM_SKY130_FD_SC_LP__A31OI_4%A3 N_A3_M1011_g N_A3_M1010_g N_A3_M1023_g
+ N_A3_M1021_g N_A3_M1027_g N_A3_M1022_g N_A3_M1029_g N_A3_M1030_g A3 A3 A3 A3
+ A3 A3 N_A3_c_126_n PM_SKY130_FD_SC_LP__A31OI_4%A3
x_PM_SKY130_FD_SC_LP__A31OI_4%A2 N_A2_M1006_g N_A2_M1005_g N_A2_M1009_g
+ N_A2_M1007_g N_A2_M1019_g N_A2_M1020_g N_A2_c_206_n N_A2_c_207_n N_A2_M1028_g
+ N_A2_M1031_g A2 A2 A2 N_A2_c_209_n PM_SKY130_FD_SC_LP__A31OI_4%A2
x_PM_SKY130_FD_SC_LP__A31OI_4%A1 N_A1_M1000_g N_A1_M1001_g N_A1_M1008_g
+ N_A1_M1004_g N_A1_M1012_g N_A1_M1016_g N_A1_M1017_g N_A1_M1018_g A1 A1 A1 A1
+ N_A1_c_298_n PM_SKY130_FD_SC_LP__A31OI_4%A1
x_PM_SKY130_FD_SC_LP__A31OI_4%B1 N_B1_M1002_g N_B1_M1013_g N_B1_M1003_g
+ N_B1_M1015_g N_B1_M1014_g N_B1_M1024_g N_B1_M1026_g N_B1_M1025_g B1 B1 B1
+ N_B1_c_386_n PM_SKY130_FD_SC_LP__A31OI_4%B1
x_PM_SKY130_FD_SC_LP__A31OI_4%A_41_367# N_A_41_367#_M1010_d N_A_41_367#_M1021_d
+ N_A_41_367#_M1030_d N_A_41_367#_M1007_s N_A_41_367#_M1031_s
+ N_A_41_367#_M1008_d N_A_41_367#_M1017_d N_A_41_367#_M1003_s
+ N_A_41_367#_M1026_s N_A_41_367#_c_456_n N_A_41_367#_c_457_n
+ N_A_41_367#_c_462_n N_A_41_367#_c_508_p N_A_41_367#_c_466_n
+ N_A_41_367#_c_505_p N_A_41_367#_c_470_n N_A_41_367#_c_509_p
+ N_A_41_367#_c_477_n N_A_41_367#_c_481_n N_A_41_367#_c_506_p
+ N_A_41_367#_c_485_n N_A_41_367#_c_487_n N_A_41_367#_c_544_p
+ N_A_41_367#_c_489_n N_A_41_367#_c_512_p N_A_41_367#_c_547_p
+ N_A_41_367#_c_491_n N_A_41_367#_c_458_n N_A_41_367#_c_459_n
+ N_A_41_367#_c_471_n N_A_41_367#_c_473_n N_A_41_367#_c_482_n
+ N_A_41_367#_c_484_n N_A_41_367#_c_510_p N_A_41_367#_c_515_p
+ PM_SKY130_FD_SC_LP__A31OI_4%A_41_367#
x_PM_SKY130_FD_SC_LP__A31OI_4%VPWR N_VPWR_M1010_s N_VPWR_M1022_s N_VPWR_M1005_d
+ N_VPWR_M1019_d N_VPWR_M1000_s N_VPWR_M1012_s N_VPWR_c_557_n N_VPWR_c_558_n
+ N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n
+ N_VPWR_c_564_n N_VPWR_c_565_n VPWR N_VPWR_c_566_n N_VPWR_c_567_n
+ N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_556_n N_VPWR_c_572_n
+ N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_575_n PM_SKY130_FD_SC_LP__A31OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A31OI_4%Y N_Y_M1001_s N_Y_M1004_s N_Y_M1018_s N_Y_M1015_s
+ N_Y_M1025_s N_Y_M1002_d N_Y_M1014_d N_Y_c_680_n N_Y_c_702_n N_Y_c_681_n
+ N_Y_c_682_n N_Y_c_683_n N_Y_c_736_n N_Y_c_684_n N_Y_c_685_n N_Y_c_686_n
+ N_Y_c_687_n N_Y_c_688_n N_Y_c_720_n N_Y_c_689_n N_Y_c_753_n Y Y Y N_Y_c_690_n
+ Y PM_SKY130_FD_SC_LP__A31OI_4%Y
x_PM_SKY130_FD_SC_LP__A31OI_4%A_27_69# N_A_27_69#_M1011_s N_A_27_69#_M1023_s
+ N_A_27_69#_M1029_s N_A_27_69#_M1009_d N_A_27_69#_M1028_d N_A_27_69#_c_808_n
+ N_A_27_69#_c_809_n N_A_27_69#_c_810_n N_A_27_69#_c_811_n N_A_27_69#_c_812_n
+ N_A_27_69#_c_813_n N_A_27_69#_c_814_n N_A_27_69#_c_843_n N_A_27_69#_c_815_n
+ N_A_27_69#_c_816_n N_A_27_69#_c_817_n N_A_27_69#_c_818_n N_A_27_69#_c_819_n
+ PM_SKY130_FD_SC_LP__A31OI_4%A_27_69#
x_PM_SKY130_FD_SC_LP__A31OI_4%VGND N_VGND_M1011_d N_VGND_M1027_d N_VGND_M1013_d
+ N_VGND_M1024_d N_VGND_c_887_n N_VGND_c_888_n N_VGND_c_889_n N_VGND_c_890_n
+ N_VGND_c_891_n VGND N_VGND_c_892_n N_VGND_c_893_n N_VGND_c_894_n
+ N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n N_VGND_c_898_n N_VGND_c_899_n
+ N_VGND_c_900_n PM_SKY130_FD_SC_LP__A31OI_4%VGND
x_PM_SKY130_FD_SC_LP__A31OI_4%A_454_69# N_A_454_69#_M1006_s N_A_454_69#_M1020_s
+ N_A_454_69#_M1001_d N_A_454_69#_M1016_d N_A_454_69#_c_997_n
+ N_A_454_69#_c_990_n N_A_454_69#_c_991_n N_A_454_69#_c_1004_n
+ N_A_454_69#_c_992_n N_A_454_69#_c_993_n N_A_454_69#_c_1022_n
+ N_A_454_69#_c_994_n N_A_454_69#_c_995_n PM_SKY130_FD_SC_LP__A31OI_4%A_454_69#
cc_1 VNB N_A3_M1011_g 0.0251004f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_2 VNB N_A3_M1023_g 0.0183221f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.765
cc_3 VNB N_A3_M1027_g 0.0183221f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.765
cc_4 VNB N_A3_M1029_g 0.0186619f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.765
cc_5 VNB A3 0.0118785f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_6 VNB N_A3_c_126_n 0.0841744f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=1.51
cc_7 VNB N_A2_M1006_g 0.0188725f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_8 VNB N_A2_M1009_g 0.0190268f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.765
cc_9 VNB N_A2_M1020_g 0.0199064f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_10 VNB N_A2_c_206_n 0.0159699f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.345
cc_11 VNB N_A2_c_207_n 0.047693f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.765
cc_12 VNB N_A2_M1028_g 0.0235315f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=1.675
cc_13 VNB N_A2_c_209_n 0.0396887f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.51
cc_14 VNB N_A1_M1001_g 0.0206035f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_15 VNB N_A1_M1004_g 0.0164242f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_16 VNB N_A1_M1016_g 0.0164463f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_17 VNB N_A1_M1018_g 0.0172741f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_18 VNB A1 0.00260148f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_19 VNB N_A1_c_298_n 0.0805982f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.51
cc_20 VNB N_B1_M1013_g 0.0194035f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_21 VNB N_B1_M1015_g 0.0190876f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_22 VNB N_B1_M1024_g 0.0190876f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_23 VNB N_B1_M1025_g 0.0259913f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_24 VNB B1 0.0131297f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_25 VNB N_B1_c_386_n 0.0729673f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.51
cc_26 VNB N_VPWR_c_556_n 0.342803f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.592
cc_27 VNB N_Y_c_680_n 0.00502388f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_28 VNB N_Y_c_681_n 0.00255168f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.765
cc_29 VNB N_Y_c_682_n 0.00226963f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_30 VNB N_Y_c_683_n 0.00553405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_684_n 0.00214825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_685_n 0.0135249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_686_n 0.0310467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_687_n 0.00227951f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.51
cc_35 VNB N_Y_c_688_n 0.00180577f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.51
cc_36 VNB N_Y_c_689_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.51
cc_37 VNB N_Y_c_690_n 0.00100488f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.592
cc_38 VNB Y 0.00391895f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.592
cc_39 VNB N_A_27_69#_c_808_n 0.0307409f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.765
cc_40 VNB N_A_27_69#_c_809_n 0.0029562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_69#_c_810_n 0.011153f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.675
cc_42 VNB N_A_27_69#_c_811_n 0.00189238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_69#_c_812_n 0.00289786f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.765
cc_44 VNB N_A_27_69#_c_813_n 0.00189149f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_45 VNB N_A_27_69#_c_814_n 0.00335977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_69#_c_815_n 0.00699647f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_47 VNB N_A_27_69#_c_816_n 0.00627741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_69#_c_817_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_69#_c_818_n 0.00169851f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_50 VNB N_A_27_69#_c_819_n 0.00306307f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_51 VNB N_VGND_c_887_n 0.00270988f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_52 VNB N_VGND_c_888_n 0.00270988f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.765
cc_53 VNB N_VGND_c_889_n 0.111453f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.675
cc_54 VNB N_VGND_c_890_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.345
cc_55 VNB N_VGND_c_891_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=1.675
cc_56 VNB N_VGND_c_892_n 0.0164926f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_57 VNB N_VGND_c_893_n 0.0146145f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_58 VNB N_VGND_c_894_n 0.0142255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_895_n 0.0162797f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.51
cc_60 VNB N_VGND_c_896_n 0.436458f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.51
cc_61 VNB N_VGND_c_897_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.51
cc_62 VNB N_VGND_c_898_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.51
cc_63 VNB N_VGND_c_899_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=1.51
cc_64 VNB N_VGND_c_900_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.51
cc_65 VNB N_A_454_69#_c_990_n 0.00294772f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.345
cc_66 VNB N_A_454_69#_c_991_n 0.00203727f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.765
cc_67 VNB N_A_454_69#_c_992_n 0.0169967f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_68 VNB N_A_454_69#_c_993_n 0.00489901f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.345
cc_69 VNB N_A_454_69#_c_994_n 0.00221189f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_70 VNB N_A_454_69#_c_995_n 0.0018161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VPB N_A3_M1010_g 0.0240279f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_72 VPB N_A3_M1021_g 0.0178551f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_73 VPB N_A3_M1022_g 0.0178551f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.465
cc_74 VPB N_A3_M1030_g 0.0180434f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_75 VPB A3 0.0204449f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.58
cc_76 VPB N_A3_c_126_n 0.0201339f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=1.51
cc_77 VPB N_A2_M1005_g 0.0180434f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_78 VPB N_A2_M1007_g 0.0181814f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_79 VPB N_A2_M1019_g 0.0233892f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.765
cc_80 VPB N_A2_c_206_n 0.00873122f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.345
cc_81 VPB N_A2_c_207_n 0.0079303f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.765
cc_82 VPB N_A2_M1031_g 0.0248575f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_83 VPB A2 0.00927925f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.58
cc_84 VPB N_A2_c_209_n 0.0119538f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.51
cc_85 VPB N_A1_M1000_g 0.0172416f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_86 VPB N_A1_M1008_g 0.0176746f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.765
cc_87 VPB N_A1_M1012_g 0.0176869f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.765
cc_88 VPB N_A1_M1017_g 0.0186962f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.765
cc_89 VPB A1 0.0113908f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_90 VPB N_A1_c_298_n 0.0166167f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.51
cc_91 VPB N_B1_M1002_g 0.0184399f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_92 VPB N_B1_M1003_g 0.0178244f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.765
cc_93 VPB N_B1_M1014_g 0.017462f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.765
cc_94 VPB N_B1_M1026_g 0.023196f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.765
cc_95 VPB B1 0.0176962f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_96 VPB N_B1_c_386_n 0.0165229f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.51
cc_97 VPB N_A_41_367#_c_456_n 0.0075508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_41_367#_c_457_n 0.0369431f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_99 VPB N_A_41_367#_c_458_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.592
cc_100 VPB N_A_41_367#_c_459_n 0.0361069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_557_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.405 $Y2=1.675
cc_102 VPB N_VPWR_c_558_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.345
cc_103 VPB N_VPWR_c_559_n 3.08929e-19 $X=-0.19 $Y=1.655 $X2=1.835 $Y2=1.675
cc_104 VPB N_VPWR_c_560_n 3.14196e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_105 VPB N_VPWR_c_561_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.58
cc_106 VPB N_VPWR_c_562_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_563_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_564_n 0.0146078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_565_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_566_n 0.0176034f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_111 VPB N_VPWR_c_567_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.51
cc_112 VPB N_VPWR_c_568_n 0.0129339f $X=-0.19 $Y=1.655 $X2=1.745 $Y2=1.51
cc_113 VPB N_VPWR_c_569_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.592
cc_114 VPB N_VPWR_c_570_n 0.0574229f $X=-0.19 $Y=1.655 $X2=1.745 $Y2=1.592
cc_115 VPB N_VPWR_c_556_n 0.0511363f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.592
cc_116 VPB N_VPWR_c_572_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_573_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_574_n 0.0198795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_575_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB Y 0.00268566f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=1.592
cc_121 N_A3_M1029_g N_A2_M1006_g 0.018756f $X=1.765 $Y=0.765 $X2=0 $Y2=0
cc_122 N_A3_M1030_g N_A2_M1005_g 0.0136235f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_123 A3 N_A2_M1005_g 0.00524682f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_124 A3 N_A2_M1007_g 0.00382709f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_125 A3 N_A2_c_207_n 0.0305596f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A3_c_126_n N_A2_c_207_n 0.0249091f $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_127 A3 A2 0.0245779f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_128 A3 N_A_41_367#_c_456_n 0.0220965f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A3_c_126_n N_A_41_367#_c_456_n 0.00127488f $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A3_M1010_g N_A_41_367#_c_462_n 0.0122595f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A3_M1021_g N_A_41_367#_c_462_n 0.0122595f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_132 A3 N_A_41_367#_c_462_n 0.0428505f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A3_c_126_n N_A_41_367#_c_462_n 5.59536e-19 $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A3_M1022_g N_A_41_367#_c_466_n 0.0122595f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A3_M1030_g N_A_41_367#_c_466_n 0.0122595f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_136 A3 N_A_41_367#_c_466_n 0.0428505f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A3_c_126_n N_A_41_367#_c_466_n 5.59536e-19 $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_138 A3 N_A_41_367#_c_470_n 0.037789f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_139 A3 N_A_41_367#_c_471_n 0.0154121f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_140 N_A3_c_126_n N_A_41_367#_c_471_n 6.32755e-19 $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_141 A3 N_A_41_367#_c_473_n 0.0154122f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A3_M1010_g N_VPWR_c_557_n 0.0163213f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A3_M1021_g N_VPWR_c_557_n 0.0144369f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A3_M1022_g N_VPWR_c_557_n 6.77662e-19 $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A3_M1021_g N_VPWR_c_558_n 6.77662e-19 $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A3_M1022_g N_VPWR_c_558_n 0.0144369f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A3_M1030_g N_VPWR_c_558_n 0.0144369f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A3_M1030_g N_VPWR_c_559_n 6.77662e-19 $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A3_M1030_g N_VPWR_c_562_n 0.00486043f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A3_M1010_g N_VPWR_c_566_n 0.00486043f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A3_M1021_g N_VPWR_c_567_n 0.00486043f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A3_M1022_g N_VPWR_c_567_n 0.00486043f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A3_M1010_g N_VPWR_c_556_n 0.00923967f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A3_M1021_g N_VPWR_c_556_n 0.00824727f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A3_M1022_g N_VPWR_c_556_n 0.00824727f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A3_M1030_g N_VPWR_c_556_n 0.0082726f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A3_M1011_g N_A_27_69#_c_808_n 0.0035087f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_158 N_A3_M1011_g N_A_27_69#_c_809_n 0.0136535f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_159 N_A3_M1023_g N_A_27_69#_c_809_n 0.0130918f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_160 A3 N_A_27_69#_c_809_n 0.0499693f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_161 N_A3_c_126_n N_A_27_69#_c_809_n 0.0041186f $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_162 A3 N_A_27_69#_c_810_n 0.0163075f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_163 N_A3_c_126_n N_A_27_69#_c_810_n 0.00320949f $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A3_M1023_g N_A_27_69#_c_811_n 8.28776e-19 $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_165 N_A3_M1027_g N_A_27_69#_c_811_n 8.28776e-19 $X=1.335 $Y=0.765 $X2=0 $Y2=0
cc_166 N_A3_M1027_g N_A_27_69#_c_812_n 0.0130918f $X=1.335 $Y=0.765 $X2=0 $Y2=0
cc_167 N_A3_M1029_g N_A_27_69#_c_812_n 0.013073f $X=1.765 $Y=0.765 $X2=0 $Y2=0
cc_168 A3 N_A_27_69#_c_812_n 0.0492169f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A3_c_126_n N_A_27_69#_c_812_n 0.00406554f $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A3_M1029_g N_A_27_69#_c_813_n 8.28776e-19 $X=1.765 $Y=0.765 $X2=0 $Y2=0
cc_171 A3 N_A_27_69#_c_814_n 0.0479359f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_172 A3 N_A_27_69#_c_817_n 0.0160407f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_173 N_A3_c_126_n N_A_27_69#_c_817_n 0.00286879f $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_174 A3 N_A_27_69#_c_818_n 0.0167221f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A3_c_126_n N_A_27_69#_c_818_n 7.49468e-19 $X=1.835 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A3_M1011_g N_VGND_c_887_n 0.0129178f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_177 N_A3_M1023_g N_VGND_c_887_n 0.0101169f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_178 N_A3_M1027_g N_VGND_c_887_n 5.0028e-19 $X=1.335 $Y=0.765 $X2=0 $Y2=0
cc_179 N_A3_M1023_g N_VGND_c_888_n 5.0028e-19 $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_180 N_A3_M1027_g N_VGND_c_888_n 0.0101169f $X=1.335 $Y=0.765 $X2=0 $Y2=0
cc_181 N_A3_M1029_g N_VGND_c_888_n 0.0103777f $X=1.765 $Y=0.765 $X2=0 $Y2=0
cc_182 N_A3_M1029_g N_VGND_c_889_n 0.00400407f $X=1.765 $Y=0.765 $X2=0 $Y2=0
cc_183 N_A3_M1011_g N_VGND_c_892_n 0.00400407f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_184 N_A3_M1023_g N_VGND_c_893_n 0.00400407f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_185 N_A3_M1027_g N_VGND_c_893_n 0.00400407f $X=1.335 $Y=0.765 $X2=0 $Y2=0
cc_186 N_A3_M1011_g N_VGND_c_896_n 0.00796025f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_187 N_A3_M1023_g N_VGND_c_896_n 0.00774504f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_188 N_A3_M1027_g N_VGND_c_896_n 0.00774504f $X=1.335 $Y=0.765 $X2=0 $Y2=0
cc_189 N_A3_M1029_g N_VGND_c_896_n 0.00775088f $X=1.765 $Y=0.765 $X2=0 $Y2=0
cc_190 N_A3_M1029_g N_A_454_69#_c_991_n 2.32983e-19 $X=1.765 $Y=0.765 $X2=0
+ $Y2=0
cc_191 N_A2_M1031_g N_A1_M1000_g 0.0201857f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_192 A2 N_A1_c_298_n 3.3544e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A2_c_209_n N_A1_c_298_n 0.0246454f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_194 N_A2_M1005_g N_A_41_367#_c_470_n 0.0122595f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A2_M1007_g N_A_41_367#_c_470_n 0.0129323f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A2_c_207_n N_A_41_367#_c_470_n 5.59536e-19 $X=3.21 $Y=1.51 $X2=0 $Y2=0
cc_197 N_A2_M1019_g N_A_41_367#_c_477_n 0.0142694f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A2_c_206_n N_A_41_367#_c_477_n 0.00359182f $X=3.57 $Y=1.51 $X2=0 $Y2=0
cc_199 N_A2_M1031_g N_A_41_367#_c_477_n 0.00934319f $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_200 A2 N_A_41_367#_c_477_n 0.083451f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_201 N_A2_M1031_g N_A_41_367#_c_481_n 0.00626615f $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_202 N_A2_c_207_n N_A_41_367#_c_482_n 0.00208463f $X=3.21 $Y=1.51 $X2=0 $Y2=0
cc_203 A2 N_A_41_367#_c_482_n 0.00597035f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_204 N_A2_M1031_g N_A_41_367#_c_484_n 0.0089909f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A2_M1005_g N_VPWR_c_558_n 6.77662e-19 $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A2_M1005_g N_VPWR_c_559_n 0.0144369f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A2_M1007_g N_VPWR_c_559_n 0.0144345f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A2_M1019_g N_VPWR_c_559_n 6.77251e-19 $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A2_M1031_g N_VPWR_c_560_n 5.8762e-19 $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A2_M1005_g N_VPWR_c_562_n 0.00486043f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A2_M1031_g N_VPWR_c_564_n 0.00585385f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A2_M1007_g N_VPWR_c_568_n 0.00486043f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A2_M1019_g N_VPWR_c_568_n 0.00486043f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A2_M1005_g N_VPWR_c_556_n 0.0082726f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A2_M1007_g N_VPWR_c_556_n 0.00824727f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A2_M1019_g N_VPWR_c_556_n 0.00819843f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A2_M1031_g N_VPWR_c_556_n 0.00749215f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A2_M1007_g N_VPWR_c_574_n 6.92339e-19 $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A2_M1019_g N_VPWR_c_574_n 0.0190023f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A2_M1031_g N_VPWR_c_574_n 0.0112763f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A2_M1031_g Y 6.59985e-19 $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A2_M1028_g N_Y_c_690_n 0.00110856f $X=3.645 $Y=0.765 $X2=0 $Y2=0
cc_223 N_A2_M1028_g Y 0.00205613f $X=3.645 $Y=0.765 $X2=0 $Y2=0
cc_224 A2 Y 0.0257635f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_225 N_A2_c_209_n Y 0.00873244f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_226 N_A2_M1006_g N_A_27_69#_c_813_n 8.28478e-19 $X=2.195 $Y=0.765 $X2=0 $Y2=0
cc_227 N_A2_M1006_g N_A_27_69#_c_814_n 0.013073f $X=2.195 $Y=0.765 $X2=0 $Y2=0
cc_228 N_A2_M1009_g N_A_27_69#_c_814_n 0.0127931f $X=2.625 $Y=0.765 $X2=0 $Y2=0
cc_229 N_A2_c_207_n N_A_27_69#_c_814_n 0.00276559f $X=3.21 $Y=1.51 $X2=0 $Y2=0
cc_230 N_A2_M1020_g N_A_27_69#_c_843_n 0.00696504f $X=3.135 $Y=0.765 $X2=0 $Y2=0
cc_231 N_A2_M1028_g N_A_27_69#_c_843_n 5.37284e-19 $X=3.645 $Y=0.765 $X2=0 $Y2=0
cc_232 N_A2_M1020_g N_A_27_69#_c_815_n 0.00966312f $X=3.135 $Y=0.765 $X2=0 $Y2=0
cc_233 N_A2_c_206_n N_A_27_69#_c_815_n 0.0044365f $X=3.57 $Y=1.51 $X2=0 $Y2=0
cc_234 N_A2_M1028_g N_A_27_69#_c_815_n 0.0143665f $X=3.645 $Y=0.765 $X2=0 $Y2=0
cc_235 A2 N_A_27_69#_c_815_n 0.0785296f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_236 N_A2_c_209_n N_A_27_69#_c_815_n 0.0105559f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_237 N_A2_M1020_g N_A_27_69#_c_819_n 0.00174458f $X=3.135 $Y=0.765 $X2=0 $Y2=0
cc_238 N_A2_c_207_n N_A_27_69#_c_819_n 0.00604839f $X=3.21 $Y=1.51 $X2=0 $Y2=0
cc_239 A2 N_A_27_69#_c_819_n 0.0129421f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_240 N_A2_M1006_g N_VGND_c_888_n 6.53017e-19 $X=2.195 $Y=0.765 $X2=0 $Y2=0
cc_241 N_A2_M1006_g N_VGND_c_889_n 0.00450424f $X=2.195 $Y=0.765 $X2=0 $Y2=0
cc_242 N_A2_M1009_g N_VGND_c_889_n 0.00291444f $X=2.625 $Y=0.765 $X2=0 $Y2=0
cc_243 N_A2_M1020_g N_VGND_c_889_n 0.0029147f $X=3.135 $Y=0.765 $X2=0 $Y2=0
cc_244 N_A2_M1028_g N_VGND_c_889_n 0.00291444f $X=3.645 $Y=0.765 $X2=0 $Y2=0
cc_245 N_A2_M1006_g N_VGND_c_896_n 0.00862457f $X=2.195 $Y=0.765 $X2=0 $Y2=0
cc_246 N_A2_M1009_g N_VGND_c_896_n 0.00403101f $X=2.625 $Y=0.765 $X2=0 $Y2=0
cc_247 N_A2_M1020_g N_VGND_c_896_n 0.00407574f $X=3.135 $Y=0.765 $X2=0 $Y2=0
cc_248 N_A2_M1028_g N_VGND_c_896_n 0.00433094f $X=3.645 $Y=0.765 $X2=0 $Y2=0
cc_249 N_A2_M1006_g N_A_454_69#_c_997_n 0.00527422f $X=2.195 $Y=0.765 $X2=0
+ $Y2=0
cc_250 N_A2_M1009_g N_A_454_69#_c_997_n 0.00697012f $X=2.625 $Y=0.765 $X2=0
+ $Y2=0
cc_251 N_A2_M1020_g N_A_454_69#_c_997_n 5.60912e-19 $X=3.135 $Y=0.765 $X2=0
+ $Y2=0
cc_252 N_A2_M1009_g N_A_454_69#_c_990_n 0.00867861f $X=2.625 $Y=0.765 $X2=0
+ $Y2=0
cc_253 N_A2_M1020_g N_A_454_69#_c_990_n 0.0120458f $X=3.135 $Y=0.765 $X2=0 $Y2=0
cc_254 N_A2_M1006_g N_A_454_69#_c_991_n 0.00344817f $X=2.195 $Y=0.765 $X2=0
+ $Y2=0
cc_255 N_A2_M1009_g N_A_454_69#_c_991_n 0.00159238f $X=2.625 $Y=0.765 $X2=0
+ $Y2=0
cc_256 N_A2_M1028_g N_A_454_69#_c_1004_n 0.0111491f $X=3.645 $Y=0.765 $X2=0
+ $Y2=0
cc_257 N_A2_M1028_g N_A_454_69#_c_992_n 0.0102755f $X=3.645 $Y=0.765 $X2=0 $Y2=0
cc_258 N_A2_M1028_g N_A_454_69#_c_994_n 0.0018274f $X=3.645 $Y=0.765 $X2=0 $Y2=0
cc_259 A1 N_B1_M1002_g 0.00547822f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_260 N_A1_M1018_g N_B1_M1013_g 0.0154989f $X=5.965 $Y=0.745 $X2=0 $Y2=0
cc_261 A1 N_B1_M1003_g 6.91425e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_262 A1 B1 0.0282902f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_263 N_A1_M1017_g N_B1_c_386_n 0.0374825f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_264 A1 N_B1_c_386_n 0.0193982f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_265 N_A1_c_298_n N_B1_c_386_n 0.0246561f $X=5.815 $Y=1.485 $X2=0 $Y2=0
cc_266 N_A1_M1000_g N_A_41_367#_c_485_n 0.0122533f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_267 N_A1_M1008_g N_A_41_367#_c_485_n 0.0122595f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A1_M1012_g N_A_41_367#_c_487_n 0.0122595f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A1_M1017_g N_A_41_367#_c_487_n 0.0122595f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_270 N_A1_M1000_g N_VPWR_c_560_n 0.0106975f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_271 N_A1_M1008_g N_VPWR_c_560_n 0.0106305f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A1_M1012_g N_VPWR_c_560_n 5.75816e-19 $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A1_M1008_g N_VPWR_c_561_n 5.75816e-19 $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_274 N_A1_M1012_g N_VPWR_c_561_n 0.0106305f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A1_M1017_g N_VPWR_c_561_n 0.011872f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A1_M1000_g N_VPWR_c_564_n 0.00486043f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A1_M1008_g N_VPWR_c_569_n 0.00486043f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_278 N_A1_M1012_g N_VPWR_c_569_n 0.00486043f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_279 N_A1_M1017_g N_VPWR_c_570_n 0.00486043f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_280 N_A1_M1000_g N_VPWR_c_556_n 0.0082726f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_281 N_A1_M1008_g N_VPWR_c_556_n 0.00824727f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_282 N_A1_M1012_g N_VPWR_c_556_n 0.00824727f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_283 N_A1_M1017_g N_VPWR_c_556_n 0.00845345f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_284 N_A1_M1001_g N_Y_c_680_n 0.00942318f $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_285 N_A1_M1004_g N_Y_c_680_n 0.0161584f $X=5.105 $Y=0.745 $X2=0 $Y2=0
cc_286 A1 N_Y_c_680_n 0.022161f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_287 N_A1_c_298_n N_Y_c_680_n 0.00387295f $X=5.815 $Y=1.485 $X2=0 $Y2=0
cc_288 N_A1_M1008_g N_Y_c_702_n 0.010446f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_289 N_A1_M1012_g N_Y_c_702_n 0.0104926f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_290 N_A1_M1017_g N_Y_c_702_n 0.0108739f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_291 A1 N_Y_c_702_n 0.101202f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_292 N_A1_c_298_n N_Y_c_702_n 0.00489787f $X=5.815 $Y=1.485 $X2=0 $Y2=0
cc_293 N_A1_M1016_g N_Y_c_681_n 0.0106492f $X=5.535 $Y=0.745 $X2=0 $Y2=0
cc_294 N_A1_M1018_g N_Y_c_681_n 0.0151126f $X=5.965 $Y=0.745 $X2=0 $Y2=0
cc_295 A1 N_Y_c_681_n 0.0442852f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_296 N_A1_c_298_n N_Y_c_681_n 0.00308478f $X=5.815 $Y=1.485 $X2=0 $Y2=0
cc_297 N_A1_M1018_g N_Y_c_682_n 0.0011129f $X=5.965 $Y=0.745 $X2=0 $Y2=0
cc_298 A1 N_Y_c_683_n 0.0215978f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_299 N_A1_M1001_g N_Y_c_687_n 9.5728e-19 $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_300 N_A1_M1004_g N_Y_c_687_n 0.00774408f $X=5.105 $Y=0.745 $X2=0 $Y2=0
cc_301 N_A1_M1016_g N_Y_c_687_n 0.00879921f $X=5.535 $Y=0.745 $X2=0 $Y2=0
cc_302 N_A1_M1018_g N_Y_c_687_n 6.26039e-19 $X=5.965 $Y=0.745 $X2=0 $Y2=0
cc_303 A1 N_Y_c_687_n 0.0275185f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_304 N_A1_c_298_n N_Y_c_687_n 0.00317902f $X=5.815 $Y=1.485 $X2=0 $Y2=0
cc_305 A1 N_Y_c_688_n 0.017785f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_306 N_A1_M1017_g N_Y_c_720_n 7.26539e-19 $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_307 A1 N_Y_c_720_n 0.0137864f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_308 N_A1_M1000_g Y 0.00761892f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_309 N_A1_M1001_g N_Y_c_690_n 0.00822886f $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_310 N_A1_M1000_g Y 0.00717106f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_311 N_A1_M1001_g Y 0.00166002f $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_312 N_A1_M1008_g Y 0.00439147f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_313 N_A1_M1004_g Y 2.18893e-19 $X=5.105 $Y=0.745 $X2=0 $Y2=0
cc_314 A1 Y 0.0291974f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_315 N_A1_c_298_n Y 0.0236034f $X=5.815 $Y=1.485 $X2=0 $Y2=0
cc_316 N_A1_M1001_g N_A_27_69#_c_815_n 6.17077e-19 $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_317 N_A1_M1001_g N_A_27_69#_c_816_n 0.00535917f $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_318 N_A1_M1001_g N_VGND_c_889_n 0.00303788f $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_319 N_A1_M1004_g N_VGND_c_889_n 0.00302501f $X=5.105 $Y=0.745 $X2=0 $Y2=0
cc_320 N_A1_M1016_g N_VGND_c_889_n 0.00302501f $X=5.535 $Y=0.745 $X2=0 $Y2=0
cc_321 N_A1_M1018_g N_VGND_c_889_n 0.00499542f $X=5.965 $Y=0.745 $X2=0 $Y2=0
cc_322 N_A1_M1018_g N_VGND_c_890_n 7.00223e-19 $X=5.965 $Y=0.745 $X2=0 $Y2=0
cc_323 N_A1_M1001_g N_VGND_c_896_n 0.00483749f $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_324 N_A1_M1004_g N_VGND_c_896_n 0.00433762f $X=5.105 $Y=0.745 $X2=0 $Y2=0
cc_325 N_A1_M1016_g N_VGND_c_896_n 0.00434671f $X=5.535 $Y=0.745 $X2=0 $Y2=0
cc_326 N_A1_M1018_g N_VGND_c_896_n 0.00991536f $X=5.965 $Y=0.745 $X2=0 $Y2=0
cc_327 N_A1_M1001_g N_A_454_69#_c_992_n 0.010103f $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_328 N_A1_M1004_g N_A_454_69#_c_993_n 0.0086703f $X=5.105 $Y=0.745 $X2=0 $Y2=0
cc_329 N_A1_M1016_g N_A_454_69#_c_993_n 0.0106826f $X=5.535 $Y=0.745 $X2=0 $Y2=0
cc_330 N_A1_M1018_g N_A_454_69#_c_993_n 0.00129509f $X=5.965 $Y=0.745 $X2=0
+ $Y2=0
cc_331 N_A1_M1001_g N_A_454_69#_c_995_n 0.0108279f $X=4.675 $Y=0.745 $X2=0 $Y2=0
cc_332 N_B1_M1002_g N_A_41_367#_c_489_n 0.0136509f $X=6.325 $Y=2.465 $X2=0 $Y2=0
cc_333 N_B1_M1003_g N_A_41_367#_c_489_n 0.0115031f $X=6.755 $Y=2.465 $X2=0 $Y2=0
cc_334 N_B1_M1014_g N_A_41_367#_c_491_n 0.0115031f $X=7.185 $Y=2.465 $X2=0 $Y2=0
cc_335 N_B1_M1026_g N_A_41_367#_c_491_n 0.0115031f $X=7.615 $Y=2.465 $X2=0 $Y2=0
cc_336 B1 N_A_41_367#_c_459_n 0.0216386f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_337 N_B1_M1002_g N_VPWR_c_561_n 0.00120156f $X=6.325 $Y=2.465 $X2=0 $Y2=0
cc_338 N_B1_M1002_g N_VPWR_c_570_n 0.00357877f $X=6.325 $Y=2.465 $X2=0 $Y2=0
cc_339 N_B1_M1003_g N_VPWR_c_570_n 0.00357877f $X=6.755 $Y=2.465 $X2=0 $Y2=0
cc_340 N_B1_M1014_g N_VPWR_c_570_n 0.00357877f $X=7.185 $Y=2.465 $X2=0 $Y2=0
cc_341 N_B1_M1026_g N_VPWR_c_570_n 0.00357877f $X=7.615 $Y=2.465 $X2=0 $Y2=0
cc_342 N_B1_M1002_g N_VPWR_c_556_n 0.00564397f $X=6.325 $Y=2.465 $X2=0 $Y2=0
cc_343 N_B1_M1003_g N_VPWR_c_556_n 0.0053512f $X=6.755 $Y=2.465 $X2=0 $Y2=0
cc_344 N_B1_M1014_g N_VPWR_c_556_n 0.0053512f $X=7.185 $Y=2.465 $X2=0 $Y2=0
cc_345 N_B1_M1026_g N_VPWR_c_556_n 0.00634361f $X=7.615 $Y=2.465 $X2=0 $Y2=0
cc_346 N_B1_M1002_g N_Y_c_702_n 0.0115313f $X=6.325 $Y=2.465 $X2=0 $Y2=0
cc_347 N_B1_M1013_g N_Y_c_682_n 0.00106024f $X=6.395 $Y=0.745 $X2=0 $Y2=0
cc_348 N_B1_M1013_g N_Y_c_683_n 0.0136107f $X=6.395 $Y=0.745 $X2=0 $Y2=0
cc_349 N_B1_M1015_g N_Y_c_683_n 0.0136351f $X=6.825 $Y=0.745 $X2=0 $Y2=0
cc_350 B1 N_Y_c_683_n 0.0141986f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_351 N_B1_c_386_n N_Y_c_683_n 0.00458192f $X=7.615 $Y=1.515 $X2=0 $Y2=0
cc_352 N_B1_M1003_g N_Y_c_736_n 0.0124938f $X=6.755 $Y=2.465 $X2=0 $Y2=0
cc_353 N_B1_M1014_g N_Y_c_736_n 0.01115f $X=7.185 $Y=2.465 $X2=0 $Y2=0
cc_354 B1 N_Y_c_736_n 0.0325079f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_355 N_B1_c_386_n N_Y_c_736_n 5.46532e-19 $X=7.615 $Y=1.515 $X2=0 $Y2=0
cc_356 N_B1_M1015_g N_Y_c_684_n 0.00105889f $X=6.825 $Y=0.745 $X2=0 $Y2=0
cc_357 N_B1_M1024_g N_Y_c_684_n 0.00105889f $X=7.255 $Y=0.745 $X2=0 $Y2=0
cc_358 N_B1_M1024_g N_Y_c_685_n 0.0136351f $X=7.255 $Y=0.745 $X2=0 $Y2=0
cc_359 N_B1_M1025_g N_Y_c_685_n 0.0143619f $X=7.685 $Y=0.745 $X2=0 $Y2=0
cc_360 B1 N_Y_c_685_n 0.0724279f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_361 N_B1_c_386_n N_Y_c_685_n 0.00277354f $X=7.615 $Y=1.515 $X2=0 $Y2=0
cc_362 N_B1_M1025_g N_Y_c_686_n 0.0035087f $X=7.685 $Y=0.745 $X2=0 $Y2=0
cc_363 N_B1_M1002_g N_Y_c_720_n 0.0102656f $X=6.325 $Y=2.465 $X2=0 $Y2=0
cc_364 N_B1_M1003_g N_Y_c_720_n 0.0107882f $X=6.755 $Y=2.465 $X2=0 $Y2=0
cc_365 N_B1_M1014_g N_Y_c_720_n 5.60744e-19 $X=7.185 $Y=2.465 $X2=0 $Y2=0
cc_366 N_B1_c_386_n N_Y_c_720_n 0.00146913f $X=7.615 $Y=1.515 $X2=0 $Y2=0
cc_367 B1 N_Y_c_689_n 0.0161047f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_368 N_B1_c_386_n N_Y_c_689_n 0.00287331f $X=7.615 $Y=1.515 $X2=0 $Y2=0
cc_369 N_B1_M1003_g N_Y_c_753_n 5.60744e-19 $X=6.755 $Y=2.465 $X2=0 $Y2=0
cc_370 N_B1_M1014_g N_Y_c_753_n 0.00995034f $X=7.185 $Y=2.465 $X2=0 $Y2=0
cc_371 N_B1_M1026_g N_Y_c_753_n 0.0106824f $X=7.615 $Y=2.465 $X2=0 $Y2=0
cc_372 B1 N_Y_c_753_n 0.023215f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_373 N_B1_c_386_n N_Y_c_753_n 6.18336e-19 $X=7.615 $Y=1.515 $X2=0 $Y2=0
cc_374 N_B1_M1013_g N_VGND_c_889_n 0.00414769f $X=6.395 $Y=0.745 $X2=0 $Y2=0
cc_375 N_B1_M1013_g N_VGND_c_890_n 0.0104336f $X=6.395 $Y=0.745 $X2=0 $Y2=0
cc_376 N_B1_M1015_g N_VGND_c_890_n 0.00997431f $X=6.825 $Y=0.745 $X2=0 $Y2=0
cc_377 N_B1_M1024_g N_VGND_c_890_n 4.56253e-19 $X=7.255 $Y=0.745 $X2=0 $Y2=0
cc_378 N_B1_M1015_g N_VGND_c_891_n 4.56253e-19 $X=6.825 $Y=0.745 $X2=0 $Y2=0
cc_379 N_B1_M1024_g N_VGND_c_891_n 0.00997431f $X=7.255 $Y=0.745 $X2=0 $Y2=0
cc_380 N_B1_M1025_g N_VGND_c_891_n 0.0125815f $X=7.685 $Y=0.745 $X2=0 $Y2=0
cc_381 N_B1_M1015_g N_VGND_c_894_n 0.00414769f $X=6.825 $Y=0.745 $X2=0 $Y2=0
cc_382 N_B1_M1024_g N_VGND_c_894_n 0.00414769f $X=7.255 $Y=0.745 $X2=0 $Y2=0
cc_383 N_B1_M1025_g N_VGND_c_895_n 0.00414769f $X=7.685 $Y=0.745 $X2=0 $Y2=0
cc_384 N_B1_M1013_g N_VGND_c_896_n 0.0078848f $X=6.395 $Y=0.745 $X2=0 $Y2=0
cc_385 N_B1_M1015_g N_VGND_c_896_n 0.00787505f $X=6.825 $Y=0.745 $X2=0 $Y2=0
cc_386 N_B1_M1024_g N_VGND_c_896_n 0.00787505f $X=7.255 $Y=0.745 $X2=0 $Y2=0
cc_387 N_B1_M1025_g N_VGND_c_896_n 0.00823375f $X=7.685 $Y=0.745 $X2=0 $Y2=0
cc_388 N_A_41_367#_c_462_n N_VPWR_M1010_s 0.00333177f $X=1.095 $Y=2.015
+ $X2=-0.19 $Y2=1.655
cc_389 N_A_41_367#_c_466_n N_VPWR_M1022_s 0.00333177f $X=1.955 $Y=2.015 $X2=0
+ $Y2=0
cc_390 N_A_41_367#_c_470_n N_VPWR_M1005_d 0.00333177f $X=2.815 $Y=2.015 $X2=0
+ $Y2=0
cc_391 N_A_41_367#_c_477_n N_VPWR_M1019_d 0.0189786f $X=4.015 $Y=2.015 $X2=0
+ $Y2=0
cc_392 N_A_41_367#_c_485_n N_VPWR_M1000_s 0.00343498f $X=5.075 $Y=2.375 $X2=0
+ $Y2=0
cc_393 N_A_41_367#_c_487_n N_VPWR_M1012_s 0.00344593f $X=5.935 $Y=2.375 $X2=0
+ $Y2=0
cc_394 N_A_41_367#_c_462_n N_VPWR_c_557_n 0.0170777f $X=1.095 $Y=2.015 $X2=0
+ $Y2=0
cc_395 N_A_41_367#_c_466_n N_VPWR_c_558_n 0.0170777f $X=1.955 $Y=2.015 $X2=0
+ $Y2=0
cc_396 N_A_41_367#_c_470_n N_VPWR_c_559_n 0.0170777f $X=2.815 $Y=2.015 $X2=0
+ $Y2=0
cc_397 N_A_41_367#_c_485_n N_VPWR_c_560_n 0.0170777f $X=5.075 $Y=2.375 $X2=0
+ $Y2=0
cc_398 N_A_41_367#_c_487_n N_VPWR_c_561_n 0.0170777f $X=5.935 $Y=2.375 $X2=0
+ $Y2=0
cc_399 N_A_41_367#_c_505_p N_VPWR_c_562_n 0.0124525f $X=2.05 $Y=2.91 $X2=0 $Y2=0
cc_400 N_A_41_367#_c_506_p N_VPWR_c_564_n 0.0134175f $X=4.295 $Y=2.47 $X2=0
+ $Y2=0
cc_401 N_A_41_367#_c_457_n N_VPWR_c_566_n 0.0178111f $X=0.33 $Y=2.91 $X2=0 $Y2=0
cc_402 N_A_41_367#_c_508_p N_VPWR_c_567_n 0.0124525f $X=1.19 $Y=2.91 $X2=0 $Y2=0
cc_403 N_A_41_367#_c_509_p N_VPWR_c_568_n 0.0124525f $X=2.91 $Y=2.91 $X2=0 $Y2=0
cc_404 N_A_41_367#_c_510_p N_VPWR_c_569_n 0.0124525f $X=5.17 $Y=2.455 $X2=0
+ $Y2=0
cc_405 N_A_41_367#_c_489_n N_VPWR_c_570_n 0.0361434f $X=6.875 $Y=2.99 $X2=0
+ $Y2=0
cc_406 N_A_41_367#_c_512_p N_VPWR_c_570_n 0.0181484f $X=6.205 $Y=2.99 $X2=0
+ $Y2=0
cc_407 N_A_41_367#_c_491_n N_VPWR_c_570_n 0.0364699f $X=7.745 $Y=2.99 $X2=0
+ $Y2=0
cc_408 N_A_41_367#_c_458_n N_VPWR_c_570_n 0.0175634f $X=7.87 $Y=2.905 $X2=0
+ $Y2=0
cc_409 N_A_41_367#_c_515_p N_VPWR_c_570_n 0.0125234f $X=6.97 $Y=2.99 $X2=0 $Y2=0
cc_410 N_A_41_367#_M1010_d N_VPWR_c_556_n 0.00371702f $X=0.205 $Y=1.835 $X2=0
+ $Y2=0
cc_411 N_A_41_367#_M1021_d N_VPWR_c_556_n 0.00536646f $X=1.05 $Y=1.835 $X2=0
+ $Y2=0
cc_412 N_A_41_367#_M1030_d N_VPWR_c_556_n 0.00536646f $X=1.91 $Y=1.835 $X2=0
+ $Y2=0
cc_413 N_A_41_367#_M1007_s N_VPWR_c_556_n 0.00536646f $X=2.77 $Y=1.835 $X2=0
+ $Y2=0
cc_414 N_A_41_367#_M1031_s N_VPWR_c_556_n 0.00386217f $X=4.17 $Y=1.835 $X2=0
+ $Y2=0
cc_415 N_A_41_367#_M1008_d N_VPWR_c_556_n 0.00536646f $X=5.03 $Y=1.835 $X2=0
+ $Y2=0
cc_416 N_A_41_367#_M1017_d N_VPWR_c_556_n 0.00441765f $X=5.89 $Y=1.835 $X2=0
+ $Y2=0
cc_417 N_A_41_367#_M1003_s N_VPWR_c_556_n 0.00223565f $X=6.83 $Y=1.835 $X2=0
+ $Y2=0
cc_418 N_A_41_367#_M1026_s N_VPWR_c_556_n 0.00215162f $X=7.69 $Y=1.835 $X2=0
+ $Y2=0
cc_419 N_A_41_367#_c_457_n N_VPWR_c_556_n 0.0100304f $X=0.33 $Y=2.91 $X2=0 $Y2=0
cc_420 N_A_41_367#_c_508_p N_VPWR_c_556_n 0.00730901f $X=1.19 $Y=2.91 $X2=0
+ $Y2=0
cc_421 N_A_41_367#_c_505_p N_VPWR_c_556_n 0.00730901f $X=2.05 $Y=2.91 $X2=0
+ $Y2=0
cc_422 N_A_41_367#_c_509_p N_VPWR_c_556_n 0.00730901f $X=2.91 $Y=2.91 $X2=0
+ $Y2=0
cc_423 N_A_41_367#_c_506_p N_VPWR_c_556_n 0.00844946f $X=4.295 $Y=2.47 $X2=0
+ $Y2=0
cc_424 N_A_41_367#_c_489_n N_VPWR_c_556_n 0.0237467f $X=6.875 $Y=2.99 $X2=0
+ $Y2=0
cc_425 N_A_41_367#_c_512_p N_VPWR_c_556_n 0.010497f $X=6.205 $Y=2.99 $X2=0 $Y2=0
cc_426 N_A_41_367#_c_491_n N_VPWR_c_556_n 0.024052f $X=7.745 $Y=2.99 $X2=0 $Y2=0
cc_427 N_A_41_367#_c_458_n N_VPWR_c_556_n 0.00970886f $X=7.87 $Y=2.905 $X2=0
+ $Y2=0
cc_428 N_A_41_367#_c_484_n N_VPWR_c_556_n 0.00465535f $X=4.405 $Y=2.38 $X2=0
+ $Y2=0
cc_429 N_A_41_367#_c_510_p N_VPWR_c_556_n 0.00730901f $X=5.17 $Y=2.455 $X2=0
+ $Y2=0
cc_430 N_A_41_367#_c_515_p N_VPWR_c_556_n 0.00738676f $X=6.97 $Y=2.99 $X2=0
+ $Y2=0
cc_431 N_A_41_367#_c_477_n N_VPWR_c_574_n 0.0537561f $X=4.015 $Y=2.015 $X2=0
+ $Y2=0
cc_432 N_A_41_367#_c_489_n N_Y_M1002_d 0.00332344f $X=6.875 $Y=2.99 $X2=0 $Y2=0
cc_433 N_A_41_367#_c_491_n N_Y_M1014_d 0.00332344f $X=7.745 $Y=2.99 $X2=0 $Y2=0
cc_434 N_A_41_367#_M1008_d N_Y_c_702_n 0.00333871f $X=5.03 $Y=1.835 $X2=0 $Y2=0
cc_435 N_A_41_367#_M1017_d N_Y_c_702_n 0.00505525f $X=5.89 $Y=1.835 $X2=0 $Y2=0
cc_436 N_A_41_367#_c_485_n N_Y_c_702_n 0.0186676f $X=5.075 $Y=2.375 $X2=0 $Y2=0
cc_437 N_A_41_367#_c_487_n N_Y_c_702_n 0.0323235f $X=5.935 $Y=2.375 $X2=0 $Y2=0
cc_438 N_A_41_367#_c_544_p N_Y_c_702_n 0.0200142f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_439 N_A_41_367#_c_510_p N_Y_c_702_n 0.0135055f $X=5.17 $Y=2.455 $X2=0 $Y2=0
cc_440 N_A_41_367#_M1003_s N_Y_c_736_n 0.00333523f $X=6.83 $Y=1.835 $X2=0 $Y2=0
cc_441 N_A_41_367#_c_547_p N_Y_c_736_n 0.0135055f $X=6.97 $Y=2.455 $X2=0 $Y2=0
cc_442 N_A_41_367#_c_489_n N_Y_c_720_n 0.0159805f $X=6.875 $Y=2.99 $X2=0 $Y2=0
cc_443 N_A_41_367#_c_491_n N_Y_c_753_n 0.0159805f $X=7.745 $Y=2.99 $X2=0 $Y2=0
cc_444 N_A_41_367#_M1031_s Y 0.00189618f $X=4.17 $Y=1.835 $X2=0 $Y2=0
cc_445 N_A_41_367#_c_484_n Y 0.0183112f $X=4.405 $Y=2.38 $X2=0 $Y2=0
cc_446 N_A_41_367#_M1031_s Y 0.0013777f $X=4.17 $Y=1.835 $X2=0 $Y2=0
cc_447 N_A_41_367#_c_470_n N_A_27_69#_c_814_n 7.37357e-19 $X=2.815 $Y=2.015
+ $X2=0 $Y2=0
cc_448 N_A_41_367#_c_470_n N_A_27_69#_c_819_n 0.00120074f $X=2.815 $Y=2.015
+ $X2=0 $Y2=0
cc_449 N_A_41_367#_c_482_n N_A_27_69#_c_819_n 0.00361646f $X=2.91 $Y=2.095 $X2=0
+ $Y2=0
cc_450 N_VPWR_c_556_n N_Y_M1002_d 0.00225186f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_451 N_VPWR_c_556_n N_Y_M1014_d 0.00225186f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_452 N_VPWR_M1000_s N_Y_c_702_n 0.00356282f $X=4.6 $Y=1.835 $X2=0 $Y2=0
cc_453 N_VPWR_M1012_s N_Y_c_702_n 0.00334301f $X=5.46 $Y=1.835 $X2=0 $Y2=0
cc_454 N_VPWR_M1000_s Y 5.21393e-19 $X=4.6 $Y=1.835 $X2=0 $Y2=0
cc_455 N_VPWR_M1000_s Y 0.00144754f $X=4.6 $Y=1.835 $X2=0 $Y2=0
cc_456 N_Y_c_690_n N_A_27_69#_c_815_n 0.0119903f $X=4.53 $Y=1.255 $X2=0 $Y2=0
cc_457 N_Y_c_690_n N_A_27_69#_c_816_n 0.0160498f $X=4.53 $Y=1.255 $X2=0 $Y2=0
cc_458 N_Y_c_683_n N_VGND_M1013_d 0.00176773f $X=6.945 $Y=1.165 $X2=0 $Y2=0
cc_459 N_Y_c_685_n N_VGND_M1024_d 0.00176773f $X=7.815 $Y=1.165 $X2=0 $Y2=0
cc_460 N_Y_c_682_n N_VGND_c_889_n 0.011926f $X=6.18 $Y=0.45 $X2=0 $Y2=0
cc_461 N_Y_c_682_n N_VGND_c_890_n 0.0247679f $X=6.18 $Y=0.45 $X2=0 $Y2=0
cc_462 N_Y_c_683_n N_VGND_c_890_n 0.0171443f $X=6.945 $Y=1.165 $X2=0 $Y2=0
cc_463 N_Y_c_684_n N_VGND_c_890_n 0.0247562f $X=7.04 $Y=0.45 $X2=0 $Y2=0
cc_464 N_Y_c_684_n N_VGND_c_891_n 0.0247562f $X=7.04 $Y=0.45 $X2=0 $Y2=0
cc_465 N_Y_c_685_n N_VGND_c_891_n 0.0171443f $X=7.815 $Y=1.165 $X2=0 $Y2=0
cc_466 N_Y_c_686_n N_VGND_c_891_n 0.0222328f $X=7.9 $Y=0.47 $X2=0 $Y2=0
cc_467 N_Y_c_684_n N_VGND_c_894_n 0.0113237f $X=7.04 $Y=0.45 $X2=0 $Y2=0
cc_468 N_Y_c_686_n N_VGND_c_895_n 0.0134916f $X=7.9 $Y=0.47 $X2=0 $Y2=0
cc_469 N_Y_c_680_n N_VGND_c_896_n 0.00110108f $X=5.155 $Y=1.047 $X2=0 $Y2=0
cc_470 N_Y_c_682_n N_VGND_c_896_n 0.00758479f $X=6.18 $Y=0.45 $X2=0 $Y2=0
cc_471 N_Y_c_684_n N_VGND_c_896_n 0.00720172f $X=7.04 $Y=0.45 $X2=0 $Y2=0
cc_472 N_Y_c_686_n N_VGND_c_896_n 0.0093995f $X=7.9 $Y=0.47 $X2=0 $Y2=0
cc_473 N_Y_c_680_n N_A_454_69#_M1001_d 0.00178913f $X=5.155 $Y=1.047 $X2=0 $Y2=0
cc_474 N_Y_c_681_n N_A_454_69#_M1016_d 0.00177483f $X=6.075 $Y=1.152 $X2=0 $Y2=0
cc_475 N_Y_M1001_s N_A_454_69#_c_992_n 0.00430028f $X=4.335 $Y=0.325 $X2=0 $Y2=0
cc_476 N_Y_c_680_n N_A_454_69#_c_992_n 5.84976e-19 $X=5.155 $Y=1.047 $X2=0 $Y2=0
cc_477 N_Y_c_690_n N_A_454_69#_c_992_n 0.0098888f $X=4.53 $Y=1.255 $X2=0 $Y2=0
cc_478 N_Y_M1004_s N_A_454_69#_c_993_n 0.00176461f $X=5.18 $Y=0.325 $X2=0 $Y2=0
cc_479 N_Y_c_680_n N_A_454_69#_c_993_n 0.00372353f $X=5.155 $Y=1.047 $X2=0 $Y2=0
cc_480 N_Y_c_681_n N_A_454_69#_c_993_n 0.00291681f $X=6.075 $Y=1.152 $X2=0 $Y2=0
cc_481 N_Y_c_682_n N_A_454_69#_c_993_n 0.00277472f $X=6.18 $Y=0.45 $X2=0 $Y2=0
cc_482 N_Y_c_687_n N_A_454_69#_c_993_n 0.0159436f $X=5.32 $Y=0.68 $X2=0 $Y2=0
cc_483 N_Y_c_681_n N_A_454_69#_c_1022_n 0.0135853f $X=6.075 $Y=1.152 $X2=0 $Y2=0
cc_484 N_Y_c_680_n N_A_454_69#_c_995_n 0.0152954f $X=5.155 $Y=1.047 $X2=0 $Y2=0
cc_485 N_A_27_69#_c_809_n N_VGND_M1011_d 0.00176461f $X=1.025 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_486 N_A_27_69#_c_812_n N_VGND_M1027_d 0.00176461f $X=1.885 $Y=1.17 $X2=0
+ $Y2=0
cc_487 N_A_27_69#_c_808_n N_VGND_c_887_n 0.0218743f $X=0.26 $Y=0.49 $X2=0 $Y2=0
cc_488 N_A_27_69#_c_809_n N_VGND_c_887_n 0.0170777f $X=1.025 $Y=1.17 $X2=0 $Y2=0
cc_489 N_A_27_69#_c_811_n N_VGND_c_887_n 0.0228652f $X=1.12 $Y=0.49 $X2=0 $Y2=0
cc_490 N_A_27_69#_c_811_n N_VGND_c_888_n 0.0228652f $X=1.12 $Y=0.49 $X2=0 $Y2=0
cc_491 N_A_27_69#_c_812_n N_VGND_c_888_n 0.0170777f $X=1.885 $Y=1.17 $X2=0 $Y2=0
cc_492 N_A_27_69#_c_813_n N_VGND_c_888_n 0.0228652f $X=1.98 $Y=0.49 $X2=0 $Y2=0
cc_493 N_A_27_69#_c_813_n N_VGND_c_889_n 0.00932149f $X=1.98 $Y=0.49 $X2=0 $Y2=0
cc_494 N_A_27_69#_c_808_n N_VGND_c_892_n 0.0122964f $X=0.26 $Y=0.49 $X2=0 $Y2=0
cc_495 N_A_27_69#_c_811_n N_VGND_c_893_n 0.00932149f $X=1.12 $Y=0.49 $X2=0 $Y2=0
cc_496 N_A_27_69#_c_808_n N_VGND_c_896_n 0.00929484f $X=0.26 $Y=0.49 $X2=0 $Y2=0
cc_497 N_A_27_69#_c_811_n N_VGND_c_896_n 0.00704609f $X=1.12 $Y=0.49 $X2=0 $Y2=0
cc_498 N_A_27_69#_c_813_n N_VGND_c_896_n 0.00704609f $X=1.98 $Y=0.49 $X2=0 $Y2=0
cc_499 N_A_27_69#_c_814_n N_A_454_69#_M1006_s 0.00176461f $X=2.755 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_500 N_A_27_69#_c_815_n N_A_454_69#_M1020_s 0.00261503f $X=3.775 $Y=1.17 $X2=0
+ $Y2=0
cc_501 N_A_27_69#_c_814_n N_A_454_69#_c_997_n 0.017036f $X=2.755 $Y=1.17 $X2=0
+ $Y2=0
cc_502 N_A_27_69#_M1009_d N_A_454_69#_c_990_n 0.00261503f $X=2.7 $Y=0.345 $X2=0
+ $Y2=0
cc_503 N_A_27_69#_c_814_n N_A_454_69#_c_990_n 0.00272017f $X=2.755 $Y=1.17 $X2=0
+ $Y2=0
cc_504 N_A_27_69#_c_843_n N_A_454_69#_c_990_n 0.0203497f $X=2.92 $Y=0.69 $X2=0
+ $Y2=0
cc_505 N_A_27_69#_c_815_n N_A_454_69#_c_990_n 0.00272017f $X=3.775 $Y=1.17 $X2=0
+ $Y2=0
cc_506 N_A_27_69#_c_813_n N_A_454_69#_c_991_n 0.0049425f $X=1.98 $Y=0.49 $X2=0
+ $Y2=0
cc_507 N_A_27_69#_c_815_n N_A_454_69#_c_1004_n 0.0217471f $X=3.775 $Y=1.17 $X2=0
+ $Y2=0
cc_508 N_A_27_69#_M1028_d N_A_454_69#_c_992_n 0.00378299f $X=3.72 $Y=0.345 $X2=0
+ $Y2=0
cc_509 N_A_27_69#_c_815_n N_A_454_69#_c_992_n 0.00272017f $X=3.775 $Y=1.17 $X2=0
+ $Y2=0
cc_510 N_A_27_69#_c_816_n N_A_454_69#_c_992_n 0.0249442f $X=3.94 $Y=0.69 $X2=0
+ $Y2=0
cc_511 N_A_27_69#_c_816_n N_A_454_69#_c_995_n 0.00219337f $X=3.94 $Y=0.69 $X2=0
+ $Y2=0
cc_512 N_VGND_c_889_n N_A_454_69#_c_990_n 0.0435927f $X=6.445 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_c_896_n N_A_454_69#_c_990_n 0.0246836f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_888_n N_A_454_69#_c_991_n 0.00219498f $X=1.55 $Y=0.47 $X2=0
+ $Y2=0
cc_515 N_VGND_c_889_n N_A_454_69#_c_991_n 0.0234284f $X=6.445 $Y=0 $X2=0 $Y2=0
cc_516 N_VGND_c_896_n N_A_454_69#_c_991_n 0.0125908f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_889_n N_A_454_69#_c_992_n 0.0720387f $X=6.445 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_896_n N_A_454_69#_c_992_n 0.0413444f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_889_n N_A_454_69#_c_993_n 0.0565048f $X=6.445 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_890_n N_A_454_69#_c_993_n 9.81589e-19 $X=6.61 $Y=0.45 $X2=0
+ $Y2=0
cc_521 N_VGND_c_896_n N_A_454_69#_c_993_n 0.0315799f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_889_n N_A_454_69#_c_994_n 0.0235159f $X=6.445 $Y=0 $X2=0 $Y2=0
cc_523 N_VGND_c_896_n N_A_454_69#_c_994_n 0.0127052f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_524 N_VGND_c_889_n N_A_454_69#_c_995_n 0.0177478f $X=6.445 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_896_n N_A_454_69#_c_995_n 0.00979598f $X=7.92 $Y=0 $X2=0 $Y2=0
