* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 Y B2 a_76_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_76_69# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR B1 a_159_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_399_367# A2 a_489_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND A2 a_76_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_76_69# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_159_367# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_489_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Y A3 a_399_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_76_69# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
