* File: sky130_fd_sc_lp__einvp_4.pex.spice
* Created: Fri Aug 28 10:33:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVP_4%TE 1 3 6 8 10 12 13 15 17 18 20 22 23 25 27
+ 28 30 31 32 33 34 35 36 37 38 44 45 49
c93 34 0 1.3382e-19 $X=2.235 $Y=1.275
c94 33 0 1.3334e-19 $X=1.805 $Y=1.275
c95 28 0 1.31521e-19 $X=2.875 $Y=1.275
c96 18 0 1.30619e-19 $X=1.73 $Y=1.275
r97 44 47 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=3.04 $Y=1.17
+ $X2=3.04 $Y2=1.275
r98 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.17 $X2=3.04 $Y2=1.17
r99 38 49 0.789345 $w=3.63e-07 $l=2.5e-08 $layer=LI1_cond $X=3.057 $Y=1.295
+ $X2=3.057 $Y2=1.32
r100 38 45 3.94672 $w=3.63e-07 $l=1.25e-07 $layer=LI1_cond $X=3.057 $Y=1.295
+ $X2=3.057 $Y2=1.17
r101 37 49 12.3102 $w=2.18e-07 $l=2.35e-07 $layer=LI1_cond $X=2.64 $Y=1.32
+ $X2=2.875 $Y2=1.32
r102 36 37 25.1442 $w=2.18e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.32
+ $X2=2.64 $Y2=1.32
r103 35 36 25.1442 $w=2.18e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.32
+ $X2=2.16 $Y2=1.32
r104 29 34 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.31 $Y=1.275
+ $X2=2.235 $Y2=1.275
r105 28 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.275
+ $X2=3.04 $Y2=1.275
r106 28 29 219.621 $w=1.8e-07 $l=5.65e-07 $layer=POLY_cond $X=2.875 $Y=1.275
+ $X2=2.31 $Y2=1.275
r107 25 34 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.235 $Y=1.185
+ $X2=2.235 $Y2=1.275
r108 25 27 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.235 $Y=1.185
+ $X2=2.235 $Y2=0.655
r109 24 33 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=1.275
+ $X2=1.805 $Y2=1.275
r110 23 34 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=1.275
+ $X2=2.235 $Y2=1.275
r111 23 24 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=2.16 $Y=1.275
+ $X2=1.88 $Y2=1.275
r112 20 33 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.805 $Y=1.185
+ $X2=1.805 $Y2=1.275
r113 20 22 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.805 $Y=1.185
+ $X2=1.805 $Y2=0.655
r114 19 32 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=1.275
+ $X2=1.375 $Y2=1.275
r115 18 33 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.73 $Y=1.275
+ $X2=1.805 $Y2=1.275
r116 18 19 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=1.73 $Y=1.275
+ $X2=1.45 $Y2=1.275
r117 15 32 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.375 $Y=1.185
+ $X2=1.375 $Y2=1.275
r118 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.375 $Y=1.185
+ $X2=1.375 $Y2=0.655
r119 14 31 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.275
+ $X2=0.945 $Y2=1.275
r120 13 32 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.3 $Y=1.275
+ $X2=1.375 $Y2=1.275
r121 13 14 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=1.3 $Y=1.275
+ $X2=1.02 $Y2=1.275
r122 10 31 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.945 $Y=1.185
+ $X2=0.945 $Y2=1.275
r123 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.945 $Y=1.185
+ $X2=0.945 $Y2=0.655
r124 9 30 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=0.59 $Y=1.275
+ $X2=0.515 $Y2=1.275
r125 8 31 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=0.87 $Y=1.275
+ $X2=0.945 $Y2=1.275
r126 8 9 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=0.87 $Y=1.275
+ $X2=0.59 $Y2=1.275
r127 4 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.515 $Y=1.365
+ $X2=0.515 $Y2=1.275
r128 4 6 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=0.515 $Y=1.365
+ $X2=0.515 $Y2=2.465
r129 1 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.515 $Y=1.185
+ $X2=0.515 $Y2=1.275
r130 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.515 $Y=1.185
+ $X2=0.515 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_4%A_35_47# 1 2 7 8 9 11 12 14 16 17 19 21 22
+ 24 26 28 29 30 33 37 41 45 46 48
c90 8 0 2.99021e-20 $X=1.345 $Y=1.65
r91 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.18
+ $Y=1.74 $X2=1.18 $Y2=1.74
r92 43 45 3.91007 $w=2.78e-07 $l=9.5e-08 $layer=LI1_cond $X=1.205 $Y=1.645
+ $X2=1.205 $Y2=1.74
r93 42 48 2.33382 $w=2.25e-07 $l=1.48e-07 $layer=LI1_cond $X=0.43 $Y=1.532
+ $X2=0.282 $Y2=1.532
r94 41 43 6.92219 $w=2.25e-07 $l=1.88202e-07 $layer=LI1_cond $X=1.065 $Y=1.532
+ $X2=1.205 $Y2=1.645
r95 41 42 32.5245 $w=2.23e-07 $l=6.35e-07 $layer=LI1_cond $X=1.065 $Y=1.532
+ $X2=0.43 $Y2=1.532
r96 37 39 36.3313 $w=2.93e-07 $l=9.3e-07 $layer=LI1_cond $X=0.282 $Y=1.98
+ $X2=0.282 $Y2=2.91
r97 35 48 4.10072 $w=2.95e-07 $l=1.13e-07 $layer=LI1_cond $X=0.282 $Y=1.645
+ $X2=0.282 $Y2=1.532
r98 35 37 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=0.282 $Y=1.645
+ $X2=0.282 $Y2=1.98
r99 31 48 4.10072 $w=2.95e-07 $l=1.12e-07 $layer=LI1_cond $X=0.282 $Y=1.42
+ $X2=0.282 $Y2=1.532
r100 31 33 39.0659 $w=2.93e-07 $l=1e-06 $layer=LI1_cond $X=0.282 $Y=1.42
+ $X2=0.282 $Y2=0.42
r101 27 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.18 $Y=1.725
+ $X2=1.18 $Y2=1.74
r102 24 26 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.135 $Y=1.725
+ $X2=3.135 $Y2=2.465
r103 23 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.78 $Y=1.65
+ $X2=2.705 $Y2=1.65
r104 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.06 $Y=1.65
+ $X2=3.135 $Y2=1.725
r105 22 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.06 $Y=1.65
+ $X2=2.78 $Y2=1.65
r106 19 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.705 $Y=1.725
+ $X2=2.705 $Y2=1.65
r107 19 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.705 $Y=1.725
+ $X2=2.705 $Y2=2.465
r108 18 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.35 $Y=1.65
+ $X2=2.275 $Y2=1.65
r109 17 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.63 $Y=1.65
+ $X2=2.705 $Y2=1.65
r110 17 18 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.63 $Y=1.65
+ $X2=2.35 $Y2=1.65
r111 14 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.275 $Y=1.725
+ $X2=2.275 $Y2=1.65
r112 14 16 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.275 $Y=1.725
+ $X2=2.275 $Y2=2.465
r113 13 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.92 $Y=1.65
+ $X2=1.845 $Y2=1.65
r114 12 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.2 $Y=1.65
+ $X2=2.275 $Y2=1.65
r115 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.2 $Y=1.65
+ $X2=1.92 $Y2=1.65
r116 9 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=1.725
+ $X2=1.845 $Y2=1.65
r117 9 11 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.845 $Y=1.725
+ $X2=1.845 $Y2=2.465
r118 8 27 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.345 $Y=1.65
+ $X2=1.18 $Y2=1.725
r119 7 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.77 $Y=1.65
+ $X2=1.845 $Y2=1.65
r120 7 8 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=1.77 $Y=1.65
+ $X2=1.345 $Y2=1.65
r121 2 39 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.835 $X2=0.3 $Y2=2.91
r122 2 37 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.835 $X2=0.3 $Y2=1.98
r123 1 33 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.175
+ $Y=0.235 $X2=0.3 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_4%A 3 7 11 15 17 18 21 25 29 33 36 38 47
r91 46 48 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.21 $Y=1.51
+ $X2=4.345 $Y2=1.51
r92 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.51 $X2=4.21 $Y2=1.51
r93 44 46 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=3.915 $Y=1.51
+ $X2=4.21 $Y2=1.51
r94 41 44 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.87 $Y=1.51
+ $X2=3.915 $Y2=1.51
r95 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.87
+ $Y=1.51 $X2=3.87 $Y2=1.51
r96 38 47 4.60977 $w=3.23e-07 $l=1.3e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.21 $Y2=1.587
r97 38 42 7.44655 $w=3.23e-07 $l=2.1e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=3.87 $Y2=1.587
r98 35 36 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.855 $Y=1.51
+ $X2=5.285 $Y2=1.51
r99 31 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.675
+ $X2=5.285 $Y2=1.51
r100 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.285 $Y=1.675
+ $X2=5.285 $Y2=2.465
r101 27 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.345
+ $X2=5.285 $Y2=1.51
r102 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.285 $Y=1.345
+ $X2=5.285 $Y2=0.765
r103 23 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.675
+ $X2=4.855 $Y2=1.51
r104 23 25 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.855 $Y=1.675
+ $X2=4.855 $Y2=2.465
r105 19 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.345
+ $X2=4.855 $Y2=1.51
r106 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.855 $Y=1.345
+ $X2=4.855 $Y2=0.765
r107 18 48 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.42 $Y=1.51
+ $X2=4.345 $Y2=1.51
r108 17 35 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.78 $Y=1.51
+ $X2=4.855 $Y2=1.51
r109 17 18 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.78 $Y=1.51
+ $X2=4.42 $Y2=1.51
r110 13 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.675
+ $X2=4.345 $Y2=1.51
r111 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.345 $Y=1.675
+ $X2=4.345 $Y2=2.465
r112 9 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.345
+ $X2=4.345 $Y2=1.51
r113 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.345 $Y=1.345
+ $X2=4.345 $Y2=0.765
r114 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.675
+ $X2=3.915 $Y2=1.51
r115 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.915 $Y=1.675
+ $X2=3.915 $Y2=2.465
r116 1 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.345
+ $X2=3.915 $Y2=1.51
r117 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.915 $Y=1.345
+ $X2=3.915 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_4%VPWR 1 2 3 12 18 24 29 30 32 33 34 36 52 53
+ 56
r70 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r72 50 53 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.52 $Y2=3.33
r73 49 52 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=5.52 $Y2=3.33
r74 49 50 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r76 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r77 44 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 41 56 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.747 $Y2=3.33
r80 41 43 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.68 $Y2=3.33
r81 39 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r82 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r83 36 56 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.747 $Y2=3.33
r84 36 38 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=3.33 $X2=0.24
+ $Y2=3.33
r85 34 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r86 34 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 32 46 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.92 $Y2=3.33
r89 31 49 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=3.12 $Y2=3.33
r90 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=2.92 $Y2=3.33
r91 29 43 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=1.68 $Y2=3.33
r92 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=2.06 $Y2=3.33
r93 28 46 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.06 $Y2=3.33
r95 24 27 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.92 $Y=2.19
+ $X2=2.92 $Y2=2.95
r96 22 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=3.33
r97 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=2.95
r98 18 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.06 $Y=2.18
+ $X2=2.06 $Y2=2.95
r99 16 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=3.245
+ $X2=2.06 $Y2=3.33
r100 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.06 $Y=3.245
+ $X2=2.06 $Y2=2.95
r101 12 15 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=0.747 $Y=1.98
+ $X2=0.747 $Y2=2.95
r102 10 56 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=3.245
+ $X2=0.747 $Y2=3.33
r103 10 15 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.747 $Y=3.245
+ $X2=0.747 $Y2=2.95
r104 3 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.835 $X2=2.92 $Y2=2.95
r105 3 24 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.835 $X2=2.92 $Y2=2.19
r106 2 21 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=2.95
r107 2 18 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=2.18
r108 1 15 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.835 $X2=0.73 $Y2=2.95
r109 1 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.835 $X2=0.73 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_4%A_301_367# 1 2 3 4 5 18 22 23 26 30 33 36 40
+ 42 44 46 48 51
c73 22 0 5.293e-19 $X=2.395 $Y=1.84
r74 44 53 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=2.905
+ $X2=5.53 $Y2=2.99
r75 44 46 39.4818 $w=2.68e-07 $l=9.25e-07 $layer=LI1_cond $X=5.53 $Y=2.905
+ $X2=5.53 $Y2=1.98
r76 43 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=2.99
+ $X2=4.6 $Y2=2.99
r77 42 53 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.395 $Y=2.99
+ $X2=5.53 $Y2=2.99
r78 42 43 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.395 $Y=2.99
+ $X2=4.765 $Y2=2.99
r79 38 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=2.905 $X2=4.6
+ $Y2=2.99
r80 38 40 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.6 $Y=2.905 $X2=4.6
+ $Y2=2.425
r81 37 50 7.27324 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=3.795 $Y=2.99
+ $X2=3.525 $Y2=2.99
r82 36 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=2.99
+ $X2=4.6 $Y2=2.99
r83 36 37 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.435 $Y=2.99
+ $X2=3.795 $Y2=2.99
r84 33 50 2.28973 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=2.905
+ $X2=3.525 $Y2=2.99
r85 33 35 20.4884 $w=5.38e-07 $l=9.25e-07 $layer=LI1_cond $X=3.525 $Y=2.905
+ $X2=3.525 $Y2=1.98
r86 32 35 1.21823 $w=5.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.525 $Y=1.925
+ $X2=3.525 $Y2=1.98
r87 31 48 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.585 $Y=1.84
+ $X2=2.49 $Y2=1.84
r88 30 32 57.0258 $w=5.9e-08 $l=3.09596e-07 $layer=LI1_cond $X=3.255 $Y=1.84
+ $X2=3.525 $Y2=1.925
r89 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.255 $Y=1.84
+ $X2=2.585 $Y2=1.84
r90 26 28 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.49 $Y=1.98
+ $X2=2.49 $Y2=2.91
r91 24 48 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=1.925
+ $X2=2.49 $Y2=1.84
r92 24 26 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=2.49 $Y=1.925
+ $X2=2.49 $Y2=1.98
r93 22 48 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.395 $Y=1.84
+ $X2=2.49 $Y2=1.84
r94 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.395 $Y=1.84
+ $X2=1.725 $Y2=1.84
r95 18 20 49.1169 $w=2.08e-07 $l=9.3e-07 $layer=LI1_cond $X=1.62 $Y=1.98
+ $X2=1.62 $Y2=2.91
r96 16 23 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.62 $Y=1.925
+ $X2=1.725 $Y2=1.84
r97 16 18 2.90476 $w=2.08e-07 $l=5.5e-08 $layer=LI1_cond $X=1.62 $Y=1.925
+ $X2=1.62 $Y2=1.98
r98 5 53 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.36
+ $Y=1.835 $X2=5.5 $Y2=2.91
r99 5 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.36
+ $Y=1.835 $X2=5.5 $Y2=1.98
r100 4 40 300 $w=1.7e-07 $l=6.74018e-07 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=1.835 $X2=4.6 $Y2=2.425
r101 3 50 200 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=3 $X=3.21
+ $Y=1.835 $X2=3.35 $Y2=2.91
r102 3 35 200 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=3 $X=3.21
+ $Y=1.835 $X2=3.35 $Y2=1.98
r103 2 28 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.835 $X2=2.49 $Y2=2.91
r104 2 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.835 $X2=2.49 $Y2=1.98
r105 1 20 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.835 $X2=1.63 $Y2=2.91
r106 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.835 $X2=1.63 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_4%Z 1 2 3 4 5 18 20 21 22 26 28 29 32 36 41 42
+ 43 47
r69 42 47 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=2.005
+ $X2=4.115 $Y2=2.09
r70 42 43 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=4.115 $Y=2.095
+ $X2=4.115 $Y2=2.405
r71 42 47 0.192074 $w=2.98e-07 $l=5e-09 $layer=LI1_cond $X=4.115 $Y=2.095
+ $X2=4.115 $Y2=2.09
r72 34 36 34.3812 $w=2.98e-07 $l=8.95e-07 $layer=LI1_cond $X=5.515 $Y=1.385
+ $X2=5.515 $Y2=0.49
r73 30 41 2.01947 $w=4.85e-07 $l=2.33666e-07 $layer=LI1_cond $X=5.08 $Y=2.09
+ $X2=4.885 $Y2=2.005
r74 30 32 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=5.08 $Y=2.09 $X2=5.08
+ $Y2=2.095
r75 29 41 2.01947 $w=4.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=1.92
+ $X2=4.885 $Y2=2.005
r76 28 34 33.1293 $w=2.32e-07 $l=6.3e-07 $layer=LI1_cond $X=4.885 $Y=1.385
+ $X2=5.515 $Y2=1.385
r77 28 29 6.42013 $w=6.78e-07 $l=3.65e-07 $layer=LI1_cond $X=4.885 $Y=1.555
+ $X2=4.885 $Y2=1.92
r78 24 28 13.4095 $w=2.32e-07 $l=2.55e-07 $layer=LI1_cond $X=4.63 $Y=1.385
+ $X2=4.885 $Y2=1.385
r79 24 26 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=4.63 $Y=1.085
+ $X2=4.63 $Y2=0.7
r80 23 42 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.265 $Y=2.005
+ $X2=4.115 $Y2=2.005
r81 22 41 5.28247 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=4.545 $Y=2.005
+ $X2=4.885 $Y2=2.005
r82 22 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.545 $Y=2.005
+ $X2=4.265 $Y2=2.005
r83 20 24 9.57122 $w=2.32e-07 $l=2.85832e-07 $layer=LI1_cond $X=4.465 $Y=1.17
+ $X2=4.63 $Y2=1.385
r84 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.465 $Y=1.17
+ $X2=3.785 $Y2=1.17
r85 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.62 $Y=1.085
+ $X2=3.785 $Y2=1.17
r86 16 18 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.62 $Y=1.085
+ $X2=3.62 $Y2=0.7
r87 5 32 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=4.93
+ $Y=1.835 $X2=5.07 $Y2=2.095
r88 4 42 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=1.835 $X2=4.13 $Y2=2.095
r89 3 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.345 $X2=5.5 $Y2=0.49
r90 2 26 91 $w=1.7e-07 $l=4.47856e-07 $layer=licon1_NDIFF $count=2 $X=4.42
+ $Y=0.345 $X2=4.63 $Y2=0.7
r91 1 18 91 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_NDIFF $count=2 $X=3.495
+ $Y=0.345 $X2=3.62 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_4%VGND 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r68 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 46 47 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r70 43 46 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.52
+ $Y2=0
r71 43 44 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r72 41 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r73 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r74 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r75 38 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r76 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r77 35 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=0.73
+ $Y2=0
r78 35 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=1.2
+ $Y2=0
r79 33 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r80 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r81 30 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.73
+ $Y2=0
r82 30 32 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.24
+ $Y2=0
r83 28 47 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=5.52
+ $Y2=0
r84 28 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r85 26 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.16
+ $Y2=0
r86 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.45
+ $Y2=0
r87 25 43 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.64
+ $Y2=0
r88 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.45
+ $Y2=0
r89 23 37 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.2
+ $Y2=0
r90 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.59
+ $Y2=0
r91 22 40 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.755 $Y=0 $X2=2.16
+ $Y2=0
r92 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.59
+ $Y2=0
r93 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0
r94 18 20 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0.44
r95 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0
r96 14 16 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0.58
r97 10 50 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r98 10 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r99 3 20 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.235 $X2=2.45 $Y2=0.44
r100 2 16 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.59 $Y2=0.58
r101 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_4%A_204_47# 1 2 3 4 15 17 18 21 23 26 27 28 31
+ 33 37 40 42
c75 17 0 2.99021e-20 $X=1.925 $Y=0.955
r76 35 37 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=5.08 $Y=0.435
+ $X2=5.08 $Y2=0.47
r77 34 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=0.35
+ $X2=4.13 $Y2=0.35
r78 33 35 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.965 $Y=0.35
+ $X2=5.08 $Y2=0.435
r79 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.965 $Y=0.35
+ $X2=4.295 $Y2=0.35
r80 29 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.435
+ $X2=4.13 $Y2=0.35
r81 29 31 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=4.13 $Y=0.435
+ $X2=4.13 $Y2=0.47
r82 27 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=0.35
+ $X2=4.13 $Y2=0.35
r83 27 28 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.965 $Y=0.35
+ $X2=3.19 $Y2=0.35
r84 25 28 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=3.015 $Y=0.435
+ $X2=3.19 $Y2=0.35
r85 25 26 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=3.015 $Y=0.435
+ $X2=3.015 $Y2=0.725
r86 24 40 4.19778 $w=2.42e-07 $l=9.5e-08 $layer=LI1_cond $X=2.115 $Y=0.882
+ $X2=2.02 $Y2=0.882
r87 23 26 19.5729 $w=3.15e-07 $l=4.67e-07 $layer=LI1_cond $X=2.548 $Y=0.882
+ $X2=3.015 $Y2=0.882
r88 23 24 15.8415 $w=3.13e-07 $l=4.33e-07 $layer=LI1_cond $X=2.548 $Y=0.882
+ $X2=2.115 $Y2=0.882
r89 19 40 2.23415 $w=1.9e-07 $l=1.57e-07 $layer=LI1_cond $X=2.02 $Y=0.725
+ $X2=2.02 $Y2=0.882
r90 19 21 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=2.02 $Y=0.725
+ $X2=2.02 $Y2=0.42
r91 17 40 4.19778 $w=2.42e-07 $l=1.26333e-07 $layer=LI1_cond $X=1.925 $Y=0.955
+ $X2=2.02 $Y2=0.882
r92 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.925 $Y=0.955
+ $X2=1.255 $Y2=0.955
r93 13 18 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.142 $Y=0.87
+ $X2=1.255 $Y2=0.955
r94 13 15 23.0489 $w=2.23e-07 $l=4.5e-07 $layer=LI1_cond $X=1.142 $Y=0.87
+ $X2=1.142 $Y2=0.42
r95 4 37 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.93
+ $Y=0.345 $X2=5.07 $Y2=0.47
r96 3 31 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.99
+ $Y=0.345 $X2=4.13 $Y2=0.47
r97 2 40 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.235 $X2=2.02 $Y2=0.875
r98 2 21 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.235 $X2=2.02 $Y2=0.42
r99 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.02
+ $Y=0.235 $X2=1.16 $Y2=0.42
.ends

