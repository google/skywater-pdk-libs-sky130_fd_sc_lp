# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__or2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__or2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.425000 2.275000 1.760000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.295000 0.545000 2.130000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.570000 0.255000 2.830000 0.735000 ;
        RECT 2.570000 0.735000 3.690000 0.905000 ;
        RECT 2.580000 1.755000 4.235000 1.945000 ;
        RECT 2.580000 1.945000 2.830000 3.075000 ;
        RECT 2.960000 0.905000 3.690000 1.065000 ;
        RECT 2.960000 1.065000 4.235000 1.245000 ;
        RECT 3.500000 0.255000 3.690000 0.735000 ;
        RECT 3.500000 1.945000 3.690000 3.075000 ;
        RECT 3.965000 1.245000 4.235000 1.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 4.320000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 4.510000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.095000  2.300000 1.045000 2.470000 ;
      RECT 0.095000  2.470000 0.355000 2.915000 ;
      RECT 0.525000  2.640000 0.855000 3.245000 ;
      RECT 0.715000  0.255000 1.045000 2.300000 ;
      RECT 1.240000  0.085000 1.570000 0.905000 ;
      RECT 1.240000  1.075000 2.790000 1.255000 ;
      RECT 1.240000  1.255000 1.415000 1.930000 ;
      RECT 1.240000  1.930000 1.570000 3.075000 ;
      RECT 1.740000  0.255000 1.965000 1.075000 ;
      RECT 2.080000  1.930000 2.410000 3.245000 ;
      RECT 2.135000  0.085000 2.400000 0.905000 ;
      RECT 2.445000  1.255000 2.790000 1.415000 ;
      RECT 2.445000  1.415000 3.795000 1.585000 ;
      RECT 3.000000  0.085000 3.330000 0.565000 ;
      RECT 3.000000  2.115000 3.330000 3.245000 ;
      RECT 3.860000  0.085000 4.190000 0.895000 ;
      RECT 3.860000  2.115000 4.190000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__or2b_4
END LIBRARY
