* File: sky130_fd_sc_lp__decap_12.pex.spice
* Created: Fri Aug 28 10:19:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAP_12%VGND 1 7 9 15 18 23 28 32 36 46 47 50 53
c29 23 0 8.49014e-20 $X=2.415 $Y=1.77
r30 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r31 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r32 47 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r33 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r34 44 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.095
+ $Y2=0
r35 44 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.52
+ $Y2=0
r36 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r37 42 43 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r38 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r39 39 42 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r40 39 40 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r42 37 39 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r43 36 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=5.095
+ $Y2=0
r44 36 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=4.56
+ $Y2=0
r45 32 43 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.56
+ $Y2=0
r46 32 40 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.2
+ $Y2=0
r47 28 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=0.36
+ $X2=5.095 $Y2=1.04
r48 26 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0.085
+ $X2=5.095 $Y2=0
r49 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.095 $Y=0.085
+ $X2=5.095 $Y2=0.36
r50 23 24 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.415
+ $Y=1.77 $X2=2.415 $Y2=1.77
r51 21 24 40.8678 $w=1.604e-06 $l=1.36e-06 $layer=POLY_cond $X=1.055 $Y=2.415
+ $X2=2.415 $Y2=2.415
r52 20 23 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=1.055 $Y=1.77
+ $X2=2.415 $Y2=1.77
r53 20 21 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.055
+ $Y=1.77 $X2=1.055 $Y2=1.77
r54 18 20 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=0.98 $Y=1.77
+ $X2=1.055 $Y2=1.77
r55 15 17 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.815 $Y=0.38
+ $X2=0.815 $Y2=1.06
r56 13 18 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=0.815 $Y=1.605
+ $X2=0.98 $Y2=1.77
r57 13 17 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.815 $Y=1.605
+ $X2=0.815 $Y2=1.06
r58 12 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r59 12 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.38
r60 7 24 6.40574 $w=1.604e-06 $l=2.24332e-07 $layer=POLY_cond $X=2.58 $Y=2.555
+ $X2=2.415 $Y2=2.415
r61 7 9 11.1507 $w=1.34e-06 $l=3.1e-07 $layer=POLY_cond $X=2.58 $Y=2.555
+ $X2=2.89 $Y2=2.555
r62 1 30 121.333 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.095 $Y2=1.04
r63 1 28 121.333 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.095 $Y2=0.36
r64 1 17 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=0.815 $Y2=1.06
r65 1 15 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=0.815 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DECAP_12%VPWR 1 11 15 22 26 29 32 37 42 52 53 56 59
c30 22 0 8.49014e-20 $X=4.79 $Y=1.51
r31 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r32 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 53 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r34 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r35 50 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.195 $Y=3.33
+ $X2=5.03 $Y2=3.33
r36 50 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.195 $Y=3.33
+ $X2=5.52 $Y2=3.33
r37 49 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r38 48 49 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r39 46 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 45 48 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r41 45 46 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 43 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r43 43 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 42 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=5.03 $Y2=3.33
r45 42 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=4.56 $Y2=3.33
r46 40 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 37 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r49 37 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 29 49 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 29 46 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 26 28 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.03 $Y=2.29
+ $X2=5.03 $Y2=2.97
r53 24 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=3.245
+ $X2=5.03 $Y2=3.33
r54 24 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.03 $Y=3.245
+ $X2=5.03 $Y2=2.97
r55 23 26 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=5.03 $Y=1.675
+ $X2=5.03 $Y2=2.29
r56 21 22 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=4.79
+ $Y=1.51 $X2=4.79 $Y2=1.51
r57 18 22 53.4994 $w=1.57e-06 $l=1.7e-06 $layer=POLY_cond $X=3.09 $Y=0.89
+ $X2=4.79 $Y2=0.89
r58 18 32 4.24848 $w=1.57e-06 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=0.89
+ $X2=2.955 $Y2=0.89
r59 17 21 58.4822 $w=3.33e-07 $l=1.7e-06 $layer=LI1_cond $X=3.09 $Y=1.507
+ $X2=4.79 $Y2=1.507
r60 17 18 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.09
+ $Y=1.51 $X2=3.09 $Y2=1.51
r61 15 23 6.81699 $w=3.35e-07 $l=2.36525e-07 $layer=LI1_cond $X=4.865 $Y=1.507
+ $X2=5.03 $Y2=1.675
r62 15 21 2.5801 $w=3.33e-07 $l=7.5e-08 $layer=LI1_cond $X=4.865 $Y=1.507
+ $X2=4.79 $Y2=1.507
r63 11 14 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.74 $Y=2.27
+ $X2=0.74 $Y2=2.95
r64 9 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245 $X2=0.74
+ $Y2=3.33
r65 9 14 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=2.95
r66 1 28 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.095 $X2=5.03 $Y2=2.97
r67 1 26 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.095 $X2=5.03 $Y2=2.29
r68 1 14 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.095 $X2=0.74 $Y2=2.95
r69 1 11 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.095 $X2=0.74 $Y2=2.27
.ends

