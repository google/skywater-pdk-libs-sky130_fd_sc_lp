* File: sky130_fd_sc_lp__and3b_m.pxi.spice
* Created: Wed Sep  2 09:32:32 2020
* 
x_PM_SKY130_FD_SC_LP__AND3B_M%A_N N_A_N_c_69_n N_A_N_M1006_g N_A_N_M1008_g
+ N_A_N_c_72_n A_N A_N A_N A_N A_N N_A_N_c_74_n PM_SKY130_FD_SC_LP__AND3B_M%A_N
x_PM_SKY130_FD_SC_LP__AND3B_M%A_110_53# N_A_110_53#_M1006_d N_A_110_53#_M1008_d
+ N_A_110_53#_c_98_n N_A_110_53#_c_99_n N_A_110_53#_c_107_n N_A_110_53#_c_108_n
+ N_A_110_53#_M1004_g N_A_110_53#_M1002_g N_A_110_53#_c_101_n
+ N_A_110_53#_c_102_n N_A_110_53#_c_103_n N_A_110_53#_c_104_n
+ N_A_110_53#_c_105_n PM_SKY130_FD_SC_LP__AND3B_M%A_110_53#
x_PM_SKY130_FD_SC_LP__AND3B_M%B N_B_M1003_g N_B_M1000_g N_B_c_155_n N_B_c_156_n
+ N_B_c_157_n B B B N_B_c_159_n PM_SKY130_FD_SC_LP__AND3B_M%B
x_PM_SKY130_FD_SC_LP__AND3B_M%C N_C_M1007_g N_C_M1005_g N_C_c_199_n N_C_c_204_n
+ C C C N_C_c_201_n PM_SKY130_FD_SC_LP__AND3B_M%C
x_PM_SKY130_FD_SC_LP__AND3B_M%A_220_53# N_A_220_53#_M1002_s N_A_220_53#_M1004_s
+ N_A_220_53#_M1000_d N_A_220_53#_c_244_n N_A_220_53#_c_240_n
+ N_A_220_53#_M1009_g N_A_220_53#_M1001_g N_A_220_53#_c_242_n
+ N_A_220_53#_c_247_n N_A_220_53#_c_248_n N_A_220_53#_c_243_n
+ N_A_220_53#_c_249_n N_A_220_53#_c_250_n N_A_220_53#_c_251_n
+ PM_SKY130_FD_SC_LP__AND3B_M%A_220_53#
x_PM_SKY130_FD_SC_LP__AND3B_M%VPWR N_VPWR_M1008_s N_VPWR_M1004_d N_VPWR_M1007_d
+ N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n
+ N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n VPWR N_VPWR_c_320_n
+ N_VPWR_c_311_n PM_SKY130_FD_SC_LP__AND3B_M%VPWR
x_PM_SKY130_FD_SC_LP__AND3B_M%X N_X_M1009_d N_X_M1001_d X X X X X X N_X_c_357_n
+ PM_SKY130_FD_SC_LP__AND3B_M%X
x_PM_SKY130_FD_SC_LP__AND3B_M%VGND N_VGND_M1006_s N_VGND_M1005_d N_VGND_c_369_n
+ N_VGND_c_370_n N_VGND_c_371_n VGND N_VGND_c_372_n N_VGND_c_373_n
+ N_VGND_c_374_n N_VGND_c_375_n PM_SKY130_FD_SC_LP__AND3B_M%VGND
cc_1 VNB N_A_N_c_69_n 0.0263701f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.288
cc_2 VNB N_A_N_M1006_g 0.0287688f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.475
cc_3 VNB N_A_N_M1008_g 0.00870147f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_4 VNB N_A_N_c_72_n 0.0373858f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_5 VNB A_N 0.00807475f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A_N_c_74_n 0.035729f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_7 VNB N_A_110_53#_c_98_n 0.00932936f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_8 VNB N_A_110_53#_c_99_n 0.0166631f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_9 VNB N_A_110_53#_M1002_g 0.0428678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_110_53#_c_101_n 0.0121271f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.005
cc_11 VNB N_A_110_53#_c_102_n 0.00223773f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=0.84
cc_12 VNB N_A_110_53#_c_103_n 0.00301901f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.295
cc_13 VNB N_A_110_53#_c_104_n 0.0169816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_110_53#_c_105_n 0.042053f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=2.035
cc_15 VNB N_B_M1000_g 0.0121375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_155_n 0.0157952f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_17 VNB N_B_c_156_n 0.0209027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_157_n 0.015314f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_19 VNB B 0.0089247f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_20 VNB N_B_c_159_n 0.016411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C_M1005_g 0.0364232f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_22 VNB N_C_c_199_n 0.0196891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB C 0.00744437f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_C_c_201_n 0.0153418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_220_53#_c_240_n 0.0523074f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_26 VNB N_A_220_53#_M1001_g 0.0345064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_220_53#_c_242_n 0.00841734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_220_53#_c_243_n 0.00283144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_311_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_357_n 0.0559937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_369_n 0.011158f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_32 VNB N_VGND_c_370_n 0.00633646f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_33 VNB N_VGND_c_371_n 0.00126149f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_VGND_c_372_n 0.057317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_373_n 0.0188381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_374_n 0.217651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_375_n 0.00473063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_N_M1008_g 0.0705536f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_39 VPB A_N 0.0423578f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_40 VPB N_A_110_53#_c_98_n 0.00198452f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_41 VPB N_A_110_53#_c_107_n 0.0204574f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.51
cc_42 VPB N_A_110_53#_c_108_n 0.0143353f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_43 VPB N_A_110_53#_M1004_g 0.0235094f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_44 VPB N_A_110_53#_c_103_n 0.0250757f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_45 VPB N_B_M1000_g 0.0304564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_C_M1007_g 0.0200301f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.84
cc_47 VPB N_C_c_199_n 0.00325954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_C_c_204_n 0.0193282f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.51
cc_49 VPB C 0.00926806f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_50 VPB N_A_220_53#_c_244_n 0.0570485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_220_53#_M1001_g 0.0667828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_220_53#_c_242_n 0.00113048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_220_53#_c_247_n 0.0183181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_220_53#_c_248_n 0.00825751f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_55 VPB N_A_220_53#_c_249_n 0.00267484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_220_53#_c_250_n 0.00243789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_220_53#_c_251_n 0.045536f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_312_n 0.010774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_313_n 0.0104735f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_60 VPB N_VPWR_c_314_n 0.0341982f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_61 VPB N_VPWR_c_315_n 0.0155838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_316_n 0.0372285f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_63 VPB N_VPWR_c_317_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_64 VPB N_VPWR_c_318_n 0.0200954f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_65 VPB N_VPWR_c_319_n 0.00370272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_320_n 0.022889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_311_n 0.0894711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_X_c_357_n 0.0401679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 N_A_N_c_72_n N_A_110_53#_c_98_n 0.00420397f $X=0.327 $Y=1.51 $X2=0 $Y2=0
cc_70 N_A_N_M1008_g N_A_110_53#_c_108_n 0.00420397f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_71 N_A_N_c_69_n N_A_110_53#_c_101_n 0.017642f $X=0.327 $Y=1.288 $X2=0 $Y2=0
cc_72 N_A_N_M1006_g N_A_110_53#_c_102_n 0.0118863f $X=0.475 $Y=0.475 $X2=0 $Y2=0
cc_73 N_A_N_c_72_n N_A_110_53#_c_103_n 0.0118863f $X=0.327 $Y=1.51 $X2=0 $Y2=0
cc_74 A_N N_A_110_53#_c_104_n 0.10308f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_75 N_A_N_c_74_n N_A_110_53#_c_104_n 0.0118863f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_76 N_A_N_M1006_g N_A_110_53#_c_105_n 0.017642f $X=0.475 $Y=0.475 $X2=0 $Y2=0
cc_77 A_N N_A_110_53#_c_105_n 4.39952e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_78 N_A_N_M1008_g N_VPWR_c_313_n 0.00463498f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_79 A_N N_VPWR_c_313_n 0.0160484f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 N_A_N_M1008_g N_VPWR_c_316_n 0.00478016f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_81 N_A_N_M1008_g N_VPWR_c_311_n 0.00983495f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_82 A_N N_VPWR_c_311_n 0.00109783f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_83 N_A_N_M1006_g N_VGND_c_370_n 0.00462473f $X=0.475 $Y=0.475 $X2=0 $Y2=0
cc_84 A_N N_VGND_c_370_n 0.0110529f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_85 N_A_N_c_74_n N_VGND_c_370_n 0.00141621f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_86 N_A_N_M1006_g N_VGND_c_372_n 0.00555245f $X=0.475 $Y=0.475 $X2=0 $Y2=0
cc_87 N_A_N_M1006_g N_VGND_c_374_n 0.012364f $X=0.475 $Y=0.475 $X2=0 $Y2=0
cc_88 A_N N_VGND_c_374_n 8.0298e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_A_N_c_74_n N_VGND_c_374_n 0.00220006f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_90 N_A_110_53#_c_98_n N_B_M1000_g 5.87802e-19 $X=1.045 $Y=1.705 $X2=0 $Y2=0
cc_91 N_A_110_53#_c_107_n N_B_M1000_g 0.0219326f $X=1.365 $Y=1.78 $X2=0 $Y2=0
cc_92 N_A_110_53#_M1002_g N_B_c_155_n 0.0406107f $X=1.445 $Y=0.475 $X2=0 $Y2=0
cc_93 N_A_110_53#_c_99_n N_B_c_156_n 0.0406107f $X=1.37 $Y=1.39 $X2=0 $Y2=0
cc_94 N_A_110_53#_M1002_g B 0.00711189f $X=1.445 $Y=0.475 $X2=0 $Y2=0
cc_95 N_A_110_53#_c_98_n N_A_220_53#_c_242_n 8.14977e-19 $X=1.045 $Y=1.705 $X2=0
+ $Y2=0
cc_96 N_A_110_53#_c_99_n N_A_220_53#_c_242_n 0.00886747f $X=1.37 $Y=1.39 $X2=0
+ $Y2=0
cc_97 N_A_110_53#_c_107_n N_A_220_53#_c_242_n 0.00500935f $X=1.365 $Y=1.78 $X2=0
+ $Y2=0
cc_98 N_A_110_53#_M1002_g N_A_220_53#_c_242_n 0.0128052f $X=1.445 $Y=0.475 $X2=0
+ $Y2=0
cc_99 N_A_110_53#_c_102_n N_A_220_53#_c_242_n 0.00707862f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_100 N_A_110_53#_c_103_n N_A_220_53#_c_242_n 0.0122553f $X=0.69 $Y=2.835 $X2=0
+ $Y2=0
cc_101 N_A_110_53#_c_104_n N_A_220_53#_c_242_n 0.0488333f $X=0.955 $Y=0.96 $X2=0
+ $Y2=0
cc_102 N_A_110_53#_c_105_n N_A_220_53#_c_242_n 0.003541f $X=0.955 $Y=0.96 $X2=0
+ $Y2=0
cc_103 N_A_110_53#_c_99_n N_A_220_53#_c_247_n 9.94864e-19 $X=1.37 $Y=1.39 $X2=0
+ $Y2=0
cc_104 N_A_110_53#_c_107_n N_A_220_53#_c_247_n 0.00352914f $X=1.365 $Y=1.78
+ $X2=0 $Y2=0
cc_105 N_A_110_53#_M1004_g N_A_220_53#_c_247_n 0.00733543f $X=1.44 $Y=2.225
+ $X2=0 $Y2=0
cc_106 N_A_110_53#_M1002_g N_A_220_53#_c_243_n 0.00292658f $X=1.445 $Y=0.475
+ $X2=0 $Y2=0
cc_107 N_A_110_53#_c_102_n N_A_220_53#_c_243_n 0.0120203f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_108 N_A_110_53#_c_105_n N_A_220_53#_c_243_n 0.00251502f $X=0.955 $Y=0.96
+ $X2=0 $Y2=0
cc_109 N_A_110_53#_c_107_n N_A_220_53#_c_249_n 0.00992614f $X=1.365 $Y=1.78
+ $X2=0 $Y2=0
cc_110 N_A_110_53#_M1004_g N_A_220_53#_c_249_n 0.00958555f $X=1.44 $Y=2.225
+ $X2=0 $Y2=0
cc_111 N_A_110_53#_c_103_n N_A_220_53#_c_249_n 0.0261169f $X=0.69 $Y=2.835 $X2=0
+ $Y2=0
cc_112 N_A_110_53#_c_103_n N_VPWR_c_313_n 0.00115095f $X=0.69 $Y=2.835 $X2=0
+ $Y2=0
cc_113 N_A_110_53#_M1004_g N_VPWR_c_314_n 0.00314874f $X=1.44 $Y=2.225 $X2=0
+ $Y2=0
cc_114 N_A_110_53#_M1004_g N_VPWR_c_316_n 0.00297774f $X=1.44 $Y=2.225 $X2=0
+ $Y2=0
cc_115 N_A_110_53#_c_103_n N_VPWR_c_316_n 0.0100892f $X=0.69 $Y=2.835 $X2=0
+ $Y2=0
cc_116 N_A_110_53#_M1004_g N_VPWR_c_311_n 0.00400849f $X=1.44 $Y=2.225 $X2=0
+ $Y2=0
cc_117 N_A_110_53#_c_103_n N_VPWR_c_311_n 0.00777327f $X=0.69 $Y=2.835 $X2=0
+ $Y2=0
cc_118 N_A_110_53#_M1002_g N_VGND_c_372_n 0.00529939f $X=1.445 $Y=0.475 $X2=0
+ $Y2=0
cc_119 N_A_110_53#_c_102_n N_VGND_c_372_n 0.00935935f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_120 N_A_110_53#_M1002_g N_VGND_c_374_n 0.0108838f $X=1.445 $Y=0.475 $X2=0
+ $Y2=0
cc_121 N_A_110_53#_c_102_n N_VGND_c_374_n 0.00777327f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_122 N_A_110_53#_c_104_n N_VGND_c_374_n 0.00903386f $X=0.955 $Y=0.96 $X2=0
+ $Y2=0
cc_123 N_A_110_53#_c_105_n N_VGND_c_374_n 5.6385e-19 $X=0.955 $Y=0.96 $X2=0
+ $Y2=0
cc_124 N_B_c_155_n N_C_M1005_g 0.0196294f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_125 B N_C_M1005_g 0.00865286f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_126 N_B_c_159_n N_C_M1005_g 0.0135986f $X=1.895 $Y=0.96 $X2=0 $Y2=0
cc_127 N_B_M1000_g N_C_c_199_n 0.00993385f $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_128 N_B_c_157_n N_C_c_199_n 0.0135986f $X=1.895 $Y=1.465 $X2=0 $Y2=0
cc_129 N_B_M1000_g N_C_c_204_n 0.0202192f $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_130 N_B_M1000_g C 0.00164048f $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_131 B C 0.0255719f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_132 N_B_c_159_n C 0.00202014f $X=1.895 $Y=0.96 $X2=0 $Y2=0
cc_133 N_B_c_156_n N_C_c_201_n 0.0135986f $X=1.895 $Y=1.3 $X2=0 $Y2=0
cc_134 N_B_M1000_g N_A_220_53#_c_242_n 0.00622295f $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_135 N_B_c_155_n N_A_220_53#_c_242_n 6.97492e-19 $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_136 B N_A_220_53#_c_242_n 0.0563916f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_137 N_B_M1000_g N_A_220_53#_c_247_n 0.0150853f $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_138 N_B_c_157_n N_A_220_53#_c_247_n 0.00391456f $X=1.895 $Y=1.465 $X2=0 $Y2=0
cc_139 B N_A_220_53#_c_247_n 0.0195355f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_140 N_B_M1000_g N_A_220_53#_c_248_n 0.00229433f $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_141 N_B_c_155_n N_A_220_53#_c_243_n 4.36821e-19 $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_142 B N_A_220_53#_c_243_n 0.00983632f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_143 N_B_M1000_g N_A_220_53#_c_249_n 5.39506e-19 $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_144 N_B_M1000_g N_VPWR_c_314_n 0.00105495f $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_145 N_B_M1000_g N_VPWR_c_318_n 0.00297774f $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_146 N_B_M1000_g N_VPWR_c_311_n 0.00400849f $X=1.87 $Y=2.225 $X2=0 $Y2=0
cc_147 N_B_c_155_n N_VGND_c_371_n 0.0018163f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_148 B N_VGND_c_371_n 0.00177802f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_149 N_B_c_155_n N_VGND_c_372_n 0.0037597f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_150 B N_VGND_c_372_n 0.00931852f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_151 N_B_c_155_n N_VGND_c_374_n 0.00542249f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_152 B N_VGND_c_374_n 0.0123305f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_153 N_B_c_159_n N_VGND_c_374_n 0.00210244f $X=1.895 $Y=0.96 $X2=0 $Y2=0
cc_154 B A_304_53# 0.00304451f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_155 B A_376_53# 0.00359473f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_156 N_C_M1007_g N_A_220_53#_c_244_n 0.00242712f $X=2.3 $Y=2.225 $X2=0 $Y2=0
cc_157 N_C_M1005_g N_A_220_53#_c_240_n 0.0276284f $X=2.345 $Y=0.475 $X2=0 $Y2=0
cc_158 C N_A_220_53#_c_240_n 0.0104433f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_159 N_C_M1007_g N_A_220_53#_M1001_g 0.014605f $X=2.3 $Y=2.225 $X2=0 $Y2=0
cc_160 N_C_c_201_n N_A_220_53#_M1001_g 0.039179f $X=2.435 $Y=1.35 $X2=0 $Y2=0
cc_161 N_C_c_204_n N_A_220_53#_c_247_n 0.00358497f $X=2.412 $Y=1.855 $X2=0 $Y2=0
cc_162 C N_A_220_53#_c_247_n 0.00651816f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_163 N_C_M1007_g N_A_220_53#_c_248_n 0.00319558f $X=2.3 $Y=2.225 $X2=0 $Y2=0
cc_164 N_C_M1007_g N_A_220_53#_c_250_n 5.48582e-19 $X=2.3 $Y=2.225 $X2=0 $Y2=0
cc_165 N_C_M1007_g N_A_220_53#_c_251_n 0.00615808f $X=2.3 $Y=2.225 $X2=0 $Y2=0
cc_166 N_C_M1007_g N_VPWR_c_315_n 0.0043911f $X=2.3 $Y=2.225 $X2=0 $Y2=0
cc_167 N_C_c_204_n N_VPWR_c_315_n 8.08513e-19 $X=2.412 $Y=1.855 $X2=0 $Y2=0
cc_168 C N_VPWR_c_315_n 0.0131759f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_169 N_C_M1007_g N_VPWR_c_311_n 3.65623e-19 $X=2.3 $Y=2.225 $X2=0 $Y2=0
cc_170 N_C_M1007_g N_X_c_357_n 0.00137009f $X=2.3 $Y=2.225 $X2=0 $Y2=0
cc_171 N_C_M1005_g N_X_c_357_n 4.31092e-19 $X=2.345 $Y=0.475 $X2=0 $Y2=0
cc_172 C N_X_c_357_n 0.0777429f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_173 N_C_c_201_n N_X_c_357_n 5.70331e-19 $X=2.435 $Y=1.35 $X2=0 $Y2=0
cc_174 N_C_M1005_g N_VGND_c_371_n 0.00998825f $X=2.345 $Y=0.475 $X2=0 $Y2=0
cc_175 C N_VGND_c_371_n 0.0132661f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_176 N_C_c_201_n N_VGND_c_371_n 5.75172e-19 $X=2.435 $Y=1.35 $X2=0 $Y2=0
cc_177 N_C_M1005_g N_VGND_c_372_n 0.00461019f $X=2.345 $Y=0.475 $X2=0 $Y2=0
cc_178 N_C_M1005_g N_VGND_c_374_n 0.00709328f $X=2.345 $Y=0.475 $X2=0 $Y2=0
cc_179 C N_VGND_c_374_n 0.00309169f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_180 N_A_220_53#_c_247_n N_VPWR_c_314_n 0.0139641f $X=1.98 $Y=1.86 $X2=0 $Y2=0
cc_181 N_A_220_53#_c_248_n N_VPWR_c_314_n 0.0264675f $X=2.085 $Y=2.16 $X2=0
+ $Y2=0
cc_182 N_A_220_53#_c_250_n N_VPWR_c_314_n 0.0105383f $X=2.145 $Y=2.94 $X2=0
+ $Y2=0
cc_183 N_A_220_53#_c_251_n N_VPWR_c_314_n 0.00588044f $X=2.145 $Y=2.94 $X2=0
+ $Y2=0
cc_184 N_A_220_53#_c_244_n N_VPWR_c_315_n 0.0219214f $X=2.81 $Y=3.03 $X2=0 $Y2=0
cc_185 N_A_220_53#_M1001_g N_VPWR_c_315_n 0.0174692f $X=2.885 $Y=2.225 $X2=0
+ $Y2=0
cc_186 N_A_220_53#_c_248_n N_VPWR_c_315_n 0.0278483f $X=2.085 $Y=2.16 $X2=0
+ $Y2=0
cc_187 N_A_220_53#_c_250_n N_VPWR_c_315_n 0.0120815f $X=2.145 $Y=2.94 $X2=0
+ $Y2=0
cc_188 N_A_220_53#_c_251_n N_VPWR_c_315_n 0.00124514f $X=2.145 $Y=2.94 $X2=0
+ $Y2=0
cc_189 N_A_220_53#_c_250_n N_VPWR_c_318_n 0.0152941f $X=2.145 $Y=2.94 $X2=0
+ $Y2=0
cc_190 N_A_220_53#_c_251_n N_VPWR_c_318_n 0.0110537f $X=2.145 $Y=2.94 $X2=0
+ $Y2=0
cc_191 N_A_220_53#_c_244_n N_VPWR_c_320_n 0.00785253f $X=2.81 $Y=3.03 $X2=0
+ $Y2=0
cc_192 N_A_220_53#_c_244_n N_VPWR_c_311_n 0.0219674f $X=2.81 $Y=3.03 $X2=0 $Y2=0
cc_193 N_A_220_53#_c_250_n N_VPWR_c_311_n 0.0104794f $X=2.145 $Y=2.94 $X2=0
+ $Y2=0
cc_194 N_A_220_53#_c_251_n N_VPWR_c_311_n 0.00782252f $X=2.145 $Y=2.94 $X2=0
+ $Y2=0
cc_195 N_A_220_53#_c_240_n N_X_c_357_n 0.0188702f $X=2.775 $Y=0.795 $X2=0 $Y2=0
cc_196 N_A_220_53#_M1001_g N_X_c_357_n 0.0431476f $X=2.885 $Y=2.225 $X2=0 $Y2=0
cc_197 N_A_220_53#_c_240_n N_VGND_c_371_n 0.0119613f $X=2.775 $Y=0.795 $X2=0
+ $Y2=0
cc_198 N_A_220_53#_c_243_n N_VGND_c_372_n 0.00998032f $X=1.305 $Y=0.51 $X2=0
+ $Y2=0
cc_199 N_A_220_53#_c_240_n N_VGND_c_373_n 0.00461019f $X=2.775 $Y=0.795 $X2=0
+ $Y2=0
cc_200 N_A_220_53#_c_240_n N_VGND_c_374_n 0.0105367f $X=2.775 $Y=0.795 $X2=0
+ $Y2=0
cc_201 N_A_220_53#_c_243_n N_VGND_c_374_n 0.0111908f $X=1.305 $Y=0.51 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_315_n N_X_c_357_n 0.0239368f $X=2.595 $Y=2.29 $X2=0 $Y2=0
cc_203 N_VPWR_c_311_n N_X_c_357_n 0.0136999f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_204 N_X_c_357_n N_VGND_c_373_n 0.0142544f $X=2.99 $Y=0.54 $X2=0 $Y2=0
cc_205 N_X_c_357_n N_VGND_c_374_n 0.0130144f $X=2.99 $Y=0.54 $X2=0 $Y2=0
