# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__sdlclkp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.925000 1.305000 1.315000 1.975000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.285000 1.855000 7.615000 2.045000 ;
        RECT 7.345000 0.255000 7.615000 1.855000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.415000 2.160000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.415000 0.840000 5.790000 1.565000 ;
        RECT 5.415000 1.565000 5.615000 1.830000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.095000  0.085000 0.425000 0.670000 ;
      RECT 0.095000  2.330000 0.415000 3.245000 ;
      RECT 0.585000  0.740000 0.820000 0.930000 ;
      RECT 0.585000  0.930000 0.755000 2.165000 ;
      RECT 0.585000  2.165000 2.135000 2.335000 ;
      RECT 0.585000  2.335000 1.215000 2.990000 ;
      RECT 0.595000  0.395000 0.820000 0.740000 ;
      RECT 0.990000  0.085000 1.250000 0.725000 ;
      RECT 1.420000  0.395000 1.715000 1.125000 ;
      RECT 1.465000  2.505000 1.795000 3.245000 ;
      RECT 1.485000  1.125000 1.715000 1.585000 ;
      RECT 1.485000  1.585000 2.525000 1.915000 ;
      RECT 1.905000  0.255000 2.235000 0.525000 ;
      RECT 1.905000  0.525000 5.245000 0.695000 ;
      RECT 1.905000  0.695000 2.235000 0.855000 ;
      RECT 1.965000  2.335000 2.135000 2.895000 ;
      RECT 1.965000  2.895000 3.135000 3.065000 ;
      RECT 2.305000  1.915000 2.525000 2.725000 ;
      RECT 2.535000  0.865000 2.865000 1.125000 ;
      RECT 2.695000  1.125000 2.865000 2.325000 ;
      RECT 2.695000  2.325000 3.135000 2.895000 ;
      RECT 3.045000  0.865000 3.545000 1.225000 ;
      RECT 3.045000  1.225000 4.560000 1.395000 ;
      RECT 3.305000  1.395000 3.545000 2.655000 ;
      RECT 3.715000  1.585000 4.040000 1.745000 ;
      RECT 3.715000  1.745000 4.900000 1.915000 ;
      RECT 3.915000  0.085000 4.245000 0.355000 ;
      RECT 4.045000  2.085000 4.490000 3.245000 ;
      RECT 4.300000  1.395000 4.560000 1.555000 ;
      RECT 4.425000  0.865000 4.900000 1.055000 ;
      RECT 4.660000  1.915000 4.900000 2.535000 ;
      RECT 4.660000  2.535000 5.955000 2.705000 ;
      RECT 4.660000  2.705000 4.920000 3.075000 ;
      RECT 4.730000  1.055000 4.900000 1.745000 ;
      RECT 4.985000  0.365000 5.245000 0.525000 ;
      RECT 5.070000  0.695000 5.245000 2.115000 ;
      RECT 5.070000  2.115000 5.460000 2.365000 ;
      RECT 5.415000  0.085000 5.745000 0.670000 ;
      RECT 5.640000  2.875000 5.970000 3.245000 ;
      RECT 5.785000  1.735000 6.715000 1.905000 ;
      RECT 5.785000  1.905000 5.955000 2.535000 ;
      RECT 6.150000  2.075000 7.115000 2.215000 ;
      RECT 6.150000  2.215000 8.045000 2.385000 ;
      RECT 6.150000  2.385000 6.410000 2.825000 ;
      RECT 6.205000  0.450000 6.535000 1.045000 ;
      RECT 6.205000  1.045000 7.115000 1.215000 ;
      RECT 6.385000  1.385000 6.715000 1.735000 ;
      RECT 6.580000  2.555000 7.185000 3.245000 ;
      RECT 6.845000  0.085000 7.175000 0.875000 ;
      RECT 6.895000  1.215000 7.115000 2.075000 ;
      RECT 7.715000  2.555000 8.045000 3.245000 ;
      RECT 7.785000  0.085000 8.045000 1.125000 ;
      RECT 7.785000  1.295000 8.045000 2.215000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__sdlclkp_2
END LIBRARY
