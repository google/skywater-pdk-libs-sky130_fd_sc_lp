* File: sky130_fd_sc_lp__invlp_2.pxi.spice
* Created: Wed Sep  2 09:57:07 2020
* 
x_PM_SKY130_FD_SC_LP__INVLP_2%A N_A_c_39_n N_A_M1001_g N_A_M1000_g N_A_c_41_n
+ N_A_M1002_g N_A_M1004_g N_A_c_44_n N_A_M1007_g N_A_M1005_g N_A_c_47_n
+ N_A_M1003_g N_A_M1006_g N_A_c_50_n N_A_c_51_n N_A_c_52_n A N_A_c_54_n
+ PM_SKY130_FD_SC_LP__INVLP_2%A
x_PM_SKY130_FD_SC_LP__INVLP_2%VPWR N_VPWR_M1000_d N_VPWR_M1003_d N_VPWR_c_116_n
+ N_VPWR_c_117_n N_VPWR_c_118_n N_VPWR_c_119_n VPWR N_VPWR_c_120_n
+ N_VPWR_c_115_n PM_SKY130_FD_SC_LP__INVLP_2%VPWR
x_PM_SKY130_FD_SC_LP__INVLP_2%A_116_367# N_A_116_367#_M1000_s
+ N_A_116_367#_M1005_d N_A_116_367#_c_161_n N_A_116_367#_c_148_n
+ N_A_116_367#_c_153_n N_A_116_367#_c_155_n N_A_116_367#_c_149_n
+ PM_SKY130_FD_SC_LP__INVLP_2%A_116_367#
x_PM_SKY130_FD_SC_LP__INVLP_2%Y N_Y_M1002_s N_Y_M1004_s Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__INVLP_2%Y
x_PM_SKY130_FD_SC_LP__INVLP_2%VGND N_VGND_M1001_d N_VGND_M1006_d N_VGND_c_196_n
+ N_VGND_c_197_n N_VGND_c_198_n N_VGND_c_199_n VGND N_VGND_c_200_n
+ N_VGND_c_201_n PM_SKY130_FD_SC_LP__INVLP_2%VGND
x_PM_SKY130_FD_SC_LP__INVLP_2%A_116_55# N_A_116_55#_M1001_s N_A_116_55#_M1007_d
+ N_A_116_55#_c_224_n N_A_116_55#_c_225_n N_A_116_55#_c_226_n
+ PM_SKY130_FD_SC_LP__INVLP_2%A_116_55#
cc_1 VNB N_A_c_39_n 0.0205056f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.225
cc_2 VNB N_A_M1000_g 0.00795969f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_3 VNB N_A_c_41_n 0.0091677f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.48
cc_4 VNB N_A_M1002_g 0.0241531f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.695
cc_5 VNB N_A_M1004_g 0.00462086f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_6 VNB N_A_c_44_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.48
cc_7 VNB N_A_M1007_g 0.0253153f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.695
cc_8 VNB N_A_M1005_g 0.00462086f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=2.465
cc_9 VNB N_A_c_47_n 0.0111229f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.48
cc_10 VNB N_A_M1003_g 0.00795969f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=2.465
cc_11 VNB N_A_M1006_g 0.0367191f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=0.695
cc_12 VNB N_A_c_50_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.48
cc_13 VNB N_A_c_51_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.48
cc_14 VNB N_A_c_52_n 0.0150011f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.48
cc_15 VNB A 0.0078043f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_A_c_54_n 0.0542323f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.39
cc_17 VNB N_VPWR_c_115_n 0.103974f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.405
cc_18 VNB N_VGND_c_196_n 0.0116259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_197_n 0.032819f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.48
cc_20 VNB N_VGND_c_198_n 0.0119539f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.695
cc_21 VNB N_VGND_c_199_n 0.0432976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_200_n 0.0366672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_201_n 0.16146f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.555
cc_24 VNB N_A_116_55#_c_224_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.48
cc_25 VNB N_A_116_55#_c_225_n 0.00406927f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.555
cc_26 VNB N_A_116_55#_c_226_n 0.00790931f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_27 VPB N_A_M1000_g 0.0265103f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_28 VPB N_A_M1004_g 0.0190413f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_29 VPB N_A_M1005_g 0.0190413f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=2.465
cc_30 VPB N_A_M1003_g 0.0271666f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=2.465
cc_31 VPB N_VPWR_c_116_n 0.0112967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_117_n 0.0535295f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.48
cc_33 VPB N_VPWR_c_118_n 0.0134631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_119_n 0.0611798f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_35 VPB N_VPWR_c_120_n 0.0345412f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=0.695
cc_36 VPB N_VPWR_c_115_n 0.0470547f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=1.405
cc_37 VPB N_A_116_367#_c_148_n 0.00261677f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.48
cc_38 VPB N_A_116_367#_c_149_n 0.00339227f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_39 N_A_M1000_g N_VPWR_c_117_n 0.023916f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_40 N_A_M1004_g N_VPWR_c_117_n 0.00109254f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_41 A N_VPWR_c_117_n 0.0202789f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_42 N_A_c_54_n N_VPWR_c_117_n 0.002285f $X=0.58 $Y=1.39 $X2=0 $Y2=0
cc_43 N_A_M1003_g N_VPWR_c_119_n 0.0294905f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_44 N_A_c_52_n N_VPWR_c_119_n 0.00105441f $X=1.83 $Y=1.48 $X2=0 $Y2=0
cc_45 N_A_M1000_g N_VPWR_c_120_n 0.00486043f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_46 N_A_M1004_g N_VPWR_c_120_n 0.00357877f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_47 N_A_M1005_g N_VPWR_c_120_n 0.00357877f $X=1.365 $Y=2.465 $X2=0 $Y2=0
cc_48 N_A_M1003_g N_VPWR_c_120_n 0.00547432f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_49 N_A_M1000_g N_VPWR_c_115_n 0.00824727f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_50 N_A_M1004_g N_VPWR_c_115_n 0.0053512f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_51 N_A_M1005_g N_VPWR_c_115_n 0.0053512f $X=1.365 $Y=2.465 $X2=0 $Y2=0
cc_52 N_A_M1003_g N_VPWR_c_115_n 0.01095f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_53 N_A_M1000_g N_A_116_367#_c_148_n 7.7109e-19 $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_54 N_A_c_41_n N_A_116_367#_c_148_n 0.00238955f $X=0.86 $Y=1.48 $X2=0 $Y2=0
cc_55 N_A_M1004_g N_A_116_367#_c_148_n 7.7109e-19 $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_56 N_A_M1004_g N_A_116_367#_c_153_n 0.0115031f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_57 N_A_M1005_g N_A_116_367#_c_153_n 0.0114565f $X=1.365 $Y=2.465 $X2=0 $Y2=0
cc_58 N_A_M1003_g N_A_116_367#_c_155_n 0.00202381f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A_M1005_g N_A_116_367#_c_149_n 7.76258e-19 $X=1.365 $Y=2.465 $X2=0 $Y2=0
cc_60 N_A_c_47_n N_A_116_367#_c_149_n 0.00238955f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_61 N_A_M1003_g N_A_116_367#_c_149_n 0.013891f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_62 N_A_c_39_n Y 0.00115202f $X=0.505 $Y=1.225 $X2=0 $Y2=0
cc_63 N_A_M1000_g Y 0.0015375f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A_M1002_g Y 0.0156977f $X=0.935 $Y=0.695 $X2=0 $Y2=0
cc_65 N_A_M1004_g Y 0.0203222f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_c_44_n Y 0.00874467f $X=1.29 $Y=1.48 $X2=0 $Y2=0
cc_67 N_A_M1007_g Y 0.0160964f $X=1.365 $Y=0.695 $X2=0 $Y2=0
cc_68 N_A_M1005_g Y 0.0203222f $X=1.365 $Y=2.465 $X2=0 $Y2=0
cc_69 N_A_M1003_g Y 0.00161469f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_M1006_g Y 0.0014821f $X=1.865 $Y=0.695 $X2=0 $Y2=0
cc_71 N_A_c_50_n Y 0.00429115f $X=0.935 $Y=1.48 $X2=0 $Y2=0
cc_72 N_A_c_51_n Y 0.00721695f $X=1.365 $Y=1.48 $X2=0 $Y2=0
cc_73 A Y 0.0110608f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_c_39_n N_VGND_c_197_n 0.0142238f $X=0.505 $Y=1.225 $X2=0 $Y2=0
cc_75 N_A_M1002_g N_VGND_c_197_n 8.80913e-19 $X=0.935 $Y=0.695 $X2=0 $Y2=0
cc_76 A N_VGND_c_197_n 0.0260923f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_54_n N_VGND_c_197_n 0.00197323f $X=0.58 $Y=1.39 $X2=0 $Y2=0
cc_78 N_A_M1006_g N_VGND_c_199_n 0.00775936f $X=1.865 $Y=0.695 $X2=0 $Y2=0
cc_79 N_A_c_39_n N_VGND_c_200_n 0.00452967f $X=0.505 $Y=1.225 $X2=0 $Y2=0
cc_80 N_A_M1002_g N_VGND_c_200_n 0.00332046f $X=0.935 $Y=0.695 $X2=0 $Y2=0
cc_81 N_A_M1007_g N_VGND_c_200_n 0.00332046f $X=1.365 $Y=0.695 $X2=0 $Y2=0
cc_82 N_A_M1006_g N_VGND_c_200_n 0.00509933f $X=1.865 $Y=0.695 $X2=0 $Y2=0
cc_83 N_A_c_39_n N_VGND_c_201_n 0.00815021f $X=0.505 $Y=1.225 $X2=0 $Y2=0
cc_84 N_A_M1002_g N_VGND_c_201_n 0.00498029f $X=0.935 $Y=0.695 $X2=0 $Y2=0
cc_85 N_A_M1007_g N_VGND_c_201_n 0.00511192f $X=1.365 $Y=0.695 $X2=0 $Y2=0
cc_86 N_A_M1006_g N_VGND_c_201_n 0.0103814f $X=1.865 $Y=0.695 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_A_116_55#_c_224_n 0.0115336f $X=0.935 $Y=0.695 $X2=0 $Y2=0
cc_88 N_A_M1007_g N_A_116_55#_c_224_n 0.0137818f $X=1.365 $Y=0.695 $X2=0 $Y2=0
cc_89 N_A_c_39_n N_A_116_55#_c_225_n 0.00113103f $X=0.505 $Y=1.225 $X2=0 $Y2=0
cc_90 N_A_c_41_n N_A_116_55#_c_225_n 0.00235845f $X=0.86 $Y=1.48 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_A_116_55#_c_225_n 8.13177e-19 $X=0.935 $Y=0.695 $X2=0 $Y2=0
cc_92 N_A_M1007_g N_A_116_55#_c_226_n 0.00376406f $X=1.365 $Y=0.695 $X2=0 $Y2=0
cc_93 N_A_c_47_n N_A_116_55#_c_226_n 0.00446702f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_94 N_A_M1006_g N_A_116_55#_c_226_n 0.0134733f $X=1.865 $Y=0.695 $X2=0 $Y2=0
cc_95 N_VPWR_c_115_n N_A_116_367#_M1000_s 0.00411415f $X=2.16 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_96 N_VPWR_c_115_n N_A_116_367#_M1005_d 0.00223562f $X=2.16 $Y=3.33 $X2=0
+ $Y2=0
cc_97 N_VPWR_c_120_n N_A_116_367#_c_161_n 0.0118138f $X=1.915 $Y=3.33 $X2=0
+ $Y2=0
cc_98 N_VPWR_c_115_n N_A_116_367#_c_161_n 0.00658808f $X=2.16 $Y=3.33 $X2=0
+ $Y2=0
cc_99 N_VPWR_c_117_n N_A_116_367#_c_148_n 0.0397536f $X=0.29 $Y=1.98 $X2=0 $Y2=0
cc_100 N_VPWR_c_120_n N_A_116_367#_c_153_n 0.0368226f $X=1.915 $Y=3.33 $X2=0
+ $Y2=0
cc_101 N_VPWR_c_115_n N_A_116_367#_c_153_n 0.024428f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_102 N_VPWR_c_120_n N_A_116_367#_c_155_n 0.0154369f $X=1.915 $Y=3.33 $X2=0
+ $Y2=0
cc_103 N_VPWR_c_115_n N_A_116_367#_c_155_n 0.00952129f $X=2.16 $Y=3.33 $X2=0
+ $Y2=0
cc_104 N_VPWR_c_119_n N_A_116_367#_c_149_n 0.0399503f $X=2.08 $Y=1.98 $X2=0
+ $Y2=0
cc_105 N_VPWR_c_115_n N_Y_M1004_s 0.00225186f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_106 N_VPWR_c_119_n N_VGND_c_199_n 0.00876255f $X=2.08 $Y=1.98 $X2=0 $Y2=0
cc_107 N_A_116_367#_c_153_n N_Y_M1004_s 0.00332344f $X=1.495 $Y=2.99 $X2=0 $Y2=0
cc_108 N_A_116_367#_c_148_n Y 0.0336606f $X=0.72 $Y=1.98 $X2=0 $Y2=0
cc_109 N_A_116_367#_c_153_n Y 0.0159805f $X=1.495 $Y=2.99 $X2=0 $Y2=0
cc_110 N_A_116_367#_c_149_n Y 0.033702f $X=1.58 $Y=1.98 $X2=0 $Y2=0
cc_111 N_A_116_367#_c_148_n N_A_116_55#_c_225_n 0.00589417f $X=0.72 $Y=1.98
+ $X2=0 $Y2=0
cc_112 N_A_116_367#_c_149_n N_A_116_55#_c_226_n 0.00859865f $X=1.58 $Y=1.98
+ $X2=0 $Y2=0
cc_113 N_Y_M1002_s N_A_116_55#_c_224_n 0.00176461f $X=1.01 $Y=0.275 $X2=0.58
+ $Y2=1.48
cc_114 Y N_A_116_55#_c_224_n 0.0160549f $X=1.115 $Y=0.84 $X2=0.58 $Y2=1.48
cc_115 Y N_A_116_55#_c_225_n 0.0200409f $X=1.115 $Y=0.84 $X2=0.935 $Y2=1.555
cc_116 Y N_A_116_55#_c_226_n 0.0210526f $X=1.115 $Y=0.84 $X2=0.935 $Y2=2.465
cc_117 N_VGND_c_200_n N_A_116_55#_c_224_n 0.0428729f $X=1.995 $Y=0 $X2=0 $Y2=0
cc_118 N_VGND_c_201_n N_A_116_55#_c_224_n 0.0241933f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_119 N_VGND_c_197_n N_A_116_55#_c_225_n 0.00697079f $X=0.29 $Y=0.42 $X2=0
+ $Y2=0
cc_120 N_VGND_c_200_n N_A_116_55#_c_225_n 0.0121867f $X=1.995 $Y=0 $X2=0 $Y2=0
cc_121 N_VGND_c_201_n N_A_116_55#_c_225_n 0.00660921f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_122 N_VGND_c_199_n N_A_116_55#_c_226_n 0.0337087f $X=2.08 $Y=0.42 $X2=0 $Y2=0
cc_123 N_VGND_c_200_n N_A_116_55#_c_226_n 0.0235688f $X=1.995 $Y=0 $X2=0 $Y2=0
cc_124 N_VGND_c_201_n N_A_116_55#_c_226_n 0.0127152f $X=2.16 $Y=0 $X2=0 $Y2=0
