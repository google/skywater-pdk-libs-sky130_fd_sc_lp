* File: sky130_fd_sc_lp__a2bb2oi_1.spice
* Created: Wed Sep  2 09:24:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2oi_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1003 N_A_113_47#_M1003_d N_A1_N_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A2_N_M1006_g N_A_113_47#_M1003_d VNB NSHORT L=0.15
+ W=0.84 AD=0.3192 AS=0.1176 PD=1.6 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_A_113_47#_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3192 PD=1.12 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5 SB=75001.2
+ A=0.126 P=1.98 MULT=1
MM1007 A_467_47# N_B2_M1007_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.84 AD=0.1596
+ AS=0.1176 PD=1.22 PS=1.12 NRD=19.284 NRS=0 M=1 R=5.6 SA=75002 SB=75000.7
+ A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g A_467_47# VNB NSHORT L=0.15 W=0.84 AD=0.2436
+ AS=0.1596 PD=2.26 PS=1.22 NRD=3.564 NRS=19.284 M=1 R=5.6 SA=75002.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1005 A_113_367# N_A1_N_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.3339 PD=1.5 PS=3.05 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_A_113_47#_M1008_d N_A2_N_M1008_g A_113_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1512 PD=3.05 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_A_381_367#_M1002_d N_A_113_47#_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.17955 AS=0.3339 PD=1.545 PS=3.05 NRD=0.7683 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_B2_M1009_g N_A_381_367#_M1002_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.252 AS=0.17955 PD=1.66 PS=1.545 NRD=10.1455 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1000 N_A_381_367#_M1000_d N_B1_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.252 PD=3.05 PS=1.66 NRD=0 NRS=8.5892 M=1 R=8.4
+ SA=75001.2 SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a2bb2oi_1.pxi.spice"
*
.ends
*
*
