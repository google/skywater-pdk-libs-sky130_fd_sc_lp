* File: sky130_fd_sc_lp__and2_lp.pxi.spice
* Created: Fri Aug 28 10:04:44 2020
* 
x_PM_SKY130_FD_SC_LP__AND2_LP%B N_B_M1008_g N_B_M1002_g N_B_M1005_g N_B_c_53_n
+ N_B_c_59_n B B B N_B_c_55_n PM_SKY130_FD_SC_LP__AND2_LP%B
x_PM_SKY130_FD_SC_LP__AND2_LP%A N_A_c_89_n N_A_M1007_g N_A_c_90_n N_A_c_96_n
+ N_A_M1004_g N_A_c_97_n N_A_c_91_n N_A_c_98_n N_A_M1003_g N_A_c_92_n N_A_c_99_n
+ A A N_A_c_94_n PM_SKY130_FD_SC_LP__AND2_LP%A
x_PM_SKY130_FD_SC_LP__AND2_LP%A_213_468# N_A_213_468#_M1007_d
+ N_A_213_468#_M1005_d N_A_213_468#_M1009_g N_A_213_468#_M1000_g
+ N_A_213_468#_M1006_g N_A_213_468#_M1001_g N_A_213_468#_c_150_n
+ N_A_213_468#_c_151_n N_A_213_468#_c_158_n N_A_213_468#_c_152_n
+ N_A_213_468#_c_153_n N_A_213_468#_c_154_n
+ PM_SKY130_FD_SC_LP__AND2_LP%A_213_468#
x_PM_SKY130_FD_SC_LP__AND2_LP%VPWR N_VPWR_M1008_s N_VPWR_M1003_d N_VPWR_c_226_n
+ N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n N_VPWR_c_230_n VPWR
+ N_VPWR_c_231_n N_VPWR_c_225_n PM_SKY130_FD_SC_LP__AND2_LP%VPWR
x_PM_SKY130_FD_SC_LP__AND2_LP%X N_X_M1001_d N_X_M1006_d X X X X X X X
+ PM_SKY130_FD_SC_LP__AND2_LP%X
x_PM_SKY130_FD_SC_LP__AND2_LP%VGND N_VGND_M1002_s N_VGND_M1000_s N_VGND_c_275_n
+ N_VGND_c_276_n VGND N_VGND_c_277_n N_VGND_c_278_n N_VGND_c_279_n
+ N_VGND_c_280_n N_VGND_c_281_n N_VGND_c_282_n PM_SKY130_FD_SC_LP__AND2_LP%VGND
cc_1 VNB N_B_M1002_g 0.0281255f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.08
cc_2 VNB N_B_c_53_n 7.45465e-19 $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2
cc_3 VNB B 0.0326678f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_B_c_55_n 0.0178016f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.645
cc_5 VNB N_A_c_89_n 0.0164208f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.15
cc_6 VNB N_A_c_90_n 0.00460665f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.48
cc_7 VNB N_A_c_91_n 0.0406366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_c_92_n 0.0339689f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.075
cc_9 VNB A 0.0180565f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_10 VNB N_A_c_94_n 0.0410085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_213_468#_M1000_g 0.0218885f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.645
cc_12 VNB N_A_213_468#_M1001_g 0.0243843f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_A_213_468#_c_150_n 0.00202741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_213_468#_c_151_n 0.0147756f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_15 VNB N_A_213_468#_c_152_n 0.00677372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_213_468#_c_153_n 0.00322564f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.815
cc_17 VNB N_A_213_468#_c_154_n 0.0851308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_225_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB X 0.0664723f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.08
cc_20 VNB N_VGND_c_275_n 0.0637196f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.15
cc_21 VNB N_VGND_c_276_n 0.0196758f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.645
cc_22 VNB N_VGND_c_277_n 0.0158267f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.075
cc_23 VNB N_VGND_c_278_n 0.0339475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_279_n 0.0298078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_280_n 0.23791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_281_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.645
cc_27 VNB N_VGND_c_282_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.815
cc_28 VPB N_B_M1008_g 0.0262787f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.55
cc_29 VPB N_B_M1005_g 0.0199715f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.55
cc_30 VPB N_B_c_53_n 0.0284933f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2
cc_31 VPB N_B_c_59_n 0.0211535f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.075
cc_32 VPB B 0.0394529f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_33 VPB N_A_c_90_n 0.0242228f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1.48
cc_34 VPB N_A_c_96_n 0.0154264f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1.08
cc_35 VPB N_A_c_97_n 0.0201198f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.15
cc_36 VPB N_A_c_98_n 0.0153012f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.645
cc_37 VPB N_A_c_99_n 0.00532081f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_38 VPB N_A_213_468#_M1009_g 0.0429083f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.15
cc_39 VPB N_A_213_468#_M1006_g 0.0472331f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.075
cc_40 VPB N_A_213_468#_c_150_n 0.00617343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_213_468#_c_158_n 0.00928467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_213_468#_c_153_n 0.00175225f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.815
cc_43 VPB N_A_213_468#_c_154_n 0.0151729f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_226_n 0.0164972f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1.08
cc_45 VPB N_VPWR_c_227_n 0.0466455f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.15
cc_46 VPB N_VPWR_c_228_n 0.0290375f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.645
cc_47 VPB N_VPWR_c_229_n 0.0364721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_230_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.075
cc_49 VPB N_VPWR_c_231_n 0.0356949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_225_n 0.0930127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB X 0.0746537f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1.08
cc_52 N_B_M1002_g N_A_c_89_n 0.0210101f $X=0.81 $Y=1.08 $X2=-0.19 $Y2=-0.245
cc_53 N_B_c_59_n N_A_c_90_n 0.0117699f $X=0.99 $Y=2.075 $X2=0 $Y2=0
cc_54 B N_A_c_90_n 0.00666703f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_55 N_B_c_55_n N_A_c_90_n 0.00889885f $X=0.72 $Y=1.645 $X2=0 $Y2=0
cc_56 B N_A_c_92_n 0.0147942f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_57 N_B_c_55_n N_A_c_92_n 0.0210101f $X=0.72 $Y=1.645 $X2=0 $Y2=0
cc_58 N_B_M1005_g N_A_c_99_n 0.0117699f $X=0.99 $Y=2.55 $X2=0 $Y2=0
cc_59 N_B_M1002_g N_A_213_468#_c_150_n 2.66747e-19 $X=0.81 $Y=1.08 $X2=0 $Y2=0
cc_60 N_B_c_59_n N_A_213_468#_c_150_n 9.18205e-19 $X=0.99 $Y=2.075 $X2=0 $Y2=0
cc_61 B N_A_213_468#_c_150_n 0.0535094f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_62 N_B_c_55_n N_A_213_468#_c_150_n 3.02549e-19 $X=0.72 $Y=1.645 $X2=0 $Y2=0
cc_63 N_B_M1008_g N_A_213_468#_c_158_n 0.00124255f $X=0.63 $Y=2.55 $X2=0 $Y2=0
cc_64 N_B_M1005_g N_A_213_468#_c_158_n 0.00883826f $X=0.99 $Y=2.55 $X2=0 $Y2=0
cc_65 B N_A_213_468#_c_158_n 0.0245604f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_66 N_B_M1002_g N_A_213_468#_c_152_n 0.0012945f $X=0.81 $Y=1.08 $X2=0 $Y2=0
cc_67 B N_A_213_468#_c_152_n 0.00545584f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_68 N_B_M1008_g N_VPWR_c_227_n 0.0137486f $X=0.63 $Y=2.55 $X2=0 $Y2=0
cc_69 N_B_M1005_g N_VPWR_c_227_n 0.00180764f $X=0.99 $Y=2.55 $X2=0 $Y2=0
cc_70 B N_VPWR_c_227_n 0.0303461f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_71 N_B_M1008_g N_VPWR_c_229_n 0.00370277f $X=0.63 $Y=2.55 $X2=0 $Y2=0
cc_72 N_B_M1005_g N_VPWR_c_229_n 0.00427474f $X=0.99 $Y=2.55 $X2=0 $Y2=0
cc_73 N_B_M1008_g N_VPWR_c_225_n 0.00407315f $X=0.63 $Y=2.55 $X2=0 $Y2=0
cc_74 N_B_M1005_g N_VPWR_c_225_n 0.00484898f $X=0.99 $Y=2.55 $X2=0 $Y2=0
cc_75 N_B_M1002_g N_VGND_c_275_n 0.0141543f $X=0.81 $Y=1.08 $X2=0 $Y2=0
cc_76 B N_VGND_c_275_n 0.0295293f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_77 N_B_c_55_n N_VGND_c_275_n 0.00490317f $X=0.72 $Y=1.645 $X2=0 $Y2=0
cc_78 N_B_M1002_g N_VGND_c_278_n 0.00255106f $X=0.81 $Y=1.08 $X2=0 $Y2=0
cc_79 N_B_M1002_g N_VGND_c_280_n 0.00341643f $X=0.81 $Y=1.08 $X2=0 $Y2=0
cc_80 N_A_c_90_n N_A_213_468#_M1009_g 0.0030445f $X=1.42 $Y=2.08 $X2=0 $Y2=0
cc_81 N_A_c_97_n N_A_213_468#_M1009_g 0.0191631f $X=1.705 $Y=2.155 $X2=0 $Y2=0
cc_82 N_A_c_91_n N_A_213_468#_M1000_g 0.00581069f $X=1.71 $Y=1.4 $X2=0 $Y2=0
cc_83 N_A_c_94_n N_A_213_468#_M1000_g 0.00482222f $X=1.68 $Y=0.515 $X2=0 $Y2=0
cc_84 N_A_c_89_n N_A_213_468#_c_150_n 0.00183833f $X=1.2 $Y=1.4 $X2=0 $Y2=0
cc_85 N_A_c_90_n N_A_213_468#_c_150_n 0.00956222f $X=1.42 $Y=2.08 $X2=0 $Y2=0
cc_86 N_A_c_96_n N_A_213_468#_c_150_n 0.00200441f $X=1.42 $Y=2.23 $X2=0 $Y2=0
cc_87 N_A_c_97_n N_A_213_468#_c_150_n 0.0080989f $X=1.705 $Y=2.155 $X2=0 $Y2=0
cc_88 N_A_c_91_n N_A_213_468#_c_150_n 0.0021284f $X=1.71 $Y=1.4 $X2=0 $Y2=0
cc_89 N_A_c_98_n N_A_213_468#_c_150_n 0.00207138f $X=1.78 $Y=2.23 $X2=0 $Y2=0
cc_90 N_A_c_92_n N_A_213_468#_c_150_n 0.0104599f $X=1.71 $Y=1.475 $X2=0 $Y2=0
cc_91 N_A_c_99_n N_A_213_468#_c_150_n 0.00192878f $X=1.42 $Y=2.155 $X2=0 $Y2=0
cc_92 N_A_c_91_n N_A_213_468#_c_151_n 0.011889f $X=1.71 $Y=1.4 $X2=0 $Y2=0
cc_93 A N_A_213_468#_c_151_n 0.00626362f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_94 N_A_c_94_n N_A_213_468#_c_151_n 0.00108337f $X=1.68 $Y=0.515 $X2=0 $Y2=0
cc_95 N_A_c_96_n N_A_213_468#_c_158_n 0.0191527f $X=1.42 $Y=2.23 $X2=0 $Y2=0
cc_96 N_A_c_97_n N_A_213_468#_c_158_n 2.11001e-19 $X=1.705 $Y=2.155 $X2=0 $Y2=0
cc_97 N_A_c_98_n N_A_213_468#_c_158_n 0.00164761f $X=1.78 $Y=2.23 $X2=0 $Y2=0
cc_98 N_A_c_89_n N_A_213_468#_c_152_n 0.00917376f $X=1.2 $Y=1.4 $X2=0 $Y2=0
cc_99 N_A_c_91_n N_A_213_468#_c_152_n 0.0128644f $X=1.71 $Y=1.4 $X2=0 $Y2=0
cc_100 N_A_c_92_n N_A_213_468#_c_152_n 0.0063659f $X=1.71 $Y=1.475 $X2=0 $Y2=0
cc_101 A N_A_213_468#_c_152_n 0.0329806f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_102 N_A_c_94_n N_A_213_468#_c_152_n 0.0024137f $X=1.68 $Y=0.515 $X2=0 $Y2=0
cc_103 N_A_c_91_n N_A_213_468#_c_153_n 0.00122938f $X=1.71 $Y=1.4 $X2=0 $Y2=0
cc_104 N_A_c_90_n N_A_213_468#_c_154_n 0.00183687f $X=1.42 $Y=2.08 $X2=0 $Y2=0
cc_105 N_A_c_91_n N_A_213_468#_c_154_n 0.0264768f $X=1.71 $Y=1.4 $X2=0 $Y2=0
cc_106 N_A_c_96_n N_VPWR_c_228_n 9.12371e-19 $X=1.42 $Y=2.23 $X2=0 $Y2=0
cc_107 N_A_c_98_n N_VPWR_c_228_n 0.0103045f $X=1.78 $Y=2.23 $X2=0 $Y2=0
cc_108 N_A_c_96_n N_VPWR_c_229_n 0.00337271f $X=1.42 $Y=2.23 $X2=0 $Y2=0
cc_109 N_A_c_98_n N_VPWR_c_229_n 0.00370277f $X=1.78 $Y=2.23 $X2=0 $Y2=0
cc_110 N_A_c_96_n N_VPWR_c_225_n 0.00484898f $X=1.42 $Y=2.23 $X2=0 $Y2=0
cc_111 N_A_c_98_n N_VPWR_c_225_n 0.00407315f $X=1.78 $Y=2.23 $X2=0 $Y2=0
cc_112 N_A_c_89_n N_VGND_c_275_n 0.00185091f $X=1.2 $Y=1.4 $X2=0 $Y2=0
cc_113 A N_VGND_c_275_n 0.018489f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_114 N_A_c_91_n N_VGND_c_276_n 0.00459435f $X=1.71 $Y=1.4 $X2=0 $Y2=0
cc_115 A N_VGND_c_276_n 0.0275242f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_116 N_A_c_94_n N_VGND_c_276_n 0.00133138f $X=1.68 $Y=0.515 $X2=0 $Y2=0
cc_117 A N_VGND_c_278_n 0.0311813f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_118 N_A_c_94_n N_VGND_c_278_n 0.00722827f $X=1.68 $Y=0.515 $X2=0 $Y2=0
cc_119 A N_VGND_c_280_n 0.0271378f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_120 N_A_c_94_n N_VGND_c_280_n 0.0105548f $X=1.68 $Y=0.515 $X2=0 $Y2=0
cc_121 N_A_213_468#_c_158_n N_VPWR_c_227_n 0.0161226f $X=1.57 $Y=2.55 $X2=0
+ $Y2=0
cc_122 N_A_213_468#_M1009_g N_VPWR_c_228_n 0.0114062f $X=2.21 $Y=2.55 $X2=0
+ $Y2=0
cc_123 N_A_213_468#_M1006_g N_VPWR_c_228_n 0.00146455f $X=2.57 $Y=2.55 $X2=0
+ $Y2=0
cc_124 N_A_213_468#_c_158_n N_VPWR_c_228_n 0.0184869f $X=1.57 $Y=2.55 $X2=0
+ $Y2=0
cc_125 N_A_213_468#_c_153_n N_VPWR_c_228_n 0.0045587f $X=2.19 $Y=1.235 $X2=0
+ $Y2=0
cc_126 N_A_213_468#_c_154_n N_VPWR_c_228_n 6.92319e-19 $X=2.57 $Y=1.405 $X2=0
+ $Y2=0
cc_127 N_A_213_468#_c_158_n N_VPWR_c_229_n 0.0141497f $X=1.57 $Y=2.55 $X2=0
+ $Y2=0
cc_128 N_A_213_468#_M1009_g N_VPWR_c_231_n 0.00370277f $X=2.21 $Y=2.55 $X2=0
+ $Y2=0
cc_129 N_A_213_468#_M1006_g N_VPWR_c_231_n 0.00151879f $X=2.57 $Y=2.55 $X2=0
+ $Y2=0
cc_130 N_A_213_468#_M1009_g N_VPWR_c_225_n 0.00407315f $X=2.21 $Y=2.55 $X2=0
+ $Y2=0
cc_131 N_A_213_468#_M1006_g N_VPWR_c_225_n 0.00100212f $X=2.57 $Y=2.55 $X2=0
+ $Y2=0
cc_132 N_A_213_468#_c_158_n N_VPWR_c_225_n 0.0193086f $X=1.57 $Y=2.55 $X2=0
+ $Y2=0
cc_133 N_A_213_468#_M1009_g X 0.00533964f $X=2.21 $Y=2.55 $X2=0 $Y2=0
cc_134 N_A_213_468#_M1000_g X 0.007102f $X=2.395 $Y=0.67 $X2=0 $Y2=0
cc_135 N_A_213_468#_M1006_g X 0.0447568f $X=2.57 $Y=2.55 $X2=0 $Y2=0
cc_136 N_A_213_468#_M1001_g X 0.0202622f $X=2.785 $Y=0.67 $X2=0 $Y2=0
cc_137 N_A_213_468#_c_153_n X 0.0542106f $X=2.19 $Y=1.235 $X2=0 $Y2=0
cc_138 N_A_213_468#_c_154_n X 0.0423435f $X=2.57 $Y=1.405 $X2=0 $Y2=0
cc_139 N_A_213_468#_c_152_n N_VGND_c_275_n 0.0149998f $X=1.655 $Y=1.08 $X2=0
+ $Y2=0
cc_140 N_A_213_468#_M1000_g N_VGND_c_276_n 0.0102448f $X=2.395 $Y=0.67 $X2=0
+ $Y2=0
cc_141 N_A_213_468#_M1001_g N_VGND_c_276_n 9.01033e-19 $X=2.785 $Y=0.67 $X2=0
+ $Y2=0
cc_142 N_A_213_468#_c_151_n N_VGND_c_276_n 5.67176e-19 $X=2.025 $Y=1.225 $X2=0
+ $Y2=0
cc_143 N_A_213_468#_c_152_n N_VGND_c_276_n 0.00225609f $X=1.655 $Y=1.08 $X2=0
+ $Y2=0
cc_144 N_A_213_468#_c_153_n N_VGND_c_276_n 0.0283019f $X=2.19 $Y=1.235 $X2=0
+ $Y2=0
cc_145 N_A_213_468#_c_154_n N_VGND_c_276_n 0.00230793f $X=2.57 $Y=1.405 $X2=0
+ $Y2=0
cc_146 N_A_213_468#_M1000_g N_VGND_c_279_n 0.00426961f $X=2.395 $Y=0.67 $X2=0
+ $Y2=0
cc_147 N_A_213_468#_M1001_g N_VGND_c_279_n 0.00375632f $X=2.785 $Y=0.67 $X2=0
+ $Y2=0
cc_148 N_A_213_468#_M1000_g N_VGND_c_280_n 0.00434697f $X=2.395 $Y=0.67 $X2=0
+ $Y2=0
cc_149 N_A_213_468#_M1001_g N_VGND_c_280_n 0.00517496f $X=2.785 $Y=0.67 $X2=0
+ $Y2=0
cc_150 N_VPWR_c_228_n X 0.0245928f $X=1.995 $Y=2.55 $X2=0 $Y2=0
cc_151 N_VPWR_c_231_n X 0.022836f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_152 N_VPWR_c_225_n X 0.0245694f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_153 X N_VGND_c_276_n 0.0181917f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_154 X N_VGND_c_279_n 0.0227539f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_155 X N_VGND_c_280_n 0.0245391f $X=2.555 $Y=0.47 $X2=0 $Y2=0
