* File: sky130_fd_sc_lp__a41oi_m.pex.spice
* Created: Wed Sep  2 09:30:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41OI_M%B1 3 4 9 13 16 17 18 19 20 21 22 23 24 25 32
r51 24 25 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=2.405
+ $X2=0.71 $Y2=2.775
r52 23 24 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=2.035
+ $X2=0.71 $Y2=2.405
r53 22 23 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=1.665
+ $X2=0.71 $Y2=2.035
r54 21 22 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=1.295
+ $X2=0.71 $Y2=1.665
r55 21 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.7
+ $Y=1.375 $X2=0.7 $Y2=1.375
r56 19 20 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=0.822 $Y=2.12
+ $X2=0.822 $Y2=2.27
r57 18 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.79 $Y=1.88
+ $X2=0.79 $Y2=2.12
r58 17 32 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.7 $Y=1.715 $X2=0.7
+ $Y2=1.375
r59 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.7 $Y=1.715
+ $X2=0.7 $Y2=1.88
r60 16 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.7 $Y=1.21 $X2=0.7
+ $Y2=1.375
r61 11 13 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.995 $Y=0.82
+ $X2=0.995 $Y2=0.445
r62 9 20 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=0.855 $Y=2.865
+ $X2=0.855 $Y2=2.27
r63 3 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.92 $Y=0.895
+ $X2=0.995 $Y2=0.82
r64 3 4 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=0.92 $Y=0.895 $X2=0.685
+ $Y2=0.895
r65 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.61 $Y=0.97
+ $X2=0.685 $Y2=0.895
r66 1 16 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.61 $Y=0.97 $X2=0.61
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_M%A1 2 5 11 12 13 14 15 16 17 22 24
r55 22 24 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.252 $Y=1.375
+ $X2=1.252 $Y2=1.21
r56 16 17 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=2.035
r57 15 16 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.22 $Y=1.295
+ $X2=1.22 $Y2=1.665
r58 15 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.24
+ $Y=1.375 $X2=1.24 $Y2=1.375
r59 14 24 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=1.355 $Y=0.915
+ $X2=1.355 $Y2=1.21
r60 13 14 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.39 $Y=0.765
+ $X2=1.39 $Y2=0.915
r61 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.425 $Y=0.445
+ $X2=1.425 $Y2=0.765
r62 5 12 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=1.285 $Y=2.865
+ $X2=1.285 $Y2=1.88
r63 2 12 40.5352 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=1.252 $Y=1.703
+ $X2=1.252 $Y2=1.88
r64 1 22 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=1.252 $Y=1.387
+ $X2=1.252 $Y2=1.375
r65 1 2 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=1.252 $Y=1.387
+ $X2=1.252 $Y2=1.703
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_M%A2 3 7 11 12 13 14 15 16 17 24
c47 12 0 1.18907e-19 $X=1.805 $Y=1.795
c48 7 0 2.08874e-19 $X=1.785 $Y=0.445
r49 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.805
+ $Y=1.29 $X2=1.805 $Y2=1.29
r50 16 17 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.742 $Y=1.665
+ $X2=1.742 $Y2=2.035
r51 15 16 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.742 $Y=1.295
+ $X2=1.742 $Y2=1.665
r52 15 25 0.195329 $w=2.93e-07 $l=5e-09 $layer=LI1_cond $X=1.742 $Y=1.295
+ $X2=1.742 $Y2=1.29
r53 14 25 14.259 $w=2.93e-07 $l=3.65e-07 $layer=LI1_cond $X=1.742 $Y=0.925
+ $X2=1.742 $Y2=1.29
r54 13 14 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.742 $Y=0.555
+ $X2=1.742 $Y2=0.925
r55 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.805 $Y=1.63
+ $X2=1.805 $Y2=1.29
r56 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.63
+ $X2=1.805 $Y2=1.795
r57 10 24 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.125
+ $X2=1.805 $Y2=1.29
r58 7 10 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.785 $Y=0.445
+ $X2=1.785 $Y2=1.125
r59 3 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.715 $Y=2.865
+ $X2=1.715 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_M%A3 3 7 11 12 13 14 15 16 22
c48 12 0 6.97821e-20 $X=2.377 $Y=2.185
r49 22 24 46.6818 $w=5.05e-07 $l=1.65e-07 $layer=POLY_cond $X=2.432 $Y=1.68
+ $X2=2.432 $Y2=1.515
r50 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.68 $X2=2.52 $Y2=1.68
r51 16 23 14.1075 $w=2.88e-07 $l=3.55e-07 $layer=LI1_cond $X=2.58 $Y=2.035
+ $X2=2.58 $Y2=1.68
r52 15 23 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=2.58 $Y=1.665
+ $X2=2.58 $Y2=1.68
r53 14 15 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.58 $Y=1.295
+ $X2=2.58 $Y2=1.665
r54 13 14 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.58 $Y=0.925
+ $X2=2.58 $Y2=1.295
r55 11 12 45.0926 $w=5.05e-07 $l=1.5e-07 $layer=POLY_cond $X=2.377 $Y=2.035
+ $X2=2.377 $Y2=2.185
r56 9 22 9.21734 $w=5.05e-07 $l=8.7e-08 $layer=POLY_cond $X=2.432 $Y=1.767
+ $X2=2.432 $Y2=1.68
r57 9 11 28.3936 $w=5.05e-07 $l=2.68e-07 $layer=POLY_cond $X=2.432 $Y=1.767
+ $X2=2.432 $Y2=2.035
r58 7 24 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.255 $Y=0.445
+ $X2=2.255 $Y2=1.515
r59 3 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.145 $Y=2.865
+ $X2=2.145 $Y2=2.185
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_M%A4 1 3 6 8 9 10 11 13 16 17 18 19 20 21 28
r43 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=2.035
+ $X2=3.105 $Y2=2.405
r44 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=1.665
+ $X2=3.105 $Y2=2.035
r45 18 19 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=1.295
+ $X2=3.105 $Y2=1.665
r46 17 18 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=0.925
+ $X2=3.105 $Y2=1.295
r47 17 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.005 $X2=3.09 $Y2=1.005
r48 15 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.09 $Y=1.345
+ $X2=3.09 $Y2=1.005
r49 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.345
+ $X2=3.09 $Y2=1.51
r50 14 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.09 $Y=0.99
+ $X2=3.09 $Y2=1.005
r51 13 16 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=3 $Y=2.395 $X2=3
+ $Y2=1.51
r52 10 14 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.925 $Y=0.915
+ $X2=3.09 $Y2=0.99
r53 10 11 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=2.925 $Y=0.915
+ $X2=2.69 $Y2=0.915
r54 8 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.925 $Y=2.47
+ $X2=3 $Y2=2.395
r55 8 9 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=2.925 $Y=2.47
+ $X2=2.65 $Y2=2.47
r56 4 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.615 $Y=0.84
+ $X2=2.69 $Y2=0.915
r57 4 6 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.615 $Y=0.84
+ $X2=2.615 $Y2=0.445
r58 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.575 $Y=2.545
+ $X2=2.65 $Y2=2.47
r59 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.575 $Y=2.545
+ $X2=2.575 $Y2=2.865
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_M%Y 1 2 7 11 13 14 15 16 17 18
c32 11 0 6.12854e-20 $X=1.21 $Y=0.51
c33 7 0 1.47589e-19 $X=1.105 $Y=0.925
r34 18 39 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.295 $Y=2.775
+ $X2=0.295 $Y2=2.8
r35 17 18 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.295 $Y=2.405
+ $X2=0.295 $Y2=2.775
r36 16 17 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.295 $Y=2.035
+ $X2=0.295 $Y2=2.405
r37 15 16 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.295 $Y=1.665
+ $X2=0.295 $Y2=2.035
r38 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.295 $Y=1.295
+ $X2=0.295 $Y2=1.665
r39 13 14 9.27226 $w=4.48e-07 $l=2.85e-07 $layer=LI1_cond $X=0.295 $Y=1.01
+ $X2=0.295 $Y2=1.295
r40 9 11 17.4286 $w=2.08e-07 $l=3.3e-07 $layer=LI1_cond $X=1.21 $Y=0.84 $X2=1.21
+ $Y2=0.51
r41 8 13 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.435 $Y=0.925
+ $X2=0.295 $Y2=0.925
r42 7 9 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.105 $Y=0.925
+ $X2=1.21 $Y2=0.84
r43 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.105 $Y=0.925
+ $X2=0.435 $Y2=0.925
r44 2 39 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=2.655 $X2=0.35 $Y2=2.8
r45 1 11 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.21 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_M%A_186_531# 1 2 3 12 14 15 18 20 22 23
c48 23 0 6.97821e-20 $X=2.79 $Y=2.52
c49 14 0 1.18907e-19 $X=1.825 $Y=2.52
r50 23 25 14.1743 $w=2.41e-07 $l=2.8e-07 $layer=LI1_cond $X=2.79 $Y=2.52
+ $X2=2.79 $Y2=2.8
r51 21 22 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.035 $Y=2.52
+ $X2=1.93 $Y2=2.52
r52 20 23 2.78154 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=2.52
+ $X2=2.79 $Y2=2.52
r53 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.625 $Y=2.52
+ $X2=2.035 $Y2=2.52
r54 16 22 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=2.605
+ $X2=1.93 $Y2=2.52
r55 16 18 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=1.93 $Y=2.605
+ $X2=1.93 $Y2=2.8
r56 14 22 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.825 $Y=2.52
+ $X2=1.93 $Y2=2.52
r57 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.825 $Y=2.52
+ $X2=1.175 $Y2=2.52
r58 10 15 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.08 $Y=2.605
+ $X2=1.175 $Y2=2.52
r59 10 12 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=1.08 $Y=2.605
+ $X2=1.08 $Y2=2.78
r60 3 25 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=2.655 $X2=2.79 $Y2=2.8
r61 2 18 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=2.655 $X2=1.93 $Y2=2.8
r62 1 12 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=2.655 $X2=1.07 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_M%VPWR 1 2 9 13 16 17 19 20 21 34 35
r43 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 19 31 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 19 20 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.35 $Y2=3.33
r54 18 34 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 18 20 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.35 $Y2=3.33
r56 16 28 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.5 $Y2=3.33
r58 15 31 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.605 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.605 $Y=3.33
+ $X2=1.5 $Y2=3.33
r60 11 20 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=3.245
+ $X2=2.35 $Y2=3.33
r61 11 13 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.35 $Y=3.245
+ $X2=2.35 $Y2=2.95
r62 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=3.245 $X2=1.5
+ $Y2=3.33
r63 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.5 $Y=3.245 $X2=1.5
+ $Y2=2.95
r64 2 13 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=2.655 $X2=2.36 $Y2=2.95
r65 1 9 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=2.655 $X2=1.5 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_M%VGND 1 2 11 15 18 19 20 30 31 34
r40 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 28 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r43 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r45 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r46 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 22 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.78
+ $Y2=0
r48 22 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.2
+ $Y2=0
r49 20 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 20 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r51 18 27 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.665 $Y=0 $X2=2.64
+ $Y2=0
r52 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.665 $Y=0 $X2=2.83
+ $Y2=0
r53 17 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.995 $Y=0 $X2=3.12
+ $Y2=0
r54 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.995 $Y=0 $X2=2.83
+ $Y2=0
r55 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.83 $Y=0.085
+ $X2=2.83 $Y2=0
r56 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.83 $Y=0.085
+ $X2=2.83 $Y2=0.38
r57 9 34 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r58 9 11 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.38
r59 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.69
+ $Y=0.235 $X2=2.83 $Y2=0.38
r60 1 11 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.655
+ $Y=0.235 $X2=0.78 $Y2=0.38
.ends

