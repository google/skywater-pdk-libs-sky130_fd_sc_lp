* NGSPICE file created from sky130_fd_sc_lp__o21a_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o21a_0 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_337_483# VPB phighvt w=640000u l=150000u
+  ad=3.84e+11p pd=3.76e+06u as=1.344e+11p ps=1.7e+06u
M1001 a_300_58# A1 VGND VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.289e+11p ps=2.77e+06u
M1002 a_300_58# B1 a_80_23# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 VPWR a_80_23# X VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1004 VGND a_80_23# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 a_337_483# A2 a_80_23# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.144e+11p ps=1.95e+06u
M1006 a_80_23# B1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_300_58# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

