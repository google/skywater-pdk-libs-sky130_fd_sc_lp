* File: sky130_fd_sc_lp__o221a_2.pxi.spice
* Created: Fri Aug 28 11:07:41 2020
* 
x_PM_SKY130_FD_SC_LP__O221A_2%C1 N_C1_c_74_n N_C1_M1001_g N_C1_M1004_g C1 C1
+ N_C1_c_77_n PM_SKY130_FD_SC_LP__O221A_2%C1
x_PM_SKY130_FD_SC_LP__O221A_2%B1 N_B1_M1002_g N_B1_M1012_g B1 N_B1_c_104_n
+ N_B1_c_107_n PM_SKY130_FD_SC_LP__O221A_2%B1
x_PM_SKY130_FD_SC_LP__O221A_2%B2 N_B2_M1005_g N_B2_M1008_g B2 N_B2_c_139_n
+ N_B2_c_140_n PM_SKY130_FD_SC_LP__O221A_2%B2
x_PM_SKY130_FD_SC_LP__O221A_2%A2 N_A2_M1009_g N_A2_c_178_n N_A2_M1003_g A2
+ N_A2_c_179_n N_A2_c_180_n PM_SKY130_FD_SC_LP__O221A_2%A2
x_PM_SKY130_FD_SC_LP__O221A_2%A1 N_A1_c_217_n N_A1_M1010_g N_A1_M1011_g A1
+ N_A1_c_215_n N_A1_c_216_n PM_SKY130_FD_SC_LP__O221A_2%A1
x_PM_SKY130_FD_SC_LP__O221A_2%A_36_67# N_A_36_67#_M1001_s N_A_36_67#_M1004_s
+ N_A_36_67#_M1008_d N_A_36_67#_M1000_g N_A_36_67#_M1007_g N_A_36_67#_M1006_g
+ N_A_36_67#_M1013_g N_A_36_67#_c_253_n N_A_36_67#_c_261_n N_A_36_67#_c_254_n
+ N_A_36_67#_c_283_n N_A_36_67#_c_263_n N_A_36_67#_c_286_n N_A_36_67#_c_295_n
+ N_A_36_67#_c_255_n N_A_36_67#_c_256_n N_A_36_67#_c_291_n N_A_36_67#_c_257_n
+ N_A_36_67#_c_258_n PM_SKY130_FD_SC_LP__O221A_2%A_36_67#
x_PM_SKY130_FD_SC_LP__O221A_2%VPWR N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_M1013_s
+ N_VPWR_c_371_n N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n VPWR
+ N_VPWR_c_375_n N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_370_n
+ PM_SKY130_FD_SC_LP__O221A_2%VPWR
x_PM_SKY130_FD_SC_LP__O221A_2%X N_X_M1000_d N_X_M1007_d N_X_c_448_n N_X_c_430_n
+ X X X X N_X_c_456_p X PM_SKY130_FD_SC_LP__O221A_2%X
x_PM_SKY130_FD_SC_LP__O221A_2%A_119_67# N_A_119_67#_M1001_d N_A_119_67#_M1005_d
+ N_A_119_67#_c_459_n N_A_119_67#_c_460_n N_A_119_67#_c_461_n
+ PM_SKY130_FD_SC_LP__O221A_2%A_119_67#
x_PM_SKY130_FD_SC_LP__O221A_2%A_205_67# N_A_205_67#_M1002_d N_A_205_67#_M1003_d
+ N_A_205_67#_c_486_n N_A_205_67#_c_483_n N_A_205_67#_c_484_n
+ N_A_205_67#_c_507_p PM_SKY130_FD_SC_LP__O221A_2%A_205_67#
x_PM_SKY130_FD_SC_LP__O221A_2%VGND N_VGND_M1003_s N_VGND_M1011_d N_VGND_M1006_s
+ N_VGND_c_510_n N_VGND_c_511_n N_VGND_c_512_n N_VGND_c_513_n VGND
+ N_VGND_c_514_n N_VGND_c_515_n N_VGND_c_516_n N_VGND_c_517_n N_VGND_c_518_n
+ N_VGND_c_519_n PM_SKY130_FD_SC_LP__O221A_2%VGND
cc_1 VNB N_C1_c_74_n 0.0204296f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.285
cc_2 VNB N_C1_M1004_g 0.00186281f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.465
cc_3 VNB C1 0.0213666f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_C1_c_77_n 0.0513853f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.45
cc_5 VNB N_B1_M1002_g 0.0207577f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.755
cc_6 VNB B1 0.00296594f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_B1_c_104_n 0.0256032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B2_M1005_g 0.0231128f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.755
cc_9 VNB N_B2_c_139_n 0.0256991f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.45
cc_10 VNB N_B2_c_140_n 0.00281736f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.45
cc_11 VNB N_A2_M1009_g 0.00309437f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.755
cc_12 VNB N_A2_c_178_n 0.0198997f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.465
cc_13 VNB N_A2_c_179_n 0.00257427f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.45
cc_14 VNB N_A2_c_180_n 0.0525762f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.45
cc_15 VNB N_A1_M1011_g 0.0259583f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.465
cc_16 VNB N_A1_c_215_n 0.033493f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.45
cc_17 VNB N_A1_c_216_n 0.00286714f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.45
cc_18 VNB N_A_36_67#_M1000_g 0.0247603f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.45
cc_19 VNB N_A_36_67#_M1006_g 0.0292438f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=1.45
cc_20 VNB N_A_36_67#_c_253_n 0.0229417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_36_67#_c_254_n 0.00344383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_36_67#_c_255_n 4.69546e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_36_67#_c_256_n 0.00731496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_36_67#_c_257_n 0.00389874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_36_67#_c_258_n 0.0351178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_370_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0163237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB X 0.0200259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_119_67#_c_459_n 0.00653972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_119_67#_c_460_n 0.00388037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_119_67#_c_461_n 0.00202279f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.45
cc_32 VNB N_A_205_67#_c_483_n 0.0210536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_510_n 0.00840949f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.45
cc_34 VNB N_VGND_c_511_n 0.0101453f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.45
cc_35 VNB N_VGND_c_512_n 0.0132347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_513_n 0.0302429f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=1.45
cc_37 VNB N_VGND_c_514_n 0.0522368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_515_n 0.0166635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_516_n 0.0165512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_517_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_518_n 0.00471252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_519_n 0.249323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_C1_M1004_g 0.0251702f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.465
cc_44 VPB C1 0.0100043f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_45 VPB B1 0.0033264f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_46 VPB N_B1_c_104_n 0.00903024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B1_c_107_n 0.0167275f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.45
cc_48 VPB N_B2_M1008_g 0.0215202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B2_c_139_n 0.00584832f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.45
cc_50 VPB N_B2_c_140_n 0.00318504f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.45
cc_51 VPB N_A2_M1009_g 0.0213802f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=0.755
cc_52 VPB N_A2_c_179_n 0.00373017f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.45
cc_53 VPB N_A1_c_217_n 0.017805f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.285
cc_54 VPB N_A1_c_215_n 0.0163611f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.45
cc_55 VPB N_A1_c_216_n 0.0029307f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.45
cc_56 VPB N_A_36_67#_M1007_g 0.020007f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.45
cc_57 VPB N_A_36_67#_M1013_g 0.0221304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_36_67#_c_261_n 0.0379094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_36_67#_c_254_n 0.00145303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_36_67#_c_263_n 0.00746105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_36_67#_c_255_n 0.00158728f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_36_67#_c_258_n 0.00490605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_371_n 0.0055721f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.45
cc_64 VPB N_VPWR_c_372_n 0.00183337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_373_n 0.0120942f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=1.45
cc_66 VPB N_VPWR_c_374_n 0.0388867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_375_n 0.0445513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_376_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_377_n 0.0265594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_378_n 0.0104351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_370_n 0.0503568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_X_c_430_n 0.0129964f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.45
cc_73 VPB X 0.00823407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 N_C1_c_74_n N_B1_M1002_g 0.0315096f $X=0.52 $Y=1.285 $X2=0 $Y2=0
cc_75 N_C1_c_77_n B1 3.66737e-19 $X=0.52 $Y=1.45 $X2=0 $Y2=0
cc_76 N_C1_c_77_n N_B1_c_104_n 0.021787f $X=0.52 $Y=1.45 $X2=0 $Y2=0
cc_77 N_C1_M1004_g N_B1_c_107_n 0.0215513f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_78 N_C1_c_74_n N_A_36_67#_c_253_n 0.00189935f $X=0.52 $Y=1.285 $X2=0 $Y2=0
cc_79 N_C1_M1004_g N_A_36_67#_c_261_n 0.0130462f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_80 N_C1_c_74_n N_A_36_67#_c_254_n 0.0103906f $X=0.52 $Y=1.285 $X2=0 $Y2=0
cc_81 N_C1_M1004_g N_A_36_67#_c_254_n 0.0122342f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_82 C1 N_A_36_67#_c_254_n 0.0396883f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_C1_c_77_n N_A_36_67#_c_254_n 0.00914022f $X=0.52 $Y=1.45 $X2=0 $Y2=0
cc_84 N_C1_M1004_g N_A_36_67#_c_263_n 0.0140797f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_85 C1 N_A_36_67#_c_263_n 0.0158959f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_C1_c_77_n N_A_36_67#_c_263_n 0.00381667f $X=0.52 $Y=1.45 $X2=0 $Y2=0
cc_87 N_C1_c_74_n N_A_36_67#_c_256_n 0.0112649f $X=0.52 $Y=1.285 $X2=0 $Y2=0
cc_88 C1 N_A_36_67#_c_256_n 0.0183859f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_C1_c_77_n N_A_36_67#_c_256_n 0.00287516f $X=0.52 $Y=1.45 $X2=0 $Y2=0
cc_90 N_C1_M1004_g N_VPWR_c_371_n 0.00430884f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_91 N_C1_M1004_g N_VPWR_c_377_n 0.00571722f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_92 N_C1_M1004_g N_VPWR_c_370_n 0.0115517f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_93 N_C1_c_74_n N_A_119_67#_c_461_n 0.00840678f $X=0.52 $Y=1.285 $X2=0 $Y2=0
cc_94 N_C1_c_74_n N_VGND_c_514_n 0.0045977f $X=0.52 $Y=1.285 $X2=0 $Y2=0
cc_95 N_C1_c_74_n N_VGND_c_519_n 0.00544919f $X=0.52 $Y=1.285 $X2=0 $Y2=0
cc_96 N_B1_M1002_g N_B2_M1005_g 0.0241897f $X=0.95 $Y=0.755 $X2=0 $Y2=0
cc_97 N_B1_c_107_n N_B2_M1008_g 0.0569516f $X=1.01 $Y=1.72 $X2=0 $Y2=0
cc_98 B1 N_B2_c_139_n 0.00292189f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_99 N_B1_c_104_n N_B2_c_139_n 0.0569516f $X=1.01 $Y=1.51 $X2=0 $Y2=0
cc_100 B1 N_B2_c_140_n 0.032719f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_101 N_B1_c_104_n N_B2_c_140_n 3.51315e-19 $X=1.01 $Y=1.51 $X2=0 $Y2=0
cc_102 N_B1_c_107_n N_A_36_67#_c_261_n 7.22817e-19 $X=1.01 $Y=1.72 $X2=0 $Y2=0
cc_103 N_B1_M1002_g N_A_36_67#_c_254_n 0.00480729f $X=0.95 $Y=0.755 $X2=0 $Y2=0
cc_104 B1 N_A_36_67#_c_254_n 0.0318797f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_105 N_B1_c_104_n N_A_36_67#_c_254_n 0.00222227f $X=1.01 $Y=1.51 $X2=0 $Y2=0
cc_106 N_B1_c_107_n N_A_36_67#_c_254_n 0.00323727f $X=1.01 $Y=1.72 $X2=0 $Y2=0
cc_107 B1 N_A_36_67#_c_283_n 0.0274216f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_B1_c_104_n N_A_36_67#_c_283_n 0.00225117f $X=1.01 $Y=1.51 $X2=0 $Y2=0
cc_109 N_B1_c_107_n N_A_36_67#_c_283_n 0.0150921f $X=1.01 $Y=1.72 $X2=0 $Y2=0
cc_110 N_B1_c_107_n N_A_36_67#_c_286_n 0.00308489f $X=1.01 $Y=1.72 $X2=0 $Y2=0
cc_111 N_B1_M1002_g N_A_36_67#_c_256_n 0.00153496f $X=0.95 $Y=0.755 $X2=0 $Y2=0
cc_112 N_B1_c_107_n N_VPWR_c_371_n 0.00430884f $X=1.01 $Y=1.72 $X2=0 $Y2=0
cc_113 N_B1_c_107_n N_VPWR_c_375_n 0.00585385f $X=1.01 $Y=1.72 $X2=0 $Y2=0
cc_114 N_B1_c_107_n N_VPWR_c_370_n 0.0107844f $X=1.01 $Y=1.72 $X2=0 $Y2=0
cc_115 N_B1_M1002_g N_A_119_67#_c_459_n 0.0111471f $X=0.95 $Y=0.755 $X2=0 $Y2=0
cc_116 N_B1_M1002_g N_A_119_67#_c_461_n 0.00761661f $X=0.95 $Y=0.755 $X2=0 $Y2=0
cc_117 B1 N_A_119_67#_c_461_n 3.55206e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_118 B1 N_A_205_67#_c_484_n 0.0178256f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_119 N_B1_c_104_n N_A_205_67#_c_484_n 0.00279068f $X=1.01 $Y=1.51 $X2=0 $Y2=0
cc_120 N_B1_M1002_g N_VGND_c_514_n 0.00298199f $X=0.95 $Y=0.755 $X2=0 $Y2=0
cc_121 N_B1_M1002_g N_VGND_c_519_n 0.00422879f $X=0.95 $Y=0.755 $X2=0 $Y2=0
cc_122 N_B2_M1008_g N_A2_M1009_g 0.00686027f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B2_c_139_n N_A2_M1009_g 0.00190368f $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_124 N_B2_c_140_n N_A2_M1009_g 4.52855e-19 $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_125 N_B2_M1008_g N_A2_c_179_n 4.06124e-19 $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B2_c_139_n N_A2_c_179_n 5.29809e-19 $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_127 N_B2_c_140_n N_A2_c_179_n 0.034084f $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_128 N_B2_M1005_g N_A2_c_180_n 0.0053678f $X=1.46 $Y=0.755 $X2=0 $Y2=0
cc_129 N_B2_c_139_n N_A2_c_180_n 0.0121868f $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_130 N_B2_c_140_n N_A2_c_180_n 0.00157844f $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_131 N_B2_M1008_g N_A_36_67#_c_283_n 0.0131379f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_132 N_B2_c_140_n N_A_36_67#_c_283_n 0.00304003f $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_133 N_B2_M1008_g N_A_36_67#_c_286_n 0.0191717f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B2_M1008_g N_A_36_67#_c_291_n 7.41524e-19 $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_135 N_B2_c_139_n N_A_36_67#_c_291_n 9.92943e-19 $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_136 N_B2_c_140_n N_A_36_67#_c_291_n 0.0222943f $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_137 N_B2_M1008_g N_VPWR_c_375_n 0.0054895f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_138 N_B2_M1008_g N_VPWR_c_370_n 0.0104939f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_139 N_B2_M1005_g N_A_119_67#_c_459_n 0.0128389f $X=1.46 $Y=0.755 $X2=0 $Y2=0
cc_140 N_B2_M1005_g N_A_119_67#_c_461_n 3.57018e-19 $X=1.46 $Y=0.755 $X2=0 $Y2=0
cc_141 N_B2_M1005_g N_A_205_67#_c_486_n 0.00966294f $X=1.46 $Y=0.755 $X2=0 $Y2=0
cc_142 N_B2_M1005_g N_A_205_67#_c_483_n 0.0135436f $X=1.46 $Y=0.755 $X2=0 $Y2=0
cc_143 N_B2_c_139_n N_A_205_67#_c_483_n 0.00394418f $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_144 N_B2_c_140_n N_A_205_67#_c_483_n 0.0236723f $X=1.55 $Y=1.5 $X2=0 $Y2=0
cc_145 N_B2_M1005_g N_A_205_67#_c_484_n 8.855e-19 $X=1.46 $Y=0.755 $X2=0 $Y2=0
cc_146 N_B2_M1005_g N_VGND_c_510_n 0.00220476f $X=1.46 $Y=0.755 $X2=0 $Y2=0
cc_147 N_B2_M1005_g N_VGND_c_514_n 0.00296932f $X=1.46 $Y=0.755 $X2=0 $Y2=0
cc_148 N_B2_M1005_g N_VGND_c_519_n 0.00463001f $X=1.46 $Y=0.755 $X2=0 $Y2=0
cc_149 N_A2_M1009_g N_A1_c_217_n 0.0499504f $X=2.23 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A2_c_178_n N_A1_M1011_g 0.0184954f $X=2.41 $Y=1.185 $X2=0 $Y2=0
cc_151 N_A2_c_179_n N_A1_c_215_n 0.00180555f $X=2.14 $Y=1.42 $X2=0 $Y2=0
cc_152 N_A2_c_180_n N_A1_c_215_n 0.0566172f $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_153 N_A2_c_179_n N_A1_c_216_n 0.0348073f $X=2.14 $Y=1.42 $X2=0 $Y2=0
cc_154 N_A2_c_180_n N_A1_c_216_n 9.51741e-19 $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_155 N_A2_M1009_g N_A_36_67#_c_286_n 0.0193517f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A2_M1009_g N_A_36_67#_c_295_n 0.00953771f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A2_c_179_n N_A_36_67#_c_295_n 0.0114625f $X=2.14 $Y=1.42 $X2=0 $Y2=0
cc_158 N_A2_c_180_n N_A_36_67#_c_295_n 0.0028079f $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_159 N_A2_M1009_g N_A_36_67#_c_291_n 0.00118794f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A2_c_179_n N_A_36_67#_c_291_n 0.0165405f $X=2.14 $Y=1.42 $X2=0 $Y2=0
cc_161 N_A2_c_180_n N_A_36_67#_c_291_n 8.12452e-19 $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_162 N_A2_M1009_g N_VPWR_c_372_n 0.00345882f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A2_M1009_g N_VPWR_c_375_n 0.00526178f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A2_M1009_g N_VPWR_c_370_n 0.009938f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A2_c_178_n N_A_205_67#_c_483_n 0.0183288f $X=2.41 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A2_c_179_n N_A_205_67#_c_483_n 0.0304993f $X=2.14 $Y=1.42 $X2=0 $Y2=0
cc_167 N_A2_c_180_n N_A_205_67#_c_483_n 0.0104406f $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_168 N_A2_c_178_n N_VGND_c_510_n 0.0114766f $X=2.41 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A2_c_178_n N_VGND_c_515_n 0.00486043f $X=2.41 $Y=1.185 $X2=0 $Y2=0
cc_170 N_A2_c_178_n N_VGND_c_519_n 0.0084429f $X=2.41 $Y=1.185 $X2=0 $Y2=0
cc_171 N_A1_M1011_g N_A_36_67#_M1000_g 0.0244283f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_172 N_A1_c_217_n N_A_36_67#_M1007_g 0.0107307f $X=2.59 $Y=1.725 $X2=0 $Y2=0
cc_173 N_A1_c_215_n N_A_36_67#_M1007_g 0.00238922f $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_174 N_A1_c_217_n N_A_36_67#_c_286_n 0.00309794f $X=2.59 $Y=1.725 $X2=0 $Y2=0
cc_175 N_A1_c_217_n N_A_36_67#_c_295_n 0.0159329f $X=2.59 $Y=1.725 $X2=0 $Y2=0
cc_176 N_A1_c_215_n N_A_36_67#_c_295_n 0.00441718f $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A1_c_216_n N_A_36_67#_c_295_n 0.0296915f $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_178 N_A1_c_217_n N_A_36_67#_c_255_n 0.00291459f $X=2.59 $Y=1.725 $X2=0 $Y2=0
cc_179 N_A1_c_215_n N_A_36_67#_c_255_n 5.73844e-19 $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A1_c_216_n N_A_36_67#_c_255_n 0.00889828f $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_181 N_A1_c_215_n N_A_36_67#_c_257_n 0.00175819f $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A1_c_216_n N_A_36_67#_c_257_n 0.0198851f $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A1_c_215_n N_A_36_67#_c_258_n 0.0175871f $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_184 N_A1_c_216_n N_A_36_67#_c_258_n 6.11811e-19 $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_185 N_A1_c_217_n N_VPWR_c_372_n 0.0227522f $X=2.59 $Y=1.725 $X2=0 $Y2=0
cc_186 N_A1_c_217_n N_VPWR_c_375_n 0.00486043f $X=2.59 $Y=1.725 $X2=0 $Y2=0
cc_187 N_A1_c_217_n N_VPWR_c_370_n 0.00818711f $X=2.59 $Y=1.725 $X2=0 $Y2=0
cc_188 N_A1_M1011_g N_A_205_67#_c_483_n 0.00147518f $X=2.915 $Y=0.655 $X2=0
+ $Y2=0
cc_189 N_A1_c_215_n N_A_205_67#_c_483_n 0.00519514f $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A1_c_216_n N_A_205_67#_c_483_n 0.0248535f $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A1_M1011_g N_VGND_c_510_n 5.84979e-19 $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A1_M1011_g N_VGND_c_511_n 0.00252456f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A1_c_215_n N_VGND_c_511_n 5.79492e-19 $X=2.86 $Y=1.51 $X2=0 $Y2=0
cc_194 N_A1_M1011_g N_VGND_c_515_n 0.00585385f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A1_M1011_g N_VGND_c_519_n 0.0107707f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A_36_67#_c_254_n N_VPWR_M1004_d 0.00129763f $X=0.63 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_197 N_A_36_67#_c_283_n N_VPWR_M1004_d 0.0090618f $X=1.51 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_36_67#_c_263_n N_VPWR_M1004_d 2.98916e-19 $X=0.715 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A_36_67#_c_295_n N_VPWR_M1010_d 0.01439f $X=3.125 $Y=2.015 $X2=0 $Y2=0
cc_200 N_A_36_67#_c_255_n N_VPWR_M1010_d 0.00139749f $X=3.21 $Y=1.93 $X2=0 $Y2=0
cc_201 N_A_36_67#_c_263_n N_VPWR_c_371_n 0.022382f $X=0.715 $Y=2.015 $X2=0 $Y2=0
cc_202 N_A_36_67#_M1007_g N_VPWR_c_372_n 0.0172839f $X=3.36 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A_36_67#_M1013_g N_VPWR_c_372_n 6.90597e-19 $X=3.79 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_A_36_67#_c_286_n N_VPWR_c_372_n 0.030927f $X=1.675 $Y=2.91 $X2=0 $Y2=0
cc_205 N_A_36_67#_c_295_n N_VPWR_c_372_n 0.0442519f $X=3.125 $Y=2.015 $X2=0
+ $Y2=0
cc_206 N_A_36_67#_c_257_n N_VPWR_c_372_n 3.97649e-19 $X=3.435 $Y=1.51 $X2=0
+ $Y2=0
cc_207 N_A_36_67#_M1007_g N_VPWR_c_374_n 7.07368e-19 $X=3.36 $Y=2.465 $X2=0
+ $Y2=0
cc_208 N_A_36_67#_M1013_g N_VPWR_c_374_n 0.0145851f $X=3.79 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A_36_67#_c_286_n N_VPWR_c_375_n 0.0438525f $X=1.675 $Y=2.91 $X2=0 $Y2=0
cc_210 N_A_36_67#_M1007_g N_VPWR_c_376_n 0.00486043f $X=3.36 $Y=2.465 $X2=0
+ $Y2=0
cc_211 N_A_36_67#_M1013_g N_VPWR_c_376_n 0.00486043f $X=3.79 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_A_36_67#_c_261_n N_VPWR_c_377_n 0.0200241f $X=0.345 $Y=2.91 $X2=0 $Y2=0
cc_213 N_A_36_67#_M1004_s N_VPWR_c_370_n 0.00215158f $X=0.22 $Y=1.835 $X2=0
+ $Y2=0
cc_214 N_A_36_67#_M1008_d N_VPWR_c_370_n 0.00505717f $X=1.535 $Y=1.835 $X2=0
+ $Y2=0
cc_215 N_A_36_67#_M1007_g N_VPWR_c_370_n 0.00824727f $X=3.36 $Y=2.465 $X2=0
+ $Y2=0
cc_216 N_A_36_67#_M1013_g N_VPWR_c_370_n 0.00824727f $X=3.79 $Y=2.465 $X2=0
+ $Y2=0
cc_217 N_A_36_67#_c_261_n N_VPWR_c_370_n 0.0120544f $X=0.345 $Y=2.91 $X2=0 $Y2=0
cc_218 N_A_36_67#_c_286_n N_VPWR_c_370_n 0.0261188f $X=1.675 $Y=2.91 $X2=0 $Y2=0
cc_219 N_A_36_67#_c_283_n A_235_367# 0.0055934f $X=1.51 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_220 N_A_36_67#_c_295_n A_461_367# 0.00518203f $X=3.125 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_221 N_A_36_67#_M1013_g N_X_c_430_n 0.0136693f $X=3.79 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A_36_67#_c_255_n N_X_c_430_n 0.00438446f $X=3.21 $Y=1.93 $X2=0 $Y2=0
cc_223 N_A_36_67#_c_257_n N_X_c_430_n 0.00880481f $X=3.435 $Y=1.51 $X2=0 $Y2=0
cc_224 N_A_36_67#_c_258_n N_X_c_430_n 0.00249365f $X=3.775 $Y=1.51 $X2=0 $Y2=0
cc_225 N_A_36_67#_M1000_g X 0.00368371f $X=3.345 $Y=0.655 $X2=0 $Y2=0
cc_226 N_A_36_67#_M1006_g X 0.0161967f $X=3.775 $Y=0.655 $X2=0 $Y2=0
cc_227 N_A_36_67#_c_257_n X 0.0128405f $X=3.435 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A_36_67#_c_258_n X 0.00258131f $X=3.775 $Y=1.51 $X2=0 $Y2=0
cc_229 N_A_36_67#_M1000_g X 5.88199e-19 $X=3.345 $Y=0.655 $X2=0 $Y2=0
cc_230 N_A_36_67#_M1007_g X 4.59752e-19 $X=3.36 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_36_67#_M1006_g X 0.00506217f $X=3.775 $Y=0.655 $X2=0 $Y2=0
cc_232 N_A_36_67#_M1013_g X 0.00615477f $X=3.79 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A_36_67#_c_255_n X 0.00536827f $X=3.21 $Y=1.93 $X2=0 $Y2=0
cc_234 N_A_36_67#_c_257_n X 0.0189016f $X=3.435 $Y=1.51 $X2=0 $Y2=0
cc_235 N_A_36_67#_c_258_n X 0.0169721f $X=3.775 $Y=1.51 $X2=0 $Y2=0
cc_236 N_A_36_67#_c_254_n N_A_119_67#_M1001_d 0.00182196f $X=0.63 $Y=1.93
+ $X2=-0.19 $Y2=-0.245
cc_237 N_A_36_67#_c_256_n N_A_119_67#_M1001_d 0.00281669f $X=0.63 $Y=0.945
+ $X2=-0.19 $Y2=-0.245
cc_238 N_A_36_67#_c_253_n N_A_119_67#_c_461_n 0.0148334f $X=0.305 $Y=0.48 $X2=0
+ $Y2=0
cc_239 N_A_36_67#_c_256_n N_A_119_67#_c_461_n 0.00652572f $X=0.63 $Y=0.945 $X2=0
+ $Y2=0
cc_240 N_A_36_67#_M1000_g N_A_205_67#_c_483_n 2.04885e-19 $X=3.345 $Y=0.655
+ $X2=0 $Y2=0
cc_241 N_A_36_67#_M1000_g N_VGND_c_511_n 0.00249047f $X=3.345 $Y=0.655 $X2=0
+ $Y2=0
cc_242 N_A_36_67#_c_257_n N_VGND_c_511_n 0.00734429f $X=3.435 $Y=1.51 $X2=0
+ $Y2=0
cc_243 N_A_36_67#_M1006_g N_VGND_c_513_n 0.00347541f $X=3.775 $Y=0.655 $X2=0
+ $Y2=0
cc_244 N_A_36_67#_c_253_n N_VGND_c_514_n 0.01317f $X=0.305 $Y=0.48 $X2=0 $Y2=0
cc_245 N_A_36_67#_M1000_g N_VGND_c_516_n 0.00585385f $X=3.345 $Y=0.655 $X2=0
+ $Y2=0
cc_246 N_A_36_67#_M1006_g N_VGND_c_516_n 0.00585385f $X=3.775 $Y=0.655 $X2=0
+ $Y2=0
cc_247 N_A_36_67#_M1000_g N_VGND_c_519_n 0.0105614f $X=3.345 $Y=0.655 $X2=0
+ $Y2=0
cc_248 N_A_36_67#_M1006_g N_VGND_c_519_n 0.0115011f $X=3.775 $Y=0.655 $X2=0
+ $Y2=0
cc_249 N_A_36_67#_c_253_n N_VGND_c_519_n 0.00965782f $X=0.305 $Y=0.48 $X2=0
+ $Y2=0
cc_250 N_A_36_67#_c_256_n N_VGND_c_519_n 0.00511012f $X=0.63 $Y=0.945 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_370_n A_235_367# 0.00899413f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_252 N_VPWR_c_370_n A_461_367# 0.00899413f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_253 N_VPWR_c_370_n N_X_M1007_d 0.00536646f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_254 N_VPWR_c_376_n N_X_c_448_n 0.0124525f $X=3.84 $Y=3.33 $X2=0 $Y2=0
cc_255 N_VPWR_c_370_n N_X_c_448_n 0.00730901f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_M1013_s N_X_c_430_n 0.00296578f $X=3.865 $Y=1.835 $X2=0 $Y2=0
cc_257 N_VPWR_c_374_n N_X_c_430_n 0.021083f $X=4.005 $Y=2.25 $X2=0 $Y2=0
cc_258 X N_A_205_67#_c_483_n 0.00242112f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_259 X N_VGND_M1006_s 0.00225342f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_260 X N_VGND_c_511_n 0.00164453f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_261 X N_VGND_c_513_n 0.0202165f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_262 N_X_c_456_p N_VGND_c_516_n 0.0149362f $X=3.56 $Y=0.42 $X2=0 $Y2=0
cc_263 N_X_M1000_d N_VGND_c_519_n 0.00293134f $X=3.42 $Y=0.235 $X2=0 $Y2=0
cc_264 N_X_c_456_p N_VGND_c_519_n 0.0100304f $X=3.56 $Y=0.42 $X2=0 $Y2=0
cc_265 N_A_119_67#_c_459_n N_A_205_67#_M1002_d 0.00261503f $X=1.57 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_266 N_A_119_67#_c_459_n N_A_205_67#_c_486_n 0.0194194f $X=1.57 $Y=0.34 $X2=0
+ $Y2=0
cc_267 N_A_119_67#_M1005_d N_A_205_67#_c_483_n 0.00488814f $X=1.535 $Y=0.335
+ $X2=0 $Y2=0
cc_268 N_A_119_67#_c_459_n N_A_205_67#_c_483_n 0.00336661f $X=1.57 $Y=0.34 $X2=0
+ $Y2=0
cc_269 N_A_119_67#_c_460_n N_A_205_67#_c_483_n 0.0199277f $X=1.675 $Y=0.66 $X2=0
+ $Y2=0
cc_270 N_A_119_67#_c_459_n N_VGND_c_510_n 0.0139f $X=1.57 $Y=0.34 $X2=0 $Y2=0
cc_271 N_A_119_67#_c_460_n N_VGND_c_510_n 0.0303028f $X=1.675 $Y=0.66 $X2=0
+ $Y2=0
cc_272 N_A_119_67#_c_459_n N_VGND_c_514_n 0.061432f $X=1.57 $Y=0.34 $X2=0 $Y2=0
cc_273 N_A_119_67#_c_461_n N_VGND_c_514_n 0.0225828f $X=0.735 $Y=0.34 $X2=0
+ $Y2=0
cc_274 N_A_119_67#_c_459_n N_VGND_c_519_n 0.0343843f $X=1.57 $Y=0.34 $X2=0 $Y2=0
cc_275 N_A_119_67#_c_461_n N_VGND_c_519_n 0.0123883f $X=0.735 $Y=0.34 $X2=0
+ $Y2=0
cc_276 N_A_205_67#_c_483_n N_VGND_M1003_s 0.00258276f $X=2.53 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_277 N_A_205_67#_c_483_n N_VGND_c_510_n 0.0220024f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_278 N_A_205_67#_c_483_n N_VGND_c_511_n 0.00533334f $X=2.53 $Y=1.08 $X2=0
+ $Y2=0
cc_279 N_A_205_67#_c_507_p N_VGND_c_515_n 0.0193226f $X=2.68 $Y=0.42 $X2=0 $Y2=0
cc_280 N_A_205_67#_M1003_d N_VGND_c_519_n 0.00440415f $X=2.485 $Y=0.235 $X2=0
+ $Y2=0
cc_281 N_A_205_67#_c_507_p N_VGND_c_519_n 0.0119743f $X=2.68 $Y=0.42 $X2=0 $Y2=0
