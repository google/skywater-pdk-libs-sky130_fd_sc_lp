* File: sky130_fd_sc_lp__buf_1.spice
* Created: Wed Sep  2 09:34:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__buf_1.pex.spice"
.subckt sky130_fd_sc_lp__buf_1  VNB VPB A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_70_237#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1694 AS=0.2226 PD=1.57333 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.4 A=0.126 P=1.98 MULT=1
MM1002 N_A_70_237#_M1002_d N_A_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0847 PD=1.37 PS=0.786667 NRD=0 NRS=41.904 M=1 R=2.8 SA=75000.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_70_237#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.25326 AS=0.3339 PD=2.12211 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.4 A=0.189 P=2.82 MULT=1
MM1000 N_A_70_237#_M1000_d N_A_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.12864 PD=1.81 PS=1.07789 NRD=0 NRS=19.2272 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__buf_1.pxi.spice"
*
.ends
*
*
