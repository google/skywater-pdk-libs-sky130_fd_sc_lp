* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_942_252# a_591_155# a_1184_60# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND a_942_252# a_1555_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_508_155# a_392_144# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_942_252# a_606_359# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND GATE_N a_113_144# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_942_252# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 Q_N a_1555_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VPWR a_1555_367# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR a_591_155# a_942_252# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND a_1555_367# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_591_155# a_162_40# a_677_155# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR GATE_N a_113_144# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_591_155# a_162_40# a_794_359# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_794_359# a_392_144# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VGND a_942_252# a_677_155# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 Q a_942_252# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_162_40# a_113_144# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_942_252# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_508_155# a_113_144# a_591_155# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1184_60# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 Q_N a_1555_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_606_359# a_113_144# a_591_155# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VGND a_942_252# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 Q a_942_252# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VGND D a_392_144# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_162_40# a_113_144# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 VPWR D a_392_144# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 VPWR a_942_252# a_1555_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
