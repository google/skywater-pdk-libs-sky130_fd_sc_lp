* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__iso1n_lp A KAGND SLEEP_B VGND VNB VPB VPWR X
X0 a_27_93# SLEEP_B a_110_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_438_93# A KAGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_340_93# A a_438_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_27_93# SLEEP_B a_154_489# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_340_489# A a_340_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 KAGND a_27_93# a_268_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 KAGND a_340_93# a_602_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_268_93# a_27_93# a_340_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_27_93# a_340_489# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR a_340_93# a_602_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_602_367# a_340_93# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_154_489# SLEEP_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_602_93# a_340_93# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_110_93# SLEEP_B KAGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
