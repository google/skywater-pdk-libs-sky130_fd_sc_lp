* File: sky130_fd_sc_lp__maj3_m.pex.spice
* Created: Wed Sep  2 09:59:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MAJ3_M%A 3 7 11 15 17 18 22
r37 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=1.07 $X2=1.16 $Y2=1.07
r38 18 23 0.714077 $w=6.68e-07 $l=4e-08 $layer=LI1_cond $X=1.2 $Y=1.24 $X2=1.16
+ $Y2=1.24
r39 17 23 7.85484 $w=6.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.72 $Y=1.24
+ $X2=1.16 $Y2=1.24
r40 13 22 86.458 $w=2.9e-07 $l=6.02993e-07 $layer=POLY_cond $X=1.35 $Y=1.575
+ $X2=1.135 $Y2=1.07
r41 13 15 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.35 $Y=1.575
+ $X2=1.35 $Y2=2.335
r42 9 22 29.9477 $w=2.9e-07 $l=2.85832e-07 $layer=POLY_cond $X=1.35 $Y=0.905
+ $X2=1.135 $Y2=1.07
r43 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.35 $Y=0.905
+ $X2=1.35 $Y2=0.495
r44 5 22 86.458 $w=2.9e-07 $l=6.02993e-07 $layer=POLY_cond $X=0.92 $Y=1.575
+ $X2=1.135 $Y2=1.07
r45 5 7 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.92 $Y=1.575 $X2=0.92
+ $Y2=2.335
r46 1 22 29.9477 $w=2.9e-07 $l=2.15e-07 $layer=POLY_cond $X=0.92 $Y=1.07
+ $X2=1.135 $Y2=1.07
r47 1 3 210.234 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.92 $Y=1.07 $X2=0.92
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_M%B 3 7 11 15 17 18 22
c44 3 0 2.1014e-20 $X=1.74 $Y=0.495
r45 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.83
+ $Y=1.07 $X2=1.83 $Y2=1.07
r46 18 23 5.89113 $w=6.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.16 $Y=1.24
+ $X2=1.83 $Y2=1.24
r47 17 23 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.68 $Y=1.24
+ $X2=1.83 $Y2=1.24
r48 13 22 86.458 $w=2.9e-07 $l=6.02993e-07 $layer=POLY_cond $X=2.17 $Y=1.575
+ $X2=1.955 $Y2=1.07
r49 13 15 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.17 $Y=1.575
+ $X2=2.17 $Y2=2.335
r50 9 22 29.9477 $w=2.9e-07 $l=2.85832e-07 $layer=POLY_cond $X=2.17 $Y=0.905
+ $X2=1.955 $Y2=1.07
r51 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.17 $Y=0.905
+ $X2=2.17 $Y2=0.495
r52 5 22 86.458 $w=2.9e-07 $l=6.02993e-07 $layer=POLY_cond $X=1.74 $Y=1.575
+ $X2=1.955 $Y2=1.07
r53 5 7 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.74 $Y=1.575 $X2=1.74
+ $Y2=2.335
r54 1 22 29.9477 $w=2.9e-07 $l=2.15e-07 $layer=POLY_cond $X=1.74 $Y=1.07
+ $X2=1.955 $Y2=1.07
r55 1 3 210.234 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.74 $Y=1.07 $X2=1.74
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_M%C 3 6 7 8 11 14 15 16 20
r54 20 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.62 $Y=2.9 $X2=2.62
+ $Y2=2.99
r55 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=2.9
+ $X2=2.62 $Y2=2.735
r56 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=2.9 $X2=2.62 $Y2=2.9
r57 16 21 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.62 $Y=2.775
+ $X2=2.62 $Y2=2.9
r58 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.405
+ $X2=2.62 $Y2=2.775
r59 14 22 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.56 $Y=2.335 $X2=2.56
+ $Y2=2.735
r60 11 14 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=2.56 $Y=0.495
+ $X2=2.56 $Y2=2.335
r61 7 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.455 $Y=2.99
+ $X2=2.62 $Y2=2.99
r62 7 8 948.617 $w=1.5e-07 $l=1.85e-06 $layer=POLY_cond $X=2.455 $Y=2.99
+ $X2=0.605 $Y2=2.99
r63 3 6 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=0.53 $Y=0.495
+ $X2=0.53 $Y2=2.335
r64 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.53 $Y=2.915
+ $X2=0.605 $Y2=2.99
r65 1 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.53 $Y=2.915 $X2=0.53
+ $Y2=2.335
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_M%A_34_57# 1 2 3 4 17 21 23 24 26 29 31 35 37
+ 39 42 43 47 48 51 54 56 60 61
c100 37 0 2.1014e-20 $X=2.455 $Y=0.64
r101 56 58 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.955 $Y=0.495
+ $X2=1.955 $Y2=0.64
r102 51 53 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.315 $Y=0.495
+ $X2=0.315 $Y2=0.725
r103 48 63 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=3.112 $Y=1.42
+ $X2=3.112 $Y2=1.255
r104 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.05
+ $Y=1.42 $X2=3.05 $Y2=1.42
r105 45 47 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.05 $Y=1.755
+ $X2=3.05 $Y2=1.42
r106 44 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=1.84
+ $X2=2.54 $Y2=1.84
r107 43 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.885 $Y=1.84
+ $X2=3.05 $Y2=1.755
r108 43 44 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.885 $Y=1.84
+ $X2=2.625 $Y2=1.84
r109 42 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=1.755
+ $X2=2.54 $Y2=1.84
r110 41 42 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.54 $Y=0.725
+ $X2=2.54 $Y2=1.755
r111 40 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=1.84
+ $X2=1.955 $Y2=1.84
r112 39 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=1.84
+ $X2=2.54 $Y2=1.84
r113 39 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.455 $Y=1.84
+ $X2=2.12 $Y2=1.84
r114 38 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=0.64
+ $X2=1.955 $Y2=0.64
r115 37 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.455 $Y=0.64
+ $X2=2.54 $Y2=0.725
r116 37 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.455 $Y=0.64
+ $X2=2.12 $Y2=0.64
r117 33 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.925
+ $X2=1.955 $Y2=1.84
r118 33 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.955 $Y=1.925
+ $X2=1.955 $Y2=2.335
r119 32 54 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.48 $Y=1.84
+ $X2=0.315 $Y2=1.84
r120 31 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=1.84
+ $X2=1.955 $Y2=1.84
r121 31 32 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.79 $Y=1.84
+ $X2=0.48 $Y2=1.84
r122 27 54 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.315 $Y=1.925
+ $X2=0.315 $Y2=1.84
r123 27 29 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.315 $Y=1.925
+ $X2=0.315 $Y2=2.335
r124 26 54 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.235 $Y=1.755
+ $X2=0.315 $Y2=1.84
r125 26 53 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.235 $Y=1.755
+ $X2=0.235 $Y2=0.725
r126 23 24 45.2433 $w=4.55e-07 $l=1.5e-07 $layer=POLY_cond $X=3.152 $Y=1.775
+ $X2=3.152 $Y2=1.925
r127 21 24 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.345 $Y=2.335
+ $X2=3.345 $Y2=1.925
r128 17 63 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.265 $Y=0.495
+ $X2=3.265 $Y2=1.255
r129 13 48 7.57836 $w=4.55e-07 $l=6.2e-08 $layer=POLY_cond $X=3.112 $Y=1.482
+ $X2=3.112 $Y2=1.42
r130 13 23 35.8139 $w=4.55e-07 $l=2.93e-07 $layer=POLY_cond $X=3.112 $Y=1.482
+ $X2=3.112 $Y2=1.775
r131 4 35 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.815
+ $Y=2.125 $X2=1.955 $Y2=2.335
r132 3 29 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.17
+ $Y=2.125 $X2=0.315 $Y2=2.335
r133 2 56 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.815
+ $Y=0.285 $X2=1.955 $Y2=0.495
r134 1 51 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.285 $X2=0.315 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_M%VPWR 1 2 9 13 15 17 22 32 33 36 39
r37 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r39 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r41 30 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.215 $Y=3.33
+ $X2=3.09 $Y2=3.33
r42 30 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=3.33
+ $X2=3.6 $Y2=3.33
r43 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r47 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.135 $Y2=3.33
r49 23 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=1.68
+ $Y2=3.33
r50 22 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.09 $Y2=3.33
r51 22 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.135 $Y2=3.33
r55 17 19 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 11 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=3.245
+ $X2=3.09 $Y2=3.33
r59 11 13 41.9489 $w=2.48e-07 $l=9.1e-07 $layer=LI1_cond $X=3.09 $Y=3.245
+ $X2=3.09 $Y2=2.335
r60 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=3.33
r61 7 9 31.7795 $w=3.28e-07 $l=9.1e-07 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=2.335
r62 2 13 600 $w=1.7e-07 $l=5.09289e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=2.125 $X2=3.05 $Y2=2.335
r63 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=2.125 $X2=1.135 $Y2=2.335
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_M%X 1 2 7 8 9 10 11 12 13 37
r15 12 13 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.56 $Y=2.335
+ $X2=3.56 $Y2=2.775
r16 11 12 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.56 $Y=2.035 $X2=3.56
+ $Y2=2.335
r17 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.56 $Y=1.665
+ $X2=3.56 $Y2=2.035
r18 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.56 $Y=1.295
+ $X2=3.56 $Y2=1.665
r19 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.56 $Y=0.925 $X2=3.56
+ $Y2=1.295
r20 8 41 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.56 $Y=0.925 $X2=3.56
+ $Y2=0.725
r21 7 41 5.25069 $w=4.08e-07 $l=1.7e-07 $layer=LI1_cond $X=3.52 $Y=0.555
+ $X2=3.52 $Y2=0.725
r22 7 37 1.6865 $w=4.08e-07 $l=6e-08 $layer=LI1_cond $X=3.52 $Y=0.555 $X2=3.52
+ $Y2=0.495
r23 2 12 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=2.125 $X2=3.56 $Y2=2.335
r24 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.34
+ $Y=0.285 $X2=3.48 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_M%VGND 1 2 9 13 16 17 18 20 33 34 37
r44 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r46 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r47 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r49 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.135
+ $Y2=0
r52 25 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.68
+ $Y2=0
r53 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r54 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.135
+ $Y2=0
r56 20 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.72
+ $Y2=0
r57 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r58 18 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r59 16 30 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.64
+ $Y2=0
r60 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.97
+ $Y2=0
r61 15 33 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.6
+ $Y2=0
r62 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=2.97
+ $Y2=0
r63 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=2.97 $Y2=0
r64 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=2.97 $Y2=0.495
r65 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0
r66 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0.495
r67 2 13 182 $w=1.7e-07 $l=4.27288e-07 $layer=licon1_NDIFF $count=1 $X=2.635
+ $Y=0.285 $X2=2.97 $Y2=0.495
r68 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.285 $X2=1.135 $Y2=0.495
.ends

