* NGSPICE file created from sky130_fd_sc_lp__o41a_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o41a_lp A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VGND A3 a_31_57# VNB nshort w=420000u l=150000u
+  ad=4.41e+11p pd=4.62e+06u as=3.696e+11p ps=4.28e+06u
M1001 X a_457_412# a_708_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1002 VGND A1 a_31_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_31_57# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_457_412# A4 a_349_412# VPB phighvt w=1e+06u l=250000u
+  ad=5.65e+11p pd=3.13e+06u as=2.9e+11p ps=2.58e+06u
M1005 X a_457_412# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=6.8e+11p ps=5.36e+06u
M1006 a_708_47# a_457_412# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_349_412# A3 a_235_412# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1008 a_137_412# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1009 a_31_57# A4 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_235_412# A2 a_137_412# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_457_412# B1 a_31_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1012 VPWR B1 a_457_412# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

