* File: sky130_fd_sc_lp__nor2b_m.pex.spice
* Created: Wed Sep  2 10:08:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2B_M%B_N 3 9 11 12 13 14 15 16 17 24
r42 24 26 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.687 $Y=1.435
+ $X2=0.687 $Y2=1.27
r43 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=1.435 $X2=0.71 $Y2=1.435
r44 16 17 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=1.665
+ $X2=0.715 $Y2=2.035
r45 16 25 14.1717 $w=1.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.715 $Y=1.665
+ $X2=0.715 $Y2=1.435
r46 15 25 8.62626 $w=1.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.715 $Y=1.295
+ $X2=0.715 $Y2=1.435
r47 14 15 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.925
+ $X2=0.715 $Y2=1.295
r48 13 14 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.555
+ $X2=0.715 $Y2=0.925
r49 11 12 42.9311 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=0.777 $Y=1.79
+ $X2=0.777 $Y2=1.94
r50 9 12 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.98 $Y=2.67 $X2=0.98
+ $Y2=1.94
r51 5 24 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.687 $Y=1.457
+ $X2=0.687 $Y2=1.435
r52 5 11 49.3865 $w=3.75e-07 $l=3.33e-07 $layer=POLY_cond $X=0.687 $Y=1.457
+ $X2=0.687 $Y2=1.79
r53 3 26 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.575 $Y=0.56
+ $X2=0.575 $Y2=1.27
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_M%A 3 5 6 8 10 11 12 15 17 18 19 20 26
c60 17 0 1.51825e-19 $X=1.2 $Y=0.925
r61 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.25
+ $Y=1.045 $X2=1.25 $Y2=1.045
r62 19 20 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.225 $Y=1.665
+ $X2=1.225 $Y2=2.035
r63 18 19 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.225 $Y=1.295
+ $X2=1.225 $Y2=1.665
r64 18 27 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=1.225 $Y=1.295
+ $X2=1.225 $Y2=1.045
r65 17 27 6.28605 $w=2.18e-07 $l=1.2e-07 $layer=LI1_cond $X=1.225 $Y=0.925
+ $X2=1.225 $Y2=1.045
r66 13 15 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.34 $Y=2.275
+ $X2=1.565 $Y2=2.275
r67 11 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.25 $Y=1.385
+ $X2=1.25 $Y2=1.045
r68 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.385
+ $X2=1.25 $Y2=1.55
r69 10 26 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=0.88
+ $X2=1.25 $Y2=1.045
r70 6 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.565 $Y=2.35
+ $X2=1.565 $Y2=2.275
r71 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.565 $Y=2.35
+ $X2=1.565 $Y2=2.67
r72 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.34 $Y=2.2 $X2=1.34
+ $Y2=2.275
r73 5 12 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.34 $Y=2.2 $X2=1.34
+ $Y2=1.55
r74 3 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.285 $Y=0.56
+ $X2=1.285 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_M%A_47_70# 1 2 8 11 15 17 20 22 23 26 27
c61 15 0 1.51825e-19 $X=1.925 $Y=2.67
r62 27 33 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.812 $Y=1.455
+ $X2=1.812 $Y2=1.29
r63 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.79
+ $Y=1.455 $X2=1.79 $Y2=1.455
r64 24 26 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.79 $Y=2.3
+ $X2=1.79 $Y2=1.455
r65 23 31 9.01297 $w=2.9e-07 $l=2.16852e-07 $layer=LI1_cond $X=0.91 $Y=2.385
+ $X2=0.745 $Y2=2.505
r66 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.705 $Y=2.385
+ $X2=1.79 $Y2=2.3
r67 22 23 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.705 $Y=2.385
+ $X2=0.91 $Y2=2.385
r68 18 31 16.6172 $w=2.9e-07 $l=4.86826e-07 $layer=LI1_cond $X=0.35 $Y=2.3
+ $X2=0.745 $Y2=2.505
r69 18 20 97.7751 $w=1.88e-07 $l=1.675e-06 $layer=LI1_cond $X=0.35 $Y=2.3
+ $X2=0.35 $Y2=0.625
r70 15 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.925 $Y=2.67
+ $X2=1.925 $Y2=1.96
r71 11 33 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.715 $Y=0.56
+ $X2=1.715 $Y2=1.29
r72 8 17 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=1.812 $Y=1.773
+ $X2=1.812 $Y2=1.96
r73 7 27 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=1.812 $Y=1.477
+ $X2=1.812 $Y2=1.455
r74 7 8 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=1.812 $Y=1.477
+ $X2=1.812 $Y2=1.773
r75 2 31 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=2.46 $X2=0.745 $Y2=2.605
r76 1 20 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.35 $X2=0.36 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_M%VPWR 1 6 8 10 17 18 21
r22 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r23 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=3.33
+ $X2=1.255 $Y2=3.33
r24 15 17 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.42 $Y=3.33
+ $X2=2.16 $Y2=3.33
r25 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=1.255 $Y2=3.33
r27 10 12 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=3.33 $X2=0.72
+ $Y2=3.33
r28 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r29 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.72
+ $Y2=3.33
r30 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r31 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=3.245
+ $X2=1.255 $Y2=3.33
r32 4 6 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.255 $Y=3.245
+ $X2=1.255 $Y2=2.755
r33 1 6 600 $w=1.7e-07 $l=3.82132e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=2.46 $X2=1.255 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_M%Y 1 2 8 9 10 14 16 17 18 19 20 21
r30 21 40 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.15 $Y=2.775
+ $X2=2.15 $Y2=2.605
r31 20 40 11.6746 $w=1.88e-07 $l=2e-07 $layer=LI1_cond $X=2.15 $Y=2.405 $X2=2.15
+ $Y2=2.605
r32 19 20 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.15 $Y=2.035
+ $X2=2.15 $Y2=2.405
r33 18 19 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.15 $Y=1.665
+ $X2=2.15 $Y2=2.035
r34 17 18 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.665
r35 16 17 11.68 $w=3.58e-07 $l=2.85e-07 $layer=LI1_cond $X=2.15 $Y=1.01 $X2=2.15
+ $Y2=1.295
r36 12 14 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=1.5 $Y=0.555 $X2=1.6
+ $Y2=0.555
r37 9 16 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.055 $Y=0.925
+ $X2=2.15 $Y2=0.925
r38 9 10 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.055 $Y=0.925
+ $X2=1.685 $Y2=0.925
r39 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=0.84
+ $X2=1.685 $Y2=0.925
r40 7 14 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.6 $Y=0.66 $X2=1.6
+ $Y2=0.555
r41 7 8 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.6 $Y=0.66 $X2=1.6
+ $Y2=0.84
r42 2 40 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2 $Y=2.46
+ $X2=2.14 $Y2=2.605
r43 1 12 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.36
+ $Y=0.35 $X2=1.5 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_M%VGND 1 2 9 13 16 17 19 20 21 31 32
r32 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r33 29 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r34 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r35 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r37 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r38 19 28 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.68
+ $Y2=0
r39 19 20 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.96
+ $Y2=0
r40 18 31 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.16
+ $Y2=0
r41 18 20 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.055 $Y=0 $X2=1.96
+ $Y2=0
r42 16 24 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r43 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.07
+ $Y2=0
r44 15 28 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.68
+ $Y2=0
r45 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.07
+ $Y2=0
r46 11 20 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r47 11 13 23.933 $w=1.88e-07 $l=4.1e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.495
r48 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r49 7 9 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0.495
r50 2 13 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.79
+ $Y=0.35 $X2=1.95 $Y2=0.495
r51 1 9 182 $w=1.7e-07 $l=4.87134e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.35 $X2=1.07 $Y2=0.495
.ends

