* File: sky130_fd_sc_lp__mux2i_4.pxi.spice
* Created: Fri Aug 28 10:45:18 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2I_4%A0 N_A0_M1005_g N_A0_M1001_g N_A0_M1020_g
+ N_A0_M1014_g N_A0_M1024_g N_A0_M1016_g N_A0_M1029_g N_A0_M1025_g A0 A0 A0
+ N_A0_c_129_n N_A0_c_130_n PM_SKY130_FD_SC_LP__MUX2I_4%A0
x_PM_SKY130_FD_SC_LP__MUX2I_4%A1 N_A1_M1002_g N_A1_M1007_g N_A1_M1013_g
+ N_A1_M1018_g N_A1_M1023_g N_A1_M1019_g N_A1_M1032_g N_A1_M1030_g A1 A1 A1
+ N_A1_c_206_n N_A1_c_207_n PM_SKY130_FD_SC_LP__MUX2I_4%A1
x_PM_SKY130_FD_SC_LP__MUX2I_4%S N_S_M1000_g N_S_M1010_g N_S_M1004_g N_S_M1012_g
+ N_S_M1017_g N_S_M1031_g N_S_M1033_g N_S_M1026_g N_S_c_276_n N_S_M1003_g
+ N_S_c_277_n N_S_M1015_g N_S_c_288_n N_S_c_278_n S S S S S S N_S_c_280_n
+ N_S_c_281_n PM_SKY130_FD_SC_LP__MUX2I_4%S
x_PM_SKY130_FD_SC_LP__MUX2I_4%A_1418_21# N_A_1418_21#_M1003_d
+ N_A_1418_21#_M1015_d N_A_1418_21#_M1006_g N_A_1418_21#_c_414_n
+ N_A_1418_21#_M1008_g N_A_1418_21#_M1009_g N_A_1418_21#_c_415_n
+ N_A_1418_21#_M1011_g N_A_1418_21#_M1027_g N_A_1418_21#_c_416_n
+ N_A_1418_21#_M1021_g N_A_1418_21#_M1028_g N_A_1418_21#_c_417_n
+ N_A_1418_21#_M1022_g N_A_1418_21#_c_408_n N_A_1418_21#_c_409_n
+ N_A_1418_21#_c_410_n N_A_1418_21#_c_486_p N_A_1418_21#_c_506_p
+ N_A_1418_21#_c_418_n N_A_1418_21#_c_419_n N_A_1418_21#_c_411_n
+ N_A_1418_21#_c_412_n N_A_1418_21#_c_413_n
+ PM_SKY130_FD_SC_LP__MUX2I_4%A_1418_21#
x_PM_SKY130_FD_SC_LP__MUX2I_4%Y N_Y_M1005_s N_Y_M1020_s N_Y_M1029_s N_Y_M1018_d
+ N_Y_M1030_d N_Y_M1001_d N_Y_M1014_d N_Y_M1025_d N_Y_M1013_d N_Y_M1032_d
+ N_Y_c_513_n N_Y_c_524_n N_Y_c_590_p N_Y_c_514_n N_Y_c_515_n N_Y_c_531_n
+ N_Y_c_521_n N_Y_c_516_n N_Y_c_560_n N_Y_c_517_n N_Y_c_518_n N_Y_c_519_n
+ N_Y_c_548_n Y N_Y_c_520_n PM_SKY130_FD_SC_LP__MUX2I_4%Y
x_PM_SKY130_FD_SC_LP__MUX2I_4%A_126_367# N_A_126_367#_M1001_s
+ N_A_126_367#_M1016_s N_A_126_367#_M1000_s N_A_126_367#_M1017_s
+ N_A_126_367#_c_640_n N_A_126_367#_c_625_n N_A_126_367#_c_662_p
+ N_A_126_367#_c_644_n N_A_126_367#_c_622_n N_A_126_367#_c_623_n
+ N_A_126_367#_c_624_n PM_SKY130_FD_SC_LP__MUX2I_4%A_126_367#
x_PM_SKY130_FD_SC_LP__MUX2I_4%A_470_367# N_A_470_367#_M1007_s
+ N_A_470_367#_M1023_s N_A_470_367#_M1008_s N_A_470_367#_M1021_s
+ N_A_470_367#_c_671_n N_A_470_367#_c_669_n N_A_470_367#_c_686_n
+ N_A_470_367#_c_676_n N_A_470_367#_c_677_n N_A_470_367#_c_691_n
+ N_A_470_367#_c_705_n N_A_470_367#_c_670_n N_A_470_367#_c_679_n
+ N_A_470_367#_c_684_n PM_SKY130_FD_SC_LP__MUX2I_4%A_470_367#
x_PM_SKY130_FD_SC_LP__MUX2I_4%VPWR N_VPWR_M1000_d N_VPWR_M1004_d N_VPWR_M1026_d
+ N_VPWR_M1011_d N_VPWR_M1022_d N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_742_n
+ N_VPWR_c_743_n VPWR N_VPWR_c_744_n N_VPWR_c_745_n N_VPWR_c_746_n
+ N_VPWR_c_747_n N_VPWR_c_748_n N_VPWR_c_749_n N_VPWR_c_739_n N_VPWR_c_751_n
+ N_VPWR_c_752_n N_VPWR_c_753_n N_VPWR_c_754_n N_VPWR_c_755_n
+ PM_SKY130_FD_SC_LP__MUX2I_4%VPWR
x_PM_SKY130_FD_SC_LP__MUX2I_4%A_110_69# N_A_110_69#_M1005_d N_A_110_69#_M1024_d
+ N_A_110_69#_M1006_s N_A_110_69#_M1027_s N_A_110_69#_c_867_n
+ N_A_110_69#_c_859_n N_A_110_69#_c_860_n N_A_110_69#_c_875_n
+ N_A_110_69#_c_861_n N_A_110_69#_c_862_n N_A_110_69#_c_863_n
+ N_A_110_69#_c_864_n N_A_110_69#_c_940_p N_A_110_69#_c_865_n
+ N_A_110_69#_c_941_p N_A_110_69#_c_866_n PM_SKY130_FD_SC_LP__MUX2I_4%A_110_69#
x_PM_SKY130_FD_SC_LP__MUX2I_4%A_470_69# N_A_470_69#_M1002_s N_A_470_69#_M1019_s
+ N_A_470_69#_M1010_s N_A_470_69#_M1031_s N_A_470_69#_c_949_n
+ N_A_470_69#_c_950_n N_A_470_69#_c_951_n N_A_470_69#_c_952_n
+ N_A_470_69#_c_959_n N_A_470_69#_c_962_n N_A_470_69#_c_965_n
+ N_A_470_69#_c_968_n PM_SKY130_FD_SC_LP__MUX2I_4%A_470_69#
x_PM_SKY130_FD_SC_LP__MUX2I_4%VGND N_VGND_M1010_d N_VGND_M1012_d N_VGND_M1033_d
+ N_VGND_M1009_d N_VGND_M1028_d N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n
+ N_VGND_c_1011_n N_VGND_c_1012_n N_VGND_c_1013_n N_VGND_c_1014_n
+ N_VGND_c_1015_n N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n
+ N_VGND_c_1019_n VGND N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n
+ N_VGND_c_1023_n N_VGND_c_1024_n PM_SKY130_FD_SC_LP__MUX2I_4%VGND
cc_1 VNB N_A0_M1005_g 0.025538f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_2 VNB N_A0_M1020_g 0.0191117f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.765
cc_3 VNB N_A0_M1024_g 0.0190879f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=0.765
cc_4 VNB N_A0_M1029_g 0.0184007f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=0.765
cc_5 VNB N_A0_c_129_n 0.0115663f $X=-0.19 $Y=-0.245 $X2=1.55 $Y2=1.51
cc_6 VNB N_A0_c_130_n 0.0775437f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.51
cc_7 VNB N_A1_M1002_g 0.0206964f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_8 VNB N_A1_M1018_g 0.0203457f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_9 VNB N_A1_M1019_g 0.0203628f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=2.465
cc_10 VNB N_A1_M1030_g 0.0234178f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.465
cc_11 VNB N_A1_c_206_n 0.00991891f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.51
cc_12 VNB N_A1_c_207_n 0.0889352f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.51
cc_13 VNB N_S_M1010_g 0.0310912f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_14 VNB N_S_M1012_g 0.0229027f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_15 VNB N_S_M1031_g 0.0229027f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=2.465
cc_16 VNB N_S_M1033_g 0.023138f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=0.765
cc_17 VNB N_S_c_276_n 0.0193851f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_S_c_277_n 0.0474653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_S_c_278_n 0.00226194f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.51
cc_20 VNB S 0.0177041f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.51
cc_21 VNB N_S_c_280_n 0.0706327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_S_c_281_n 0.00355698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_1418_21#_M1006_g 0.0228952f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.345
cc_24 VNB N_A_1418_21#_M1009_g 0.0227036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_1418_21#_M1027_g 0.0226963f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=2.465
cc_26 VNB N_A_1418_21#_M1028_g 0.0229962f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.465
cc_27 VNB N_A_1418_21#_c_408_n 0.00103041f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_28 VNB N_A_1418_21#_c_409_n 0.0019826f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.51
cc_29 VNB N_A_1418_21#_c_410_n 0.00237512f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.51
cc_30 VNB N_A_1418_21#_c_411_n 0.0247561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_1418_21#_c_412_n 0.0235668f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.587
cc_32 VNB N_A_1418_21#_c_413_n 0.0733075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_513_n 0.00249281f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_34 VNB N_Y_c_514_n 0.00330243f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_35 VNB N_Y_c_515_n 0.00440725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_516_n 0.00379012f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.51
cc_37 VNB N_Y_c_517_n 0.00224921f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.587
cc_38 VNB N_Y_c_518_n 0.0152383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_519_n 0.00238675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_520_n 0.00333866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VPWR_c_739_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_110_69#_c_859_n 0.00458861f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.345
cc_43 VNB N_A_110_69#_c_860_n 0.00203674f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=0.765
cc_44 VNB N_A_110_69#_c_861_n 0.0131582f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.675
cc_45 VNB N_A_110_69#_c_862_n 0.0114714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_110_69#_c_863_n 0.042375f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.345
cc_47 VNB N_A_110_69#_c_864_n 0.00391207f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=0.765
cc_48 VNB N_A_110_69#_c_865_n 0.0118262f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.465
cc_49 VNB N_A_110_69#_c_866_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_50 VNB N_A_470_69#_c_949_n 0.0251624f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.675
cc_51 VNB N_A_470_69#_c_950_n 0.0108348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_470_69#_c_951_n 0.0041456f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.675
cc_53 VNB N_A_470_69#_c_952_n 0.0042908f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=2.465
cc_54 VNB N_VGND_c_1008_n 0.00430043f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=0.765
cc_55 VNB N_VGND_c_1009_n 0.0174138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1010_n 0.00372238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1011_n 0.00178362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1012_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1013_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1014_n 0.123701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1015_n 0.00362784f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_62 VNB N_VGND_c_1016_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.51
cc_63 VNB N_VGND_c_1017_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.51
cc_64 VNB N_VGND_c_1018_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.51
cc_65 VNB N_VGND_c_1019_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.51
cc_66 VNB N_VGND_c_1020_n 0.0173211f $X=-0.19 $Y=-0.245 $X2=1.55 $Y2=1.51
cc_67 VNB N_VGND_c_1021_n 0.0235776f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.587
cc_68 VNB N_VGND_c_1022_n 0.488862f $X=-0.19 $Y=-0.245 $X2=1.55 $Y2=1.587
cc_69 VNB N_VGND_c_1023_n 0.00362451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1024_n 0.00378455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VPB N_A0_M1001_g 0.0244533f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_72 VPB N_A0_M1014_g 0.0181378f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_73 VPB N_A0_M1016_g 0.0181378f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=2.465
cc_74 VPB N_A0_M1025_g 0.0190451f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=2.465
cc_75 VPB N_A0_c_129_n 0.0174544f $X=-0.19 $Y=1.655 $X2=1.55 $Y2=1.51
cc_76 VPB N_A0_c_130_n 0.0161279f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=1.51
cc_77 VPB N_A1_M1007_g 0.0190426f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_78 VPB N_A1_M1013_g 0.0180542f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.765
cc_79 VPB N_A1_M1023_g 0.0180542f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=0.765
cc_80 VPB N_A1_M1032_g 0.0227262f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=0.765
cc_81 VPB N_A1_c_206_n 0.0103211f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=1.51
cc_82 VPB N_A1_c_207_n 0.022189f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=1.51
cc_83 VPB N_S_M1000_g 0.0224653f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_84 VPB N_S_M1004_g 0.017193f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.765
cc_85 VPB N_S_M1017_g 0.0174281f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=0.765
cc_86 VPB N_S_M1026_g 0.0174489f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=2.465
cc_87 VPB N_S_c_277_n 0.00631588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_S_M1015_g 0.0221029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_S_c_288_n 0.00950074f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_S_c_278_n 0.00189476f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.51
cc_91 VPB S 0.0246203f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=1.51
cc_92 VPB N_S_c_280_n 0.0130822f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_S_c_281_n 0.00129169f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_1418_21#_c_414_n 0.0155329f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.765
cc_95 VPB N_A_1418_21#_c_415_n 0.017003f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=0.765
cc_96 VPB N_A_1418_21#_c_416_n 0.0170041f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=1.345
cc_97 VPB N_A_1418_21#_c_417_n 0.0159622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_1418_21#_c_418_n 0.00636377f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=1.51
cc_99 VPB N_A_1418_21#_c_419_n 0.0441363f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.51
cc_100 VPB N_A_1418_21#_c_412_n 0.00890909f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.587
cc_101 VPB N_A_1418_21#_c_413_n 0.0258564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_Y_c_521_n 0.0149845f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.51
cc_103 VPB N_Y_c_518_n 0.00957929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_126_367#_c_622_n 0.0109459f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=0.765
cc_105 VPB N_A_126_367#_c_623_n 0.0177068f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=2.465
cc_106 VPB N_A_126_367#_c_624_n 0.0189931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_470_367#_c_669_n 0.0243943f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.345
cc_108 VPB N_A_470_367#_c_670_n 0.00988841f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_109 VPB N_VPWR_c_740_n 3.31199e-19 $X=-0.19 $Y=1.655 $X2=1.415 $Y2=0.765
cc_110 VPB N_VPWR_c_741_n 3.25996e-19 $X=-0.19 $Y=1.655 $X2=1.415 $Y2=2.465
cc_111 VPB N_VPWR_c_742_n 0.00493241f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=0.765
cc_112 VPB N_VPWR_c_743_n 0.00251047f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=2.465
cc_113 VPB N_VPWR_c_744_n 0.131688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_745_n 0.0166969f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.51
cc_115 VPB N_VPWR_c_746_n 0.0130051f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.51
cc_116 VPB N_VPWR_c_747_n 0.0150899f $X=-0.19 $Y=1.655 $X2=1.55 $Y2=1.51
cc_117 VPB N_VPWR_c_748_n 0.018457f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.587
cc_118 VPB N_VPWR_c_749_n 0.0164495f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.587
cc_119 VPB N_VPWR_c_739_n 0.0612538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_751_n 0.0150851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_752_n 0.00436274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_753_n 0.00436274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_754_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_755_n 0.00414668f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 N_A0_M1029_g N_A1_M1002_g 0.0355293f $X=1.845 $Y=0.765 $X2=0 $Y2=0
cc_126 N_A0_M1025_g N_A1_M1007_g 0.0355293f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A0_c_130_n N_A1_c_206_n 0.00105815f $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_128 N_A0_c_129_n N_A1_c_207_n 0.00104983f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A0_c_130_n N_A1_c_207_n 0.0355293f $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A0_M1005_g N_Y_c_513_n 0.00350469f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_131 N_A0_c_129_n N_Y_c_524_n 0.0156951f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A0_c_130_n N_Y_c_524_n 3.83932e-19 $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_133 N_A0_M1005_g N_Y_c_514_n 0.013408f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_134 N_A0_M1020_g N_Y_c_514_n 0.0113303f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_135 N_A0_c_129_n N_Y_c_514_n 0.0485315f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_136 N_A0_c_130_n N_Y_c_514_n 0.00364629f $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_137 N_A0_c_129_n N_Y_c_515_n 0.0161224f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_138 N_A0_M1001_g N_Y_c_531_n 0.0130544f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A0_M1014_g N_Y_c_531_n 0.0130078f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A0_c_129_n N_Y_c_531_n 0.0417123f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_141 N_A0_c_130_n N_Y_c_531_n 5.68911e-19 $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_142 N_A0_M1016_g N_Y_c_521_n 0.0110437f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A0_M1025_g N_Y_c_521_n 0.012798f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A0_c_129_n N_Y_c_521_n 0.0272288f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_145 N_A0_c_130_n N_Y_c_521_n 5.77374e-19 $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_146 N_A0_M1024_g N_Y_c_516_n 0.0127418f $X=1.415 $Y=0.765 $X2=0 $Y2=0
cc_147 N_A0_M1029_g N_Y_c_516_n 0.0150214f $X=1.845 $Y=0.765 $X2=0 $Y2=0
cc_148 N_A0_c_129_n N_Y_c_516_n 0.0256582f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A0_c_130_n N_Y_c_516_n 0.00248147f $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A0_M1020_g N_Y_c_519_n 4.11272e-19 $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_151 N_A0_M1024_g N_Y_c_519_n 0.00756439f $X=1.415 $Y=0.765 $X2=0 $Y2=0
cc_152 N_A0_M1029_g N_Y_c_519_n 8.93811e-19 $X=1.845 $Y=0.765 $X2=0 $Y2=0
cc_153 N_A0_c_129_n N_Y_c_519_n 0.0261235f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_154 N_A0_c_130_n N_Y_c_519_n 0.00491511f $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A0_c_129_n N_Y_c_548_n 0.0139322f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_156 N_A0_c_130_n N_Y_c_548_n 6.47588e-19 $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A0_M1024_g N_Y_c_520_n 6.11822e-19 $X=1.415 $Y=0.765 $X2=0 $Y2=0
cc_158 N_A0_M1029_g N_Y_c_520_n 0.00545809f $X=1.845 $Y=0.765 $X2=0 $Y2=0
cc_159 N_A0_c_129_n N_Y_c_520_n 0.00337525f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A0_c_130_n N_Y_c_520_n 0.00686853f $X=1.845 $Y=1.51 $X2=0 $Y2=0
cc_161 N_A0_M1014_g N_A_126_367#_c_625_n 0.0129895f $X=0.985 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A0_M1016_g N_A_126_367#_c_625_n 0.0107022f $X=1.415 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A0_M1025_g N_A_126_367#_c_623_n 0.0132528f $X=1.845 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A0_M1001_g N_VPWR_c_744_n 0.00585385f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A0_M1014_g N_VPWR_c_744_n 0.00382632f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A0_M1016_g N_VPWR_c_744_n 0.00382632f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A0_M1025_g N_VPWR_c_744_n 0.00585385f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A0_M1001_g N_VPWR_c_739_n 0.0120577f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A0_M1014_g N_VPWR_c_739_n 0.0055144f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A0_M1016_g N_VPWR_c_739_n 0.0055144f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A0_M1025_g N_VPWR_c_739_n 0.0110081f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A0_M1005_g N_A_110_69#_c_867_n 0.00523186f $X=0.475 $Y=0.765 $X2=0
+ $Y2=0
cc_173 N_A0_M1020_g N_A_110_69#_c_867_n 0.00664098f $X=0.905 $Y=0.765 $X2=0
+ $Y2=0
cc_174 N_A0_M1024_g N_A_110_69#_c_867_n 5.84315e-19 $X=1.415 $Y=0.765 $X2=0
+ $Y2=0
cc_175 N_A0_M1020_g N_A_110_69#_c_859_n 0.00938101f $X=0.905 $Y=0.765 $X2=0
+ $Y2=0
cc_176 N_A0_M1024_g N_A_110_69#_c_859_n 0.0121498f $X=1.415 $Y=0.765 $X2=0 $Y2=0
cc_177 N_A0_M1029_g N_A_110_69#_c_859_n 0.00602332f $X=1.845 $Y=0.765 $X2=0
+ $Y2=0
cc_178 N_A0_M1005_g N_A_110_69#_c_860_n 0.00592745f $X=0.475 $Y=0.765 $X2=0
+ $Y2=0
cc_179 N_A0_M1020_g N_A_110_69#_c_860_n 0.00166018f $X=0.905 $Y=0.765 $X2=0
+ $Y2=0
cc_180 N_A0_M1029_g N_A_110_69#_c_875_n 0.00372352f $X=1.845 $Y=0.765 $X2=0
+ $Y2=0
cc_181 N_A0_M1029_g N_A_110_69#_c_861_n 0.00826878f $X=1.845 $Y=0.765 $X2=0
+ $Y2=0
cc_182 N_A0_M1005_g N_VGND_c_1014_n 0.00450424f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_183 N_A0_M1020_g N_VGND_c_1014_n 0.00291444f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_184 N_A0_M1024_g N_VGND_c_1014_n 0.0029147f $X=1.415 $Y=0.765 $X2=0 $Y2=0
cc_185 N_A0_M1029_g N_VGND_c_1014_n 0.00332982f $X=1.845 $Y=0.765 $X2=0 $Y2=0
cc_186 N_A0_M1005_g N_VGND_c_1022_n 0.00883394f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_187 N_A0_M1020_g N_VGND_c_1022_n 0.00403101f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_188 N_A0_M1024_g N_VGND_c_1022_n 0.00403103f $X=1.415 $Y=0.765 $X2=0 $Y2=0
cc_189 N_A0_M1029_g N_VGND_c_1022_n 0.00447438f $X=1.845 $Y=0.765 $X2=0 $Y2=0
cc_190 N_A1_M1007_g N_Y_c_521_n 0.0121462f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A1_M1013_g N_Y_c_521_n 0.00871272f $X=2.705 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A1_M1023_g N_Y_c_521_n 0.00871272f $X=3.135 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A1_M1032_g N_Y_c_521_n 0.00871272f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A1_c_206_n N_Y_c_521_n 0.0922055f $X=3.61 $Y=1.51 $X2=0 $Y2=0
cc_195 N_A1_c_207_n N_Y_c_521_n 0.00938937f $X=3.885 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A1_M1002_g N_Y_c_560_n 0.0112623f $X=2.275 $Y=0.765 $X2=0 $Y2=0
cc_197 N_A1_M1018_g N_Y_c_560_n 0.0101957f $X=2.865 $Y=0.765 $X2=0 $Y2=0
cc_198 N_A1_M1019_g N_Y_c_560_n 0.0101957f $X=3.295 $Y=0.765 $X2=0 $Y2=0
cc_199 N_A1_M1030_g N_Y_c_560_n 0.0144905f $X=3.885 $Y=0.765 $X2=0 $Y2=0
cc_200 N_A1_c_206_n N_Y_c_560_n 0.0972461f $X=3.61 $Y=1.51 $X2=0 $Y2=0
cc_201 N_A1_c_207_n N_Y_c_560_n 0.0042625f $X=3.885 $Y=1.51 $X2=0 $Y2=0
cc_202 N_A1_M1032_g N_Y_c_518_n 0.00353704f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A1_M1030_g N_Y_c_518_n 0.0155398f $X=3.885 $Y=0.765 $X2=0 $Y2=0
cc_204 N_A1_c_206_n N_Y_c_518_n 0.0214314f $X=3.61 $Y=1.51 $X2=0 $Y2=0
cc_205 N_A1_M1002_g N_Y_c_520_n 0.00827979f $X=2.275 $Y=0.765 $X2=0 $Y2=0
cc_206 N_A1_M1018_g N_Y_c_520_n 9.18514e-19 $X=2.865 $Y=0.765 $X2=0 $Y2=0
cc_207 N_A1_c_206_n N_Y_c_520_n 0.0107665f $X=3.61 $Y=1.51 $X2=0 $Y2=0
cc_208 N_A1_c_207_n N_Y_c_520_n 0.00511949f $X=3.885 $Y=1.51 $X2=0 $Y2=0
cc_209 N_A1_M1007_g N_A_126_367#_c_623_n 0.0154538f $X=2.275 $Y=2.465 $X2=0
+ $Y2=0
cc_210 N_A1_M1013_g N_A_126_367#_c_623_n 0.010883f $X=2.705 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A1_M1023_g N_A_126_367#_c_623_n 0.010883f $X=3.135 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A1_M1032_g N_A_126_367#_c_623_n 0.013045f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A1_M1013_g N_A_470_367#_c_671_n 0.0156515f $X=2.705 $Y=2.465 $X2=0
+ $Y2=0
cc_214 N_A1_M1023_g N_A_470_367#_c_671_n 0.0156046f $X=3.135 $Y=2.465 $X2=0
+ $Y2=0
cc_215 N_A1_M1032_g N_A_470_367#_c_669_n 0.0113549f $X=3.565 $Y=2.465 $X2=0
+ $Y2=0
cc_216 N_A1_M1007_g N_VPWR_c_744_n 0.00585385f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A1_M1013_g N_VPWR_c_744_n 0.00357877f $X=2.705 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A1_M1023_g N_VPWR_c_744_n 0.00357877f $X=3.135 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A1_M1032_g N_VPWR_c_744_n 0.00408809f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A1_M1007_g N_VPWR_c_739_n 0.0110081f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A1_M1013_g N_VPWR_c_739_n 0.00542194f $X=2.705 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A1_M1023_g N_VPWR_c_739_n 0.00542194f $X=3.135 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A1_M1032_g N_VPWR_c_739_n 0.00718256f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A1_M1002_g N_A_110_69#_c_859_n 6.08975e-19 $X=2.275 $Y=0.765 $X2=0
+ $Y2=0
cc_225 N_A1_M1002_g N_A_110_69#_c_875_n 8.26284e-19 $X=2.275 $Y=0.765 $X2=0
+ $Y2=0
cc_226 N_A1_M1002_g N_A_110_69#_c_861_n 0.0124015f $X=2.275 $Y=0.765 $X2=0 $Y2=0
cc_227 N_A1_M1018_g N_A_110_69#_c_861_n 0.0112681f $X=2.865 $Y=0.765 $X2=0 $Y2=0
cc_228 N_A1_M1019_g N_A_110_69#_c_861_n 0.0112681f $X=3.295 $Y=0.765 $X2=0 $Y2=0
cc_229 N_A1_M1030_g N_A_110_69#_c_861_n 0.0132234f $X=3.885 $Y=0.765 $X2=0 $Y2=0
cc_230 N_A1_M1030_g N_A_110_69#_c_862_n 0.00295605f $X=3.885 $Y=0.765 $X2=0
+ $Y2=0
cc_231 N_A1_M1002_g N_A_470_69#_c_949_n 0.0022355f $X=2.275 $Y=0.765 $X2=0 $Y2=0
cc_232 N_A1_M1018_g N_A_470_69#_c_949_n 0.0110236f $X=2.865 $Y=0.765 $X2=0 $Y2=0
cc_233 N_A1_M1019_g N_A_470_69#_c_949_n 0.0114012f $X=3.295 $Y=0.765 $X2=0 $Y2=0
cc_234 N_A1_M1030_g N_A_470_69#_c_949_n 0.0138062f $X=3.885 $Y=0.765 $X2=0 $Y2=0
cc_235 N_A1_M1002_g N_VGND_c_1014_n 0.00341315f $X=2.275 $Y=0.765 $X2=0 $Y2=0
cc_236 N_A1_M1018_g N_VGND_c_1014_n 0.0029147f $X=2.865 $Y=0.765 $X2=0 $Y2=0
cc_237 N_A1_M1019_g N_VGND_c_1014_n 0.0029147f $X=3.295 $Y=0.765 $X2=0 $Y2=0
cc_238 N_A1_M1030_g N_VGND_c_1014_n 0.0029147f $X=3.885 $Y=0.765 $X2=0 $Y2=0
cc_239 N_A1_M1002_g N_VGND_c_1022_n 0.0046539f $X=2.275 $Y=0.765 $X2=0 $Y2=0
cc_240 N_A1_M1018_g N_VGND_c_1022_n 0.00406937f $X=2.865 $Y=0.765 $X2=0 $Y2=0
cc_241 N_A1_M1019_g N_VGND_c_1022_n 0.00406937f $X=3.295 $Y=0.765 $X2=0 $Y2=0
cc_242 N_A1_M1030_g N_VGND_c_1022_n 0.0043693f $X=3.885 $Y=0.765 $X2=0 $Y2=0
cc_243 N_S_M1033_g N_A_1418_21#_M1006_g 0.0167479f $X=6.735 $Y=0.655 $X2=0 $Y2=0
cc_244 N_S_M1026_g N_A_1418_21#_c_414_n 0.029401f $X=6.745 $Y=2.465 $X2=0 $Y2=0
cc_245 N_S_c_288_n N_A_1418_21#_c_414_n 0.0116353f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_246 N_S_c_288_n N_A_1418_21#_c_415_n 0.0112519f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_247 N_S_c_288_n N_A_1418_21#_c_416_n 0.0112926f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_248 N_S_c_276_n N_A_1418_21#_M1028_g 0.0241795f $X=8.885 $Y=1.185 $X2=0 $Y2=0
cc_249 N_S_c_277_n N_A_1418_21#_M1028_g 2.84688e-19 $X=9.075 $Y=1.665 $X2=0
+ $Y2=0
cc_250 N_S_c_288_n N_A_1418_21#_c_417_n 0.0145464f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_251 N_S_c_277_n N_A_1418_21#_c_408_n 6.23007e-19 $X=9.075 $Y=1.665 $X2=0
+ $Y2=0
cc_252 N_S_c_288_n N_A_1418_21#_c_408_n 0.104029f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_253 N_S_c_278_n N_A_1418_21#_c_408_n 0.0160161f $X=9.075 $Y=1.5 $X2=0 $Y2=0
cc_254 N_S_c_281_n N_A_1418_21#_c_408_n 0.0160454f $X=7.045 $Y=1.68 $X2=0 $Y2=0
cc_255 N_S_c_276_n N_A_1418_21#_c_409_n 0.00202605f $X=8.885 $Y=1.185 $X2=0
+ $Y2=0
cc_256 N_S_c_277_n N_A_1418_21#_c_409_n 2.31177e-19 $X=9.075 $Y=1.665 $X2=0
+ $Y2=0
cc_257 N_S_c_278_n N_A_1418_21#_c_409_n 0.00605901f $X=9.075 $Y=1.5 $X2=0 $Y2=0
cc_258 N_S_c_276_n N_A_1418_21#_c_410_n 0.0156693f $X=8.885 $Y=1.185 $X2=0 $Y2=0
cc_259 N_S_c_277_n N_A_1418_21#_c_410_n 0.00972587f $X=9.075 $Y=1.665 $X2=0
+ $Y2=0
cc_260 N_S_c_288_n N_A_1418_21#_c_410_n 0.00393234f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_261 N_S_c_278_n N_A_1418_21#_c_410_n 0.0240873f $X=9.075 $Y=1.5 $X2=0 $Y2=0
cc_262 N_S_c_277_n N_A_1418_21#_c_418_n 0.0017498f $X=9.075 $Y=1.665 $X2=0 $Y2=0
cc_263 N_S_c_276_n N_A_1418_21#_c_412_n 3.54886e-19 $X=8.885 $Y=1.185 $X2=0
+ $Y2=0
cc_264 N_S_c_277_n N_A_1418_21#_c_412_n 0.0127183f $X=9.075 $Y=1.665 $X2=0 $Y2=0
cc_265 N_S_M1015_g N_A_1418_21#_c_412_n 0.00345176f $X=9.075 $Y=2.465 $X2=0
+ $Y2=0
cc_266 N_S_c_278_n N_A_1418_21#_c_412_n 0.0332794f $X=9.075 $Y=1.5 $X2=0 $Y2=0
cc_267 N_S_c_277_n N_A_1418_21#_c_413_n 0.0142424f $X=9.075 $Y=1.665 $X2=0 $Y2=0
cc_268 N_S_M1015_g N_A_1418_21#_c_413_n 0.0234664f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_269 N_S_c_288_n N_A_1418_21#_c_413_n 0.0134225f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_270 N_S_c_278_n N_A_1418_21#_c_413_n 0.00475226f $X=9.075 $Y=1.5 $X2=0 $Y2=0
cc_271 N_S_c_280_n N_A_1418_21#_c_413_n 0.0474369f $X=6.735 $Y=1.51 $X2=0 $Y2=0
cc_272 N_S_c_281_n N_A_1418_21#_c_413_n 0.00754377f $X=7.045 $Y=1.68 $X2=0 $Y2=0
cc_273 S N_Y_c_518_n 0.0353042f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_274 N_S_M1000_g N_A_126_367#_c_622_n 0.0167022f $X=5.435 $Y=2.465 $X2=0 $Y2=0
cc_275 N_S_M1004_g N_A_126_367#_c_622_n 0.0126273f $X=5.865 $Y=2.465 $X2=0 $Y2=0
cc_276 N_S_M1017_g N_A_126_367#_c_622_n 0.0127182f $X=6.295 $Y=2.465 $X2=0 $Y2=0
cc_277 N_S_c_280_n N_A_126_367#_c_622_n 0.00161383f $X=6.735 $Y=1.51 $X2=0 $Y2=0
cc_278 S N_A_126_367#_c_623_n 3.97915e-19 $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_279 S N_A_126_367#_c_624_n 0.164846f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_280 N_S_c_288_n N_A_470_367#_M1008_s 0.00176891f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_281 N_S_c_288_n N_A_470_367#_M1021_s 0.00176461f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_282 N_S_c_288_n N_A_470_367#_c_676_n 0.0401176f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_283 N_S_c_288_n N_A_470_367#_c_677_n 0.0179918f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_284 N_S_M1000_g N_A_470_367#_c_670_n 0.00387508f $X=5.435 $Y=2.465 $X2=0
+ $Y2=0
cc_285 N_S_M1000_g N_A_470_367#_c_679_n 0.0135488f $X=5.435 $Y=2.465 $X2=0 $Y2=0
cc_286 N_S_M1004_g N_A_470_367#_c_679_n 0.0116931f $X=5.865 $Y=2.465 $X2=0 $Y2=0
cc_287 N_S_M1017_g N_A_470_367#_c_679_n 0.0118131f $X=6.295 $Y=2.465 $X2=0 $Y2=0
cc_288 N_S_M1026_g N_A_470_367#_c_679_n 0.0140451f $X=6.745 $Y=2.465 $X2=0 $Y2=0
cc_289 S N_A_470_367#_c_679_n 0.00527679f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_290 N_S_M1026_g N_A_470_367#_c_684_n 0.00747147f $X=6.745 $Y=2.465 $X2=0
+ $Y2=0
cc_291 N_S_c_281_n N_A_470_367#_c_684_n 0.0401176f $X=7.045 $Y=1.68 $X2=0 $Y2=0
cc_292 N_S_c_281_n N_VPWR_M1026_d 0.00179873f $X=7.045 $Y=1.68 $X2=0 $Y2=0
cc_293 N_S_c_288_n N_VPWR_M1011_d 0.00395655f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_294 N_S_c_288_n N_VPWR_M1022_d 0.0010795f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_295 N_S_c_278_n N_VPWR_M1022_d 9.94388e-19 $X=9.075 $Y=1.5 $X2=0 $Y2=0
cc_296 N_S_M1000_g N_VPWR_c_740_n 0.00146468f $X=5.435 $Y=2.465 $X2=0 $Y2=0
cc_297 N_S_M1004_g N_VPWR_c_740_n 0.0088668f $X=5.865 $Y=2.465 $X2=0 $Y2=0
cc_298 N_S_M1017_g N_VPWR_c_740_n 0.00847294f $X=6.295 $Y=2.465 $X2=0 $Y2=0
cc_299 N_S_M1026_g N_VPWR_c_740_n 0.0011721f $X=6.745 $Y=2.465 $X2=0 $Y2=0
cc_300 N_S_M1017_g N_VPWR_c_741_n 0.0011721f $X=6.295 $Y=2.465 $X2=0 $Y2=0
cc_301 N_S_M1026_g N_VPWR_c_741_n 0.00843718f $X=6.745 $Y=2.465 $X2=0 $Y2=0
cc_302 N_S_c_277_n N_VPWR_c_743_n 2.78893e-19 $X=9.075 $Y=1.665 $X2=0 $Y2=0
cc_303 N_S_M1015_g N_VPWR_c_743_n 0.0156403f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_304 N_S_c_288_n N_VPWR_c_743_n 0.00799911f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_305 N_S_c_278_n N_VPWR_c_743_n 0.00942265f $X=9.075 $Y=1.5 $X2=0 $Y2=0
cc_306 N_S_M1000_g N_VPWR_c_745_n 0.00428022f $X=5.435 $Y=2.465 $X2=0 $Y2=0
cc_307 N_S_M1004_g N_VPWR_c_745_n 0.00355956f $X=5.865 $Y=2.465 $X2=0 $Y2=0
cc_308 N_S_M1017_g N_VPWR_c_746_n 0.00355956f $X=6.295 $Y=2.465 $X2=0 $Y2=0
cc_309 N_S_M1026_g N_VPWR_c_746_n 0.00355956f $X=6.745 $Y=2.465 $X2=0 $Y2=0
cc_310 N_S_M1015_g N_VPWR_c_749_n 0.00486043f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_311 N_S_M1000_g N_VPWR_c_739_n 0.00744823f $X=5.435 $Y=2.465 $X2=0 $Y2=0
cc_312 N_S_M1004_g N_VPWR_c_739_n 0.00423262f $X=5.865 $Y=2.465 $X2=0 $Y2=0
cc_313 N_S_M1017_g N_VPWR_c_739_n 0.00428782f $X=6.295 $Y=2.465 $X2=0 $Y2=0
cc_314 N_S_M1026_g N_VPWR_c_739_n 0.00428782f $X=6.745 $Y=2.465 $X2=0 $Y2=0
cc_315 N_S_M1015_g N_VPWR_c_739_n 0.00922386f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_316 N_S_M1000_g N_VPWR_c_751_n 0.00637672f $X=5.435 $Y=2.465 $X2=0 $Y2=0
cc_317 S N_A_110_69#_c_861_n 3.13109e-19 $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_318 N_S_M1010_g N_A_110_69#_c_863_n 0.0125321f $X=5.445 $Y=0.655 $X2=0 $Y2=0
cc_319 N_S_M1012_g N_A_110_69#_c_863_n 0.0104915f $X=5.875 $Y=0.655 $X2=0 $Y2=0
cc_320 N_S_M1031_g N_A_110_69#_c_863_n 0.0104915f $X=6.305 $Y=0.655 $X2=0 $Y2=0
cc_321 N_S_M1033_g N_A_110_69#_c_863_n 0.0142626f $X=6.735 $Y=0.655 $X2=0 $Y2=0
cc_322 N_S_c_288_n N_A_110_69#_c_863_n 0.00349173f $X=8.855 $Y=1.86 $X2=0 $Y2=0
cc_323 S N_A_110_69#_c_863_n 0.188221f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_324 N_S_c_280_n N_A_110_69#_c_863_n 0.00749652f $X=6.735 $Y=1.51 $X2=0 $Y2=0
cc_325 S N_A_110_69#_c_864_n 0.015193f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_326 N_S_M1010_g N_A_470_69#_c_950_n 0.00265741f $X=5.445 $Y=0.655 $X2=0 $Y2=0
cc_327 N_S_M1010_g N_A_470_69#_c_951_n 0.0107124f $X=5.445 $Y=0.655 $X2=0 $Y2=0
cc_328 N_S_M1010_g N_A_470_69#_c_959_n 0.00592348f $X=5.445 $Y=0.655 $X2=0 $Y2=0
cc_329 N_S_M1012_g N_A_470_69#_c_959_n 0.00545927f $X=5.875 $Y=0.655 $X2=0 $Y2=0
cc_330 N_S_M1031_g N_A_470_69#_c_959_n 4.9709e-19 $X=6.305 $Y=0.655 $X2=0 $Y2=0
cc_331 N_S_M1012_g N_A_470_69#_c_962_n 0.0088372f $X=5.875 $Y=0.655 $X2=0 $Y2=0
cc_332 N_S_M1031_g N_A_470_69#_c_962_n 0.00955415f $X=6.305 $Y=0.655 $X2=0 $Y2=0
cc_333 N_S_M1033_g N_A_470_69#_c_962_n 0.00205832f $X=6.735 $Y=0.655 $X2=0 $Y2=0
cc_334 N_S_M1012_g N_A_470_69#_c_965_n 5.22552e-19 $X=5.875 $Y=0.655 $X2=0 $Y2=0
cc_335 N_S_M1031_g N_A_470_69#_c_965_n 0.00627821f $X=6.305 $Y=0.655 $X2=0 $Y2=0
cc_336 N_S_M1033_g N_A_470_69#_c_965_n 0.00503721f $X=6.735 $Y=0.655 $X2=0 $Y2=0
cc_337 N_S_M1010_g N_A_470_69#_c_968_n 7.14816e-19 $X=5.445 $Y=0.655 $X2=0 $Y2=0
cc_338 N_S_M1012_g N_A_470_69#_c_968_n 7.14816e-19 $X=5.875 $Y=0.655 $X2=0 $Y2=0
cc_339 N_S_M1010_g N_VGND_c_1008_n 0.00322927f $X=5.445 $Y=0.655 $X2=0 $Y2=0
cc_340 N_S_M1010_g N_VGND_c_1009_n 0.00430034f $X=5.445 $Y=0.655 $X2=0 $Y2=0
cc_341 N_S_M1012_g N_VGND_c_1009_n 0.00430034f $X=5.875 $Y=0.655 $X2=0 $Y2=0
cc_342 N_S_M1012_g N_VGND_c_1010_n 0.00153274f $X=5.875 $Y=0.655 $X2=0 $Y2=0
cc_343 N_S_M1031_g N_VGND_c_1010_n 0.00153274f $X=6.305 $Y=0.655 $X2=0 $Y2=0
cc_344 N_S_M1033_g N_VGND_c_1011_n 0.00157435f $X=6.735 $Y=0.655 $X2=0 $Y2=0
cc_345 N_S_c_276_n N_VGND_c_1013_n 0.0116893f $X=8.885 $Y=1.185 $X2=0 $Y2=0
cc_346 N_S_M1031_g N_VGND_c_1020_n 0.00427134f $X=6.305 $Y=0.655 $X2=0 $Y2=0
cc_347 N_S_M1033_g N_VGND_c_1020_n 0.0054895f $X=6.735 $Y=0.655 $X2=0 $Y2=0
cc_348 N_S_c_276_n N_VGND_c_1021_n 0.00486043f $X=8.885 $Y=1.185 $X2=0 $Y2=0
cc_349 N_S_M1010_g N_VGND_c_1022_n 0.00720467f $X=5.445 $Y=0.655 $X2=0 $Y2=0
cc_350 N_S_M1012_g N_VGND_c_1022_n 0.00590497f $X=5.875 $Y=0.655 $X2=0 $Y2=0
cc_351 N_S_M1031_g N_VGND_c_1022_n 0.0058261f $X=6.305 $Y=0.655 $X2=0 $Y2=0
cc_352 N_S_M1033_g N_VGND_c_1022_n 0.00979102f $X=6.735 $Y=0.655 $X2=0 $Y2=0
cc_353 N_S_c_276_n N_VGND_c_1022_n 0.00934144f $X=8.885 $Y=1.185 $X2=0 $Y2=0
cc_354 N_A_1418_21#_c_415_n N_A_470_367#_c_686_n 0.00469909f $X=7.605 $Y=1.725
+ $X2=0 $Y2=0
cc_355 N_A_1418_21#_c_415_n N_A_470_367#_c_676_n 0.0112141f $X=7.605 $Y=1.725
+ $X2=0 $Y2=0
cc_356 N_A_1418_21#_c_416_n N_A_470_367#_c_676_n 0.0112141f $X=8.195 $Y=1.725
+ $X2=0 $Y2=0
cc_357 N_A_1418_21#_c_416_n N_A_470_367#_c_677_n 0.00103713f $X=8.195 $Y=1.725
+ $X2=0 $Y2=0
cc_358 N_A_1418_21#_c_417_n N_A_470_367#_c_677_n 0.00216754f $X=8.625 $Y=1.725
+ $X2=0 $Y2=0
cc_359 N_A_1418_21#_c_415_n N_A_470_367#_c_691_n 6.57491e-19 $X=7.605 $Y=1.725
+ $X2=0 $Y2=0
cc_360 N_A_1418_21#_c_416_n N_A_470_367#_c_691_n 0.0105817f $X=8.195 $Y=1.725
+ $X2=0 $Y2=0
cc_361 N_A_1418_21#_c_417_n N_A_470_367#_c_691_n 0.00810575f $X=8.625 $Y=1.725
+ $X2=0 $Y2=0
cc_362 N_A_1418_21#_c_414_n N_A_470_367#_c_684_n 0.0186874f $X=7.175 $Y=1.725
+ $X2=0 $Y2=0
cc_363 N_A_1418_21#_c_415_n N_A_470_367#_c_684_n 0.00725838f $X=7.605 $Y=1.725
+ $X2=0 $Y2=0
cc_364 N_A_1418_21#_c_416_n N_A_470_367#_c_684_n 5.80303e-19 $X=8.195 $Y=1.725
+ $X2=0 $Y2=0
cc_365 N_A_1418_21#_c_414_n N_VPWR_c_741_n 0.00686775f $X=7.175 $Y=1.725 $X2=0
+ $Y2=0
cc_366 N_A_1418_21#_c_415_n N_VPWR_c_741_n 4.90758e-19 $X=7.605 $Y=1.725 $X2=0
+ $Y2=0
cc_367 N_A_1418_21#_c_415_n N_VPWR_c_742_n 0.00566219f $X=7.605 $Y=1.725 $X2=0
+ $Y2=0
cc_368 N_A_1418_21#_c_416_n N_VPWR_c_742_n 0.00708091f $X=8.195 $Y=1.725 $X2=0
+ $Y2=0
cc_369 N_A_1418_21#_c_417_n N_VPWR_c_743_n 0.00294729f $X=8.625 $Y=1.725 $X2=0
+ $Y2=0
cc_370 N_A_1418_21#_c_414_n N_VPWR_c_747_n 0.00355956f $X=7.175 $Y=1.725 $X2=0
+ $Y2=0
cc_371 N_A_1418_21#_c_415_n N_VPWR_c_747_n 0.00533193f $X=7.605 $Y=1.725 $X2=0
+ $Y2=0
cc_372 N_A_1418_21#_c_416_n N_VPWR_c_748_n 0.00534242f $X=8.195 $Y=1.725 $X2=0
+ $Y2=0
cc_373 N_A_1418_21#_c_417_n N_VPWR_c_748_n 0.00549284f $X=8.625 $Y=1.725 $X2=0
+ $Y2=0
cc_374 N_A_1418_21#_c_419_n N_VPWR_c_749_n 0.0217539f $X=9.29 $Y=2.01 $X2=0
+ $Y2=0
cc_375 N_A_1418_21#_M1015_d N_VPWR_c_739_n 0.00371702f $X=9.15 $Y=1.835 $X2=0
+ $Y2=0
cc_376 N_A_1418_21#_c_414_n N_VPWR_c_739_n 0.00415754f $X=7.175 $Y=1.725 $X2=0
+ $Y2=0
cc_377 N_A_1418_21#_c_415_n N_VPWR_c_739_n 0.00987153f $X=7.605 $Y=1.725 $X2=0
+ $Y2=0
cc_378 N_A_1418_21#_c_416_n N_VPWR_c_739_n 0.00991768f $X=8.195 $Y=1.725 $X2=0
+ $Y2=0
cc_379 N_A_1418_21#_c_417_n N_VPWR_c_739_n 0.00983896f $X=8.625 $Y=1.725 $X2=0
+ $Y2=0
cc_380 N_A_1418_21#_c_419_n N_VPWR_c_739_n 0.0121687f $X=9.29 $Y=2.01 $X2=0
+ $Y2=0
cc_381 N_A_1418_21#_M1006_g N_A_110_69#_c_863_n 0.0159373f $X=7.165 $Y=0.655
+ $X2=0 $Y2=0
cc_382 N_A_1418_21#_c_408_n N_A_110_69#_c_863_n 0.00423349f $X=8.505 $Y=1.51
+ $X2=0 $Y2=0
cc_383 N_A_1418_21#_M1009_g N_A_110_69#_c_865_n 0.0143861f $X=7.595 $Y=0.655
+ $X2=0 $Y2=0
cc_384 N_A_1418_21#_M1027_g N_A_110_69#_c_865_n 0.013983f $X=8.025 $Y=0.655
+ $X2=0 $Y2=0
cc_385 N_A_1418_21#_M1028_g N_A_110_69#_c_865_n 0.00139645f $X=8.455 $Y=0.655
+ $X2=0 $Y2=0
cc_386 N_A_1418_21#_c_408_n N_A_110_69#_c_865_n 0.0625611f $X=8.505 $Y=1.51
+ $X2=0 $Y2=0
cc_387 N_A_1418_21#_c_409_n N_A_110_69#_c_865_n 0.00641961f $X=8.59 $Y=1.415
+ $X2=0 $Y2=0
cc_388 N_A_1418_21#_c_486_p N_A_110_69#_c_865_n 0.00797592f $X=8.675 $Y=1.075
+ $X2=0 $Y2=0
cc_389 N_A_1418_21#_c_413_n N_A_110_69#_c_865_n 0.00550397f $X=8.455 $Y=1.535
+ $X2=0 $Y2=0
cc_390 N_A_1418_21#_c_408_n N_A_110_69#_c_866_n 0.0154426f $X=8.505 $Y=1.51
+ $X2=0 $Y2=0
cc_391 N_A_1418_21#_c_413_n N_A_110_69#_c_866_n 0.00264307f $X=8.455 $Y=1.535
+ $X2=0 $Y2=0
cc_392 N_A_1418_21#_c_410_n N_VGND_M1028_d 8.1997e-19 $X=9.005 $Y=1.075 $X2=0
+ $Y2=0
cc_393 N_A_1418_21#_c_486_p N_VGND_M1028_d 9.71089e-19 $X=8.675 $Y=1.075 $X2=0
+ $Y2=0
cc_394 N_A_1418_21#_M1006_g N_VGND_c_1011_n 0.0105367f $X=7.165 $Y=0.655 $X2=0
+ $Y2=0
cc_395 N_A_1418_21#_M1009_g N_VGND_c_1011_n 6.2955e-19 $X=7.595 $Y=0.655 $X2=0
+ $Y2=0
cc_396 N_A_1418_21#_M1006_g N_VGND_c_1012_n 6.05521e-19 $X=7.165 $Y=0.655 $X2=0
+ $Y2=0
cc_397 N_A_1418_21#_M1009_g N_VGND_c_1012_n 0.00996875f $X=7.595 $Y=0.655 $X2=0
+ $Y2=0
cc_398 N_A_1418_21#_M1027_g N_VGND_c_1012_n 0.00996875f $X=8.025 $Y=0.655 $X2=0
+ $Y2=0
cc_399 N_A_1418_21#_M1028_g N_VGND_c_1012_n 6.05521e-19 $X=8.455 $Y=0.655 $X2=0
+ $Y2=0
cc_400 N_A_1418_21#_M1027_g N_VGND_c_1013_n 6.0835e-19 $X=8.025 $Y=0.655 $X2=0
+ $Y2=0
cc_401 N_A_1418_21#_M1028_g N_VGND_c_1013_n 0.00993814f $X=8.455 $Y=0.655 $X2=0
+ $Y2=0
cc_402 N_A_1418_21#_c_410_n N_VGND_c_1013_n 0.00812698f $X=9.005 $Y=1.075 $X2=0
+ $Y2=0
cc_403 N_A_1418_21#_c_486_p N_VGND_c_1013_n 0.00985537f $X=8.675 $Y=1.075 $X2=0
+ $Y2=0
cc_404 N_A_1418_21#_M1006_g N_VGND_c_1016_n 0.00486043f $X=7.165 $Y=0.655 $X2=0
+ $Y2=0
cc_405 N_A_1418_21#_M1009_g N_VGND_c_1016_n 0.00486043f $X=7.595 $Y=0.655 $X2=0
+ $Y2=0
cc_406 N_A_1418_21#_M1027_g N_VGND_c_1018_n 0.00486043f $X=8.025 $Y=0.655 $X2=0
+ $Y2=0
cc_407 N_A_1418_21#_M1028_g N_VGND_c_1018_n 0.00486043f $X=8.455 $Y=0.655 $X2=0
+ $Y2=0
cc_408 N_A_1418_21#_c_506_p N_VGND_c_1021_n 0.0135387f $X=9.1 $Y=0.42 $X2=0
+ $Y2=0
cc_409 N_A_1418_21#_M1003_d N_VGND_c_1022_n 0.00444756f $X=8.96 $Y=0.235 $X2=0
+ $Y2=0
cc_410 N_A_1418_21#_M1006_g N_VGND_c_1022_n 0.00824727f $X=7.165 $Y=0.655 $X2=0
+ $Y2=0
cc_411 N_A_1418_21#_M1009_g N_VGND_c_1022_n 0.00824727f $X=7.595 $Y=0.655 $X2=0
+ $Y2=0
cc_412 N_A_1418_21#_M1027_g N_VGND_c_1022_n 0.00824727f $X=8.025 $Y=0.655 $X2=0
+ $Y2=0
cc_413 N_A_1418_21#_M1028_g N_VGND_c_1022_n 0.00824727f $X=8.455 $Y=0.655 $X2=0
+ $Y2=0
cc_414 N_A_1418_21#_c_506_p N_VGND_c_1022_n 0.00769778f $X=9.1 $Y=0.42 $X2=0
+ $Y2=0
cc_415 N_Y_c_531_n N_A_126_367#_M1001_s 0.00341063f $X=1.115 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_416 N_Y_c_521_n N_A_126_367#_M1016_s 0.00337374f $X=4.095 $Y=2.02 $X2=0 $Y2=0
cc_417 N_Y_c_531_n N_A_126_367#_c_640_n 0.0129246f $X=1.115 $Y=2.015 $X2=0 $Y2=0
cc_418 N_Y_M1014_d N_A_126_367#_c_625_n 0.00380104f $X=1.06 $Y=1.835 $X2=0 $Y2=0
cc_419 N_Y_c_521_n N_A_126_367#_c_625_n 0.00322336f $X=4.095 $Y=2.02 $X2=0 $Y2=0
cc_420 N_Y_c_548_n N_A_126_367#_c_625_n 0.0123171f $X=1.2 $Y=2.095 $X2=0 $Y2=0
cc_421 N_Y_c_521_n N_A_126_367#_c_644_n 0.0135413f $X=4.095 $Y=2.02 $X2=0 $Y2=0
cc_422 N_Y_M1025_d N_A_126_367#_c_623_n 0.00814987f $X=1.92 $Y=1.835 $X2=0 $Y2=0
cc_423 N_Y_M1013_d N_A_126_367#_c_623_n 0.00345391f $X=2.78 $Y=1.835 $X2=0 $Y2=0
cc_424 N_Y_M1032_d N_A_126_367#_c_623_n 0.00509067f $X=3.64 $Y=1.835 $X2=0 $Y2=0
cc_425 N_Y_c_521_n N_A_126_367#_c_623_n 0.143676f $X=4.095 $Y=2.02 $X2=0 $Y2=0
cc_426 N_Y_c_521_n N_A_126_367#_c_624_n 0.00935508f $X=4.095 $Y=2.02 $X2=0 $Y2=0
cc_427 N_Y_c_521_n N_A_470_367#_M1007_s 0.00384139f $X=4.095 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_428 N_Y_c_521_n N_A_470_367#_M1023_s 0.00334197f $X=4.095 $Y=2.02 $X2=0 $Y2=0
cc_429 N_Y_M1013_d N_A_470_367#_c_671_n 0.00342769f $X=2.78 $Y=1.835 $X2=0 $Y2=0
cc_430 N_Y_M1032_d N_A_470_367#_c_669_n 0.00617422f $X=3.64 $Y=1.835 $X2=0 $Y2=0
cc_431 N_Y_c_590_p N_VPWR_c_744_n 0.00699362f $X=0.34 $Y=2.775 $X2=0 $Y2=0
cc_432 N_Y_M1001_d N_VPWR_c_739_n 0.00495509f $X=0.215 $Y=1.835 $X2=0 $Y2=0
cc_433 N_Y_M1014_d N_VPWR_c_739_n 0.00240554f $X=1.06 $Y=1.835 $X2=0 $Y2=0
cc_434 N_Y_M1025_d N_VPWR_c_739_n 0.0119922f $X=1.92 $Y=1.835 $X2=0 $Y2=0
cc_435 N_Y_M1013_d N_VPWR_c_739_n 0.00225186f $X=2.78 $Y=1.835 $X2=0 $Y2=0
cc_436 N_Y_M1032_d N_VPWR_c_739_n 0.00272831f $X=3.64 $Y=1.835 $X2=0 $Y2=0
cc_437 N_Y_c_590_p N_VPWR_c_739_n 0.00676664f $X=0.34 $Y=2.775 $X2=0 $Y2=0
cc_438 N_Y_c_514_n N_A_110_69#_M1005_d 0.00176461f $X=1.035 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_439 N_Y_c_516_n N_A_110_69#_M1024_d 0.00179194f $X=1.895 $Y=1.105 $X2=0 $Y2=0
cc_440 N_Y_c_514_n N_A_110_69#_c_867_n 0.0170147f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_441 N_Y_M1020_s N_A_110_69#_c_859_n 0.00269203f $X=0.98 $Y=0.345 $X2=0 $Y2=0
cc_442 N_Y_c_514_n N_A_110_69#_c_859_n 0.00292119f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_443 N_Y_c_516_n N_A_110_69#_c_859_n 0.0036223f $X=1.895 $Y=1.105 $X2=0 $Y2=0
cc_444 N_Y_c_519_n N_A_110_69#_c_859_n 0.0196117f $X=1.2 $Y=0.72 $X2=0 $Y2=0
cc_445 N_Y_c_513_n N_A_110_69#_c_860_n 0.00593039f $X=0.26 $Y=0.49 $X2=0 $Y2=0
cc_446 N_Y_c_516_n N_A_110_69#_c_875_n 0.01562f $X=1.895 $Y=1.105 $X2=0 $Y2=0
cc_447 N_Y_M1029_s N_A_110_69#_c_861_n 0.00462143f $X=1.92 $Y=0.345 $X2=0 $Y2=0
cc_448 N_Y_M1018_d N_A_110_69#_c_861_n 0.00336136f $X=2.94 $Y=0.345 $X2=0 $Y2=0
cc_449 N_Y_M1030_d N_A_110_69#_c_861_n 0.00572184f $X=3.96 $Y=0.345 $X2=0 $Y2=0
cc_450 N_Y_c_516_n N_A_110_69#_c_861_n 0.00701411f $X=1.895 $Y=1.105 $X2=0 $Y2=0
cc_451 N_Y_c_560_n N_A_110_69#_c_861_n 0.103149f $X=4.095 $Y=1.065 $X2=0 $Y2=0
cc_452 N_Y_c_517_n N_A_110_69#_c_861_n 0.013893f $X=4.18 $Y=1.165 $X2=0 $Y2=0
cc_453 N_Y_c_520_n N_A_110_69#_c_861_n 0.0188996f $X=2.06 $Y=1.06 $X2=0 $Y2=0
cc_454 N_Y_c_517_n N_A_110_69#_c_862_n 0.00888518f $X=4.18 $Y=1.165 $X2=0 $Y2=0
cc_455 N_Y_c_517_n N_A_110_69#_c_864_n 0.00809565f $X=4.18 $Y=1.165 $X2=0 $Y2=0
cc_456 N_Y_c_518_n N_A_110_69#_c_864_n 0.00645203f $X=4.18 $Y=1.93 $X2=0 $Y2=0
cc_457 N_Y_c_560_n N_A_470_69#_M1002_s 0.00777701f $X=4.095 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_458 N_Y_c_560_n N_A_470_69#_M1019_s 0.00726934f $X=4.095 $Y=1.065 $X2=0 $Y2=0
cc_459 N_Y_M1018_d N_A_470_69#_c_949_n 0.00177781f $X=2.94 $Y=0.345 $X2=0 $Y2=0
cc_460 N_Y_M1030_d N_A_470_69#_c_949_n 0.00307529f $X=3.96 $Y=0.345 $X2=0 $Y2=0
cc_461 N_Y_c_513_n N_VGND_c_1014_n 0.00932149f $X=0.26 $Y=0.49 $X2=0 $Y2=0
cc_462 N_Y_c_513_n N_VGND_c_1022_n 0.00704609f $X=0.26 $Y=0.49 $X2=0 $Y2=0
cc_463 N_A_126_367#_c_623_n N_A_470_367#_M1007_s 0.00345391f $X=4.445 $Y=2.232
+ $X2=-0.19 $Y2=1.655
cc_464 N_A_126_367#_c_623_n N_A_470_367#_M1023_s 0.00345391f $X=4.445 $Y=2.232
+ $X2=0 $Y2=0
cc_465 N_A_126_367#_c_623_n N_A_470_367#_c_671_n 0.0705349f $X=4.445 $Y=2.232
+ $X2=0 $Y2=0
cc_466 N_A_126_367#_c_622_n N_A_470_367#_c_669_n 0.00970899f $X=6.51 $Y=2.17
+ $X2=0 $Y2=0
cc_467 N_A_126_367#_c_624_n N_A_470_367#_c_705_n 0.0705349f $X=4.615 $Y=2.232
+ $X2=0 $Y2=0
cc_468 N_A_126_367#_c_622_n N_A_470_367#_c_670_n 0.0139246f $X=6.51 $Y=2.17
+ $X2=0 $Y2=0
cc_469 N_A_126_367#_M1000_s N_A_470_367#_c_679_n 0.00472599f $X=5.51 $Y=1.835
+ $X2=0 $Y2=0
cc_470 N_A_126_367#_M1017_s N_A_470_367#_c_679_n 0.00529539f $X=6.37 $Y=1.835
+ $X2=0 $Y2=0
cc_471 N_A_126_367#_c_622_n N_A_470_367#_c_679_n 0.0974402f $X=6.51 $Y=2.17
+ $X2=0 $Y2=0
cc_472 N_A_126_367#_c_622_n N_VPWR_M1000_d 0.0114006f $X=6.51 $Y=2.17 $X2=-0.19
+ $Y2=1.655
cc_473 N_A_126_367#_c_622_n N_VPWR_M1004_d 0.00343187f $X=6.51 $Y=2.17 $X2=0
+ $Y2=0
cc_474 N_A_126_367#_c_625_n N_VPWR_c_744_n 0.0270087f $X=1.525 $Y=2.865 $X2=0
+ $Y2=0
cc_475 N_A_126_367#_c_662_p N_VPWR_c_744_n 0.0073172f $X=0.875 $Y=2.865 $X2=0
+ $Y2=0
cc_476 N_A_126_367#_M1001_s N_VPWR_c_739_n 0.00360224f $X=0.63 $Y=1.835 $X2=0
+ $Y2=0
cc_477 N_A_126_367#_M1016_s N_VPWR_c_739_n 0.00360224f $X=1.49 $Y=1.835 $X2=0
+ $Y2=0
cc_478 N_A_126_367#_M1000_s N_VPWR_c_739_n 0.00333718f $X=5.51 $Y=1.835 $X2=0
+ $Y2=0
cc_479 N_A_126_367#_M1017_s N_VPWR_c_739_n 0.00357554f $X=6.37 $Y=1.835 $X2=0
+ $Y2=0
cc_480 N_A_126_367#_c_625_n N_VPWR_c_739_n 0.0286432f $X=1.525 $Y=2.865 $X2=0
+ $Y2=0
cc_481 N_A_126_367#_c_662_p N_VPWR_c_739_n 0.00761013f $X=0.875 $Y=2.865 $X2=0
+ $Y2=0
cc_482 N_A_470_367#_c_670_n N_VPWR_M1000_d 0.00227007f $X=4.88 $Y=2.59 $X2=-0.19
+ $Y2=1.655
cc_483 N_A_470_367#_c_679_n N_VPWR_M1000_d 0.0106494f $X=6.88 $Y=2.395 $X2=-0.19
+ $Y2=1.655
cc_484 N_A_470_367#_c_679_n N_VPWR_M1004_d 0.00347121f $X=6.88 $Y=2.395 $X2=0
+ $Y2=0
cc_485 N_A_470_367#_c_684_n N_VPWR_M1026_d 0.00843151f $X=7.565 $Y=2.395 $X2=0
+ $Y2=0
cc_486 N_A_470_367#_c_676_n N_VPWR_M1011_d 0.00728226f $X=8.235 $Y=2.2 $X2=0
+ $Y2=0
cc_487 N_A_470_367#_c_679_n N_VPWR_c_740_n 0.016098f $X=6.88 $Y=2.395 $X2=0
+ $Y2=0
cc_488 N_A_470_367#_c_679_n N_VPWR_c_741_n 0.017195f $X=6.88 $Y=2.395 $X2=0
+ $Y2=0
cc_489 N_A_470_367#_c_676_n N_VPWR_c_742_n 0.0265229f $X=8.235 $Y=2.2 $X2=0
+ $Y2=0
cc_490 N_A_470_367#_c_671_n N_VPWR_c_744_n 0.0630289f $X=3.233 $Y=2.852 $X2=0
+ $Y2=0
cc_491 N_A_470_367#_c_669_n N_VPWR_c_744_n 0.0296608f $X=4.795 $Y=2.715 $X2=0
+ $Y2=0
cc_492 N_A_470_367#_c_670_n N_VPWR_c_744_n 0.00347758f $X=4.88 $Y=2.59 $X2=0
+ $Y2=0
cc_493 N_A_470_367#_c_679_n N_VPWR_c_745_n 0.00919442f $X=6.88 $Y=2.395 $X2=0
+ $Y2=0
cc_494 N_A_470_367#_c_679_n N_VPWR_c_746_n 0.00804859f $X=6.88 $Y=2.395 $X2=0
+ $Y2=0
cc_495 N_A_470_367#_c_686_n N_VPWR_c_747_n 0.0148797f $X=7.39 $Y=2.9 $X2=0 $Y2=0
cc_496 N_A_470_367#_c_684_n N_VPWR_c_747_n 0.00253472f $X=7.565 $Y=2.395 $X2=0
+ $Y2=0
cc_497 N_A_470_367#_c_691_n N_VPWR_c_748_n 0.0184348f $X=8.41 $Y=2.96 $X2=0
+ $Y2=0
cc_498 N_A_470_367#_M1007_s N_VPWR_c_739_n 0.0034694f $X=2.35 $Y=1.835 $X2=0
+ $Y2=0
cc_499 N_A_470_367#_M1023_s N_VPWR_c_739_n 0.00232694f $X=3.21 $Y=1.835 $X2=0
+ $Y2=0
cc_500 N_A_470_367#_M1008_s N_VPWR_c_739_n 0.00241223f $X=7.25 $Y=1.835 $X2=0
+ $Y2=0
cc_501 N_A_470_367#_M1021_s N_VPWR_c_739_n 0.00223819f $X=8.27 $Y=1.835 $X2=0
+ $Y2=0
cc_502 N_A_470_367#_c_671_n N_VPWR_c_739_n 0.0397493f $X=3.233 $Y=2.852 $X2=0
+ $Y2=0
cc_503 N_A_470_367#_c_669_n N_VPWR_c_739_n 0.0407555f $X=4.795 $Y=2.715 $X2=0
+ $Y2=0
cc_504 N_A_470_367#_c_686_n N_VPWR_c_739_n 0.0099921f $X=7.39 $Y=2.9 $X2=0 $Y2=0
cc_505 N_A_470_367#_c_691_n N_VPWR_c_739_n 0.0126656f $X=8.41 $Y=2.96 $X2=0
+ $Y2=0
cc_506 N_A_470_367#_c_670_n N_VPWR_c_739_n 0.00473969f $X=4.88 $Y=2.59 $X2=0
+ $Y2=0
cc_507 N_A_470_367#_c_679_n N_VPWR_c_739_n 0.0357396f $X=6.88 $Y=2.395 $X2=0
+ $Y2=0
cc_508 N_A_470_367#_c_684_n N_VPWR_c_739_n 0.00443271f $X=7.565 $Y=2.395 $X2=0
+ $Y2=0
cc_509 N_A_470_367#_c_670_n N_VPWR_c_751_n 0.00181629f $X=4.88 $Y=2.59 $X2=0
+ $Y2=0
cc_510 N_A_470_367#_c_679_n N_VPWR_c_751_n 0.0140043f $X=6.88 $Y=2.395 $X2=0
+ $Y2=0
cc_511 N_A_110_69#_c_861_n N_A_470_69#_M1002_s 0.00727881f $X=4.445 $Y=0.71
+ $X2=-0.19 $Y2=-0.245
cc_512 N_A_110_69#_c_861_n N_A_470_69#_M1019_s 0.00727881f $X=4.445 $Y=0.71
+ $X2=0 $Y2=0
cc_513 N_A_110_69#_c_859_n N_A_470_69#_c_949_n 0.00454351f $X=1.535 $Y=0.355
+ $X2=0 $Y2=0
cc_514 N_A_110_69#_c_861_n N_A_470_69#_c_949_n 0.130081f $X=4.445 $Y=0.71 $X2=0
+ $Y2=0
cc_515 N_A_110_69#_c_863_n N_A_470_69#_c_949_n 0.00554476f $X=7.285 $Y=1.16
+ $X2=0 $Y2=0
cc_516 N_A_110_69#_c_861_n N_A_470_69#_c_950_n 0.00888527f $X=4.445 $Y=0.71
+ $X2=0 $Y2=0
cc_517 N_A_110_69#_c_863_n N_A_470_69#_c_951_n 0.0364744f $X=7.285 $Y=1.16 $X2=0
+ $Y2=0
cc_518 N_A_110_69#_c_861_n N_A_470_69#_c_952_n 0.00539716f $X=4.445 $Y=0.71
+ $X2=0 $Y2=0
cc_519 N_A_110_69#_c_862_n N_A_470_69#_c_952_n 0.00888527f $X=4.53 $Y=1.075
+ $X2=0 $Y2=0
cc_520 N_A_110_69#_c_863_n N_A_470_69#_c_952_n 0.0143046f $X=7.285 $Y=1.16 $X2=0
+ $Y2=0
cc_521 N_A_110_69#_c_863_n N_A_470_69#_c_962_n 0.0551461f $X=7.285 $Y=1.16 $X2=0
+ $Y2=0
cc_522 N_A_110_69#_c_863_n N_A_470_69#_c_968_n 0.0214932f $X=7.285 $Y=1.16 $X2=0
+ $Y2=0
cc_523 N_A_110_69#_c_863_n N_VGND_c_1011_n 0.0180835f $X=7.285 $Y=1.16 $X2=0
+ $Y2=0
cc_524 N_A_110_69#_c_865_n N_VGND_c_1012_n 0.0154179f $X=8.145 $Y=1.16 $X2=0
+ $Y2=0
cc_525 N_A_110_69#_c_859_n N_VGND_c_1014_n 0.0616577f $X=1.535 $Y=0.355 $X2=0
+ $Y2=0
cc_526 N_A_110_69#_c_860_n N_VGND_c_1014_n 0.0234016f $X=0.855 $Y=0.355 $X2=0
+ $Y2=0
cc_527 N_A_110_69#_c_861_n N_VGND_c_1014_n 0.00925261f $X=4.445 $Y=0.71 $X2=0
+ $Y2=0
cc_528 N_A_110_69#_c_940_p N_VGND_c_1016_n 0.0124525f $X=7.38 $Y=0.42 $X2=0
+ $Y2=0
cc_529 N_A_110_69#_c_941_p N_VGND_c_1018_n 0.0124525f $X=8.24 $Y=0.42 $X2=0
+ $Y2=0
cc_530 N_A_110_69#_M1006_s N_VGND_c_1022_n 0.00536646f $X=7.24 $Y=0.235 $X2=0
+ $Y2=0
cc_531 N_A_110_69#_M1027_s N_VGND_c_1022_n 0.00536646f $X=8.1 $Y=0.235 $X2=0
+ $Y2=0
cc_532 N_A_110_69#_c_859_n N_VGND_c_1022_n 0.0343288f $X=1.535 $Y=0.355 $X2=0
+ $Y2=0
cc_533 N_A_110_69#_c_860_n N_VGND_c_1022_n 0.0125857f $X=0.855 $Y=0.355 $X2=0
+ $Y2=0
cc_534 N_A_110_69#_c_861_n N_VGND_c_1022_n 0.0200897f $X=4.445 $Y=0.71 $X2=0
+ $Y2=0
cc_535 N_A_110_69#_c_940_p N_VGND_c_1022_n 0.00730901f $X=7.38 $Y=0.42 $X2=0
+ $Y2=0
cc_536 N_A_110_69#_c_941_p N_VGND_c_1022_n 0.00730901f $X=8.24 $Y=0.42 $X2=0
+ $Y2=0
cc_537 N_A_470_69#_c_951_n N_VGND_M1010_d 0.00542469f $X=5.495 $Y=0.82 $X2=-0.19
+ $Y2=-0.245
cc_538 N_A_470_69#_c_962_n N_VGND_M1012_d 0.00335437f $X=6.355 $Y=0.82 $X2=0
+ $Y2=0
cc_539 N_A_470_69#_c_949_n N_VGND_c_1008_n 0.0167481f $X=4.795 $Y=0.355 $X2=0
+ $Y2=0
cc_540 N_A_470_69#_c_950_n N_VGND_c_1008_n 0.00816573f $X=4.88 $Y=0.735 $X2=0
+ $Y2=0
cc_541 N_A_470_69#_c_951_n N_VGND_c_1008_n 0.0138809f $X=5.495 $Y=0.82 $X2=0
+ $Y2=0
cc_542 N_A_470_69#_c_951_n N_VGND_c_1009_n 0.00196209f $X=5.495 $Y=0.82 $X2=0
+ $Y2=0
cc_543 N_A_470_69#_c_959_n N_VGND_c_1009_n 0.0118985f $X=5.66 $Y=0.45 $X2=0
+ $Y2=0
cc_544 N_A_470_69#_c_962_n N_VGND_c_1009_n 0.00196209f $X=6.355 $Y=0.82 $X2=0
+ $Y2=0
cc_545 N_A_470_69#_c_962_n N_VGND_c_1010_n 0.0130182f $X=6.355 $Y=0.82 $X2=0
+ $Y2=0
cc_546 N_A_470_69#_c_949_n N_VGND_c_1014_n 0.165859f $X=4.795 $Y=0.355 $X2=0
+ $Y2=0
cc_547 N_A_470_69#_c_951_n N_VGND_c_1014_n 0.0024983f $X=5.495 $Y=0.82 $X2=0
+ $Y2=0
cc_548 N_A_470_69#_c_962_n N_VGND_c_1020_n 0.00196209f $X=6.355 $Y=0.82 $X2=0
+ $Y2=0
cc_549 N_A_470_69#_c_965_n N_VGND_c_1020_n 0.0188748f $X=6.52 $Y=0.42 $X2=0
+ $Y2=0
cc_550 N_A_470_69#_M1002_s N_VGND_c_1022_n 0.00235918f $X=2.35 $Y=0.345 $X2=0
+ $Y2=0
cc_551 N_A_470_69#_M1019_s N_VGND_c_1022_n 0.00235918f $X=3.37 $Y=0.345 $X2=0
+ $Y2=0
cc_552 N_A_470_69#_M1010_s N_VGND_c_1022_n 0.00233619f $X=5.52 $Y=0.235 $X2=0
+ $Y2=0
cc_553 N_A_470_69#_M1031_s N_VGND_c_1022_n 0.00223559f $X=6.38 $Y=0.235 $X2=0
+ $Y2=0
cc_554 N_A_470_69#_c_949_n N_VGND_c_1022_n 0.0947194f $X=4.795 $Y=0.355 $X2=0
+ $Y2=0
cc_555 N_A_470_69#_c_951_n N_VGND_c_1022_n 0.00906049f $X=5.495 $Y=0.82 $X2=0
+ $Y2=0
cc_556 N_A_470_69#_c_959_n N_VGND_c_1022_n 0.011818f $X=5.66 $Y=0.45 $X2=0 $Y2=0
cc_557 N_A_470_69#_c_962_n N_VGND_c_1022_n 0.00835756f $X=6.355 $Y=0.82 $X2=0
+ $Y2=0
cc_558 N_A_470_69#_c_965_n N_VGND_c_1022_n 0.012371f $X=6.52 $Y=0.42 $X2=0 $Y2=0
