* File: sky130_fd_sc_lp__a22oi_4.spice
* Created: Fri Aug 28 09:55:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22oi_4.pex.spice"
.subckt sky130_fd_sc_lp__a22oi_4  VNB VPB B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1009 N_A_63_65#_M1009_d N_B2_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1010 N_A_63_65#_M1010_d N_B2_M1010_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1018 N_A_63_65#_M1010_d N_B2_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1028 N_A_63_65#_M1028_d N_B2_M1028_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1428 AS=0.1176 PD=1.18 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5 SB=75002
+ A=0.126 P=1.98 MULT=1
MM1001 N_A_63_65#_M1028_d N_B1_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1428 AS=0.1176 PD=1.18 PS=1.12 NRD=8.568 NRS=0 M=1 R=5.6 SA=75002
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1011 N_A_63_65#_M1011_d N_B1_M1011_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1020 N_A_63_65#_M1011_d N_B1_M1020_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1024 N_A_63_65#_M1024_d N_B1_M1024_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_867_47#_M1004_d N_A1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_867_47#_M1005_d N_A1_M1005_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1021 N_A_867_47#_M1005_d N_A1_M1021_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1022 N_A_867_47#_M1022_d N_A1_M1022_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_867_47#_M1022_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1002_d N_A2_M1012_g N_A_867_47#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1014_d N_A2_M1014_g N_A_867_47#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1031 N_VGND_M1014_d N_A2_M1031_g N_A_867_47#_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_Y_M1006_d N_B2_M1006_g N_A_89_367#_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75006.9 A=0.189 P=2.82 MULT=1
MM1015 N_Y_M1006_d N_B2_M1015_g N_A_89_367#_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75006.4 A=0.189 P=2.82 MULT=1
MM1023 N_Y_M1023_d N_B2_M1023_g N_A_89_367#_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1 SB=75006
+ A=0.189 P=2.82 MULT=1
MM1027 N_Y_M1023_d N_B2_M1027_g N_A_89_367#_M1027_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75005.6 A=0.189 P=2.82 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_A_89_367#_M1027_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75005.1 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1000_d N_B1_M1008_g N_A_89_367#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2268 PD=1.54 PS=1.62 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75002.3
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1016 N_Y_M1016_d N_B1_M1016_g N_A_89_367#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2268 PD=1.54 PS=1.62 NRD=0 NRS=4.6886 M=1 R=8.4 SA=75002.8
+ SB=75004.2 A=0.189 P=2.82 MULT=1
MM1019 N_Y_M1016_d N_B1_M1019_g N_A_89_367#_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.24255 PD=1.54 PS=1.645 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75003.3
+ SB=75003.8 A=0.189 P=2.82 MULT=1
MM1013 N_A_89_367#_M1019_s N_A1_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.24255 AS=0.1764 PD=1.645 PS=1.54 NRD=8.5892 NRS=0 M=1 R=8.4 SA=75003.8
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1017 N_A_89_367#_M1017_d N_A1_M1017_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1026 N_A_89_367#_M1017_d N_A1_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.20475 PD=1.54 PS=1.585 NRD=0 NRS=0 M=1 R=8.4 SA=75004.7
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1030 N_A_89_367#_M1030_d N_A1_M1030_g N_VPWR_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.20475 PD=1.54 PS=1.585 NRD=0 NRS=7.0329 M=1 R=8.4 SA=75005.1
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_89_367#_M1030_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1003_d N_A2_M1007_g N_A_89_367#_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006 SB=75001.1
+ A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1025_d N_A2_M1025_g N_A_89_367#_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1029 N_VPWR_M1025_d N_A2_M1029_g N_A_89_367#_M1029_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75006.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.9271 P=20.81
*
.include "sky130_fd_sc_lp__a22oi_4.pxi.spice"
*
.ends
*
*
