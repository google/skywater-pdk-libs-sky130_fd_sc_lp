* NGSPICE file created from sky130_fd_sc_lp__dlygate4s18_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlygate4s18_1 A VGND VNB VPB VPWR X
M1000 a_288_52# a_27_52# VGND VNB nshort w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=6.867e+11p ps=5.26e+06u
M1001 X a_405_136# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1002 X a_405_136# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=7.98e+11p ps=6.1e+06u
M1003 VPWR A a_27_52# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 a_288_52# a_27_52# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 VGND A a_27_52# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 VGND a_288_52# a_405_136# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 VPWR a_288_52# a_405_136# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

