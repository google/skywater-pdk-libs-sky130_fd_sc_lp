* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux4_lp A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_114_47# a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_320_366# S1 a_684_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_470_57# S0 a_1692_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 X a_84_21# a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1600_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND S0 a_1860_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND A3 a_915_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_245_411# a_946_317# a_1112_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_245_411# a_320_366# a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_1414_47# S0 a_470_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_245_411# S0 a_1210_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_1210_419# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_915_101# S0 a_245_411# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_470_57# a_946_317# a_1600_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VPWR A1 a_1433_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 VPWR S0 a_946_317# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_1433_419# a_946_317# a_470_57# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X18 a_245_411# S1 a_84_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND A1 a_1414_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_84_21# a_320_366# a_470_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_84_21# S1 a_470_57# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_684_101# S1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_1860_47# S0 a_946_317# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR A3 a_898_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 a_320_366# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X26 a_1112_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_898_419# a_946_317# a_245_411# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X28 a_1692_419# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
