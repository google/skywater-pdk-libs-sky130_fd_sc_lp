* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
X0 VPWR C_N a_206_51# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_1139_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR A a_1139_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND a_37_51# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 Y a_206_51# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_37_51# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND a_206_51# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 Y a_37_51# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_347_349# a_206_51# a_774_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_347_349# a_37_51# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_774_349# B a_1139_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_1139_367# B a_774_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_347_349# a_206_51# a_774_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_774_349# a_206_51# a_347_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_774_349# a_206_51# a_347_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VGND C_N a_206_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_1139_367# B a_774_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND a_37_51# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 Y a_37_51# a_347_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 Y a_206_51# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_774_349# B a_1139_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VPWR A a_1139_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 a_1139_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 Y a_37_51# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 VGND a_206_51# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 a_37_51# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 a_347_349# a_37_51# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 Y a_37_51# a_347_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
