* File: sky130_fd_sc_lp__decapkapwr_12.pxi.spice
* Created: Fri Aug 28 10:20:20 2020
* 
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_12%VGND N_VGND_M1000_s N_VGND_c_27_n
+ N_VGND_M1001_g N_VGND_c_28_n N_VGND_c_29_n N_VGND_c_30_n N_VGND_c_31_n VGND
+ N_VGND_c_32_n N_VGND_c_33_n N_VGND_c_34_n N_VGND_c_35_n N_VGND_c_36_n
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_12%VGND
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_12%KAPWR N_KAPWR_M1001_s N_KAPWR_c_63_n
+ N_KAPWR_c_64_n N_KAPWR_c_73_n N_KAPWR_c_60_n N_KAPWR_c_61_n N_KAPWR_c_67_n
+ N_KAPWR_c_68_n KAPWR N_KAPWR_M1000_g N_KAPWR_c_69_n
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_12%KAPWR
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_12%VPWR VPWR N_VPWR_c_99_n VPWR
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_12%VPWR
cc_1 VNB N_VGND_c_27_n 0.0434284f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=2.555
cc_2 VNB N_VGND_c_28_n 0.0651019f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=0.38
cc_3 VNB N_VGND_c_29_n 0.00211035f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.77
cc_4 VNB N_VGND_c_30_n 4.23625e-19 $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.77
cc_5 VNB N_VGND_c_31_n 0.0371702f $X=-0.19 $Y=-0.245 $X2=5.095 $Y2=0.36
cc_6 VNB N_VGND_c_32_n 0.12354f $X=-0.19 $Y=-0.245 $X2=4.93 $Y2=0
cc_7 VNB N_VGND_c_33_n 0.0180543f $X=-0.19 $Y=-0.245 $X2=5.52 $Y2=0
cc_8 VNB N_VGND_c_34_n 0.327077f $X=-0.19 $Y=-0.245 $X2=5.52 $Y2=0
cc_9 VNB N_VGND_c_35_n 0.0279619f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_10 VNB N_VGND_c_36_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=5.04 $Y2=0
cc_11 VNB N_KAPWR_c_60_n 0.0262142f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=0.38
cc_12 VNB N_KAPWR_c_61_n 0.213478f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.77
cc_13 VNB N_KAPWR_M1000_g 0.167743f $X=-0.19 $Y=-0.245 $X2=5.095 $Y2=1.04
cc_14 VNB VPWR 0.243291f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.235
cc_15 VPB N_VGND_c_27_n 0.403619f $X=-0.19 $Y=1.655 $X2=2.58 $Y2=2.555
cc_16 VPB N_VGND_c_29_n 0.0140672f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.77
cc_17 VPB N_VGND_c_30_n 0.00875776f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=1.77
cc_18 VPB N_KAPWR_c_63_n 0.00922717f $X=-0.19 $Y=1.655 $X2=2.89 $Y2=2.595
cc_19 VPB N_KAPWR_c_64_n 0.023615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_20 VPB N_KAPWR_c_60_n 0.0010232f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=0.38
cc_21 VPB N_KAPWR_c_61_n 0.0404704f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=1.77
cc_22 VPB N_KAPWR_c_67_n 0.00878569f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=1.77
cc_23 VPB N_KAPWR_c_68_n 0.0468814f $X=-0.19 $Y=1.655 $X2=5.095 $Y2=0.085
cc_24 VPB N_KAPWR_c_69_n 0.0691955f $X=-0.19 $Y=1.655 $X2=4.56 $Y2=0
cc_25 VPB VPWR 0.0517013f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.235
cc_26 VPB N_VPWR_c_99_n 0.153085f $X=-0.19 $Y=1.655 $X2=2.89 $Y2=2.555
cc_27 N_VGND_c_27_n N_KAPWR_c_63_n 0.00685959f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_28 N_VGND_c_27_n N_KAPWR_c_64_n 0.0280564f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_29 N_VGND_c_29_n N_KAPWR_c_64_n 0.0205458f $X=0.98 $Y=1.77 $X2=0 $Y2=0
cc_30 N_VGND_c_27_n N_KAPWR_c_73_n 0.237984f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_31 N_VGND_c_27_n N_KAPWR_c_60_n 0.0149963f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_32 N_VGND_c_30_n N_KAPWR_c_60_n 0.00324791f $X=2.415 $Y=1.77 $X2=0 $Y2=0
cc_33 N_VGND_c_31_n N_KAPWR_c_60_n 0.0180876f $X=5.095 $Y=0.36 $X2=0 $Y2=0
cc_34 N_VGND_c_27_n N_KAPWR_c_61_n 0.151712f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_35 N_VGND_c_31_n N_KAPWR_c_61_n 0.0510144f $X=5.095 $Y=0.36 $X2=0 $Y2=0
cc_36 N_VGND_c_34_n N_KAPWR_c_61_n 0.123649f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_37 N_VGND_c_27_n N_KAPWR_c_67_n 0.00731334f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_38 N_VGND_c_27_n N_KAPWR_c_68_n 0.0438461f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_39 N_VGND_c_27_n N_KAPWR_M1000_g 0.119822f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_40 N_VGND_c_28_n N_KAPWR_M1000_g 0.0654854f $X=0.815 $Y=0.38 $X2=0 $Y2=0
cc_41 N_VGND_c_30_n N_KAPWR_M1000_g 0.0121106f $X=2.415 $Y=1.77 $X2=0 $Y2=0
cc_42 N_VGND_c_32_n N_KAPWR_M1000_g 0.154094f $X=4.93 $Y=0 $X2=0 $Y2=0
cc_43 N_VGND_c_34_n N_KAPWR_M1000_g 0.11988f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_44 N_VGND_c_27_n N_KAPWR_c_69_n 0.196513f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_45 N_VGND_c_27_n VPWR 0.0885427f $X=2.58 $Y=2.555 $X2=-0.19 $Y2=-0.245
cc_46 N_VGND_c_27_n N_VPWR_c_99_n 0.103539f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_47 N_KAPWR_M1001_s VPWR 0.00234386f $X=0.615 $Y=2.095 $X2=-0.19 $Y2=-0.245
cc_48 N_KAPWR_c_63_n VPWR 0.00306712f $X=0.74 $Y=2.675 $X2=-0.19 $Y2=-0.245
cc_49 N_KAPWR_c_73_n VPWR 0.0220134f $X=4.865 $Y=2.81 $X2=-0.19 $Y2=-0.245
cc_50 N_KAPWR_c_67_n VPWR 0.00305163f $X=5.03 $Y=2.675 $X2=-0.19 $Y2=-0.245
cc_51 N_KAPWR_c_69_n VPWR 0.600777f $X=5.015 $Y=2.81 $X2=-0.19 $Y2=-0.245
cc_52 N_KAPWR_c_63_n N_VPWR_c_99_n 0.0212079f $X=0.74 $Y=2.675 $X2=0 $Y2=0
cc_53 N_KAPWR_c_73_n N_VPWR_c_99_n 0.143201f $X=4.865 $Y=2.81 $X2=0 $Y2=0
cc_54 N_KAPWR_c_67_n N_VPWR_c_99_n 0.0211263f $X=5.03 $Y=2.675 $X2=0 $Y2=0
cc_55 N_KAPWR_c_69_n N_VPWR_c_99_n 0.0153779f $X=5.015 $Y=2.81 $X2=0 $Y2=0
