* File: sky130_fd_sc_lp__ha_m.pxi.spice
* Created: Wed Sep  2 09:54:51 2020
* 
x_PM_SKY130_FD_SC_LP__HA_M%A_80_60# N_A_80_60#_M1011_s N_A_80_60#_M1003_d
+ N_A_80_60#_M1001_g N_A_80_60#_c_101_n N_A_80_60#_c_102_n N_A_80_60#_c_103_n
+ N_A_80_60#_M1002_g N_A_80_60#_c_97_n N_A_80_60#_c_98_n N_A_80_60#_c_106_n
+ N_A_80_60#_c_107_n N_A_80_60#_c_99_n N_A_80_60#_c_109_n N_A_80_60#_c_110_n
+ N_A_80_60#_c_120_p N_A_80_60#_c_132_p N_A_80_60#_c_100_n N_A_80_60#_c_111_n
+ PM_SKY130_FD_SC_LP__HA_M%A_80_60#
x_PM_SKY130_FD_SC_LP__HA_M%A_249_212# N_A_249_212#_M1005_s N_A_249_212#_M1013_d
+ N_A_249_212#_M1011_g N_A_249_212#_c_189_n N_A_249_212#_M1003_g
+ N_A_249_212#_c_191_n N_A_249_212#_M1010_g N_A_249_212#_M1004_g
+ N_A_249_212#_c_179_n N_A_249_212#_c_180_n N_A_249_212#_c_194_n
+ N_A_249_212#_c_181_n N_A_249_212#_c_182_n N_A_249_212#_c_183_n
+ N_A_249_212#_c_196_n N_A_249_212#_c_184_n N_A_249_212#_c_185_n
+ N_A_249_212#_c_186_n N_A_249_212#_c_187_n N_A_249_212#_c_188_n
+ N_A_249_212#_c_198_n PM_SKY130_FD_SC_LP__HA_M%A_249_212#
x_PM_SKY130_FD_SC_LP__HA_M%B N_B_M1006_g N_B_c_298_n N_B_M1012_g N_B_c_306_n
+ N_B_M1013_g N_B_M1005_g N_B_c_300_n N_B_c_308_n N_B_c_301_n N_B_c_302_n
+ N_B_c_309_n N_B_c_340_n N_B_c_303_n B PM_SKY130_FD_SC_LP__HA_M%B
x_PM_SKY130_FD_SC_LP__HA_M%A N_A_c_378_n N_A_M1007_g N_A_c_379_n N_A_c_380_n
+ N_A_M1009_g N_A_c_382_n N_A_c_383_n N_A_c_384_n N_A_M1000_g N_A_M1008_g A
+ N_A_c_386_n PM_SKY130_FD_SC_LP__HA_M%A
x_PM_SKY130_FD_SC_LP__HA_M%SUM N_SUM_M1001_s N_SUM_M1002_s N_SUM_c_446_n SUM SUM
+ SUM SUM SUM SUM SUM PM_SKY130_FD_SC_LP__HA_M%SUM
x_PM_SKY130_FD_SC_LP__HA_M%VPWR N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_M1008_d
+ N_VPWR_c_471_n N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_475_n
+ N_VPWR_c_476_n N_VPWR_c_477_n VPWR N_VPWR_c_478_n N_VPWR_c_479_n
+ N_VPWR_c_470_n N_VPWR_c_481_n PM_SKY130_FD_SC_LP__HA_M%VPWR
x_PM_SKY130_FD_SC_LP__HA_M%COUT N_COUT_M1010_d N_COUT_M1004_d COUT COUT COUT
+ COUT COUT COUT COUT PM_SKY130_FD_SC_LP__HA_M%COUT
x_PM_SKY130_FD_SC_LP__HA_M%VGND N_VGND_M1001_d N_VGND_M1006_d N_VGND_M1000_d
+ N_VGND_c_542_n N_VGND_c_543_n VGND N_VGND_c_544_n N_VGND_c_545_n
+ N_VGND_c_546_n N_VGND_c_547_n N_VGND_c_548_n N_VGND_c_549_n N_VGND_c_550_n
+ N_VGND_c_551_n PM_SKY130_FD_SC_LP__HA_M%VGND
x_PM_SKY130_FD_SC_LP__HA_M%A_301_47# N_A_301_47#_M1011_d N_A_301_47#_M1007_d
+ N_A_301_47#_c_595_n N_A_301_47#_c_596_n N_A_301_47#_c_597_n
+ PM_SKY130_FD_SC_LP__HA_M%A_301_47#
cc_1 VNB N_A_80_60#_M1001_g 0.0592011f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_2 VNB N_A_80_60#_c_97_n 0.00682989f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.615
cc_3 VNB N_A_80_60#_c_98_n 0.032832f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.615
cc_4 VNB N_A_80_60#_c_99_n 0.0226877f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.95
cc_5 VNB N_A_80_60#_c_100_n 0.0098814f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=0.51
cc_6 VNB N_A_249_212#_M1011_g 0.036639f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_7 VNB N_A_249_212#_M1010_g 0.046205f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.615
cc_8 VNB N_A_249_212#_c_179_n 0.0268083f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.95
cc_9 VNB N_A_249_212#_c_180_n 0.00613729f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=2.035
cc_10 VNB N_A_249_212#_c_181_n 0.00117897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_249_212#_c_182_n 0.0203806f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=0.51
cc_12 VNB N_A_249_212#_c_183_n 0.0168386f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=0.51
cc_13 VNB N_A_249_212#_c_184_n 0.00490232f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=2.035
cc_14 VNB N_A_249_212#_c_185_n 0.00383177f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.45
cc_15 VNB N_A_249_212#_c_186_n 0.00599907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_249_212#_c_187_n 0.0114484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_249_212#_c_188_n 0.00844873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_M1006_g 0.0651268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_c_298_n 0.00769642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_M1005_g 0.0195694f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.045
cc_21 VNB N_B_c_300_n 0.00328608f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=2.53
cc_22 VNB N_B_c_301_n 0.0445222f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.615
cc_23 VNB N_B_c_302_n 0.00860446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_303_n 0.00149679f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.36
cc_25 VNB N_A_c_378_n 0.0171616f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=0.235
cc_26 VNB N_A_c_379_n 0.0267479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_c_380_n 0.0558024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_M1009_g 0.0154485f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_29 VNB N_A_c_382_n 0.0358373f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.677
cc_30 VNB N_A_c_383_n 0.0680944f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.97
cc_31 VNB N_A_c_384_n 0.00989713f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.045
cc_32 VNB N_A_M1000_g 0.057976f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=2.53
cc_33 VNB N_A_c_386_n 0.00495698f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.035
cc_34 VNB SUM 0.0488112f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.677
cc_35 VNB N_VPWR_c_470_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB COUT 0.0422515f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.45
cc_37 VNB N_VGND_c_542_n 0.011586f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.97
cc_38 VNB N_VGND_c_543_n 0.0202292f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=2.53
cc_39 VNB N_VGND_c_544_n 0.0193716f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.615
cc_40 VNB N_VGND_c_545_n 0.0326235f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.035
cc_41 VNB N_VGND_c_546_n 0.0504619f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.12
cc_42 VNB N_VGND_c_547_n 0.0203686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_548_n 0.278917f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=2.035
cc_44 VNB N_VGND_c_549_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_550_n 0.0116582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_551_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_301_47#_c_595_n 0.00986895f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.45
cc_48 VNB N_A_301_47#_c_596_n 0.00836207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_301_47#_c_597_n 0.00150115f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=2.12
cc_50 VPB N_A_80_60#_c_101_n 0.0301299f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.97
cc_51 VPB N_A_80_60#_c_102_n 0.0229948f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.045
cc_52 VPB N_A_80_60#_c_103_n 0.0248633f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.045
cc_53 VPB N_A_80_60#_M1002_g 0.0273905f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=2.53
cc_54 VPB N_A_80_60#_c_98_n 0.00220214f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.615
cc_55 VPB N_A_80_60#_c_106_n 0.00408807f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.035
cc_56 VPB N_A_80_60#_c_107_n 0.00216294f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=2.035
cc_57 VPB N_A_80_60#_c_99_n 0.00487477f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.95
cc_58 VPB N_A_80_60#_c_109_n 0.0121853f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=2.035
cc_59 VPB N_A_80_60#_c_110_n 0.00199972f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.36
cc_60 VPB N_A_80_60#_c_111_n 0.00114618f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=2.035
cc_61 VPB N_A_249_212#_c_189_n 0.0184766f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.97
cc_62 VPB N_A_249_212#_M1003_g 0.0195432f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=2.12
cc_63 VPB N_A_249_212#_c_191_n 0.0443438f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=2.53
cc_64 VPB N_A_249_212#_M1010_g 0.0415069f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.615
cc_65 VPB N_A_249_212#_c_180_n 0.0101021f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=2.035
cc_66 VPB N_A_249_212#_c_194_n 0.0274766f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.36
cc_67 VPB N_A_249_212#_c_183_n 0.00586579f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=0.51
cc_68 VPB N_A_249_212#_c_196_n 0.00101985f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=0.51
cc_69 VPB N_A_249_212#_c_186_n 0.0122782f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_249_212#_c_198_n 0.0461866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_B_c_298_n 0.0534362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_B_M1012_g 0.0206078f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.45
cc_73 VPB N_B_c_306_n 0.0205692f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.64
cc_74 VPB N_B_c_300_n 0.00280318f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=2.53
cc_75 VPB N_B_c_308_n 0.0243112f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.615
cc_76 VPB N_B_c_309_n 0.0207542f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.035
cc_77 VPB N_B_c_303_n 0.0035103f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.36
cc_78 VPB N_A_M1009_g 0.0494948f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.64
cc_79 VPB N_A_M1000_g 0.02983f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=2.53
cc_80 VPB N_SUM_c_446_n 0.0160571f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.64
cc_81 VPB SUM 0.0421237f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.677
cc_82 VPB SUM 0.0230255f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=2.53
cc_83 VPB N_VPWR_c_471_n 0.0252144f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.97
cc_84 VPB N_VPWR_c_472_n 0.0264172f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=2.53
cc_85 VPB N_VPWR_c_473_n 0.0171033f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.615
cc_86 VPB N_VPWR_c_474_n 0.0364187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_475_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.035
cc_88 VPB N_VPWR_c_476_n 0.0400815f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=0.675
cc_89 VPB N_VPWR_c_477_n 0.00632158f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.95
cc_90 VPB N_VPWR_c_478_n 0.0249566f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.45
cc_91 VPB N_VPWR_c_479_n 0.0203686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_470_n 0.116287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_481_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB COUT 0.0425212f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.45
cc_95 N_A_80_60#_c_99_n N_A_249_212#_M1011_g 0.0115024f $X=1.06 $Y=1.95 $X2=0
+ $Y2=0
cc_96 N_A_80_60#_c_100_n N_A_249_212#_M1011_g 4.43596e-19 $X=1.215 $Y=0.51 $X2=0
+ $Y2=0
cc_97 N_A_80_60#_c_101_n N_A_249_212#_c_189_n 0.00326993f $X=0.627 $Y=1.97 $X2=0
+ $Y2=0
cc_98 N_A_80_60#_c_102_n N_A_249_212#_c_189_n 0.00705855f $X=1.065 $Y=2.045
+ $X2=0 $Y2=0
cc_99 N_A_80_60#_c_99_n N_A_249_212#_c_189_n 0.00447058f $X=1.06 $Y=1.95 $X2=0
+ $Y2=0
cc_100 N_A_80_60#_c_109_n N_A_249_212#_c_189_n 0.00556739f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_101 N_A_80_60#_M1002_g N_A_249_212#_M1003_g 0.0112436f $X=1.14 $Y=2.53 $X2=0
+ $Y2=0
cc_102 N_A_80_60#_c_110_n N_A_249_212#_M1003_g 0.00538443f $X=1.765 $Y=2.36
+ $X2=0 $Y2=0
cc_103 N_A_80_60#_c_120_p N_A_249_212#_M1003_g 0.00782229f $X=1.85 $Y=2.465
+ $X2=0 $Y2=0
cc_104 N_A_80_60#_c_98_n N_A_249_212#_c_179_n 0.00348877f $X=0.69 $Y=1.615 $X2=0
+ $Y2=0
cc_105 N_A_80_60#_c_101_n N_A_249_212#_c_180_n 0.00348877f $X=0.627 $Y=1.97
+ $X2=0 $Y2=0
cc_106 N_A_80_60#_c_109_n N_A_249_212#_c_180_n 0.00377636f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_107 N_A_80_60#_M1002_g N_A_249_212#_c_194_n 0.00705855f $X=1.14 $Y=2.53 $X2=0
+ $Y2=0
cc_108 N_A_80_60#_c_109_n N_A_249_212#_c_194_n 0.0156497f $X=1.68 $Y=2.035 $X2=0
+ $Y2=0
cc_109 N_A_80_60#_c_110_n N_A_249_212#_c_194_n 0.0020618f $X=1.765 $Y=2.36 $X2=0
+ $Y2=0
cc_110 N_A_80_60#_c_99_n N_A_249_212#_c_181_n 0.0341905f $X=1.06 $Y=1.95 $X2=0
+ $Y2=0
cc_111 N_A_80_60#_M1001_g N_A_249_212#_c_182_n 0.00386146f $X=0.475 $Y=0.64
+ $X2=0 $Y2=0
cc_112 N_A_80_60#_c_99_n N_A_249_212#_c_182_n 0.00725983f $X=1.06 $Y=1.95 $X2=0
+ $Y2=0
cc_113 N_A_80_60#_c_100_n N_A_249_212#_c_182_n 0.00192551f $X=1.215 $Y=0.51
+ $X2=0 $Y2=0
cc_114 N_A_80_60#_c_109_n N_A_249_212#_c_183_n 0.0225855f $X=1.68 $Y=2.035 $X2=0
+ $Y2=0
cc_115 N_A_80_60#_c_132_p N_A_249_212#_c_183_n 0.00420091f $X=1.96 $Y=2.465
+ $X2=0 $Y2=0
cc_116 N_A_80_60#_c_99_n N_A_249_212#_c_196_n 0.0129659f $X=1.06 $Y=1.95 $X2=0
+ $Y2=0
cc_117 N_A_80_60#_c_109_n N_A_249_212#_c_196_n 0.010897f $X=1.68 $Y=2.035 $X2=0
+ $Y2=0
cc_118 N_A_80_60#_c_109_n N_B_c_298_n 0.00184719f $X=1.68 $Y=2.035 $X2=0 $Y2=0
cc_119 N_A_80_60#_c_110_n N_B_c_298_n 7.89749e-19 $X=1.765 $Y=2.36 $X2=0 $Y2=0
cc_120 N_A_80_60#_c_132_p N_B_c_298_n 0.00453717f $X=1.96 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_80_60#_c_110_n N_B_M1012_g 0.00298567f $X=1.765 $Y=2.36 $X2=0 $Y2=0
cc_122 N_A_80_60#_c_132_p N_B_M1012_g 0.0050279f $X=1.96 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_80_60#_c_109_n N_B_c_309_n 0.0144263f $X=1.68 $Y=2.035 $X2=0 $Y2=0
cc_124 N_A_80_60#_c_132_p N_B_c_309_n 0.00354063f $X=1.96 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_80_60#_c_132_p N_A_M1009_g 8.63719e-19 $X=1.96 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_80_60#_c_102_n N_SUM_c_446_n 3.84218e-19 $X=1.065 $Y=2.045 $X2=0
+ $Y2=0
cc_127 N_A_80_60#_c_103_n N_SUM_c_446_n 0.011498f $X=0.855 $Y=2.045 $X2=0 $Y2=0
cc_128 N_A_80_60#_M1002_g N_SUM_c_446_n 0.00754051f $X=1.14 $Y=2.53 $X2=0 $Y2=0
cc_129 N_A_80_60#_c_106_n N_SUM_c_446_n 0.00822156f $X=0.975 $Y=2.035 $X2=0
+ $Y2=0
cc_130 N_A_80_60#_c_107_n N_SUM_c_446_n 0.00802704f $X=0.775 $Y=2.035 $X2=0
+ $Y2=0
cc_131 N_A_80_60#_c_111_n N_SUM_c_446_n 0.00381747f $X=1.06 $Y=2.035 $X2=0 $Y2=0
cc_132 N_A_80_60#_M1001_g SUM 0.031151f $X=0.475 $Y=0.64 $X2=0 $Y2=0
cc_133 N_A_80_60#_c_101_n SUM 0.0107398f $X=0.627 $Y=1.97 $X2=0 $Y2=0
cc_134 N_A_80_60#_c_103_n SUM 0.00614085f $X=0.855 $Y=2.045 $X2=0 $Y2=0
cc_135 N_A_80_60#_M1002_g SUM 0.00748519f $X=1.14 $Y=2.53 $X2=0 $Y2=0
cc_136 N_A_80_60#_c_97_n SUM 0.034006f $X=0.69 $Y=1.615 $X2=0 $Y2=0
cc_137 N_A_80_60#_c_98_n SUM 0.00838967f $X=0.69 $Y=1.615 $X2=0 $Y2=0
cc_138 N_A_80_60#_c_107_n SUM 0.0128825f $X=0.775 $Y=2.035 $X2=0 $Y2=0
cc_139 N_A_80_60#_c_99_n SUM 0.0219618f $X=1.06 $Y=1.95 $X2=0 $Y2=0
cc_140 N_A_80_60#_M1002_g N_VPWR_c_471_n 0.00141408f $X=1.14 $Y=2.53 $X2=0 $Y2=0
cc_141 N_A_80_60#_c_109_n N_VPWR_c_471_n 0.0109284f $X=1.68 $Y=2.035 $X2=0 $Y2=0
cc_142 N_A_80_60#_c_120_p N_VPWR_c_471_n 0.00952264f $X=1.85 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_80_60#_c_132_p N_VPWR_c_472_n 0.00211665f $X=1.96 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_80_60#_M1002_g N_VPWR_c_474_n 0.00415805f $X=1.14 $Y=2.53 $X2=0 $Y2=0
cc_145 N_A_80_60#_c_120_p N_VPWR_c_476_n 0.00210502f $X=1.85 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_80_60#_c_132_p N_VPWR_c_476_n 0.00317676f $X=1.96 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_80_60#_M1002_g N_VPWR_c_470_n 0.00479212f $X=1.14 $Y=2.53 $X2=0 $Y2=0
cc_148 N_A_80_60#_c_120_p N_VPWR_c_470_n 0.00447421f $X=1.85 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_80_60#_c_132_p N_VPWR_c_470_n 0.00715072f $X=1.96 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_80_60#_M1001_g N_VGND_c_542_n 0.00509177f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_151 N_A_80_60#_c_99_n N_VGND_c_542_n 0.00465097f $X=1.06 $Y=1.95 $X2=0 $Y2=0
cc_152 N_A_80_60#_c_100_n N_VGND_c_542_n 0.0249227f $X=1.215 $Y=0.51 $X2=0 $Y2=0
cc_153 N_A_80_60#_M1001_g N_VGND_c_544_n 0.00511809f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_154 N_A_80_60#_c_100_n N_VGND_c_545_n 0.0137343f $X=1.215 $Y=0.51 $X2=0 $Y2=0
cc_155 N_A_80_60#_M1011_s N_VGND_c_548_n 0.00413758f $X=1.09 $Y=0.235 $X2=0
+ $Y2=0
cc_156 N_A_80_60#_M1001_g N_VGND_c_548_n 0.00526787f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_157 N_A_80_60#_c_100_n N_VGND_c_548_n 0.0117432f $X=1.215 $Y=0.51 $X2=0 $Y2=0
cc_158 N_A_80_60#_c_99_n N_A_301_47#_c_596_n 0.00382969f $X=1.06 $Y=1.95 $X2=0
+ $Y2=0
cc_159 N_A_80_60#_c_100_n N_A_301_47#_c_596_n 0.00114009f $X=1.215 $Y=0.51 $X2=0
+ $Y2=0
cc_160 N_A_249_212#_M1011_g N_B_M1006_g 0.0286724f $X=1.43 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_249_212#_c_181_n N_B_M1006_g 0.00203421f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_162 N_A_249_212#_c_182_n N_B_M1006_g 0.0233717f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_163 N_A_249_212#_c_183_n N_B_M1006_g 0.0101958f $X=2.61 $Y=1.645 $X2=0 $Y2=0
cc_164 N_A_249_212#_c_184_n N_B_M1006_g 8.05945e-19 $X=2.695 $Y=1.56 $X2=0 $Y2=0
cc_165 N_A_249_212#_c_185_n N_B_M1006_g 0.00108249f $X=2.78 $Y=1.03 $X2=0 $Y2=0
cc_166 N_A_249_212#_c_189_n N_B_c_298_n 0.00672917f $X=1.5 $Y=2.035 $X2=0 $Y2=0
cc_167 N_A_249_212#_c_180_n N_B_c_298_n 0.0233717f $X=1.41 $Y=1.73 $X2=0 $Y2=0
cc_168 N_A_249_212#_c_194_n N_B_c_298_n 0.00999437f $X=1.745 $Y=2.11 $X2=0 $Y2=0
cc_169 N_A_249_212#_c_183_n N_B_c_298_n 0.0166438f $X=2.61 $Y=1.645 $X2=0 $Y2=0
cc_170 N_A_249_212#_c_194_n N_B_M1012_g 0.0165305f $X=1.745 $Y=2.11 $X2=0 $Y2=0
cc_171 N_A_249_212#_c_186_n N_B_c_306_n 0.0125387f $X=3.575 $Y=2.29 $X2=0 $Y2=0
cc_172 N_A_249_212#_c_184_n N_B_M1005_g 0.00202473f $X=2.695 $Y=1.56 $X2=0 $Y2=0
cc_173 N_A_249_212#_c_186_n N_B_M1005_g 0.00660054f $X=3.575 $Y=2.29 $X2=0 $Y2=0
cc_174 N_A_249_212#_c_188_n N_B_M1005_g 0.0160324f $X=3.635 $Y=0.955 $X2=0 $Y2=0
cc_175 N_A_249_212#_c_186_n N_B_c_300_n 0.00668744f $X=3.575 $Y=2.29 $X2=0 $Y2=0
cc_176 N_A_249_212#_c_186_n N_B_c_308_n 0.00825612f $X=3.575 $Y=2.29 $X2=0 $Y2=0
cc_177 N_A_249_212#_c_184_n N_B_c_301_n 0.0040207f $X=2.695 $Y=1.56 $X2=0 $Y2=0
cc_178 N_A_249_212#_c_187_n N_B_c_301_n 0.0142101f $X=3.05 $Y=0.955 $X2=0 $Y2=0
cc_179 N_A_249_212#_c_186_n N_B_c_302_n 0.0134734f $X=3.575 $Y=2.29 $X2=0 $Y2=0
cc_180 N_A_249_212#_c_189_n N_B_c_309_n 2.89893e-19 $X=1.5 $Y=2.035 $X2=0 $Y2=0
cc_181 N_A_249_212#_c_183_n N_B_c_309_n 0.05345f $X=2.61 $Y=1.645 $X2=0 $Y2=0
cc_182 N_A_249_212#_c_186_n N_B_c_340_n 0.0167127f $X=3.575 $Y=2.29 $X2=0 $Y2=0
cc_183 N_A_249_212#_c_183_n N_B_c_303_n 0.014439f $X=2.61 $Y=1.645 $X2=0 $Y2=0
cc_184 N_A_249_212#_c_184_n N_B_c_303_n 0.0191031f $X=2.695 $Y=1.56 $X2=0 $Y2=0
cc_185 N_A_249_212#_c_186_n N_B_c_303_n 0.0448328f $X=3.575 $Y=2.29 $X2=0 $Y2=0
cc_186 N_A_249_212#_c_187_n N_B_c_303_n 0.0259311f $X=3.05 $Y=0.955 $X2=0 $Y2=0
cc_187 N_A_249_212#_c_185_n N_A_c_379_n 0.00280351f $X=2.78 $Y=1.03 $X2=0 $Y2=0
cc_188 N_A_249_212#_c_187_n N_A_c_379_n 0.0101396f $X=3.05 $Y=0.955 $X2=0 $Y2=0
cc_189 N_A_249_212#_c_188_n N_A_c_379_n 0.00439539f $X=3.635 $Y=0.955 $X2=0
+ $Y2=0
cc_190 N_A_249_212#_c_183_n N_A_c_380_n 0.00891601f $X=2.61 $Y=1.645 $X2=0 $Y2=0
cc_191 N_A_249_212#_c_184_n N_A_c_380_n 0.00689847f $X=2.695 $Y=1.56 $X2=0 $Y2=0
cc_192 N_A_249_212#_c_185_n N_A_c_380_n 0.00375731f $X=2.78 $Y=1.03 $X2=0 $Y2=0
cc_193 N_A_249_212#_c_183_n N_A_M1009_g 0.0108295f $X=2.61 $Y=1.645 $X2=0 $Y2=0
cc_194 N_A_249_212#_c_184_n N_A_M1009_g 0.00509516f $X=2.695 $Y=1.56 $X2=0 $Y2=0
cc_195 N_A_249_212#_c_188_n N_A_c_383_n 0.0106646f $X=3.635 $Y=0.955 $X2=0 $Y2=0
cc_196 N_A_249_212#_c_191_n N_A_M1000_g 0.00948934f $X=4.24 $Y=2.88 $X2=0 $Y2=0
cc_197 N_A_249_212#_M1010_g N_A_M1000_g 0.0557734f $X=4.315 $Y=0.835 $X2=0 $Y2=0
cc_198 N_A_249_212#_c_186_n N_A_M1000_g 0.0176378f $X=3.575 $Y=2.29 $X2=0 $Y2=0
cc_199 N_A_249_212#_c_188_n N_A_M1000_g 0.00200793f $X=3.635 $Y=0.955 $X2=0
+ $Y2=0
cc_200 N_A_249_212#_c_181_n N_A_c_386_n 0.0095845f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_201 N_A_249_212#_c_183_n N_A_c_386_n 0.0259917f $X=2.61 $Y=1.645 $X2=0 $Y2=0
cc_202 N_A_249_212#_c_184_n N_A_c_386_n 0.0186968f $X=2.695 $Y=1.56 $X2=0 $Y2=0
cc_203 N_A_249_212#_c_185_n N_A_c_386_n 0.00521892f $X=2.78 $Y=1.03 $X2=0 $Y2=0
cc_204 N_A_249_212#_M1003_g N_VPWR_c_471_n 0.00785705f $X=1.745 $Y=2.53 $X2=0
+ $Y2=0
cc_205 N_A_249_212#_c_194_n N_VPWR_c_471_n 0.00145115f $X=1.745 $Y=2.11 $X2=0
+ $Y2=0
cc_206 N_A_249_212#_c_186_n N_VPWR_c_472_n 0.0259578f $X=3.575 $Y=2.29 $X2=0
+ $Y2=0
cc_207 N_A_249_212#_c_198_n N_VPWR_c_472_n 0.0079729f $X=3.8 $Y=2.94 $X2=0 $Y2=0
cc_208 N_A_249_212#_c_191_n N_VPWR_c_473_n 0.017918f $X=4.24 $Y=2.88 $X2=0 $Y2=0
cc_209 N_A_249_212#_M1010_g N_VPWR_c_473_n 0.00618526f $X=4.315 $Y=0.835 $X2=0
+ $Y2=0
cc_210 N_A_249_212#_c_186_n N_VPWR_c_473_n 0.041109f $X=3.575 $Y=2.29 $X2=0
+ $Y2=0
cc_211 N_A_249_212#_c_198_n N_VPWR_c_473_n 0.00455944f $X=3.8 $Y=2.94 $X2=0
+ $Y2=0
cc_212 N_A_249_212#_M1003_g N_VPWR_c_476_n 0.00348772f $X=1.745 $Y=2.53 $X2=0
+ $Y2=0
cc_213 N_A_249_212#_c_191_n N_VPWR_c_478_n 0.00502584f $X=4.24 $Y=2.88 $X2=0
+ $Y2=0
cc_214 N_A_249_212#_c_186_n N_VPWR_c_478_n 0.0167839f $X=3.575 $Y=2.29 $X2=0
+ $Y2=0
cc_215 N_A_249_212#_c_198_n N_VPWR_c_478_n 0.0059602f $X=3.8 $Y=2.94 $X2=0 $Y2=0
cc_216 N_A_249_212#_c_191_n N_VPWR_c_479_n 0.00624401f $X=4.24 $Y=2.88 $X2=0
+ $Y2=0
cc_217 N_A_249_212#_M1003_g N_VPWR_c_470_n 0.00479212f $X=1.745 $Y=2.53 $X2=0
+ $Y2=0
cc_218 N_A_249_212#_c_191_n N_VPWR_c_470_n 0.0117606f $X=4.24 $Y=2.88 $X2=0
+ $Y2=0
cc_219 N_A_249_212#_c_186_n N_VPWR_c_470_n 0.0108843f $X=3.575 $Y=2.29 $X2=0
+ $Y2=0
cc_220 N_A_249_212#_c_198_n N_VPWR_c_470_n 0.00813556f $X=3.8 $Y=2.94 $X2=0
+ $Y2=0
cc_221 N_A_249_212#_M1010_g COUT 0.0447188f $X=4.315 $Y=0.835 $X2=0 $Y2=0
cc_222 N_A_249_212#_c_186_n COUT 0.0287885f $X=3.575 $Y=2.29 $X2=0 $Y2=0
cc_223 N_A_249_212#_c_188_n COUT 0.00231043f $X=3.635 $Y=0.955 $X2=0 $Y2=0
cc_224 N_A_249_212#_M1011_g N_VGND_c_542_n 0.00438568f $X=1.43 $Y=0.445 $X2=0
+ $Y2=0
cc_225 N_A_249_212#_M1010_g N_VGND_c_543_n 0.00104922f $X=4.315 $Y=0.835 $X2=0
+ $Y2=0
cc_226 N_A_249_212#_M1011_g N_VGND_c_545_n 0.00585385f $X=1.43 $Y=0.445 $X2=0
+ $Y2=0
cc_227 N_A_249_212#_M1010_g N_VGND_c_547_n 0.00415323f $X=4.315 $Y=0.835 $X2=0
+ $Y2=0
cc_228 N_A_249_212#_M1011_g N_VGND_c_548_n 0.0124078f $X=1.43 $Y=0.445 $X2=0
+ $Y2=0
cc_229 N_A_249_212#_M1010_g N_VGND_c_548_n 0.00469432f $X=4.315 $Y=0.835 $X2=0
+ $Y2=0
cc_230 N_A_249_212#_c_188_n N_VGND_c_548_n 0.025146f $X=3.635 $Y=0.955 $X2=0
+ $Y2=0
cc_231 N_A_249_212#_M1011_g N_A_301_47#_c_596_n 0.00115186f $X=1.43 $Y=0.445
+ $X2=0 $Y2=0
cc_232 N_A_249_212#_c_182_n N_A_301_47#_c_596_n 0.00135605f $X=1.41 $Y=1.225
+ $X2=0 $Y2=0
cc_233 N_A_249_212#_c_185_n N_A_301_47#_c_597_n 0.0131159f $X=2.78 $Y=1.03 $X2=0
+ $Y2=0
cc_234 N_A_249_212#_c_188_n A_720_125# 0.00123774f $X=3.635 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_235 N_B_M1006_g N_A_c_378_n 0.0258072f $X=1.86 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_236 N_B_c_301_n N_A_c_379_n 0.00208957f $X=3.45 $Y=1.38 $X2=0 $Y2=0
cc_237 N_B_M1006_g N_A_c_380_n 0.0174568f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_238 N_B_c_298_n N_A_c_380_n 0.00398663f $X=2.175 $Y=2.16 $X2=0 $Y2=0
cc_239 N_B_c_301_n N_A_c_380_n 0.0160409f $X=3.45 $Y=1.38 $X2=0 $Y2=0
cc_240 N_B_c_303_n N_A_c_380_n 2.83371e-19 $X=3.125 $Y=1.38 $X2=0 $Y2=0
cc_241 N_B_M1006_g N_A_M1009_g 0.0039992f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_242 N_B_c_298_n N_A_M1009_g 0.0282093f $X=2.175 $Y=2.16 $X2=0 $Y2=0
cc_243 N_B_M1012_g N_A_M1009_g 0.0291686f $X=2.175 $Y=2.53 $X2=0 $Y2=0
cc_244 N_B_c_308_n N_A_M1009_g 0.0204443f $X=3.525 $Y=1.83 $X2=0 $Y2=0
cc_245 N_B_c_309_n N_A_M1009_g 0.017241f $X=2.96 $Y=2.015 $X2=0 $Y2=0
cc_246 N_B_c_303_n N_A_M1009_g 0.00564383f $X=3.125 $Y=1.38 $X2=0 $Y2=0
cc_247 N_B_M1005_g N_A_c_382_n 0.0119958f $X=3.525 $Y=0.835 $X2=0 $Y2=0
cc_248 N_B_M1005_g N_A_c_383_n 0.00857118f $X=3.525 $Y=0.835 $X2=0 $Y2=0
cc_249 N_B_c_306_n N_A_M1000_g 0.0105699f $X=3.265 $Y=1.905 $X2=0 $Y2=0
cc_250 N_B_M1005_g N_A_M1000_g 0.0832681f $X=3.525 $Y=0.835 $X2=0 $Y2=0
cc_251 N_B_M1006_g N_A_c_386_n 0.00377373f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_252 N_B_c_298_n N_A_c_386_n 6.16164e-19 $X=2.175 $Y=2.16 $X2=0 $Y2=0
cc_253 N_B_c_309_n N_VPWR_M1009_d 0.00233754f $X=2.96 $Y=2.015 $X2=0 $Y2=0
cc_254 N_B_c_340_n N_VPWR_M1009_d 0.00347798f $X=3.125 $Y=1.91 $X2=0 $Y2=0
cc_255 N_B_c_306_n N_VPWR_c_472_n 9.2134e-19 $X=3.265 $Y=1.905 $X2=0 $Y2=0
cc_256 N_B_c_309_n N_VPWR_c_472_n 0.00789408f $X=2.96 $Y=2.015 $X2=0 $Y2=0
cc_257 N_B_c_340_n N_VPWR_c_472_n 0.00812836f $X=3.125 $Y=1.91 $X2=0 $Y2=0
cc_258 N_B_M1012_g N_VPWR_c_476_n 0.00418997f $X=2.175 $Y=2.53 $X2=0 $Y2=0
cc_259 N_B_c_306_n N_VPWR_c_478_n 0.00297774f $X=3.265 $Y=1.905 $X2=0 $Y2=0
cc_260 N_B_M1012_g N_VPWR_c_470_n 0.00479212f $X=2.175 $Y=2.53 $X2=0 $Y2=0
cc_261 N_B_c_306_n N_VPWR_c_470_n 0.00400849f $X=3.265 $Y=1.905 $X2=0 $Y2=0
cc_262 N_B_M1006_g N_VGND_c_545_n 0.00419075f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_263 N_B_M1006_g N_VGND_c_548_n 0.006227f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_264 N_B_M1005_g N_VGND_c_548_n 9.49986e-19 $X=3.525 $Y=0.835 $X2=0 $Y2=0
cc_265 N_B_M1006_g N_VGND_c_550_n 0.00423616f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_266 N_B_M1006_g N_A_301_47#_c_595_n 0.0153982f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_267 N_B_M1006_g N_A_301_47#_c_596_n 2.71441e-19 $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_268 N_A_M1009_g N_VPWR_c_472_n 0.0137849f $X=2.645 $Y=2.53 $X2=0 $Y2=0
cc_269 N_A_M1000_g N_VPWR_c_473_n 0.00100512f $X=3.885 $Y=0.835 $X2=0 $Y2=0
cc_270 N_A_M1009_g N_VPWR_c_476_n 0.00434252f $X=2.645 $Y=2.53 $X2=0 $Y2=0
cc_271 N_A_M1009_g N_VPWR_c_470_n 0.00479212f $X=2.645 $Y=2.53 $X2=0 $Y2=0
cc_272 N_A_M1000_g COUT 0.00224589f $X=3.885 $Y=0.835 $X2=0 $Y2=0
cc_273 N_A_c_383_n N_VGND_c_543_n 0.0186992f $X=3.81 $Y=0.18 $X2=0 $Y2=0
cc_274 N_A_c_378_n N_VGND_c_546_n 0.00419075f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_275 N_A_c_379_n N_VGND_c_546_n 4.70115e-19 $X=2.865 $Y=0.84 $X2=0 $Y2=0
cc_276 N_A_c_384_n N_VGND_c_546_n 0.0403985f $X=3.015 $Y=0.18 $X2=0 $Y2=0
cc_277 N_A_c_378_n N_VGND_c_548_n 0.00635917f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_278 N_A_c_383_n N_VGND_c_548_n 0.0361099f $X=3.81 $Y=0.18 $X2=0 $Y2=0
cc_279 N_A_c_384_n N_VGND_c_548_n 0.0102835f $X=3.015 $Y=0.18 $X2=0 $Y2=0
cc_280 N_A_c_378_n N_VGND_c_550_n 0.00423616f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_281 N_A_c_378_n N_A_301_47#_c_595_n 0.0139628f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_282 N_A_c_380_n N_A_301_47#_c_595_n 0.00460692f $X=2.645 $Y=1.405 $X2=0 $Y2=0
cc_283 N_A_c_386_n N_A_301_47#_c_595_n 0.0183815f $X=2.345 $Y=1.215 $X2=0 $Y2=0
cc_284 N_A_c_378_n N_A_301_47#_c_597_n 3.20799e-19 $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_285 N_A_c_379_n N_A_301_47#_c_597_n 0.00564389f $X=2.865 $Y=0.84 $X2=0 $Y2=0
cc_286 N_A_c_380_n N_A_301_47#_c_597_n 3.35749e-19 $X=2.645 $Y=1.405 $X2=0 $Y2=0
cc_287 N_A_c_382_n N_A_301_47#_c_597_n 0.0102212f $X=2.94 $Y=0.765 $X2=0 $Y2=0
cc_288 N_SUM_c_446_n N_VPWR_c_471_n 0.0192235f $X=0.925 $Y=2.595 $X2=0 $Y2=0
cc_289 N_SUM_c_446_n N_VPWR_c_474_n 0.0189623f $X=0.925 $Y=2.595 $X2=0 $Y2=0
cc_290 SUM N_VPWR_c_474_n 0.00987967f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_291 N_SUM_c_446_n N_VPWR_c_470_n 0.0221316f $X=0.925 $Y=2.595 $X2=0 $Y2=0
cc_292 SUM N_VPWR_c_470_n 0.0112661f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_293 SUM N_VGND_c_544_n 0.00871478f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_294 SUM N_VGND_c_548_n 0.0111671f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_295 N_VPWR_c_473_n COUT 0.0255623f $X=4.1 $Y=2.29 $X2=0 $Y2=0
cc_296 N_VPWR_c_479_n COUT 0.00653615f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_297 N_VPWR_c_470_n COUT 0.0074472f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_298 COUT N_VGND_c_543_n 0.00936443f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_299 COUT N_VGND_c_547_n 0.00653615f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_300 COUT N_VGND_c_548_n 0.0074472f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_301 N_VGND_c_548_n N_A_301_47#_M1011_d 0.00366446f $X=4.56 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_302 N_VGND_c_548_n N_A_301_47#_M1007_d 0.00288373f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_303 N_VGND_M1006_d N_A_301_47#_c_595_n 0.00364078f $X=1.935 $Y=0.235 $X2=0
+ $Y2=0
cc_304 N_VGND_c_545_n N_A_301_47#_c_595_n 0.00366601f $X=1.99 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_c_546_n N_A_301_47#_c_595_n 0.00366601f $X=3.995 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_c_548_n N_A_301_47#_c_595_n 0.0142336f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_550_n N_A_301_47#_c_595_n 0.023293f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_308 N_VGND_c_545_n N_A_301_47#_c_596_n 0.00809875f $X=1.99 $Y=0 $X2=0 $Y2=0
cc_309 N_VGND_c_548_n N_A_301_47#_c_596_n 0.00758505f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_546_n N_A_301_47#_c_597_n 0.00850877f $X=3.995 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_548_n N_A_301_47#_c_597_n 0.00758505f $X=4.56 $Y=0 $X2=0 $Y2=0
