* File: sky130_fd_sc_lp__a21o_1.pxi.spice
* Created: Wed Sep  2 09:19:55 2020
* 
x_PM_SKY130_FD_SC_LP__A21O_1%A_80_237# N_A_80_237#_M1003_d N_A_80_237#_M1001_s
+ N_A_80_237#_M1007_g N_A_80_237#_c_50_n N_A_80_237#_M1000_g N_A_80_237#_c_51_n
+ N_A_80_237#_c_52_n N_A_80_237#_c_53_n N_A_80_237#_c_57_n N_A_80_237#_c_58_n
+ N_A_80_237#_c_99_p N_A_80_237#_c_54_n PM_SKY130_FD_SC_LP__A21O_1%A_80_237#
x_PM_SKY130_FD_SC_LP__A21O_1%B1 N_B1_M1003_g N_B1_M1001_g B1 N_B1_c_104_n
+ N_B1_c_105_n PM_SKY130_FD_SC_LP__A21O_1%B1
x_PM_SKY130_FD_SC_LP__A21O_1%A1 N_A1_M1002_g N_A1_M1006_g A1 A1 A1 N_A1_c_142_n
+ N_A1_c_143_n PM_SKY130_FD_SC_LP__A21O_1%A1
x_PM_SKY130_FD_SC_LP__A21O_1%A2 N_A2_M1005_g N_A2_M1004_g A2 N_A2_c_177_n
+ N_A2_c_178_n PM_SKY130_FD_SC_LP__A21O_1%A2
x_PM_SKY130_FD_SC_LP__A21O_1%X N_X_M1000_s N_X_M1007_s X X X X X X X N_X_c_198_n
+ PM_SKY130_FD_SC_LP__A21O_1%X
x_PM_SKY130_FD_SC_LP__A21O_1%VPWR N_VPWR_M1007_d N_VPWR_M1006_d N_VPWR_c_211_n
+ N_VPWR_c_212_n VPWR N_VPWR_c_213_n N_VPWR_c_214_n N_VPWR_c_215_n
+ N_VPWR_c_210_n N_VPWR_c_217_n N_VPWR_c_218_n PM_SKY130_FD_SC_LP__A21O_1%VPWR
x_PM_SKY130_FD_SC_LP__A21O_1%A_300_367# N_A_300_367#_M1001_d
+ N_A_300_367#_M1004_d N_A_300_367#_c_265_n N_A_300_367#_c_249_n
+ N_A_300_367#_c_250_n N_A_300_367#_c_251_n
+ PM_SKY130_FD_SC_LP__A21O_1%A_300_367#
x_PM_SKY130_FD_SC_LP__A21O_1%VGND N_VGND_M1000_d N_VGND_M1005_d N_VGND_c_271_n
+ N_VGND_c_272_n N_VGND_c_273_n VGND N_VGND_c_274_n N_VGND_c_275_n
+ N_VGND_c_276_n N_VGND_c_277_n PM_SKY130_FD_SC_LP__A21O_1%VGND
cc_1 VNB N_A_80_237#_M1007_g 0.00896044f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB N_A_80_237#_c_50_n 0.0215218f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.185
cc_3 VNB N_A_80_237#_c_51_n 0.0123297f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.515
cc_4 VNB N_A_80_237#_c_52_n 0.0019435f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.92
cc_5 VNB N_A_80_237#_c_53_n 0.0117164f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.07
cc_6 VNB N_A_80_237#_c_54_n 0.0484052f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.35
cc_7 VNB N_B1_M1003_g 0.0281418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_104_n 0.0293204f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.655
cc_9 VNB N_B1_c_105_n 0.00377017f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.655
cc_10 VNB N_A1_M1006_g 0.00802835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A1 0.0024827f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_12 VNB A1 0.00767634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_142_n 0.0309799f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.92
cc_14 VNB N_A1_c_143_n 0.0187028f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.07
cc_15 VNB N_A2_M1004_g 0.0119208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A2 0.0163382f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_17 VNB N_A2_c_177_n 0.0383763f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.185
cc_18 VNB N_A2_c_178_n 0.0225381f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.655
cc_19 VNB N_X_c_198_n 0.0614634f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.985
cc_20 VNB N_VPWR_c_210_n 0.123877f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=2.01
cc_21 VNB N_VGND_c_271_n 0.00203511f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_22 VNB N_VGND_c_272_n 0.0110036f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.185
cc_23 VNB N_VGND_c_273_n 0.0331498f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.655
cc_24 VNB N_VGND_c_274_n 0.015535f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.07
cc_25 VNB N_VGND_c_275_n 0.0309273f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.985
cc_26 VNB N_VGND_c_276_n 0.0108457f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.35
cc_27 VNB N_VGND_c_277_n 0.168858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A_80_237#_M1007_g 0.0258819f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_29 VPB N_A_80_237#_c_52_n 0.00534499f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.92
cc_30 VPB N_A_80_237#_c_57_n 0.0152569f $X=-0.19 $Y=1.655 $X2=1.18 $Y2=2.1
cc_31 VPB N_A_80_237#_c_58_n 0.0101063f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=2.91
cc_32 VPB N_B1_M1001_g 0.0233498f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.515
cc_33 VPB N_B1_c_104_n 0.00802101f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.655
cc_34 VPB N_B1_c_105_n 0.00442997f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.655
cc_35 VPB N_A1_M1006_g 0.0198757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A2_M1004_g 0.0255526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_X_c_198_n 0.0565224f $X=-0.19 $Y=1.655 $X2=1.555 $Y2=0.985
cc_38 VPB N_VPWR_c_211_n 0.0106971f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_39 VPB N_VPWR_c_212_n 0.00561552f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.655
cc_40 VPB N_VPWR_c_213_n 0.0153759f $X=-0.19 $Y=1.655 $X2=1.18 $Y2=2.91
cc_41 VPB N_VPWR_c_214_n 0.0308098f $X=-0.19 $Y=1.655 $X2=1.555 $Y2=0.42
cc_42 VPB N_VPWR_c_215_n 0.0180549f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_210_n 0.0537057f $X=-0.19 $Y=1.655 $X2=1.18 $Y2=2.01
cc_44 VPB N_VPWR_c_217_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.35
cc_45 VPB N_VPWR_c_218_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.35
cc_46 VPB N_A_300_367#_c_249_n 0.0144956f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.655
cc_47 VPB N_A_300_367#_c_250_n 0.0050726f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.515
cc_48 VPB N_A_300_367#_c_251_n 0.0470363f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=1.07
cc_49 N_A_80_237#_c_50_n N_B1_M1003_g 0.00512052f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_50 N_A_80_237#_c_51_n N_B1_M1003_g 0.00158409f $X=0.8 $Y=1.515 $X2=0 $Y2=0
cc_51 N_A_80_237#_c_53_n N_B1_M1003_g 0.0155486f $X=1.39 $Y=1.07 $X2=0 $Y2=0
cc_52 N_A_80_237#_c_54_n N_B1_M1003_g 0.00586378f $X=0.69 $Y=1.35 $X2=0 $Y2=0
cc_53 N_A_80_237#_c_52_n N_B1_M1001_g 0.00273921f $X=0.8 $Y=1.92 $X2=0 $Y2=0
cc_54 N_A_80_237#_M1007_g N_B1_c_104_n 0.00213849f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_55 N_A_80_237#_c_52_n N_B1_c_104_n 5.21031e-19 $X=0.8 $Y=1.92 $X2=0 $Y2=0
cc_56 N_A_80_237#_c_53_n N_B1_c_104_n 0.0061827f $X=1.39 $Y=1.07 $X2=0 $Y2=0
cc_57 N_A_80_237#_c_57_n N_B1_c_104_n 0.00105054f $X=1.18 $Y=2.1 $X2=0 $Y2=0
cc_58 N_A_80_237#_c_54_n N_B1_c_104_n 0.00937535f $X=0.69 $Y=1.35 $X2=0 $Y2=0
cc_59 N_A_80_237#_c_51_n N_B1_c_105_n 0.013605f $X=0.8 $Y=1.515 $X2=0 $Y2=0
cc_60 N_A_80_237#_c_52_n N_B1_c_105_n 0.0185927f $X=0.8 $Y=1.92 $X2=0 $Y2=0
cc_61 N_A_80_237#_c_53_n N_B1_c_105_n 0.0228593f $X=1.39 $Y=1.07 $X2=0 $Y2=0
cc_62 N_A_80_237#_c_57_n N_B1_c_105_n 0.0199357f $X=1.18 $Y=2.1 $X2=0 $Y2=0
cc_63 N_A_80_237#_c_54_n N_B1_c_105_n 5.73063e-19 $X=0.69 $Y=1.35 $X2=0 $Y2=0
cc_64 N_A_80_237#_c_53_n A1 0.00558588f $X=1.39 $Y=1.07 $X2=0 $Y2=0
cc_65 N_A_80_237#_c_53_n N_A1_c_143_n 0.00121953f $X=1.39 $Y=1.07 $X2=0 $Y2=0
cc_66 N_A_80_237#_c_50_n N_X_c_198_n 0.00506418f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_67 N_A_80_237#_c_51_n N_X_c_198_n 0.0337182f $X=0.8 $Y=1.515 $X2=0 $Y2=0
cc_68 N_A_80_237#_c_52_n N_X_c_198_n 0.0164966f $X=0.8 $Y=1.92 $X2=0 $Y2=0
cc_69 N_A_80_237#_c_54_n N_X_c_198_n 0.0204002f $X=0.69 $Y=1.35 $X2=0 $Y2=0
cc_70 N_A_80_237#_c_52_n N_VPWR_M1007_d 0.00172644f $X=0.8 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A_80_237#_c_57_n N_VPWR_M1007_d 0.0044012f $X=1.18 $Y=2.1 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_80_237#_M1007_g N_VPWR_c_211_n 0.020417f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A_80_237#_c_57_n N_VPWR_c_211_n 0.0114373f $X=1.18 $Y=2.1 $X2=0 $Y2=0
cc_74 N_A_80_237#_c_58_n N_VPWR_c_211_n 0.0610596f $X=1.21 $Y=2.91 $X2=0 $Y2=0
cc_75 N_A_80_237#_M1007_g N_VPWR_c_213_n 0.00486043f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_76 N_A_80_237#_c_58_n N_VPWR_c_214_n 0.0181659f $X=1.21 $Y=2.91 $X2=0 $Y2=0
cc_77 N_A_80_237#_M1001_s N_VPWR_c_210_n 0.00336915f $X=1.085 $Y=1.835 $X2=0
+ $Y2=0
cc_78 N_A_80_237#_M1007_g N_VPWR_c_210_n 0.00917987f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_79 N_A_80_237#_c_58_n N_VPWR_c_210_n 0.0104192f $X=1.21 $Y=2.91 $X2=0 $Y2=0
cc_80 N_A_80_237#_c_52_n N_A_300_367#_c_250_n 0.00297956f $X=0.8 $Y=1.92 $X2=0
+ $Y2=0
cc_81 N_A_80_237#_c_53_n N_A_300_367#_c_250_n 0.00511699f $X=1.39 $Y=1.07 $X2=0
+ $Y2=0
cc_82 N_A_80_237#_c_51_n N_VGND_M1000_d 0.00312785f $X=0.8 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_83 N_A_80_237#_c_53_n N_VGND_M1000_d 0.00281447f $X=1.39 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_80_237#_c_50_n N_VGND_c_271_n 0.0130406f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_85 N_A_80_237#_c_51_n N_VGND_c_271_n 0.0221701f $X=0.8 $Y=1.515 $X2=0 $Y2=0
cc_86 N_A_80_237#_c_53_n N_VGND_c_271_n 0.0223333f $X=1.39 $Y=1.07 $X2=0 $Y2=0
cc_87 N_A_80_237#_c_54_n N_VGND_c_271_n 0.00175095f $X=0.69 $Y=1.35 $X2=0 $Y2=0
cc_88 N_A_80_237#_c_50_n N_VGND_c_274_n 0.00486043f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_89 N_A_80_237#_c_99_p N_VGND_c_275_n 0.0214254f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_90 N_A_80_237#_M1003_d N_VGND_c_277_n 0.00547617f $X=1.345 $Y=0.235 $X2=0
+ $Y2=0
cc_91 N_A_80_237#_c_50_n N_VGND_c_277_n 0.00918457f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_92 N_A_80_237#_c_99_p N_VGND_c_277_n 0.0127519f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_93 N_B1_c_104_n N_A1_M1006_g 0.0260695f $X=1.29 $Y=1.51 $X2=0 $Y2=0
cc_94 N_B1_c_105_n N_A1_M1006_g 8.9055e-19 $X=1.29 $Y=1.51 $X2=0 $Y2=0
cc_95 N_B1_M1003_g A1 9.10057e-19 $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_96 N_B1_c_104_n A1 6.82046e-19 $X=1.29 $Y=1.51 $X2=0 $Y2=0
cc_97 N_B1_c_105_n A1 0.00729005f $X=1.29 $Y=1.51 $X2=0 $Y2=0
cc_98 N_B1_c_104_n N_A1_c_142_n 0.00917207f $X=1.29 $Y=1.51 $X2=0 $Y2=0
cc_99 N_B1_M1003_g N_A1_c_143_n 0.0221412f $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_100 N_B1_M1001_g N_VPWR_c_211_n 0.00355208f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_101 N_B1_M1001_g N_VPWR_c_214_n 0.00585385f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_102 N_B1_M1001_g N_VPWR_c_210_n 0.0120903f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_103 N_B1_M1001_g N_A_300_367#_c_250_n 0.00191686f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_B1_c_105_n N_A_300_367#_c_250_n 0.00548086f $X=1.29 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B1_M1003_g N_VGND_c_271_n 0.0123281f $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_106 N_B1_M1003_g N_VGND_c_275_n 0.00486043f $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_107 N_B1_M1003_g N_VGND_c_277_n 0.00865379f $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_108 N_A1_M1006_g N_A2_M1004_g 0.019289f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_109 A1 A2 0.0273822f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A1_c_142_n A2 2.5152e-19 $X=1.905 $Y=1.35 $X2=0 $Y2=0
cc_111 A1 N_A2_c_177_n 0.00264386f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_112 N_A1_c_142_n N_A2_c_177_n 0.0172946f $X=1.905 $Y=1.35 $X2=0 $Y2=0
cc_113 A1 N_A2_c_178_n 0.00749311f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_114 N_A1_c_143_n N_A2_c_178_n 0.0228977f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_115 N_A1_M1006_g N_VPWR_c_212_n 0.00355081f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A1_M1006_g N_VPWR_c_214_n 0.00585385f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A1_M1006_g N_VPWR_c_210_n 0.0108498f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A1_M1006_g N_A_300_367#_c_249_n 0.0148391f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_119 A1 N_A_300_367#_c_249_n 0.0384945f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_120 N_A1_c_142_n N_A_300_367#_c_249_n 0.0040593f $X=1.905 $Y=1.35 $X2=0 $Y2=0
cc_121 A1 N_A_300_367#_c_250_n 4.21667e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A1_c_143_n N_VGND_c_271_n 0.00109708f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_123 N_A1_c_143_n N_VGND_c_273_n 0.00146738f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_124 A1 N_VGND_c_275_n 0.0140182f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_125 N_A1_c_143_n N_VGND_c_275_n 0.00585385f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_126 A1 N_VGND_c_277_n 0.0116227f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_127 N_A1_c_143_n N_VGND_c_277_n 0.011501f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_128 A1 A_378_47# 0.0148429f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_129 N_A2_M1004_g N_VPWR_c_212_n 0.00362135f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A2_M1004_g N_VPWR_c_215_n 0.00585385f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A2_M1004_g N_VPWR_c_210_n 0.0117482f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A2_M1004_g N_A_300_367#_c_249_n 0.0199708f $X=2.385 $Y=2.465 $X2=0
+ $Y2=0
cc_133 A2 N_A_300_367#_c_249_n 0.0285587f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A2_c_177_n N_A_300_367#_c_249_n 0.00500857f $X=2.51 $Y=1.35 $X2=0 $Y2=0
cc_135 A2 N_VGND_c_273_n 0.0248549f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_136 N_A2_c_177_n N_VGND_c_273_n 0.00483488f $X=2.51 $Y=1.35 $X2=0 $Y2=0
cc_137 N_A2_c_178_n N_VGND_c_273_n 0.0186921f $X=2.492 $Y=1.185 $X2=0 $Y2=0
cc_138 N_A2_c_178_n N_VGND_c_275_n 0.00486043f $X=2.492 $Y=1.185 $X2=0 $Y2=0
cc_139 N_A2_c_178_n N_VGND_c_277_n 0.00870566f $X=2.492 $Y=1.185 $X2=0 $Y2=0
cc_140 N_X_c_198_n N_VPWR_c_213_n 0.0178111f $X=0.265 $Y=0.42 $X2=0 $Y2=0
cc_141 N_X_M1007_s N_VPWR_c_210_n 0.00371702f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_142 N_X_c_198_n N_VPWR_c_210_n 0.0100304f $X=0.265 $Y=0.42 $X2=0 $Y2=0
cc_143 N_X_c_198_n N_VGND_c_274_n 0.0179921f $X=0.265 $Y=0.42 $X2=0 $Y2=0
cc_144 N_X_M1000_s N_VGND_c_277_n 0.00389096f $X=0.14 $Y=0.235 $X2=0 $Y2=0
cc_145 N_X_c_198_n N_VGND_c_277_n 0.0100304f $X=0.265 $Y=0.42 $X2=0 $Y2=0
cc_146 N_VPWR_c_210_n N_A_300_367#_M1001_d 0.00536646f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_147 N_VPWR_c_210_n N_A_300_367#_M1004_d 0.00215158f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_148 N_VPWR_c_214_n N_A_300_367#_c_265_n 0.0124525f $X=1.96 $Y=3.33 $X2=0
+ $Y2=0
cc_149 N_VPWR_c_210_n N_A_300_367#_c_265_n 0.00730372f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_150 N_VPWR_M1006_d N_A_300_367#_c_249_n 0.00284866f $X=1.93 $Y=1.835 $X2=0
+ $Y2=0
cc_151 N_VPWR_c_212_n N_A_300_367#_c_249_n 0.0216414f $X=2.125 $Y=2.11 $X2=0
+ $Y2=0
cc_152 N_VPWR_c_215_n N_A_300_367#_c_251_n 0.0194077f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_153 N_VPWR_c_210_n N_A_300_367#_c_251_n 0.0117799f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_154 N_VGND_c_277_n A_378_47# 0.00720532f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
