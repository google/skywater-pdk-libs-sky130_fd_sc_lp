* NGSPICE file created from sky130_fd_sc_lp__nor2_8.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor2_8 A B VGND VNB VPB VPWR Y
M1000 VPWR A a_47_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.4112e+12p pd=1.232e+07u as=3.1374e+12p ps=2.766e+07u
M1001 a_47_367# B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.4112e+12p ps=1.232e+07u
M1002 Y B a_47_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B VGND VNB nshort w=840000u l=150000u
+  ad=1.8816e+12p pd=1.792e+07u as=2.1e+12p ps=2.012e+07u
M1004 VPWR A a_47_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_47_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_47_367# B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_47_367# B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A a_47_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_47_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B a_47_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_47_367# B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND B Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_47_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B a_47_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_47_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND B Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y B a_47_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND B Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_47_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

