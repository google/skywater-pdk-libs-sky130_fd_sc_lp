* File: sky130_fd_sc_lp__and3_2.pex.spice
* Created: Wed Sep  2 09:31:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3_2%A 1 3 4 6 10 12 13 16 17
r35 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.1 $X2=0.275 $Y2=1.1
r36 13 17 0.820838 $w=5.08e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.27
+ $X2=0.275 $Y2=1.27
r37 12 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.275 $Y=1.44
+ $X2=0.275 $Y2=1.1
r38 8 16 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.275 $Y=0.915
+ $X2=0.275 $Y2=1.1
r39 8 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.275 $Y=0.84
+ $X2=0.545 $Y2=0.84
r40 4 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.545 $Y=0.765
+ $X2=0.545 $Y2=0.84
r41 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.545 $Y=0.765
+ $X2=0.545 $Y2=0.445
r42 1 12 66.2088 $w=2.73e-07 $l=4.64354e-07 $layer=POLY_cond $X=0.475 $Y=1.815
+ $X2=0.275 $Y2=1.44
r43 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=1.815
+ $X2=0.475 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_2%B 3 7 9 12 13
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.815 $Y=1.29
+ $X2=0.815 $Y2=1.455
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.815 $Y=1.29
+ $X2=0.815 $Y2=1.125
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.815
+ $Y=1.29 $X2=0.815 $Y2=1.29
r37 9 13 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=1.29
+ $X2=0.815 $Y2=1.29
r38 7 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.905 $Y=2.135
+ $X2=0.905 $Y2=1.455
r39 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.905 $Y=0.445
+ $X2=0.905 $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_2%C 3 7 9 12 13
c39 13 0 8.10772e-20 $X=1.355 $Y=1.35
r40 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=1.515
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=1.185
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.355
+ $Y=1.35 $X2=1.355 $Y2=1.35
r43 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=1.35
+ $X2=1.355 $Y2=1.35
r44 7 15 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.41 $Y=2.135
+ $X2=1.41 $Y2=1.515
r45 3 14 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.265 $Y=0.445
+ $X2=1.265 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_2%A_27_385# 1 2 3 12 16 18 22 26 28 31 35 37 38
+ 39 40 43 45 48 49 51 54
c109 12 0 8.10772e-20 $X=1.935 $Y=0.655
r110 54 55 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.895 $Y=1.35
+ $X2=1.895 $Y2=1.275
r111 52 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.44
+ $X2=1.895 $Y2=1.605
r112 52 54 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.895 $Y=1.44
+ $X2=1.895 $Y2=1.35
r113 51 53 18.3262 $w=2.33e-07 $l=3.5e-07 $layer=LI1_cond $X=1.837 $Y=1.44
+ $X2=1.837 $Y2=1.79
r114 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.895
+ $Y=1.44 $X2=1.895 $Y2=1.44
r115 48 51 9.55378 $w=2.33e-07 $l=1.9139e-07 $layer=LI1_cond $X=1.78 $Y=1.275
+ $X2=1.837 $Y2=1.44
r116 47 48 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.78 $Y=0.845
+ $X2=1.78 $Y2=1.275
r117 46 49 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.29 $Y=1.79
+ $X2=1.14 $Y2=1.79
r118 45 53 2.58477 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.695 $Y=1.79
+ $X2=1.837 $Y2=1.79
r119 45 46 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.695 $Y=1.79
+ $X2=1.29 $Y2=1.79
r120 41 49 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.875
+ $X2=1.14 $Y2=1.79
r121 41 43 9.98784 $w=2.98e-07 $l=2.6e-07 $layer=LI1_cond $X=1.14 $Y=1.875
+ $X2=1.14 $Y2=2.135
r122 39 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.695 $Y=0.76
+ $X2=1.78 $Y2=0.845
r123 39 40 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=1.695 $Y=0.76
+ $X2=0.495 $Y2=0.76
r124 37 49 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.99 $Y=1.79
+ $X2=1.14 $Y2=1.79
r125 37 38 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.99 $Y=1.79 $X2=0.39
+ $Y2=1.79
r126 33 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.33 $Y=0.675
+ $X2=0.495 $Y2=0.76
r127 33 35 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.33 $Y=0.675
+ $X2=0.33 $Y2=0.42
r128 29 38 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=0.242 $Y=1.875
+ $X2=0.39 $Y2=1.79
r129 29 31 10.1571 $w=2.93e-07 $l=2.6e-07 $layer=LI1_cond $X=0.242 $Y=1.875
+ $X2=0.242 $Y2=2.135
r130 24 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.365 $Y=1.425
+ $X2=2.365 $Y2=1.35
r131 24 26 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.365 $Y=1.425
+ $X2=2.365 $Y2=2.465
r132 20 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.365 $Y=1.275
+ $X2=2.365 $Y2=1.35
r133 20 22 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.365 $Y=1.275
+ $X2=2.365 $Y2=0.655
r134 19 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.35
+ $X2=1.895 $Y2=1.35
r135 18 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.29 $Y=1.35
+ $X2=2.365 $Y2=1.35
r136 18 19 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.29 $Y=1.35
+ $X2=2.06 $Y2=1.35
r137 16 57 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.935 $Y=2.465
+ $X2=1.935 $Y2=1.605
r138 12 55 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.935 $Y=0.655
+ $X2=1.935 $Y2=1.275
r139 3 43 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.925 $X2=1.155 $Y2=2.135
r140 2 31 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.925 $X2=0.26 $Y2=2.135
r141 1 35 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.235 $X2=0.33 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_2%VPWR 1 2 3 12 16 20 22 26 28 33 38 44 47 51
r34 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 42 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 39 47 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=1.855 $Y=3.33
+ $X2=1.657 $Y2=3.33
r41 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.855 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 38 50 4.09051 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.5 $Y=3.33 $X2=2.69
+ $Y2=3.33
r43 38 41 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.5 $Y=3.33 $X2=2.16
+ $Y2=3.33
r44 37 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 34 44 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.82 $Y=3.33 $X2=0.69
+ $Y2=3.33
r47 34 36 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 33 47 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=1.46 $Y=3.33
+ $X2=1.657 $Y2=3.33
r49 33 36 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.46 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 28 44 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.69
+ $Y2=3.33
r53 28 30 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r54 26 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 26 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 22 25 42.995 $w=2.58e-07 $l=9.7e-07 $layer=LI1_cond $X=2.63 $Y=1.98 $X2=2.63
+ $Y2=2.95
r57 20 50 3.12171 $w=2.6e-07 $l=1.11018e-07 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.69 $Y2=3.33
r58 20 25 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=2.95
r59 16 19 12.2538 $w=3.93e-07 $l=4.2e-07 $layer=LI1_cond $X=1.657 $Y=2.13
+ $X2=1.657 $Y2=2.55
r60 14 47 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.657 $Y=3.245
+ $X2=1.657 $Y2=3.33
r61 14 19 20.2772 $w=3.93e-07 $l=6.95e-07 $layer=LI1_cond $X=1.657 $Y=3.245
+ $X2=1.657 $Y2=2.55
r62 10 44 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r63 10 12 45.8761 $w=2.58e-07 $l=1.035e-06 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.21
r64 3 25 400 $w=1.7e-07 $l=1.18998e-06 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.835 $X2=2.595 $Y2=2.95
r65 3 22 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.835 $X2=2.595 $Y2=1.98
r66 2 19 300 $w=1.7e-07 $l=7.33144e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.925 $X2=1.72 $Y2=2.55
r67 2 16 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.925 $X2=1.625 $Y2=2.13
r68 1 12 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.925 $X2=0.69 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_2%X 1 2 9 13 14 15 16 24 34
r32 21 24 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=2.182 $Y=1.962
+ $X2=2.182 $Y2=1.98
r33 16 31 5.27389 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=2.182 $Y=2.775
+ $X2=2.182 $Y2=2.91
r34 15 16 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.182 $Y=2.405
+ $X2=2.182 $Y2=2.775
r35 14 21 0.234395 $w=2.93e-07 $l=6e-09 $layer=LI1_cond $X=2.182 $Y=1.956
+ $X2=2.182 $Y2=1.962
r36 14 34 7.24732 $w=2.93e-07 $l=1.41e-07 $layer=LI1_cond $X=2.182 $Y=1.956
+ $X2=2.182 $Y2=1.815
r37 14 15 14.22 $w=2.93e-07 $l=3.64e-07 $layer=LI1_cond $X=2.182 $Y=2.041
+ $X2=2.182 $Y2=2.405
r38 14 24 2.38302 $w=2.93e-07 $l=6.1e-08 $layer=LI1_cond $X=2.182 $Y=2.041
+ $X2=2.182 $Y2=1.98
r39 13 34 44.3636 $w=1.78e-07 $l=7.2e-07 $layer=LI1_cond $X=2.24 $Y=1.095
+ $X2=2.24 $Y2=1.815
r40 7 13 6.93297 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=2.197 $Y=0.963
+ $X2=2.197 $Y2=1.095
r41 7 9 23.6142 $w=2.63e-07 $l=5.43e-07 $layer=LI1_cond $X=2.197 $Y=0.963
+ $X2=2.197 $Y2=0.42
r42 2 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.15 $Y2=2.91
r43 2 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.15 $Y2=1.98
r44 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.235 $X2=2.15 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_2%VGND 1 2 9 11 13 15 17 25 31 35
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r39 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r40 29 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r41 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 26 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.61
+ $Y2=0
r43 26 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=2.16
+ $Y2=0
r44 25 34 4.09051 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.69
+ $Y2=0
r45 25 28 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.16
+ $Y2=0
r46 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 20 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r48 19 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r49 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.61
+ $Y2=0
r51 17 23 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.2
+ $Y2=0
r52 15 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r53 15 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r54 11 34 3.12171 $w=2.6e-07 $l=1.11018e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.69 $Y2=0
r55 11 13 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.38
r56 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=0.085 $X2=1.61
+ $Y2=0
r57 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.61 $Y=0.085
+ $X2=1.61 $Y2=0.38
r58 2 13 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.44
+ $Y=0.235 $X2=2.595 $Y2=0.38
r59 1 9 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.235 $X2=1.61 $Y2=0.38
.ends

