* File: sky130_fd_sc_lp__xnor2_0.pxi.spice
* Created: Wed Sep  2 10:39:54 2020
* 
x_PM_SKY130_FD_SC_LP__XNOR2_0%A N_A_M1006_g N_A_M1000_g N_A_c_74_n N_A_c_75_n
+ N_A_c_76_n N_A_c_77_n N_A_M1003_g N_A_M1005_g N_A_c_88_n N_A_c_89_n N_A_c_79_n
+ N_A_c_80_n N_A_c_81_n N_A_c_82_n A A N_A_c_84_n N_A_c_85_n
+ PM_SKY130_FD_SC_LP__XNOR2_0%A
x_PM_SKY130_FD_SC_LP__XNOR2_0%B N_B_c_157_n N_B_M1001_g N_B_M1004_g N_B_M1007_g
+ N_B_M1009_g N_B_c_159_n N_B_c_166_n B B N_B_c_161_n N_B_c_162_n
+ PM_SKY130_FD_SC_LP__XNOR2_0%B
x_PM_SKY130_FD_SC_LP__XNOR2_0%A_143_487# N_A_143_487#_M1001_d
+ N_A_143_487#_M1000_d N_A_143_487#_M1008_g N_A_143_487#_M1002_g
+ N_A_143_487#_c_238_n N_A_143_487#_c_232_n N_A_143_487#_c_233_n
+ N_A_143_487#_c_285_p N_A_143_487#_c_234_n N_A_143_487#_c_240_n
+ N_A_143_487#_c_241_n N_A_143_487#_c_270_n N_A_143_487#_c_235_n
+ N_A_143_487#_c_243_n N_A_143_487#_c_236_n N_A_143_487#_c_244_n
+ PM_SKY130_FD_SC_LP__XNOR2_0%A_143_487#
x_PM_SKY130_FD_SC_LP__XNOR2_0%VPWR N_VPWR_M1000_s N_VPWR_M1004_d N_VPWR_M1008_d
+ N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n VPWR N_VPWR_c_314_n
+ N_VPWR_c_324_n PM_SKY130_FD_SC_LP__XNOR2_0%VPWR
x_PM_SKY130_FD_SC_LP__XNOR2_0%Y N_Y_M1002_d N_Y_M1007_d N_Y_c_362_n N_Y_c_359_n
+ N_Y_c_360_n N_Y_c_356_n Y Y Y N_Y_c_358_n PM_SKY130_FD_SC_LP__XNOR2_0%Y
x_PM_SKY130_FD_SC_LP__XNOR2_0%VGND N_VGND_M1006_s N_VGND_M1003_d N_VGND_c_397_n
+ N_VGND_c_398_n N_VGND_c_399_n VGND N_VGND_c_400_n N_VGND_c_401_n
+ N_VGND_c_402_n N_VGND_c_403_n PM_SKY130_FD_SC_LP__XNOR2_0%VGND
x_PM_SKY130_FD_SC_LP__XNOR2_0%A_300_60# N_A_300_60#_M1003_s N_A_300_60#_M1009_d
+ N_A_300_60#_c_436_n N_A_300_60#_c_437_n N_A_300_60#_c_438_n
+ N_A_300_60#_c_439_n PM_SKY130_FD_SC_LP__XNOR2_0%A_300_60#
cc_1 VNB N_A_M1006_g 0.0285484f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.095
cc_2 VNB N_A_c_74_n 0.0198258f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=0.83
cc_3 VNB N_A_c_75_n 0.0208217f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.905
cc_4 VNB N_A_c_76_n 0.00959019f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.905
cc_5 VNB N_A_c_77_n 0.0179119f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.83
cc_6 VNB N_A_M1005_g 0.0346092f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.755
cc_7 VNB N_A_c_79_n 0.00446978f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.905
cc_8 VNB N_A_c_80_n 0.00758209f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.43
cc_9 VNB N_A_c_81_n 0.00531388f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.385
cc_10 VNB N_A_c_82_n 0.00767297f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.35
cc_11 VNB A 0.0145658f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_12 VNB N_A_c_84_n 0.0117329f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.74
cc_13 VNB N_A_c_85_n 0.0509065f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=0.35
cc_14 VNB N_B_c_157_n 0.018243f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.575
cc_15 VNB N_B_M1009_g 0.0365168f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.51
cc_16 VNB N_B_c_159_n 0.0149611f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.755
cc_17 VNB B 0.0147277f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.575
cc_18 VNB N_B_c_161_n 0.0143144f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.905
cc_19 VNB N_B_c_162_n 0.0481013f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.385
cc_20 VNB N_A_143_487#_c_232_n 0.021261f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.755
cc_21 VNB N_A_143_487#_c_233_n 0.0220633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_143_487#_c_234_n 0.00187771f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.905
cc_23 VNB N_A_143_487#_c_235_n 0.0537954f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_143_487#_c_236_n 0.00515713f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.74
cc_25 VNB N_VPWR_c_314_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_356_n 0.012834f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.83
cc_27 VNB Y 0.0151727f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.98
cc_28 VNB N_Y_c_358_n 0.0365709f $X=-0.19 $Y=-0.245 $X2=0.467 $Y2=2.095
cc_29 VNB N_VGND_c_397_n 0.0106171f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.755
cc_30 VNB N_VGND_c_398_n 0.0552944f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=0.515
cc_31 VNB N_VGND_c_399_n 0.00709023f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.83
cc_32 VNB N_VGND_c_400_n 0.0396683f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.755
cc_33 VNB N_VGND_c_401_n 0.0338082f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.43
cc_34 VNB N_VGND_c_402_n 0.208451f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.385
cc_35 VNB N_VGND_c_403_n 0.00490486f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_36 VNB N_A_300_60#_c_436_n 0.00194462f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=0.515
cc_37 VNB N_A_300_60#_c_437_n 0.0123577f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.905
cc_38 VNB N_A_300_60#_c_438_n 0.002985f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.905
cc_39 VNB N_A_300_60#_c_439_n 0.00191629f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.51
cc_40 VPB N_A_M1000_g 0.0276139f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.755
cc_41 VPB N_A_M1005_g 0.0484744f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.755
cc_42 VPB N_A_c_88_n 0.0291007f $X=-0.19 $Y=1.655 $X2=0.467 $Y2=2.095
cc_43 VPB N_A_c_89_n 0.0296577f $X=-0.19 $Y=1.655 $X2=0.467 $Y2=2.245
cc_44 VPB A 0.0364893f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_45 VPB N_A_c_84_n 0.00700725f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.74
cc_46 VPB N_B_M1004_g 0.0309034f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.755
cc_47 VPB N_B_M1007_g 0.0373138f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=0.83
cc_48 VPB N_B_c_159_n 0.0038376f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.755
cc_49 VPB N_B_c_166_n 0.0143144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB B 0.0122887f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.575
cc_51 VPB N_B_c_162_n 0.0501761f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.385
cc_52 VPB N_A_143_487#_M1008_g 0.0226974f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=0.515
cc_53 VPB N_A_143_487#_c_238_n 0.0224888f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=0.98
cc_54 VPB N_A_143_487#_c_234_n 0.00420373f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=0.905
cc_55 VPB N_A_143_487#_c_240_n 0.0142644f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.515
cc_56 VPB N_A_143_487#_c_241_n 0.0125999f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.385
cc_57 VPB N_A_143_487#_c_235_n 0.0368889f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_58 VPB N_A_143_487#_c_243_n 0.00516886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_143_487#_c_244_n 0.00566703f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=0.35
cc_60 VPB N_VPWR_c_315_n 0.0154735f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=0.83
cc_61 VPB N_VPWR_c_316_n 0.0307707f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=0.905
cc_62 VPB N_VPWR_c_317_n 0.0155083f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=0.51
cc_63 VPB N_VPWR_c_318_n 0.00460443f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.755
cc_64 VPB N_VPWR_c_319_n 0.0198782f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.095
cc_65 VPB N_VPWR_c_320_n 0.0109393f $X=-0.19 $Y=1.655 $X2=0.467 $Y2=2.245
cc_66 VPB N_VPWR_c_321_n 0.0267876f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=0.905
cc_67 VPB N_VPWR_c_322_n 0.00555175f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.515
cc_68 VPB N_VPWR_c_314_n 0.0675921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_324_n 0.0110305f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=0.35
cc_70 VPB N_Y_c_359_n 0.0176741f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.905
cc_71 VPB N_Y_c_360_n 0.00245069f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=0.905
cc_72 VPB N_Y_c_356_n 0.035368f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=0.83
cc_73 N_A_M1006_g N_B_c_157_n 0.0486639f $X=0.475 $Y=1.095 $X2=-0.19 $Y2=-0.245
cc_74 N_A_c_74_n N_B_c_157_n 0.00662657f $X=1.325 $Y=0.83 $X2=-0.19 $Y2=-0.245
cc_75 N_A_c_80_n N_B_c_157_n 0.00515877f $X=0.63 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_76 N_A_c_82_n N_B_c_157_n 0.00570962f $X=1.175 $Y=0.35 $X2=-0.19 $Y2=-0.245
cc_77 N_A_M1005_g N_B_M1004_g 0.0121323f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_78 N_A_c_89_n N_B_M1004_g 0.020633f $X=0.467 $Y=2.245 $X2=0 $Y2=0
cc_79 N_A_c_77_n N_B_M1009_g 0.0299823f $X=1.84 $Y=0.83 $X2=0 $Y2=0
cc_80 N_A_c_75_n B 0.00146537f $X=1.765 $Y=0.905 $X2=0 $Y2=0
cc_81 N_A_c_76_n B 0.00137233f $X=1.4 $Y=0.905 $X2=0 $Y2=0
cc_82 N_A_M1005_g B 0.0328595f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_83 N_A_M1005_g N_B_c_161_n 0.121873f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_84 N_A_c_76_n N_B_c_162_n 0.00855299f $X=1.4 $Y=0.905 $X2=0 $Y2=0
cc_85 N_A_M1005_g N_B_c_162_n 0.0423731f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_86 A N_B_c_162_n 0.00298259f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_87 N_A_c_84_n N_B_c_162_n 0.0122857f $X=0.385 $Y=1.74 $X2=0 $Y2=0
cc_88 N_A_M1005_g N_A_143_487#_c_234_n 0.00174409f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_89 N_A_c_89_n N_A_143_487#_c_234_n 0.00169761f $X=0.467 $Y=2.245 $X2=0 $Y2=0
cc_90 A N_A_143_487#_c_234_n 0.0641201f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_91 N_A_c_84_n N_A_143_487#_c_234_n 0.00131823f $X=0.385 $Y=1.74 $X2=0 $Y2=0
cc_92 N_A_M1005_g N_A_143_487#_c_240_n 0.0149773f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_93 N_A_M1000_g N_A_143_487#_c_243_n 0.00509387f $X=0.64 $Y=2.755 $X2=0 $Y2=0
cc_94 N_A_M1006_g N_A_143_487#_c_236_n 4.96905e-19 $X=0.475 $Y=1.095 $X2=0 $Y2=0
cc_95 N_A_c_76_n N_A_143_487#_c_236_n 6.39892e-19 $X=1.4 $Y=0.905 $X2=0 $Y2=0
cc_96 N_A_M1005_g N_A_143_487#_c_236_n 0.00504967f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_97 N_A_c_80_n N_A_143_487#_c_236_n 0.0230135f $X=0.63 $Y=1.43 $X2=0 $Y2=0
cc_98 N_A_c_82_n N_A_143_487#_c_236_n 0.0123447f $X=1.175 $Y=0.35 $X2=0 $Y2=0
cc_99 N_A_c_85_n N_A_143_487#_c_236_n 0.00400941f $X=1.325 $Y=0.35 $X2=0 $Y2=0
cc_100 N_A_M1005_g N_A_143_487#_c_244_n 0.00487833f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_101 N_A_M1000_g N_VPWR_c_316_n 0.0105077f $X=0.64 $Y=2.755 $X2=0 $Y2=0
cc_102 N_A_c_89_n N_VPWR_c_316_n 0.00238144f $X=0.467 $Y=2.245 $X2=0 $Y2=0
cc_103 A N_VPWR_c_316_n 0.0274416f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_104 N_A_M1000_g N_VPWR_c_317_n 0.00544562f $X=0.64 $Y=2.755 $X2=0 $Y2=0
cc_105 N_A_M1005_g N_VPWR_c_318_n 0.0159513f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_106 N_A_M1005_g N_VPWR_c_321_n 0.00469214f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_107 N_A_M1000_g N_VPWR_c_314_n 0.00951556f $X=0.64 $Y=2.755 $X2=0 $Y2=0
cc_108 N_A_M1005_g N_VPWR_c_314_n 0.00810928f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_109 N_A_M1005_g N_Y_c_362_n 0.00124905f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_110 N_A_M1005_g N_Y_c_360_n 6.69631e-19 $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_111 N_A_M1006_g N_VGND_c_398_n 0.00329965f $X=0.475 $Y=1.095 $X2=0 $Y2=0
cc_112 N_A_c_80_n N_VGND_c_398_n 0.0410951f $X=0.63 $Y=1.43 $X2=0 $Y2=0
cc_113 N_A_c_81_n N_VGND_c_398_n 0.022733f $X=0.715 $Y=0.385 $X2=0 $Y2=0
cc_114 A N_VGND_c_398_n 0.0242278f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_115 N_A_c_84_n N_VGND_c_398_n 7.79026e-19 $X=0.385 $Y=1.74 $X2=0 $Y2=0
cc_116 N_A_c_85_n N_VGND_c_398_n 0.00179084f $X=1.325 $Y=0.35 $X2=0 $Y2=0
cc_117 N_A_c_77_n N_VGND_c_399_n 0.00271771f $X=1.84 $Y=0.83 $X2=0 $Y2=0
cc_118 N_A_c_82_n N_VGND_c_399_n 0.00206613f $X=1.175 $Y=0.35 $X2=0 $Y2=0
cc_119 N_A_M1006_g N_VGND_c_400_n 0.00292802f $X=0.475 $Y=1.095 $X2=0 $Y2=0
cc_120 N_A_c_77_n N_VGND_c_400_n 0.00522039f $X=1.84 $Y=0.83 $X2=0 $Y2=0
cc_121 N_A_c_81_n N_VGND_c_400_n 0.0121867f $X=0.715 $Y=0.385 $X2=0 $Y2=0
cc_122 N_A_c_82_n N_VGND_c_400_n 0.0404267f $X=1.175 $Y=0.35 $X2=0 $Y2=0
cc_123 N_A_c_85_n N_VGND_c_400_n 0.00840857f $X=1.325 $Y=0.35 $X2=0 $Y2=0
cc_124 N_A_M1006_g N_VGND_c_402_n 0.0039117f $X=0.475 $Y=1.095 $X2=0 $Y2=0
cc_125 N_A_c_75_n N_VGND_c_402_n 4.30519e-19 $X=1.765 $Y=0.905 $X2=0 $Y2=0
cc_126 N_A_c_77_n N_VGND_c_402_n 0.00584136f $X=1.84 $Y=0.83 $X2=0 $Y2=0
cc_127 N_A_c_81_n N_VGND_c_402_n 0.00660921f $X=0.715 $Y=0.385 $X2=0 $Y2=0
cc_128 N_A_c_82_n N_VGND_c_402_n 0.0222082f $X=1.175 $Y=0.35 $X2=0 $Y2=0
cc_129 N_A_c_85_n N_VGND_c_402_n 0.0132523f $X=1.325 $Y=0.35 $X2=0 $Y2=0
cc_130 N_A_c_75_n N_A_300_60#_c_436_n 0.00450001f $X=1.765 $Y=0.905 $X2=0 $Y2=0
cc_131 N_A_c_77_n N_A_300_60#_c_436_n 0.00176547f $X=1.84 $Y=0.83 $X2=0 $Y2=0
cc_132 N_A_c_82_n N_A_300_60#_c_436_n 0.01363f $X=1.175 $Y=0.35 $X2=0 $Y2=0
cc_133 N_A_c_85_n N_A_300_60#_c_436_n 0.00930062f $X=1.325 $Y=0.35 $X2=0 $Y2=0
cc_134 N_A_c_75_n N_A_300_60#_c_437_n 4.17754e-19 $X=1.765 $Y=0.905 $X2=0 $Y2=0
cc_135 N_A_M1005_g N_A_300_60#_c_437_n 0.00454396f $X=1.84 $Y=2.755 $X2=0 $Y2=0
cc_136 N_A_c_79_n N_A_300_60#_c_437_n 0.00705259f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_137 N_A_c_75_n N_A_300_60#_c_438_n 0.00902957f $X=1.765 $Y=0.905 $X2=0 $Y2=0
cc_138 N_B_M1007_g N_A_143_487#_c_238_n 0.0190484f $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_139 N_B_M1009_g N_A_143_487#_c_232_n 0.0176362f $X=2.27 $Y=0.51 $X2=0 $Y2=0
cc_140 N_B_c_157_n N_A_143_487#_c_234_n 0.0041379f $X=0.835 $Y=1.425 $X2=0 $Y2=0
cc_141 N_B_M1004_g N_A_143_487#_c_234_n 0.00617077f $X=1.07 $Y=2.755 $X2=0 $Y2=0
cc_142 B N_A_143_487#_c_234_n 0.0558044f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_143 N_B_c_162_n N_A_143_487#_c_234_n 0.0325996f $X=1.07 $Y=1.76 $X2=0 $Y2=0
cc_144 N_B_M1004_g N_A_143_487#_c_240_n 0.00527632f $X=1.07 $Y=2.755 $X2=0 $Y2=0
cc_145 B N_A_143_487#_c_240_n 0.0376148f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_146 N_B_c_162_n N_A_143_487#_c_240_n 0.00831901f $X=1.07 $Y=1.76 $X2=0 $Y2=0
cc_147 N_B_M1007_g N_A_143_487#_c_241_n 0.0134887f $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_148 N_B_c_166_n N_A_143_487#_c_241_n 0.00123455f $X=2.29 $Y=1.89 $X2=0 $Y2=0
cc_149 B N_A_143_487#_c_241_n 0.0287202f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_B_M1007_g N_A_143_487#_c_270_n 9.84104e-19 $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_151 N_B_c_159_n N_A_143_487#_c_270_n 4.12227e-19 $X=2.29 $Y=1.725 $X2=0 $Y2=0
cc_152 B N_A_143_487#_c_270_n 0.0214283f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_153 N_B_M1007_g N_A_143_487#_c_235_n 0.00763521f $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_154 N_B_M1009_g N_A_143_487#_c_235_n 0.00955303f $X=2.27 $Y=0.51 $X2=0 $Y2=0
cc_155 B N_A_143_487#_c_235_n 0.0026068f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_156 N_B_c_161_n N_A_143_487#_c_235_n 0.0408791f $X=2.29 $Y=1.385 $X2=0 $Y2=0
cc_157 N_B_M1004_g N_A_143_487#_c_243_n 0.0103648f $X=1.07 $Y=2.755 $X2=0 $Y2=0
cc_158 N_B_c_162_n N_A_143_487#_c_243_n 0.00354294f $X=1.07 $Y=1.76 $X2=0 $Y2=0
cc_159 N_B_c_157_n N_A_143_487#_c_236_n 0.00365601f $X=0.835 $Y=1.425 $X2=0
+ $Y2=0
cc_160 B N_A_143_487#_c_236_n 0.00202474f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_161 N_B_c_162_n N_A_143_487#_c_236_n 0.00394938f $X=1.07 $Y=1.76 $X2=0 $Y2=0
cc_162 N_B_M1007_g N_A_143_487#_c_244_n 0.00463967f $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_163 B N_A_143_487#_c_244_n 0.0164344f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_164 N_B_M1004_g N_VPWR_c_316_n 6.10799e-19 $X=1.07 $Y=2.755 $X2=0 $Y2=0
cc_165 N_B_M1004_g N_VPWR_c_317_n 0.00565115f $X=1.07 $Y=2.755 $X2=0 $Y2=0
cc_166 N_B_M1004_g N_VPWR_c_318_n 0.00315148f $X=1.07 $Y=2.755 $X2=0 $Y2=0
cc_167 N_B_M1007_g N_VPWR_c_318_n 0.00251318f $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_168 N_B_M1007_g N_VPWR_c_321_n 0.00559492f $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_169 N_B_M1004_g N_VPWR_c_314_n 0.0111464f $X=1.07 $Y=2.755 $X2=0 $Y2=0
cc_170 N_B_M1007_g N_VPWR_c_314_n 0.0104996f $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_171 N_B_M1007_g N_Y_c_362_n 0.0067136f $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_172 N_B_M1007_g N_Y_c_360_n 0.00302297f $X=2.2 $Y=2.755 $X2=0 $Y2=0
cc_173 B N_Y_c_356_n 0.00522175f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_174 B Y 0.0084821f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_175 N_B_M1009_g N_Y_c_358_n 0.00123474f $X=2.27 $Y=0.51 $X2=0 $Y2=0
cc_176 N_B_M1009_g N_VGND_c_399_n 0.00325556f $X=2.27 $Y=0.51 $X2=0 $Y2=0
cc_177 N_B_M1009_g N_VGND_c_401_n 0.00522039f $X=2.27 $Y=0.51 $X2=0 $Y2=0
cc_178 N_B_M1009_g N_VGND_c_402_n 0.00562511f $X=2.27 $Y=0.51 $X2=0 $Y2=0
cc_179 N_B_M1009_g N_A_300_60#_c_437_n 0.0123545f $X=2.27 $Y=0.51 $X2=0 $Y2=0
cc_180 B N_A_300_60#_c_437_n 0.0534965f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_181 N_B_c_161_n N_A_300_60#_c_437_n 0.00132478f $X=2.29 $Y=1.385 $X2=0 $Y2=0
cc_182 N_B_c_157_n N_A_300_60#_c_438_n 2.63194e-19 $X=0.835 $Y=1.425 $X2=0 $Y2=0
cc_183 B N_A_300_60#_c_438_n 0.0183398f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_184 N_B_c_162_n N_A_300_60#_c_438_n 2.2172e-19 $X=1.07 $Y=1.76 $X2=0 $Y2=0
cc_185 N_B_M1009_g N_A_300_60#_c_439_n 0.00182871f $X=2.27 $Y=0.51 $X2=0 $Y2=0
cc_186 N_A_143_487#_c_243_n N_VPWR_c_316_n 0.00163258f $X=0.932 $Y=2.35 $X2=0
+ $Y2=0
cc_187 N_A_143_487#_c_285_p N_VPWR_c_317_n 0.0137139f $X=0.855 $Y=2.56 $X2=0
+ $Y2=0
cc_188 N_A_143_487#_c_240_n N_VPWR_c_318_n 0.0473322f $X=1.93 $Y=2.35 $X2=0
+ $Y2=0
cc_189 N_A_143_487#_M1008_g N_VPWR_c_319_n 0.00458904f $X=2.65 $Y=2.755 $X2=0
+ $Y2=0
cc_190 N_A_143_487#_M1008_g N_VPWR_c_321_n 0.00414311f $X=2.65 $Y=2.755 $X2=0
+ $Y2=0
cc_191 N_A_143_487#_M1008_g N_VPWR_c_314_n 0.00687257f $X=2.65 $Y=2.755 $X2=0
+ $Y2=0
cc_192 N_A_143_487#_c_285_p N_VPWR_c_314_n 0.0095959f $X=0.855 $Y=2.56 $X2=0
+ $Y2=0
cc_193 N_A_143_487#_c_244_n A_383_487# 0.00704584f $X=2.015 $Y=2.15 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_143_487#_M1008_g N_Y_c_362_n 0.0105461f $X=2.65 $Y=2.755 $X2=0 $Y2=0
cc_195 N_A_143_487#_M1008_g N_Y_c_359_n 0.0107211f $X=2.65 $Y=2.755 $X2=0 $Y2=0
cc_196 N_A_143_487#_c_238_n N_Y_c_359_n 0.00874248f $X=2.787 $Y=2.28 $X2=0 $Y2=0
cc_197 N_A_143_487#_c_241_n N_Y_c_359_n 0.0252238f $X=2.67 $Y=2.15 $X2=0 $Y2=0
cc_198 N_A_143_487#_M1008_g N_Y_c_360_n 0.00109181f $X=2.65 $Y=2.755 $X2=0 $Y2=0
cc_199 N_A_143_487#_c_241_n N_Y_c_360_n 0.0274138f $X=2.67 $Y=2.15 $X2=0 $Y2=0
cc_200 N_A_143_487#_c_244_n N_Y_c_360_n 0.00239713f $X=2.015 $Y=2.15 $X2=0 $Y2=0
cc_201 N_A_143_487#_M1008_g N_Y_c_356_n 0.00341538f $X=2.65 $Y=2.755 $X2=0 $Y2=0
cc_202 N_A_143_487#_c_241_n N_Y_c_356_n 0.0135424f $X=2.67 $Y=2.15 $X2=0 $Y2=0
cc_203 N_A_143_487#_c_270_n N_Y_c_356_n 0.0368657f $X=2.835 $Y=1.73 $X2=0 $Y2=0
cc_204 N_A_143_487#_c_235_n N_Y_c_356_n 0.0237967f $X=2.835 $Y=1.73 $X2=0 $Y2=0
cc_205 N_A_143_487#_c_270_n Y 0.0140534f $X=2.835 $Y=1.73 $X2=0 $Y2=0
cc_206 N_A_143_487#_c_235_n Y 0.0207439f $X=2.835 $Y=1.73 $X2=0 $Y2=0
cc_207 N_A_143_487#_c_232_n N_Y_c_358_n 0.00794661f $X=2.812 $Y=0.83 $X2=0 $Y2=0
cc_208 N_A_143_487#_c_233_n N_Y_c_358_n 0.0126779f $X=2.812 $Y=0.98 $X2=0 $Y2=0
cc_209 N_A_143_487#_c_235_n N_Y_c_358_n 0.00770982f $X=2.835 $Y=1.73 $X2=0 $Y2=0
cc_210 N_A_143_487#_c_232_n N_VGND_c_401_n 0.0049163f $X=2.812 $Y=0.83 $X2=0
+ $Y2=0
cc_211 N_A_143_487#_c_232_n N_VGND_c_402_n 0.0100091f $X=2.812 $Y=0.83 $X2=0
+ $Y2=0
cc_212 N_A_143_487#_c_233_n N_A_300_60#_c_437_n 0.00124872f $X=2.812 $Y=0.98
+ $X2=0 $Y2=0
cc_213 N_A_143_487#_c_235_n N_A_300_60#_c_437_n 4.8637e-19 $X=2.835 $Y=1.73
+ $X2=0 $Y2=0
cc_214 N_A_143_487#_c_236_n N_A_300_60#_c_438_n 0.00608607f $X=1.05 $Y=1.095
+ $X2=0 $Y2=0
cc_215 N_A_143_487#_c_232_n N_A_300_60#_c_439_n 9.86554e-19 $X=2.812 $Y=0.83
+ $X2=0 $Y2=0
cc_216 N_VPWR_c_318_n N_Y_c_362_n 0.0142493f $X=1.625 $Y=2.77 $X2=0 $Y2=0
cc_217 N_VPWR_c_321_n N_Y_c_362_n 0.014327f $X=2.77 $Y=3.33 $X2=0 $Y2=0
cc_218 N_VPWR_c_314_n N_Y_c_362_n 0.0122422f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_219 N_VPWR_M1008_d N_Y_c_359_n 0.00281787f $X=2.725 $Y=2.435 $X2=0 $Y2=0
cc_220 N_VPWR_c_319_n N_Y_c_359_n 0.0220376f $X=2.865 $Y=2.91 $X2=0 $Y2=0
cc_221 N_VPWR_c_320_n N_Y_c_359_n 0.00327508f $X=3.06 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_321_n N_Y_c_359_n 0.00187826f $X=2.77 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_c_314_n N_Y_c_359_n 0.0106656f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_224 N_Y_c_358_n N_VGND_c_401_n 0.0219794f $X=2.915 $Y=0.51 $X2=0 $Y2=0
cc_225 N_Y_c_358_n N_VGND_c_402_n 0.0190611f $X=2.915 $Y=0.51 $X2=0 $Y2=0
cc_226 N_Y_c_358_n N_A_300_60#_c_437_n 0.0164965f $X=2.915 $Y=0.51 $X2=0 $Y2=0
cc_227 N_Y_c_358_n N_A_300_60#_c_439_n 0.0249171f $X=2.915 $Y=0.51 $X2=0 $Y2=0
cc_228 N_VGND_c_400_n N_A_300_60#_c_436_n 0.0098153f $X=1.925 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_c_402_n N_A_300_60#_c_436_n 0.00900613f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_399_n N_A_300_60#_c_437_n 0.0167125f $X=2.055 $Y=0.51 $X2=0
+ $Y2=0
cc_231 N_VGND_c_402_n N_A_300_60#_c_437_n 0.0104618f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_401_n N_A_300_60#_c_439_n 0.00881347f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_402_n N_A_300_60#_c_439_n 0.0084502f $X=3.12 $Y=0 $X2=0 $Y2=0
