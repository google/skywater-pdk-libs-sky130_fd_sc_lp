* File: sky130_fd_sc_lp__o21ai_0.pxi.spice
* Created: Wed Sep  2 10:15:50 2020
* 
x_PM_SKY130_FD_SC_LP__O21AI_0%A1 N_A1_c_51_n N_A1_c_58_n N_A1_c_59_n
+ N_A1_M1002_g N_A1_c_60_n N_A1_M1003_g N_A1_c_53_n N_A1_c_54_n A1 A1 A1
+ N_A1_c_55_n N_A1_c_56_n PM_SKY130_FD_SC_LP__O21AI_0%A1
x_PM_SKY130_FD_SC_LP__O21AI_0%A2 N_A2_c_94_n N_A2_M1005_g N_A2_M1004_g
+ N_A2_c_100_n A2 A2 A2 N_A2_c_97_n PM_SKY130_FD_SC_LP__O21AI_0%A2
x_PM_SKY130_FD_SC_LP__O21AI_0%B1 N_B1_M1000_g N_B1_c_143_n N_B1_M1001_g
+ N_B1_c_145_n B1 B1 N_B1_c_141_n N_B1_c_142_n PM_SKY130_FD_SC_LP__O21AI_0%B1
x_PM_SKY130_FD_SC_LP__O21AI_0%VPWR N_VPWR_M1003_s N_VPWR_M1001_d N_VPWR_c_173_n
+ N_VPWR_c_174_n N_VPWR_c_175_n N_VPWR_c_176_n VPWR N_VPWR_c_177_n
+ N_VPWR_c_172_n PM_SKY130_FD_SC_LP__O21AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O21AI_0%Y N_Y_M1000_d N_Y_M1004_d N_Y_c_198_n N_Y_c_199_n
+ N_Y_c_200_n N_Y_c_201_n Y Y N_Y_c_204_n Y PM_SKY130_FD_SC_LP__O21AI_0%Y
x_PM_SKY130_FD_SC_LP__O21AI_0%A_39_47# N_A_39_47#_M1002_s N_A_39_47#_M1005_d
+ N_A_39_47#_c_235_n N_A_39_47#_c_236_n N_A_39_47#_c_237_n N_A_39_47#_c_238_n
+ PM_SKY130_FD_SC_LP__O21AI_0%A_39_47#
x_PM_SKY130_FD_SC_LP__O21AI_0%VGND N_VGND_M1002_d N_VGND_c_265_n VGND
+ N_VGND_c_266_n N_VGND_c_267_n N_VGND_c_268_n N_VGND_c_269_n
+ PM_SKY130_FD_SC_LP__O21AI_0%VGND
cc_1 VNB N_A1_c_51_n 0.00394182f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.155
cc_2 VNB N_A1_M1002_g 0.0248134f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.445
cc_3 VNB N_A1_c_53_n 0.0360149f $X=-0.19 $Y=-0.245 $X2=0.367 $Y2=1.005
cc_4 VNB N_A1_c_54_n 0.0207833f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.605
cc_5 VNB N_A1_c_55_n 0.0464259f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.1
cc_6 VNB N_A1_c_56_n 3.10515e-19 $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.1
cc_7 VNB N_A2_c_94_n 0.0158058f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.155
cc_8 VNB N_A2_M1005_g 0.0408348f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.855
cc_9 VNB A2 0.00628158f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.005
cc_10 VNB N_A2_c_97_n 0.0190451f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_11 VNB N_B1_M1000_g 0.0629793f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.23
cc_12 VNB N_B1_c_141_n 0.022889f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_13 VNB N_B1_c_142_n 0.0123442f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_VPWR_c_172_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_198_n 0.00626956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_199_n 0.0127268f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.305
cc_17 VNB N_Y_c_200_n 0.00318978f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.735
cc_18 VNB N_Y_c_201_n 0.0390672f $X=-0.19 $Y=-0.245 $X2=0.367 $Y2=0.855
cc_19 VNB N_A_39_47#_c_235_n 0.0153392f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.305
cc_20 VNB N_A_39_47#_c_236_n 0.0116793f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.735
cc_21 VNB N_A_39_47#_c_237_n 0.00917553f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.005
cc_22 VNB N_A_39_47#_c_238_n 3.26325e-19 $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.44
cc_23 VNB N_VGND_c_265_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.445
cc_24 VNB N_VGND_c_266_n 0.0166947f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.735
cc_25 VNB N_VGND_c_267_n 0.0277357f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_26 VNB N_VGND_c_268_n 0.13243f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_27 VNB N_VGND_c_269_n 0.0043639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A1_c_51_n 0.0415925f $X=-0.19 $Y=1.655 $X2=0.2 $Y2=2.155
cc_29 VPB N_A1_c_58_n 0.0276347f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.23
cc_30 VPB N_A1_c_59_n 0.0163313f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=2.23
cc_31 VPB N_A1_c_60_n 0.0208199f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.305
cc_32 VPB N_A1_c_56_n 0.00428927f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.1
cc_33 VPB N_A2_c_94_n 0.00562302f $X=-0.19 $Y=1.655 $X2=0.2 $Y2=2.155
cc_34 VPB N_A2_M1004_g 0.0377417f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.305
cc_35 VPB N_A2_c_100_n 0.0203371f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.735
cc_36 VPB A2 0.0132147f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.005
cc_37 VPB N_B1_c_143_n 0.0254125f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.445
cc_38 VPB N_B1_M1001_g 0.0339983f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.305
cc_39 VPB N_B1_c_145_n 0.0233302f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.735
cc_40 VPB N_B1_c_141_n 4.4119e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_41 VPB N_B1_c_142_n 0.0255856f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_42 VPB N_VPWR_c_173_n 0.0138329f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.445
cc_43 VPB N_VPWR_c_174_n 0.0327068f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.305
cc_44 VPB N_VPWR_c_175_n 0.0119904f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.735
cc_45 VPB N_VPWR_c_176_n 0.0346192f $X=-0.19 $Y=1.655 $X2=0.367 $Y2=0.855
cc_46 VPB N_VPWR_c_177_n 0.0271245f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_47 VPB N_VPWR_c_172_n 0.062488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_Y_c_198_n 0.0110911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB Y 0.00203831f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.44
cc_50 VPB N_Y_c_204_n 0.00485884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 N_A1_c_51_n N_A2_c_94_n 0.00874958f $X=0.2 $Y=2.155 $X2=0 $Y2=0
cc_52 N_A1_c_54_n N_A2_c_94_n 0.0108965f $X=0.29 $Y=1.605 $X2=0 $Y2=0
cc_53 N_A1_c_56_n N_A2_c_94_n 0.0010601f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_54 N_A1_M1002_g N_A2_M1005_g 0.0252811f $X=0.535 $Y=0.445 $X2=0 $Y2=0
cc_55 N_A1_c_55_n N_A2_M1005_g 0.00620083f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_56 N_A1_c_56_n N_A2_M1005_g 6.03808e-19 $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_57 N_A1_c_51_n N_A2_M1004_g 0.00348165f $X=0.2 $Y=2.155 $X2=0 $Y2=0
cc_58 N_A1_c_58_n N_A2_M1004_g 0.0531675f $X=0.5 $Y=2.23 $X2=0 $Y2=0
cc_59 N_A1_c_56_n N_A2_M1004_g 4.89102e-19 $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_60 N_A1_c_51_n A2 0.00134602f $X=0.2 $Y=2.155 $X2=0 $Y2=0
cc_61 N_A1_c_58_n A2 0.0013458f $X=0.5 $Y=2.23 $X2=0 $Y2=0
cc_62 N_A1_c_55_n A2 0.00323719f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_63 N_A1_c_56_n A2 0.0820913f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_64 N_A1_c_55_n N_A2_c_97_n 0.0108965f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_65 N_A1_c_56_n N_A2_c_97_n 4.10574e-19 $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_66 N_A1_c_59_n N_VPWR_c_174_n 0.00883951f $X=0.275 $Y=2.23 $X2=0 $Y2=0
cc_67 N_A1_c_60_n N_VPWR_c_174_n 0.0181618f $X=0.575 $Y=2.305 $X2=0 $Y2=0
cc_68 N_A1_c_56_n N_VPWR_c_174_n 0.0168461f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_69 N_A1_c_60_n N_VPWR_c_177_n 0.00452967f $X=0.575 $Y=2.305 $X2=0 $Y2=0
cc_70 N_A1_c_60_n N_VPWR_c_172_n 0.00809218f $X=0.575 $Y=2.305 $X2=0 $Y2=0
cc_71 N_A1_c_60_n Y 0.00168372f $X=0.575 $Y=2.305 $X2=0 $Y2=0
cc_72 N_A1_c_60_n N_Y_c_204_n 6.13655e-19 $X=0.575 $Y=2.305 $X2=0 $Y2=0
cc_73 N_A1_M1002_g N_A_39_47#_c_235_n 8.56298e-19 $X=0.535 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A1_M1002_g N_A_39_47#_c_236_n 0.0168305f $X=0.535 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A1_c_53_n N_A_39_47#_c_236_n 0.00149195f $X=0.367 $Y=1.005 $X2=0 $Y2=0
cc_76 N_A1_c_56_n N_A_39_47#_c_236_n 0.00307848f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_77 N_A1_c_53_n N_A_39_47#_c_237_n 0.00853498f $X=0.367 $Y=1.005 $X2=0 $Y2=0
cc_78 N_A1_c_56_n N_A_39_47#_c_237_n 0.0228447f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_79 N_A1_M1002_g N_VGND_c_265_n 0.00920213f $X=0.535 $Y=0.445 $X2=0 $Y2=0
cc_80 N_A1_M1002_g N_VGND_c_266_n 0.00358332f $X=0.535 $Y=0.445 $X2=0 $Y2=0
cc_81 N_A1_M1002_g N_VGND_c_268_n 0.00533413f $X=0.535 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A1_c_53_n N_VGND_c_268_n 7.84805e-19 $X=0.367 $Y=1.005 $X2=0 $Y2=0
cc_83 N_A2_M1005_g N_B1_M1000_g 0.0171395f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_84 A2 N_B1_M1000_g 4.44047e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A2_c_94_n N_B1_c_143_n 0.0171395f $X=0.855 $Y=1.73 $X2=0 $Y2=0
cc_86 N_A2_M1004_g N_B1_M1001_g 0.0171395f $X=0.965 $Y=2.735 $X2=0 $Y2=0
cc_87 N_A2_c_100_n N_B1_c_145_n 0.0171395f $X=0.855 $Y=1.915 $X2=0 $Y2=0
cc_88 N_A2_c_97_n N_B1_c_141_n 0.0171395f $X=0.835 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A2_M1004_g N_VPWR_c_174_n 0.00278661f $X=0.965 $Y=2.735 $X2=0 $Y2=0
cc_90 N_A2_M1004_g N_VPWR_c_177_n 0.00511358f $X=0.965 $Y=2.735 $X2=0 $Y2=0
cc_91 N_A2_M1004_g N_VPWR_c_172_n 0.00961121f $X=0.965 $Y=2.735 $X2=0 $Y2=0
cc_92 A2 N_Y_c_198_n 0.0590924f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A2_c_97_n N_Y_c_198_n 0.0102144f $X=0.835 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A2_M1005_g N_Y_c_200_n 0.00142265f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_95 A2 N_Y_c_200_n 0.0135822f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_96 A2 N_Y_c_201_n 6.01403e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A2_M1004_g Y 0.010254f $X=0.965 $Y=2.735 $X2=0 $Y2=0
cc_98 N_A2_M1004_g N_Y_c_204_n 0.00615898f $X=0.965 $Y=2.735 $X2=0 $Y2=0
cc_99 N_A2_M1005_g N_A_39_47#_c_236_n 0.015461f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_100 A2 N_A_39_47#_c_236_n 0.018383f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A2_c_97_n N_A_39_47#_c_236_n 0.00104593f $X=0.835 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A2_M1005_g N_A_39_47#_c_238_n 3.24738e-19 $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_103 N_A2_M1005_g N_VGND_c_265_n 0.00820137f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A2_M1005_g N_VGND_c_267_n 0.00358332f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A2_M1005_g N_VGND_c_268_n 0.00430105f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_106 N_B1_M1001_g N_VPWR_c_176_n 0.00486495f $X=1.395 $Y=2.735 $X2=0 $Y2=0
cc_107 N_B1_c_145_n N_VPWR_c_176_n 0.0014227f $X=1.51 $Y=2.14 $X2=0 $Y2=0
cc_108 N_B1_c_142_n N_VPWR_c_176_n 0.0194068f $X=1.535 $Y=1.635 $X2=0 $Y2=0
cc_109 N_B1_M1001_g N_VPWR_c_177_n 0.00525604f $X=1.395 $Y=2.735 $X2=0 $Y2=0
cc_110 N_B1_M1001_g N_VPWR_c_172_n 0.0106161f $X=1.395 $Y=2.735 $X2=0 $Y2=0
cc_111 N_B1_M1000_g N_Y_c_198_n 0.0129635f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_112 N_B1_c_142_n N_Y_c_198_n 0.0494154f $X=1.535 $Y=1.635 $X2=0 $Y2=0
cc_113 N_B1_M1000_g N_Y_c_199_n 0.0199704f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_114 N_B1_c_141_n N_Y_c_199_n 0.00176764f $X=1.535 $Y=1.635 $X2=0 $Y2=0
cc_115 N_B1_c_142_n N_Y_c_199_n 0.0275488f $X=1.535 $Y=1.635 $X2=0 $Y2=0
cc_116 N_B1_M1000_g N_Y_c_201_n 0.016238f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_117 N_B1_M1001_g Y 0.00624832f $X=1.395 $Y=2.735 $X2=0 $Y2=0
cc_118 N_B1_M1001_g N_Y_c_204_n 0.00792625f $X=1.395 $Y=2.735 $X2=0 $Y2=0
cc_119 N_B1_M1000_g N_A_39_47#_c_236_n 0.00154364f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_120 N_B1_M1000_g N_A_39_47#_c_238_n 2.26018e-19 $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_121 N_B1_M1000_g N_VGND_c_265_n 0.00124917f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_122 N_B1_M1000_g N_VGND_c_267_n 0.00585385f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B1_M1000_g N_VGND_c_268_n 0.0120598f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_124 N_VPWR_c_174_n Y 0.0187899f $X=0.36 $Y=2.56 $X2=0 $Y2=0
cc_125 N_VPWR_c_176_n Y 0.0229504f $X=1.61 $Y=2.56 $X2=0 $Y2=0
cc_126 N_VPWR_c_177_n Y 0.0226628f $X=1.505 $Y=3.33 $X2=0 $Y2=0
cc_127 N_VPWR_c_172_n Y 0.0121892f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_128 N_VPWR_c_174_n N_Y_c_204_n 0.00269259f $X=0.36 $Y=2.56 $X2=0 $Y2=0
cc_129 N_VPWR_c_176_n N_Y_c_204_n 0.00396258f $X=1.61 $Y=2.56 $X2=0 $Y2=0
cc_130 N_Y_c_199_n N_A_39_47#_c_236_n 0.00294647f $X=1.49 $Y=1.205 $X2=0 $Y2=0
cc_131 N_Y_c_200_n N_A_39_47#_c_236_n 0.0112096f $X=1.27 $Y=1.205 $X2=0 $Y2=0
cc_132 N_Y_c_201_n N_A_39_47#_c_236_n 0.0141076f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_133 N_Y_c_201_n N_A_39_47#_c_238_n 0.0157113f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_134 N_Y_c_201_n N_VGND_c_267_n 0.0161226f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_135 N_Y_M1000_d N_VGND_c_268_n 0.00289872f $X=1.47 $Y=0.235 $X2=0 $Y2=0
cc_136 N_Y_c_201_n N_VGND_c_268_n 0.0108688f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A_39_47#_c_236_n N_VGND_c_265_n 0.02032f $X=1.085 $Y=0.76 $X2=0 $Y2=0
cc_138 N_A_39_47#_c_235_n N_VGND_c_266_n 0.0151488f $X=0.32 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A_39_47#_c_236_n N_VGND_c_266_n 0.00260179f $X=1.085 $Y=0.76 $X2=0
+ $Y2=0
cc_140 N_A_39_47#_c_236_n N_VGND_c_267_n 0.00260179f $X=1.085 $Y=0.76 $X2=0
+ $Y2=0
cc_141 N_A_39_47#_c_238_n N_VGND_c_267_n 0.011992f $X=1.18 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_39_47#_M1002_s N_VGND_c_268_n 0.00234689f $X=0.195 $Y=0.235 $X2=0
+ $Y2=0
cc_143 N_A_39_47#_M1005_d N_VGND_c_268_n 0.00243138f $X=1.04 $Y=0.235 $X2=0
+ $Y2=0
cc_144 N_A_39_47#_c_235_n N_VGND_c_268_n 0.00985676f $X=0.32 $Y=0.445 $X2=0
+ $Y2=0
cc_145 N_A_39_47#_c_236_n N_VGND_c_268_n 0.00957128f $X=1.085 $Y=0.76 $X2=0
+ $Y2=0
cc_146 N_A_39_47#_c_238_n N_VGND_c_268_n 0.00890164f $X=1.18 $Y=0.445 $X2=0
+ $Y2=0
