* File: sky130_fd_sc_lp__a221oi_lp.spice
* Created: Fri Aug 28 09:53:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a221oi_lp.pex.spice"
.subckt sky130_fd_sc_lp__a221oi_lp  VNB VPB B2 B1 A1 A2 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1008 A_155_48# N_B2_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.7
+ A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1009_d N_B1_M1009_g A_155_48# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0504 PD=0.81 PS=0.66 NRD=31.428 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1001 A_341_48# N_A1_M1001_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g A_341_48# VNB NSHORT L=0.15 W=0.42 AD=0.147
+ AS=0.0504 PD=1.12 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1006 A_589_48# N_C1_M1006_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.147 PD=0.63 PS=1.12 NRD=14.28 NRS=120 M=1 R=2.8 SA=75002.4 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g A_589_48# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_163_412#_M1010_d N_B2_M1010_g N_A_56_412#_M1010_s VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_163_412#_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=1.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1002 N_A_163_412#_M1002_d N_A2_M1002_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=1.57 NRD=0 NRS=57.13 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1007 N_A_56_412#_M1007_d N_B1_M1007_g N_A_163_412#_M1002_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1004 N_Y_M1004_d N_C1_M1004_g N_A_56_412#_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX11_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a221oi_lp.pxi.spice"
*
.ends
*
*
