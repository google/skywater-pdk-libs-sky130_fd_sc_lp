* File: sky130_fd_sc_lp__and2b_2.pex.spice
* Created: Fri Aug 28 10:05:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2B_2%A_N 3 7 8 9 13 15
c29 13 0 1.94138e-19 $X=0.525 $Y=1.375
c30 8 0 3.93152e-20 $X=0.72 $Y=1.295
r31 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.375
+ $X2=0.525 $Y2=1.54
r32 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.375
+ $X2=0.525 $Y2=1.21
r33 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.375 $X2=0.525 $Y2=1.375
r34 9 14 7.22631 $w=4.78e-07 $l=2.9e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.375
r35 8 14 1.99346 $w=4.78e-07 $l=8e-08 $layer=LI1_cond $X=0.68 $Y=1.295 $X2=0.68
+ $Y2=1.375
r36 7 15 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.59 $Y=0.875
+ $X2=0.59 $Y2=1.21
r37 3 16 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.48 $Y=2.045
+ $X2=0.48 $Y2=1.54
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_2%A_186_239# 1 2 9 11 13 16 20 24 25 27 28 31
+ 33 36 37 41
c84 33 0 1.62043e-19 $X=2.905 $Y=1.71
c85 11 0 3.93152e-20 $X=1.18 $Y=1.195
r86 44 45 41.8061 $w=2.94e-07 $l=2.55e-07 $layer=POLY_cond $X=1.18 $Y=1.435
+ $X2=1.435 $Y2=1.435
r87 39 41 9.71075 $w=3.03e-07 $l=2.57e-07 $layer=LI1_cond $X=2.775 $Y=0.877
+ $X2=3.032 $Y2=0.877
r88 35 41 1.80741 $w=2.55e-07 $l=1.53e-07 $layer=LI1_cond $X=3.032 $Y=1.03
+ $X2=3.032 $Y2=0.877
r89 35 36 26.8903 $w=2.53e-07 $l=5.95e-07 $layer=LI1_cond $X=3.032 $Y=1.03
+ $X2=3.032 $Y2=1.625
r90 34 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.44 $Y=1.71
+ $X2=2.345 $Y2=1.71
r91 33 36 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=2.905 $Y=1.71
+ $X2=3.032 $Y2=1.625
r92 33 34 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.905 $Y=1.71
+ $X2=2.44 $Y2=1.71
r93 29 37 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=1.795
+ $X2=2.345 $Y2=1.71
r94 29 31 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=2.345 $Y=1.795
+ $X2=2.345 $Y2=2.045
r95 27 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.25 $Y=1.71
+ $X2=2.345 $Y2=1.71
r96 27 28 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.25 $Y=1.71
+ $X2=1.735 $Y2=1.71
r97 25 45 22.1327 $w=2.94e-07 $l=1.35e-07 $layer=POLY_cond $X=1.57 $Y=1.435
+ $X2=1.435 $Y2=1.435
r98 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.51 $X2=1.57 $Y2=1.51
r99 22 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.61 $Y=1.625
+ $X2=1.735 $Y2=1.71
r100 22 24 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=1.61 $Y=1.625
+ $X2=1.61 $Y2=1.51
r101 18 25 6.55782 $w=2.94e-07 $l=4e-08 $layer=POLY_cond $X=1.61 $Y=1.435
+ $X2=1.57 $Y2=1.435
r102 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.61 $Y=1.345
+ $X2=1.61 $Y2=0.665
r103 14 45 18.4939 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.435 $Y=1.675
+ $X2=1.435 $Y2=1.435
r104 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.435 $Y=1.675
+ $X2=1.435 $Y2=2.465
r105 11 44 18.4939 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.18 $Y=1.195
+ $X2=1.18 $Y2=1.435
r106 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.18 $Y=1.195
+ $X2=1.18 $Y2=0.665
r107 7 44 28.6905 $w=2.94e-07 $l=1.75e-07 $layer=POLY_cond $X=1.005 $Y=1.435
+ $X2=1.18 $Y2=1.435
r108 7 9 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=1.005 $Y=1.495
+ $X2=1.005 $Y2=2.465
r109 2 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.205
+ $Y=1.835 $X2=2.345 $Y2=2.045
r110 1 39 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.635
+ $Y=0.665 $X2=2.775 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_2%B 3 7 8 9 13 15
r39 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.36
+ $X2=2.11 $Y2=1.525
r40 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.36
+ $X2=2.11 $Y2=1.195
r41 8 9 23.9527 $w=2.53e-07 $l=5.3e-07 $layer=LI1_cond $X=2.11 $Y=1.327 $X2=2.64
+ $Y2=1.327
r42 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.36 $X2=2.11 $Y2=1.36
r43 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.2 $Y=0.875 $X2=2.2
+ $Y2=1.195
r44 3 16 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.13 $Y=2.045
+ $X2=2.13 $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_2%A_28_367# 1 2 10 13 16 18 19 21 29 33
c58 16 0 1.62043e-19 $X=2.575 $Y=1.345
r59 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=0.39
+ $X2=2.65 $Y2=0.555
r60 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=0.39 $X2=2.65 $Y2=0.39
r61 26 29 3.57655 $w=2.88e-07 $l=9e-08 $layer=LI1_cond $X=0.175 $Y=2.065
+ $X2=0.265 $Y2=2.065
r62 24 25 8.11487 $w=4.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.305 $Y=0.875
+ $X2=0.305 $Y2=1.015
r63 21 24 6.83426 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.305 $Y=0.62
+ $X2=0.305 $Y2=0.875
r64 20 21 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.52 $Y=0.62
+ $X2=0.305 $Y2=0.62
r65 19 32 16.933 $w=3.45e-07 $l=4.54643e-07 $layer=LI1_cond $X=2.26 $Y=0.62
+ $X2=2.65 $Y2=0.48
r66 19 20 113.519 $w=1.68e-07 $l=1.74e-06 $layer=LI1_cond $X=2.26 $Y=0.62
+ $X2=0.52 $Y2=0.62
r67 18 26 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.175 $Y=1.92
+ $X2=0.175 $Y2=2.065
r68 18 25 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=0.175 $Y=1.92
+ $X2=0.175 $Y2=1.015
r69 15 16 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.575 $Y=1.195
+ $X2=2.575 $Y2=1.345
r70 13 16 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=2.56 $Y=2.045 $X2=2.56
+ $Y2=1.345
r71 10 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.56 $Y=0.875
+ $X2=2.56 $Y2=1.195
r72 10 36 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.56 $Y=0.875
+ $X2=2.56 $Y2=0.555
r73 2 29 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.045
r74 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.23
+ $Y=0.665 $X2=0.355 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_2%VPWR 1 2 3 12 18 22 26 28 30 35 42 43 46 49
+ 52
r33 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 43 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 40 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.94 $Y=3.33
+ $X2=2.775 $Y2=3.33
r38 40 42 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.94 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 39 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r41 36 46 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.92 $Y=3.33 $X2=0.76
+ $Y2=3.33
r42 36 38 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.92 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 35 49 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.782 $Y2=3.33
r44 35 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 30 46 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.6 $Y=3.33 $X2=0.76
+ $Y2=3.33
r48 30 32 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=3.33 $X2=0.24
+ $Y2=3.33
r49 28 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 28 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 24 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=3.245
+ $X2=2.775 $Y2=3.33
r53 24 26 40.8593 $w=3.28e-07 $l=1.17e-06 $layer=LI1_cond $X=2.775 $Y=3.245
+ $X2=2.775 $Y2=2.075
r54 23 49 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=2.08 $Y=3.33
+ $X2=1.782 $Y2=3.33
r55 22 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=2.775 $Y2=3.33
r56 22 23 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=2.08 $Y2=3.33
r57 18 21 8.04086 $w=5.93e-07 $l=4e-07 $layer=LI1_cond $X=1.782 $Y=2.05
+ $X2=1.782 $Y2=2.45
r58 16 49 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.782 $Y=3.245
+ $X2=1.782 $Y2=3.33
r59 16 21 15.9812 $w=5.93e-07 $l=7.95e-07 $layer=LI1_cond $X=1.782 $Y=3.245
+ $X2=1.782 $Y2=2.45
r60 12 15 14.7657 $w=3.18e-07 $l=4.1e-07 $layer=LI1_cond $X=0.76 $Y=2.085
+ $X2=0.76 $Y2=2.495
r61 10 46 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=3.33
r62 10 15 27.0104 $w=3.18e-07 $l=7.5e-07 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=2.495
r63 3 26 600 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.835 $X2=2.775 $Y2=2.075
r64 2 21 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=1.51
+ $Y=1.835 $X2=1.65 $Y2=2.45
r65 2 18 600 $w=1.7e-07 $l=5.01099e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.835 $X2=1.915 $Y2=2.05
r66 1 15 300 $w=1.7e-07 $l=7.6857e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.835 $X2=0.79 $Y2=2.495
r67 1 12 600 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.835 $X2=0.695 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_2%X 1 2 11 13 14 15 16 17
c24 13 0 1.94138e-19 $X=1.2 $Y=1.295
r25 17 35 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=1.202 $Y=2.775
+ $X2=1.202 $Y2=2.91
r26 16 17 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.202 $Y=2.405
+ $X2=1.202 $Y2=2.775
r27 15 16 21.7684 $w=2.23e-07 $l=4.25e-07 $layer=LI1_cond $X=1.202 $Y=1.98
+ $X2=1.202 $Y2=2.405
r28 14 15 16.1342 $w=2.23e-07 $l=3.15e-07 $layer=LI1_cond $X=1.202 $Y=1.665
+ $X2=1.202 $Y2=1.98
r29 13 14 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.202 $Y=1.295
+ $X2=1.202 $Y2=1.665
r30 8 13 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.202 $Y=1.125
+ $X2=1.202 $Y2=1.295
r31 7 11 8.89686 $w=2.48e-07 $l=1.93e-07 $layer=LI1_cond $X=1.202 $Y=1 $X2=1.395
+ $Y2=1
r32 7 8 1.37548 $w=2.25e-07 $l=1.25e-07 $layer=LI1_cond $X=1.202 $Y=1 $X2=1.202
+ $Y2=1.125
r33 2 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.22 $Y2=2.91
r34 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.22 $Y2=1.98
r35 1 11 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=1.255
+ $Y=0.245 $X2=1.395 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_2%VGND 1 2 9 10 16 26 27 30
r30 30 34 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.885
+ $Y2=0.26
r31 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r32 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r33 24 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r34 23 26 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r35 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r36 18 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=0.885
+ $Y2=0
r37 18 20 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=1.68
+ $Y2=0
r38 16 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r39 16 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r40 16 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r41 12 23 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.16
+ $Y2=0
r42 10 20 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.68
+ $Y2=0
r43 9 14 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.905
+ $Y2=0.26
r44 9 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=2.07
+ $Y2=0
r45 9 10 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.74
+ $Y2=0
r46 2 14 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.245 $X2=1.905 $Y2=0.26
r47 1 34 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=0.665
+ $Y=0.665 $X2=0.885 $Y2=0.26
.ends

