* File: sky130_fd_sc_lp__o41a_m.pxi.spice
* Created: Wed Sep  2 10:27:55 2020
* 
x_PM_SKY130_FD_SC_LP__O41A_M%A_80_21# N_A_80_21#_M1009_s N_A_80_21#_M1007_d
+ N_A_80_21#_M1006_g N_A_80_21#_c_92_n N_A_80_21#_M1002_g N_A_80_21#_c_94_n
+ N_A_80_21#_c_95_n N_A_80_21#_c_96_n N_A_80_21#_c_97_n N_A_80_21#_c_98_n
+ N_A_80_21#_c_103_n N_A_80_21#_c_104_n N_A_80_21#_c_99_n N_A_80_21#_c_105_n
+ N_A_80_21#_c_100_n PM_SKY130_FD_SC_LP__O41A_M%A_80_21#
x_PM_SKY130_FD_SC_LP__O41A_M%B1 N_B1_M1007_g N_B1_M1009_g N_B1_c_167_n
+ N_B1_c_172_n N_B1_c_173_n N_B1_c_168_n B1 B1 B1 N_B1_c_174_n
+ PM_SKY130_FD_SC_LP__O41A_M%B1
x_PM_SKY130_FD_SC_LP__O41A_M%A4 N_A4_c_219_n N_A4_M1003_g N_A4_M1001_g
+ N_A4_c_227_n N_A4_c_220_n N_A4_c_221_n A4 A4 A4 A4 A4 N_A4_c_223_n
+ N_A4_c_224_n PM_SKY130_FD_SC_LP__O41A_M%A4
x_PM_SKY130_FD_SC_LP__O41A_M%A3 N_A3_M1004_g N_A3_M1008_g N_A3_c_275_n
+ N_A3_c_276_n A3 A3 A3 A3 N_A3_c_278_n PM_SKY130_FD_SC_LP__O41A_M%A3
x_PM_SKY130_FD_SC_LP__O41A_M%A2 N_A2_M1010_g N_A2_M1000_g N_A2_c_321_n
+ N_A2_c_322_n A2 A2 A2 A2 N_A2_c_319_n PM_SKY130_FD_SC_LP__O41A_M%A2
x_PM_SKY130_FD_SC_LP__O41A_M%A1 N_A1_c_368_n N_A1_M1011_g N_A1_c_369_n
+ N_A1_c_370_n N_A1_M1005_g N_A1_c_365_n N_A1_c_366_n N_A1_c_372_n A1 A1 A1 A1
+ N_A1_c_374_n PM_SKY130_FD_SC_LP__O41A_M%A1
x_PM_SKY130_FD_SC_LP__O41A_M%X N_X_M1006_s N_X_M1002_s X X X X X N_X_c_404_n X
+ N_X_c_406_n PM_SKY130_FD_SC_LP__O41A_M%X
x_PM_SKY130_FD_SC_LP__O41A_M%VPWR N_VPWR_M1002_d N_VPWR_M1011_d N_VPWR_c_421_n
+ N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_424_n VPWR N_VPWR_c_425_n
+ N_VPWR_c_426_n N_VPWR_c_420_n N_VPWR_c_428_n PM_SKY130_FD_SC_LP__O41A_M%VPWR
x_PM_SKY130_FD_SC_LP__O41A_M%VGND N_VGND_M1006_d N_VGND_M1001_d N_VGND_M1000_d
+ N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n
+ N_VGND_c_477_n N_VGND_c_478_n VGND N_VGND_c_479_n N_VGND_c_480_n
+ N_VGND_c_481_n N_VGND_c_482_n PM_SKY130_FD_SC_LP__O41A_M%VGND
x_PM_SKY130_FD_SC_LP__O41A_M%A_300_51# N_A_300_51#_M1009_d N_A_300_51#_M1008_d
+ N_A_300_51#_M1005_d N_A_300_51#_c_529_n N_A_300_51#_c_530_n
+ N_A_300_51#_c_531_n N_A_300_51#_c_532_n N_A_300_51#_c_533_n
+ N_A_300_51#_c_534_n N_A_300_51#_c_535_n PM_SKY130_FD_SC_LP__O41A_M%A_300_51#
cc_1 VNB N_A_80_21#_c_92_n 0.0239125f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.238
cc_2 VNB N_A_80_21#_M1002_g 0.014714f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.885
cc_3 VNB N_A_80_21#_c_94_n 0.0292158f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.435
cc_4 VNB N_A_80_21#_c_95_n 0.00206039f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_5 VNB N_A_80_21#_c_96_n 0.0236002f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_6 VNB N_A_80_21#_c_97_n 0.0132837f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.81
cc_7 VNB N_A_80_21#_c_98_n 0.00165376f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.81
cc_8 VNB N_A_80_21#_c_99_n 9.78793e-19 $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.53
cc_9 VNB N_A_80_21#_c_100_n 0.0231723f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=0.765
cc_10 VNB N_B1_M1009_g 0.0216272f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_11 VNB N_B1_c_167_n 0.03633f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.435
cc_12 VNB N_B1_c_168_n 0.0286522f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.895
cc_13 VNB B1 0.00518501f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_14 VNB N_A4_c_219_n 0.0188733f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=2.675
cc_15 VNB N_A4_c_220_n 0.0162771f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.885
cc_16 VNB N_A4_c_221_n 0.0130957f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.885
cc_17 VNB A4 0.00132294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A4_c_223_n 0.020126f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.725
cc_19 VNB N_A4_c_224_n 0.0162722f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.53
cc_20 VNB N_A3_M1008_g 0.0348337f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_21 VNB N_A3_c_275_n 0.0234776f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.238
cc_22 VNB N_A3_c_276_n 3.47302e-19 $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.435
cc_23 VNB A3 0.0014048f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.885
cc_24 VNB N_A3_c_278_n 0.0165463f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.81
cc_25 VNB N_A2_M1000_g 0.0521953f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_26 VNB A2 0.0084058f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.885
cc_27 VNB N_A2_c_319_n 0.0158031f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.81
cc_28 VNB N_A1_M1005_g 0.043663f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_29 VNB N_A1_c_365_n 0.0324743f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.885
cc_30 VNB N_A1_c_366_n 0.0243252f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.895
cc_31 VNB A1 0.0263625f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_32 VNB N_X_c_404_n 0.0491632f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_33 VNB N_VPWR_c_420_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=0.93
cc_34 VNB N_VGND_c_472_n 0.00495479f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.435
cc_35 VNB N_VGND_c_473_n 0.00495206f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.435
cc_36 VNB N_VGND_c_474_n 0.00495206f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_37 VNB N_VGND_c_475_n 0.0320583f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.81
cc_38 VNB N_VGND_c_476_n 0.00401244f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.53
cc_39 VNB N_VGND_c_477_n 0.0174548f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.725
cc_40 VNB N_VGND_c_478_n 0.00401244f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.53
cc_41 VNB N_VGND_c_479_n 0.0189732f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=2.615
cc_42 VNB N_VGND_c_480_n 0.0253882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_481_n 0.23625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_482_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_300_51#_c_529_n 0.00100113f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.435
cc_46 VNB N_A_300_51#_c_530_n 0.00994006f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.885
cc_47 VNB N_A_300_51#_c_531_n 0.0028056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_300_51#_c_532_n 0.00114865f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.445
cc_49 VNB N_A_300_51#_c_533_n 0.0194167f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_50 VNB N_A_300_51#_c_534_n 0.00317049f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.53
cc_51 VNB N_A_300_51#_c_535_n 0.0067463f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.725
cc_52 VPB N_A_80_21#_M1002_g 0.0753931f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.885
cc_53 VPB N_A_80_21#_c_95_n 0.00738931f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.93
cc_54 VPB N_A_80_21#_c_103_n 0.0182952f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=2.53
cc_55 VPB N_A_80_21#_c_104_n 0.00205971f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.53
cc_56 VPB N_A_80_21#_c_105_n 9.7767e-19 $X=-0.19 $Y=1.655 $X2=1.33 $Y2=2.82
cc_57 VPB N_B1_M1007_g 0.027292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_B1_c_167_n 9.40404e-19 $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.435
cc_59 VPB N_B1_c_172_n 0.0230837f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.885
cc_60 VPB N_B1_c_173_n 0.0158081f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.885
cc_61 VPB N_B1_c_174_n 0.0163775f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=0.725
cc_62 VPB N_A4_c_219_n 0.00302549f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=2.675
cc_63 VPB N_A4_M1003_g 0.0527979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A4_c_227_n 0.021813f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.435
cc_65 VPB A4 0.00680737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A3_M1004_g 0.0565156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A3_c_276_n 0.0183998f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.435
cc_68 VPB A3 0.00661342f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.885
cc_69 VPB N_A2_M1010_g 0.0342961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A2_c_321_n 0.0316978f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_71 VPB N_A2_c_322_n 0.02747f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.238
cc_72 VPB A2 0.00993929f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.885
cc_73 VPB N_A2_c_319_n 0.00101463f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.81
cc_74 VPB N_A1_c_368_n 0.0207587f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=0.255
cc_75 VPB N_A1_c_369_n 0.0528667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A1_c_370_n 0.00651614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A1_c_366_n 9.11448e-19 $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.895
cc_78 VPB N_A1_c_372_n 0.0484921f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.445
cc_79 VPB A1 0.0331466f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.93
cc_80 VPB N_A1_c_374_n 0.0191013f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=0.53
cc_81 VPB N_X_c_404_n 0.0559233f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.93
cc_82 VPB N_X_c_406_n 0.0113339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_421_n 0.00482922f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_84 VPB N_VPWR_c_422_n 0.0127533f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.885
cc_85 VPB N_VPWR_c_423_n 0.0231054f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.435
cc_86 VPB N_VPWR_c_424_n 0.00362661f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.895
cc_87 VPB N_VPWR_c_425_n 0.0567279f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=2.53
cc_88 VPB N_VPWR_c_426_n 0.0210774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_420_n 0.0571955f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=0.93
cc_90 VPB N_VPWR_c_428_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 N_A_80_21#_M1002_g N_B1_M1007_g 0.0240613f $X=0.67 $Y=2.885 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_95_n N_B1_M1007_g 5.81548e-19 $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_103_n N_B1_M1007_g 0.0119095f $X=1.225 $Y=2.53 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_105_n N_B1_M1007_g 0.00147946f $X=1.33 $Y=2.82 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_96_n N_B1_M1009_g 7.6453e-19 $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_97_n N_B1_M1009_g 0.0016851f $X=1.105 $Y=0.81 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_99_n N_B1_M1009_g 0.00116361f $X=1.21 $Y=0.53 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_92_n N_B1_c_167_n 0.0114718f $X=0.597 $Y=1.238 $X2=0 $Y2=0
cc_99 N_A_80_21#_M1002_g N_B1_c_167_n 0.00614442f $X=0.67 $Y=2.885 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_95_n N_B1_c_167_n 4.33687e-19 $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_103_n N_B1_c_173_n 0.00521921f $X=1.225 $Y=2.53 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_95_n N_B1_c_168_n 0.00166978f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_96_n N_B1_c_168_n 0.0114718f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_97_n N_B1_c_168_n 0.0112675f $X=1.105 $Y=0.81 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_92_n B1 0.00193259f $X=0.597 $Y=1.238 $X2=0 $Y2=0
cc_106 N_A_80_21#_M1002_g B1 0.00359122f $X=0.67 $Y=2.885 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_95_n B1 0.059048f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_97_n B1 0.0174857f $X=1.105 $Y=0.81 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_103_n B1 0.0249264f $X=1.225 $Y=2.53 $X2=0 $Y2=0
cc_110 N_A_80_21#_M1002_g N_B1_c_174_n 0.039167f $X=0.67 $Y=2.885 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_95_n N_B1_c_174_n 0.00250158f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_103_n N_A4_M1003_g 0.00139033f $X=1.225 $Y=2.53 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_105_n N_A4_M1003_g 0.00340664f $X=1.33 $Y=2.82 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_103_n A4 0.0131381f $X=1.225 $Y=2.53 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_105_n A4 0.0166463f $X=1.33 $Y=2.82 $X2=0 $Y2=0
cc_116 N_A_80_21#_M1002_g N_X_c_404_n 0.0119249f $X=0.67 $Y=2.885 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_95_n N_X_c_404_n 0.111727f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_98_n N_X_c_404_n 0.0131664f $X=0.715 $Y=0.81 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_104_n N_X_c_404_n 0.0139873f $X=0.715 $Y=2.53 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_100_n N_X_c_404_n 0.0221785f $X=0.597 $Y=0.765 $X2=0 $Y2=0
cc_121 N_A_80_21#_M1002_g N_X_c_406_n 0.00286108f $X=0.67 $Y=2.885 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_104_n N_X_c_406_n 0.00371979f $X=0.715 $Y=2.53 $X2=0 $Y2=0
cc_123 N_A_80_21#_M1002_g N_VPWR_c_421_n 0.00277144f $X=0.67 $Y=2.885 $X2=0
+ $Y2=0
cc_124 N_A_80_21#_c_103_n N_VPWR_c_421_n 0.01326f $X=1.225 $Y=2.53 $X2=0 $Y2=0
cc_125 N_A_80_21#_M1002_g N_VPWR_c_423_n 0.00425667f $X=0.67 $Y=2.885 $X2=0
+ $Y2=0
cc_126 N_A_80_21#_c_103_n N_VPWR_c_423_n 0.00124851f $X=1.225 $Y=2.53 $X2=0
+ $Y2=0
cc_127 N_A_80_21#_c_104_n N_VPWR_c_423_n 0.00142127f $X=0.715 $Y=2.53 $X2=0
+ $Y2=0
cc_128 N_A_80_21#_c_103_n N_VPWR_c_425_n 0.00335002f $X=1.225 $Y=2.53 $X2=0
+ $Y2=0
cc_129 N_A_80_21#_c_105_n N_VPWR_c_425_n 0.00777502f $X=1.33 $Y=2.82 $X2=0 $Y2=0
cc_130 N_A_80_21#_M1007_d N_VPWR_c_420_n 0.00548586f $X=1.19 $Y=2.675 $X2=0
+ $Y2=0
cc_131 N_A_80_21#_M1002_g N_VPWR_c_420_n 0.00695851f $X=0.67 $Y=2.885 $X2=0
+ $Y2=0
cc_132 N_A_80_21#_c_103_n N_VPWR_c_420_n 0.00836575f $X=1.225 $Y=2.53 $X2=0
+ $Y2=0
cc_133 N_A_80_21#_c_104_n N_VPWR_c_420_n 0.00238635f $X=0.715 $Y=2.53 $X2=0
+ $Y2=0
cc_134 N_A_80_21#_c_105_n N_VPWR_c_420_n 0.00691106f $X=1.33 $Y=2.82 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_96_n N_VGND_c_472_n 0.00139794f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_97_n N_VGND_c_472_n 0.00594593f $X=1.105 $Y=0.81 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_98_n N_VGND_c_472_n 0.0099165f $X=0.715 $Y=0.81 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_99_n N_VGND_c_472_n 0.0086771f $X=1.21 $Y=0.53 $X2=0 $Y2=0
cc_139 N_A_80_21#_c_100_n N_VGND_c_472_n 0.00460896f $X=0.597 $Y=0.765 $X2=0
+ $Y2=0
cc_140 N_A_80_21#_c_97_n N_VGND_c_475_n 0.00469837f $X=1.105 $Y=0.81 $X2=0 $Y2=0
cc_141 N_A_80_21#_c_99_n N_VGND_c_475_n 0.00797539f $X=1.21 $Y=0.53 $X2=0 $Y2=0
cc_142 N_A_80_21#_c_98_n N_VGND_c_479_n 6.60115e-19 $X=0.715 $Y=0.81 $X2=0 $Y2=0
cc_143 N_A_80_21#_c_100_n N_VGND_c_479_n 0.00580462f $X=0.597 $Y=0.765 $X2=0
+ $Y2=0
cc_144 N_A_80_21#_c_97_n N_VGND_c_481_n 0.00860138f $X=1.105 $Y=0.81 $X2=0 $Y2=0
cc_145 N_A_80_21#_c_98_n N_VGND_c_481_n 0.00165007f $X=0.715 $Y=0.81 $X2=0 $Y2=0
cc_146 N_A_80_21#_c_99_n N_VGND_c_481_n 0.00754715f $X=1.21 $Y=0.53 $X2=0 $Y2=0
cc_147 N_A_80_21#_c_100_n N_VGND_c_481_n 0.012818f $X=0.597 $Y=0.765 $X2=0 $Y2=0
cc_148 N_A_80_21#_c_97_n N_A_300_51#_c_529_n 0.00139521f $X=1.105 $Y=0.81 $X2=0
+ $Y2=0
cc_149 N_A_80_21#_c_99_n N_A_300_51#_c_529_n 0.00314476f $X=1.21 $Y=0.53 $X2=0
+ $Y2=0
cc_150 N_A_80_21#_c_97_n N_A_300_51#_c_531_n 0.0113496f $X=1.105 $Y=0.81 $X2=0
+ $Y2=0
cc_151 N_B1_c_174_n N_A4_c_219_n 0.0169535f $X=1.12 $Y=1.84 $X2=0 $Y2=0
cc_152 N_B1_M1007_g N_A4_M1003_g 0.0214361f $X=1.115 $Y=2.885 $X2=0 $Y2=0
cc_153 N_B1_c_173_n N_A4_M1003_g 0.0169535f $X=1.12 $Y=2.345 $X2=0 $Y2=0
cc_154 N_B1_c_172_n N_A4_c_227_n 0.0169535f $X=1.12 $Y=2.18 $X2=0 $Y2=0
cc_155 N_B1_M1009_g N_A4_c_220_n 0.0142081f $X=1.425 $Y=0.465 $X2=0 $Y2=0
cc_156 N_B1_M1009_g N_A4_c_221_n 0.00589822f $X=1.425 $Y=0.465 $X2=0 $Y2=0
cc_157 N_B1_M1007_g A4 7.20149e-19 $X=1.115 $Y=2.885 $X2=0 $Y2=0
cc_158 N_B1_c_167_n A4 0.00344495f $X=1.12 $Y=1.675 $X2=0 $Y2=0
cc_159 B1 A4 0.0464531f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_160 N_B1_c_167_n N_A4_c_223_n 0.0169535f $X=1.12 $Y=1.675 $X2=0 $Y2=0
cc_161 N_B1_c_168_n N_A4_c_223_n 3.7023e-19 $X=1.425 $Y=0.895 $X2=0 $Y2=0
cc_162 B1 N_A4_c_223_n 0.00380839f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_163 N_B1_c_167_n N_A4_c_224_n 0.00831692f $X=1.12 $Y=1.675 $X2=0 $Y2=0
cc_164 N_B1_c_168_n N_A4_c_224_n 0.00589822f $X=1.425 $Y=0.895 $X2=0 $Y2=0
cc_165 N_B1_M1007_g N_VPWR_c_421_n 0.00279837f $X=1.115 $Y=2.885 $X2=0 $Y2=0
cc_166 N_B1_M1007_g N_VPWR_c_425_n 0.00436487f $X=1.115 $Y=2.885 $X2=0 $Y2=0
cc_167 N_B1_M1007_g N_VPWR_c_420_n 0.00616409f $X=1.115 $Y=2.885 $X2=0 $Y2=0
cc_168 N_B1_M1009_g N_VGND_c_472_n 0.00451066f $X=1.425 $Y=0.465 $X2=0 $Y2=0
cc_169 N_B1_M1009_g N_VGND_c_475_n 0.00565115f $X=1.425 $Y=0.465 $X2=0 $Y2=0
cc_170 N_B1_M1009_g N_VGND_c_481_n 0.0119838f $X=1.425 $Y=0.465 $X2=0 $Y2=0
cc_171 N_B1_c_168_n N_VGND_c_481_n 7.33874e-19 $X=1.425 $Y=0.895 $X2=0 $Y2=0
cc_172 N_B1_M1009_g N_A_300_51#_c_529_n 5.68223e-19 $X=1.425 $Y=0.465 $X2=0
+ $Y2=0
cc_173 N_B1_M1009_g N_A_300_51#_c_531_n 0.00200864f $X=1.425 $Y=0.465 $X2=0
+ $Y2=0
cc_174 N_A4_M1003_g N_A3_M1004_g 0.034324f $X=1.57 $Y=2.885 $X2=0 $Y2=0
cc_175 N_A4_c_227_n N_A3_M1004_g 0.0114158f $X=1.677 $Y=1.88 $X2=0 $Y2=0
cc_176 A4 N_A3_M1004_g 0.0110045f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A4_c_220_n N_A3_M1008_g 0.0213215f $X=1.82 $Y=0.785 $X2=0 $Y2=0
cc_178 N_A4_c_224_n N_A3_M1008_g 0.00867821f $X=1.677 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A4_c_223_n N_A3_c_275_n 0.0114158f $X=1.68 $Y=1.375 $X2=0 $Y2=0
cc_180 N_A4_c_219_n N_A3_c_276_n 0.0114158f $X=1.677 $Y=1.698 $X2=0 $Y2=0
cc_181 N_A4_M1003_g A3 6.588e-19 $X=1.57 $Y=2.885 $X2=0 $Y2=0
cc_182 A4 A3 0.0574397f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A4_c_224_n A3 0.0029498f $X=1.677 $Y=1.21 $X2=0 $Y2=0
cc_184 A4 N_A3_c_278_n 0.00200475f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A4_c_224_n N_A3_c_278_n 0.0114158f $X=1.677 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A4_M1003_g N_VPWR_c_425_n 0.00524368f $X=1.57 $Y=2.885 $X2=0 $Y2=0
cc_187 A4 N_VPWR_c_425_n 0.00401892f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A4_M1003_g N_VPWR_c_420_n 0.00969422f $X=1.57 $Y=2.885 $X2=0 $Y2=0
cc_189 A4 N_VPWR_c_420_n 0.00549302f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_190 A4 A_329_535# 0.00329307f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_191 N_A4_c_220_n N_VGND_c_473_n 0.002825f $X=1.82 $Y=0.785 $X2=0 $Y2=0
cc_192 N_A4_c_220_n N_VGND_c_475_n 0.0042337f $X=1.82 $Y=0.785 $X2=0 $Y2=0
cc_193 N_A4_c_220_n N_VGND_c_481_n 0.00594773f $X=1.82 $Y=0.785 $X2=0 $Y2=0
cc_194 N_A4_c_220_n N_A_300_51#_c_529_n 9.4709e-19 $X=1.82 $Y=0.785 $X2=0 $Y2=0
cc_195 N_A4_c_220_n N_A_300_51#_c_530_n 0.00519604f $X=1.82 $Y=0.785 $X2=0 $Y2=0
cc_196 N_A4_c_221_n N_A_300_51#_c_530_n 0.0113981f $X=1.82 $Y=0.935 $X2=0 $Y2=0
cc_197 A4 N_A_300_51#_c_530_n 9.07762e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_198 N_A4_c_221_n N_A_300_51#_c_531_n 0.00263664f $X=1.82 $Y=0.935 $X2=0 $Y2=0
cc_199 A4 N_A_300_51#_c_531_n 0.00847662f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_200 N_A4_c_223_n N_A_300_51#_c_531_n 0.00331588f $X=1.68 $Y=1.375 $X2=0 $Y2=0
cc_201 N_A3_M1008_g N_A2_M1000_g 0.0315424f $X=2.285 $Y=0.465 $X2=0 $Y2=0
cc_202 A3 N_A2_M1000_g 9.49498e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A3_c_278_n N_A2_M1000_g 0.0117705f $X=2.235 $Y=1.31 $X2=0 $Y2=0
cc_204 N_A3_M1004_g N_A2_c_321_n 0.0739769f $X=2.145 $Y=2.885 $X2=0 $Y2=0
cc_205 A3 N_A2_c_321_n 0.00297013f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_206 N_A3_M1004_g N_A2_c_322_n 0.00615982f $X=2.145 $Y=2.885 $X2=0 $Y2=0
cc_207 N_A3_c_276_n N_A2_c_322_n 0.0117705f $X=2.235 $Y=1.815 $X2=0 $Y2=0
cc_208 A3 N_A2_c_322_n 7.72746e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_209 N_A3_M1004_g A2 0.00118062f $X=2.145 $Y=2.885 $X2=0 $Y2=0
cc_210 A3 A2 0.0788053f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_211 N_A3_c_278_n A2 0.0043091f $X=2.235 $Y=1.31 $X2=0 $Y2=0
cc_212 N_A3_c_275_n N_A2_c_319_n 0.0117705f $X=2.235 $Y=1.65 $X2=0 $Y2=0
cc_213 N_A3_M1004_g N_VPWR_c_425_n 0.00585385f $X=2.145 $Y=2.885 $X2=0 $Y2=0
cc_214 N_A3_M1004_g N_VPWR_c_420_n 0.00690179f $X=2.145 $Y=2.885 $X2=0 $Y2=0
cc_215 A3 N_VPWR_c_420_n 0.0084721f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_216 N_A3_M1008_g N_VGND_c_473_n 0.00153867f $X=2.285 $Y=0.465 $X2=0 $Y2=0
cc_217 N_A3_M1008_g N_VGND_c_477_n 0.0042337f $X=2.285 $Y=0.465 $X2=0 $Y2=0
cc_218 N_A3_M1008_g N_VGND_c_481_n 0.00594773f $X=2.285 $Y=0.465 $X2=0 $Y2=0
cc_219 N_A3_M1008_g N_A_300_51#_c_530_n 0.01371f $X=2.285 $Y=0.465 $X2=0 $Y2=0
cc_220 A3 N_A_300_51#_c_530_n 0.0150352f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_221 N_A3_c_278_n N_A_300_51#_c_530_n 0.00244198f $X=2.235 $Y=1.31 $X2=0 $Y2=0
cc_222 N_A3_M1008_g N_A_300_51#_c_532_n 9.4709e-19 $X=2.285 $Y=0.465 $X2=0 $Y2=0
cc_223 N_A3_c_278_n N_A_300_51#_c_535_n 2.1956e-19 $X=2.235 $Y=1.31 $X2=0 $Y2=0
cc_224 N_A2_M1010_g N_A1_c_370_n 0.0533082f $X=2.505 $Y=2.885 $X2=0 $Y2=0
cc_225 N_A2_c_321_n N_A1_c_370_n 0.0110256f $X=2.505 $Y=2.13 $X2=0 $Y2=0
cc_226 A2 N_A1_c_370_n 0.00708722f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_227 N_A2_M1000_g N_A1_M1005_g 0.0379811f $X=2.715 $Y=0.465 $X2=0 $Y2=0
cc_228 A2 N_A1_c_365_n 5.66509e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_229 N_A2_M1000_g N_A1_c_366_n 0.00275047f $X=2.715 $Y=0.465 $X2=0 $Y2=0
cc_230 A2 N_A1_c_366_n 0.00355534f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_231 N_A2_c_319_n N_A1_c_366_n 0.00840193f $X=2.805 $Y=1.67 $X2=0 $Y2=0
cc_232 N_A2_M1010_g N_A1_c_372_n 0.00122454f $X=2.505 $Y=2.885 $X2=0 $Y2=0
cc_233 N_A2_c_321_n N_A1_c_372_n 0.00898995f $X=2.505 $Y=2.13 $X2=0 $Y2=0
cc_234 A2 N_A1_c_372_n 0.00146166f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_235 N_A2_M1000_g A1 4.12109e-19 $X=2.715 $Y=0.465 $X2=0 $Y2=0
cc_236 A2 A1 0.0433212f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_237 N_A2_c_319_n A1 0.00249759f $X=2.805 $Y=1.67 $X2=0 $Y2=0
cc_238 N_A2_c_322_n N_A1_c_374_n 0.00840193f $X=2.805 $Y=2.055 $X2=0 $Y2=0
cc_239 N_A2_M1010_g N_VPWR_c_422_n 0.00238543f $X=2.505 $Y=2.885 $X2=0 $Y2=0
cc_240 N_A2_M1010_g N_VPWR_c_425_n 0.00585385f $X=2.505 $Y=2.885 $X2=0 $Y2=0
cc_241 N_A2_M1010_g N_VPWR_c_420_n 0.00993297f $X=2.505 $Y=2.885 $X2=0 $Y2=0
cc_242 A2 N_VPWR_c_420_n 0.0121826f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_243 N_A2_M1000_g N_VGND_c_474_n 0.00153867f $X=2.715 $Y=0.465 $X2=0 $Y2=0
cc_244 N_A2_M1000_g N_VGND_c_477_n 0.0042337f $X=2.715 $Y=0.465 $X2=0 $Y2=0
cc_245 N_A2_M1000_g N_VGND_c_481_n 0.00594773f $X=2.715 $Y=0.465 $X2=0 $Y2=0
cc_246 N_A2_M1000_g N_A_300_51#_c_532_n 9.4709e-19 $X=2.715 $Y=0.465 $X2=0 $Y2=0
cc_247 N_A2_M1000_g N_A_300_51#_c_533_n 0.0129107f $X=2.715 $Y=0.465 $X2=0 $Y2=0
cc_248 A2 N_A_300_51#_c_533_n 0.0150212f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_249 N_A2_c_319_n N_A_300_51#_c_533_n 0.00251178f $X=2.805 $Y=1.67 $X2=0 $Y2=0
cc_250 A2 N_A_300_51#_c_535_n 0.00307299f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_251 N_A1_c_368_n N_VPWR_c_422_n 0.0107354f $X=2.865 $Y=2.565 $X2=0 $Y2=0
cc_252 N_A1_c_369_n N_VPWR_c_422_n 0.00959211f $X=3.29 $Y=2.49 $X2=0 $Y2=0
cc_253 N_A1_c_368_n N_VPWR_c_425_n 0.00486043f $X=2.865 $Y=2.565 $X2=0 $Y2=0
cc_254 N_A1_c_369_n N_VPWR_c_426_n 0.00723527f $X=3.29 $Y=2.49 $X2=0 $Y2=0
cc_255 N_A1_c_368_n N_VPWR_c_420_n 0.00525025f $X=2.865 $Y=2.565 $X2=0 $Y2=0
cc_256 N_A1_c_369_n N_VPWR_c_420_n 0.00978923f $X=3.29 $Y=2.49 $X2=0 $Y2=0
cc_257 A1 N_VPWR_c_420_n 0.0116364f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_258 N_A1_M1005_g N_VGND_c_474_n 0.002825f $X=3.145 $Y=0.465 $X2=0 $Y2=0
cc_259 N_A1_M1005_g N_VGND_c_480_n 0.0042337f $X=3.145 $Y=0.465 $X2=0 $Y2=0
cc_260 N_A1_M1005_g N_VGND_c_481_n 0.00692566f $X=3.145 $Y=0.465 $X2=0 $Y2=0
cc_261 N_A1_M1005_g N_A_300_51#_c_533_n 0.0174965f $X=3.145 $Y=0.465 $X2=0 $Y2=0
cc_262 N_A1_c_365_n N_A_300_51#_c_533_n 0.00809352f $X=3.365 $Y=1.19 $X2=0 $Y2=0
cc_263 A1 N_A_300_51#_c_533_n 0.00556566f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_264 N_A1_M1005_g N_A_300_51#_c_534_n 0.0020107f $X=3.145 $Y=0.465 $X2=0 $Y2=0
cc_265 N_X_c_406_n N_VPWR_c_423_n 0.0196527f $X=0.455 $Y=2.9 $X2=0 $Y2=0
cc_266 N_X_M1002_s N_VPWR_c_420_n 0.00220403f $X=0.33 $Y=2.675 $X2=0 $Y2=0
cc_267 N_X_c_406_n N_VPWR_c_420_n 0.0166278f $X=0.455 $Y=2.9 $X2=0 $Y2=0
cc_268 N_X_c_404_n N_VGND_c_479_n 0.00877924f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_269 N_X_M1006_s N_VGND_c_481_n 0.0042053f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_270 N_X_c_404_n N_VGND_c_481_n 0.00770513f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_271 N_VPWR_c_420_n A_329_535# 0.0142521f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_272 N_VPWR_c_420_n A_444_535# 0.00620535f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_273 N_VPWR_c_420_n A_516_535# 0.00307853f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_274 N_VGND_c_475_n N_A_300_51#_c_529_n 0.00760345f $X=1.965 $Y=0 $X2=0 $Y2=0
cc_275 N_VGND_c_481_n N_A_300_51#_c_529_n 0.00755664f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_473_n N_A_300_51#_c_530_n 0.0140329f $X=2.07 $Y=0.4 $X2=0 $Y2=0
cc_277 N_VGND_c_475_n N_A_300_51#_c_530_n 0.0029308f $X=1.965 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_477_n N_A_300_51#_c_530_n 0.0029308f $X=2.825 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_481_n N_A_300_51#_c_530_n 0.0109017f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_477_n N_A_300_51#_c_532_n 0.00760345f $X=2.825 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_481_n N_A_300_51#_c_532_n 0.00755664f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_474_n N_A_300_51#_c_533_n 0.0140329f $X=2.93 $Y=0.4 $X2=0 $Y2=0
cc_283 N_VGND_c_477_n N_A_300_51#_c_533_n 0.0029308f $X=2.825 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_480_n N_A_300_51#_c_533_n 0.0029308f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_481_n N_A_300_51#_c_533_n 0.0109017f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_480_n N_A_300_51#_c_534_n 0.00799446f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_c_481_n N_A_300_51#_c_534_n 0.00755664f $X=3.6 $Y=0 $X2=0 $Y2=0
