# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a21oi_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a21oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.200000 3.230000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.375000 1.765000 1.615000 ;
        RECT 0.105000 1.615000 3.675000 1.785000 ;
        RECT 3.400000 1.345000 3.675000 1.615000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.425000 5.235000 1.760000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.646400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.820000 0.820000 4.260000 1.030000 ;
        RECT 4.055000 1.930000 5.585000 2.100000 ;
        RECT 4.055000 2.100000 4.295000 2.735000 ;
        RECT 4.060000 0.255000 4.260000 0.820000 ;
        RECT 4.070000 1.030000 4.260000 1.085000 ;
        RECT 4.070000 1.085000 5.585000 1.255000 ;
        RECT 4.910000 2.100000 5.155000 2.735000 ;
        RECT 4.940000 0.255000 5.130000 1.085000 ;
        RECT 5.415000 1.255000 5.585000 1.930000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.760000 0.085000 ;
        RECT 0.100000  0.085000 0.390000 1.095000 ;
        RECT 0.960000  0.085000 1.290000 0.865000 ;
        RECT 3.560000  0.085000 3.890000 0.650000 ;
        RECT 4.440000  0.085000 4.770000 0.915000 ;
        RECT 5.300000  0.085000 5.630000 0.915000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 5.760000 3.415000 ;
        RECT 0.530000 2.295000 0.860000 3.245000 ;
        RECT 1.390000 2.295000 1.720000 3.245000 ;
        RECT 2.250000 2.295000 2.580000 3.245000 ;
        RECT 3.110000 2.295000 3.440000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.100000 1.955000 3.885000 2.125000 ;
      RECT 0.100000 2.125000 0.360000 3.075000 ;
      RECT 0.560000 0.255000 0.790000 1.035000 ;
      RECT 0.560000 1.035000 1.650000 1.205000 ;
      RECT 1.030000 2.125000 1.220000 3.075000 ;
      RECT 1.460000 0.255000 3.380000 0.640000 ;
      RECT 1.460000 0.640000 1.650000 1.035000 ;
      RECT 1.900000 2.125000 2.080000 3.075000 ;
      RECT 2.750000 2.125000 2.940000 3.075000 ;
      RECT 3.610000 2.125000 3.885000 2.905000 ;
      RECT 3.610000 2.905000 5.630000 3.075000 ;
      RECT 4.465000 2.270000 4.740000 2.905000 ;
      RECT 5.325000 2.270000 5.630000 2.905000 ;
  END
END sky130_fd_sc_lp__a21oi_4
