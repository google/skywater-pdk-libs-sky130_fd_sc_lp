* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and2_lp2 A B VGND VNB VPB VPWR X
M1000 VPWR a_99_21# X VPB phighvt w=1e+06u l=250000u
+  ad=5.65e+11p pd=5.13e+06u as=2.85e+11p ps=2.57e+06u
M1001 a_129_47# a_99_21# X VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1002 a_99_21# A a_287_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1003 a_287_47# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1004 a_99_21# B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=3.1e+11p pd=2.62e+06u as=0p ps=0u
M1005 VPWR A a_99_21# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_99_21# a_129_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
