* File: sky130_fd_sc_lp__nand4b_lp.pex.spice
* Created: Fri Aug 28 10:51:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4B_LP%A_87_231# 1 2 7 9 13 15 19 23 27 34 35 36
c73 36 0 9.80814e-20 $X=3.067 $Y=0.91
r74 34 35 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.027 $Y=2.19
+ $X2=3.027 $Y2=2.025
r75 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.7
+ $Y=0.99 $X2=0.7 $Y2=0.99
r76 27 30 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.7 $Y=0.91 $X2=0.7
+ $Y2=0.99
r77 25 36 3.70735 $w=2.5e-07 $l=1.39155e-07 $layer=LI1_cond $X=3.17 $Y=0.995
+ $X2=3.067 $Y2=0.91
r78 25 35 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.17 $Y=0.995
+ $X2=3.17 $Y2=2.025
r79 21 36 3.70735 $w=2.5e-07 $l=9.53677e-08 $layer=LI1_cond $X=3.045 $Y=0.825
+ $X2=3.067 $Y2=0.91
r80 21 23 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.045 $Y=0.825
+ $X2=3.045 $Y2=0.47
r81 17 34 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=3.027 $Y=2.252
+ $X2=3.027 $Y2=2.19
r82 17 19 17.0343 $w=4.53e-07 $l=6.48e-07 $layer=LI1_cond $X=3.027 $Y=2.252
+ $X2=3.027 $Y2=2.9
r83 16 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=0.91
+ $X2=0.7 $Y2=0.91
r84 15 36 2.76166 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.88 $Y=0.91
+ $X2=3.067 $Y2=0.91
r85 15 16 131.46 $w=1.68e-07 $l=2.015e-06 $layer=LI1_cond $X=2.88 $Y=0.91
+ $X2=0.865 $Y2=0.91
r86 11 31 38.5326 $w=3.08e-07 $l=2.24332e-07 $layer=POLY_cond $X=0.79 $Y=0.825
+ $X2=0.65 $Y2=0.99
r87 11 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.79 $Y=0.825
+ $X2=0.79 $Y2=0.445
r88 7 31 47.2339 $w=3.08e-07 $l=3.31964e-07 $layer=POLY_cond $X=0.56 $Y=1.28
+ $X2=0.65 $Y2=0.99
r89 7 9 314.294 $w=2.5e-07 $l=1.265e-06 $layer=POLY_cond $X=0.56 $Y=1.28
+ $X2=0.56 $Y2=2.545
r90 2 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=2.045 $X2=2.965 $Y2=2.19
r91 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=2.045 $X2=2.965 $Y2=2.9
r92 1 23 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.905
+ $Y=0.235 $X2=3.045 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_LP%B 3 7 9 12 13
r44 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.615
+ $X2=1.09 $Y2=1.45
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.615 $X2=1.09 $Y2=1.615
r46 9 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=1.09 $Y2=1.615
r47 7 14 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.18 $Y=0.445
+ $X2=1.18 $Y2=1.45
r48 1 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.78
+ $X2=1.09 $Y2=1.615
r49 1 3 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.09 $Y=1.78 $X2=1.09
+ $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_LP%C 3 7 11 12 13 14 18
c45 12 0 1.99507e-19 $X=1.63 $Y=1.845
r46 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=1.295
+ $X2=1.63 $Y2=1.665
r47 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.34 $X2=1.63 $Y2=1.34
r48 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.63 $Y=1.68
+ $X2=1.63 $Y2=1.34
r49 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.68
+ $X2=1.63 $Y2=1.845
r50 10 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.175
+ $X2=1.63 $Y2=1.34
r51 7 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.62 $Y=2.545 $X2=1.62
+ $Y2=1.845
r52 3 10 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.57 $Y=0.445
+ $X2=1.57 $Y2=1.175
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_LP%D 1 3 8 12 15 16 17 18 19 23
c47 17 0 1.47526e-19 $X=2.17 $Y=1.845
r48 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=1.295
+ $X2=2.17 $Y2=1.665
r49 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.17
+ $Y=1.34 $X2=2.17 $Y2=1.34
r50 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.17 $Y=1.68
+ $X2=2.17 $Y2=1.34
r51 16 17 31.2043 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.68
+ $X2=2.17 $Y2=1.845
r52 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.175
+ $X2=2.17 $Y2=1.34
r53 10 12 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.96 $Y=0.805
+ $X2=2.08 $Y2=0.805
r54 8 17 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.15 $Y=2.545 $X2=2.15
+ $Y2=1.845
r55 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.08 $Y=0.88 $X2=2.08
+ $Y2=0.805
r56 4 15 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.08 $Y=0.88
+ $X2=2.08 $Y2=1.175
r57 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=0.73 $X2=1.96
+ $Y2=0.805
r58 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.96 $Y=0.73 $X2=1.96
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_LP%A_N 1 3 8 10 12 16 19 20 21 22 23 27
c50 27 0 9.80814e-20 $X=2.74 $Y=1.34
c51 8 0 4.74694e-20 $X=2.7 $Y=2.545
r52 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.74
+ $Y=1.34 $X2=2.74 $Y2=1.34
r53 23 28 9.85642 $w=3.78e-07 $l=3.25e-07 $layer=LI1_cond $X=2.715 $Y=1.665
+ $X2=2.715 $Y2=1.34
r54 22 28 1.36474 $w=3.78e-07 $l=4.5e-08 $layer=LI1_cond $X=2.715 $Y=1.295
+ $X2=2.715 $Y2=1.34
r55 20 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.74 $Y=1.68
+ $X2=2.74 $Y2=1.34
r56 20 21 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.68
+ $X2=2.74 $Y2=1.845
r57 19 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.175
+ $X2=2.74 $Y2=1.34
r58 15 16 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.65 $Y=0.805
+ $X2=2.83 $Y2=0.805
r59 13 15 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.47 $Y=0.805
+ $X2=2.65 $Y2=0.805
r60 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.83 $Y=0.73
+ $X2=2.83 $Y2=0.805
r61 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.83 $Y=0.73 $X2=2.83
+ $Y2=0.445
r62 8 21 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.7 $Y=2.545 $X2=2.7
+ $Y2=1.845
r63 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.65 $Y=0.88 $X2=2.65
+ $Y2=0.805
r64 4 19 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.65 $Y=0.88
+ $X2=2.65 $Y2=1.175
r65 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.47 $Y=0.73 $X2=2.47
+ $Y2=0.805
r66 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.47 $Y=0.73 $X2=2.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_LP%VPWR 1 2 3 10 12 14 18 22 27 28 29 36 37
+ 43
r51 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 31 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=3.33
+ $X2=1.355 $Y2=3.33
r58 31 33 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.52 $Y=3.33 $X2=2.16
+ $Y2=3.33
r59 29 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 29 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 27 33 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.25 $Y=3.33 $X2=2.16
+ $Y2=3.33
r62 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=2.415 $Y2=3.33
r63 26 36 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.58 $Y=3.33
+ $X2=3.12 $Y2=3.33
r64 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=3.33
+ $X2=2.415 $Y2=3.33
r65 22 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.415 $Y=2.19
+ $X2=2.415 $Y2=2.9
r66 20 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=3.245
+ $X2=2.415 $Y2=3.33
r67 20 25 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.415 $Y=3.245
+ $X2=2.415 $Y2=2.9
r68 16 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=3.33
r69 16 18 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=2.54
r70 15 40 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=3.33 $X2=0.23
+ $Y2=3.33
r71 14 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=3.33
+ $X2=1.355 $Y2=3.33
r72 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.19 $Y=3.33
+ $X2=0.46 $Y2=3.33
r73 10 40 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.23 $Y2=3.33
r74 10 12 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.475
r75 3 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=2.045 $X2=2.415 $Y2=2.9
r76 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=2.045 $X2=2.415 $Y2=2.19
r77 2 18 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=1.215
+ $Y=2.045 $X2=1.355 $Y2=2.54
r78 1 12 300 $w=1.7e-07 $l=4.97242e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.045 $X2=0.295 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_LP%Y 1 2 3 10 11 14 16 18 20 23 28 31 32
c60 18 0 1.94995e-19 $X=1.885 $Y=2.195
c61 16 0 1.99507e-19 $X=1.72 $Y=2.11
r62 31 32 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r63 26 32 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=1.96
+ $X2=0.24 $Y2=1.665
r64 23 31 32.569 $w=2.28e-07 $l=6.5e-07 $layer=LI1_cond $X=0.24 $Y=0.645
+ $X2=0.24 $Y2=1.295
r65 23 25 14.4929 $w=2.82e-07 $l=4.19375e-07 $layer=LI1_cond $X=0.24 $Y=0.645
+ $X2=0.575 $Y2=0.455
r66 18 30 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=2.195
+ $X2=1.885 $Y2=2.11
r67 18 20 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.885 $Y=2.195
+ $X2=1.885 $Y2=2.9
r68 17 28 8.61065 $w=1.7e-07 $l=1.80748e-07 $layer=LI1_cond $X=0.99 $Y=2.11
+ $X2=0.825 $Y2=2.077
r69 16 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=2.11
+ $X2=1.885 $Y2=2.11
r70 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.72 $Y=2.11
+ $X2=0.99 $Y2=2.11
r71 12 28 0.89609 $w=3.3e-07 $l=1.18e-07 $layer=LI1_cond $X=0.825 $Y=2.195
+ $X2=0.825 $Y2=2.077
r72 12 14 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.825 $Y=2.195
+ $X2=0.825 $Y2=2.9
r73 11 26 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=2.045
+ $X2=0.24 $Y2=1.96
r74 10 28 8.61065 $w=1.7e-07 $l=1.80291e-07 $layer=LI1_cond $X=0.66 $Y=2.045
+ $X2=0.825 $Y2=2.077
r75 10 11 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.66 $Y=2.045
+ $X2=0.355 $Y2=2.045
r76 3 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=2.045 $X2=1.885 $Y2=2.19
r77 3 20 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=2.045 $X2=1.885 $Y2=2.9
r78 2 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.045 $X2=0.825 $Y2=2.19
r79 2 14 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.045 $X2=0.825 $Y2=2.9
r80 1 25 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=0.43
+ $Y=0.235 $X2=0.575 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_LP%VGND 1 6 8 10 20 21 24
r37 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r39 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.175
+ $Y2=0
r41 18 20 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=3.12
+ $Y2=0
r42 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r43 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.175
+ $Y2=0
r45 10 16 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.68
+ $Y2=0
r46 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r47 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r48 8 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r49 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0
r50 4 6 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0.43
r51 1 6 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.035
+ $Y=0.235 $X2=2.175 $Y2=0.43
.ends

