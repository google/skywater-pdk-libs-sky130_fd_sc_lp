* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__ebufn_8 A TE_B VGND VNB VPB VPWR Z
X0 a_27_47# a_84_21# Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 Z a_84_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_27_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_27_47# a_84_21# Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_27_47# a_772_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_27_47# a_84_21# Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND a_772_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VPWR TE_B a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND a_772_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 Z a_84_21# a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_27_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_27_47# a_772_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VPWR TE_B a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_27_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_772_21# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR TE_B a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_27_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 Z a_84_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_27_367# a_84_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_27_367# a_84_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VPWR TE_B a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VPWR A a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_772_21# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 Z a_84_21# a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_27_367# a_84_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_27_47# a_84_21# Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 VGND A a_84_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 Z a_84_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_84_21# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 VGND a_772_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 Z a_84_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 a_27_47# a_772_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 a_27_47# a_772_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 a_84_21# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 VGND a_772_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 a_27_367# a_84_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 Z a_84_21# a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 Z a_84_21# a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
