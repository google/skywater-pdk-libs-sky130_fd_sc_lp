* File: sky130_fd_sc_lp__nor2_lp.pex.spice
* Created: Fri Aug 28 10:54:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2_LP%A 3 7 9 13 16 18 19 20 21 32
r37 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.485
+ $Y=1.345 $X2=0.485 $Y2=1.345
r38 20 21 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=2.035
r39 20 33 5.39078 $w=7.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=1.345
r40 19 33 0.842309 $w=7.08e-07 $l=5e-08 $layer=LI1_cond $X=0.48 $Y=1.295
+ $X2=0.48 $Y2=1.345
r41 17 32 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.485 $Y=1.685
+ $X2=0.485 $Y2=1.345
r42 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.685
+ $X2=0.485 $Y2=1.85
r43 15 32 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.485 $Y=1.33
+ $X2=0.485 $Y2=1.345
r44 15 16 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=0.485 $Y=1.33
+ $X2=0.485 $Y2=1.255
r45 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.965 $Y=1.18
+ $X2=0.965 $Y2=0.77
r46 10 16 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=1.255
+ $X2=0.485 $Y2=1.255
r47 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.89 $Y=1.255
+ $X2=0.965 $Y2=1.18
r48 9 10 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.89 $Y=1.255
+ $X2=0.65 $Y2=1.255
r49 7 18 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.575 $Y=2.66
+ $X2=0.575 $Y2=1.85
r50 1 16 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.575 $Y=1.18
+ $X2=0.485 $Y2=1.255
r51 1 3 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.575 $Y=1.18
+ $X2=0.575 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_LP%B 3 5 6 9 11 15 17 20 21 22 23 24 25 42
r41 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.875
+ $Y=1.345 $X2=1.875 $Y2=1.345
r42 24 25 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.405
+ $X2=1.92 $Y2=2.775
r43 23 24 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=1.92 $Y2=2.405
r44 22 23 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=1.665
+ $X2=1.92 $Y2=2.035
r45 22 43 5.39078 $w=7.08e-07 $l=3.2e-07 $layer=LI1_cond $X=1.92 $Y=1.665
+ $X2=1.92 $Y2=1.345
r46 21 43 0.842309 $w=7.08e-07 $l=5e-08 $layer=LI1_cond $X=1.92 $Y=1.295
+ $X2=1.92 $Y2=1.345
r47 20 42 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.875 $Y=1.7
+ $X2=1.875 $Y2=1.345
r48 19 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.18
+ $X2=1.875 $Y2=1.345
r49 15 19 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.785 $Y=0.77
+ $X2=1.785 $Y2=1.18
r50 12 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.47 $Y=1.775
+ $X2=1.395 $Y2=1.775
r51 11 20 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.71 $Y=1.775
+ $X2=1.875 $Y2=1.7
r52 11 12 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.71 $Y=1.775
+ $X2=1.47 $Y2=1.775
r53 7 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=1.7
+ $X2=1.395 $Y2=1.775
r54 7 9 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=1.395 $Y=1.7 $X2=1.395
+ $Y2=0.77
r55 5 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.32 $Y=1.775
+ $X2=1.395 $Y2=1.775
r56 5 6 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.32 $Y=1.775 $X2=1.04
+ $Y2=1.775
r57 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.965 $Y=1.85
+ $X2=1.04 $Y2=1.775
r58 1 3 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.965 $Y=1.85 $X2=0.965
+ $Y2=2.66
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_LP%VPB__2 1 4 6 8 15 16
r18 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r19 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r20 13 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r21 12 15 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r22 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r23 10 19 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.262 $Y2=3.33
r24 10 12 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 8 16 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r26 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.72
+ $Y2=3.33
r27 4 19 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.262 $Y2=3.33
r28 4 6 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.36 $Y2=2.66
r29 1 6 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=2.45 $X2=0.36 $Y2=2.66
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_LP%Y 1 2 7 8 9 10 11 12 13
r24 13 37 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.18 $Y=2.775
+ $X2=1.18 $Y2=2.66
r25 12 37 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.18 $Y=2.405
+ $X2=1.18 $Y2=2.66
r26 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=2.035
+ $X2=1.18 $Y2=2.405
r27 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=2.035
r28 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=1.295
+ $X2=1.18 $Y2=1.665
r29 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=0.925 $X2=1.18
+ $Y2=1.295
r30 8 25 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.18 $Y=0.925
+ $X2=1.18 $Y2=0.77
r31 7 25 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.18 $Y=0.555
+ $X2=1.18 $Y2=0.77
r32 2 37 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=2.45 $X2=1.18 $Y2=2.66
r33 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.56 $X2=1.18 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_LP%VNB__2 1 2 7 9 11 13 15 17 30
r26 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r29 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r30 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r31 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r32 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r33 18 26 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.262
+ $Y2=0
r34 18 20 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.72
+ $Y2=0
r35 17 29 4.52492 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2.117
+ $Y2=0
r36 17 23 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.68
+ $Y2=0
r37 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r38 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r39 11 29 3.24126 $w=3.3e-07 $l=1.53734e-07 $layer=LI1_cond $X=2 $Y=0.085
+ $X2=2.117 $Y2=0
r40 11 13 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0.77
r41 7 26 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.262 $Y2=0
r42 7 9 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.36 $Y2=0.77
r43 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.56 $X2=2 $Y2=0.77
r44 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.56 $X2=0.36 $Y2=0.77
.ends

