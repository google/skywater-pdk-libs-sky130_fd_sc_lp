* File: sky130_fd_sc_lp__sdfbbn_1.spice
* Created: Fri Aug 28 11:27:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfbbn_1.pex.spice"
.subckt sky130_fd_sc_lp__sdfbbn_1  VNB VPB SCD D SCE CLK_N SET_B RESET_B VPWR
+ Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* CLK_N	CLK_N
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1032 A_122_119# N_SCD_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1012 N_A_200_119#_M1012_d N_SCE_M1012_g A_122_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=1.428 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1007 A_314_119# N_D_M1007_g N_A_200_119#_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1029 AS=0.0882 PD=0.91 PS=0.84 NRD=54.276 NRS=38.568 M=1 R=2.8 SA=75001.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_328_429#_M1013_g A_314_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1428 AS=0.1029 PD=1.1 PS=0.91 NRD=47.136 NRS=54.276 M=1 R=2.8 SA=75001.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 N_A_328_429#_M1010_d N_SCE_M1010_g N_VGND_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1533 AS=0.1428 PD=1.57 PS=1.1 NRD=22.848 NRS=67.14 M=1 R=2.8
+ SA=75002.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1015 N_A_838_50#_M1015_d N_CLK_N_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.1533 PD=1.41 PS=1.57 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75000.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1039 N_VGND_M1039_d N_A_838_50#_M1039_g N_A_995_66#_M1039_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1491 AS=0.1239 PD=1.55 PS=1.43 NRD=19.992 NRS=2.856 M=1 R=2.8
+ SA=75000.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1005 N_A_1295_379#_M1005_d N_A_995_66#_M1005_g N_A_200_119#_M1005_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.133875 AS=0.1197 PD=1.09 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1028 A_1439_104# N_A_838_50#_M1028_g N_A_1295_379#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.133875 PD=0.84 PS=1.09 NRD=44.28 NRS=58.56 M=1 R=2.8
+ SA=75000.8 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1040 N_VGND_M1040_d N_A_1445_324#_M1040_g A_1439_104# VNB NSHORT L=0.15 W=0.42
+ AD=0.212714 AS=0.0882 PD=1.24415 PS=0.84 NRD=128.988 NRS=44.28 M=1 R=2.8
+ SA=75001.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1035 N_A_1752_60#_M1035_d N_SET_B_M1035_g N_VGND_M1040_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0912 AS=0.324136 PD=0.925 PS=1.89585 NRD=0 NRS=81.552 M=1
+ R=4.26667 SA=75001.8 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1000 N_A_1445_324#_M1000_d N_A_1295_379#_M1000_g N_A_1752_60#_M1035_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.185287 AS=0.0912 PD=1.41 PS=0.925 NRD=43.968
+ NRS=0.936 M=1 R=4.26667 SA=75002.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1008 N_A_1752_60#_M1008_d N_A_1926_21#_M1008_g N_A_1445_324#_M1000_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1824 AS=0.185287 PD=1.85 PS=1.41 NRD=0 NRS=43.968
+ M=1 R=4.26667 SA=75002.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1027 A_2198_119# N_A_1445_324#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1136 AS=0.1824 PD=0.995 PS=1.85 NRD=22.968 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1016 N_A_2299_119#_M1016_d N_A_838_50#_M1016_g A_2198_119# VNB NSHORT L=0.15
+ W=0.64 AD=0.129147 AS=0.1136 PD=1.20755 PS=0.995 NRD=0 NRS=22.968 M=1
+ R=4.26667 SA=75000.7 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1014 A_2401_163# N_A_995_66#_M1014_g N_A_2299_119#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=24.276 M=1
+ R=2.8 SA=75001.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_2449_137#_M1025_g A_2401_163# VNB NSHORT L=0.15 W=0.42
+ AD=0.166792 AS=0.0504 PD=1.21245 PS=0.66 NRD=97.74 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1022 N_A_2636_119#_M1022_d N_SET_B_M1022_g N_VGND_M1025_d VNB NSHORT L=0.15
+ W=0.64 AD=0.177775 AS=0.254158 PD=1.335 PS=1.84755 NRD=41.76 NRS=64.14 M=1
+ R=4.26667 SA=75001.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1036 N_A_2449_137#_M1036_d N_A_2299_119#_M1036_g N_A_2636_119#_M1022_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.176325 AS=0.177775 PD=1.325 PS=1.335 NRD=14.988
+ NRS=41.76 M=1 R=4.26667 SA=75002.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1017 N_A_2636_119#_M1017_d N_A_1926_21#_M1017_g N_A_2449_137#_M1036_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1824 AS=0.176325 PD=1.85 PS=1.325 NRD=0 NRS=15.936
+ M=1 R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_RESET_B_M1006_g N_A_1926_21#_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1021 N_Q_N_M1021_d N_A_2449_137#_M1021_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1806 PD=2.25 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1041 N_VGND_M1041_d N_A_2449_137#_M1041_g N_A_3279_367#_M1041_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0805 AS=0.1197 PD=0.776667 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1023 N_Q_M1023_d N_A_3279_367#_M1023_g N_VGND_M1041_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.161 PD=2.25 PS=1.55333 NRD=0 NRS=6.42 M=1 R=5.6 SA=75000.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1024 N_VPWR_M1024_d N_SCD_M1024_g N_A_27_474#_M1024_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1042 A_200_474# N_SCE_M1042_g N_VPWR_M1024_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1046 N_A_200_119#_M1046_d N_D_M1046_g A_200_474# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1031 N_A_27_474#_M1031_d N_A_328_429#_M1031_g N_A_200_119#_M1046_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1792 AS=0.0896 PD=1.84 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1047 N_A_328_429#_M1047_d N_SCE_M1047_g N_VPWR_M1047_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.352 PD=1.85 PS=2.38 NRD=0 NRS=83.0946 M=1 R=4.26667
+ SA=75000.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1029 N_A_838_50#_M1029_d N_CLK_N_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1792 AS=0.3552 PD=1.84 PS=2.39 NRD=0 NRS=83.0946 M=1 R=4.26667
+ SA=75000.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_VPWR_M1018_d N_A_838_50#_M1018_g N_A_995_66#_M1018_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.37 AS=0.1792 PD=3.01 PS=1.84 NRD=161.008 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1033 N_A_1295_379#_M1033_d N_A_838_50#_M1033_g N_A_200_119#_M1033_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0756 AS=0.1176 PD=0.78 PS=1.4 NRD=37.5088 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75004.9 A=0.063 P=1.14 MULT=1
MM1034 A_1397_379# N_A_995_66#_M1034_g N_A_1295_379#_M1033_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1445_324#_M1009_g A_1397_379# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.2345 AS=0.0504 PD=1.43333 PS=0.66 NRD=236.085 NRS=30.4759 M=1
+ R=2.8 SA=75001.1 SB=75004 A=0.063 P=1.14 MULT=1
MM1030 N_A_1445_324#_M1030_d N_SET_B_M1030_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.4179 AS=0.469 PD=1.835 PS=2.86667 NRD=167.667 NRS=18.7544 M=1
+ R=5.6 SA=75001.4 SB=75003.4 A=0.126 P=1.98 MULT=1
MM1001 A_1996_379# N_A_1295_379#_M1001_g N_A_1445_324#_M1030_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1008 AS=0.4179 PD=1.08 PS=1.835 NRD=15.2281 NRS=0 M=1 R=5.6
+ SA=75002.6 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_1926_21#_M1003_g A_1996_379# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1974 AS=0.1008 PD=1.31 PS=1.08 NRD=0 NRS=15.2281 M=1 R=5.6 SA=75003
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1043 A_2198_379# N_A_1445_324#_M1043_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.166862 AS=0.1974 PD=1.44 PS=1.31 NRD=33.687 NRS=44.5417 M=1 R=5.6
+ SA=75003.6 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1038 N_A_2299_119#_M1038_d N_A_995_66#_M1038_g A_2198_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1799 AS=0.166862 PD=1.6 PS=1.44 NRD=0 NRS=33.687 M=1 R=5.6
+ SA=75002.6 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1026 A_2401_506# N_A_838_50#_M1026_g N_A_2299_119#_M1038_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.13965 AS=0.08995 PD=1.085 PS=0.8 NRD=130.158 NRS=74.6433 M=1 R=2.8
+ SA=75002 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1037 N_VPWR_M1037_d N_A_2449_137#_M1037_g A_2401_506# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1218 AS=0.13965 PD=0.953333 PS=1.085 NRD=145.386 NRS=130.158 M=1
+ R=2.8 SA=75002.9 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1011 N_A_2449_137#_M1011_d N_SET_B_M1011_g N_VPWR_M1037_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1176 AS=0.2436 PD=1.12 PS=1.90667 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1045 A_2798_451# N_A_2299_119#_M1045_g N_A_2449_137#_M1011_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.0882 AS=0.1176 PD=1.05 PS=1.12 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75002.3 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1044 N_VPWR_M1044_d N_A_1926_21#_M1044_g A_2798_451# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75002.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1019 N_VPWR_M1019_d N_RESET_B_M1019_g N_A_1926_21#_M1019_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.137128 AS=0.1792 PD=1.09137 PS=1.84 NRD=49.0136 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1020 N_Q_N_M1020_d N_A_2449_137#_M1020_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3528 AS=0.269972 PD=3.08 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A_2449_137#_M1002_g N_A_3279_367#_M1002_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.137128 AS=0.1824 PD=1.09137 PS=1.85 NRD=25.3933 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1004 N_Q_M1004_d N_A_3279_367#_M1004_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.269972 PD=3.09 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX48_noxref VNB VPB NWDIODE A=33.8311 P=40.01
c_187 VNB 0 2.08564e-19 $X=0 $Y=0
c_348 VPB 0 3.7507e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfbbn_1.pxi.spice"
*
.ends
*
*
