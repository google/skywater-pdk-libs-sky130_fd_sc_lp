* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
X0 a_27_51# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_486_65# B a_217_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_697_69# C a_486_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_486_65# C a_697_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_217_65# B a_486_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_217_65# a_27_51# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_27_51# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_697_69# D VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND D a_697_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Y a_27_51# a_217_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 Y a_27_51# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VPWR a_27_51# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
