# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__maj3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__maj3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.180000 1.415000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.180000 2.305000 1.515000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.180000 0.905000 1.515000 ;
        RECT 0.735000 1.515000 0.905000 2.225000 ;
        RECT 0.735000 2.225000 2.655000 2.395000 ;
        RECT 2.485000 1.275000 2.980000 1.605000 ;
        RECT 2.485000 1.605000 2.655000 2.225000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.209600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.345000 1.785000 5.155000 1.955000 ;
        RECT 3.345000 1.955000 3.675000 3.065000 ;
        RECT 3.510000 0.265000 3.680000 0.925000 ;
        RECT 3.510000 0.925000 5.155000 1.095000 ;
        RECT 4.325000 0.265000 4.655000 0.925000 ;
        RECT 4.365000 1.955000 4.695000 3.065000 ;
        RECT 4.925000 1.095000 5.155000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 5.280000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 5.470000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.090000  0.830000 3.330000 1.000000 ;
      RECT 0.090000  1.000000 0.260000 1.795000 ;
      RECT 0.090000  1.795000 0.555000 3.065000 ;
      RECT 0.315000  0.265000 0.645000 0.830000 ;
      RECT 1.135000  0.085000 1.465000 0.650000 ;
      RECT 1.135000  2.575000 1.465000 3.245000 ;
      RECT 1.625000  1.000000 1.795000 1.795000 ;
      RECT 1.625000  1.795000 2.285000 2.045000 ;
      RECT 1.955000  0.295000 2.285000 0.830000 ;
      RECT 2.775000  0.085000 3.105000 0.650000 ;
      RECT 2.835000  1.795000 3.165000 3.245000 ;
      RECT 3.160000  1.000000 3.330000 1.275000 ;
      RECT 3.160000  1.275000 4.670000 1.605000 ;
      RECT 3.855000  2.135000 4.185000 3.245000 ;
      RECT 3.860000  0.085000 4.110000 0.745000 ;
      RECT 4.835000  0.085000 5.165000 0.745000 ;
      RECT 4.875000  2.135000 5.125000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_lp__maj3_4
END LIBRARY
