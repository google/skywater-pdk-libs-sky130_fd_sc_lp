* File: sky130_fd_sc_lp__dfrtp_2.pex.spice
* Created: Fri Aug 28 10:22:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFRTP_2%CLK 3 7 11 12 13 14 18 19
c36 18 0 6.65401e-20 $X=0.385 $Y=1.615
r37 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r38 13 14 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=2.035
r39 13 19 1.82927 $w=3.13e-07 $l=5e-08 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=1.615
r40 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.955
+ $X2=0.385 $Y2=1.615
r41 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.955
+ $X2=0.385 $Y2=2.12
r42 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.45
+ $X2=0.385 $Y2=1.615
r43 7 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.475 $Y=2.64
+ $X2=0.475 $Y2=2.12
r44 3 10 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=0.475 $Y=0.715
+ $X2=0.475 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%A_27_101# 1 2 8 11 15 18 22 25 29 30 33 37
+ 39 40 42 45 46 48 49 50 52 53 54 56 57 60 61 62 64 65 66 69 70 74 75 78 79 80
+ 83 87 91 92 94 96 103
c277 103 0 2.74955e-19 $X=7.01 $Y=0.515
c278 91 0 1.88632e-19 $X=3.415 $Y=0.362
c279 87 0 1.69354e-20 $X=3.3 $Y=1.3
c280 79 0 1.63461e-19 $X=0.895 $Y=1.185
c281 57 0 1.55293e-19 $X=4.05 $Y=0.362
c282 54 0 4.28297e-20 $X=2.58 $Y=0.362
c283 52 0 1.92879e-19 $X=2.495 $Y=0.87
c284 39 0 6.65401e-20 $X=0.665 $Y=1.185
r285 87 97 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.3 $X2=3.3
+ $Y2=1.465
r286 87 96 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.3 $X2=3.3
+ $Y2=1.135
r287 86 87 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.3
+ $Y=1.3 $X2=3.3 $Y2=1.3
r288 83 94 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.972 $Y=1.2
+ $X2=0.972 $Y2=1.035
r289 82 84 18.1207 $w=4.58e-07 $l=5.05e-07 $layer=LI1_cond $X=0.895 $Y=1.2
+ $X2=0.895 $Y2=1.705
r290 82 83 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=1.2 $X2=0.955 $Y2=1.2
r291 79 82 0.390026 $w=4.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.895 $Y=1.185
+ $X2=0.895 $Y2=1.2
r292 79 80 7.19996 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=1.185
+ $X2=0.895 $Y2=1.1
r293 75 103 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.01 $Y=0.35
+ $X2=7.01 $Y2=0.515
r294 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.01
+ $Y=0.35 $X2=7.01 $Y2=0.35
r295 72 92 5.28824 $w=1.75e-07 $l=9e-08 $layer=LI1_cond $X=6.355 $Y=0.345
+ $X2=6.265 $Y2=0.345
r296 72 74 40.3586 $w=1.78e-07 $l=6.55e-07 $layer=LI1_cond $X=6.355 $Y=0.345
+ $X2=7.01 $Y2=0.345
r297 70 100 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.26 $Y=1.91
+ $X2=6.26 $Y2=2.075
r298 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.26
+ $Y=1.91 $X2=6.26 $Y2=1.91
r299 67 92 1.24132 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=6.265 $Y=0.435
+ $X2=6.265 $Y2=0.345
r300 67 69 90.8838 $w=1.78e-07 $l=1.475e-06 $layer=LI1_cond $X=6.265 $Y=0.435
+ $X2=6.265 $Y2=1.91
r301 65 92 5.28824 $w=1.75e-07 $l=9.24662e-08 $layer=LI1_cond $X=6.175 $Y=0.34
+ $X2=6.265 $Y2=0.345
r302 65 66 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.175 $Y=0.34
+ $X2=5.655 $Y2=0.34
r303 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.57 $Y=0.425
+ $X2=5.655 $Y2=0.34
r304 63 64 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.57 $Y=0.425
+ $X2=5.57 $Y2=0.805
r305 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.485 $Y=0.89
+ $X2=5.57 $Y2=0.805
r306 61 62 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=5.485 $Y=0.89
+ $X2=4.22 $Y2=0.89
r307 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.135 $Y=0.805
+ $X2=4.22 $Y2=0.89
r308 59 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.135 $Y=0.47
+ $X2=4.135 $Y2=0.805
r309 58 91 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=0.362
+ $X2=3.415 $Y2=0.362
r310 57 59 6.93832 $w=2.15e-07 $l=1.44375e-07 $layer=LI1_cond $X=4.05 $Y=0.362
+ $X2=4.135 $Y2=0.47
r311 57 58 29.4811 $w=2.13e-07 $l=5.5e-07 $layer=LI1_cond $X=4.05 $Y=0.362
+ $X2=3.5 $Y2=0.362
r312 56 86 5.40943 $w=2.43e-07 $l=1.15e-07 $layer=LI1_cond $X=3.415 $Y=1.262
+ $X2=3.3 $Y2=1.262
r313 55 91 2.20034 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=3.415 $Y=0.47
+ $X2=3.415 $Y2=0.362
r314 55 56 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=0.47
+ $X2=3.415 $Y2=1.14
r315 53 91 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=0.362
+ $X2=3.415 $Y2=0.362
r316 53 54 40.2015 $w=2.13e-07 $l=7.5e-07 $layer=LI1_cond $X=3.33 $Y=0.362
+ $X2=2.58 $Y2=0.362
r317 51 54 6.93832 $w=2.15e-07 $l=1.44375e-07 $layer=LI1_cond $X=2.495 $Y=0.47
+ $X2=2.58 $Y2=0.362
r318 51 52 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.495 $Y=0.47
+ $X2=2.495 $Y2=0.87
r319 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.41 $Y=0.955
+ $X2=2.495 $Y2=0.87
r320 49 50 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.41 $Y=0.955
+ $X2=1.825 $Y2=0.955
r321 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.74 $Y=0.87
+ $X2=1.825 $Y2=0.955
r322 47 48 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.74 $Y=0.425
+ $X2=1.74 $Y2=0.87
r323 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.655 $Y=0.34
+ $X2=1.74 $Y2=0.425
r324 45 46 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.655 $Y=0.34
+ $X2=1.125 $Y2=0.34
r325 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.04 $Y=0.425
+ $X2=1.125 $Y2=0.34
r326 43 80 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.04 $Y=0.425
+ $X2=1.04 $Y2=1.1
r327 42 84 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.75 $Y=2.3
+ $X2=0.75 $Y2=1.705
r328 39 79 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.665 $Y=1.185
+ $X2=0.895 $Y2=1.185
r329 39 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.665 $Y=1.185
+ $X2=0.39 $Y2=1.185
r330 38 78 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.355 $Y=2.385
+ $X2=0.225 $Y2=2.385
r331 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=2.385
+ $X2=0.75 $Y2=2.3
r332 37 38 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.665 $Y=2.385
+ $X2=0.355 $Y2=2.385
r333 31 40 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=0.242 $Y=1.1
+ $X2=0.39 $Y2=1.185
r334 31 33 15.0404 $w=2.93e-07 $l=3.85e-07 $layer=LI1_cond $X=0.242 $Y=1.1
+ $X2=0.242 $Y2=0.715
r335 29 103 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.92 $Y=0.835
+ $X2=6.92 $Y2=0.515
r336 25 100 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.185 $Y=2.675
+ $X2=6.185 $Y2=2.075
r337 22 96 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.28 $Y=0.805
+ $X2=3.28 $Y2=1.135
r338 18 97 728.128 $w=1.5e-07 $l=1.42e-06 $layer=POLY_cond $X=3.26 $Y=2.885
+ $X2=3.26 $Y2=1.465
r339 15 94 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.08 $Y=0.715
+ $X2=1.08 $Y2=1.035
r340 11 30 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=0.905 $Y=2.64
+ $X2=0.905 $Y2=1.705
r341 8 30 43.7733 $w=3.65e-07 $l=1.82e-07 $layer=POLY_cond $X=0.972 $Y=1.523
+ $X2=0.972 $Y2=1.705
r342 7 83 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.972 $Y=1.217
+ $X2=0.972 $Y2=1.2
r343 7 8 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=0.972 $Y=1.217
+ $X2=0.972 $Y2=1.523
r344 2 78 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.26 $Y2=2.465
r345 1 33 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.505 $X2=0.26 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%D 3 5 6 9 14 15 18
c57 15 0 7.22623e-20 $X=2.16 $Y=1.295
r58 15 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.16
+ $Y=1.375 $X2=2.16 $Y2=1.375
r59 13 18 49.3587 $w=4e-07 $l=3.55e-07 $layer=POLY_cond $X=2.195 $Y=1.73
+ $X2=2.195 $Y2=1.375
r60 13 14 43.5898 $w=4e-07 $l=1.5e-07 $layer=POLY_cond $X=2.215 $Y=1.73
+ $X2=2.215 $Y2=1.88
r61 11 18 2.08558 $w=4e-07 $l=1.5e-08 $layer=POLY_cond $X=2.195 $Y=1.36
+ $X2=2.195 $Y2=1.375
r62 7 9 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.85 $Y=1.21 $X2=2.85
+ $Y2=0.805
r63 6 11 34.8994 $w=1.5e-07 $l=2.34521e-07 $layer=POLY_cond $X=2.395 $Y=1.285
+ $X2=2.195 $Y2=1.36
r64 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.775 $Y=1.285
+ $X2=2.85 $Y2=1.21
r65 5 6 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.775 $Y=1.285
+ $X2=2.395 $Y2=1.285
r66 3 14 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=2.36 $Y=2.885
+ $X2=2.36 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%A_196_464# 1 2 9 11 13 17 19 20 23 27 30 34
+ 37 38 39 44 45 49 50 51 52 55 61 65 66 72
c227 66 0 2.0317e-19 $X=6.96 $Y=1.62
c228 52 0 3.19907e-19 $X=3.745 $Y=1.665
c229 27 0 1.54549e-19 $X=6.88 $Y=2.125
c230 11 0 1.78156e-19 $X=3.98 $Y=1.205
r231 80 82 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.385 $Y=1.665
+ $X2=1.39 $Y2=1.665
r232 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.84
+ $Y=1.65 $X2=3.84 $Y2=1.65
r233 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.96
+ $Y=1.62 $X2=6.96 $Y2=1.62
r234 61 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.665
+ $X2=6.96 $Y2=1.665
r235 59 72 13.6503 $w=1.93e-07 $l=2.4e-07 $layer=LI1_cond $X=3.6 $Y=1.652
+ $X2=3.84 $Y2=1.652
r236 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=1.665
+ $X2=3.6 $Y2=1.665
r237 55 82 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.39 $Y2=1.665
r238 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.665
r239 52 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=1.665
+ $X2=3.6 $Y2=1.665
r240 51 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=1.665
+ $X2=6.96 $Y2=1.665
r241 51 52 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.815 $Y=1.665
+ $X2=3.745 $Y2=1.665
r242 50 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.825 $Y=1.665
+ $X2=1.68 $Y2=1.665
r243 49 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.455 $Y=1.665
+ $X2=3.6 $Y2=1.665
r244 49 50 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=3.455 $Y=1.665
+ $X2=1.825 $Y2=1.665
r245 45 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=2.09
+ $X2=2.81 $Y2=2.255
r246 44 47 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=2.775 $Y=2.09
+ $X2=2.775 $Y2=2.17
r247 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=2.09 $X2=2.81 $Y2=2.09
r248 39 42 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.475 $Y=2.17
+ $X2=1.385 $Y2=2.17
r249 38 47 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.645 $Y=2.17
+ $X2=2.775 $Y2=2.17
r250 38 39 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=2.645 $Y=2.17
+ $X2=1.475 $Y2=2.17
r251 37 42 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=2.085
+ $X2=1.385 $Y2=2.17
r252 36 80 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=1.83
+ $X2=1.385 $Y2=1.665
r253 36 37 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=1.385 $Y=1.83
+ $X2=1.385 $Y2=2.085
r254 32 82 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.5
+ $X2=1.39 $Y2=1.665
r255 32 34 43.1962 $w=1.88e-07 $l=7.4e-07 $layer=LI1_cond $X=1.39 $Y=1.5
+ $X2=1.39 $Y2=0.76
r256 28 42 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.155 $Y=2.17
+ $X2=1.385 $Y2=2.17
r257 28 30 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.155 $Y=2.255
+ $X2=1.155 $Y2=2.465
r258 26 65 28.3893 $w=4.9e-07 $l=2.6e-07 $layer=POLY_cond $X=6.88 $Y=1.88
+ $X2=6.88 $Y2=1.62
r259 26 27 54.9885 $w=4.9e-07 $l=2.45e-07 $layer=POLY_cond $X=6.88 $Y=1.88
+ $X2=6.88 $Y2=2.125
r260 25 65 9.28112 $w=4.9e-07 $l=8.5e-08 $layer=POLY_cond $X=6.88 $Y=1.535
+ $X2=6.88 $Y2=1.62
r261 23 27 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.71 $Y=2.885
+ $X2=6.71 $Y2=2.125
r262 19 25 184.911 $w=6.6e-08 $l=2.8e-07 $layer=POLY_cond $X=6.635 $Y=1.46
+ $X2=6.88 $Y2=1.535
r263 19 20 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=6.635 $Y=1.46
+ $X2=6.375 $Y2=1.46
r264 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.3 $Y=1.385
+ $X2=6.375 $Y2=1.46
r265 15 17 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=6.3 $Y=1.385
+ $X2=6.3 $Y2=0.635
r266 11 71 91.2799 $w=2.59e-07 $l=4.99199e-07 $layer=POLY_cond $X=3.98 $Y=1.205
+ $X2=3.865 $Y2=1.65
r267 11 13 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.98 $Y=1.205
+ $X2=3.98 $Y2=0.805
r268 9 69 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.79 $Y=2.885
+ $X2=2.79 $Y2=2.255
r269 2 30 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.32 $X2=1.12 $Y2=2.465
r270 1 34 182 $w=1.7e-07 $l=3.53483e-07 $layer=licon1_NDIFF $count=1 $X=1.155
+ $Y=0.505 $X2=1.39 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%A_709_411# 1 2 9 11 12 13 14 17 19 26 30 32
+ 33
c87 33 0 1.54549e-19 $X=5.965 $Y=2.405
c88 30 0 1.772e-19 $X=5.915 $Y=1.585
c89 19 0 1.58556e-19 $X=5.825 $Y=1.585
c90 17 0 1.55293e-19 $X=4.34 $Y=0.805
c91 14 0 1.20958e-19 $X=4.29 $Y=2.055
c92 9 0 2.69181e-19 $X=3.62 $Y=2.885
r93 32 33 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.965 $Y=2.57
+ $X2=5.965 $Y2=2.405
r94 28 30 5.28824 $w=1.75e-07 $l=9.24662e-08 $layer=LI1_cond $X=5.92 $Y=1.675
+ $X2=5.915 $Y2=1.585
r95 28 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.92 $Y=1.675
+ $X2=5.92 $Y2=2.405
r96 24 30 5.28824 $w=1.75e-07 $l=9e-08 $layer=LI1_cond $X=5.915 $Y=1.495
+ $X2=5.915 $Y2=1.585
r97 24 26 45.2879 $w=1.78e-07 $l=7.35e-07 $layer=LI1_cond $X=5.915 $Y=1.495
+ $X2=5.915 $Y2=0.76
r98 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.43
+ $Y=1.58 $X2=4.43 $Y2=1.58
r99 19 30 1.24132 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=5.825 $Y=1.585
+ $X2=5.915 $Y2=1.585
r100 19 21 85.9545 $w=1.78e-07 $l=1.395e-06 $layer=LI1_cond $X=5.825 $Y=1.585
+ $X2=4.43 $Y2=1.585
r101 15 22 38.8075 $w=3.52e-07 $l=1.94808e-07 $layer=POLY_cond $X=4.34 $Y=1.415
+ $X2=4.405 $Y2=1.58
r102 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.34 $Y=1.415
+ $X2=4.34 $Y2=0.805
r103 13 22 38.8075 $w=3.52e-07 $l=2.14942e-07 $layer=POLY_cond $X=4.29 $Y=1.745
+ $X2=4.405 $Y2=1.58
r104 13 14 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=4.29 $Y=1.745
+ $X2=4.29 $Y2=2.055
r105 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.215 $Y=2.13
+ $X2=4.29 $Y2=2.055
r106 11 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=4.215 $Y=2.13
+ $X2=3.695 $Y2=2.13
r107 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.62 $Y=2.205
+ $X2=3.695 $Y2=2.13
r108 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.62 $Y=2.205
+ $X2=3.62 $Y2=2.885
r109 2 32 600 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=2.255 $X2=5.97 $Y2=2.57
r110 1 26 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=5.77
+ $Y=0.315 $X2=5.91 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%RESET_B 2 3 4 7 11 13 15 17 19 23 25 28 32
+ 36 38 40 44 47 48 54 55 56 58 60 61 62 65 67 70 71 73 74
c228 71 0 1.88119e-19 $X=8.2 $Y=1.83
c229 44 0 8.34918e-21 $X=8.2 $Y=1.815
c230 40 0 1.58556e-19 $X=4.895 $Y=1.215
c231 38 0 4.28297e-20 $X=2.34 $Y=0.18
c232 36 0 1.05727e-20 $X=1.93 $Y=2.195
c233 11 0 6.16896e-20 $X=2.34 $Y=0.6
c234 2 0 3.56339e-19 $X=1.68 $Y=2.12
r235 71 78 1.30009 $w=4.58e-07 $l=5e-08 $layer=LI1_cond $X=8.265 $Y=1.83
+ $X2=8.265 $Y2=1.88
r236 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.2
+ $Y=1.83 $X2=8.2 $Y2=1.83
r237 67 78 4.03026 $w=4.58e-07 $l=1.55e-07 $layer=LI1_cond $X=8.265 $Y=2.035
+ $X2=8.265 $Y2=1.88
r238 63 65 13.0115 $w=3.08e-07 $l=3.5e-07 $layer=LI1_cond $X=6.95 $Y=2.45
+ $X2=7.3 $Y2=2.45
r239 61 78 3.85449 $w=2.7e-07 $l=2.3e-07 $layer=LI1_cond $X=8.035 $Y=1.88
+ $X2=8.265 $Y2=1.88
r240 61 62 27.744 $w=2.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.035 $Y=1.88
+ $X2=7.385 $Y2=1.88
r241 60 65 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.3 $Y=2.295
+ $X2=7.3 $Y2=2.45
r242 59 62 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.3 $Y=2.015
+ $X2=7.385 $Y2=1.88
r243 59 60 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.3 $Y=2.015
+ $X2=7.3 $Y2=2.295
r244 57 63 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=6.95 $Y=2.605
+ $X2=6.95 $Y2=2.45
r245 57 58 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.95 $Y=2.605
+ $X2=6.95 $Y2=2.905
r246 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.865 $Y=2.99
+ $X2=6.95 $Y2=2.905
r247 55 56 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=6.865 $Y=2.99
+ $X2=5.665 $Y2=2.99
r248 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.58 $Y=2.905
+ $X2=5.665 $Y2=2.99
r249 53 54 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.58 $Y=2.565
+ $X2=5.58 $Y2=2.905
r250 51 74 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.76 $Y=2.4
+ $X2=4.91 $Y2=2.4
r251 51 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.76 $Y=2.4
+ $X2=4.595 $Y2=2.4
r252 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.76
+ $Y=2.4 $X2=4.76 $Y2=2.4
r253 48 53 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.495 $Y=2.4
+ $X2=5.58 $Y2=2.565
r254 48 50 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=5.495 $Y=2.4
+ $X2=4.76 $Y2=2.4
r255 46 70 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.2 $Y=2.17 $X2=8.2
+ $Y2=1.83
r256 46 47 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.2 $Y=2.17
+ $X2=8.2 $Y2=2.335
r257 44 70 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.2 $Y=1.815
+ $X2=8.2 $Y2=1.83
r258 41 44 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.89 $Y=1.74
+ $X2=8.2 $Y2=1.74
r259 39 40 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.895 $Y=1.065
+ $X2=4.895 $Y2=1.215
r260 34 36 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.68 $Y=2.195
+ $X2=1.93 $Y2=2.195
r261 32 47 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=8.22 $Y=2.885
+ $X2=8.22 $Y2=2.335
r262 26 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.89 $Y=1.665
+ $X2=7.89 $Y2=1.74
r263 26 28 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.89 $Y=1.665
+ $X2=7.89 $Y2=0.835
r264 25 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.91 $Y=2.235
+ $X2=4.91 $Y2=2.4
r265 25 40 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=4.91 $Y=2.235
+ $X2=4.91 $Y2=1.215
r266 23 39 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.88 $Y=0.745
+ $X2=4.88 $Y2=1.065
r267 20 23 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=4.88 $Y=0.255
+ $X2=4.88 $Y2=0.745
r268 19 73 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.15 $Y=2.49
+ $X2=4.595 $Y2=2.49
r269 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.075 $Y=2.565
+ $X2=4.15 $Y2=2.49
r270 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.075 $Y=2.565
+ $X2=4.075 $Y2=2.885
r271 14 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.415 $Y=0.18
+ $X2=2.34 $Y2=0.18
r272 13 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.805 $Y=0.18
+ $X2=4.88 $Y2=0.255
r273 13 14 1225.51 $w=1.5e-07 $l=2.39e-06 $layer=POLY_cond $X=4.805 $Y=0.18
+ $X2=2.415 $Y2=0.18
r274 9 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.34 $Y=0.255
+ $X2=2.34 $Y2=0.18
r275 9 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.34 $Y=0.255
+ $X2=2.34 $Y2=0.6
r276 5 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.93 $Y=2.27
+ $X2=1.93 $Y2=2.195
r277 5 7 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.93 $Y=2.27
+ $X2=1.93 $Y2=2.885
r278 3 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.265 $Y=0.18
+ $X2=2.34 $Y2=0.18
r279 3 4 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.265 $Y=0.18
+ $X2=1.755 $Y2=0.18
r280 2 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.68 $Y=2.12
+ $X2=1.68 $Y2=2.195
r281 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.68 $Y=0.255
+ $X2=1.755 $Y2=0.18
r282 1 2 956.309 $w=1.5e-07 $l=1.865e-06 $layer=POLY_cond $X=1.68 $Y=0.255
+ $X2=1.68 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%A_573_535# 1 2 3 11 12 14 17 19 24 25 26 29
+ 31 33 38 42 43 45 49
c126 43 0 1.772e-19 $X=5.48 $Y=1.93
c127 29 0 1.69354e-20 $X=3.765 $Y=0.805
c128 26 0 1.24911e-19 $X=3.585 $Y=2.07
r129 43 51 16.3698 $w=2.65e-07 $l=9e-08 $layer=POLY_cond $X=5.48 $Y=1.93
+ $X2=5.39 $Y2=1.93
r130 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.48
+ $Y=1.93 $X2=5.48 $Y2=1.93
r131 40 45 5.65194 $w=2.6e-07 $l=3.07002e-07 $layer=LI1_cond $X=4.455 $Y=1.955
+ $X2=4.165 $Y2=1.92
r132 40 42 53.6934 $w=2.18e-07 $l=1.025e-06 $layer=LI1_cond $X=4.455 $Y=1.955
+ $X2=5.48 $Y2=1.955
r133 36 45 0.952445 $w=2.9e-07 $l=3.65377e-07 $layer=LI1_cond $X=4.31 $Y=2.22
+ $X2=4.165 $Y2=1.92
r134 36 38 26.4267 $w=2.88e-07 $l=6.65e-07 $layer=LI1_cond $X=4.31 $Y=2.22
+ $X2=4.31 $Y2=2.885
r135 34 49 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.48 $Y=1.23
+ $X2=5.695 $Y2=1.23
r136 34 46 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.48 $Y=1.23 $X2=5.39
+ $Y2=1.23
r137 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.48
+ $Y=1.23 $X2=5.48 $Y2=1.23
r138 31 33 98.5859 $w=1.78e-07 $l=1.6e-06 $layer=LI1_cond $X=3.88 $Y=1.235
+ $X2=5.48 $Y2=1.235
r139 27 31 6.86909 $w=1.8e-07 $l=1.43091e-07 $layer=LI1_cond $X=3.775 $Y=1.145
+ $X2=3.88 $Y2=1.235
r140 27 29 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=3.775 $Y=1.145
+ $X2=3.775 $Y2=0.805
r141 25 45 5.65194 $w=2.6e-07 $l=1.5e-07 $layer=LI1_cond $X=4.165 $Y=2.07
+ $X2=4.165 $Y2=1.92
r142 25 26 22.2806 $w=2.98e-07 $l=5.8e-07 $layer=LI1_cond $X=4.165 $Y=2.07
+ $X2=3.585 $Y2=2.07
r143 23 26 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.5 $Y=2.22
+ $X2=3.585 $Y2=2.07
r144 23 24 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.5 $Y=2.22
+ $X2=3.5 $Y2=2.765
r145 19 24 7.39867 $w=2.85e-07 $l=1.79538e-07 $layer=LI1_cond $X=3.415 $Y=2.907
+ $X2=3.5 $Y2=2.765
r146 19 21 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.415 $Y=2.907
+ $X2=3.045 $Y2=2.907
r147 15 43 50.0189 $w=2.65e-07 $l=3.47851e-07 $layer=POLY_cond $X=5.755 $Y=2.095
+ $X2=5.48 $Y2=1.93
r148 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.755 $Y=2.095
+ $X2=5.755 $Y2=2.675
r149 12 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.065
+ $X2=5.695 $Y2=1.23
r150 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.695 $Y=1.065
+ $X2=5.695 $Y2=0.635
r151 11 51 16.0701 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.39 $Y=1.765
+ $X2=5.39 $Y2=1.93
r152 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.39 $Y=1.395
+ $X2=5.39 $Y2=1.23
r153 10 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.39 $Y=1.395
+ $X2=5.39 $Y2=1.765
r154 3 38 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.15
+ $Y=2.675 $X2=4.29 $Y2=2.885
r155 2 21 600 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_PDIFF $count=1 $X=2.865
+ $Y=2.675 $X2=3.045 $Y2=2.885
r156 1 29 182 $w=1.7e-07 $l=5.04182e-07 $layer=licon1_NDIFF $count=1 $X=3.355
+ $Y=0.595 $X2=3.765 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%A_1399_473# 1 2 9 12 15 17 21 23 25 26 28 30
+ 31 36 42
c117 31 0 1.30728e-19 $X=7.66 $Y=2.35
c118 30 0 8.34918e-21 $X=7.66 $Y=2.35
c119 28 0 5.67188e-20 $X=9.11 $Y=2.175
c120 12 0 2.53085e-19 $X=7.145 $Y=2.44
c121 9 0 1.10105e-19 $X=7.07 $Y=2.885
r122 41 42 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.46 $Y=2.35
+ $X2=7.385 $Y2=2.35
r123 36 38 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=8.465 $Y=0.835
+ $X2=8.465 $Y2=1.07
r124 31 41 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=7.66 $Y=2.35 $X2=7.46
+ $Y2=2.35
r125 30 33 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=7.7 $Y=2.35 $X2=7.7
+ $Y2=2.52
r126 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.66
+ $Y=2.35 $X2=7.66 $Y2=2.35
r127 27 28 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=9.11 $Y=1.155
+ $X2=9.11 $Y2=2.175
r128 26 40 20.6253 $w=2.57e-07 $l=4.84665e-07 $layer=LI1_cond $X=8.835 $Y=2.26
+ $X2=8.43 $Y2=2.435
r129 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.025 $Y=2.26
+ $X2=9.11 $Y2=2.175
r130 25 26 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.025 $Y=2.26
+ $X2=8.835 $Y2=2.26
r131 24 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.63 $Y=1.07
+ $X2=8.465 $Y2=1.07
r132 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.025 $Y=1.07
+ $X2=9.11 $Y2=1.155
r133 23 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.025 $Y=1.07
+ $X2=8.63 $Y2=1.07
r134 19 40 2.20825 $w=2e-07 $l=1.7e-07 $layer=LI1_cond $X=8.43 $Y=2.605 $X2=8.43
+ $Y2=2.435
r135 19 21 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=8.43 $Y=2.605
+ $X2=8.43 $Y2=2.885
r136 18 33 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.825 $Y=2.52
+ $X2=7.7 $Y2=2.52
r137 17 40 6.14668 $w=2.57e-07 $l=1.36015e-07 $layer=LI1_cond $X=8.33 $Y=2.52
+ $X2=8.43 $Y2=2.435
r138 17 18 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=8.33 $Y=2.52
+ $X2=7.825 $Y2=2.52
r139 13 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=2.185
+ $X2=7.46 $Y2=2.35
r140 13 15 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=7.46 $Y=2.185
+ $X2=7.46 $Y2=0.835
r141 12 42 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.145 $Y=2.44
+ $X2=7.385 $Y2=2.44
r142 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.07 $Y=2.515
+ $X2=7.145 $Y2=2.44
r143 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.07 $Y=2.515
+ $X2=7.07 $Y2=2.885
r144 2 21 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.295
+ $Y=2.675 $X2=8.435 $Y2=2.885
r145 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.325
+ $Y=0.625 $X2=8.465 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%A_1252_451# 1 2 9 11 12 15 17 21 24 27 31 33
+ 34 37 41 44 45 47 54 56 57 62 63
c148 57 0 1.25078e-19 $X=7.31 $Y=1.14
c149 54 0 2.76228e-19 $X=6.61 $Y=2.57
c150 44 0 1.64396e-19 $X=6.61 $Y=2.405
c151 21 0 5.33327e-20 $X=9.52 $Y=0.445
c152 12 0 1.88119e-19 $X=8.325 $Y=1.35
r153 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.77
+ $Y=1.49 $X2=8.77 $Y2=1.49
r154 57 59 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.31 $Y=1.14
+ $X2=7.31 $Y2=1.41
r155 52 54 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.4 $Y=2.57
+ $X2=6.61 $Y2=2.57
r156 48 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=1.41
+ $X2=7.31 $Y2=1.41
r157 47 62 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.685 $Y=1.41
+ $X2=8.77 $Y2=1.41
r158 47 48 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=8.685 $Y=1.41
+ $X2=7.395 $Y2=1.41
r159 46 56 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.775 $Y=1.14
+ $X2=6.65 $Y2=1.14
r160 45 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.225 $Y=1.14
+ $X2=7.31 $Y2=1.14
r161 45 46 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.225 $Y=1.14
+ $X2=6.775 $Y2=1.14
r162 44 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.61 $Y=2.405
+ $X2=6.61 $Y2=2.57
r163 43 56 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=6.61 $Y=1.225
+ $X2=6.65 $Y2=1.14
r164 43 44 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=6.61 $Y=1.225
+ $X2=6.61 $Y2=2.405
r165 39 56 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.65 $Y=1.055
+ $X2=6.65 $Y2=1.14
r166 39 41 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.65 $Y=1.055
+ $X2=6.65 $Y2=0.77
r167 35 37 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=9.52 $Y=1.83 $X2=9.6
+ $Y2=1.83
r168 32 63 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=8.77 $Y=1.425
+ $X2=8.77 $Y2=1.49
r169 32 33 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.77 $Y=1.425
+ $X2=8.77 $Y2=1.35
r170 30 63 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=8.77 $Y=1.845
+ $X2=8.77 $Y2=1.49
r171 30 31 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=8.755 $Y=1.845
+ $X2=8.755 $Y2=1.995
r172 25 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.6 $Y=1.905
+ $X2=9.6 $Y2=1.83
r173 25 27 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=9.6 $Y=1.905
+ $X2=9.6 $Y2=2.775
r174 24 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.52 $Y=1.755
+ $X2=9.52 $Y2=1.83
r175 23 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.52 $Y=1.425
+ $X2=9.52 $Y2=1.35
r176 23 24 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=9.52 $Y=1.425
+ $X2=9.52 $Y2=1.755
r177 19 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.52 $Y=1.275
+ $X2=9.52 $Y2=1.35
r178 19 21 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.52 $Y=1.275
+ $X2=9.52 $Y2=0.445
r179 18 33 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.935 $Y=1.35
+ $X2=8.77 $Y2=1.35
r180 17 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.445 $Y=1.35
+ $X2=9.52 $Y2=1.35
r181 17 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=9.445 $Y=1.35
+ $X2=8.935 $Y2=1.35
r182 15 31 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=8.65 $Y=2.885
+ $X2=8.65 $Y2=1.995
r183 11 33 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.605 $Y=1.35
+ $X2=8.77 $Y2=1.35
r184 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=8.605 $Y=1.35
+ $X2=8.325 $Y2=1.35
r185 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.25 $Y=1.275
+ $X2=8.325 $Y2=1.35
r186 7 9 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.25 $Y=1.275
+ $X2=8.25 $Y2=0.835
r187 2 52 600 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_PDIFF $count=1 $X=6.26
+ $Y=2.255 $X2=6.4 $Y2=2.57
r188 1 41 182 $w=1.7e-07 $l=5.60312e-07 $layer=licon1_NDIFF $count=1 $X=6.375
+ $Y=0.315 $X2=6.61 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%A_1836_47# 1 2 9 12 14 16 18 21 23 26 31 36
+ 41 44 45 46 47 48
c85 47 0 5.67188e-20 $X=9.995 $Y=1.26
r86 47 48 32.0796 $w=3.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.995 $Y=1.26
+ $X2=9.995 $Y2=1.185
r87 44 45 5.40936 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=9.387 $Y=2.61
+ $X2=9.387 $Y2=2.515
r88 37 50 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.995 $Y=1.35
+ $X2=9.995 $Y2=1.515
r89 37 47 13.1721 $w=3.8e-07 $l=9e-08 $layer=POLY_cond $X=9.995 $Y=1.35
+ $X2=9.995 $Y2=1.26
r90 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.97
+ $Y=1.35 $X2=9.97 $Y2=1.35
r91 34 46 0.718145 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=9.555 $Y=1.35
+ $X2=9.46 $Y2=1.35
r92 34 36 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=9.555 $Y=1.35
+ $X2=9.97 $Y2=1.35
r93 32 46 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.46 $Y=1.515
+ $X2=9.46 $Y2=1.35
r94 32 45 58.3732 $w=1.88e-07 $l=1e-06 $layer=LI1_cond $X=9.46 $Y=1.515 $X2=9.46
+ $Y2=2.515
r95 31 46 8.26956 $w=1.8e-07 $l=1.69926e-07 $layer=LI1_cond $X=9.45 $Y=1.185
+ $X2=9.46 $Y2=1.35
r96 30 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.45 $Y=0.815
+ $X2=9.45 $Y2=0.73
r97 30 31 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.45 $Y=0.815
+ $X2=9.45 $Y2=1.185
r98 24 41 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=9.27 $Y=0.73
+ $X2=9.45 $Y2=0.73
r99 24 26 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=9.27 $Y=0.645 $X2=9.27
+ $Y2=0.445
r100 19 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.54 $Y=1.335
+ $X2=10.54 $Y2=1.26
r101 19 21 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=10.54 $Y=1.335
+ $X2=10.54 $Y2=2.465
r102 16 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.54 $Y=1.185
+ $X2=10.54 $Y2=1.26
r103 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.54 $Y=1.185
+ $X2=10.54 $Y2=0.655
r104 15 47 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.185 $Y=1.26
+ $X2=9.995 $Y2=1.26
r105 14 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.465 $Y=1.26
+ $X2=10.54 $Y2=1.26
r106 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.465 $Y=1.26
+ $X2=10.185 $Y2=1.26
r107 12 50 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=10.11 $Y=2.465
+ $X2=10.11 $Y2=1.515
r108 9 48 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.11 $Y=0.655
+ $X2=10.11 $Y2=1.185
r109 2 44 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=9.26
+ $Y=2.455 $X2=9.385 $Y2=2.61
r110 1 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.18
+ $Y=0.235 $X2=9.305 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51 53
+ 58 59 61 62 63 65 70 95 100 105 111 114 119 122 124 127 131
r157 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r158 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r159 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r160 121 122 10.4169 $w=6.38e-07 $l=1.65e-07 $layer=LI1_cond $X=7.995 $Y=3.095
+ $X2=8.16 $Y2=3.095
r161 117 121 1.40165 $w=6.38e-07 $l=7.5e-08 $layer=LI1_cond $X=7.92 $Y=3.095
+ $X2=7.995 $Y2=3.095
r162 117 119 20.6957 $w=6.38e-07 $l=7.15e-07 $layer=LI1_cond $X=7.92 $Y=3.095
+ $X2=7.205 $Y2=3.095
r163 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r164 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r165 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r166 109 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r167 109 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r168 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r169 106 127 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=10.06 $Y=3.33
+ $X2=9.892 $Y2=3.33
r170 106 108 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=10.06 $Y=3.33
+ $X2=10.32 $Y2=3.33
r171 105 130 4.39729 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=10.625 $Y=3.33
+ $X2=10.832 $Y2=3.33
r172 105 108 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.625 $Y=3.33
+ $X2=10.32 $Y2=3.33
r173 104 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r174 104 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r175 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r176 101 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=8.865 $Y2=3.33
r177 101 103 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=9.36 $Y2=3.33
r178 100 127 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=9.725 $Y=3.33
+ $X2=9.892 $Y2=3.33
r179 100 103 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.725 $Y=3.33
+ $X2=9.36 $Y2=3.33
r180 99 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r181 99 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r182 98 122 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=8.16 $Y2=3.33
r183 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r184 95 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.7 $Y=3.33
+ $X2=8.865 $Y2=3.33
r185 95 98 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.7 $Y=3.33 $X2=8.4
+ $Y2=3.33
r186 94 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r187 93 119 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.205 $Y2=3.33
r188 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r189 90 93 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=6.96 $Y2=3.33
r190 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r191 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r192 83 86 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r193 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r194 81 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r195 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r196 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r197 78 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r198 77 80 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r199 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r200 75 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=3.33
+ $X2=2.145 $Y2=3.33
r201 75 77 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.31 $Y=3.33
+ $X2=2.64 $Y2=3.33
r202 74 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r203 74 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r204 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r205 71 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r206 71 73 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r207 70 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=3.33
+ $X2=2.145 $Y2=3.33
r208 70 73 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.98 $Y=3.33 $X2=1.68
+ $Y2=3.33
r209 68 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r210 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r211 65 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r212 65 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r213 63 94 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.96 $Y2=3.33
r214 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r215 63 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r216 61 86 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.065 $Y=3.33
+ $X2=5.04 $Y2=3.33
r217 61 62 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.065 $Y=3.33
+ $X2=5.195 $Y2=3.33
r218 60 90 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.325 $Y=3.33
+ $X2=5.52 $Y2=3.33
r219 60 62 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.325 $Y=3.33
+ $X2=5.195 $Y2=3.33
r220 58 80 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.6 $Y2=3.33
r221 58 59 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.875 $Y2=3.33
r222 57 83 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=3.33
+ $X2=4.08 $Y2=3.33
r223 57 59 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.995 $Y=3.33
+ $X2=3.875 $Y2=3.33
r224 53 56 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=10.772 $Y=1.98
+ $X2=10.772 $Y2=2.95
r225 51 130 3.08023 $w=2.95e-07 $l=1.11018e-07 $layer=LI1_cond $X=10.772
+ $Y=3.245 $X2=10.832 $Y2=3.33
r226 51 56 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=10.772 $Y=3.245
+ $X2=10.772 $Y2=2.95
r227 47 50 33.3692 $w=3.33e-07 $l=9.7e-07 $layer=LI1_cond $X=9.892 $Y=1.98
+ $X2=9.892 $Y2=2.95
r228 45 127 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=9.892 $Y=3.245
+ $X2=9.892 $Y2=3.33
r229 45 50 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=9.892 $Y=3.245
+ $X2=9.892 $Y2=2.95
r230 41 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.865 $Y=3.245
+ $X2=8.865 $Y2=3.33
r231 41 43 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=8.865 $Y=3.245
+ $X2=8.865 $Y2=2.885
r232 37 62 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.195 $Y=3.245
+ $X2=5.195 $Y2=3.33
r233 37 39 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=5.195 $Y=3.245
+ $X2=5.195 $Y2=2.9
r234 33 59 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=3.245
+ $X2=3.875 $Y2=3.33
r235 33 35 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=3.875 $Y=3.245
+ $X2=3.875 $Y2=2.885
r236 29 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=3.245
+ $X2=2.145 $Y2=3.33
r237 29 31 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.145 $Y=3.245
+ $X2=2.145 $Y2=2.885
r238 25 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r239 25 27 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.765
r240 8 56 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=10.615
+ $Y=1.835 $X2=10.755 $Y2=2.95
r241 8 53 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.615
+ $Y=1.835 $X2=10.755 $Y2=1.98
r242 7 50 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=9.675
+ $Y=2.455 $X2=9.815 $Y2=2.95
r243 7 47 300 $w=1.7e-07 $l=5.74565e-07 $layer=licon1_PDIFF $count=2 $X=9.675
+ $Y=2.455 $X2=9.895 $Y2=1.98
r244 6 43 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.725
+ $Y=2.675 $X2=8.865 $Y2=2.885
r245 5 121 300 $w=1.7e-07 $l=9.4921e-07 $layer=licon1_PDIFF $count=2 $X=7.145
+ $Y=2.675 $X2=7.995 $Y2=2.885
r246 4 39 600 $w=1.7e-07 $l=7.13828e-07 $layer=licon1_PDIFF $count=1 $X=5.085
+ $Y=2.255 $X2=5.23 $Y2=2.9
r247 3 35 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=3.695
+ $Y=2.675 $X2=3.86 $Y2=2.885
r248 2 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.005
+ $Y=2.675 $X2=2.145 $Y2=2.885
r249 1 27 600 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.32 $X2=0.69 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%A_318_535# 1 2 3 12 14 15 18 20 23 25 26 30
+ 34
c84 34 0 3.77105e-19 $X=3.16 $Y=1.65
c85 20 0 1.4427e-19 $X=3.075 $Y=2.51
r86 32 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.87 $Y=1.65
+ $X2=3.16 $Y2=1.65
r87 27 30 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.87 $Y=0.805
+ $X2=3.065 $Y2=0.805
r88 24 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=1.735
+ $X2=3.16 $Y2=1.65
r89 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.16 $Y=1.735
+ $X2=3.16 $Y2=2.425
r90 23 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.565
+ $X2=2.87 $Y2=1.65
r91 22 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=0.97
+ $X2=2.87 $Y2=0.805
r92 22 23 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.87 $Y=0.97
+ $X2=2.87 $Y2=1.565
r93 21 26 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.7 $Y=2.51 $X2=2.59
+ $Y2=2.51
r94 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.075 $Y=2.51
+ $X2=3.16 $Y2=2.425
r95 20 21 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.075 $Y=2.51
+ $X2=2.7 $Y2=2.51
r96 16 26 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=2.595
+ $X2=2.59 $Y2=2.51
r97 16 18 15.1913 $w=2.18e-07 $l=2.9e-07 $layer=LI1_cond $X=2.59 $Y=2.595
+ $X2=2.59 $Y2=2.885
r98 14 26 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.48 $Y=2.51 $X2=2.59
+ $Y2=2.51
r99 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.48 $Y=2.51
+ $X2=1.81 $Y2=2.51
r100 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.68 $Y=2.595
+ $X2=1.81 $Y2=2.51
r101 10 12 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=2.595
+ $X2=1.68 $Y2=2.885
r102 3 18 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=2.675 $X2=2.575 $Y2=2.885
r103 2 12 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=2.675 $X2=1.715 $Y2=2.885
r104 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.925
+ $Y=0.595 $X2=3.065 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%Q 1 2 7 8 9 10 11 12 13 22
c18 22 0 5.33327e-20 $X=10.325 $Y=0.42
r19 13 40 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=10.342 $Y=2.775
+ $X2=10.342 $Y2=2.91
r20 12 13 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=10.342 $Y=2.405
+ $X2=10.342 $Y2=2.775
r21 11 12 19.9757 $w=2.23e-07 $l=3.9e-07 $layer=LI1_cond $X=10.342 $Y=2.015
+ $X2=10.342 $Y2=2.405
r22 10 11 17.9269 $w=2.23e-07 $l=3.5e-07 $layer=LI1_cond $X=10.342 $Y=1.665
+ $X2=10.342 $Y2=2.015
r23 9 10 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=10.342 $Y=1.295
+ $X2=10.342 $Y2=1.665
r24 8 9 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=10.342 $Y=0.925
+ $X2=10.342 $Y2=1.295
r25 7 8 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=10.342 $Y=0.555
+ $X2=10.342 $Y2=0.925
r26 7 22 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=10.342 $Y=0.555
+ $X2=10.342 $Y2=0.42
r27 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.185
+ $Y=1.835 $X2=10.325 $Y2=2.91
r28 2 11 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=10.185
+ $Y=1.835 $X2=10.325 $Y2=2.015
r29 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=10.185
+ $Y=0.235 $X2=10.325 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_2%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 47 48 49 51 56 71 78 84 87 91 98
r120 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r121 94 95 3.73559 $w=4.88e-07 $l=1.15e-07 $layer=LI1_cond $X=9.815 $Y=0.36
+ $X2=9.815 $Y2=0.475
r122 91 94 8.78751 $w=4.88e-07 $l=3.6e-07 $layer=LI1_cond $X=9.815 $Y=0
+ $X2=9.815 $Y2=0.36
r123 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r124 87 88 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r125 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r126 82 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r127 82 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r128 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r129 79 91 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=10.06 $Y=0
+ $X2=9.815 $Y2=0
r130 79 81 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=10.06 $Y=0
+ $X2=10.32 $Y2=0
r131 78 97 4.39729 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=10.625 $Y=0
+ $X2=10.832 $Y2=0
r132 78 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.625 $Y=0
+ $X2=10.32 $Y2=0
r133 77 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r134 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r135 74 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.36 $Y2=0
r136 73 76 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.36
+ $Y2=0
r137 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r138 71 91 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=9.57 $Y=0 $X2=9.815
+ $Y2=0
r139 71 76 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.57 $Y=0 $X2=9.36
+ $Y2=0
r140 70 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r141 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r142 66 69 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r143 64 88 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=2.16 $Y2=0
r144 63 64 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r145 61 87 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.117
+ $Y2=0
r146 61 63 182.674 $w=1.68e-07 $l=2.8e-06 $layer=LI1_cond $X=2.24 $Y=0 $X2=5.04
+ $Y2=0
r147 60 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r148 60 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r149 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r150 57 84 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.785 $Y=0
+ $X2=0.672 $Y2=0
r151 57 59 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=0.785 $Y=0
+ $X2=1.68 $Y2=0
r152 56 87 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=1.995 $Y=0
+ $X2=2.117 $Y2=0
r153 56 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=0
+ $X2=1.68 $Y2=0
r154 54 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r155 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r156 51 84 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.672
+ $Y2=0
r157 51 53 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r158 49 70 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=7.44 $Y2=0
r159 49 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r160 49 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r161 47 69 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=7.51 $Y=0 $X2=7.44
+ $Y2=0
r162 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.51 $Y=0 $X2=7.675
+ $Y2=0
r163 46 73 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.84 $Y=0 $X2=7.92
+ $Y2=0
r164 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.84 $Y=0 $X2=7.675
+ $Y2=0
r165 44 63 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.045 $Y=0 $X2=5.04
+ $Y2=0
r166 44 45 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.045 $Y=0 $X2=5.18
+ $Y2=0
r167 43 66 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.315 $Y=0
+ $X2=5.52 $Y2=0
r168 43 45 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.18
+ $Y2=0
r169 39 97 3.08023 $w=2.95e-07 $l=1.11018e-07 $layer=LI1_cond $X=10.772 $Y=0.085
+ $X2=10.832 $Y2=0
r170 39 41 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=10.772 $Y=0.085
+ $X2=10.772 $Y2=0.38
r171 37 95 13.9592 $w=3.53e-07 $l=4.3e-07 $layer=LI1_cond $X=9.882 $Y=0.905
+ $X2=9.882 $Y2=0.475
r172 31 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.675 $Y=0.085
+ $X2=7.675 $Y2=0
r173 31 33 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=7.675 $Y=0.085
+ $X2=7.675 $Y2=0.785
r174 27 45 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=0.085
+ $X2=5.18 $Y2=0
r175 27 29 16.433 $w=2.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.18 $Y=0.085
+ $X2=5.18 $Y2=0.47
r176 23 87 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.117 $Y=0.085
+ $X2=2.117 $Y2=0
r177 23 25 21.1673 $w=2.43e-07 $l=4.5e-07 $layer=LI1_cond $X=2.117 $Y=0.085
+ $X2=2.117 $Y2=0.535
r178 19 84 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.672 $Y=0.085
+ $X2=0.672 $Y2=0
r179 19 21 32.2684 $w=2.23e-07 $l=6.3e-07 $layer=LI1_cond $X=0.672 $Y=0.085
+ $X2=0.672 $Y2=0.715
r180 6 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.615
+ $Y=0.235 $X2=10.755 $Y2=0.38
r181 5 94 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=9.595
+ $Y=0.235 $X2=9.735 $Y2=0.36
r182 5 37 182 $w=1.7e-07 $l=8.06164e-07 $layer=licon1_NDIFF $count=1 $X=9.595
+ $Y=0.235 $X2=9.895 $Y2=0.905
r183 4 33 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.535
+ $Y=0.625 $X2=7.675 $Y2=0.785
r184 3 29 182 $w=1.7e-07 $l=2.85657e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.535 $X2=5.21 $Y2=0.47
r185 2 25 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.39 $X2=2.125 $Y2=0.535
r186 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.505 $X2=0.69 $Y2=0.715
.ends

