* File: sky130_fd_sc_lp__a221oi_1.spice
* Created: Fri Aug 28 09:53:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a221oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a221oi_1  VNB VPB C1 B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_C1_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2667 AS=0.2226 PD=1.475 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1001 A_300_47# N_B2_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.2667 PD=1.05 PS=1.475 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g A_300_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=7.848 NRS=7.14 M=1 R=5.6 SA=75001.3 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1005 A_480_47# N_A1_M1005_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.1638 PD=1.23 PS=1.23 NRD=19.992 NRS=7.848 M=1 R=5.6 SA=75001.9 SB=75000.7
+ A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g A_480_47# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6 SA=75002.4 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1009 N_A_110_367#_M1009_d N_C1_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1004 N_A_110_367#_M1004_d N_B2_M1004_g N_A_217_367#_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.189 AS=0.3339 PD=1.56 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1006 N_A_217_367#_M1006_d N_B1_M1006_g N_A_110_367#_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2079 AS=0.189 PD=1.59 PS=1.56 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75000.6 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_217_367#_M1006_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.2079 PD=1.62 PS=1.59 NRD=5.4569 NRS=7.8012 M=1 R=8.4
+ SA=75001.1 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1002 N_A_217_367#_M1002_d N_A2_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2268 PD=3.05 PS=1.62 NRD=0 NRS=7.0329 M=1 R=8.4
+ SA=75001.6 SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a221oi_1.pxi.spice"
*
.ends
*
*
