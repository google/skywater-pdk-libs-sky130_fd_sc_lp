* File: sky130_fd_sc_lp__a22o_4.pex.spice
* Created: Wed Sep  2 09:22:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22O_4%A_103_263# 1 2 3 4 15 19 23 27 31 35 39 43 45
+ 54 56 57 58 61 62 65 69 71 73 75 89
c156 71 0 1.14977e-19 $X=3.3 $Y=2.12
c157 43 0 1.4432e-19 $X=2.58 $Y=0.655
r158 86 87 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.13 $Y=1.48 $X2=2.15
+ $Y2=1.48
r159 85 86 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.72 $Y=1.48
+ $X2=2.13 $Y2=1.48
r160 84 85 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.7 $Y=1.48 $X2=1.72
+ $Y2=1.48
r161 83 84 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.29 $Y=1.48
+ $X2=1.7 $Y2=1.48
r162 82 83 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.27 $Y=1.48 $X2=1.29
+ $Y2=1.48
r163 81 82 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.84 $Y=1.48
+ $X2=1.27 $Y2=1.48
r164 75 77 2.46952 $w=2.78e-07 $l=6e-08 $layer=LI1_cond $X=5.625 $Y=0.865
+ $X2=5.625 $Y2=0.925
r165 66 71 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.395 $Y=2.045
+ $X2=3.3 $Y2=2.045
r166 65 73 3.89832 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=4.065 $Y=2.045
+ $X2=4.18 $Y2=2.045
r167 65 66 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.065 $Y=2.045
+ $X2=3.395 $Y2=2.045
r168 61 71 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.205 $Y=2.045
+ $X2=3.3 $Y2=2.045
r169 61 62 24.9545 $w=1.78e-07 $l=4.05e-07 $layer=LI1_cond $X=3.205 $Y=2.045
+ $X2=2.8 $Y2=2.045
r170 58 60 49.1169 $w=2.08e-07 $l=9.3e-07 $layer=LI1_cond $X=2.8 $Y=0.925
+ $X2=3.73 $Y2=0.925
r171 57 77 2.424 $w=2.1e-07 $l=1.4e-07 $layer=LI1_cond $X=5.485 $Y=0.925
+ $X2=5.625 $Y2=0.925
r172 57 60 92.6883 $w=2.08e-07 $l=1.755e-06 $layer=LI1_cond $X=5.485 $Y=0.925
+ $X2=3.73 $Y2=0.925
r173 56 62 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.715 $Y=1.955
+ $X2=2.8 $Y2=2.045
r174 55 69 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.715 $Y=1.585
+ $X2=2.715 $Y2=1.485
r175 55 56 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.715 $Y=1.585
+ $X2=2.715 $Y2=1.955
r176 54 69 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.715 $Y=1.385
+ $X2=2.715 $Y2=1.485
r177 53 58 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.715 $Y=1.03
+ $X2=2.8 $Y2=0.925
r178 53 54 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.715 $Y=1.03
+ $X2=2.715 $Y2=1.385
r179 52 89 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=2.38 $Y=1.48 $X2=2.58
+ $Y2=1.48
r180 52 87 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.38 $Y=1.48
+ $X2=2.15 $Y2=1.48
r181 51 52 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.38
+ $Y=1.48 $X2=2.38 $Y2=1.48
r182 48 81 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.68 $Y=1.48
+ $X2=0.84 $Y2=1.48
r183 47 51 94.2727 $w=1.98e-07 $l=1.7e-06 $layer=LI1_cond $X=0.68 $Y=1.485
+ $X2=2.38 $Y2=1.485
r184 47 48 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=0.68
+ $Y=1.48 $X2=0.68 $Y2=1.48
r185 45 69 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=1.485
+ $X2=2.715 $Y2=1.485
r186 45 51 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=2.63 $Y=1.485
+ $X2=2.38 $Y2=1.485
r187 41 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.315
+ $X2=2.58 $Y2=1.48
r188 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.58 $Y=1.315
+ $X2=2.58 $Y2=0.655
r189 37 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.315
+ $X2=2.15 $Y2=1.48
r190 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.315
+ $X2=2.15 $Y2=0.655
r191 33 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.645
+ $X2=2.13 $Y2=1.48
r192 33 35 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.13 $Y=1.645
+ $X2=2.13 $Y2=2.465
r193 29 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.72 $Y=1.315
+ $X2=1.72 $Y2=1.48
r194 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.72 $Y=1.315
+ $X2=1.72 $Y2=0.655
r195 25 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.645
+ $X2=1.7 $Y2=1.48
r196 25 27 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.7 $Y=1.645
+ $X2=1.7 $Y2=2.465
r197 21 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.315
+ $X2=1.29 $Y2=1.48
r198 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.29 $Y=1.315
+ $X2=1.29 $Y2=0.655
r199 17 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.27 $Y=1.645
+ $X2=1.27 $Y2=1.48
r200 17 19 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.27 $Y=1.645
+ $X2=1.27 $Y2=2.465
r201 13 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.645
+ $X2=0.84 $Y2=1.48
r202 13 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.84 $Y=1.645
+ $X2=0.84 $Y2=2.465
r203 4 73 300 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=2 $X=4.02
+ $Y=1.835 $X2=4.16 $Y2=2.13
r204 3 71 300 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=2 $X=3.16
+ $Y=1.835 $X2=3.3 $Y2=2.12
r205 2 75 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.235 $X2=5.6 $Y2=0.865
r206 1 60 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.235 $X2=3.73 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%B2 3 7 11 15 17 20 21 25 28 29
c88 29 0 1.30656e-19 $X=3.065 $Y=1.51
c89 28 0 1.14977e-19 $X=3.065 $Y=1.51
c90 20 0 1.30739e-19 $X=4.395 $Y=1.51
c91 11 0 1.15476e-19 $X=4.375 $Y=0.655
r92 28 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.51
+ $X2=3.065 $Y2=1.675
r93 28 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.51
+ $X2=3.065 $Y2=1.345
r94 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.065
+ $Y=1.51 $X2=3.065 $Y2=1.51
r95 25 39 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=3.1 $Y=1.665 $X2=3.1
+ $Y2=1.7
r96 25 29 6.87033 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=3.1 $Y=1.665
+ $X2=3.1 $Y2=1.51
r97 21 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.51
+ $X2=4.395 $Y2=1.675
r98 21 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.51
+ $X2=4.395 $Y2=1.345
r99 20 23 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.395 $Y=1.51
+ $X2=4.395 $Y2=1.7
r100 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=1.51 $X2=4.395 $Y2=1.51
r101 18 39 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.23 $Y=1.7 $X2=3.1
+ $Y2=1.7
r102 17 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=1.7
+ $X2=4.395 $Y2=1.7
r103 17 18 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=4.23 $Y=1.7 $X2=3.23
+ $Y2=1.7
r104 15 34 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.375 $Y=2.465
+ $X2=4.375 $Y2=1.675
r105 11 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.375 $Y=0.655
+ $X2=4.375 $Y2=1.345
r106 7 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.085 $Y=2.465
+ $X2=3.085 $Y2=1.675
r107 3 30 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.085 $Y=0.655
+ $X2=3.085 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%B1 1 3 6 8 10 13 15 21 22
c51 13 0 1.30739e-19 $X=3.945 $Y=2.465
c52 6 0 1.30656e-19 $X=3.515 $Y=2.465
r53 20 22 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.72 $Y=1.35
+ $X2=3.945 $Y2=1.35
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.72
+ $Y=1.35 $X2=3.72 $Y2=1.35
r55 17 20 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.515 $Y=1.35
+ $X2=3.72 $Y2=1.35
r56 15 21 5.64462 $w=2.43e-07 $l=1.2e-07 $layer=LI1_cond $X=3.6 $Y=1.322
+ $X2=3.72 $Y2=1.322
r57 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.515
+ $X2=3.945 $Y2=1.35
r58 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.945 $Y=1.515
+ $X2=3.945 $Y2=2.465
r59 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.185
+ $X2=3.945 $Y2=1.35
r60 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.945 $Y=1.185
+ $X2=3.945 $Y2=0.655
r61 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.515 $Y=1.515
+ $X2=3.515 $Y2=1.35
r62 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.515 $Y=1.515
+ $X2=3.515 $Y2=2.465
r63 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.515 $Y=1.185
+ $X2=3.515 $Y2=1.35
r64 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.515 $Y=1.185
+ $X2=3.515 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%A2 3 7 11 15 17 20 21 25 26 36 39
c69 20 0 1.53398e-19 $X=4.935 $Y=1.51
r70 33 36 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.245 $Y=1.375
+ $X2=6.45 $Y2=1.375
r71 26 39 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=1.7 $X2=6.45
+ $Y2=1.615
r72 26 39 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=6.45 $Y=1.597
+ $X2=6.45 $Y2=1.615
r73 25 26 10.5466 $w=3.28e-07 $l=3.02e-07 $layer=LI1_cond $X=6.45 $Y=1.295
+ $X2=6.45 $Y2=1.597
r74 25 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.375 $X2=6.45 $Y2=1.375
r75 21 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.51
+ $X2=4.935 $Y2=1.675
r76 21 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.51
+ $X2=4.935 $Y2=1.345
r77 20 23 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.935 $Y=1.51
+ $X2=4.935 $Y2=1.7
r78 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.51 $X2=4.935 $Y2=1.51
r79 18 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.1 $Y=1.7 $X2=4.935
+ $Y2=1.7
r80 17 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.285 $Y=1.7
+ $X2=6.45 $Y2=1.7
r81 17 18 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=6.285 $Y=1.7
+ $X2=5.1 $Y2=1.7
r82 13 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.54
+ $X2=6.245 $Y2=1.375
r83 13 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=6.245 $Y=1.54
+ $X2=6.245 $Y2=2.465
r84 9 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.21
+ $X2=6.245 $Y2=1.375
r85 9 11 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.245 $Y=1.21
+ $X2=6.245 $Y2=0.655
r86 7 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.955 $Y=0.655
+ $X2=4.955 $Y2=1.345
r87 3 32 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.875 $Y=2.465
+ $X2=4.875 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%A1 1 3 6 8 10 13 15 16 24
c49 6 0 1.53398e-19 $X=5.385 $Y=2.465
r50 22 24 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=5.595 $Y=1.35
+ $X2=5.815 $Y2=1.35
r51 19 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.385 $Y=1.35
+ $X2=5.595 $Y2=1.35
r52 15 16 22.5785 $w=2.43e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.322 $X2=6
+ $Y2=1.322
r53 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.595
+ $Y=1.35 $X2=5.595 $Y2=1.35
r54 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.515
+ $X2=5.815 $Y2=1.35
r55 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.815 $Y=1.515
+ $X2=5.815 $Y2=2.465
r56 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.185
+ $X2=5.815 $Y2=1.35
r57 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.815 $Y=1.185
+ $X2=5.815 $Y2=0.655
r58 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.515
+ $X2=5.385 $Y2=1.35
r59 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.385 $Y=1.515
+ $X2=5.385 $Y2=2.465
r60 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.185
+ $X2=5.385 $Y2=1.35
r61 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.385 $Y=1.185
+ $X2=5.385 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%VPWR 1 2 3 4 5 18 24 30 36 40 43 44 46 47 49
+ 50 51 63 67 74 75 78 81
r95 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r96 78 79 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r97 75 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r98 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r99 72 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=6.03 $Y2=3.33
r100 72 74 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 71 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r102 71 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r104 68 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.295 $Y=3.33
+ $X2=5.13 $Y2=3.33
r105 68 70 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.295 $Y=3.33
+ $X2=5.52 $Y2=3.33
r106 67 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=3.33
+ $X2=6.03 $Y2=3.33
r107 67 70 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.865 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 65 66 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 63 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.965 $Y=3.33
+ $X2=5.13 $Y2=3.33
r110 63 65 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=4.965 $Y=3.33
+ $X2=2.64 $Y2=3.33
r111 62 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r113 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r114 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 55 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r116 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r117 51 79 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=5.04 $Y2=3.33
r118 51 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 49 61 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.22 $Y=3.33 $X2=2.16
+ $Y2=3.33
r120 49 50 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.22 $Y=3.33
+ $X2=2.34 $Y2=3.33
r121 48 65 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.46 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 48 50 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.46 $Y=3.33
+ $X2=2.34 $Y2=3.33
r123 46 58 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.485 $Y2=3.33
r125 45 61 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=1.485 $Y2=3.33
r127 43 54 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.24 $Y2=3.33
r128 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.625 $Y2=3.33
r129 42 58 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.79 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=3.33
+ $X2=0.625 $Y2=3.33
r131 38 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=3.245
+ $X2=6.03 $Y2=3.33
r132 38 40 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=6.03 $Y=3.245
+ $X2=6.03 $Y2=2.38
r133 34 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.13 $Y=3.245
+ $X2=5.13 $Y2=3.33
r134 34 36 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=5.13 $Y=3.245
+ $X2=5.13 $Y2=2.38
r135 30 33 46.5779 $w=2.38e-07 $l=9.7e-07 $layer=LI1_cond $X=2.34 $Y=1.98
+ $X2=2.34 $Y2=2.95
r136 28 50 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=3.245
+ $X2=2.34 $Y2=3.33
r137 28 33 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.34 $Y=3.245
+ $X2=2.34 $Y2=2.95
r138 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.485 $Y=2.18
+ $X2=1.485 $Y2=2.95
r139 22 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=3.245
+ $X2=1.485 $Y2=3.33
r140 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.485 $Y=3.245
+ $X2=1.485 $Y2=2.95
r141 18 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.625 $Y=2.18
+ $X2=0.625 $Y2=2.95
r142 16 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.625 $Y=3.245
+ $X2=0.625 $Y2=3.33
r143 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.625 $Y=3.245
+ $X2=0.625 $Y2=2.95
r144 5 40 300 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=2 $X=5.89
+ $Y=1.835 $X2=6.03 $Y2=2.38
r145 4 36 300 $w=1.7e-07 $l=6.2859e-07 $layer=licon1_PDIFF $count=2 $X=4.95
+ $Y=1.835 $X2=5.13 $Y2=2.38
r146 3 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.205
+ $Y=1.835 $X2=2.345 $Y2=2.95
r147 3 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.205
+ $Y=1.835 $X2=2.345 $Y2=1.98
r148 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=1.835 $X2=1.485 $Y2=2.95
r149 2 24 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=1.835 $X2=1.485 $Y2=2.18
r150 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.5
+ $Y=1.835 $X2=0.625 $Y2=2.95
r151 1 18 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.5
+ $Y=1.835 $X2=0.625 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%X 1 2 3 4 13 14 15 19 23 27 29 33 39 42 43 44
+ 45 46 47 61
r60 59 61 3.76308 $w=2.43e-07 $l=8e-08 $layer=LI1_cond $X=0.222 $Y=1.215
+ $X2=0.222 $Y2=1.295
r61 46 53 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.262 $Y=1.13
+ $X2=0.262 $Y2=1.045
r62 46 59 3.29812 $w=2.85e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.262 $Y=1.13
+ $X2=0.222 $Y2=1.215
r63 46 47 17.3102 $w=2.43e-07 $l=3.68e-07 $layer=LI1_cond $X=0.222 $Y=1.297
+ $X2=0.222 $Y2=1.665
r64 46 61 0.094077 $w=2.43e-07 $l=2e-09 $layer=LI1_cond $X=0.222 $Y=1.297
+ $X2=0.222 $Y2=1.295
r65 45 53 4.25517 $w=3.23e-07 $l=1.2e-07 $layer=LI1_cond $X=0.262 $Y=0.925
+ $X2=0.262 $Y2=1.045
r66 44 45 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.262 $Y=0.555
+ $X2=0.262 $Y2=0.925
r67 41 47 4.23346 $w=2.43e-07 $l=9e-08 $layer=LI1_cond $X=0.222 $Y=1.755
+ $X2=0.222 $Y2=1.665
r68 37 39 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=2.365 $Y=1.045
+ $X2=2.365 $Y2=0.42
r69 33 35 46.5988 $w=2.28e-07 $l=9.3e-07 $layer=LI1_cond $X=1.935 $Y=1.98
+ $X2=1.935 $Y2=2.91
r70 31 33 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.935 $Y=1.925
+ $X2=1.935 $Y2=1.98
r71 30 43 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.59 $Y=1.13 $X2=1.5
+ $Y2=1.13
r72 29 37 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.27 $Y=1.13
+ $X2=2.365 $Y2=1.045
r73 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.27 $Y=1.13
+ $X2=1.59 $Y2=1.13
r74 25 43 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=1.045 $X2=1.5
+ $Y2=1.13
r75 25 27 38.5101 $w=1.78e-07 $l=6.25e-07 $layer=LI1_cond $X=1.5 $Y=1.045
+ $X2=1.5 $Y2=0.42
r76 24 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.15 $Y=1.84
+ $X2=1.055 $Y2=1.84
r77 23 31 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.82 $Y=1.84
+ $X2=1.935 $Y2=1.925
r78 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.82 $Y=1.84
+ $X2=1.15 $Y2=1.84
r79 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.055 $Y=1.98
+ $X2=1.055 $Y2=2.91
r80 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=1.925
+ $X2=1.055 $Y2=1.84
r81 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.055 $Y=1.925
+ $X2=1.055 $Y2=1.98
r82 16 46 3.25423 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=0.425 $Y=1.13
+ $X2=0.262 $Y2=1.13
r83 15 43 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.41 $Y=1.13 $X2=1.5
+ $Y2=1.13
r84 15 16 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=1.41 $Y=1.13
+ $X2=0.425 $Y2=1.13
r85 14 41 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.345 $Y=1.84
+ $X2=0.222 $Y2=1.755
r86 13 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.96 $Y=1.84
+ $X2=1.055 $Y2=1.84
r87 13 14 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.96 $Y=1.84
+ $X2=0.345 $Y2=1.84
r88 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.775
+ $Y=1.835 $X2=1.915 $Y2=2.91
r89 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.775
+ $Y=1.835 $X2=1.915 $Y2=1.98
r90 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.915
+ $Y=1.835 $X2=1.055 $Y2=2.91
r91 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.915
+ $Y=1.835 $X2=1.055 $Y2=1.98
r92 2 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.225
+ $Y=0.235 $X2=2.365 $Y2=0.42
r93 1 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.365
+ $Y=0.235 $X2=1.505 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%A_549_367# 1 2 3 4 5 18 20 21 24 26 28 32 36
+ 38 40 42 44 48
r65 40 50 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.495 $Y=2.125
+ $X2=6.495 $Y2=2.04
r66 40 42 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=6.495 $Y=2.125
+ $X2=6.495 $Y2=2.91
r67 39 48 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.695 $Y=2.04
+ $X2=5.58 $Y2=2.04
r68 38 50 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.365 $Y=2.04
+ $X2=6.495 $Y2=2.04
r69 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.365 $Y=2.04
+ $X2=5.695 $Y2=2.04
r70 34 48 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=2.125
+ $X2=5.58 $Y2=2.04
r71 34 36 39.3334 $w=2.28e-07 $l=7.85e-07 $layer=LI1_cond $X=5.58 $Y=2.125
+ $X2=5.58 $Y2=2.91
r72 33 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=2.04
+ $X2=4.63 $Y2=2.04
r73 32 48 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.465 $Y=2.04
+ $X2=5.58 $Y2=2.04
r74 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.465 $Y=2.04
+ $X2=4.795 $Y2=2.04
r75 29 31 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.63 $Y=2.905
+ $X2=4.63 $Y2=2.48
r76 28 46 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=2.125 $X2=4.63
+ $Y2=2.04
r77 28 31 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.63 $Y=2.125
+ $X2=4.63 $Y2=2.48
r78 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=2.99
+ $X2=3.73 $Y2=2.99
r79 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.465 $Y=2.99
+ $X2=4.63 $Y2=2.905
r80 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.465 $Y=2.99
+ $X2=3.895 $Y2=2.99
r81 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=2.905
+ $X2=3.73 $Y2=2.99
r82 22 24 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=3.73 $Y=2.905
+ $X2=3.73 $Y2=2.39
r83 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.565 $Y=2.99
+ $X2=3.73 $Y2=2.99
r84 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.565 $Y=2.99
+ $X2=3.035 $Y2=2.99
r85 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.87 $Y=2.905
+ $X2=3.035 $Y2=2.99
r86 16 18 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=2.87 $Y=2.905
+ $X2=2.87 $Y2=2.39
r87 5 50 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.12
r88 5 42 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.91
r89 4 48 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.12
r90 4 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.91
r91 3 46 600 $w=1.7e-07 $l=2.80936e-07 $layer=licon1_PDIFF $count=1 $X=4.45
+ $Y=1.835 $X2=4.63 $Y2=2.04
r92 3 31 300 $w=1.7e-07 $l=7.29469e-07 $layer=licon1_PDIFF $count=2 $X=4.45
+ $Y=1.835 $X2=4.63 $Y2=2.48
r93 2 24 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=3.59
+ $Y=1.835 $X2=3.73 $Y2=2.39
r94 1 18 300 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.835 $X2=2.87 $Y2=2.39
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%VGND 1 2 3 4 5 18 22 24 28 32 34 36 39 40 41
+ 42 43 52 60 69 72 76
r90 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r91 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r92 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r93 67 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r94 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r95 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r96 64 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r97 63 66 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6 $Y2=0
r98 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r99 61 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.775 $Y=0 $X2=4.61
+ $Y2=0
r100 61 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.775 $Y=0
+ $X2=5.04 $Y2=0
r101 60 75 4.40761 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.527 $Y2=0
r102 60 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.335 $Y=0 $X2=6
+ $Y2=0
r103 59 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r104 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r105 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r106 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r107 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r108 53 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=2.795
+ $Y2=0
r109 53 55 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=3.12
+ $Y2=0
r110 52 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.445 $Y=0 $X2=4.61
+ $Y2=0
r111 52 58 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.445 $Y=0
+ $X2=4.08 $Y2=0
r112 51 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r113 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r114 47 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r115 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r116 43 59 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r117 43 56 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r118 41 50 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.77 $Y=0 $X2=1.68
+ $Y2=0
r119 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=1.935
+ $Y2=0
r120 39 46 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.72
+ $Y2=0
r121 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.075
+ $Y2=0
r122 38 50 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.68
+ $Y2=0
r123 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.075
+ $Y2=0
r124 34 75 3.03023 $w=2.9e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.48 $Y=0.085
+ $X2=6.527 $Y2=0
r125 34 36 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=6.48 $Y=0.085
+ $X2=6.48 $Y2=0.38
r126 30 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=0.085
+ $X2=4.61 $Y2=0
r127 30 32 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.61 $Y=0.085 $X2=4.61
+ $Y2=0.485
r128 26 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0
r129 26 28 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0.565
r130 25 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=1.935
+ $Y2=0
r131 24 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.795
+ $Y2=0
r132 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.1
+ $Y2=0
r133 20 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.935 $Y=0.085
+ $X2=1.935 $Y2=0
r134 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.935 $Y=0.085
+ $X2=1.935 $Y2=0.36
r135 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.075 $Y=0.085
+ $X2=1.075 $Y2=0
r136 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.075 $Y=0.085
+ $X2=1.075 $Y2=0.38
r137 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.32
+ $Y=0.235 $X2=6.46 $Y2=0.38
r138 4 32 182 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_NDIFF $count=1 $X=4.45
+ $Y=0.235 $X2=4.61 $Y2=0.485
r139 3 28 182 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_NDIFF $count=1 $X=2.655
+ $Y=0.235 $X2=2.795 $Y2=0.565
r140 2 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.795
+ $Y=0.235 $X2=1.935 $Y2=0.36
r141 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.95
+ $Y=0.235 $X2=1.075 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%A_632_47# 1 2 11
c11 11 0 1.4432e-19 $X=4.16 $Y=0.485
r12 8 11 25.0912 $w=3.93e-07 $l=8.6e-07 $layer=LI1_cond $X=3.3 $Y=0.452 $X2=4.16
+ $Y2=0.452
r13 2 11 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=4.02
+ $Y=0.235 $X2=4.16 $Y2=0.485
r14 1 8 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.16
+ $Y=0.235 $X2=3.3 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_4%A_1006_47# 1 2 7 9 11 16
c19 16 0 1.15476e-19 $X=5.315 $Y=0.452
r20 14 16 5.30602 $w=3.93e-07 $l=1.45e-07 $layer=LI1_cond $X=5.17 $Y=0.452
+ $X2=5.315 $Y2=0.452
r21 9 18 3.75662 $w=2.3e-07 $l=1.38e-07 $layer=LI1_cond $X=6.05 $Y=0.53 $X2=6.05
+ $Y2=0.392
r22 9 11 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.05 $Y=0.53
+ $X2=6.05 $Y2=0.865
r23 7 18 3.13051 $w=2.75e-07 $l=1.15e-07 $layer=LI1_cond $X=5.935 $Y=0.392
+ $X2=6.05 $Y2=0.392
r24 7 16 25.9824 $w=2.73e-07 $l=6.2e-07 $layer=LI1_cond $X=5.935 $Y=0.392
+ $X2=5.315 $Y2=0.392
r25 2 18 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.89
+ $Y=0.235 $X2=6.03 $Y2=0.42
r26 2 11 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=5.89
+ $Y=0.235 $X2=6.03 $Y2=0.865
r27 1 14 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.235 $X2=5.17 $Y2=0.485
.ends

