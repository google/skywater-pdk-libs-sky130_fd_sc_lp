* File: sky130_fd_sc_lp__nand4_0.pex.spice
* Created: Wed Sep  2 10:05:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4_0%D 3 7 12 13 14 15 16 17 23
r33 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.32 $X2=0.63 $Y2=1.32
r34 16 17 7.02459 $w=6.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.4 $Y=1.665 $X2=0.4
+ $Y2=2.035
r35 16 24 6.54995 $w=6.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.4 $Y=1.665
+ $X2=0.4 $Y2=1.32
r36 15 24 0.474634 $w=6.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.4 $Y=1.295
+ $X2=0.4 $Y2=1.32
r37 14 15 7.02459 $w=6.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.4 $Y=0.925 $X2=0.4
+ $Y2=1.295
r38 12 23 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.63 $Y=1.675
+ $X2=0.63 $Y2=1.32
r39 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.7 $Y=1.675 $X2=0.7
+ $Y2=1.825
r40 10 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.155
+ $X2=0.63 $Y2=1.32
r41 7 13 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.86 $Y=2.63
+ $X2=0.86 $Y2=1.825
r42 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.72 $Y=0.445
+ $X2=0.72 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_0%C 3 6 9 10 11 12 13 14 15 21
c47 11 0 3.44906e-20 $X=1.2 $Y=1.435
r48 14 15 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.192 $Y=1.295
+ $X2=1.192 $Y2=1.665
r49 13 14 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.192 $Y=0.925
+ $X2=1.192 $Y2=1.295
r50 13 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2 $Y=0.93
+ $X2=1.2 $Y2=0.93
r51 12 13 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.192 $Y=0.555
+ $X2=1.192 $Y2=0.925
r52 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.2 $Y=1.27 $X2=1.2
+ $Y2=0.93
r53 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.27 $X2=1.2
+ $Y2=1.435
r54 9 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=0.765 $X2=1.2
+ $Y2=0.93
r55 6 11 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=1.29 $Y=2.63
+ $X2=1.29 $Y2=1.435
r56 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.11 $Y=0.445 $X2=1.11
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_0%B 3 6 9 10 11 12 13 14 15 21
c49 11 0 1.77399e-19 $X=1.77 $Y=1.435
r50 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.77
+ $Y=0.93 $X2=1.77 $Y2=0.93
r51 14 15 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.687 $Y=1.295
+ $X2=1.687 $Y2=1.665
r52 14 22 12.5565 $w=3.33e-07 $l=3.65e-07 $layer=LI1_cond $X=1.687 $Y=1.295
+ $X2=1.687 $Y2=0.93
r53 13 22 0.172006 $w=3.33e-07 $l=5e-09 $layer=LI1_cond $X=1.687 $Y=0.925
+ $X2=1.687 $Y2=0.93
r54 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.687 $Y=0.555
+ $X2=1.687 $Y2=0.925
r55 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.77 $Y=1.27
+ $X2=1.77 $Y2=0.93
r56 10 11 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.27
+ $X2=1.77 $Y2=1.435
r57 9 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=0.765
+ $X2=1.77 $Y2=0.93
r58 6 11 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=1.72 $Y=2.63
+ $X2=1.72 $Y2=1.435
r59 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.68 $Y=0.445 $X2=1.68
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_0%A 3 7 10 13 17 18 19 20 21 26
r43 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.34
+ $Y=1.005 $X2=2.34 $Y2=1.005
r44 20 21 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.225 $Y=1.295
+ $X2=2.225 $Y2=1.665
r45 20 27 8.35521 $w=3.98e-07 $l=2.9e-07 $layer=LI1_cond $X=2.225 $Y=1.295
+ $X2=2.225 $Y2=1.005
r46 19 27 2.30489 $w=3.98e-07 $l=8e-08 $layer=LI1_cond $X=2.225 $Y=0.925
+ $X2=2.225 $Y2=1.005
r47 17 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.34 $Y=1.345
+ $X2=2.34 $Y2=1.005
r48 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=1.345
+ $X2=2.34 $Y2=1.51
r49 16 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=0.84
+ $X2=2.34 $Y2=1.005
r50 11 13 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=2.15 $Y=1.75 $X2=2.25
+ $Y2=1.75
r51 10 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.25 $Y=1.675
+ $X2=2.25 $Y2=1.75
r52 10 18 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.675
+ $X2=2.25 $Y2=1.51
r53 7 16 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.84
r54 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.15 $Y=1.825
+ $X2=2.15 $Y2=1.75
r55 1 3 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=2.15 $Y=1.825
+ $X2=2.15 $Y2=2.63
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_0%VPWR 1 2 3 12 16 20 23 24 26 27 29 30 31 44
+ 45
r36 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 42 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 35 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 31 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 31 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 29 41 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 29 30 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.382 $Y2=3.33
r46 28 44 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.53 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 28 30 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.53 $Y=3.33
+ $X2=2.382 $Y2=3.33
r48 26 38 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.375 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 26 27 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.375 $Y=3.33
+ $X2=1.505 $Y2=3.33
r50 25 41 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 25 27 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=1.505 $Y2=3.33
r52 23 34 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 23 24 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.48 $Y=3.33
+ $X2=0.627 $Y2=3.33
r54 22 38 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.775 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 22 24 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.775 $Y=3.33
+ $X2=0.627 $Y2=3.33
r56 18 30 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.382 $Y=3.245
+ $X2=2.382 $Y2=3.33
r57 18 20 30.4714 $w=2.93e-07 $l=7.8e-07 $layer=LI1_cond $X=2.382 $Y=3.245
+ $X2=2.382 $Y2=2.465
r58 14 27 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=3.245
+ $X2=1.505 $Y2=3.33
r59 14 16 34.5733 $w=2.58e-07 $l=7.8e-07 $layer=LI1_cond $X=1.505 $Y=3.245
+ $X2=1.505 $Y2=2.465
r60 10 24 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.627 $Y=3.245
+ $X2=0.627 $Y2=3.33
r61 10 12 30.862 $w=2.93e-07 $l=7.9e-07 $layer=LI1_cond $X=0.627 $Y=3.245
+ $X2=0.627 $Y2=2.455
r62 3 20 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=2.31 $X2=2.365 $Y2=2.465
r63 2 16 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1.365
+ $Y=2.31 $X2=1.505 $Y2=2.465
r64 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.52
+ $Y=2.31 $X2=0.645 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_0%Y 1 2 3 10 12 16 19 21 22 26 28 29 30 31
c52 21 0 2.1189e-19 $X=1.805 $Y=2.025
r53 29 36 3.8266 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=1.075 $Y=2.025
+ $X2=1.205 $Y2=2.025
r54 29 30 22.974 $w=2.08e-07 $l=4.35e-07 $layer=LI1_cond $X=1.245 $Y=2.025
+ $X2=1.68 $Y2=2.025
r55 29 36 2.11255 $w=2.08e-07 $l=4e-08 $layer=LI1_cond $X=1.245 $Y=2.025
+ $X2=1.205 $Y2=2.025
r56 28 31 22.974 $w=2.08e-07 $l=4.35e-07 $layer=LI1_cond $X=2.595 $Y=2.025
+ $X2=2.16 $Y2=2.025
r57 24 26 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.485 $Y=0.445
+ $X2=2.695 $Y2=0.445
r58 21 30 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=2.025
+ $X2=1.68 $Y2=2.025
r59 21 22 6.1471 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=1.805 $Y=2.025
+ $X2=1.935 $Y2=2.025
r60 20 31 5.01732 $w=2.08e-07 $l=9.5e-08 $layer=LI1_cond $X=2.065 $Y=2.025
+ $X2=2.16 $Y2=2.025
r61 20 22 6.1471 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=2.065 $Y=2.025
+ $X2=1.935 $Y2=2.025
r62 19 28 6.82177 $w=2.1e-07 $l=1.46714e-07 $layer=LI1_cond $X=2.695 $Y=1.92
+ $X2=2.595 $Y2=2.025
r63 18 26 3.66692 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0.61
+ $X2=2.695 $Y2=0.445
r64 18 19 72.6455 $w=1.98e-07 $l=1.31e-06 $layer=LI1_cond $X=2.695 $Y=0.61
+ $X2=2.695 $Y2=1.92
r65 14 22 0.586024 $w=2.6e-07 $l=1.05e-07 $layer=LI1_cond $X=1.935 $Y=2.13
+ $X2=1.935 $Y2=2.025
r66 14 16 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=1.935 $Y=2.13
+ $X2=1.935 $Y2=2.455
r67 10 29 3.09071 $w=2.6e-07 $l=1.05e-07 $layer=LI1_cond $X=1.075 $Y=2.13
+ $X2=1.075 $Y2=2.025
r68 10 12 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=1.075 $Y=2.13
+ $X2=1.075 $Y2=2.455
r69 3 16 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.795
+ $Y=2.31 $X2=1.935 $Y2=2.455
r70 2 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.935
+ $Y=2.31 $X2=1.075 $Y2=2.455
r71 1 24 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.485 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_0%VGND 1 6 9 10 11 21 22
r34 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 18 21 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r36 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r37 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r38 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 11 22 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r40 11 19 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r41 9 14 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.24
+ $Y2=0
r42 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.505
+ $Y2=0
r43 8 18 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.72
+ $Y2=0
r44 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.505
+ $Y2=0
r45 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0
r46 4 6 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0.445
r47 1 6 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.38
+ $Y=0.235 $X2=0.505 $Y2=0.445
.ends

