* File: sky130_fd_sc_lp__o21ba_m.spice
* Created: Fri Aug 28 11:06:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ba_m.pex.spice"
.subckt sky130_fd_sc_lp__o21ba_m  VNB VPB B1_N A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_88_41#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0875 AS=0.1113 PD=0.81 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_256_79#_M1008_d N_B1_N_M1008_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.175 PD=2.21 PS=1.62 NRD=0 NRS=10.704 M=1 R=5.6
+ SA=75000.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_500_49#_M1007_d N_A_256_79#_M1007_g N_A_88_41#_M1007_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_500_49#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_500_49#_M1006_d N_A1_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_88_41#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=46.886 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_256_79#_M1005_d N_B1_N_M1005_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.4 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1009 N_A_88_41#_M1009_d N_A_256_79#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_532_535# N_A2_M1003_g N_A_88_41#_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_532_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_42 VNB 0 7.45681e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o21ba_m.pxi.spice"
*
.ends
*
*
