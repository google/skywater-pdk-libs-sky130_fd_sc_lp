* File: sky130_fd_sc_lp__and2_1.pxi.spice
* Created: Wed Sep  2 09:30:14 2020
* 
x_PM_SKY130_FD_SC_LP__AND2_1%A N_A_M1005_g N_A_M1000_g N_A_c_42_n N_A_c_43_n A A
+ PM_SKY130_FD_SC_LP__AND2_1%A
x_PM_SKY130_FD_SC_LP__AND2_1%B N_B_M1003_g N_B_M1002_g B N_B_c_70_n
+ PM_SKY130_FD_SC_LP__AND2_1%B
x_PM_SKY130_FD_SC_LP__AND2_1%A_92_131# N_A_92_131#_M1005_s N_A_92_131#_M1000_d
+ N_A_92_131#_c_102_n N_A_92_131#_M1004_g N_A_92_131#_M1001_g
+ N_A_92_131#_c_104_n N_A_92_131#_c_105_n N_A_92_131#_c_106_n
+ N_A_92_131#_c_124_n N_A_92_131#_c_107_n N_A_92_131#_c_130_n
+ N_A_92_131#_c_108_n PM_SKY130_FD_SC_LP__AND2_1%A_92_131#
x_PM_SKY130_FD_SC_LP__AND2_1%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_c_154_n
+ N_VPWR_c_155_n N_VPWR_c_156_n N_VPWR_c_157_n VPWR N_VPWR_c_158_n
+ N_VPWR_c_159_n N_VPWR_c_153_n N_VPWR_c_161_n PM_SKY130_FD_SC_LP__AND2_1%VPWR
x_PM_SKY130_FD_SC_LP__AND2_1%X N_X_M1004_d N_X_M1001_d X X X X X X X N_X_c_179_n
+ X PM_SKY130_FD_SC_LP__AND2_1%X
x_PM_SKY130_FD_SC_LP__AND2_1%VGND N_VGND_M1003_d N_VGND_c_194_n N_VGND_c_195_n
+ N_VGND_c_196_n VGND N_VGND_c_197_n N_VGND_c_198_n
+ PM_SKY130_FD_SC_LP__AND2_1%VGND
cc_1 VNB N_A_M1005_g 0.0367591f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.865
cc_2 VNB N_A_c_42_n 0.0403612f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.585
cc_3 VNB N_A_c_43_n 0.00772691f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.585
cc_4 VNB A 0.0106608f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_5 VNB N_B_M1003_g 0.0280506f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.865
cc_6 VNB B 0.00278986f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.585
cc_7 VNB N_B_c_70_n 0.0195823f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_A_92_131#_c_102_n 0.0227717f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=2.12
cc_9 VNB N_A_92_131#_M1001_g 0.00774838f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_10 VNB N_A_92_131#_c_104_n 0.0181712f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.585
cc_11 VNB N_A_92_131#_c_105_n 0.0209253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_92_131#_c_106_n 0.00948307f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.62
cc_13 VNB N_A_92_131#_c_107_n 8.92909e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_92_131#_c_108_n 0.0397139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_153_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB X 0.0347025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_X_c_179_n 0.0371756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_194_n 0.0169651f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=2.12
cc_19 VNB N_VGND_c_195_n 0.0393651f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_20 VNB N_VGND_c_196_n 0.00711353f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_21 VNB N_VGND_c_197_n 0.0228166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_198_n 0.180133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VPB N_A_M1000_g 0.0285196f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=2.12
cc_24 VPB N_A_c_42_n 0.0270256f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.585
cc_25 VPB N_A_c_43_n 0.00311897f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.585
cc_26 VPB A 0.00780986f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_27 VPB N_B_M1002_g 0.0245771f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=2.12
cc_28 VPB B 0.00353188f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.585
cc_29 VPB N_B_c_70_n 0.0111564f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_30 VPB N_A_92_131#_M1001_g 0.0251035f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_31 VPB N_A_92_131#_c_107_n 0.00171437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_154_n 0.0790481f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.585
cc_33 VPB N_VPWR_c_155_n 0.0286917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_156_n 0.0155085f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.585
cc_35 VPB N_VPWR_c_157_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.585
cc_36 VPB N_VPWR_c_158_n 0.0252349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_159_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_153_n 0.0839304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_161_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB X 0.0570099f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 N_A_M1005_g N_B_M1003_g 0.0385507f $X=0.8 $Y=0.865 $X2=0 $Y2=0
cc_42 N_A_M1000_g N_B_M1002_g 0.0148899f $X=0.8 $Y=2.12 $X2=0 $Y2=0
cc_43 N_A_c_43_n B 0.00170498f $X=0.8 $Y=1.585 $X2=0 $Y2=0
cc_44 A B 0.021968f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_45 N_A_c_43_n N_B_c_70_n 0.0385507f $X=0.8 $Y=1.585 $X2=0 $Y2=0
cc_46 A N_B_c_70_n 2.84444e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_47 N_A_M1005_g N_A_92_131#_c_104_n 0.00963054f $X=0.8 $Y=0.865 $X2=0 $Y2=0
cc_48 N_A_M1005_g N_A_92_131#_c_105_n 0.0107543f $X=0.8 $Y=0.865 $X2=0 $Y2=0
cc_49 A N_A_92_131#_c_105_n 0.00802377f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_50 N_A_M1005_g N_A_92_131#_c_106_n 0.0041813f $X=0.8 $Y=0.865 $X2=0 $Y2=0
cc_51 N_A_c_42_n N_A_92_131#_c_106_n 0.00767773f $X=0.725 $Y=1.585 $X2=0 $Y2=0
cc_52 A N_A_92_131#_c_106_n 0.0270225f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_53 N_A_M1000_g N_VPWR_c_154_n 0.010786f $X=0.8 $Y=2.12 $X2=0 $Y2=0
cc_54 N_A_c_42_n N_VPWR_c_154_n 0.00674338f $X=0.725 $Y=1.585 $X2=0 $Y2=0
cc_55 A N_VPWR_c_154_n 0.0207706f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_56 N_A_M1000_g N_VPWR_c_153_n 0.00316838f $X=0.8 $Y=2.12 $X2=0 $Y2=0
cc_57 N_A_M1005_g N_VGND_c_194_n 0.00163759f $X=0.8 $Y=0.865 $X2=0 $Y2=0
cc_58 N_A_M1005_g N_VGND_c_195_n 0.00385987f $X=0.8 $Y=0.865 $X2=0 $Y2=0
cc_59 N_A_M1005_g N_VGND_c_198_n 0.0046122f $X=0.8 $Y=0.865 $X2=0 $Y2=0
cc_60 N_B_M1003_g N_A_92_131#_c_102_n 0.0197486f $X=1.16 $Y=0.865 $X2=0 $Y2=0
cc_61 B N_A_92_131#_M1001_g 5.92497e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_62 N_B_c_70_n N_A_92_131#_M1001_g 0.0184849f $X=1.25 $Y=1.585 $X2=0 $Y2=0
cc_63 N_B_M1003_g N_A_92_131#_c_104_n 0.00161163f $X=1.16 $Y=0.865 $X2=0 $Y2=0
cc_64 N_B_M1003_g N_A_92_131#_c_105_n 0.0141493f $X=1.16 $Y=0.865 $X2=0 $Y2=0
cc_65 B N_A_92_131#_c_105_n 0.0292343f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_66 N_B_c_70_n N_A_92_131#_c_105_n 0.005019f $X=1.25 $Y=1.585 $X2=0 $Y2=0
cc_67 N_B_M1002_g N_A_92_131#_c_124_n 0.0131851f $X=1.34 $Y=2.12 $X2=0 $Y2=0
cc_68 B N_A_92_131#_c_124_n 0.0118793f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_69 N_B_M1003_g N_A_92_131#_c_107_n 5.74481e-19 $X=1.16 $Y=0.865 $X2=0 $Y2=0
cc_70 N_B_M1002_g N_A_92_131#_c_107_n 0.00383496f $X=1.34 $Y=2.12 $X2=0 $Y2=0
cc_71 B N_A_92_131#_c_107_n 0.019799f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_72 N_B_c_70_n N_A_92_131#_c_107_n 0.00139158f $X=1.25 $Y=1.585 $X2=0 $Y2=0
cc_73 B N_A_92_131#_c_130_n 0.0150534f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_74 N_B_c_70_n N_A_92_131#_c_130_n 0.00110608f $X=1.25 $Y=1.585 $X2=0 $Y2=0
cc_75 N_B_c_70_n N_A_92_131#_c_108_n 0.00636686f $X=1.25 $Y=1.585 $X2=0 $Y2=0
cc_76 N_B_M1002_g N_VPWR_c_154_n 7.80451e-19 $X=1.34 $Y=2.12 $X2=0 $Y2=0
cc_77 N_B_M1002_g N_VPWR_c_155_n 0.00486239f $X=1.34 $Y=2.12 $X2=0 $Y2=0
cc_78 N_B_M1002_g N_VPWR_c_153_n 0.00377188f $X=1.34 $Y=2.12 $X2=0 $Y2=0
cc_79 N_B_M1003_g N_VGND_c_194_n 0.0107701f $X=1.16 $Y=0.865 $X2=0 $Y2=0
cc_80 N_B_M1003_g N_VGND_c_195_n 0.00332367f $X=1.16 $Y=0.865 $X2=0 $Y2=0
cc_81 N_B_M1003_g N_VGND_c_198_n 0.00387424f $X=1.16 $Y=0.865 $X2=0 $Y2=0
cc_82 N_A_92_131#_c_124_n N_VPWR_M1002_d 0.0090375f $X=1.625 $Y=2.005 $X2=0
+ $Y2=0
cc_83 N_A_92_131#_c_107_n N_VPWR_M1002_d 0.00125488f $X=1.79 $Y=1.35 $X2=0 $Y2=0
cc_84 N_A_92_131#_M1001_g N_VPWR_c_155_n 0.019459f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_92_131#_c_124_n N_VPWR_c_155_n 0.0234822f $X=1.625 $Y=2.005 $X2=0
+ $Y2=0
cc_86 N_A_92_131#_M1001_g N_VPWR_c_159_n 0.00486043f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_87 N_A_92_131#_M1001_g N_VPWR_c_153_n 0.00917987f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_88 N_A_92_131#_c_102_n X 0.0042636f $X=1.7 $Y=1.185 $X2=0 $Y2=0
cc_89 N_A_92_131#_c_105_n X 0.0142103f $X=1.625 $Y=1.235 $X2=0 $Y2=0
cc_90 N_A_92_131#_c_107_n X 0.0422131f $X=1.79 $Y=1.35 $X2=0 $Y2=0
cc_91 N_A_92_131#_c_108_n X 0.019007f $X=1.925 $Y=1.35 $X2=0 $Y2=0
cc_92 N_A_92_131#_c_102_n N_X_c_179_n 0.010948f $X=1.7 $Y=1.185 $X2=0 $Y2=0
cc_93 N_A_92_131#_c_105_n N_X_c_179_n 0.0086126f $X=1.625 $Y=1.235 $X2=0 $Y2=0
cc_94 N_A_92_131#_c_108_n N_X_c_179_n 0.00638032f $X=1.925 $Y=1.35 $X2=0 $Y2=0
cc_95 N_A_92_131#_c_102_n N_VGND_c_194_n 0.00701211f $X=1.7 $Y=1.185 $X2=0 $Y2=0
cc_96 N_A_92_131#_c_104_n N_VGND_c_194_n 0.0094508f $X=0.585 $Y=0.865 $X2=0
+ $Y2=0
cc_97 N_A_92_131#_c_105_n N_VGND_c_194_n 0.0271794f $X=1.625 $Y=1.235 $X2=0
+ $Y2=0
cc_98 N_A_92_131#_c_104_n N_VGND_c_195_n 0.00500197f $X=0.585 $Y=0.865 $X2=0
+ $Y2=0
cc_99 N_A_92_131#_c_102_n N_VGND_c_197_n 0.0054895f $X=1.7 $Y=1.185 $X2=0 $Y2=0
cc_100 N_A_92_131#_c_102_n N_VGND_c_198_n 0.0121525f $X=1.7 $Y=1.185 $X2=0 $Y2=0
cc_101 N_A_92_131#_c_104_n N_VGND_c_198_n 0.0094007f $X=0.585 $Y=0.865 $X2=0
+ $Y2=0
cc_102 N_VPWR_c_153_n N_X_M1001_d 0.00371702f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_103 N_VPWR_c_159_n X 0.018528f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_104 N_VPWR_c_153_n X 0.0104192f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_105 N_X_c_179_n N_VGND_c_197_n 0.0378518f $X=1.915 $Y=0.38 $X2=0 $Y2=0
cc_106 N_X_M1004_d N_VGND_c_198_n 0.00240292f $X=1.775 $Y=0.235 $X2=0 $Y2=0
cc_107 N_X_c_179_n N_VGND_c_198_n 0.0217051f $X=1.915 $Y=0.38 $X2=0 $Y2=0
