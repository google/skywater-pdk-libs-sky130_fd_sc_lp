* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor2_4 A B VGND VNB VPB VPWR Y
X0 Y a_808_39# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR A a_808_39# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR a_808_39# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_808_39# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 Y a_808_39# a_31_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 Y B a_110_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_110_367# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_31_65# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_808_39# B a_1235_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VGND B a_31_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VGND A a_1235_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_110_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_31_65# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_808_39# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VPWR a_808_39# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_808_39# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 Y a_808_39# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VGND A a_31_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_1235_65# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VPWR A a_110_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 Y B a_110_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_31_65# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_110_367# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_1235_65# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VGND A a_1235_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 VPWR B a_808_39# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_808_39# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VGND A a_31_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_31_65# a_808_39# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 a_31_65# a_808_39# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 a_110_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 VPWR A a_808_39# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 VPWR B a_808_39# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 Y a_808_39# a_31_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 a_1235_65# B a_808_39# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 a_31_65# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 a_808_39# B a_1235_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X37 VGND B a_31_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 a_1235_65# B a_808_39# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 VPWR A a_110_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
