* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 a_196_128# SCE a_124_128# VNB nshort w=420000u l=150000u
+  ad=4.311e+11p pd=3.75e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_1912_463# a_871_47# a_1810_463# VPB phighvt w=420000u l=150000u
+  ad=3.969e+11p pd=3.84e+06u as=2.95e+11p ps=3.19e+06u
M1002 a_1912_463# a_871_47# a_1847_125# VNB nshort w=640000u l=150000u
+  ad=4.629e+11p pd=2.95e+06u as=1.344e+11p ps=1.7e+06u
M1003 a_282_128# D a_196_128# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_1263_31# a_1135_57# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.239e+11p pd=1.43e+06u as=2.11845e+12p ps=1.749e+07u
M1005 VGND a_1912_463# a_2598_153# VNB nshort w=420000u l=150000u
+  ad=1.4032e+12p pd=1.305e+07u as=1.113e+11p ps=1.37e+06u
M1006 a_2116_125# a_702_47# a_1912_463# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1007 a_1847_125# a_1135_57# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_1912_463# a_2598_153# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1009 a_27_408# a_324_102# a_196_128# VPB phighvt w=640000u l=150000u
+  ad=3.392e+11p pd=3.62e+06u as=3.609e+11p ps=3.43e+06u
M1010 VPWR a_2158_231# a_1810_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_2158_231# a_1912_463# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1012 VGND SET_B a_2224_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1013 VPWR SCD a_27_408# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_124_128# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_2598_153# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1016 a_871_47# a_702_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1017 a_1703_379# a_702_47# a_1912_463# VPB phighvt w=840000u l=150000u
+  ad=4.44375e+11p pd=4.42e+06u as=0p ps=0u
M1018 a_1135_57# a_702_47# a_196_128# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1019 a_1221_57# a_871_47# a_1135_57# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1020 VPWR SET_B a_1263_31# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND SET_B a_1502_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.512e+11p ps=1.56e+06u
M1022 VGND a_1263_31# a_1221_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1135_57# a_871_47# a_196_128# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1024 a_2224_125# a_2158_231# a_2116_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND CLK a_702_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1026 a_324_102# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1027 VPWR CLK a_702_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.459e+11p ps=2.7e+06u
M1028 a_1221_463# a_702_47# a_1135_57# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1029 a_1703_379# a_1135_57# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Q a_2598_153# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1031 a_2158_231# a_1912_463# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1032 VPWR a_1263_31# a_1221_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_196_408# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1034 VGND a_324_102# a_282_128# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1912_463# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_196_128# D a_196_408# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_871_47# a_702_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1038 a_324_102# SCE VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1039 a_1502_125# a_1135_57# a_1263_31# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends
