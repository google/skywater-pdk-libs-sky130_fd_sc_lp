* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor2_0 A B VGND VNB VPB VPWR Y
X0 a_143_487# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VPWR A a_383_487# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_383_487# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_300_60# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_110_177# B a_143_487# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND A a_110_177# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND B a_300_60# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_300_60# a_143_487# Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR A a_143_487# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 Y a_143_487# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
