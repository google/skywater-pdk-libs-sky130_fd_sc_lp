* File: sky130_fd_sc_lp__and4b_lp.spice
* Created: Wed Sep  2 09:33:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4b_lp.pex.spice"
.subckt sky130_fd_sc_lp__and4b_lp  VNB VPB D C B A_N X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A_N	A_N
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1006 A_114_47# N_A_84_21#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_84_21#_M1012_g A_114_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.0441 PD=0.72 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 A_276_47# N_D_M1000_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.063 PD=0.66 PS=0.72 NRD=18.564 NRS=5.712 M=1 R=2.8 SA=75001 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1001 A_354_47# N_C_M1001_g A_276_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.4 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1002 A_432_47# N_B_M1002_g A_354_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_84_21#_M1010_d N_A_480_21#_M1010_g A_432_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 A_708_47# N_A_N_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_480_21#_M1003_d N_A_N_M1003_g A_708_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_84_21#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1013 N_A_84_21#_M1013_d N_D_M1013_g N_VPWR_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_C_M1009_g N_A_84_21#_M1013_d VPB PHIGHVT L=0.25 W=1
+ AD=0.15 AS=0.14 PD=1.3 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1011 N_A_84_21#_M1011_d N_B_M1011_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.15 PD=1.28 PS=1.3 NRD=0 NRS=3.9203 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A_480_21#_M1007_g N_A_84_21#_M1011_d VPB PHIGHVT L=0.25
+ W=1 AD=0.28 AS=0.14 PD=1.56 PS=1.28 NRD=7.8603 NRS=0 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1005 N_A_480_21#_M1005_d N_A_N_M1005_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.28 PD=2.57 PS=1.56 NRD=0 NRS=47.28 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__and4b_lp.pxi.spice"
*
.ends
*
*
