* File: sky130_fd_sc_lp__isolatch_lp.pex.spice
* Created: Fri Aug 28 10:42:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%D 3 7 9 10 14 15 17 18 26
c54 26 0 1.57135e-19 $X=0.66 $Y=1.42
c55 14 0 1.83485e-19 $X=0.42 $Y=2.35
c56 7 0 7.93832e-20 $X=1.085 $Y=0.835
r57 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.66
+ $Y=1.42 $X2=0.66 $Y2=1.42
r58 18 27 1.36695 $w=5.23e-07 $l=6e-08 $layer=LI1_cond $X=0.72 $Y=1.517 $X2=0.66
+ $Y2=1.517
r59 17 29 2.30558 $w=5.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.21 $Y=1.517
+ $X2=0.295 $Y2=1.517
r60 17 27 7.97386 $w=5.23e-07 $l=3.5e-07 $layer=LI1_cond $X=0.31 $Y=1.517
+ $X2=0.66 $Y2=1.517
r61 17 29 0.341737 $w=5.23e-07 $l=1.5e-08 $layer=LI1_cond $X=0.31 $Y=1.517
+ $X2=0.295 $Y2=1.517
r62 15 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=2.35
+ $X2=0.42 $Y2=2.515
r63 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.42
+ $Y=2.35 $X2=0.42 $Y2=2.35
r64 11 14 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.21 $Y=2.35
+ $X2=0.42 $Y2=2.35
r65 10 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.21 $Y=2.185
+ $X2=0.21 $Y2=2.35
r66 9 17 7.13375 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.21 $Y=1.78 $X2=0.21
+ $Y2=1.517
r67 9 10 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.21 $Y=1.78
+ $X2=0.21 $Y2=2.185
r68 5 26 71.1285 $w=2.88e-07 $l=5.09166e-07 $layer=POLY_cond $X=1.085 $Y=1.215
+ $X2=0.66 $Y2=1.4
r69 5 7 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.085 $Y=1.215
+ $X2=1.085 $Y2=0.835
r70 3 24 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.51 $Y=2.885
+ $X2=0.51 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_36_73# 1 2 9 13 17 19 20 21 22 24 25
+ 26 28 29 30 33 43
c129 21 0 1.57135e-19 $X=1.24 $Y=2.12
c130 17 0 7.93832e-20 $X=0.325 $Y=0.575
r131 42 43 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=1.475 $Y=1.77
+ $X2=1.925 $Y2=1.77
r132 39 42 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.35 $Y=1.77
+ $X2=1.475 $Y2=1.77
r133 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.35
+ $Y=1.77 $X2=1.35 $Y2=1.77
r134 33 35 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=3.17 $Y=2.22
+ $X2=3.17 $Y2=2.9
r135 31 33 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=3.17 $Y=1.955
+ $X2=3.17 $Y2=2.22
r136 29 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.045 $Y=1.87
+ $X2=3.17 $Y2=1.955
r137 29 30 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.045 $Y=1.87
+ $X2=2.345 $Y2=1.87
r138 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.26 $Y=1.955
+ $X2=2.345 $Y2=1.87
r139 27 28 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.26 $Y=1.955
+ $X2=2.26 $Y2=2.905
r140 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.175 $Y=2.99
+ $X2=2.26 $Y2=2.905
r141 25 26 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.175 $Y=2.99
+ $X2=1.325 $Y2=2.99
r142 24 38 6.64448 $w=3.41e-07 $l=1.28452e-07 $layer=LI1_cond $X=1.27 $Y=1.67
+ $X2=1.335 $Y2=1.77
r143 23 24 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.27 $Y=1.085
+ $X2=1.27 $Y2=1.67
r144 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.24 $Y=2.905
+ $X2=1.325 $Y2=2.99
r145 21 38 15.5888 $w=3.41e-07 $l=3.94652e-07 $layer=LI1_cond $X=1.24 $Y=2.12
+ $X2=1.335 $Y2=1.77
r146 21 22 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.24 $Y=2.12
+ $X2=1.24 $Y2=2.905
r147 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.185 $Y=1
+ $X2=1.27 $Y2=1.085
r148 19 20 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.185 $Y=1
+ $X2=0.41 $Y2=1
r149 15 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.285 $Y=0.915
+ $X2=0.41 $Y2=1
r150 15 17 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.285 $Y=0.915
+ $X2=0.285 $Y2=0.575
r151 11 43 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.935
+ $X2=1.925 $Y2=1.77
r152 11 13 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.925 $Y=1.935
+ $X2=1.925 $Y2=2.595
r153 7 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.605
+ $X2=1.475 $Y2=1.77
r154 7 9 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.475 $Y=1.605
+ $X2=1.475 $Y2=0.835
r155 2 35 400 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=3.07
+ $Y=2.095 $X2=3.21 $Y2=2.9
r156 2 33 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.07
+ $Y=2.095 $X2=3.21 $Y2=2.22
r157 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.365 $X2=0.325 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_21_179# 1 2 8 9 10 11 12 16 17 18 20
+ 21 22 25 30 33 35 39 42 46 48 51 52 54 56
c159 52 0 1.43968e-19 $X=2.08 $Y=1.06
c160 25 0 1.83485e-19 $X=1.33 $Y=2.885
r161 54 55 11.6304 $w=2.57e-07 $l=2.45e-07 $layer=LI1_cond $X=3.855 $Y=1.45
+ $X2=4.1 $Y2=1.45
r162 52 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.08 $Y=1.06
+ $X2=2.08 $Y2=0.895
r163 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.06 $X2=2.08 $Y2=1.06
r164 46 56 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4.14 $Y=2.18
+ $X2=4.14 $Y2=2.055
r165 46 48 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=4.14 $Y=2.18 $X2=4.14
+ $Y2=2.22
r166 44 55 3.1561 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=1.615 $X2=4.1
+ $Y2=1.45
r167 44 56 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.1 $Y=1.615
+ $X2=4.1 $Y2=2.055
r168 40 54 0.884329 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=1.285
+ $X2=3.855 $Y2=1.45
r169 40 42 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=3.855 $Y=1.285
+ $X2=3.855 $Y2=0.76
r170 39 62 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.985 $Y=1.45
+ $X2=2.985 $Y2=1.615
r171 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.985
+ $Y=1.45 $X2=2.985 $Y2=1.45
r172 36 51 20.8684 $w=2.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.08 $Y=1.45
+ $X2=2.08 $Y2=1.06
r173 36 38 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=2.245 $Y=1.45
+ $X2=2.985 $Y2=1.45
r174 35 54 5.25093 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=3.73 $Y=1.45
+ $X2=3.855 $Y2=1.45
r175 35 38 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=3.73 $Y=1.45
+ $X2=2.985 $Y2=1.45
r176 33 62 243.485 $w=2.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.945 $Y=2.595
+ $X2=2.945 $Y2=1.615
r177 30 58 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.02 $Y=0.575
+ $X2=2.02 $Y2=0.895
r178 27 30 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.02 $Y=0.255
+ $X2=2.02 $Y2=0.575
r179 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.33 $Y=2.325
+ $X2=1.33 $Y2=2.885
r180 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.255 $Y=2.25
+ $X2=1.33 $Y2=2.325
r181 21 22 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.255 $Y=2.25
+ $X2=0.945 $Y2=2.25
r182 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.87 $Y=2.175
+ $X2=0.945 $Y2=2.25
r183 19 20 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=0.87 $Y=1.975
+ $X2=0.87 $Y2=2.175
r184 17 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.945 $Y=0.18
+ $X2=2.02 $Y2=0.255
r185 17 18 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=1.945 $Y=0.18
+ $X2=0.615 $Y2=0.18
r186 14 16 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=0.895
+ $X2=0.54 $Y2=0.575
r187 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.54 $Y=0.255
+ $X2=0.615 $Y2=0.18
r188 13 16 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=0.255
+ $X2=0.54 $Y2=0.575
r189 11 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.795 $Y=1.9
+ $X2=0.87 $Y2=1.975
r190 11 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.795 $Y=1.9
+ $X2=0.255 $Y2=1.9
r191 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.465 $Y=0.97
+ $X2=0.54 $Y2=0.895
r192 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.465 $Y=0.97
+ $X2=0.255 $Y2=0.97
r193 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.18 $Y=1.825
+ $X2=0.255 $Y2=1.9
r194 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.18 $Y=1.045
+ $X2=0.255 $Y2=0.97
r195 7 8 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.18 $Y=1.045
+ $X2=0.18 $Y2=1.825
r196 2 48 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=2.075 $X2=4.18 $Y2=2.22
r197 1 42 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=3.75
+ $Y=0.465 $X2=3.895 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_458_293# 1 2 9 11 13 16 18 20 21 25 26
+ 27 28 30 33 34 36 37 39 40 41 44 47 49 51
c149 49 0 5.82594e-20 $X=5.5 $Y=2.08
c150 41 0 1.57765e-19 $X=4.605 $Y=2.035
c151 34 0 5.8299e-20 $X=3.68 $Y=1.95
c152 30 0 1.35042e-19 $X=3.68 $Y=1.785
c153 26 0 1.51853e-19 $X=2.447 $Y=1.615
r154 51 53 9.2829 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=5.562 $Y=0.61
+ $X2=5.562 $Y2=0.775
r155 47 49 3.70735 $w=2.5e-07 $l=1.3625e-07 $layer=LI1_cond $X=5.58 $Y=1.915
+ $X2=5.5 $Y2=2.017
r156 47 53 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=5.58 $Y=1.915
+ $X2=5.58 $Y2=0.775
r157 42 49 3.70735 $w=2.5e-07 $l=1.03e-07 $layer=LI1_cond $X=5.5 $Y=2.12 $X2=5.5
+ $Y2=2.017
r158 42 44 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=5.5 $Y=2.12 $X2=5.5
+ $Y2=2.79
r159 40 49 2.76166 $w=1.7e-07 $l=1.73767e-07 $layer=LI1_cond $X=5.335 $Y=2.035
+ $X2=5.5 $Y2=2.017
r160 40 41 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.335 $Y=2.035
+ $X2=4.605 $Y2=2.035
r161 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.52 $Y=2.12
+ $X2=4.605 $Y2=2.035
r162 38 39 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=4.52 $Y=2.12
+ $X2=4.52 $Y2=2.905
r163 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=2.99
+ $X2=4.52 $Y2=2.905
r164 36 37 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.435 $Y=2.99
+ $X2=3.845 $Y2=2.99
r165 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.68
+ $Y=1.95 $X2=3.68 $Y2=1.95
r166 31 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.68 $Y=2.905
+ $X2=3.845 $Y2=2.99
r167 31 33 33.351 $w=3.28e-07 $l=9.55e-07 $layer=LI1_cond $X=3.68 $Y=2.905
+ $X2=3.68 $Y2=1.95
r168 30 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.785
+ $X2=3.68 $Y2=1.95
r169 25 26 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.447 $Y=1.465
+ $X2=2.447 $Y2=1.615
r170 23 30 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.59 $Y=1.045
+ $X2=3.59 $Y2=1.785
r171 22 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.995 $Y=0.97
+ $X2=2.92 $Y2=0.97
r172 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.515 $Y=0.97
+ $X2=3.59 $Y2=1.045
r173 21 22 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.515 $Y=0.97
+ $X2=2.995 $Y2=0.97
r174 18 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.92 $Y=0.895
+ $X2=2.92 $Y2=0.97
r175 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.92 $Y=0.895
+ $X2=2.92 $Y2=0.575
r176 17 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.605 $Y=0.97
+ $X2=2.53 $Y2=0.97
r177 16 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.845 $Y=0.97
+ $X2=2.92 $Y2=0.97
r178 16 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.845 $Y=0.97
+ $X2=2.605 $Y2=0.97
r179 14 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.53 $Y=1.045
+ $X2=2.53 $Y2=0.97
r180 14 25 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.53 $Y=1.045
+ $X2=2.53 $Y2=1.465
r181 11 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.53 $Y=0.895
+ $X2=2.53 $Y2=0.97
r182 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.53 $Y=0.895
+ $X2=2.53 $Y2=0.575
r183 9 26 243.485 $w=2.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.415 $Y=2.595
+ $X2=2.415 $Y2=1.615
r184 2 49 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.935 $X2=5.5 $Y2=2.08
r185 2 44 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.935 $X2=5.5 $Y2=2.79
r186 1 51 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.465 $X2=5.545 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%SLEEP_B 3 5 6 9 11 13 15
c52 15 0 1.35042e-19 $X=4.56 $Y=1.665
c53 11 0 1.57765e-19 $X=4.51 $Y=1.78
r54 17 19 37.4369 $w=3.09e-07 $l=2.4e-07 $layer=POLY_cond $X=4.52 $Y=1.375
+ $X2=4.52 $Y2=1.615
r55 15 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.52
+ $Y=1.615 $X2=4.52 $Y2=1.615
r56 11 19 38.532 $w=3.09e-07 $l=1.69926e-07 $layer=POLY_cond $X=4.51 $Y=1.78
+ $X2=4.52 $Y2=1.615
r57 11 13 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.51 $Y=1.78
+ $X2=4.51 $Y2=2.395
r58 7 17 24.4932 $w=3.09e-07 $l=9.68246e-08 $layer=POLY_cond $X=4.47 $Y=1.3
+ $X2=4.52 $Y2=1.375
r59 7 9 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=4.47 $Y=1.3 $X2=4.47
+ $Y2=0.675
r60 5 17 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.375
+ $X2=4.52 $Y2=1.375
r61 5 6 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.355 $Y=1.375
+ $X2=4.185 $Y2=1.375
r62 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.11 $Y=1.3
+ $X2=4.185 $Y2=1.375
r63 1 3 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=4.11 $Y=1.3 $X2=4.11
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_281_535# 1 2 9 13 15 16 18 21 23 27 29
+ 31 32 34 36 42 43 45 48 51 52 53 55 56 57 59 60 61 65 66 72 75 78 79
c187 75 0 1.51853e-19 $X=1.77 $Y=1.415
c188 51 0 1.43968e-19 $X=2.5 $Y=0.945
c189 27 0 5.82594e-20 $X=6.295 $Y=2.435
r190 78 79 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.06
+ $Y=1.24 $X2=5.06 $Y2=1.24
r191 73 75 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.66 $Y=1.415
+ $X2=1.77 $Y2=1.415
r192 71 72 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0.535
+ $X2=1.97 $Y2=0.535
r193 68 71 4.39748 $w=3.78e-07 $l=1.45e-07 $layer=LI1_cond $X=1.66 $Y=0.535
+ $X2=1.805 $Y2=0.535
r194 65 66 10.2717 $w=3.58e-07 $l=2.2e-07 $layer=LI1_cond $X=1.675 $Y=2.51
+ $X2=1.675 $Y2=2.29
r195 60 78 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=1.16
+ $X2=5.06 $Y2=1.16
r196 60 61 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.895 $Y=1.16
+ $X2=4.32 $Y2=1.16
r197 59 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.235 $Y=1.075
+ $X2=4.32 $Y2=1.16
r198 58 59 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.235 $Y=0.425
+ $X2=4.235 $Y2=1.075
r199 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.15 $Y=0.34
+ $X2=4.235 $Y2=0.425
r200 56 57 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.15 $Y=0.34
+ $X2=3.56 $Y2=0.34
r201 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.475 $Y=0.425
+ $X2=3.56 $Y2=0.34
r202 54 55 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.475 $Y=0.425
+ $X2=3.475 $Y2=0.945
r203 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.39 $Y=1.03
+ $X2=3.475 $Y2=0.945
r204 52 53 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=3.39 $Y=1.03
+ $X2=2.585 $Y2=1.03
r205 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.5 $Y=0.945
+ $X2=2.585 $Y2=1.03
r206 50 51 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.5 $Y=0.725
+ $X2=2.5 $Y2=0.945
r207 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.415 $Y=0.64
+ $X2=2.5 $Y2=0.725
r208 48 72 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.415 $Y=0.64
+ $X2=1.97 $Y2=0.64
r209 46 75 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=1.5
+ $X2=1.77 $Y2=1.415
r210 46 66 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.77 $Y=1.5
+ $X2=1.77 $Y2=2.29
r211 45 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=1.33
+ $X2=1.66 $Y2=1.415
r212 44 68 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.66 $Y=0.725
+ $X2=1.66 $Y2=0.535
r213 44 45 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.66 $Y=0.725
+ $X2=1.66 $Y2=1.33
r214 40 79 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.06 $Y=1.225
+ $X2=5.06 $Y2=1.24
r215 40 41 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.06 $Y=1.15
+ $X2=5.33 $Y2=1.15
r216 37 40 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.97 $Y=1.15 $X2=5.06
+ $Y2=1.15
r217 34 36 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.705 $Y=1.425
+ $X2=6.705 $Y2=1.095
r218 33 43 15.684 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=6.42 $Y=1.5
+ $X2=6.295 $Y2=1.5
r219 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.63 $Y=1.5
+ $X2=6.705 $Y2=1.425
r220 32 33 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.63 $Y=1.5
+ $X2=6.42 $Y2=1.5
r221 29 43 8.77658 $w=1.5e-07 $l=9.68246e-08 $layer=POLY_cond $X=6.345 $Y=1.425
+ $X2=6.295 $Y2=1.5
r222 29 31 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.345 $Y=1.425
+ $X2=6.345 $Y2=1.095
r223 25 43 8.77658 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.295 $Y=1.575
+ $X2=6.295 $Y2=1.5
r224 25 27 213.67 $w=2.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.295 $Y=1.575
+ $X2=6.295 $Y2=2.435
r225 24 42 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=5.89 $Y=1.5
+ $X2=5.765 $Y2=1.5
r226 23 43 15.684 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=6.17 $Y=1.5
+ $X2=6.295 $Y2=1.5
r227 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.17 $Y=1.5
+ $X2=5.89 $Y2=1.5
r228 19 42 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=5.765 $Y=1.575
+ $X2=5.765 $Y2=1.5
r229 19 21 213.67 $w=2.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.765 $Y=1.575
+ $X2=5.765 $Y2=2.435
r230 18 42 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=5.715 $Y=1.425
+ $X2=5.765 $Y2=1.5
r231 17 18 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.715 $Y=1.225
+ $X2=5.715 $Y2=1.425
r232 16 41 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.405 $Y=1.15
+ $X2=5.33 $Y2=1.15
r233 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.64 $Y=1.15
+ $X2=5.715 $Y2=1.225
r234 15 16 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.64 $Y=1.15
+ $X2=5.405 $Y2=1.15
r235 11 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.33 $Y=1.075
+ $X2=5.33 $Y2=1.15
r236 11 13 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.33 $Y=1.075
+ $X2=5.33 $Y2=0.675
r237 7 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.97 $Y=1.075
+ $X2=4.97 $Y2=1.15
r238 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.97 $Y=1.075 $X2=4.97
+ $Y2=0.675
r239 2 65 600 $w=1.7e-07 $l=3.27261e-07 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=2.675 $X2=1.66 $Y2=2.51
r240 1 71 182 $w=1.7e-07 $l=2.96606e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.625 $X2=1.805 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%VPWR 1 4 6 8 15 16
r53 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 15 16 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r55 13 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 12 15 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r57 12 13 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 10 19 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=3.33 $X2=0.23
+ $Y2=3.33
r59 10 12 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 8 16 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r61 8 13 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 4 19 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.23 $Y2=3.33
r63 4 6 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.9
r64 1 6 600 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.675 $X2=0.295 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%KAPWR 1 2 3 10 13 21 28 33
c66 33 0 5.8299e-20 $X=6 $Y=2.82
r67 31 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=2.82 $X2=6
+ $Y2=2.82
r68 28 31 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.03 $Y=2.08 $X2=6.03
+ $Y2=2.79
r69 25 33 0.52469 $w=2.7e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=2.81 $X2=6
+ $Y2=2.81
r70 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.82
+ $X2=5.04 $Y2=2.82
r71 21 24 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=4.965 $Y=2.51
+ $X2=4.965 $Y2=2.82
r72 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=2.82
+ $X2=2.64 $Y2=2.82
r73 13 16 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=2.68 $Y=2.22 $X2=2.68
+ $Y2=2.82
r74 10 25 0.787035 $w=2.7e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=2.81
+ $X2=5.04 $Y2=2.81
r75 10 17 0.52469 $w=2.7e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=2.81 $X2=2.64
+ $Y2=2.81
r76 3 31 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=1.935 $X2=6.03 $Y2=2.79
r77 3 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=1.935 $X2=6.03 $Y2=2.08
r78 2 21 600 $w=1.7e-07 $l=5.86217e-07 $layer=licon1_PDIFF $count=1 $X=4.585
+ $Y=2.075 $X2=4.94 $Y2=2.51
r79 1 16 400 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=2.095 $X2=2.68 $Y2=2.9
r80 1 13 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=2.095 $X2=2.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%Q 1 2 7 8 9 10 11
r14 31 33 13.3735 $w=6.33e-07 $l=7.1e-07 $layer=LI1_cond $X=6.767 $Y=2.08
+ $X2=6.767 $Y2=2.79
r15 11 31 0.847615 $w=6.33e-07 $l=4.5e-08 $layer=LI1_cond $X=6.767 $Y=2.035
+ $X2=6.767 $Y2=2.08
r16 10 11 6.96928 $w=6.33e-07 $l=3.7e-07 $layer=LI1_cond $X=6.767 $Y=1.665
+ $X2=6.767 $Y2=2.035
r17 9 10 6.96928 $w=6.33e-07 $l=3.7e-07 $layer=LI1_cond $X=6.767 $Y=1.295
+ $X2=6.767 $Y2=1.665
r18 9 23 3.76718 $w=6.33e-07 $l=2e-07 $layer=LI1_cond $X=6.767 $Y=1.295
+ $X2=6.767 $Y2=1.095
r19 8 23 3.2021 $w=6.33e-07 $l=1.7e-07 $layer=LI1_cond $X=6.767 $Y=0.925
+ $X2=6.767 $Y2=1.095
r20 7 8 6.96928 $w=6.33e-07 $l=3.7e-07 $layer=LI1_cond $X=6.767 $Y=0.555
+ $X2=6.767 $Y2=0.925
r21 2 33 400 $w=1.7e-07 $l=9.47497e-07 $layer=licon1_PDIFF $count=1 $X=6.42
+ $Y=1.935 $X2=6.615 $Y2=2.79
r22 2 31 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=6.42
+ $Y=1.935 $X2=6.615 $Y2=2.08
r23 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.78
+ $Y=0.885 $X2=6.92 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_LP__ISOLATCH_LP%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39
+ 54 60 61 64 67 70
r79 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r80 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r81 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r82 61 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6
+ $Y2=0
r83 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r84 58 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.28 $Y=0 $X2=6.115
+ $Y2=0
r85 58 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.28 $Y=0 $X2=6.96
+ $Y2=0
r86 57 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r87 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r88 54 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.95 $Y=0 $X2=6.115
+ $Y2=0
r89 54 56 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=5.95 $Y=0 $X2=5.04
+ $Y2=0
r90 53 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r91 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r92 49 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r93 47 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.095
+ $Y2=0
r94 47 49 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.6
+ $Y2=0
r95 46 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r96 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r97 43 46 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r98 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r99 42 45 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r100 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r101 40 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=0.755
+ $Y2=0
r102 40 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=1.2
+ $Y2=0
r103 39 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=3.095
+ $Y2=0
r104 39 45 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=2.64
+ $Y2=0
r105 37 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r106 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r107 34 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.59 $Y=0 $X2=0.755
+ $Y2=0
r108 34 36 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.59 $Y=0 $X2=0.24
+ $Y2=0
r109 32 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r110 32 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r111 32 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r112 30 52 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.56
+ $Y2=0
r113 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.725
+ $Y2=0
r114 29 56 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.85 $Y=0 $X2=5.04
+ $Y2=0
r115 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.85 $Y=0 $X2=4.725
+ $Y2=0
r116 25 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.115 $Y=0.085
+ $X2=6.115 $Y2=0
r117 25 27 37.5417 $w=3.28e-07 $l=1.075e-06 $layer=LI1_cond $X=6.115 $Y=0.085
+ $X2=6.115 $Y2=1.16
r118 21 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.725 $Y=0.085
+ $X2=4.725 $Y2=0
r119 21 23 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=4.725 $Y=0.085
+ $X2=4.725 $Y2=0.675
r120 17 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0
r121 17 19 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0.56
r122 13 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r123 13 15 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.545
r124 4 27 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=5.97
+ $Y=0.885 $X2=6.115 $Y2=1.16
r125 3 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.545
+ $Y=0.465 $X2=4.685 $Y2=0.675
r126 2 19 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.365 $X2=3.135 $Y2=0.56
r127 1 15 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.365 $X2=0.755 $Y2=0.545
.ends

