* File: sky130_fd_sc_lp__bufkapwr_1.spice
* Created: Wed Sep  2 09:35:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__bufkapwr_1.pex.spice"
.subckt sky130_fd_sc_lp__bufkapwr_1  VNB VPB A X KAPWR VGND VPWR
* 
* VGND	VGND
* KAPWR	KAPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_69_161#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.1113 PD=0.75 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_69_161#_M1002_d N_A_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0693 PD=1.37 PS=0.75 NRD=0 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_KAPWR_M1003_d N_A_69_161#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_A_69_161#_M1000_d N_A_M1000_g N_KAPWR_M1003_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__bufkapwr_1.pxi.spice"
*
.ends
*
*
