* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_103_263# B1 a_549_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR A2 a_549_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 X a_103_263# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND A2 a_1006_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND a_103_263# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 X a_103_263# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_632_47# B1 a_103_263# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_549_367# B1 a_103_263# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_103_263# B1 a_632_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 X a_103_263# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR a_103_263# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_632_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VGND B2 a_632_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VPWR a_103_263# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_549_367# B2 a_103_263# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_103_263# B2 a_549_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_1006_47# A1 a_103_263# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_549_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_549_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VGND a_103_263# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VPWR A1 a_549_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 X a_103_263# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_103_263# A1 a_1006_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_1006_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
