* File: sky130_fd_sc_lp__a211o_0.pex.spice
* Created: Wed Sep  2 09:17:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211O_0%A_80_172# 1 2 3 11 14 18 20 23 27 29 35 39
+ 42 43 44 45 47 48
c93 43 0 1.26458e-19 $X=0.59 $Y=1.025
r94 47 48 9.92865 $w=5.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.817 $Y=2.555
+ $X2=2.817 $Y2=2.39
r95 43 51 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.025
+ $X2=0.577 $Y2=0.86
r96 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.025 $X2=0.59 $Y2=1.025
r97 37 39 13.4452 $w=2.98e-07 $l=3.5e-07 $layer=LI1_cond $X=3.04 $Y=0.86
+ $X2=3.04 $Y2=0.51
r98 36 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=0.945
+ $X2=2.62 $Y2=0.945
r99 35 37 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.89 $Y=0.945
+ $X2=3.04 $Y2=0.86
r100 35 36 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.89 $Y=0.945
+ $X2=2.705 $Y2=0.945
r101 31 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.03
+ $X2=2.62 $Y2=0.945
r102 31 48 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.62 $Y=1.03
+ $X2=2.62 $Y2=2.39
r103 30 44 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.96 $Y=0.945
+ $X2=1.81 $Y2=0.945
r104 29 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=0.945
+ $X2=2.62 $Y2=0.945
r105 29 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.535 $Y=0.945
+ $X2=1.96 $Y2=0.945
r106 25 44 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0.86 $X2=1.81
+ $Y2=0.945
r107 25 27 13.4452 $w=2.98e-07 $l=3.5e-07 $layer=LI1_cond $X=1.81 $Y=0.86
+ $X2=1.81 $Y2=0.51
r108 24 42 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.755 $Y=0.945
+ $X2=0.63 $Y2=0.945
r109 23 44 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.66 $Y=0.945
+ $X2=1.81 $Y2=0.945
r110 23 24 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.66 $Y=0.945
+ $X2=0.755 $Y2=0.945
r111 18 51 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.48 $Y=0.51
+ $X2=0.48 $Y2=0.86
r112 14 20 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=0.475 $Y=2.52
+ $X2=0.475 $Y2=1.53
r113 11 20 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.577 $Y=1.353
+ $X2=0.577 $Y2=1.53
r114 10 43 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.577 $Y=1.037
+ $X2=0.577 $Y2=1.025
r115 10 11 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.577 $Y=1.037
+ $X2=0.577 $Y2=1.353
r116 3 47 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.795
+ $Y=2.41 $X2=2.935 $Y2=2.555
r117 2 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.885
+ $Y=0.3 $X2=3.025 $Y2=0.51
r118 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.3 $X2=1.825 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_0%A2 3 6 9 13 14 17 19 20 24
r52 19 20 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=1.295
+ $X2=1.17 $Y2=1.665
r53 19 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=1.375 $X2=1.16 $Y2=1.375
r54 15 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.25 $Y=2.205
+ $X2=1.46 $Y2=2.205
r55 13 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.16 $Y=1.715
+ $X2=1.16 $Y2=1.375
r56 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.715
+ $X2=1.16 $Y2=1.88
r57 12 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.21
+ $X2=1.16 $Y2=1.375
r58 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.46 $Y=2.28 $X2=1.46
+ $Y2=2.205
r59 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.46 $Y=2.28 $X2=1.46
+ $Y2=2.73
r60 6 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.25 $Y=2.13 $X2=1.25
+ $Y2=2.205
r61 6 14 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.25 $Y=2.13 $X2=1.25
+ $Y2=1.88
r62 3 12 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=1.25 $Y=0.51 $X2=1.25
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_0%A1 3 6 8 11 13 16 18 19 23
c49 18 0 1.08716e-19 $X=1.68 $Y=1.295
c50 16 0 1.19954e-19 $X=1.93 $Y=2.195
c51 11 0 2.70489e-20 $X=1.93 $Y=2.73
c52 3 0 5.48067e-20 $X=1.61 $Y=0.51
r53 23 25 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.385
+ $X2=1.715 $Y2=1.22
r54 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=1.385 $X2=1.73 $Y2=1.385
r55 19 24 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=1.682 $Y=1.665
+ $X2=1.682 $Y2=1.385
r56 18 24 3.40065 $w=3.03e-07 $l=9e-08 $layer=LI1_cond $X=1.682 $Y=1.295
+ $X2=1.682 $Y2=1.385
r57 14 16 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.82 $Y=2.195
+ $X2=1.93 $Y2=2.195
r58 9 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.93 $Y=2.27 $X2=1.93
+ $Y2=2.195
r59 9 11 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.93 $Y=2.27 $X2=1.93
+ $Y2=2.73
r60 8 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.82 $Y=2.12 $X2=1.82
+ $Y2=2.195
r61 8 13 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.82 $Y=2.12 $X2=1.82
+ $Y2=1.89
r62 6 13 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.715 $Y=1.71
+ $X2=1.715 $Y2=1.89
r63 5 23 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.715 $Y=1.4
+ $X2=1.715 $Y2=1.385
r64 5 6 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.715 $Y=1.4 $X2=1.715
+ $Y2=1.71
r65 3 25 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.61 $Y=0.51 $X2=1.61
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_0%B1 1 3 8 12 15 16 17 18 19 23
c46 18 0 5.48067e-20 $X=2.16 $Y=1.295
c47 15 0 5.95004e-20 $X=2.27 $Y=1.21
c48 8 0 4.92156e-20 $X=2.36 $Y=2.73
r49 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.27
+ $Y=1.375 $X2=2.27 $Y2=1.375
r50 19 24 9.28357 $w=3.58e-07 $l=2.9e-07 $layer=LI1_cond $X=2.185 $Y=1.665
+ $X2=2.185 $Y2=1.375
r51 18 24 2.56098 $w=3.58e-07 $l=8e-08 $layer=LI1_cond $X=2.185 $Y=1.295
+ $X2=2.185 $Y2=1.375
r52 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.27 $Y=1.715
+ $X2=2.27 $Y2=1.375
r53 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.715
+ $X2=2.27 $Y2=1.88
r54 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.21
+ $X2=2.27 $Y2=1.375
r55 10 12 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.04 $Y=0.905
+ $X2=2.18 $Y2=0.905
r56 8 17 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=2.36 $Y=2.73 $X2=2.36
+ $Y2=1.88
r57 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.18 $Y=0.98 $X2=2.18
+ $Y2=0.905
r58 4 15 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.18 $Y=0.98 $X2=2.18
+ $Y2=1.21
r59 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.04 $Y=0.83 $X2=2.04
+ $Y2=0.905
r60 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.04 $Y=0.83 $X2=2.04
+ $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_0%C1 3 7 9 10 11 16
c27 16 0 1.79838e-19 $X=2.97 $Y=1.375
r28 16 19 83.3779 $w=4.9e-07 $l=5.05e-07 $layer=POLY_cond $X=2.89 $Y=1.375
+ $X2=2.89 $Y2=1.88
r29 16 18 46.2534 $w=4.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=1.375
+ $X2=2.89 $Y2=1.21
r30 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.97
+ $Y=1.375 $X2=2.97 $Y2=1.375
r31 10 11 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.075 $Y=1.665
+ $X2=3.075 $Y2=2.035
r32 10 17 8.35521 $w=3.98e-07 $l=2.9e-07 $layer=LI1_cond $X=3.075 $Y=1.665
+ $X2=3.075 $Y2=1.375
r33 9 17 2.30489 $w=3.98e-07 $l=8e-08 $layer=LI1_cond $X=3.075 $Y=1.295
+ $X2=3.075 $Y2=1.375
r34 7 18 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=2.81 $Y=0.51 $X2=2.81
+ $Y2=1.21
r35 3 19 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=2.72 $Y=2.73 $X2=2.72
+ $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_0%X 1 2 7 8 9 10 11 12 13 35
r15 32 35 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=0.24 $Y=2.325
+ $X2=0.24 $Y2=2.345
r16 12 32 0.119218 $w=2.88e-07 $l=3e-09 $layer=LI1_cond $X=0.24 $Y=2.322
+ $X2=0.24 $Y2=2.325
r17 12 46 6.01966 $w=2.88e-07 $l=1.42e-07 $layer=LI1_cond $X=0.24 $Y=2.322
+ $X2=0.24 $Y2=2.18
r18 12 13 14.6241 $w=2.88e-07 $l=3.68e-07 $layer=LI1_cond $X=0.24 $Y=2.407
+ $X2=0.24 $Y2=2.775
r19 12 35 2.46384 $w=2.88e-07 $l=6.2e-08 $layer=LI1_cond $X=0.24 $Y=2.407
+ $X2=0.24 $Y2=2.345
r20 11 46 6.96268 $w=2.38e-07 $l=1.45e-07 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=2.18
r21 10 11 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=1.665
+ $X2=0.215 $Y2=2.035
r22 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=1.295
+ $X2=0.215 $Y2=1.665
r23 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=0.925
+ $X2=0.215 $Y2=1.295
r24 8 44 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=0.215 $Y=0.925
+ $X2=0.215 $Y2=0.675
r25 7 44 6.88038 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=0.242 $Y=0.51
+ $X2=0.242 $Y2=0.675
r26 2 35 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.2 $X2=0.26 $Y2=2.345
r27 1 7 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.3 $X2=0.265 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_0%VPWR 1 2 9 13 15 17 22 32 33 36 39
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r45 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 27 39 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.84 $Y=3.33
+ $X2=1.695 $Y2=3.33
r47 27 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.84 $Y=3.33 $X2=2.16
+ $Y2=3.33
r48 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 23 36 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.705 $Y2=3.33
r51 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 22 39 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.695 $Y2=3.33
r53 22 25 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.55 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 17 36 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.705 $Y2=3.33
r57 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 15 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 15 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 11 39 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=3.245
+ $X2=1.695 $Y2=3.33
r62 11 13 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=1.695 $Y=3.245
+ $X2=1.695 $Y2=2.565
r63 7 36 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=3.245
+ $X2=0.705 $Y2=3.33
r64 7 9 34.5733 $w=2.98e-07 $l=9e-07 $layer=LI1_cond $X=0.705 $Y=3.245 $X2=0.705
+ $Y2=2.345
r65 2 13 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=2.41 $X2=1.685 $Y2=2.565
r66 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.2 $X2=0.69 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_0%A_224_482# 1 2 9 11 12 15
c33 9 0 1.47003e-19 $X=1.245 $Y=2.555
r34 13 15 14.1337 $w=2.63e-07 $l=3.25e-07 $layer=LI1_cond $X=2.142 $Y=2.23
+ $X2=2.142 $Y2=2.555
r35 11 13 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=2.01 $Y=2.145
+ $X2=2.142 $Y2=2.23
r36 11 12 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.01 $Y=2.145
+ $X2=1.38 $Y2=2.145
r37 7 12 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.23 $Y=2.23
+ $X2=1.38 $Y2=2.145
r38 7 9 12.4848 $w=2.98e-07 $l=3.25e-07 $layer=LI1_cond $X=1.23 $Y=2.23 $X2=1.23
+ $Y2=2.555
r39 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.005
+ $Y=2.41 $X2=2.145 $Y2=2.555
r40 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.12
+ $Y=2.41 $X2=1.245 $Y2=2.555
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_0%VGND 1 2 7 9 14 21 22 26 33
c40 33 0 1.79838e-19 $X=2.16 $Y=0
c41 22 0 1.26458e-19 $X=3.12 $Y=0
r42 33 36 10.339 $w=5.88e-07 $l=5.1e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.425
+ $Y2=0.51
r43 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 26 29 9.53125 $w=6.38e-07 $l=5.1e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.88
+ $Y2=0.51
r45 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 22 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r47 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 19 33 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.425
+ $Y2=0
r49 19 21 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=3.12
+ $Y2=0
r50 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 17 26 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=0.88
+ $Y2=0
r52 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 14 33 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=2.425
+ $Y2=0
r54 14 17 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=1.2
+ $Y2=0
r55 12 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r56 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 9 26 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.88
+ $Y2=0
r58 9 11 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r59 7 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r60 7 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r61 2 36 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=2.115 $Y=0.3
+ $X2=2.595 $Y2=0.51
r62 1 29 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=0.555 $Y=0.3
+ $X2=1.035 $Y2=0.51
.ends

