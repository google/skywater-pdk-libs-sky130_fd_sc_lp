* File: sky130_fd_sc_lp__o2111ai_1.spice
* Created: Fri Aug 28 11:00:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111ai_1.pex.spice"
.subckt sky130_fd_sc_lp__o2111ai_1  VNB VPB D1 C1 B1 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1002 A_181_47# N_D1_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84 AD=0.1218
+ AS=0.5082 PD=1.13 PS=2.89 NRD=12.852 NRS=48.564 M=1 R=5.6 SA=75000.5
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1003 A_269_47# N_C1_M1003_g A_181_47# VNB NSHORT L=0.15 W=0.84 AD=0.1302
+ AS=0.1218 PD=1.15 PS=1.13 NRD=14.28 NRS=12.852 M=1 R=5.6 SA=75001 SB=75001.8
+ A=0.126 P=1.98 MULT=1
MM1007 N_A_361_47#_M1007_d N_B1_M1007_g A_269_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.168 AS=0.1302 PD=1.24 PS=1.15 NRD=8.568 NRS=14.28 M=1 R=5.6 SA=75001.4
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_361_47#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1764 AS=0.168 PD=1.26 PS=1.24 NRD=9.996 NRS=8.568 M=1 R=5.6 SA=75002
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1008 N_A_361_47#_M1008_d N_A1_M1008_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1764 PD=2.21 PS=1.26 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1009_d N_D1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.3339 PD=1.65 PS=3.05 NRD=8.5892 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_C1_M1005_g N_Y_M1009_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.252 AS=0.2457 PD=1.66 PS=1.65 NRD=9.3772 NRS=8.5892 M=1 R=8.4 SA=75000.7
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.252 PD=1.68 PS=1.66 NRD=10.1455 NRS=9.3772 M=1 R=8.4 SA=75001.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1000 A_513_367# N_A2_M1000_g N_Y_M1006_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.2646 PD=1.47 PS=1.68 NRD=7.8012 NRS=11.7215 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_513_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75002.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o2111ai_1.pxi.spice"
*
.ends
*
*
