# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a31oi_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a31oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.875000 1.425000 6.565000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.930000 1.425000 4.165000 1.760000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.425000 2.725000 1.760000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.750000 1.425000 8.060000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.856400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 0.840000 5.485000 1.050000 ;
        RECT 4.355000 1.050000 6.275000 1.075000 ;
        RECT 4.355000 1.075000 8.065000 1.255000 ;
        RECT 4.355000 1.255000 4.705000 1.950000 ;
        RECT 4.355000 1.950000 7.565000 2.120000 ;
        RECT 5.155000 0.595000 5.485000 0.840000 ;
        RECT 6.075000 0.285000 6.275000 1.050000 ;
        RECT 6.375000 2.120000 6.705000 2.735000 ;
        RECT 6.945000 0.285000 7.135000 1.075000 ;
        RECT 7.235000 2.120000 7.565000 2.735000 ;
        RECT 7.815000 0.305000 8.065000 1.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.095000  0.325000 0.345000 1.085000 ;
      RECT 0.095000  1.085000 4.105000 1.255000 ;
      RECT 0.165000  1.930000 4.185000 2.100000 ;
      RECT 0.165000  2.100000 0.425000 3.075000 ;
      RECT 0.525000  0.085000 0.855000 0.915000 ;
      RECT 0.595000  2.270000 0.925000 3.245000 ;
      RECT 1.025000  0.325000 1.215000 1.085000 ;
      RECT 1.095000  2.100000 1.285000 3.075000 ;
      RECT 1.385000  0.085000 1.715000 0.915000 ;
      RECT 1.455000  2.270000 1.785000 3.245000 ;
      RECT 1.885000  0.325000 2.075000 1.085000 ;
      RECT 1.955000  2.100000 2.145000 3.075000 ;
      RECT 2.245000  0.255000 5.855000 0.425000 ;
      RECT 2.245000  0.425000 2.575000 0.915000 ;
      RECT 2.315000  2.270000 2.645000 3.245000 ;
      RECT 2.755000  0.595000 3.085000 1.085000 ;
      RECT 2.815000  2.100000 3.005000 3.075000 ;
      RECT 3.175000  2.270000 3.845000 2.640000 ;
      RECT 3.175000  2.640000 4.015000 3.245000 ;
      RECT 3.265000  0.425000 3.595000 0.915000 ;
      RECT 3.775000  0.595000 4.105000 1.085000 ;
      RECT 4.015000  2.100000 4.185000 2.290000 ;
      RECT 4.015000  2.290000 6.205000 2.460000 ;
      RECT 4.015000  2.460000 4.405000 2.470000 ;
      RECT 4.185000  2.470000 4.405000 3.075000 ;
      RECT 4.575000  2.630000 4.905000 3.245000 ;
      RECT 4.725000  0.425000 4.985000 0.670000 ;
      RECT 5.075000  2.460000 5.265000 3.075000 ;
      RECT 5.435000  2.630000 5.765000 3.245000 ;
      RECT 5.655000  0.425000 5.855000 0.880000 ;
      RECT 5.935000  2.460000 6.205000 2.905000 ;
      RECT 5.935000  2.905000 7.995000 3.075000 ;
      RECT 6.445000  0.085000 6.775000 0.905000 ;
      RECT 6.875000  2.290000 7.065000 2.905000 ;
      RECT 7.305000  0.085000 7.635000 0.905000 ;
      RECT 7.745000  1.950000 7.995000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__a31oi_4
