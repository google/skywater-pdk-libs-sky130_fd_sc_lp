* File: sky130_fd_sc_lp__a211oi_4.pxi.spice
* Created: Fri Aug 28 09:48:31 2020
* 
x_PM_SKY130_FD_SC_LP__A211OI_4%A2 N_A2_M1006_g N_A2_c_126_n N_A2_M1004_g
+ N_A2_M1008_g N_A2_c_127_n N_A2_M1009_g N_A2_M1023_g N_A2_c_128_n N_A2_M1012_g
+ N_A2_M1026_g N_A2_M1018_g N_A2_c_120_n N_A2_c_121_n N_A2_c_122_n N_A2_c_123_n
+ N_A2_c_124_n A2 A2 A2 N_A2_c_125_n PM_SKY130_FD_SC_LP__A211OI_4%A2
x_PM_SKY130_FD_SC_LP__A211OI_4%A1 N_A1_c_226_n N_A1_M1002_g N_A1_M1005_g
+ N_A1_c_228_n N_A1_M1003_g N_A1_M1016_g N_A1_c_230_n N_A1_M1015_g N_A1_M1025_g
+ N_A1_c_232_n N_A1_M1024_g N_A1_M1027_g A1 A1 A1 N_A1_c_235_n
+ PM_SKY130_FD_SC_LP__A211OI_4%A1
x_PM_SKY130_FD_SC_LP__A211OI_4%B1 N_B1_c_302_n N_B1_M1011_g N_B1_M1007_g
+ N_B1_c_304_n N_B1_M1020_g N_B1_M1017_g N_B1_c_306_n N_B1_M1029_g N_B1_M1019_g
+ N_B1_M1031_g N_B1_M1028_g N_B1_c_309_n N_B1_c_310_n N_B1_c_311_n B1 B1 B1
+ N_B1_c_312_n N_B1_c_313_n N_B1_c_314_n N_B1_c_315_n
+ PM_SKY130_FD_SC_LP__A211OI_4%B1
x_PM_SKY130_FD_SC_LP__A211OI_4%C1 N_C1_M1000_g N_C1_M1010_g N_C1_M1001_g
+ N_C1_M1013_g N_C1_M1014_g N_C1_M1021_g N_C1_M1022_g N_C1_M1030_g N_C1_c_423_n
+ C1 C1 N_C1_c_424_n N_C1_c_430_n C1 N_C1_c_431_n
+ PM_SKY130_FD_SC_LP__A211OI_4%C1
x_PM_SKY130_FD_SC_LP__A211OI_4%A_45_367# N_A_45_367#_M1004_s N_A_45_367#_M1009_s
+ N_A_45_367#_M1005_d N_A_45_367#_M1025_d N_A_45_367#_M1018_s
+ N_A_45_367#_M1017_d N_A_45_367#_M1028_d N_A_45_367#_c_513_n
+ N_A_45_367#_c_514_n N_A_45_367#_c_521_n N_A_45_367#_c_573_p
+ N_A_45_367#_c_525_n N_A_45_367#_c_570_p N_A_45_367#_c_527_n
+ N_A_45_367#_c_571_p N_A_45_367#_c_528_n N_A_45_367#_c_515_n
+ N_A_45_367#_c_535_n N_A_45_367#_c_516_n N_A_45_367#_c_550_n
+ N_A_45_367#_c_598_p N_A_45_367#_c_517_n N_A_45_367#_c_518_n
+ N_A_45_367#_c_536_n N_A_45_367#_c_538_n N_A_45_367#_c_539_n
+ PM_SKY130_FD_SC_LP__A211OI_4%A_45_367#
x_PM_SKY130_FD_SC_LP__A211OI_4%VPWR N_VPWR_M1004_d N_VPWR_M1012_d N_VPWR_M1016_s
+ N_VPWR_M1027_s N_VPWR_c_607_n N_VPWR_c_608_n N_VPWR_c_609_n N_VPWR_c_610_n
+ N_VPWR_c_611_n N_VPWR_c_612_n N_VPWR_c_613_n N_VPWR_c_614_n VPWR
+ N_VPWR_c_615_n N_VPWR_c_616_n N_VPWR_c_617_n N_VPWR_c_606_n N_VPWR_c_619_n
+ N_VPWR_c_620_n PM_SKY130_FD_SC_LP__A211OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A211OI_4%A_826_367# N_A_826_367#_M1007_s
+ N_A_826_367#_M1019_s N_A_826_367#_M1013_d N_A_826_367#_M1030_d
+ N_A_826_367#_c_724_n N_A_826_367#_c_716_n N_A_826_367#_c_706_n
+ PM_SKY130_FD_SC_LP__A211OI_4%A_826_367#
x_PM_SKY130_FD_SC_LP__A211OI_4%Y N_Y_M1002_d N_Y_M1015_d N_Y_M1011_s N_Y_M1029_s
+ N_Y_M1001_s N_Y_M1022_s N_Y_M1010_s N_Y_M1021_s N_Y_c_737_n N_Y_c_749_n
+ N_Y_c_753_n N_Y_c_755_n N_Y_c_756_n N_Y_c_796_n N_Y_c_757_n N_Y_c_734_n
+ N_Y_c_762_n N_Y_c_732_n N_Y_c_733_n N_Y_c_770_n N_Y_c_772_n N_Y_c_736_n
+ N_Y_c_774_n Y Y N_Y_c_738_n N_Y_c_782_n Y N_Y_c_784_n
+ PM_SKY130_FD_SC_LP__A211OI_4%Y
x_PM_SKY130_FD_SC_LP__A211OI_4%VGND N_VGND_M1006_d N_VGND_M1008_d N_VGND_M1026_d
+ N_VGND_M1020_d N_VGND_M1000_d N_VGND_M1014_d N_VGND_M1031_d N_VGND_c_874_n
+ N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n N_VGND_c_879_n
+ N_VGND_c_880_n N_VGND_c_881_n N_VGND_c_882_n N_VGND_c_883_n N_VGND_c_884_n
+ N_VGND_c_885_n N_VGND_c_886_n VGND N_VGND_c_887_n N_VGND_c_888_n
+ N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n
+ N_VGND_c_894_n PM_SKY130_FD_SC_LP__A211OI_4%VGND
x_PM_SKY130_FD_SC_LP__A211OI_4%A_114_47# N_A_114_47#_M1006_s N_A_114_47#_M1023_s
+ N_A_114_47#_M1003_s N_A_114_47#_M1024_s N_A_114_47#_c_1024_n
+ N_A_114_47#_c_1000_n N_A_114_47#_c_1001_n N_A_114_47#_c_1029_n
+ N_A_114_47#_c_1011_n PM_SKY130_FD_SC_LP__A211OI_4%A_114_47#
cc_1 VNB N_A2_M1006_g 0.0303822f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_2 VNB N_A2_M1008_g 0.0207302f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_3 VNB N_A2_M1023_g 0.0209089f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_4 VNB N_A2_M1026_g 0.022222f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=0.655
cc_5 VNB N_A2_M1018_g 0.00246836f $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=2.465
cc_6 VNB N_A2_c_120_n 0.00979837f $X=-0.19 $Y=-0.245 $X2=3.385 $Y2=1.7
cc_7 VNB N_A2_c_121_n 0.0125848f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.565
cc_8 VNB N_A2_c_122_n 0.00414641f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.565
cc_9 VNB N_A2_c_123_n 0.00711214f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.44
cc_10 VNB N_A2_c_124_n 0.0291039f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.44
cc_11 VNB N_A2_c_125_n 0.0834601f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.51
cc_12 VNB N_A1_c_226_n 0.0163563f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.295
cc_13 VNB N_A1_M1005_g 0.00692979f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.465
cc_14 VNB N_A1_c_228_n 0.016096f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.295
cc_15 VNB N_A1_M1016_g 0.00672302f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.465
cc_16 VNB N_A1_c_230_n 0.0161006f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.295
cc_17 VNB N_A1_M1025_g 0.00672351f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.465
cc_18 VNB N_A1_c_232_n 0.0163339f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.275
cc_19 VNB N_A1_M1027_g 0.00672313f $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=2.465
cc_20 VNB A1 0.00994797f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.7
cc_21 VNB N_A1_c_235_n 0.0822154f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.51
cc_22 VNB N_B1_c_302_n 0.0173848f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.295
cc_23 VNB N_B1_M1007_g 0.00708397f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.465
cc_24 VNB N_B1_c_304_n 0.0159959f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.295
cc_25 VNB N_B1_M1017_g 0.00706879f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.465
cc_26 VNB N_B1_c_306_n 0.0158746f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.295
cc_27 VNB N_B1_M1019_g 0.0072382f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.465
cc_28 VNB N_B1_M1028_g 0.00816598f $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=2.465
cc_29 VNB N_B1_c_309_n 0.0246274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B1_c_310_n 0.00319455f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.7
cc_31 VNB N_B1_c_311_n 0.0351341f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.44
cc_32 VNB N_B1_c_312_n 0.0552944f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.46
cc_33 VNB N_B1_c_313_n 0.0196933f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.44
cc_34 VNB N_B1_c_314_n 0.00122075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B1_c_315_n 0.0115546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_C1_M1000_g 0.0230646f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_37 VNB N_C1_M1001_g 0.0229169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_C1_M1014_g 0.0229376f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.725
cc_39 VNB N_C1_M1022_g 0.0231597f $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=2.465
cc_40 VNB N_C1_c_423_n 0.00227206f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_41 VNB N_C1_c_424_n 0.0656779f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.605
cc_42 VNB N_VPWR_c_606_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_43 VNB N_Y_c_732_n 0.0110697f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.46
cc_44 VNB N_Y_c_733_n 0.035571f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.44
cc_45 VNB N_VGND_c_874_n 0.0116397f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.275
cc_46 VNB N_VGND_c_875_n 0.0398592f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=0.655
cc_47 VNB N_VGND_c_876_n 4.04385e-19 $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=2.465
cc_48 VNB N_VGND_c_877_n 0.00223571f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.565
cc_49 VNB N_VGND_c_878_n 0.0150706f $X=-0.19 $Y=-0.245 $X2=3.572 $Y2=1.44
cc_50 VNB N_VGND_c_879_n 0.00180145f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_51 VNB N_VGND_c_880_n 0.016693f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_52 VNB N_VGND_c_881_n 0.003699f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=1.51
cc_53 VNB N_VGND_c_882_n 0.003699f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.51
cc_54 VNB N_VGND_c_883_n 0.0144677f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.51
cc_55 VNB N_VGND_c_884_n 0.0175966f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.46
cc_56 VNB N_VGND_c_885_n 0.0167176f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.51
cc_57 VNB N_VGND_c_886_n 0.00362148f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.44
cc_58 VNB N_VGND_c_887_n 0.0146078f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_59 VNB N_VGND_c_888_n 0.0503823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_889_n 0.0167176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_890_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_891_n 0.00510459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_892_n 0.00375705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_893_n 0.00362148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_894_n 0.369885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_114_47#_c_1000_n 0.00644838f $X=-0.19 $Y=-0.245 $X2=1.355
+ $Y2=0.655
cc_67 VNB N_A_114_47#_c_1001_n 0.0029808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VPB N_A2_c_126_n 0.0205699f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.725
cc_69 VPB N_A2_c_127_n 0.0155213f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=1.725
cc_70 VPB N_A2_c_128_n 0.0156216f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.725
cc_71 VPB N_A2_M1018_g 0.0203235f $X=-0.19 $Y=1.655 $X2=3.625 $Y2=2.465
cc_72 VPB N_A2_c_120_n 0.0104693f $X=-0.19 $Y=1.655 $X2=3.385 $Y2=1.7
cc_73 VPB N_A2_c_121_n 0.0158326f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.565
cc_74 VPB N_A2_c_122_n 0.00135408f $X=-0.19 $Y=1.655 $X2=1.645 $Y2=1.565
cc_75 VPB N_A2_c_123_n 0.00154208f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=1.44
cc_76 VPB N_A2_c_125_n 0.02946f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.51
cc_77 VPB N_A1_M1005_g 0.0186439f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.465
cc_78 VPB N_A1_M1016_g 0.0185384f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=2.465
cc_79 VPB N_A1_M1025_g 0.0185384f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=2.465
cc_80 VPB N_A1_M1027_g 0.0192323f $X=-0.19 $Y=1.655 $X2=3.625 $Y2=2.465
cc_81 VPB N_B1_M1007_g 0.0188405f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.465
cc_82 VPB N_B1_M1017_g 0.018695f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=2.465
cc_83 VPB N_B1_M1019_g 0.0201142f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=2.465
cc_84 VPB N_B1_M1028_g 0.0238645f $X=-0.19 $Y=1.655 $X2=3.625 $Y2=2.465
cc_85 VPB N_C1_M1010_g 0.0186966f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.465
cc_86 VPB N_C1_M1013_g 0.0180114f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.295
cc_87 VPB N_C1_M1021_g 0.0183567f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=0.655
cc_88 VPB N_C1_M1030_g 0.018829f $X=-0.19 $Y=1.655 $X2=1.645 $Y2=1.7
cc_89 VPB N_C1_c_424_n 0.0123221f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=1.605
cc_90 VPB N_C1_c_430_n 0.00375605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_C1_c_431_n 0.00144106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_45_367#_c_513_n 0.0074281f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=1.275
cc_93 VPB N_A_45_367#_c_514_n 0.0360021f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=0.655
cc_94 VPB N_A_45_367#_c_515_n 0.00882678f $X=-0.19 $Y=1.655 $X2=0.285 $Y2=1.46
cc_95 VPB N_A_45_367#_c_516_n 0.00691676f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=1.51
cc_96 VPB N_A_45_367#_c_517_n 0.0171381f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=1.605
cc_97 VPB N_A_45_367#_c_518_n 0.0188366f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_607_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.295
cc_99 VPB N_VPWR_c_608_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.725
cc_100 VPB N_VPWR_c_609_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=3.505 $Y2=0.655
cc_101 VPB N_VPWR_c_610_n 0.00269808f $X=-0.19 $Y=1.655 $X2=3.625 $Y2=2.465
cc_102 VPB N_VPWR_c_611_n 0.0129398f $X=-0.19 $Y=1.655 $X2=3.385 $Y2=1.7
cc_103 VPB N_VPWR_c_612_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.645 $Y2=1.7
cc_104 VPB N_VPWR_c_613_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.645 $Y2=1.565
cc_105 VPB N_VPWR_c_614_n 0.00510509f $X=-0.19 $Y=1.655 $X2=3.572 $Y2=1.44
cc_106 VPB N_VPWR_c_615_n 0.0182398f $X=-0.19 $Y=1.655 $X2=3.385 $Y2=1.7
cc_107 VPB N_VPWR_c_616_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_617_n 0.101229f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=1.605
cc_109 VPB N_VPWR_c_606_n 0.054076f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.565
cc_110 VPB N_VPWR_c_619_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.285 $Y2=1.565
cc_111 VPB N_VPWR_c_620_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.565
cc_112 VPB N_Y_c_734_n 0.0221367f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.51
cc_113 VPB N_Y_c_733_n 0.0080893f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=1.44
cc_114 VPB N_Y_c_736_n 0.00211871f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.565
cc_115 N_A2_M1023_g N_A1_c_226_n 0.0216329f $X=1.355 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A2_c_120_n N_A1_M1005_g 0.0121258f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_117 N_A2_c_125_n N_A1_M1005_g 0.0420027f $X=1.355 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A2_c_120_n N_A1_M1016_g 0.0104926f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_119 N_A2_c_120_n N_A1_M1025_g 0.0104926f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_120 N_A2_M1026_g N_A1_c_232_n 0.0339739f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_121 N_A2_M1018_g N_A1_M1027_g 0.0328896f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A2_c_120_n N_A1_M1027_g 0.0108404f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_123 N_A2_M1023_g A1 5.46055e-19 $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_124 N_A2_M1026_g A1 0.00260553f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_125 N_A2_c_120_n A1 0.0992879f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_126 N_A2_c_122_n A1 0.0080292f $X=1.645 $Y=1.565 $X2=0 $Y2=0
cc_127 N_A2_c_123_n A1 0.0146163f $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_128 N_A2_c_125_n A1 3.8895e-19 $X=1.355 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A2_M1026_g N_A1_c_235_n 0.00927116f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_130 N_A2_c_120_n N_A1_c_235_n 0.0107818f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_131 N_A2_c_122_n N_A1_c_235_n 0.00597338f $X=1.645 $Y=1.565 $X2=0 $Y2=0
cc_132 N_A2_c_123_n N_A1_c_235_n 0.00467357f $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_133 N_A2_c_124_n N_A1_c_235_n 0.0152234f $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_134 N_A2_c_125_n N_A1_c_235_n 0.0120781f $X=1.355 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A2_M1026_g N_B1_c_302_n 0.0302003f $X=3.505 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A2_M1018_g N_B1_M1007_g 0.0222767f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A2_c_123_n N_B1_M1007_g 8.25545e-19 $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_138 N_A2_c_123_n N_B1_c_312_n 6.51285e-19 $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_139 N_A2_c_124_n N_B1_c_312_n 0.0205965f $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_140 N_A2_M1026_g N_B1_c_314_n 3.36652e-19 $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_141 N_A2_c_123_n N_B1_c_314_n 0.0160652f $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_142 N_A2_c_124_n N_B1_c_314_n 2.99365e-19 $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_143 N_A2_c_121_n N_A_45_367#_c_513_n 0.0225542f $X=1.425 $Y=1.565 $X2=0 $Y2=0
cc_144 N_A2_c_125_n N_A_45_367#_c_513_n 0.00171925f $X=1.355 $Y=1.51 $X2=0 $Y2=0
cc_145 N_A2_c_126_n N_A_45_367#_c_521_n 0.0122595f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_146 N_A2_c_127_n N_A_45_367#_c_521_n 0.0122595f $X=0.995 $Y=1.725 $X2=0 $Y2=0
cc_147 N_A2_c_121_n N_A_45_367#_c_521_n 0.0439805f $X=1.425 $Y=1.565 $X2=0 $Y2=0
cc_148 N_A2_c_125_n N_A_45_367#_c_521_n 5.937e-19 $X=1.355 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A2_c_128_n N_A_45_367#_c_525_n 0.0122129f $X=1.425 $Y=1.725 $X2=0 $Y2=0
cc_150 N_A2_c_121_n N_A_45_367#_c_525_n 0.042487f $X=1.425 $Y=1.565 $X2=0 $Y2=0
cc_151 N_A2_c_120_n N_A_45_367#_c_527_n 0.0402256f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_152 N_A2_M1018_g N_A_45_367#_c_528_n 0.0140754f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A2_c_120_n N_A_45_367#_c_528_n 0.0223559f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_154 N_A2_c_123_n N_A_45_367#_c_528_n 0.0164233f $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_155 N_A2_c_124_n N_A_45_367#_c_528_n 4.54826e-19 $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_156 N_A2_M1018_g N_A_45_367#_c_515_n 0.00234732f $X=3.625 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A2_c_123_n N_A_45_367#_c_515_n 0.009699f $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_158 N_A2_c_124_n N_A_45_367#_c_515_n 6.33571e-19 $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_159 N_A2_M1018_g N_A_45_367#_c_535_n 0.0114257f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A2_c_121_n N_A_45_367#_c_536_n 0.015747f $X=1.425 $Y=1.565 $X2=0 $Y2=0
cc_161 N_A2_c_125_n N_A_45_367#_c_536_n 6.70625e-19 $X=1.355 $Y=1.51 $X2=0 $Y2=0
cc_162 N_A2_c_120_n N_A_45_367#_c_538_n 0.0146339f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_163 N_A2_c_120_n N_A_45_367#_c_539_n 0.0146339f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_164 N_A2_c_126_n N_VPWR_c_607_n 0.0159947f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_165 N_A2_c_127_n N_VPWR_c_607_n 0.0141241f $X=0.995 $Y=1.725 $X2=0 $Y2=0
cc_166 N_A2_c_128_n N_VPWR_c_607_n 6.7059e-19 $X=1.425 $Y=1.725 $X2=0 $Y2=0
cc_167 N_A2_c_127_n N_VPWR_c_608_n 6.7059e-19 $X=0.995 $Y=1.725 $X2=0 $Y2=0
cc_168 N_A2_c_128_n N_VPWR_c_608_n 0.014044f $X=1.425 $Y=1.725 $X2=0 $Y2=0
cc_169 N_A2_M1018_g N_VPWR_c_610_n 0.00404015f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A2_c_126_n N_VPWR_c_615_n 0.00486043f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_171 N_A2_c_127_n N_VPWR_c_616_n 0.00486043f $X=0.995 $Y=1.725 $X2=0 $Y2=0
cc_172 N_A2_c_128_n N_VPWR_c_616_n 0.00486043f $X=1.425 $Y=1.725 $X2=0 $Y2=0
cc_173 N_A2_M1018_g N_VPWR_c_617_n 0.00579312f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A2_c_126_n N_VPWR_c_606_n 0.00925455f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_175 N_A2_c_127_n N_VPWR_c_606_n 0.00824727f $X=0.995 $Y=1.725 $X2=0 $Y2=0
cc_176 N_A2_c_128_n N_VPWR_c_606_n 0.00824727f $X=1.425 $Y=1.725 $X2=0 $Y2=0
cc_177 N_A2_M1018_g N_VPWR_c_606_n 0.0105917f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A2_M1026_g N_Y_c_737_n 5.38418e-19 $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_179 N_A2_M1026_g N_Y_c_738_n 0.0165399f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_180 N_A2_c_120_n N_Y_c_738_n 0.0038797f $X=3.385 $Y=1.7 $X2=0 $Y2=0
cc_181 N_A2_c_123_n N_Y_c_738_n 0.0184933f $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_182 N_A2_c_124_n N_Y_c_738_n 0.00101829f $X=3.595 $Y=1.44 $X2=0 $Y2=0
cc_183 N_A2_M1006_g N_VGND_c_875_n 0.00712852f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_184 N_A2_c_121_n N_VGND_c_875_n 0.018958f $X=1.425 $Y=1.565 $X2=0 $Y2=0
cc_185 N_A2_c_125_n N_VGND_c_875_n 0.00732517f $X=1.355 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A2_M1006_g N_VGND_c_876_n 6.26215e-19 $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_187 N_A2_M1008_g N_VGND_c_876_n 0.0102463f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A2_M1023_g N_VGND_c_876_n 0.0113462f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A2_M1026_g N_VGND_c_877_n 0.00921419f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_190 N_A2_M1006_g N_VGND_c_887_n 0.00585385f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A2_M1008_g N_VGND_c_887_n 0.00486043f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A2_M1023_g N_VGND_c_888_n 0.00486043f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A2_M1026_g N_VGND_c_888_n 0.00367409f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A2_M1006_g N_VGND_c_894_n 0.0114597f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A2_M1008_g N_VGND_c_894_n 0.00824727f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A2_M1023_g N_VGND_c_894_n 0.0082726f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_197 N_A2_M1026_g N_VGND_c_894_n 0.00438943f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_198 N_A2_M1008_g N_A_114_47#_c_1000_n 0.0131979f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_199 N_A2_M1023_g N_A_114_47#_c_1000_n 0.0131442f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_200 N_A2_c_121_n N_A_114_47#_c_1000_n 0.0502727f $X=1.425 $Y=1.565 $X2=0
+ $Y2=0
cc_201 N_A2_c_122_n N_A_114_47#_c_1000_n 0.0153543f $X=1.645 $Y=1.565 $X2=0
+ $Y2=0
cc_202 N_A2_c_125_n N_A_114_47#_c_1000_n 0.00396262f $X=1.355 $Y=1.51 $X2=0
+ $Y2=0
cc_203 N_A2_M1006_g N_A_114_47#_c_1001_n 0.00283166f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_204 N_A2_c_121_n N_A_114_47#_c_1001_n 0.0189283f $X=1.425 $Y=1.565 $X2=0
+ $Y2=0
cc_205 N_A2_c_125_n N_A_114_47#_c_1001_n 0.00280626f $X=1.355 $Y=1.51 $X2=0
+ $Y2=0
cc_206 N_A1_M1005_g N_A_45_367#_c_525_n 0.0122129f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A1_M1016_g N_A_45_367#_c_527_n 0.0122595f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A1_M1025_g N_A_45_367#_c_527_n 0.0122595f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A1_M1027_g N_A_45_367#_c_528_n 0.0124907f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A1_M1027_g N_A_45_367#_c_535_n 5.95673e-19 $X=3.145 $Y=2.465 $X2=0
+ $Y2=0
cc_211 N_A1_M1005_g N_VPWR_c_608_n 0.014044f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A1_M1016_g N_VPWR_c_608_n 6.7059e-19 $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A1_M1005_g N_VPWR_c_609_n 6.7059e-19 $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A1_M1016_g N_VPWR_c_609_n 0.0142444f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A1_M1025_g N_VPWR_c_609_n 0.0142444f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A1_M1027_g N_VPWR_c_609_n 6.7059e-19 $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A1_M1025_g N_VPWR_c_610_n 6.7059e-19 $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A1_M1027_g N_VPWR_c_610_n 0.014138f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A1_M1005_g N_VPWR_c_611_n 0.00486043f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A1_M1016_g N_VPWR_c_611_n 0.00486043f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A1_M1025_g N_VPWR_c_613_n 0.00486043f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A1_M1027_g N_VPWR_c_613_n 0.00486043f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A1_M1005_g N_VPWR_c_606_n 0.00824727f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A1_M1016_g N_VPWR_c_606_n 0.00824727f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A1_M1025_g N_VPWR_c_606_n 0.00824727f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A1_M1027_g N_VPWR_c_606_n 0.00824727f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_227 N_A1_c_226_n N_Y_c_738_n 0.00320348f $X=1.785 $Y=1.185 $X2=0 $Y2=0
cc_228 N_A1_c_228_n N_Y_c_738_n 0.0107125f $X=2.215 $Y=1.185 $X2=0 $Y2=0
cc_229 N_A1_c_230_n N_Y_c_738_n 0.0107125f $X=2.645 $Y=1.185 $X2=0 $Y2=0
cc_230 N_A1_c_232_n N_Y_c_738_n 0.0106424f $X=3.075 $Y=1.185 $X2=0 $Y2=0
cc_231 A1 N_Y_c_738_n 0.0894862f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_232 N_A1_c_235_n N_Y_c_738_n 0.00249708f $X=3.075 $Y=1.35 $X2=0 $Y2=0
cc_233 N_A1_c_226_n N_VGND_c_876_n 0.00109252f $X=1.785 $Y=1.185 $X2=0 $Y2=0
cc_234 N_A1_c_232_n N_VGND_c_877_n 0.00109496f $X=3.075 $Y=1.185 $X2=0 $Y2=0
cc_235 N_A1_c_226_n N_VGND_c_888_n 0.00357877f $X=1.785 $Y=1.185 $X2=0 $Y2=0
cc_236 N_A1_c_228_n N_VGND_c_888_n 0.00357877f $X=2.215 $Y=1.185 $X2=0 $Y2=0
cc_237 N_A1_c_230_n N_VGND_c_888_n 0.00357877f $X=2.645 $Y=1.185 $X2=0 $Y2=0
cc_238 N_A1_c_232_n N_VGND_c_888_n 0.00357877f $X=3.075 $Y=1.185 $X2=0 $Y2=0
cc_239 N_A1_c_226_n N_VGND_c_894_n 0.00537654f $X=1.785 $Y=1.185 $X2=0 $Y2=0
cc_240 N_A1_c_228_n N_VGND_c_894_n 0.0053512f $X=2.215 $Y=1.185 $X2=0 $Y2=0
cc_241 N_A1_c_230_n N_VGND_c_894_n 0.0053512f $X=2.645 $Y=1.185 $X2=0 $Y2=0
cc_242 N_A1_c_232_n N_VGND_c_894_n 0.00537654f $X=3.075 $Y=1.185 $X2=0 $Y2=0
cc_243 N_A1_c_226_n N_A_114_47#_c_1000_n 0.00317585f $X=1.785 $Y=1.185 $X2=0
+ $Y2=0
cc_244 N_A1_c_226_n N_A_114_47#_c_1011_n 0.0160765f $X=1.785 $Y=1.185 $X2=0
+ $Y2=0
cc_245 N_A1_c_228_n N_A_114_47#_c_1011_n 0.0118112f $X=2.215 $Y=1.185 $X2=0
+ $Y2=0
cc_246 N_A1_c_230_n N_A_114_47#_c_1011_n 0.0118112f $X=2.645 $Y=1.185 $X2=0
+ $Y2=0
cc_247 N_A1_c_232_n N_A_114_47#_c_1011_n 0.0119021f $X=3.075 $Y=1.185 $X2=0
+ $Y2=0
cc_248 N_B1_c_306_n N_C1_M1000_g 0.0173611f $X=4.905 $Y=1.185 $X2=0 $Y2=0
cc_249 N_B1_c_309_n N_C1_M1000_g 0.0131381f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_250 N_B1_c_312_n N_C1_M1000_g 0.0119099f $X=4.905 $Y=1.35 $X2=0 $Y2=0
cc_251 N_B1_c_315_n N_C1_M1000_g 0.00616608f $X=5.18 $Y=1.3 $X2=0 $Y2=0
cc_252 N_B1_M1019_g N_C1_M1010_g 0.0534654f $X=4.915 $Y=2.465 $X2=0 $Y2=0
cc_253 N_B1_c_309_n N_C1_M1001_g 0.0104915f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_254 N_B1_c_309_n N_C1_M1014_g 0.010445f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_255 N_B1_c_309_n N_C1_M1022_g 0.0104313f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_256 N_B1_c_310_n N_C1_M1022_g 6.79925e-19 $X=7.11 $Y=1.17 $X2=0 $Y2=0
cc_257 N_B1_c_313_n N_C1_M1022_g 0.0248915f $X=7.145 $Y=1.185 $X2=0 $Y2=0
cc_258 N_B1_M1028_g N_C1_c_423_n 7.98556e-19 $X=7.065 $Y=2.465 $X2=0 $Y2=0
cc_259 N_B1_c_310_n N_C1_c_423_n 0.00481725f $X=7.11 $Y=1.17 $X2=0 $Y2=0
cc_260 N_B1_c_311_n N_C1_c_423_n 3.41346e-19 $X=7.145 $Y=1.35 $X2=0 $Y2=0
cc_261 N_B1_M1019_g N_C1_c_424_n 0.0119099f $X=4.915 $Y=2.465 $X2=0 $Y2=0
cc_262 N_B1_M1028_g N_C1_c_424_n 0.0617309f $X=7.065 $Y=2.465 $X2=0 $Y2=0
cc_263 N_B1_c_309_n N_C1_c_424_n 0.00781256f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_264 N_B1_c_310_n N_C1_c_424_n 7.20151e-19 $X=7.11 $Y=1.17 $X2=0 $Y2=0
cc_265 N_B1_c_311_n N_C1_c_424_n 0.00856044f $X=7.145 $Y=1.35 $X2=0 $Y2=0
cc_266 N_B1_c_309_n N_C1_c_430_n 0.0990958f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_267 N_B1_c_312_n N_C1_c_430_n 0.0012497f $X=4.905 $Y=1.35 $X2=0 $Y2=0
cc_268 N_B1_c_315_n N_C1_c_430_n 0.00784469f $X=5.18 $Y=1.3 $X2=0 $Y2=0
cc_269 N_B1_M1007_g N_A_45_367#_c_516_n 0.014305f $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_270 N_B1_M1017_g N_A_45_367#_c_516_n 0.014305f $X=4.485 $Y=2.465 $X2=0 $Y2=0
cc_271 N_B1_M1019_g N_A_45_367#_c_516_n 0.00317938f $X=4.915 $Y=2.465 $X2=0
+ $Y2=0
cc_272 N_B1_c_312_n N_A_45_367#_c_516_n 0.0049322f $X=4.905 $Y=1.35 $X2=0 $Y2=0
cc_273 N_B1_c_314_n N_A_45_367#_c_516_n 0.0572923f $X=4.895 $Y=1.3 $X2=0 $Y2=0
cc_274 N_B1_M1019_g N_A_45_367#_c_550_n 0.0159045f $X=4.915 $Y=2.465 $X2=0 $Y2=0
cc_275 N_B1_M1028_g N_A_45_367#_c_550_n 0.0129371f $X=7.065 $Y=2.465 $X2=0 $Y2=0
cc_276 N_B1_M1028_g N_A_45_367#_c_517_n 0.00279257f $X=7.065 $Y=2.465 $X2=0
+ $Y2=0
cc_277 N_B1_M1028_g N_A_45_367#_c_518_n 0.00554108f $X=7.065 $Y=2.465 $X2=0
+ $Y2=0
cc_278 N_B1_M1007_g N_VPWR_c_617_n 0.00585385f $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_279 N_B1_M1017_g N_VPWR_c_617_n 0.00357877f $X=4.485 $Y=2.465 $X2=0 $Y2=0
cc_280 N_B1_M1019_g N_VPWR_c_617_n 0.00357877f $X=4.915 $Y=2.465 $X2=0 $Y2=0
cc_281 N_B1_M1028_g N_VPWR_c_617_n 0.00440697f $X=7.065 $Y=2.465 $X2=0 $Y2=0
cc_282 N_B1_M1007_g N_VPWR_c_606_n 0.0107906f $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_283 N_B1_M1017_g N_VPWR_c_606_n 0.0053512f $X=4.485 $Y=2.465 $X2=0 $Y2=0
cc_284 N_B1_M1019_g N_VPWR_c_606_n 0.00537654f $X=4.915 $Y=2.465 $X2=0 $Y2=0
cc_285 N_B1_M1028_g N_VPWR_c_606_n 0.00717334f $X=7.065 $Y=2.465 $X2=0 $Y2=0
cc_286 N_B1_M1017_g N_A_826_367#_c_706_n 0.0169181f $X=4.485 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_B1_M1019_g N_A_826_367#_c_706_n 0.0118112f $X=4.915 $Y=2.465 $X2=0
+ $Y2=0
cc_288 N_B1_c_302_n N_Y_c_737_n 0.00828106f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_289 N_B1_c_306_n N_Y_c_749_n 0.00959712f $X=4.905 $Y=1.185 $X2=0 $Y2=0
cc_290 N_B1_c_312_n N_Y_c_749_n 3.15467e-19 $X=4.905 $Y=1.35 $X2=0 $Y2=0
cc_291 N_B1_c_314_n N_Y_c_749_n 0.00663174f $X=4.895 $Y=1.3 $X2=0 $Y2=0
cc_292 N_B1_c_315_n N_Y_c_749_n 0.00437842f $X=5.18 $Y=1.3 $X2=0 $Y2=0
cc_293 N_B1_c_304_n N_Y_c_753_n 4.4915e-19 $X=4.475 $Y=1.185 $X2=0 $Y2=0
cc_294 N_B1_c_306_n N_Y_c_753_n 0.00671598f $X=4.905 $Y=1.185 $X2=0 $Y2=0
cc_295 N_B1_c_309_n N_Y_c_755_n 0.033448f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_296 N_B1_M1019_g N_Y_c_756_n 6.24983e-19 $X=4.915 $Y=2.465 $X2=0 $Y2=0
cc_297 N_B1_c_309_n N_Y_c_757_n 0.033448f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_298 N_B1_M1028_g N_Y_c_734_n 0.0137731f $X=7.065 $Y=2.465 $X2=0 $Y2=0
cc_299 N_B1_c_309_n N_Y_c_734_n 0.0088927f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_300 N_B1_c_310_n N_Y_c_734_n 0.0124059f $X=7.11 $Y=1.17 $X2=0 $Y2=0
cc_301 N_B1_c_311_n N_Y_c_734_n 0.00299594f $X=7.145 $Y=1.35 $X2=0 $Y2=0
cc_302 N_B1_c_313_n N_Y_c_762_n 0.0112832f $X=7.145 $Y=1.185 $X2=0 $Y2=0
cc_303 N_B1_c_310_n N_Y_c_732_n 0.0157764f $X=7.11 $Y=1.17 $X2=0 $Y2=0
cc_304 N_B1_c_311_n N_Y_c_732_n 0.00288645f $X=7.145 $Y=1.35 $X2=0 $Y2=0
cc_305 N_B1_c_313_n N_Y_c_732_n 0.01056f $X=7.145 $Y=1.185 $X2=0 $Y2=0
cc_306 N_B1_M1028_g N_Y_c_733_n 0.00919683f $X=7.065 $Y=2.465 $X2=0 $Y2=0
cc_307 N_B1_c_310_n N_Y_c_733_n 0.0321355f $X=7.11 $Y=1.17 $X2=0 $Y2=0
cc_308 N_B1_c_311_n N_Y_c_733_n 0.00803689f $X=7.145 $Y=1.35 $X2=0 $Y2=0
cc_309 N_B1_c_313_n N_Y_c_733_n 0.00569489f $X=7.145 $Y=1.185 $X2=0 $Y2=0
cc_310 N_B1_c_306_n N_Y_c_770_n 7.62368e-19 $X=4.905 $Y=1.185 $X2=0 $Y2=0
cc_311 N_B1_c_315_n N_Y_c_770_n 0.0229533f $X=5.18 $Y=1.3 $X2=0 $Y2=0
cc_312 N_B1_c_309_n N_Y_c_772_n 0.0217194f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_313 N_B1_M1028_g N_Y_c_736_n 9.1526e-19 $X=7.065 $Y=2.465 $X2=0 $Y2=0
cc_314 N_B1_c_309_n N_Y_c_774_n 0.0198615f $X=6.98 $Y=1.17 $X2=0 $Y2=0
cc_315 N_B1_c_310_n N_Y_c_774_n 0.00195878f $X=7.11 $Y=1.17 $X2=0 $Y2=0
cc_316 N_B1_c_313_n N_Y_c_774_n 7.1616e-19 $X=7.145 $Y=1.185 $X2=0 $Y2=0
cc_317 N_B1_c_302_n Y 0.00327998f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_318 N_B1_c_312_n Y 0.00240375f $X=4.905 $Y=1.35 $X2=0 $Y2=0
cc_319 N_B1_c_314_n Y 0.0187698f $X=4.895 $Y=1.3 $X2=0 $Y2=0
cc_320 N_B1_c_302_n N_Y_c_738_n 0.00954049f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_321 N_B1_c_314_n N_Y_c_738_n 0.00478478f $X=4.895 $Y=1.3 $X2=0 $Y2=0
cc_322 N_B1_c_304_n N_Y_c_782_n 0.0127252f $X=4.475 $Y=1.185 $X2=0 $Y2=0
cc_323 N_B1_c_314_n N_Y_c_782_n 0.0209479f $X=4.895 $Y=1.3 $X2=0 $Y2=0
cc_324 N_B1_c_306_n N_Y_c_784_n 0.00279843f $X=4.905 $Y=1.185 $X2=0 $Y2=0
cc_325 N_B1_c_312_n N_Y_c_784_n 0.00199064f $X=4.905 $Y=1.35 $X2=0 $Y2=0
cc_326 N_B1_c_302_n N_VGND_c_877_n 0.00453051f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_327 N_B1_c_302_n N_VGND_c_878_n 0.00406904f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_328 N_B1_c_304_n N_VGND_c_878_n 0.00364083f $X=4.475 $Y=1.185 $X2=0 $Y2=0
cc_329 N_B1_c_302_n N_VGND_c_879_n 4.8729e-19 $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_330 N_B1_c_304_n N_VGND_c_879_n 0.00724225f $X=4.475 $Y=1.185 $X2=0 $Y2=0
cc_331 N_B1_c_306_n N_VGND_c_879_n 0.00157435f $X=4.905 $Y=1.185 $X2=0 $Y2=0
cc_332 N_B1_c_306_n N_VGND_c_880_n 0.00426006f $X=4.905 $Y=1.185 $X2=0 $Y2=0
cc_333 N_B1_c_313_n N_VGND_c_884_n 0.00327088f $X=7.145 $Y=1.185 $X2=0 $Y2=0
cc_334 N_B1_c_313_n N_VGND_c_889_n 0.00428252f $X=7.145 $Y=1.185 $X2=0 $Y2=0
cc_335 N_B1_c_302_n N_VGND_c_894_n 0.00610132f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_336 N_B1_c_304_n N_VGND_c_894_n 0.00430165f $X=4.475 $Y=1.185 $X2=0 $Y2=0
cc_337 N_B1_c_306_n N_VGND_c_894_n 0.00583081f $X=4.905 $Y=1.185 $X2=0 $Y2=0
cc_338 N_B1_c_313_n N_VGND_c_894_n 0.00691896f $X=7.145 $Y=1.185 $X2=0 $Y2=0
cc_339 N_C1_c_430_n N_A_45_367#_c_516_n 0.00216323f $X=5.975 $Y=1.595 $X2=0
+ $Y2=0
cc_340 N_C1_M1010_g N_A_45_367#_c_550_n 0.0166995f $X=5.345 $Y=2.465 $X2=0 $Y2=0
cc_341 N_C1_M1013_g N_A_45_367#_c_550_n 0.0136548f $X=5.775 $Y=2.465 $X2=0 $Y2=0
cc_342 N_C1_M1021_g N_A_45_367#_c_550_n 0.0136547f $X=6.205 $Y=2.465 $X2=0 $Y2=0
cc_343 N_C1_M1030_g N_A_45_367#_c_550_n 0.0141382f $X=6.635 $Y=2.465 $X2=0 $Y2=0
cc_344 N_C1_c_430_n N_A_45_367#_c_550_n 0.00124371f $X=5.975 $Y=1.595 $X2=0
+ $Y2=0
cc_345 N_C1_M1030_g N_A_45_367#_c_517_n 7.53175e-19 $X=6.635 $Y=2.465 $X2=0
+ $Y2=0
cc_346 N_C1_M1030_g N_A_45_367#_c_518_n 7.36266e-19 $X=6.635 $Y=2.465 $X2=0
+ $Y2=0
cc_347 N_C1_M1010_g N_VPWR_c_617_n 0.00357877f $X=5.345 $Y=2.465 $X2=0 $Y2=0
cc_348 N_C1_M1013_g N_VPWR_c_617_n 0.00357877f $X=5.775 $Y=2.465 $X2=0 $Y2=0
cc_349 N_C1_M1021_g N_VPWR_c_617_n 0.00357877f $X=6.205 $Y=2.465 $X2=0 $Y2=0
cc_350 N_C1_M1030_g N_VPWR_c_617_n 0.00357877f $X=6.635 $Y=2.465 $X2=0 $Y2=0
cc_351 N_C1_M1010_g N_VPWR_c_606_n 0.00537654f $X=5.345 $Y=2.465 $X2=0 $Y2=0
cc_352 N_C1_M1013_g N_VPWR_c_606_n 0.0053512f $X=5.775 $Y=2.465 $X2=0 $Y2=0
cc_353 N_C1_M1021_g N_VPWR_c_606_n 0.0053512f $X=6.205 $Y=2.465 $X2=0 $Y2=0
cc_354 N_C1_M1030_g N_VPWR_c_606_n 0.00537654f $X=6.635 $Y=2.465 $X2=0 $Y2=0
cc_355 N_C1_M1010_g N_A_826_367#_c_706_n 0.0119021f $X=5.345 $Y=2.465 $X2=0
+ $Y2=0
cc_356 N_C1_M1013_g N_A_826_367#_c_706_n 0.0119021f $X=5.775 $Y=2.465 $X2=0
+ $Y2=0
cc_357 N_C1_M1021_g N_A_826_367#_c_706_n 0.0118112f $X=6.205 $Y=2.465 $X2=0
+ $Y2=0
cc_358 N_C1_M1030_g N_A_826_367#_c_706_n 0.0119021f $X=6.635 $Y=2.465 $X2=0
+ $Y2=0
cc_359 N_C1_M1000_g N_Y_c_753_n 0.00638313f $X=5.335 $Y=0.655 $X2=0 $Y2=0
cc_360 N_C1_M1001_g N_Y_c_753_n 4.66504e-19 $X=5.765 $Y=0.655 $X2=0 $Y2=0
cc_361 N_C1_M1000_g N_Y_c_755_n 0.00886808f $X=5.335 $Y=0.655 $X2=0 $Y2=0
cc_362 N_C1_M1001_g N_Y_c_755_n 0.00886808f $X=5.765 $Y=0.655 $X2=0 $Y2=0
cc_363 N_C1_M1010_g N_Y_c_756_n 0.0045107f $X=5.345 $Y=2.465 $X2=0 $Y2=0
cc_364 N_C1_M1013_g N_Y_c_756_n 0.00952341f $X=5.775 $Y=2.465 $X2=0 $Y2=0
cc_365 N_C1_M1021_g N_Y_c_756_n 0.0102006f $X=6.205 $Y=2.465 $X2=0 $Y2=0
cc_366 N_C1_c_423_n N_Y_c_756_n 0.00694943f $X=6.535 $Y=1.51 $X2=0 $Y2=0
cc_367 N_C1_c_424_n N_Y_c_756_n 0.0011477f $X=6.635 $Y=1.51 $X2=0 $Y2=0
cc_368 N_C1_c_430_n N_Y_c_756_n 0.0495681f $X=5.975 $Y=1.595 $X2=0 $Y2=0
cc_369 N_C1_M1000_g N_Y_c_796_n 5.25357e-19 $X=5.335 $Y=0.655 $X2=0 $Y2=0
cc_370 N_C1_M1001_g N_Y_c_796_n 0.00674009f $X=5.765 $Y=0.655 $X2=0 $Y2=0
cc_371 N_C1_M1014_g N_Y_c_796_n 0.00674041f $X=6.195 $Y=0.655 $X2=0 $Y2=0
cc_372 N_C1_M1022_g N_Y_c_796_n 5.68592e-19 $X=6.625 $Y=0.655 $X2=0 $Y2=0
cc_373 N_C1_M1014_g N_Y_c_757_n 0.00886808f $X=6.195 $Y=0.655 $X2=0 $Y2=0
cc_374 N_C1_M1022_g N_Y_c_757_n 0.00886808f $X=6.625 $Y=0.655 $X2=0 $Y2=0
cc_375 N_C1_M1030_g N_Y_c_734_n 0.00750487f $X=6.635 $Y=2.465 $X2=0 $Y2=0
cc_376 N_C1_c_423_n N_Y_c_734_n 0.00656934f $X=6.535 $Y=1.51 $X2=0 $Y2=0
cc_377 N_C1_M1014_g N_Y_c_762_n 5.68592e-19 $X=6.195 $Y=0.655 $X2=0 $Y2=0
cc_378 N_C1_M1022_g N_Y_c_762_n 0.00673209f $X=6.625 $Y=0.655 $X2=0 $Y2=0
cc_379 N_C1_M1000_g N_Y_c_770_n 0.00106715f $X=5.335 $Y=0.655 $X2=0 $Y2=0
cc_380 N_C1_M1001_g N_Y_c_772_n 7.17169e-19 $X=5.765 $Y=0.655 $X2=0 $Y2=0
cc_381 N_C1_M1014_g N_Y_c_772_n 7.17169e-19 $X=6.195 $Y=0.655 $X2=0 $Y2=0
cc_382 N_C1_M1021_g N_Y_c_736_n 5.2288e-19 $X=6.205 $Y=2.465 $X2=0 $Y2=0
cc_383 N_C1_M1030_g N_Y_c_736_n 0.00633007f $X=6.635 $Y=2.465 $X2=0 $Y2=0
cc_384 N_C1_c_423_n N_Y_c_736_n 0.0228039f $X=6.535 $Y=1.51 $X2=0 $Y2=0
cc_385 N_C1_c_424_n N_Y_c_736_n 0.00240338f $X=6.635 $Y=1.51 $X2=0 $Y2=0
cc_386 N_C1_M1022_g N_Y_c_774_n 7.17169e-19 $X=6.625 $Y=0.655 $X2=0 $Y2=0
cc_387 N_C1_M1000_g N_VGND_c_880_n 0.00428252f $X=5.335 $Y=0.655 $X2=0 $Y2=0
cc_388 N_C1_M1000_g N_VGND_c_881_n 0.00153274f $X=5.335 $Y=0.655 $X2=0 $Y2=0
cc_389 N_C1_M1001_g N_VGND_c_881_n 0.00153274f $X=5.765 $Y=0.655 $X2=0 $Y2=0
cc_390 N_C1_M1014_g N_VGND_c_882_n 0.00153274f $X=6.195 $Y=0.655 $X2=0 $Y2=0
cc_391 N_C1_M1022_g N_VGND_c_882_n 0.00153274f $X=6.625 $Y=0.655 $X2=0 $Y2=0
cc_392 N_C1_M1001_g N_VGND_c_885_n 0.00428252f $X=5.765 $Y=0.655 $X2=0 $Y2=0
cc_393 N_C1_M1014_g N_VGND_c_885_n 0.00428252f $X=6.195 $Y=0.655 $X2=0 $Y2=0
cc_394 N_C1_M1022_g N_VGND_c_889_n 0.00428252f $X=6.625 $Y=0.655 $X2=0 $Y2=0
cc_395 N_C1_M1000_g N_VGND_c_894_n 0.00587209f $X=5.335 $Y=0.655 $X2=0 $Y2=0
cc_396 N_C1_M1001_g N_VGND_c_894_n 0.00584676f $X=5.765 $Y=0.655 $X2=0 $Y2=0
cc_397 N_C1_M1014_g N_VGND_c_894_n 0.00584676f $X=6.195 $Y=0.655 $X2=0 $Y2=0
cc_398 N_C1_M1022_g N_VGND_c_894_n 0.00587209f $X=6.625 $Y=0.655 $X2=0 $Y2=0
cc_399 N_A_45_367#_c_521_n N_VPWR_M1004_d 0.00332334f $X=1.115 $Y=2.04 $X2=-0.19
+ $Y2=1.655
cc_400 N_A_45_367#_c_525_n N_VPWR_M1012_d 0.00352229f $X=1.975 $Y=2.04 $X2=0
+ $Y2=0
cc_401 N_A_45_367#_c_527_n N_VPWR_M1016_s 0.00339614f $X=2.835 $Y=2.04 $X2=0
+ $Y2=0
cc_402 N_A_45_367#_c_528_n N_VPWR_M1027_s 0.00448943f $X=3.695 $Y=2.04 $X2=0
+ $Y2=0
cc_403 N_A_45_367#_c_521_n N_VPWR_c_607_n 0.0170777f $X=1.115 $Y=2.04 $X2=0
+ $Y2=0
cc_404 N_A_45_367#_c_525_n N_VPWR_c_608_n 0.0170777f $X=1.975 $Y=2.04 $X2=0
+ $Y2=0
cc_405 N_A_45_367#_c_527_n N_VPWR_c_609_n 0.0170777f $X=2.835 $Y=2.04 $X2=0
+ $Y2=0
cc_406 N_A_45_367#_c_528_n N_VPWR_c_610_n 0.0193595f $X=3.695 $Y=2.04 $X2=0
+ $Y2=0
cc_407 N_A_45_367#_c_570_p N_VPWR_c_611_n 0.0124525f $X=2.07 $Y=2.91 $X2=0 $Y2=0
cc_408 N_A_45_367#_c_571_p N_VPWR_c_613_n 0.0124525f $X=2.93 $Y=2.9 $X2=0 $Y2=0
cc_409 N_A_45_367#_c_514_n N_VPWR_c_615_n 0.0178111f $X=0.35 $Y=2.91 $X2=0 $Y2=0
cc_410 N_A_45_367#_c_573_p N_VPWR_c_616_n 0.0124525f $X=1.21 $Y=2.91 $X2=0 $Y2=0
cc_411 N_A_45_367#_c_535_n N_VPWR_c_617_n 0.0146794f $X=3.84 $Y=2.45 $X2=0 $Y2=0
cc_412 N_A_45_367#_c_550_n N_VPWR_c_617_n 0.00203954f $X=7.135 $Y=2.45 $X2=0
+ $Y2=0
cc_413 N_A_45_367#_c_518_n N_VPWR_c_617_n 0.0187054f $X=7.3 $Y=2.95 $X2=0 $Y2=0
cc_414 N_A_45_367#_M1004_s N_VPWR_c_606_n 0.00371702f $X=0.225 $Y=1.835 $X2=0
+ $Y2=0
cc_415 N_A_45_367#_M1009_s N_VPWR_c_606_n 0.00536646f $X=1.07 $Y=1.835 $X2=0
+ $Y2=0
cc_416 N_A_45_367#_M1005_d N_VPWR_c_606_n 0.00536646f $X=1.93 $Y=1.835 $X2=0
+ $Y2=0
cc_417 N_A_45_367#_M1025_d N_VPWR_c_606_n 0.00536646f $X=2.79 $Y=1.835 $X2=0
+ $Y2=0
cc_418 N_A_45_367#_M1018_s N_VPWR_c_606_n 0.00345315f $X=3.7 $Y=1.835 $X2=0
+ $Y2=0
cc_419 N_A_45_367#_M1017_d N_VPWR_c_606_n 0.00225186f $X=4.56 $Y=1.835 $X2=0
+ $Y2=0
cc_420 N_A_45_367#_M1028_d N_VPWR_c_606_n 0.00232623f $X=7.14 $Y=1.835 $X2=0
+ $Y2=0
cc_421 N_A_45_367#_c_514_n N_VPWR_c_606_n 0.0100304f $X=0.35 $Y=2.91 $X2=0 $Y2=0
cc_422 N_A_45_367#_c_573_p N_VPWR_c_606_n 0.00730901f $X=1.21 $Y=2.91 $X2=0
+ $Y2=0
cc_423 N_A_45_367#_c_570_p N_VPWR_c_606_n 0.00730901f $X=2.07 $Y=2.91 $X2=0
+ $Y2=0
cc_424 N_A_45_367#_c_571_p N_VPWR_c_606_n 0.00730901f $X=2.93 $Y=2.9 $X2=0 $Y2=0
cc_425 N_A_45_367#_c_535_n N_VPWR_c_606_n 0.00955018f $X=3.84 $Y=2.45 $X2=0
+ $Y2=0
cc_426 N_A_45_367#_c_550_n N_VPWR_c_606_n 0.0072215f $X=7.135 $Y=2.45 $X2=0
+ $Y2=0
cc_427 N_A_45_367#_c_518_n N_VPWR_c_606_n 0.012538f $X=7.3 $Y=2.95 $X2=0 $Y2=0
cc_428 N_A_45_367#_c_516_n N_A_826_367#_M1007_s 0.00176461f $X=4.595 $Y=1.79
+ $X2=-0.19 $Y2=1.655
cc_429 N_A_45_367#_c_550_n N_A_826_367#_M1019_s 0.008388f $X=7.135 $Y=2.45 $X2=0
+ $Y2=0
cc_430 N_A_45_367#_c_550_n N_A_826_367#_M1013_d 0.00350157f $X=7.135 $Y=2.45
+ $X2=0 $Y2=0
cc_431 N_A_45_367#_c_550_n N_A_826_367#_M1030_d 0.00423004f $X=7.135 $Y=2.45
+ $X2=0 $Y2=0
cc_432 N_A_45_367#_c_516_n N_A_826_367#_c_716_n 0.0135055f $X=4.595 $Y=1.79
+ $X2=0 $Y2=0
cc_433 N_A_45_367#_M1017_d N_A_826_367#_c_706_n 0.00339199f $X=4.56 $Y=1.835
+ $X2=0 $Y2=0
cc_434 N_A_45_367#_c_550_n N_A_826_367#_c_706_n 0.116126f $X=7.135 $Y=2.45 $X2=0
+ $Y2=0
cc_435 N_A_45_367#_c_598_p N_A_826_367#_c_706_n 0.0136347f $X=4.805 $Y=2.45
+ $X2=0 $Y2=0
cc_436 N_A_45_367#_c_550_n N_Y_M1010_s 0.00350157f $X=7.135 $Y=2.45 $X2=0 $Y2=0
cc_437 N_A_45_367#_c_550_n N_Y_M1021_s 0.00349756f $X=7.135 $Y=2.45 $X2=0 $Y2=0
cc_438 N_A_45_367#_c_550_n N_Y_c_756_n 0.0461014f $X=7.135 $Y=2.45 $X2=0 $Y2=0
cc_439 N_A_45_367#_M1028_d N_Y_c_734_n 0.00333692f $X=7.14 $Y=1.835 $X2=0 $Y2=0
cc_440 N_A_45_367#_c_550_n N_Y_c_734_n 0.0170575f $X=7.135 $Y=2.45 $X2=0 $Y2=0
cc_441 N_A_45_367#_c_517_n N_Y_c_734_n 0.0217862f $X=7.3 $Y=2.575 $X2=0 $Y2=0
cc_442 N_A_45_367#_c_550_n N_Y_c_736_n 0.0163324f $X=7.135 $Y=2.45 $X2=0 $Y2=0
cc_443 N_VPWR_c_606_n N_A_826_367#_M1007_s 0.00341839f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_444 N_VPWR_c_606_n N_A_826_367#_M1019_s 0.00223577f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_606_n N_A_826_367#_M1013_d 0.00223577f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_606_n N_A_826_367#_M1030_d 0.00236437f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_617_n N_A_826_367#_c_724_n 0.0132331f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_606_n N_A_826_367#_c_724_n 0.00816431f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_617_n N_A_826_367#_c_706_n 0.148245f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_450 N_VPWR_c_606_n N_A_826_367#_c_706_n 0.0942853f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_606_n N_Y_M1010_s 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_452 N_VPWR_c_606_n N_Y_M1021_s 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_453 N_A_826_367#_c_706_n N_Y_M1010_s 0.00339639f $X=6.85 $Y=2.91 $X2=0 $Y2=0
cc_454 N_A_826_367#_c_706_n N_Y_M1021_s 0.00339639f $X=6.85 $Y=2.91 $X2=4.475
+ $Y2=1.185
cc_455 N_A_826_367#_M1013_d N_Y_c_756_n 0.00340276f $X=5.85 $Y=1.835 $X2=3.995
+ $Y2=1.21
cc_456 N_A_826_367#_M1030_d N_Y_c_734_n 0.00244731f $X=6.71 $Y=1.835 $X2=4.145
+ $Y2=1.35
cc_457 N_Y_c_738_n N_VGND_M1026_d 0.0109946f $X=4.055 $Y=0.882 $X2=0 $Y2=0
cc_458 N_Y_c_749_n N_VGND_M1020_d 0.00109633f $X=4.955 $Y=0.82 $X2=0 $Y2=0
cc_459 N_Y_c_784_n N_VGND_M1020_d 0.00363871f $X=4.725 $Y=0.867 $X2=0 $Y2=0
cc_460 N_Y_c_755_n N_VGND_M1000_d 0.00335318f $X=5.815 $Y=0.83 $X2=0 $Y2=0
cc_461 N_Y_c_757_n N_VGND_M1014_d 0.00335318f $X=6.675 $Y=0.83 $X2=0 $Y2=0
cc_462 N_Y_c_732_n N_VGND_M1031_d 0.00753544f $X=7.41 $Y=0.83 $X2=0 $Y2=0
cc_463 N_Y_c_737_n N_VGND_c_877_n 0.0254367f $X=4.26 $Y=0.42 $X2=0 $Y2=0
cc_464 N_Y_c_738_n N_VGND_c_877_n 0.02177f $X=4.055 $Y=0.882 $X2=0 $Y2=0
cc_465 N_Y_c_737_n N_VGND_c_878_n 0.0184149f $X=4.26 $Y=0.42 $X2=0 $Y2=0
cc_466 N_Y_c_738_n N_VGND_c_878_n 0.00188421f $X=4.055 $Y=0.882 $X2=0 $Y2=0
cc_467 N_Y_c_782_n N_VGND_c_878_n 0.00206327f $X=4.583 $Y=0.867 $X2=0 $Y2=0
cc_468 N_Y_c_782_n N_VGND_c_879_n 0.0150767f $X=4.583 $Y=0.867 $X2=0 $Y2=0
cc_469 N_Y_c_749_n N_VGND_c_880_n 0.00201785f $X=4.955 $Y=0.82 $X2=0 $Y2=0
cc_470 N_Y_c_753_n N_VGND_c_880_n 0.0188913f $X=5.12 $Y=0.37 $X2=0 $Y2=0
cc_471 N_Y_c_755_n N_VGND_c_880_n 0.00191958f $X=5.815 $Y=0.83 $X2=0 $Y2=0
cc_472 N_Y_c_755_n N_VGND_c_881_n 0.0130506f $X=5.815 $Y=0.83 $X2=0 $Y2=0
cc_473 N_Y_c_757_n N_VGND_c_882_n 0.0130506f $X=6.675 $Y=0.83 $X2=0 $Y2=0
cc_474 N_Y_c_732_n N_VGND_c_883_n 0.00237918f $X=7.41 $Y=0.83 $X2=0 $Y2=0
cc_475 N_Y_c_732_n N_VGND_c_884_n 0.0197079f $X=7.41 $Y=0.83 $X2=0 $Y2=0
cc_476 N_Y_c_755_n N_VGND_c_885_n 0.00191958f $X=5.815 $Y=0.83 $X2=0 $Y2=0
cc_477 N_Y_c_796_n N_VGND_c_885_n 0.0188913f $X=5.98 $Y=0.37 $X2=0 $Y2=0
cc_478 N_Y_c_757_n N_VGND_c_885_n 0.00191958f $X=6.675 $Y=0.83 $X2=0 $Y2=0
cc_479 N_Y_c_738_n N_VGND_c_888_n 0.00192662f $X=4.055 $Y=0.882 $X2=0 $Y2=0
cc_480 N_Y_c_757_n N_VGND_c_889_n 0.00191958f $X=6.675 $Y=0.83 $X2=0 $Y2=0
cc_481 N_Y_c_762_n N_VGND_c_889_n 0.0188913f $X=6.84 $Y=0.37 $X2=0 $Y2=0
cc_482 N_Y_c_732_n N_VGND_c_889_n 0.00191958f $X=7.41 $Y=0.83 $X2=0 $Y2=0
cc_483 N_Y_M1002_d N_VGND_c_894_n 0.00225186f $X=1.86 $Y=0.235 $X2=0 $Y2=0
cc_484 N_Y_M1015_d N_VGND_c_894_n 0.00225186f $X=2.72 $Y=0.235 $X2=0 $Y2=0
cc_485 N_Y_M1011_s N_VGND_c_894_n 0.00244361f $X=4.12 $Y=0.235 $X2=0 $Y2=0
cc_486 N_Y_M1029_s N_VGND_c_894_n 0.00223559f $X=4.98 $Y=0.235 $X2=0 $Y2=0
cc_487 N_Y_M1001_s N_VGND_c_894_n 0.00223559f $X=5.84 $Y=0.235 $X2=0 $Y2=0
cc_488 N_Y_M1022_s N_VGND_c_894_n 0.00223559f $X=6.7 $Y=0.235 $X2=0 $Y2=0
cc_489 N_Y_c_737_n N_VGND_c_894_n 0.0112195f $X=4.26 $Y=0.42 $X2=0 $Y2=0
cc_490 N_Y_c_749_n N_VGND_c_894_n 0.00387795f $X=4.955 $Y=0.82 $X2=0 $Y2=0
cc_491 N_Y_c_753_n N_VGND_c_894_n 0.012376f $X=5.12 $Y=0.37 $X2=0 $Y2=0
cc_492 N_Y_c_755_n N_VGND_c_894_n 0.00827851f $X=5.815 $Y=0.83 $X2=0 $Y2=0
cc_493 N_Y_c_796_n N_VGND_c_894_n 0.012376f $X=5.98 $Y=0.37 $X2=0 $Y2=0
cc_494 N_Y_c_757_n N_VGND_c_894_n 0.00827851f $X=6.675 $Y=0.83 $X2=0 $Y2=0
cc_495 N_Y_c_762_n N_VGND_c_894_n 0.012376f $X=6.84 $Y=0.37 $X2=0 $Y2=0
cc_496 N_Y_c_732_n N_VGND_c_894_n 0.00885552f $X=7.41 $Y=0.83 $X2=0 $Y2=0
cc_497 N_Y_c_738_n N_VGND_c_894_n 0.0117371f $X=4.055 $Y=0.882 $X2=0 $Y2=0
cc_498 N_Y_c_782_n N_VGND_c_894_n 0.00498915f $X=4.583 $Y=0.867 $X2=0 $Y2=0
cc_499 N_Y_c_738_n N_A_114_47#_M1003_s 0.00331384f $X=4.055 $Y=0.882 $X2=0 $Y2=0
cc_500 N_Y_c_738_n N_A_114_47#_M1024_s 0.0058129f $X=4.055 $Y=0.882 $X2=0 $Y2=0
cc_501 N_Y_M1002_d N_A_114_47#_c_1011_n 0.00330327f $X=1.86 $Y=0.235 $X2=0 $Y2=0
cc_502 N_Y_M1015_d N_A_114_47#_c_1011_n 0.00330327f $X=2.72 $Y=0.235 $X2=0 $Y2=0
cc_503 N_Y_c_738_n N_A_114_47#_c_1011_n 0.0840442f $X=4.055 $Y=0.882 $X2=0 $Y2=0
cc_504 N_VGND_c_894_n N_A_114_47#_M1006_s 0.00432284f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_505 N_VGND_c_894_n N_A_114_47#_M1023_s 0.00376627f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_506 N_VGND_c_894_n N_A_114_47#_M1003_s 0.00223577f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_507 N_VGND_c_894_n N_A_114_47#_M1024_s 0.00247154f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_508 N_VGND_c_887_n N_A_114_47#_c_1024_n 0.0135169f $X=0.975 $Y=0 $X2=0 $Y2=0
cc_509 N_VGND_c_894_n N_A_114_47#_c_1024_n 0.00847534f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_510 N_VGND_M1008_d N_A_114_47#_c_1000_n 0.00176461f $X=1 $Y=0.235 $X2=0 $Y2=0
cc_511 N_VGND_c_876_n N_A_114_47#_c_1000_n 0.0170777f $X=1.14 $Y=0.38 $X2=0
+ $Y2=0
cc_512 N_VGND_c_875_n N_A_114_47#_c_1001_n 0.00166817f $X=0.28 $Y=0.38 $X2=0
+ $Y2=0
cc_513 N_VGND_c_888_n N_A_114_47#_c_1029_n 0.0125234f $X=3.555 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_894_n N_A_114_47#_c_1029_n 0.00738676f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_515 N_VGND_c_888_n N_A_114_47#_c_1011_n 0.0985947f $X=3.555 $Y=0 $X2=0 $Y2=0
cc_516 N_VGND_c_894_n N_A_114_47#_c_1011_n 0.062601f $X=7.44 $Y=0 $X2=0 $Y2=0
