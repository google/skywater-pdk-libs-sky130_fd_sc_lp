* File: sky130_fd_sc_lp__a22o_2.pxi.spice
* Created: Fri Aug 28 09:54:07 2020
* 
x_PM_SKY130_FD_SC_LP__A22O_2%A_94_249# N_A_94_249#_M1000_d N_A_94_249#_M1007_d
+ N_A_94_249#_M1010_s N_A_94_249#_M1004_d N_A_94_249#_M1008_g
+ N_A_94_249#_M1001_g N_A_94_249#_M1011_g N_A_94_249#_M1002_g N_A_94_249#_c_72_n
+ N_A_94_249#_c_73_n N_A_94_249#_c_74_n N_A_94_249#_c_75_n N_A_94_249#_c_76_n
+ N_A_94_249#_c_77_n N_A_94_249#_c_111_p N_A_94_249#_c_83_n N_A_94_249#_c_78_n
+ N_A_94_249#_c_84_n N_A_94_249#_c_85_n N_A_94_249#_c_79_n
+ PM_SKY130_FD_SC_LP__A22O_2%A_94_249#
x_PM_SKY130_FD_SC_LP__A22O_2%A2 N_A2_M1009_g N_A2_M1005_g A2 N_A2_c_185_n
+ N_A2_c_186_n PM_SKY130_FD_SC_LP__A22O_2%A2
x_PM_SKY130_FD_SC_LP__A22O_2%A1 N_A1_M1000_g N_A1_M1003_g A1 A1 N_A1_c_225_n
+ N_A1_c_226_n PM_SKY130_FD_SC_LP__A22O_2%A1
x_PM_SKY130_FD_SC_LP__A22O_2%B2 N_B2_M1010_g N_B2_M1006_g B2 N_B2_c_261_n
+ PM_SKY130_FD_SC_LP__A22O_2%B2
x_PM_SKY130_FD_SC_LP__A22O_2%B1 N_B1_M1007_g N_B1_M1004_g B1 N_B1_c_294_n
+ N_B1_c_295_n PM_SKY130_FD_SC_LP__A22O_2%B1
x_PM_SKY130_FD_SC_LP__A22O_2%VPWR N_VPWR_M1008_s N_VPWR_M1011_s N_VPWR_M1003_d
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n VPWR
+ N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_319_n N_VPWR_c_328_n
+ N_VPWR_c_329_n PM_SKY130_FD_SC_LP__A22O_2%VPWR
x_PM_SKY130_FD_SC_LP__A22O_2%X N_X_M1001_d N_X_M1008_d N_X_c_373_n N_X_c_370_n
+ N_X_c_372_n X X N_X_c_385_n X PM_SKY130_FD_SC_LP__A22O_2%X
x_PM_SKY130_FD_SC_LP__A22O_2%A_326_367# N_A_326_367#_M1009_d
+ N_A_326_367#_M1010_d N_A_326_367#_c_402_n N_A_326_367#_c_405_n
+ N_A_326_367#_c_397_n N_A_326_367#_c_411_n N_A_326_367#_c_406_n
+ PM_SKY130_FD_SC_LP__A22O_2%A_326_367#
x_PM_SKY130_FD_SC_LP__A22O_2%VGND N_VGND_M1001_s N_VGND_M1002_s N_VGND_M1006_s
+ N_VGND_c_425_n N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n
+ VGND N_VGND_c_430_n N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n
+ N_VGND_c_434_n PM_SKY130_FD_SC_LP__A22O_2%VGND
cc_1 VNB N_A_94_249#_M1008_g 0.0191811f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_2 VNB N_A_94_249#_M1001_g 0.0249119f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.665
cc_3 VNB N_A_94_249#_M1011_g 0.00419036f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_4 VNB N_A_94_249#_M1002_g 0.0195466f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=0.665
cc_5 VNB N_A_94_249#_c_72_n 0.00714787f $X=-0.19 $Y=-0.245 $X2=2.035 $Y2=1.08
cc_6 VNB N_A_94_249#_c_73_n 0.00748998f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.08
cc_7 VNB N_A_94_249#_c_74_n 0.00854602f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=0.42
cc_8 VNB N_A_94_249#_c_75_n 0.0110752f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.93
cc_9 VNB N_A_94_249#_c_76_n 0.0177756f $X=-0.19 $Y=-0.245 $X2=3.385 $Y2=1.08
cc_10 VNB N_A_94_249#_c_77_n 0.0170393f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=1.08
cc_11 VNB N_A_94_249#_c_78_n 0.0288914f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=0.42
cc_12 VNB N_A_94_249#_c_79_n 0.0504198f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.41
cc_13 VNB N_A2_M1005_g 0.0244635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_185_n 0.024295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_186_n 0.00450243f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.395
cc_16 VNB N_A1_M1000_g 0.0277014f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=1.835
cc_17 VNB N_A1_c_225_n 0.033248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_226_n 0.0017619f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.245
cc_19 VNB N_B2_M1006_g 0.0264832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B2 0.00344711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B2_c_261_n 0.0259318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_M1007_g 0.0275273f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=1.835
cc_23 VNB N_B1_M1004_g 0.00179535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_c_294_n 0.0485726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_c_295_n 0.0116455f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_26 VNB N_VPWR_c_319_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=0.42
cc_27 VNB N_X_c_370_n 0.00283128f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_28 VNB N_VGND_c_425_n 0.0115378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_426_n 0.049327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_427_n 0.021138f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_31 VNB N_VGND_c_428_n 0.00599595f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.665
cc_32 VNB N_VGND_c_429_n 0.00852114f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_33 VNB N_VGND_c_430_n 0.03125f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=0.665
cc_34 VNB N_VGND_c_431_n 0.0270663f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=0.42
cc_35 VNB N_VGND_c_432_n 0.2205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_433_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=2.035
cc_37 VNB N_VGND_c_434_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=0.995
cc_38 VPB N_A_94_249#_M1008_g 0.0270105f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_39 VPB N_A_94_249#_M1011_g 0.0213298f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_40 VPB N_A_94_249#_c_75_n 0.00495342f $X=-0.19 $Y=1.655 $X2=2.535 $Y2=1.93
cc_41 VPB N_A_94_249#_c_83_n 0.00401936f $X=-0.19 $Y=1.655 $X2=2.62 $Y2=2.035
cc_42 VPB N_A_94_249#_c_84_n 0.00920755f $X=-0.19 $Y=1.655 $X2=3.615 $Y2=2.14
cc_43 VPB N_A_94_249#_c_85_n 0.0354376f $X=-0.19 $Y=1.655 $X2=3.58 $Y2=2.475
cc_44 VPB N_A2_M1009_g 0.0200159f $X=-0.19 $Y=1.655 $X2=2.595 $Y2=1.835
cc_45 VPB N_A2_c_185_n 0.00677079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A2_c_186_n 0.00500967f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.395
cc_47 VPB N_A1_M1003_g 0.0225735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A1_c_225_n 0.00964859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A1_c_226_n 0.00128511f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.245
cc_50 VPB N_B2_M1010_g 0.0226133f $X=-0.19 $Y=1.655 $X2=2.595 $Y2=1.835
cc_51 VPB B2 0.00377335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_B2_c_261_n 0.0063256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_B1_M1004_g 0.0263397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B1_c_295_n 0.00645499f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_55 VPB N_VPWR_c_320_n 0.012247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_321_n 0.0475609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_322_n 0.00495383f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=0.665
cc_58 VPB N_VPWR_c_323_n 0.00908224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_324_n 0.0184717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_325_n 0.0155889f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=0.42
cc_61 VPB N_VPWR_c_326_n 0.0433388f $X=-0.19 $Y=1.655 $X2=3.55 $Y2=0.995
cc_62 VPB N_VPWR_c_319_n 0.0503575f $X=-0.19 $Y=1.655 $X2=3.55 $Y2=0.42
cc_63 VPB N_VPWR_c_328_n 0.00631677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_329_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=1.41
cc_65 VPB N_X_c_370_n 4.76728e-19 $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_66 VPB N_X_c_372_n 0.00200272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_326_367#_c_397_n 0.0116489f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_68 N_A_94_249#_M1011_g N_A2_M1009_g 0.0323512f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_69 N_A_94_249#_M1002_g N_A2_M1005_g 0.0260771f $X=1.05 $Y=0.665 $X2=0 $Y2=0
cc_70 N_A_94_249#_c_72_n N_A2_M1005_g 0.015296f $X=2.035 $Y=1.08 $X2=0 $Y2=0
cc_71 N_A_94_249#_c_73_n N_A2_M1005_g 0.00380458f $X=1.28 $Y=1.08 $X2=0 $Y2=0
cc_72 N_A_94_249#_c_74_n N_A2_M1005_g 0.00246041f $X=2.2 $Y=0.42 $X2=0 $Y2=0
cc_73 N_A_94_249#_c_79_n N_A2_M1005_g 0.00262218f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_94_249#_M1011_g N_A2_c_185_n 0.0037549f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_75 N_A_94_249#_c_72_n N_A2_c_185_n 0.00369309f $X=2.035 $Y=1.08 $X2=0 $Y2=0
cc_76 N_A_94_249#_c_73_n N_A2_c_185_n 0.00162646f $X=1.28 $Y=1.08 $X2=0 $Y2=0
cc_77 N_A_94_249#_c_79_n N_A2_c_185_n 0.0142478f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_94_249#_M1011_g N_A2_c_186_n 0.0019789f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A_94_249#_c_72_n N_A2_c_186_n 0.0320324f $X=2.035 $Y=1.08 $X2=0 $Y2=0
cc_80 N_A_94_249#_c_73_n N_A2_c_186_n 0.0196499f $X=1.28 $Y=1.08 $X2=0 $Y2=0
cc_81 N_A_94_249#_c_72_n N_A1_M1000_g 0.0144354f $X=2.035 $Y=1.08 $X2=0 $Y2=0
cc_82 N_A_94_249#_c_74_n N_A1_M1000_g 0.0155222f $X=2.2 $Y=0.42 $X2=0 $Y2=0
cc_83 N_A_94_249#_c_75_n N_A1_M1000_g 0.00486772f $X=2.535 $Y=1.93 $X2=0 $Y2=0
cc_84 N_A_94_249#_c_77_n N_A1_M1000_g 0.00326747f $X=2.62 $Y=1.08 $X2=0 $Y2=0
cc_85 N_A_94_249#_c_75_n N_A1_M1003_g 0.00116202f $X=2.535 $Y=1.93 $X2=0 $Y2=0
cc_86 N_A_94_249#_c_83_n N_A1_M1003_g 0.00110295f $X=2.62 $Y=2.035 $X2=0 $Y2=0
cc_87 N_A_94_249#_c_75_n N_A1_c_225_n 0.00298958f $X=2.535 $Y=1.93 $X2=0 $Y2=0
cc_88 N_A_94_249#_c_77_n N_A1_c_225_n 0.00429125f $X=2.62 $Y=1.08 $X2=0 $Y2=0
cc_89 N_A_94_249#_c_75_n N_A1_c_226_n 0.0374933f $X=2.535 $Y=1.93 $X2=0 $Y2=0
cc_90 N_A_94_249#_c_77_n N_A1_c_226_n 0.0143698f $X=2.62 $Y=1.08 $X2=0 $Y2=0
cc_91 N_A_94_249#_c_83_n N_A1_c_226_n 0.0153595f $X=2.62 $Y=2.035 $X2=0 $Y2=0
cc_92 N_A_94_249#_c_75_n N_B2_M1010_g 0.00475552f $X=2.535 $Y=1.93 $X2=0 $Y2=0
cc_93 N_A_94_249#_c_111_p N_B2_M1010_g 0.00952237f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A_94_249#_c_74_n N_B2_M1006_g 0.00303731f $X=2.2 $Y=0.42 $X2=0 $Y2=0
cc_95 N_A_94_249#_c_75_n N_B2_M1006_g 0.00546311f $X=2.535 $Y=1.93 $X2=0 $Y2=0
cc_96 N_A_94_249#_c_76_n N_B2_M1006_g 0.0159399f $X=3.385 $Y=1.08 $X2=0 $Y2=0
cc_97 N_A_94_249#_c_78_n N_B2_M1006_g 0.00240096f $X=3.55 $Y=0.42 $X2=0 $Y2=0
cc_98 N_A_94_249#_c_75_n B2 0.0312891f $X=2.535 $Y=1.93 $X2=0 $Y2=0
cc_99 N_A_94_249#_c_76_n B2 0.0304463f $X=3.385 $Y=1.08 $X2=0 $Y2=0
cc_100 N_A_94_249#_c_111_p B2 0.0268858f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_101 N_A_94_249#_c_75_n N_B2_c_261_n 0.00288855f $X=2.535 $Y=1.93 $X2=0 $Y2=0
cc_102 N_A_94_249#_c_76_n N_B2_c_261_n 0.00520773f $X=3.385 $Y=1.08 $X2=0 $Y2=0
cc_103 N_A_94_249#_c_111_p N_B2_c_261_n 0.00274772f $X=3.485 $Y=2.035 $X2=0
+ $Y2=0
cc_104 N_A_94_249#_c_76_n N_B1_M1007_g 0.0166797f $X=3.385 $Y=1.08 $X2=0 $Y2=0
cc_105 N_A_94_249#_c_78_n N_B1_M1007_g 0.0148243f $X=3.55 $Y=0.42 $X2=0 $Y2=0
cc_106 N_A_94_249#_c_111_p N_B1_M1004_g 0.0164129f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A_94_249#_c_76_n N_B1_c_294_n 0.00779116f $X=3.385 $Y=1.08 $X2=0 $Y2=0
cc_108 N_A_94_249#_c_84_n N_B1_c_294_n 0.00131037f $X=3.615 $Y=2.14 $X2=0 $Y2=0
cc_109 N_A_94_249#_c_76_n N_B1_c_295_n 0.0238681f $X=3.385 $Y=1.08 $X2=0 $Y2=0
cc_110 N_A_94_249#_c_111_p N_B1_c_295_n 0.00560783f $X=3.485 $Y=2.035 $X2=0
+ $Y2=0
cc_111 N_A_94_249#_c_84_n N_B1_c_295_n 0.0213876f $X=3.615 $Y=2.14 $X2=0 $Y2=0
cc_112 N_A_94_249#_M1008_g N_VPWR_c_321_n 0.00459557f $X=0.545 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_94_249#_M1011_g N_VPWR_c_322_n 0.0103438f $X=0.975 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_94_249#_c_73_n N_VPWR_c_322_n 0.00980784f $X=1.28 $Y=1.08 $X2=0 $Y2=0
cc_115 N_A_94_249#_c_79_n N_VPWR_c_322_n 3.94633e-19 $X=0.995 $Y=1.41 $X2=0
+ $Y2=0
cc_116 N_A_94_249#_M1008_g N_VPWR_c_324_n 0.00564131f $X=0.545 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_94_249#_M1011_g N_VPWR_c_324_n 0.00541359f $X=0.975 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_94_249#_c_85_n N_VPWR_c_326_n 0.0178111f $X=3.58 $Y=2.475 $X2=0 $Y2=0
cc_119 N_A_94_249#_M1010_s N_VPWR_c_319_n 0.00395695f $X=2.595 $Y=1.835 $X2=0
+ $Y2=0
cc_120 N_A_94_249#_M1004_d N_VPWR_c_319_n 0.00371702f $X=3.44 $Y=1.835 $X2=0
+ $Y2=0
cc_121 N_A_94_249#_M1008_g N_VPWR_c_319_n 0.011156f $X=0.545 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_A_94_249#_M1011_g N_VPWR_c_319_n 0.0100721f $X=0.975 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_94_249#_c_85_n N_VPWR_c_319_n 0.0100304f $X=3.58 $Y=2.475 $X2=0 $Y2=0
cc_124 N_A_94_249#_M1008_g N_X_c_373_n 0.0163267f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_94_249#_M1011_g N_X_c_373_n 0.0143022f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_94_249#_M1008_g N_X_c_370_n 0.0178257f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_94_249#_M1001_g N_X_c_370_n 0.00838459f $X=0.62 $Y=0.665 $X2=0 $Y2=0
cc_128 N_A_94_249#_M1011_g N_X_c_370_n 0.00256499f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A_94_249#_M1002_g N_X_c_370_n 8.84541e-19 $X=1.05 $Y=0.665 $X2=0 $Y2=0
cc_130 N_A_94_249#_c_73_n N_X_c_370_n 0.0307257f $X=1.28 $Y=1.08 $X2=0 $Y2=0
cc_131 N_A_94_249#_c_79_n N_X_c_370_n 0.0141736f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_94_249#_M1008_g N_X_c_372_n 0.0104993f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A_94_249#_M1011_g N_X_c_372_n 0.00527327f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A_94_249#_c_73_n N_X_c_372_n 0.00152786f $X=1.28 $Y=1.08 $X2=0 $Y2=0
cc_135 N_A_94_249#_c_79_n N_X_c_372_n 0.00642683f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_94_249#_M1001_g N_X_c_385_n 0.0126056f $X=0.62 $Y=0.665 $X2=0 $Y2=0
cc_137 N_A_94_249#_M1001_g X 0.00317896f $X=0.62 $Y=0.665 $X2=0 $Y2=0
cc_138 N_A_94_249#_c_73_n X 0.00139996f $X=1.28 $Y=1.08 $X2=0 $Y2=0
cc_139 N_A_94_249#_c_79_n X 0.00424802f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_94_249#_c_111_p N_A_326_367#_M1010_d 0.0043882f $X=3.485 $Y=2.035
+ $X2=0 $Y2=0
cc_141 N_A_94_249#_M1010_s N_A_326_367#_c_397_n 0.00714407f $X=2.595 $Y=1.835
+ $X2=0 $Y2=0
cc_142 N_A_94_249#_c_111_p N_A_326_367#_c_397_n 0.039493f $X=3.485 $Y=2.035
+ $X2=0 $Y2=0
cc_143 N_A_94_249#_c_83_n N_A_326_367#_c_397_n 0.0141892f $X=2.62 $Y=2.035 $X2=0
+ $Y2=0
cc_144 N_A_94_249#_c_72_n N_VGND_M1002_s 0.00253506f $X=2.035 $Y=1.08 $X2=0
+ $Y2=0
cc_145 N_A_94_249#_c_73_n N_VGND_M1002_s 0.00107981f $X=1.28 $Y=1.08 $X2=0 $Y2=0
cc_146 N_A_94_249#_c_76_n N_VGND_M1006_s 0.00284759f $X=3.385 $Y=1.08 $X2=0
+ $Y2=0
cc_147 N_A_94_249#_M1001_g N_VGND_c_426_n 0.0211007f $X=0.62 $Y=0.665 $X2=0
+ $Y2=0
cc_148 N_A_94_249#_M1001_g N_VGND_c_427_n 0.00389872f $X=0.62 $Y=0.665 $X2=0
+ $Y2=0
cc_149 N_A_94_249#_M1002_g N_VGND_c_427_n 0.00575161f $X=1.05 $Y=0.665 $X2=0
+ $Y2=0
cc_150 N_A_94_249#_M1002_g N_VGND_c_428_n 0.00650772f $X=1.05 $Y=0.665 $X2=0
+ $Y2=0
cc_151 N_A_94_249#_c_72_n N_VGND_c_428_n 0.0172929f $X=2.035 $Y=1.08 $X2=0 $Y2=0
cc_152 N_A_94_249#_c_73_n N_VGND_c_428_n 0.0087438f $X=1.28 $Y=1.08 $X2=0 $Y2=0
cc_153 N_A_94_249#_c_74_n N_VGND_c_429_n 0.0384285f $X=2.2 $Y=0.42 $X2=0 $Y2=0
cc_154 N_A_94_249#_c_77_n N_VGND_c_429_n 0.0219041f $X=2.62 $Y=1.08 $X2=0 $Y2=0
cc_155 N_A_94_249#_c_78_n N_VGND_c_429_n 0.0190707f $X=3.55 $Y=0.42 $X2=0 $Y2=0
cc_156 N_A_94_249#_c_74_n N_VGND_c_430_n 0.0210467f $X=2.2 $Y=0.42 $X2=0 $Y2=0
cc_157 N_A_94_249#_c_78_n N_VGND_c_431_n 0.0210467f $X=3.55 $Y=0.42 $X2=0 $Y2=0
cc_158 N_A_94_249#_M1000_d N_VGND_c_432_n 0.00212301f $X=2.06 $Y=0.245 $X2=0
+ $Y2=0
cc_159 N_A_94_249#_M1007_d N_VGND_c_432_n 0.00212301f $X=3.41 $Y=0.245 $X2=0
+ $Y2=0
cc_160 N_A_94_249#_M1001_g N_VGND_c_432_n 0.00731027f $X=0.62 $Y=0.665 $X2=0
+ $Y2=0
cc_161 N_A_94_249#_M1002_g N_VGND_c_432_n 0.0110395f $X=1.05 $Y=0.665 $X2=0
+ $Y2=0
cc_162 N_A_94_249#_c_74_n N_VGND_c_432_n 0.0125689f $X=2.2 $Y=0.42 $X2=0 $Y2=0
cc_163 N_A_94_249#_c_78_n N_VGND_c_432_n 0.0125689f $X=3.55 $Y=0.42 $X2=0 $Y2=0
cc_164 N_A_94_249#_c_72_n A_340_49# 0.00366293f $X=2.035 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A_94_249#_c_76_n A_610_49# 0.00366293f $X=3.385 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A2_M1005_g N_A1_M1000_g 0.0478662f $X=1.625 $Y=0.665 $X2=0 $Y2=0
cc_167 N_A2_M1009_g N_A1_M1003_g 0.0177062f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A2_c_185_n N_A1_c_225_n 0.0478662f $X=1.535 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A2_c_186_n N_A1_c_225_n 0.00326328f $X=1.535 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A2_M1009_g N_A1_c_226_n 7.94492e-19 $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A2_c_185_n N_A1_c_226_n 2.38276e-19 $X=1.535 $Y=1.51 $X2=0 $Y2=0
cc_172 N_A2_c_186_n N_A1_c_226_n 0.0314963f $X=1.535 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A2_M1009_g N_VPWR_c_322_n 0.00891046f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A2_c_185_n N_VPWR_c_322_n 0.00228522f $X=1.535 $Y=1.51 $X2=0 $Y2=0
cc_175 N_A2_M1009_g N_VPWR_c_323_n 6.09324e-19 $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A2_M1009_g N_VPWR_c_325_n 0.0054895f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A2_M1009_g N_VPWR_c_319_n 0.0102827f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A2_M1009_g N_X_c_372_n 9.81338e-19 $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A2_M1009_g N_A_326_367#_c_402_n 0.00463867f $X=1.555 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A2_c_185_n N_A_326_367#_c_402_n 3.01661e-19 $X=1.535 $Y=1.51 $X2=0
+ $Y2=0
cc_181 N_A2_c_186_n N_A_326_367#_c_402_n 0.0204033f $X=1.535 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A2_M1009_g N_A_326_367#_c_405_n 0.00658865f $X=1.555 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A2_M1009_g N_A_326_367#_c_406_n 0.00178332f $X=1.555 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A2_M1005_g N_VGND_c_428_n 0.00670511f $X=1.625 $Y=0.665 $X2=0 $Y2=0
cc_185 N_A2_M1005_g N_VGND_c_430_n 0.00575161f $X=1.625 $Y=0.665 $X2=0 $Y2=0
cc_186 N_A2_M1005_g N_VGND_c_432_n 0.0108887f $X=1.625 $Y=0.665 $X2=0 $Y2=0
cc_187 N_A1_c_225_n N_B2_c_261_n 0.00804278f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_188 N_A1_c_226_n N_VPWR_M1003_d 0.00467613f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_189 N_A1_M1003_g N_VPWR_c_323_n 0.0125581f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A1_M1003_g N_VPWR_c_325_n 0.00486043f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A1_M1003_g N_VPWR_c_319_n 0.00458726f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A1_M1003_g N_A_326_367#_c_397_n 0.0161222f $X=1.985 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_A1_c_225_n N_A_326_367#_c_397_n 0.00233696f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_194 N_A1_c_226_n N_A_326_367#_c_397_n 0.0106372f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_195 N_A1_M1000_g N_VGND_c_429_n 0.00334368f $X=1.985 $Y=0.665 $X2=0 $Y2=0
cc_196 N_A1_M1000_g N_VGND_c_430_n 0.00539298f $X=1.985 $Y=0.665 $X2=0 $Y2=0
cc_197 N_A1_M1000_g N_VGND_c_432_n 0.0111162f $X=1.985 $Y=0.665 $X2=0 $Y2=0
cc_198 N_B2_M1006_g N_B1_M1007_g 0.040645f $X=2.975 $Y=0.665 $X2=0 $Y2=0
cc_199 N_B2_M1010_g N_B1_M1004_g 0.0361215f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_200 B2 N_B1_c_294_n 0.00364369f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_201 N_B2_c_261_n N_B1_c_294_n 0.0526347f $X=2.885 $Y=1.51 $X2=0 $Y2=0
cc_202 B2 N_B1_c_295_n 0.0291532f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_203 N_B2_c_261_n N_B1_c_295_n 2.45272e-19 $X=2.885 $Y=1.51 $X2=0 $Y2=0
cc_204 N_B2_M1010_g N_VPWR_c_323_n 0.00949594f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B2_M1010_g N_VPWR_c_326_n 0.0054895f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_206 N_B2_M1010_g N_VPWR_c_319_n 0.00771417f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B2_M1010_g N_A_326_367#_c_397_n 0.0114464f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_208 N_B2_M1010_g N_A_326_367#_c_411_n 0.0170121f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_209 N_B2_M1006_g N_VGND_c_429_n 0.0154267f $X=2.975 $Y=0.665 $X2=0 $Y2=0
cc_210 N_B2_M1006_g N_VGND_c_431_n 0.00477554f $X=2.975 $Y=0.665 $X2=0 $Y2=0
cc_211 N_B2_M1006_g N_VGND_c_432_n 0.00814835f $X=2.975 $Y=0.665 $X2=0 $Y2=0
cc_212 N_B1_M1004_g N_VPWR_c_326_n 0.0054895f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_213 N_B1_M1004_g N_VPWR_c_319_n 0.0108708f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_214 N_B1_M1004_g N_A_326_367#_c_397_n 0.00216614f $X=3.365 $Y=2.465 $X2=0
+ $Y2=0
cc_215 N_B1_M1004_g N_A_326_367#_c_411_n 0.00693633f $X=3.365 $Y=2.465 $X2=0
+ $Y2=0
cc_216 N_B1_M1007_g N_VGND_c_429_n 0.00269887f $X=3.335 $Y=0.665 $X2=0 $Y2=0
cc_217 N_B1_M1007_g N_VGND_c_431_n 0.00539298f $X=3.335 $Y=0.665 $X2=0 $Y2=0
cc_218 N_B1_M1007_g N_VGND_c_432_n 0.0107763f $X=3.335 $Y=0.665 $X2=0 $Y2=0
cc_219 N_VPWR_c_319_n N_X_M1008_d 0.00223559f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_220 N_VPWR_c_324_n N_X_c_373_n 0.0185828f $X=1.1 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_319_n N_X_c_373_n 0.0122144f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_319_n N_A_326_367#_M1009_d 0.00252567f $X=3.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_223 N_VPWR_c_319_n N_A_326_367#_M1010_d 0.00223559f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_325_n N_A_326_367#_c_405_n 0.015688f $X=2.035 $Y=3.33 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_319_n N_A_326_367#_c_405_n 0.00984745f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_226 N_VPWR_M1003_d N_A_326_367#_c_397_n 0.00561481f $X=2.06 $Y=1.835 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_323_n N_A_326_367#_c_397_n 0.021538f $X=2.2 $Y=2.765 $X2=0 $Y2=0
cc_228 N_VPWR_c_319_n N_A_326_367#_c_397_n 0.0255918f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_229 N_VPWR_c_323_n N_A_326_367#_c_411_n 0.0126246f $X=2.2 $Y=2.765 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_326_n N_A_326_367#_c_411_n 0.0189236f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_231 N_VPWR_c_319_n N_A_326_367#_c_411_n 0.0123859f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_232 N_VPWR_c_319_n N_A_326_367#_c_406_n 7.67545e-19 $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_233 N_X_c_385_n N_VGND_c_426_n 0.0656374f $X=0.835 $Y=0.42 $X2=0 $Y2=0
cc_234 N_X_c_385_n N_VGND_c_427_n 0.0228601f $X=0.835 $Y=0.42 $X2=0 $Y2=0
cc_235 N_X_M1001_d N_VGND_c_432_n 0.00345315f $X=0.695 $Y=0.245 $X2=0 $Y2=0
cc_236 N_X_c_385_n N_VGND_c_432_n 0.0136664f $X=0.835 $Y=0.42 $X2=0 $Y2=0
cc_237 N_VGND_c_432_n A_340_49# 0.00899413f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_238 N_VGND_c_432_n A_610_49# 0.00899413f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
