* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand3b_2 A_N B C VGND VNB VPB VPWR Y
M1000 Y a_55_155# a_332_71# VNB nshort w=840000u l=150000u
+  ad=3.948e+11p pd=2.62e+06u as=5.376e+11p ps=4.64e+06u
M1001 Y C VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0584e+12p pd=9.24e+06u as=1.8291e+12p ps=1.313e+07u
M1002 Y a_55_155# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_332_71# a_55_155# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A_N a_55_155# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 a_246_71# C VGND VNB nshort w=840000u l=150000u
+  ad=5.04e+11p pd=4.56e+06u as=4.977e+11p ps=4.67e+06u
M1006 VPWR C Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C a_246_71# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_246_71# B a_332_71# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A_N a_55_155# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1010 a_332_71# B a_246_71# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_55_155# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
