* NGSPICE file created from sky130_fd_sc_lp__ha_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__ha_m A B VGND VNB VPB VPWR COUT SUM
M1000 VGND A a_720_125# VNB nshort w=420000u l=150000u
+  ad=4.224e+11p pd=4.55e+06u as=8.82e+10p ps=1.26e+06u
M1001 VGND a_80_60# SUM VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1002 VPWR a_80_60# SUM VPB phighvt w=420000u l=150000u
+  ad=5.8235e+11p pd=5.54e+06u as=1.113e+11p ps=1.37e+06u
M1003 a_80_60# a_249_212# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1004 COUT a_249_212# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 a_720_125# B a_249_212# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.512e+11p ps=1.56e+06u
M1006 VGND B a_301_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.289e+11p ps=2.77e+06u
M1007 a_301_47# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A a_249_212# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.974e+11p ps=1.78e+06u
M1009 VPWR A a_450_464# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1010 COUT a_249_212# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 a_301_47# a_249_212# a_80_60# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 a_450_464# B a_80_60# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_249_212# B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

