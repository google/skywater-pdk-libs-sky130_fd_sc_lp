* File: sky130_fd_sc_lp__nand3_1.spice
* Created: Wed Sep  2 10:04:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand3_1.pex.spice"
.subckt sky130_fd_sc_lp__nand3_1  VNB VPB C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1005 A_141_76# N_C_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.2226 PD=1.08 PS=2.21 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2 SB=75001.4
+ A=0.126 P=1.98 MULT=1
MM1004 A_219_76# N_B_M1004_g A_141_76# VNB NSHORT L=0.15 W=0.84 AD=0.1764
+ AS=0.1008 PD=1.26 PS=1.08 NRD=22.14 NRS=9.276 M=1 R=5.6 SA=75000.6 SB=75001
+ A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g A_219_76# VNB NSHORT L=0.15 W=0.84 AD=0.4284
+ AS=0.1764 PD=2.7 PS=1.26 NRD=30.708 NRS=22.14 M=1 R=5.6 SA=75001.1 SB=75000.4
+ A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.378 PD=1.54 PS=3.12 NRD=0 NRS=5.4569 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_B_M1002_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2394 AS=0.1764 PD=1.64 PS=1.54 NRD=8.5892 NRS=0 M=1 R=8.4 SA=75000.7
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2394 PD=3.05 PS=1.64 NRD=0 NRS=7.0329 M=1 R=8.4 SA=75001.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__nand3_1.pxi.spice"
*
.ends
*
*
