* File: sky130_fd_sc_lp__o21a_0.pex.spice
* Created: Wed Sep  2 10:15:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21A_0%A_80_23# 1 2 9 11 14 16 17 18 19 21 22 25 29
+ 33 35
c71 33 0 1.36625e-19 $X=0.59 $Y=0.94
c72 19 0 8.64221e-20 $X=1.105 $Y=0.865
r73 33 35 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=0.94
+ $X2=0.577 $Y2=0.775
r74 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=0.94 $X2=0.59 $Y2=0.94
r75 27 29 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=1.3 $Y=2.215
+ $X2=1.3 $Y2=2.56
r76 23 25 13.2051 $w=2.38e-07 $l=2.75e-07 $layer=LI1_cond $X=1.225 $Y=0.775
+ $X2=1.225 $Y2=0.5
r77 21 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.175 $Y=2.13
+ $X2=1.3 $Y2=2.215
r78 21 22 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.175 $Y=2.13
+ $X2=0.755 $Y2=2.13
r79 20 32 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=0.755 $Y=0.865
+ $X2=0.63 $Y2=0.865
r80 19 23 6.999 $w=1.8e-07 $l=1.58745e-07 $layer=LI1_cond $X=1.105 $Y=0.865
+ $X2=1.225 $Y2=0.775
r81 19 20 21.5657 $w=1.78e-07 $l=3.5e-07 $layer=LI1_cond $X=1.105 $Y=0.865
+ $X2=0.755 $Y2=0.865
r82 18 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.63 $Y=2.045
+ $X2=0.755 $Y2=2.13
r83 17 32 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=0.63 $Y=0.955 $X2=0.63
+ $Y2=0.865
r84 17 18 50.2465 $w=2.48e-07 $l=1.09e-06 $layer=LI1_cond $X=0.63 $Y=0.955
+ $X2=0.63 $Y2=2.045
r85 14 16 661.468 $w=1.5e-07 $l=1.29e-06 $layer=POLY_cond $X=0.64 $Y=2.735
+ $X2=0.64 $Y2=1.445
r86 11 16 43.0294 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.577 $Y=1.268
+ $X2=0.577 $Y2=1.445
r87 10 33 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.577 $Y=0.952
+ $X2=0.577 $Y2=0.94
r88 10 11 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.577 $Y=0.952
+ $X2=0.577 $Y2=1.268
r89 9 35 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.455
+ $X2=0.475 $Y2=0.775
r90 2 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.2
+ $Y=2.415 $X2=1.34 $Y2=2.56
r91 1 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.29 $X2=1.21 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_0%B1 3 7 9 11 12 13 16 18 19 23
c53 16 0 1.15274e-19 $X=1.425 $Y=0.895
r54 18 19 11.6802 $w=3.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.18 $Y=1.29
+ $X2=1.18 $Y2=1.665
r55 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=1.29 $X2=1.16 $Y2=1.29
r56 14 16 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.25 $Y=0.895
+ $X2=1.425 $Y2=0.895
r57 12 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.16 $Y=1.63
+ $X2=1.16 $Y2=1.29
r58 12 13 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.63
+ $X2=1.16 $Y2=1.795
r59 11 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.125
+ $X2=1.16 $Y2=1.29
r60 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=0.82
+ $X2=1.425 $Y2=0.895
r61 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.425 $Y=0.82
+ $X2=1.425 $Y2=0.5
r62 5 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.25 $Y=0.97 $X2=1.25
+ $Y2=0.895
r63 5 11 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.25 $Y=0.97
+ $X2=1.25 $Y2=1.125
r64 3 13 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.125 $Y=2.735 $X2=1.125
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_0%A2 2 5 9 11 12 13 14 15 16 23
c48 23 0 9.26367e-20 $X=1.73 $Y=1.375
c49 9 0 8.64221e-20 $X=1.855 $Y=0.5
r50 23 25 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.732 $Y=1.375
+ $X2=1.732 $Y2=1.21
r51 15 16 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=2.405
+ $X2=1.717 $Y2=2.775
r52 14 15 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=2.035
+ $X2=1.717 $Y2=2.405
r53 13 14 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=1.665
+ $X2=1.717 $Y2=2.035
r54 12 13 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=1.295
+ $X2=1.717 $Y2=1.665
r55 12 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=1.375 $X2=1.73 $Y2=1.375
r56 9 25 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.855 $Y=0.5
+ $X2=1.855 $Y2=1.21
r57 5 11 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.61 $Y=2.735
+ $X2=1.61 $Y2=1.88
r58 2 11 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=1.732 $Y=1.683
+ $X2=1.732 $Y2=1.88
r59 1 23 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=1.732 $Y=1.407
+ $X2=1.732 $Y2=1.375
r60 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=1.732 $Y=1.407
+ $X2=1.732 $Y2=1.683
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_0%A1 3 7 12 16 17 18 23
r29 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.335
+ $Y=1.72 $X2=2.335 $Y2=1.72
r30 18 24 6.91311 $w=5.43e-07 $l=3.15e-07 $layer=LI1_cond $X=2.282 $Y=2.035
+ $X2=2.282 $Y2=1.72
r31 17 24 1.20705 $w=5.43e-07 $l=5.5e-08 $layer=LI1_cond $X=2.282 $Y=1.665
+ $X2=2.282 $Y2=1.72
r32 16 17 8.12016 $w=5.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.282 $Y=1.295
+ $X2=2.282 $Y2=1.665
r33 15 23 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.555
+ $X2=2.335 $Y2=1.72
r34 12 23 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=2.335 $Y=2.12
+ $X2=2.335 $Y2=1.72
r35 9 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.97 $Y=2.195
+ $X2=2.335 $Y2=2.195
r36 7 15 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=2.285 $Y=0.5
+ $X2=2.285 $Y2=1.555
r37 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.97 $Y=2.27 $X2=1.97
+ $Y2=2.195
r38 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.97 $Y=2.27 $X2=1.97
+ $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_0%X 1 2 9 12 13 14 15 16 32
r17 32 33 2.9837 $w=4.78e-07 $l=1e-08 $layer=LI1_cond $X=0.325 $Y=2.405
+ $X2=0.325 $Y2=2.395
r18 16 36 5.35743 $w=4.78e-07 $l=2.15e-07 $layer=LI1_cond $X=0.325 $Y=2.775
+ $X2=0.325 $Y2=2.56
r19 15 36 2.94036 $w=4.78e-07 $l=1.18e-07 $layer=LI1_cond $X=0.325 $Y=2.442
+ $X2=0.325 $Y2=2.56
r20 15 32 0.921977 $w=4.78e-07 $l=3.7e-08 $layer=LI1_cond $X=0.325 $Y=2.442
+ $X2=0.325 $Y2=2.405
r21 15 33 1.75171 $w=2.48e-07 $l=3.8e-08 $layer=LI1_cond $X=0.21 $Y=2.357
+ $X2=0.21 $Y2=2.395
r22 14 15 14.8435 $w=2.48e-07 $l=3.22e-07 $layer=LI1_cond $X=0.21 $Y=2.035
+ $X2=0.21 $Y2=2.357
r23 13 14 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=2.035
r24 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.295
+ $X2=0.21 $Y2=1.665
r25 11 12 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=0.21 $Y=0.605
+ $X2=0.21 $Y2=1.295
r26 9 11 6.55995 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.242 $Y=0.44
+ $X2=0.242 $Y2=0.605
r27 2 36 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.3
+ $Y=2.415 $X2=0.425 $Y2=2.56
r28 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.245 $X2=0.26 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_0%VPWR 1 2 9 13 16 17 18 24 30 31 34
r35 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.185 $Y2=3.33
r39 28 30 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.02 $Y=3.33
+ $X2=2.185 $Y2=3.33
r43 24 26 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.02 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 18 22 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 16 21 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 16 17 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.87 $Y2=3.33
r49 15 26 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 15 17 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.87 $Y2=3.33
r51 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=3.245
+ $X2=2.185 $Y2=3.33
r52 11 13 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.185 $Y=3.245
+ $X2=2.185 $Y2=2.56
r53 7 17 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=3.33
r54 7 9 29.2379 $w=2.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=2.56
r55 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=2.415 $X2=2.185 $Y2=2.56
r56 1 9 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.715
+ $Y=2.415 $X2=0.9 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_0%VGND 1 2 9 13 16 17 18 20 30 31 34
c37 31 0 1.15274e-19 $X=2.64 $Y=0
c38 20 0 1.36625e-19 $X=0.57 $Y=0
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r42 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r43 25 34 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.712
+ $Y2=0
r44 25 27 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.68
+ $Y2=0
r45 23 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r46 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 20 34 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.712
+ $Y2=0
r48 20 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.24
+ $Y2=0
r49 18 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r50 18 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r51 16 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.68
+ $Y2=0
r52 16 17 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.07
+ $Y2=0
r53 15 30 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.64
+ $Y2=0
r54 15 17 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.07
+ $Y2=0
r55 11 17 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0
r56 11 13 17.7135 $w=2.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0.5
r57 7 34 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0
r58 7 9 14.355 $w=2.83e-07 $l=3.55e-07 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0.44
r59 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.29 $X2=2.07 $Y2=0.5
r60 1 9 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.245 $X2=0.69 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_0%A_300_58# 1 2 9 11 12 15
c25 11 0 9.26367e-20 $X=2.375 $Y=0.92
r26 13 15 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.52 $Y=0.835
+ $X2=2.52 $Y2=0.5
r27 11 13 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.375 $Y=0.92
+ $X2=2.52 $Y2=0.835
r28 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.375 $Y=0.92
+ $X2=1.765 $Y2=0.92
r29 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.64 $Y=0.835
+ $X2=1.765 $Y2=0.92
r30 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.64 $Y=0.835
+ $X2=1.64 $Y2=0.5
r31 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.29 $X2=2.5 $Y2=0.5
r32 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.29 $X2=1.64 $Y2=0.5
.ends

