* File: sky130_fd_sc_lp__o31a_2.pxi.spice
* Created: Wed Sep  2 10:24:37 2020
* 
x_PM_SKY130_FD_SC_LP__O31A_2%A_85_21# N_A_85_21#_M1003_d N_A_85_21#_M1005_d
+ N_A_85_21#_c_64_n N_A_85_21#_M1010_g N_A_85_21#_M1002_g N_A_85_21#_c_66_n
+ N_A_85_21#_M1011_g N_A_85_21#_M1008_g N_A_85_21#_c_68_n N_A_85_21#_c_69_n
+ N_A_85_21#_c_140_p N_A_85_21#_c_70_n N_A_85_21#_c_110_p N_A_85_21#_c_71_n
+ N_A_85_21#_c_72_n N_A_85_21#_c_73_n N_A_85_21#_c_74_n N_A_85_21#_c_103_p
+ N_A_85_21#_c_75_n PM_SKY130_FD_SC_LP__O31A_2%A_85_21#
x_PM_SKY130_FD_SC_LP__O31A_2%A1 N_A1_M1007_g N_A1_M1001_g A1 A1 A1 A1
+ N_A1_c_165_n N_A1_c_166_n A1 PM_SKY130_FD_SC_LP__O31A_2%A1
x_PM_SKY130_FD_SC_LP__O31A_2%A2 N_A2_M1006_g N_A2_M1000_g A2 A2 A2 A2
+ N_A2_c_209_n N_A2_c_212_n PM_SKY130_FD_SC_LP__O31A_2%A2
x_PM_SKY130_FD_SC_LP__O31A_2%A3 N_A3_M1005_g N_A3_M1004_g A3 N_A3_c_242_n
+ N_A3_c_243_n PM_SKY130_FD_SC_LP__O31A_2%A3
x_PM_SKY130_FD_SC_LP__O31A_2%B1 N_B1_M1003_g N_B1_M1009_g B1 N_B1_c_276_n
+ PM_SKY130_FD_SC_LP__O31A_2%B1
x_PM_SKY130_FD_SC_LP__O31A_2%VPWR N_VPWR_M1002_d N_VPWR_M1008_d N_VPWR_M1009_d
+ N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n N_VPWR_c_308_n N_VPWR_c_309_n
+ N_VPWR_c_310_n VPWR N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_304_n
+ N_VPWR_c_314_n PM_SKY130_FD_SC_LP__O31A_2%VPWR
x_PM_SKY130_FD_SC_LP__O31A_2%X N_X_M1010_s N_X_M1002_s X X X X X X X N_X_c_353_n
+ X PM_SKY130_FD_SC_LP__O31A_2%X
x_PM_SKY130_FD_SC_LP__O31A_2%VGND N_VGND_M1010_d N_VGND_M1011_d N_VGND_M1000_d
+ N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n
+ N_VGND_c_386_n VGND N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n
+ N_VGND_c_390_n PM_SKY130_FD_SC_LP__O31A_2%VGND
x_PM_SKY130_FD_SC_LP__O31A_2%A_355_47# N_A_355_47#_M1007_d N_A_355_47#_M1004_d
+ N_A_355_47#_c_439_n N_A_355_47#_c_443_n N_A_355_47#_c_440_n
+ N_A_355_47#_c_441_n N_A_355_47#_c_447_n PM_SKY130_FD_SC_LP__O31A_2%A_355_47#
cc_1 VNB N_A_85_21#_c_64_n 0.0215279f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_2 VNB N_A_85_21#_M1002_g 0.0106048f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.465
cc_3 VNB N_A_85_21#_c_66_n 0.0177327f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.185
cc_4 VNB N_A_85_21#_M1008_g 0.00784791f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.465
cc_5 VNB N_A_85_21#_c_68_n 0.00407386f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.35
cc_6 VNB N_A_85_21#_c_69_n 0.0729787f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.35
cc_7 VNB N_A_85_21#_c_70_n 0.0149562f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.09
cc_8 VNB N_A_85_21#_c_71_n 0.00994307f $X=-0.19 $Y=-0.245 $X2=3.39 $Y2=1.005
cc_9 VNB N_A_85_21#_c_72_n 0.0285946f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=0.42
cc_10 VNB N_A_85_21#_c_73_n 0.00621528f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=1.105
cc_11 VNB N_A_85_21#_c_74_n 0.00476225f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.105
cc_12 VNB N_A_85_21#_c_75_n 0.00384551f $X=-0.19 $Y=-0.245 $X2=2.917 $Y2=1.93
cc_13 VNB N_A1_M1007_g 0.0278603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_165_n 0.0246834f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.465
cc_15 VNB N_A1_c_166_n 0.00207116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_M1000_g 0.025042f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_17 VNB N_A2_c_209_n 0.0257976f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.465
cc_18 VNB N_A3_M1004_g 0.0248639f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_19 VNB N_A3_c_242_n 0.0259195f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.465
cc_20 VNB N_A3_c_243_n 0.00100522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_M1003_g 0.033049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB B1 0.0198394f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_23 VNB N_B1_c_276_n 0.0372306f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.185
cc_24 VNB N_VPWR_c_304_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_353_n 0.0028991f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.35
cc_26 VNB N_VGND_c_381_n 0.0113184f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.515
cc_27 VNB N_VGND_c_382_n 0.0484565f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.465
cc_28 VNB N_VGND_c_383_n 0.00372231f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.655
cc_29 VNB N_VGND_c_384_n 4.2118e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_385_n 0.0162836f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.35
cc_31 VNB N_VGND_c_386_n 0.00436333f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.35
cc_32 VNB N_VGND_c_387_n 0.0156137f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.12
cc_33 VNB N_VGND_c_388_n 0.0345135f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=1.105
cc_34 VNB N_VGND_c_389_n 0.218205f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.105
cc_35 VNB N_VGND_c_390_n 0.0104501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_A_85_21#_M1002_g 0.0264965f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.465
cc_37 VPB N_A_85_21#_M1008_g 0.022304f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.465
cc_38 VPB N_A_85_21#_c_75_n 0.00147446f $X=-0.19 $Y=1.655 $X2=2.917 $Y2=1.93
cc_39 VPB N_A1_M1001_g 0.01917f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.185
cc_40 VPB A1 0.00278174f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.655
cc_41 VPB N_A1_c_165_n 0.00650311f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.465
cc_42 VPB N_A1_c_166_n 0.00303419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A2_M1006_g 0.0187009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A2_c_209_n 0.00647392f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.465
cc_45 VPB N_A2_c_212_n 0.00135437f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.465
cc_46 VPB N_A3_M1005_g 0.0211196f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A3_c_242_n 0.00617499f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.465
cc_48 VPB N_A3_c_243_n 0.00254201f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B1_M1009_g 0.0247497f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.185
cc_50 VPB B1 0.0153109f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.655
cc_51 VPB N_B1_c_276_n 0.0133238f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.185
cc_52 VPB N_VPWR_c_305_n 0.0123094f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.515
cc_53 VPB N_VPWR_c_306_n 0.064594f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.465
cc_54 VPB N_VPWR_c_307_n 0.00847352f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.465
cc_55 VPB N_VPWR_c_308_n 0.0468692f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.35
cc_56 VPB N_VPWR_c_309_n 0.0531442f $X=-0.19 $Y=1.655 $X2=1.93 $Y2=1.09
cc_57 VPB N_VPWR_c_310_n 0.00420242f $X=-0.19 $Y=1.655 $X2=2.917 $Y2=2.137
cc_58 VPB N_VPWR_c_311_n 0.0183613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_312_n 0.0124854f $X=-0.19 $Y=1.655 $X2=3.39 $Y2=1.09
cc_60 VPB N_VPWR_c_304_n 0.055674f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_314_n 0.0047828f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.35
cc_62 VPB X 0.00305456f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.515
cc_63 VPB N_X_c_353_n 3.66861e-19 $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.35
cc_64 N_A_85_21#_c_66_n N_A1_M1007_g 0.00732805f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_65 N_A_85_21#_c_68_n N_A1_M1007_g 8.06595e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_66 N_A_85_21#_c_69_n N_A1_M1007_g 0.00568669f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_67 N_A_85_21#_c_73_n N_A1_M1007_g 0.0130834f $X=1.76 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_85_21#_c_74_n N_A1_M1007_g 0.00466644f $X=1.93 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A_85_21#_M1008_g N_A1_M1001_g 0.0207853f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_85_21#_M1008_g A1 0.00288892f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_71 N_A_85_21#_M1008_g N_A1_c_165_n 0.00441116f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_72 N_A_85_21#_c_68_n N_A1_c_165_n 7.03201e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_73 N_A_85_21#_c_69_n N_A1_c_165_n 0.0112341f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_74 N_A_85_21#_c_73_n N_A1_c_165_n 0.0041938f $X=1.76 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_85_21#_M1008_g N_A1_c_166_n 6.22181e-19 $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_76 N_A_85_21#_c_68_n N_A1_c_166_n 0.00876587f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_77 N_A_85_21#_c_69_n N_A1_c_166_n 5.64994e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_78 N_A_85_21#_c_73_n N_A1_c_166_n 0.0286508f $X=1.76 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_85_21#_c_70_n N_A2_M1000_g 0.011003f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_80 N_A_85_21#_c_74_n N_A2_M1000_g 7.88849e-19 $X=1.93 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A_85_21#_c_70_n N_A2_c_209_n 0.00471777f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_82 N_A_85_21#_c_70_n N_A2_c_212_n 0.0226002f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_83 N_A_85_21#_c_75_n N_A2_c_212_n 0.00529995f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_84 N_A_85_21#_c_75_n N_A3_M1005_g 0.0018621f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_85 N_A_85_21#_c_70_n N_A3_M1004_g 0.0107724f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_86 N_A_85_21#_c_75_n N_A3_M1004_g 0.00333584f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_87 N_A_85_21#_c_70_n N_A3_c_242_n 0.00342488f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_88 N_A_85_21#_c_103_p N_A3_c_242_n 0.0032981f $X=2.875 $Y=2.095 $X2=0 $Y2=0
cc_89 N_A_85_21#_c_75_n N_A3_c_242_n 0.00200461f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_90 N_A_85_21#_c_70_n N_A3_c_243_n 0.0192331f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_91 N_A_85_21#_c_103_p N_A3_c_243_n 0.00528262f $X=2.875 $Y=2.095 $X2=0 $Y2=0
cc_92 N_A_85_21#_c_75_n N_A3_c_243_n 0.0301899f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_93 N_A_85_21#_c_71_n N_B1_M1003_g 0.0167221f $X=3.39 $Y=1.005 $X2=0 $Y2=0
cc_94 N_A_85_21#_c_75_n N_B1_M1003_g 0.00882031f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_95 N_A_85_21#_c_110_p N_B1_M1009_g 0.0131688f $X=2.875 $Y=2.91 $X2=0 $Y2=0
cc_96 N_A_85_21#_c_103_p N_B1_M1009_g 0.00269421f $X=2.875 $Y=2.095 $X2=0 $Y2=0
cc_97 N_A_85_21#_c_75_n N_B1_M1009_g 0.0104173f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_98 N_A_85_21#_c_71_n B1 0.0164155f $X=3.39 $Y=1.005 $X2=0 $Y2=0
cc_99 N_A_85_21#_c_75_n B1 0.0286136f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_100 N_A_85_21#_c_71_n N_B1_c_276_n 0.00820138f $X=3.39 $Y=1.005 $X2=0 $Y2=0
cc_101 N_A_85_21#_c_75_n N_B1_c_276_n 0.00797462f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_102 N_A_85_21#_M1002_g N_VPWR_c_306_n 0.00885808f $X=0.535 $Y=2.465 $X2=0
+ $Y2=0
cc_103 N_A_85_21#_M1008_g N_VPWR_c_307_n 0.0172761f $X=0.965 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_A_85_21#_c_68_n N_VPWR_c_307_n 0.00718631f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_105 N_A_85_21#_c_69_n N_VPWR_c_307_n 9.42641e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_106 N_A_85_21#_c_73_n N_VPWR_c_307_n 0.00408014f $X=1.76 $Y=1.105 $X2=0 $Y2=0
cc_107 N_A_85_21#_c_75_n N_VPWR_c_308_n 0.0883576f $X=2.917 $Y=1.93 $X2=0 $Y2=0
cc_108 N_A_85_21#_c_110_p N_VPWR_c_309_n 0.0261633f $X=2.875 $Y=2.91 $X2=0 $Y2=0
cc_109 N_A_85_21#_M1002_g N_VPWR_c_311_n 0.00564131f $X=0.535 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_85_21#_M1008_g N_VPWR_c_311_n 0.0054895f $X=0.965 $Y=2.465 $X2=0
+ $Y2=0
cc_111 N_A_85_21#_M1005_d N_VPWR_c_304_n 0.00439065f $X=2.675 $Y=1.835 $X2=0
+ $Y2=0
cc_112 N_A_85_21#_M1002_g N_VPWR_c_304_n 0.0110936f $X=0.535 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_85_21#_M1008_g N_VPWR_c_304_n 0.0105673f $X=0.965 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_85_21#_c_110_p N_VPWR_c_304_n 0.0157133f $X=2.875 $Y=2.91 $X2=0 $Y2=0
cc_115 N_A_85_21#_M1002_g X 0.00715749f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_85_21#_M1008_g X 0.00595538f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_85_21#_M1002_g X 0.0140624f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_85_21#_M1008_g X 0.0156202f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_85_21#_c_64_n N_X_c_353_n 0.00314882f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_120 N_A_85_21#_M1002_g N_X_c_353_n 0.008786f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_85_21#_c_66_n N_X_c_353_n 0.0014112f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_122 N_A_85_21#_M1008_g N_X_c_353_n 0.00248806f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_85_21#_c_68_n N_X_c_353_n 0.0220423f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_124 N_A_85_21#_c_69_n N_X_c_353_n 0.0293729f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_125 N_A_85_21#_c_140_p N_X_c_353_n 0.0121102f $X=1.235 $Y=1.12 $X2=0 $Y2=0
cc_126 N_A_85_21#_c_140_p N_VGND_M1011_d 0.00188328f $X=1.235 $Y=1.12 $X2=0
+ $Y2=0
cc_127 N_A_85_21#_c_73_n N_VGND_M1011_d 0.00359398f $X=1.76 $Y=1.105 $X2=0 $Y2=0
cc_128 N_A_85_21#_c_70_n N_VGND_M1000_d 0.00176891f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_129 N_A_85_21#_c_64_n N_VGND_c_382_n 0.00689436f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_130 N_A_85_21#_c_64_n N_VGND_c_383_n 6.51537e-19 $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_131 N_A_85_21#_c_66_n N_VGND_c_383_n 0.0111209f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_132 N_A_85_21#_c_69_n N_VGND_c_383_n 0.0011379f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_133 N_A_85_21#_c_140_p N_VGND_c_383_n 0.0167321f $X=1.235 $Y=1.12 $X2=0 $Y2=0
cc_134 N_A_85_21#_c_73_n N_VGND_c_383_n 0.0270559f $X=1.76 $Y=1.105 $X2=0 $Y2=0
cc_135 N_A_85_21#_c_64_n N_VGND_c_387_n 0.00585385f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_136 N_A_85_21#_c_66_n N_VGND_c_387_n 0.00505556f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_137 N_A_85_21#_c_72_n N_VGND_c_388_n 0.0178111f $X=3.355 $Y=0.42 $X2=0 $Y2=0
cc_138 N_A_85_21#_M1003_d N_VGND_c_389_n 0.00371702f $X=3.215 $Y=0.235 $X2=0
+ $Y2=0
cc_139 N_A_85_21#_c_64_n N_VGND_c_389_n 0.0115325f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_140 N_A_85_21#_c_66_n N_VGND_c_389_n 0.00855618f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_141 N_A_85_21#_c_72_n N_VGND_c_389_n 0.0100304f $X=3.355 $Y=0.42 $X2=0 $Y2=0
cc_142 N_A_85_21#_c_70_n N_A_355_47#_M1007_d 0.00156264f $X=2.955 $Y=1.09
+ $X2=-0.19 $Y2=-0.245
cc_143 N_A_85_21#_c_74_n N_A_355_47#_M1007_d 0.00104699f $X=1.93 $Y=1.105
+ $X2=-0.19 $Y2=-0.245
cc_144 N_A_85_21#_c_70_n N_A_355_47#_M1004_d 0.0019347f $X=2.955 $Y=1.09 $X2=0
+ $Y2=0
cc_145 N_A_85_21#_c_71_n N_A_355_47#_M1004_d 5.634e-19 $X=3.39 $Y=1.005 $X2=0
+ $Y2=0
cc_146 N_A_85_21#_c_74_n N_A_355_47#_c_439_n 0.0209088f $X=1.93 $Y=1.105 $X2=0
+ $Y2=0
cc_147 N_A_85_21#_c_70_n N_A_355_47#_c_440_n 0.0323912f $X=2.955 $Y=1.09 $X2=0
+ $Y2=0
cc_148 N_A_85_21#_c_70_n N_A_355_47#_c_441_n 0.0207563f $X=2.955 $Y=1.09 $X2=0
+ $Y2=0
cc_149 N_A1_M1001_g N_A2_M1006_g 0.0571581f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_150 A1 N_A2_M1006_g 0.00268365f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A1_M1007_g N_A2_M1000_g 0.0294622f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_152 N_A1_c_165_n N_A2_c_209_n 0.0571581f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_153 N_A1_c_166_n N_A2_c_209_n 0.00268365f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_154 N_A1_c_165_n N_A2_c_212_n 0.00182591f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A1_c_166_n N_A2_c_212_n 0.0780236f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_156 A1 N_VPWR_M1008_d 0.0111664f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A1_M1001_g N_VPWR_c_307_n 0.00898558f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_158 A1 N_VPWR_c_307_n 0.0875853f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_159 N_A1_M1001_g N_VPWR_c_309_n 0.00383378f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_160 A1 N_VPWR_c_309_n 0.00897846f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_161 N_A1_M1001_g N_VPWR_c_304_n 0.00599137f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_162 A1 N_VPWR_c_304_n 0.00967541f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_163 A1 X 0.0037137f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A1_c_166_n N_X_c_353_n 0.00452578f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A1_M1007_g N_VGND_c_383_n 0.00219585f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_166 N_A1_M1007_g N_VGND_c_384_n 4.55611e-19 $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_167 N_A1_M1007_g N_VGND_c_385_n 0.00564131f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A1_M1007_g N_VGND_c_389_n 0.0109563f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_169 N_A1_M1007_g N_A_355_47#_c_439_n 0.00188832f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_170 N_A1_M1007_g N_A_355_47#_c_443_n 0.00418638f $X=1.7 $Y=0.655 $X2=0 $Y2=0
cc_171 N_A2_M1006_g N_A3_M1005_g 0.0421157f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A2_c_212_n N_A3_M1005_g 0.0119019f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A2_M1000_g N_A3_M1004_g 0.0419786f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A2_c_209_n N_A3_c_242_n 0.0203109f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_175 N_A2_c_212_n N_A3_c_242_n 0.00104487f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A2_c_209_n N_A3_c_243_n 0.00126086f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A2_c_212_n N_A3_c_243_n 0.0236232f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_178 N_A2_M1006_g N_VPWR_c_309_n 0.00384725f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A2_c_212_n N_VPWR_c_309_n 0.0111904f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A2_M1006_g N_VPWR_c_304_n 0.00563009f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A2_c_212_n N_VPWR_c_304_n 0.011126f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A2_c_212_n A_427_367# 0.015501f $X=2.15 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_183 N_A2_M1000_g N_VGND_c_384_n 0.00704326f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_184 N_A2_M1000_g N_VGND_c_385_n 0.0035715f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_185 N_A2_M1000_g N_VGND_c_389_n 0.00447519f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_186 N_A2_M1000_g N_A_355_47#_c_440_n 0.0120633f $X=2.21 $Y=0.655 $X2=0 $Y2=0
cc_187 N_A3_M1004_g N_B1_M1003_g 0.0283256f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A3_M1005_g N_B1_M1009_g 0.0238891f $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A3_c_243_n N_B1_M1009_g 2.11552e-19 $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A3_c_242_n N_B1_c_276_n 0.02049f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A3_c_243_n N_B1_c_276_n 2.96922e-19 $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_192 N_A3_M1005_g N_VPWR_c_309_n 0.00585385f $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A3_M1005_g N_VPWR_c_304_n 0.011557f $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A3_M1004_g N_VGND_c_384_n 0.00793352f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A3_M1004_g N_VGND_c_388_n 0.0035715f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A3_M1004_g N_VGND_c_389_n 0.00445236f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_197 N_A3_M1004_g N_A_355_47#_c_440_n 0.0120146f $X=2.64 $Y=0.655 $X2=0 $Y2=0
cc_198 N_B1_M1009_g N_VPWR_c_308_n 0.00937945f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_199 B1 N_VPWR_c_308_n 0.0184088f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_200 N_B1_c_276_n N_VPWR_c_308_n 0.00173378f $X=3.39 $Y=1.51 $X2=0 $Y2=0
cc_201 N_B1_M1009_g N_VPWR_c_309_n 0.00495816f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B1_M1009_g N_VPWR_c_304_n 0.0099189f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B1_M1003_g N_VGND_c_384_n 9.91773e-19 $X=3.14 $Y=0.655 $X2=0 $Y2=0
cc_204 N_B1_M1003_g N_VGND_c_388_n 0.0054895f $X=3.14 $Y=0.655 $X2=0 $Y2=0
cc_205 N_B1_M1003_g N_VGND_c_389_n 0.011185f $X=3.14 $Y=0.655 $X2=0 $Y2=0
cc_206 N_B1_M1003_g N_A_355_47#_c_441_n 0.00214936f $X=3.14 $Y=0.655 $X2=0 $Y2=0
cc_207 N_B1_M1003_g N_A_355_47#_c_447_n 0.00455395f $X=3.14 $Y=0.655 $X2=0 $Y2=0
cc_208 N_VPWR_c_304_n N_X_M1002_s 0.00223559f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_209 N_VPWR_c_306_n X 0.0477854f $X=0.32 $Y=1.98 $X2=0 $Y2=0
cc_210 N_VPWR_c_307_n X 0.0873179f $X=1.27 $Y=1.985 $X2=0 $Y2=0
cc_211 N_VPWR_c_311_n X 0.0182419f $X=1.105 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_304_n X 0.0120429f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_304_n A_355_367# 0.00766008f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_214 N_VPWR_c_304_n A_427_367# 0.0105905f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_215 N_X_c_353_n N_VGND_c_382_n 0.00134887f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_216 N_X_c_353_n N_VGND_c_387_n 0.0135169f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_217 N_X_M1010_s N_VGND_c_389_n 0.00432284f $X=0.575 $Y=0.235 $X2=0 $Y2=0
cc_218 N_X_c_353_n N_VGND_c_389_n 0.00847534f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_219 N_VGND_c_389_n N_A_355_47#_M1007_d 0.00305995f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_220 N_VGND_c_389_n N_A_355_47#_M1004_d 0.00297953f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_c_385_n N_A_355_47#_c_443_n 0.0204214f $X=2.26 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_389_n N_A_355_47#_c_443_n 0.0125622f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_M1000_d N_A_355_47#_c_440_n 0.00347417f $X=2.285 $Y=0.235 $X2=0
+ $Y2=0
cc_224 N_VGND_c_384_n N_A_355_47#_c_440_n 0.0161464f $X=2.425 $Y=0.37 $X2=0
+ $Y2=0
cc_225 N_VGND_c_385_n N_A_355_47#_c_440_n 0.00230386f $X=2.26 $Y=0 $X2=0 $Y2=0
cc_226 N_VGND_c_388_n N_A_355_47#_c_440_n 0.00230386f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_227 N_VGND_c_389_n N_A_355_47#_c_440_n 0.00966916f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_388_n N_A_355_47#_c_447_n 0.0204003f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_c_389_n N_A_355_47#_c_447_n 0.0125165f $X=3.6 $Y=0 $X2=0 $Y2=0
