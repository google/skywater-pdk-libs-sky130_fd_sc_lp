* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor3_lp A B C VGND VNB VPB VPWR Y
X0 a_395_409# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_489_57# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_173_57# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND B a_331_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_331_57# B Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y C a_297_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 Y C a_173_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_297_409# B a_395_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 Y A a_489_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
