# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__dlymetal6s6s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dlymetal6s6s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.315000 0.550000 1.765000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.960000 2.320000 4.205000 2.490000 ;
        RECT 3.840000 1.920000 4.205000 2.320000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 4.320000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 4.510000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.095000  0.700000 0.390000 0.975000 ;
      RECT 0.095000  0.975000 0.890000 1.145000 ;
      RECT 0.095000  1.935000 0.890000 2.160000 ;
      RECT 0.095000  2.160000 0.425000 2.225000 ;
      RECT 0.585000  0.085000 0.915000 0.805000 ;
      RECT 0.585000  2.330000 0.880000 3.245000 ;
      RECT 0.720000  1.145000 0.890000 1.275000 ;
      RECT 0.720000  1.275000 1.010000 1.605000 ;
      RECT 0.720000  1.605000 0.890000 1.935000 ;
      RECT 1.060000  1.835000 1.350000 3.075000 ;
      RECT 1.085000  0.255000 1.350000 1.075000 ;
      RECT 1.180000  1.075000 1.350000 1.315000 ;
      RECT 1.180000  1.315000 1.990000 1.605000 ;
      RECT 1.180000  1.605000 1.350000 1.835000 ;
      RECT 1.535000  0.700000 1.830000 0.975000 ;
      RECT 1.535000  0.975000 2.330000 1.145000 ;
      RECT 1.535000  1.895000 2.330000 2.160000 ;
      RECT 1.535000  2.160000 1.865000 2.225000 ;
      RECT 2.025000  0.085000 2.355000 0.805000 ;
      RECT 2.025000  2.330000 2.320000 3.245000 ;
      RECT 2.160000  1.145000 2.330000 1.275000 ;
      RECT 2.160000  1.275000 2.450000 1.605000 ;
      RECT 2.160000  1.605000 2.330000 1.895000 ;
      RECT 2.500000  1.835000 2.790000 3.075000 ;
      RECT 2.525000  0.255000 2.790000 1.075000 ;
      RECT 2.620000  1.075000 2.790000 1.315000 ;
      RECT 2.620000  1.315000 3.430000 1.605000 ;
      RECT 2.620000  1.605000 2.790000 1.835000 ;
      RECT 2.975000  0.700000 3.270000 0.975000 ;
      RECT 2.975000  0.975000 3.770000 1.145000 ;
      RECT 2.975000  1.895000 3.770000 2.160000 ;
      RECT 2.975000  2.160000 3.305000 2.225000 ;
      RECT 3.465000  0.085000 3.795000 0.805000 ;
      RECT 3.465000  2.330000 3.760000 3.245000 ;
      RECT 3.600000  1.145000 3.770000 1.275000 ;
      RECT 3.600000  1.275000 3.890000 1.605000 ;
      RECT 3.600000  1.605000 3.770000 1.895000 ;
      RECT 3.940000  1.835000 4.235000 3.075000 ;
      RECT 3.965000  0.255000 4.235000 1.075000 ;
      RECT 4.060000  1.075000 4.235000 1.835000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.095000  1.950000 1.265000 2.120000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.535000  1.950000 2.705000 2.120000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.975000  1.950000 4.145000 2.120000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
    LAYER met1 ;
      RECT 0.960000 1.920000 1.325000 2.150000 ;
      RECT 2.400000 1.920000 2.765000 2.150000 ;
  END
END sky130_fd_sc_lp__dlymetal6s6s_1
END LIBRARY
