# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.210000 2.325000 1.880000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.230000 0.255000 10.455000 3.075000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.625000 2.235000 5.665000 2.565000 ;
        RECT 5.495000 2.565000 5.665000 2.905000 ;
        RECT 5.495000 2.905000 7.035000 3.075000 ;
        RECT 6.865000 2.295000 7.385000 2.605000 ;
        RECT 6.865000 2.605000 7.035000 2.905000 ;
        RECT 7.215000 1.745000 8.495000 2.015000 ;
        RECT 7.215000 2.015000 7.385000 2.295000 ;
        RECT 8.035000 2.015000 8.495000 2.255000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.450000 0.470000 2.120000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.095000  0.545000  0.390000 1.100000 ;
      RECT  0.095000  1.100000  1.125000 1.270000 ;
      RECT  0.095000  2.300000  0.835000 2.470000 ;
      RECT  0.095000  2.470000  0.355000 2.970000 ;
      RECT  0.525000  2.640000  0.855000 3.245000 ;
      RECT  0.560000  0.085000  0.785000 0.880000 ;
      RECT  0.665000  1.270000  1.125000 1.705000 ;
      RECT  0.665000  1.705000  0.835000 2.300000 ;
      RECT  0.955000  0.255000  1.825000 0.425000 ;
      RECT  0.955000  0.425000  1.125000 1.100000 ;
      RECT  1.025000  2.085000  2.905000 2.255000 ;
      RECT  1.025000  2.255000  1.285000 2.970000 ;
      RECT  1.295000  0.595000  1.485000 1.500000 ;
      RECT  1.295000  1.500000  1.825000 1.830000 ;
      RECT  1.295000  1.830000  1.475000 2.085000 ;
      RECT  1.550000  2.425000  3.245000 2.595000 ;
      RECT  1.550000  2.595000  1.810000 3.050000 ;
      RECT  1.655000  0.425000  1.825000 0.870000 ;
      RECT  1.655000  0.870000  2.580000 1.040000 ;
      RECT  1.980000  2.765000  2.310000 3.245000 ;
      RECT  1.995000  0.085000  2.240000 0.700000 ;
      RECT  2.410000  0.255000  4.220000 0.470000 ;
      RECT  2.410000  0.470000  2.580000 0.870000 ;
      RECT  2.480000  2.595000  2.700000 3.050000 ;
      RECT  2.645000  1.925000  2.905000 2.085000 ;
      RECT  2.785000  0.640000  3.160000 0.970000 ;
      RECT  2.785000  0.970000  2.955000 1.565000 ;
      RECT  2.785000  1.565000  3.245000 1.735000 ;
      RECT  2.870000  2.765000  3.585000 3.050000 ;
      RECT  3.075000  1.735000  3.245000 2.425000 ;
      RECT  3.135000  1.140000  3.500000 1.385000 ;
      RECT  3.330000  0.470000  3.500000 1.140000 ;
      RECT  3.415000  1.555000  4.005000 1.750000 ;
      RECT  3.415000  1.920000  5.645000 2.065000 ;
      RECT  3.415000  2.065000  4.455000 2.220000 ;
      RECT  3.415000  2.220000  3.585000 2.765000 ;
      RECT  3.670000  0.640000  3.880000 1.145000 ;
      RECT  3.670000  1.145000  5.645000 1.325000 ;
      RECT  3.755000  2.720000  3.995000 3.245000 ;
      RECT  4.050000  0.470000  4.220000 0.805000 ;
      RECT  4.050000  0.805000  5.655000 0.975000 ;
      RECT  4.165000  2.220000  4.455000 3.050000 ;
      RECT  4.185000  1.845000  5.645000 1.920000 ;
      RECT  4.265000  1.495000  6.005000 1.675000 ;
      RECT  5.045000  0.085000  5.315000 0.635000 ;
      RECT  5.065000  2.735000  5.325000 3.245000 ;
      RECT  5.485000  0.255000  7.175000 0.425000 ;
      RECT  5.485000  0.425000  5.655000 0.805000 ;
      RECT  5.825000  0.595000  6.005000 1.495000 ;
      RECT  5.835000  1.675000  6.005000 2.405000 ;
      RECT  5.835000  2.405000  6.095000 2.735000 ;
      RECT  6.175000  0.425000  7.175000 0.435000 ;
      RECT  6.175000  0.435000  6.355000 2.075000 ;
      RECT  6.265000  2.405000  6.695000 2.735000 ;
      RECT  6.525000  0.605000  6.775000 1.055000 ;
      RECT  6.525000  1.055000  7.395000 1.225000 ;
      RECT  6.525000  1.225000  6.695000 2.405000 ;
      RECT  6.865000  1.455000  7.045000 2.125000 ;
      RECT  7.205000  2.775000  8.160000 3.245000 ;
      RECT  7.225000  1.225000  7.395000 1.325000 ;
      RECT  7.225000  1.325000  8.855000 1.495000 ;
      RECT  7.510000  0.085000  7.840000 0.885000 ;
      RECT  7.575000  2.185000  7.825000 2.435000 ;
      RECT  7.575000  2.435000  8.835000 2.605000 ;
      RECT  8.300000  0.670000  8.630000 0.985000 ;
      RECT  8.300000  0.985000  9.195000 1.155000 ;
      RECT  8.330000  2.605000  8.530000 3.050000 ;
      RECT  8.665000  2.175000  9.195000 2.345000 ;
      RECT  8.665000  2.345000  8.835000 2.435000 ;
      RECT  8.685000  1.495000  8.855000 1.995000 ;
      RECT  8.700000  2.775000  9.030000 3.245000 ;
      RECT  9.025000  1.155000  9.195000 2.175000 ;
      RECT  9.140000  0.255000  9.400000 0.645000 ;
      RECT  9.140000  0.645000  9.535000 0.815000 ;
      RECT  9.220000  2.515000  9.555000 3.075000 ;
      RECT  9.365000  0.815000  9.535000 1.185000 ;
      RECT  9.365000  1.185000 10.060000 1.515000 ;
      RECT  9.365000  1.515000  9.555000 2.515000 ;
      RECT  9.570000  0.085000 10.060000 0.475000 ;
      RECT  9.705000  0.475000 10.060000 1.015000 ;
      RECT  9.725000  1.815000 10.060000 3.245000 ;
      RECT 10.625000  0.085000 10.920000 1.095000 ;
      RECT 10.625000  1.815000 10.920000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  1.580000  1.765000 1.750000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  1.580000  3.685000 1.750000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  1.580000  7.045000 1.750000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
    LAYER met1 ;
      RECT 1.535000 1.550000 1.825000 1.595000 ;
      RECT 1.535000 1.595000 7.105000 1.735000 ;
      RECT 1.535000 1.735000 1.825000 1.780000 ;
      RECT 3.455000 1.550000 3.745000 1.595000 ;
      RECT 3.455000 1.735000 3.745000 1.780000 ;
      RECT 6.815000 1.550000 7.105000 1.595000 ;
      RECT 6.815000 1.735000 7.105000 1.780000 ;
  END
END sky130_fd_sc_lp__dfrtp_2
END LIBRARY
