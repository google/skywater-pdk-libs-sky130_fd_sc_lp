* File: sky130_fd_sc_lp__mux4_2.pex.spice
* Created: Wed Sep  2 10:01:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX4_2%A_80_293# 1 2 9 11 12 13 15 16 19 23 27 28
c61 28 0 4.91358e-20 $X=0.905 $Y=1.49
r62 23 27 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.73 $Y=2.17
+ $X2=1.73 $Y2=1.825
r63 20 28 42.1207 $w=5.55e-07 $l=4.85e-07 $layer=POLY_cond $X=1.39 $Y=1.49
+ $X2=0.905 $Y2=1.49
r64 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.39
+ $Y=1.32 $X2=1.39 $Y2=1.32
r65 17 27 8.3845 $w=5.98e-07 $l=3e-07 $layer=LI1_cond $X=1.595 $Y=1.525
+ $X2=1.595 $Y2=1.825
r66 17 19 4.0866 $w=5.98e-07 $l=2.05e-07 $layer=LI1_cond $X=1.595 $Y=1.525
+ $X2=1.595 $Y2=1.32
r67 16 26 3.66473 $w=5.16e-07 $l=2.10178e-07 $layer=LI1_cond $X=1.595 $Y=1.115
+ $X2=1.725 $Y2=0.96
r68 16 19 4.0866 $w=5.98e-07 $l=2.05e-07 $layer=LI1_cond $X=1.595 $Y=1.115
+ $X2=1.595 $Y2=1.32
r69 13 28 34.0645 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.905 $Y=1.155
+ $X2=0.905 $Y2=1.49
r70 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.905 $Y=1.155
+ $X2=0.905 $Y2=0.835
r71 11 28 35.559 $w=5.55e-07 $l=9.68246e-08 $layer=POLY_cond $X=0.83 $Y=1.54
+ $X2=0.905 $Y2=1.49
r72 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.54
+ $X2=0.55 $Y2=1.54
r73 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=1.615
+ $X2=0.55 $Y2=1.54
r74 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.475 $Y=1.615
+ $X2=0.475 $Y2=2.305
r75 2 23 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=2.025 $X2=1.73 $Y2=2.17
r76 1 26 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.655 $X2=1.99 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%S1 3 5 6 7 9 10 11 15 19 20 21 28 29
c78 29 0 7.78613e-20 $X=2.32 $Y=1.45
r79 27 29 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.16 $Y=1.45
+ $X2=2.32 $Y2=1.45
r80 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.45 $X2=2.16 $Y2=1.45
r81 24 27 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.04 $Y=1.45
+ $X2=2.16 $Y2=1.45
r82 20 21 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=2.035
r83 20 28 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=1.45
r84 17 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.285
+ $X2=2.32 $Y2=1.45
r85 17 19 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.32 $Y=1.285
+ $X2=2.32 $Y2=0.865
r86 16 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.32 $Y=0.255
+ $X2=2.32 $Y2=0.865
r87 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.04 $Y=2.735
+ $X2=2.04 $Y2=2.095
r88 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.615
+ $X2=2.04 $Y2=1.45
r89 12 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.04 $Y=1.615
+ $X2=2.04 $Y2=2.095
r90 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.965 $Y=2.81
+ $X2=2.04 $Y2=2.735
r91 10 11 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=1.965 $Y=2.81
+ $X2=0.98 $Y2=2.81
r92 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=2.735
+ $X2=0.98 $Y2=2.81
r93 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.905 $Y=2.735
+ $X2=0.905 $Y2=2.305
r94 5 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.245 $Y=0.18
+ $X2=2.32 $Y2=0.255
r95 5 6 869.138 $w=1.5e-07 $l=1.695e-06 $layer=POLY_cond $X=2.245 $Y=0.18
+ $X2=0.55 $Y2=0.18
r96 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=0.255
+ $X2=0.55 $Y2=0.18
r97 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.475 $Y=0.255
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%A_110_125# 1 2 9 11 13 16 18 20 23 27 28 29
+ 33 36 43
r92 43 44 5.95062 $w=3.24e-07 $l=4e-08 $layer=POLY_cond $X=3.335 $Y=1.352
+ $X2=3.375 $Y2=1.352
r93 42 43 58.0185 $w=3.24e-07 $l=3.9e-07 $layer=POLY_cond $X=2.945 $Y=1.352
+ $X2=3.335 $Y2=1.352
r94 41 42 5.95062 $w=3.24e-07 $l=4e-08 $layer=POLY_cond $X=2.905 $Y=1.352
+ $X2=2.945 $Y2=1.352
r95 36 38 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.55 $Y=0.41 $X2=1.55
+ $Y2=0.61
r96 34 41 20.0833 $w=3.24e-07 $l=1.35e-07 $layer=POLY_cond $X=2.77 $Y=1.352
+ $X2=2.905 $Y2=1.352
r97 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.35 $X2=2.77 $Y2=1.35
r98 31 33 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=2.73 $Y=0.695
+ $X2=2.73 $Y2=1.35
r99 30 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0.61
+ $X2=1.55 $Y2=0.61
r100 29 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.605 $Y=0.61
+ $X2=2.73 $Y2=0.695
r101 29 30 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=2.605 $Y=0.61
+ $X2=1.635 $Y2=0.61
r102 27 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=0.41
+ $X2=1.55 $Y2=0.41
r103 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.465 $Y=0.41
+ $X2=0.775 $Y2=0.41
r104 23 25 67.837 $w=2.18e-07 $l=1.295e-06 $layer=LI1_cond $X=0.665 $Y=0.835
+ $X2=0.665 $Y2=2.13
r105 21 28 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.665 $Y=0.495
+ $X2=0.775 $Y2=0.41
r106 21 23 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=0.665 $Y=0.495
+ $X2=0.665 $Y2=0.835
r107 18 44 20.7868 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=3.375 $Y=1.185
+ $X2=3.375 $Y2=1.352
r108 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.375 $Y=1.185
+ $X2=3.375 $Y2=0.655
r109 14 43 20.7868 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=3.335 $Y=1.52
+ $X2=3.335 $Y2=1.352
r110 14 16 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=3.335 $Y=1.52
+ $X2=3.335 $Y2=2.405
r111 11 42 20.7868 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=2.945 $Y=1.185
+ $X2=2.945 $Y2=1.352
r112 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.945 $Y=1.185
+ $X2=2.945 $Y2=0.655
r113 7 41 20.7868 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=2.905 $Y=1.52
+ $X2=2.905 $Y2=1.352
r114 7 9 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=2.905 $Y=1.52
+ $X2=2.905 $Y2=2.405
r115 2 25 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.985 $X2=0.69 $Y2=2.13
r116 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.625 $X2=0.69 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%A3 3 7 9 10 11 22
c40 22 0 1.49142e-19 $X=3.96 $Y=1.35
c41 7 0 5.31684e-20 $X=4.05 $Y=0.805
c42 3 0 2.41342e-21 $X=4.01 $Y=2.415
r43 22 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.96 $Y=1.35
+ $X2=3.96 $Y2=1.515
r44 22 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.96 $Y=1.35
+ $X2=3.96 $Y2=1.185
r45 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.96
+ $Y=1.35 $X2=3.96 $Y2=1.35
r46 10 11 5.98039 $w=7.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.795 $Y=1.665
+ $X2=3.795 $Y2=2.035
r47 10 23 5.09141 $w=7.38e-07 $l=3.15e-07 $layer=LI1_cond $X=3.795 $Y=1.665
+ $X2=3.795 $Y2=1.35
r48 9 23 0.888977 $w=7.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.795 $Y=1.295
+ $X2=3.795 $Y2=1.35
r49 7 24 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4.05 $Y=0.805
+ $X2=4.05 $Y2=1.185
r50 3 25 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=4.01 $Y=2.415 $X2=4.01
+ $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%A_859_351# 1 2 9 13 14 17 21 23 24 27 29 30
+ 31 34 35 36 39 43 45 49 53 55 56 59 61 63 64
c160 56 0 1.52601e-19 $X=6.907 $Y=0.985
c161 55 0 6.87706e-20 $X=6.907 $Y=1.07
c162 27 0 5.31684e-20 $X=6.83 $Y=0.805
c163 24 0 3.51732e-20 $X=6.475 $Y=1.46
c164 17 0 5.31684e-20 $X=4.84 $Y=0.805
c165 14 0 3.60778e-20 $X=4.485 $Y=1.46
r166 63 64 9.42615 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=8.227 $Y=2.24
+ $X2=8.227 $Y2=2.075
r167 59 72 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=6.85 $Y=1.315
+ $X2=6.85 $Y2=1.46
r168 59 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.85 $Y=1.315
+ $X2=6.85 $Y2=1.15
r169 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.315 $X2=6.85 $Y2=1.315
r170 55 58 6.34491 $w=4.43e-07 $l=2.45e-07 $layer=LI1_cond $X=6.907 $Y=1.07
+ $X2=6.907 $Y2=1.315
r171 55 56 6.78944 $w=4.43e-07 $l=8.5e-08 $layer=LI1_cond $X=6.907 $Y=1.07
+ $X2=6.907 $Y2=0.985
r172 53 68 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=4.86 $Y=1.315
+ $X2=4.86 $Y2=1.46
r173 53 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.86 $Y=1.315
+ $X2=4.86 $Y2=1.15
r174 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.86
+ $Y=1.315 $X2=4.86 $Y2=1.315
r175 49 52 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.86 $Y=1.08
+ $X2=4.86 $Y2=1.315
r176 47 64 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.385 $Y=1.155
+ $X2=8.385 $Y2=2.075
r177 46 61 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.11 $Y=1.07
+ $X2=7.98 $Y2=1.07
r178 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.3 $Y=1.07
+ $X2=8.385 $Y2=1.155
r179 45 46 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=8.3 $Y=1.07
+ $X2=8.11 $Y2=1.07
r180 41 61 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=0.985
+ $X2=7.98 $Y2=1.07
r181 41 43 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=7.98 $Y=0.985
+ $X2=7.98 $Y2=0.805
r182 40 55 6.43131 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=7.13 $Y=1.07
+ $X2=6.907 $Y2=1.07
r183 39 61 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.85 $Y=1.07
+ $X2=7.98 $Y2=1.07
r184 39 40 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.85 $Y=1.07
+ $X2=7.13 $Y2=1.07
r185 37 56 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.045 $Y=0.435
+ $X2=7.045 $Y2=0.985
r186 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.96 $Y=0.35
+ $X2=7.045 $Y2=0.435
r187 35 36 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=6.96 $Y=0.35
+ $X2=6.155 $Y2=0.35
r188 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.07 $Y=0.435
+ $X2=6.155 $Y2=0.35
r189 33 34 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.07 $Y=0.435
+ $X2=6.07 $Y2=0.995
r190 32 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=1.08
+ $X2=4.86 $Y2=1.08
r191 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.985 $Y=1.08
+ $X2=6.07 $Y2=0.995
r192 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.985 $Y=1.08
+ $X2=5.025 $Y2=1.08
r193 29 30 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=4.39 $Y=1.755
+ $X2=4.39 $Y2=1.905
r194 27 71 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.83 $Y=0.805
+ $X2=6.83 $Y2=1.15
r195 23 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.685 $Y=1.46
+ $X2=6.85 $Y2=1.46
r196 23 24 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.685 $Y=1.46
+ $X2=6.475 $Y2=1.46
r197 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.4 $Y=1.535
+ $X2=6.475 $Y2=1.46
r198 19 21 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=6.4 $Y=1.535
+ $X2=6.4 $Y2=2.415
r199 17 67 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.84 $Y=0.805
+ $X2=4.84 $Y2=1.15
r200 13 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.695 $Y=1.46
+ $X2=4.86 $Y2=1.46
r201 13 14 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.695 $Y=1.46
+ $X2=4.485 $Y2=1.46
r202 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.41 $Y=1.535
+ $X2=4.485 $Y2=1.46
r203 11 29 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=4.41 $Y=1.535
+ $X2=4.41 $Y2=1.755
r204 9 30 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.37 $Y=2.415
+ $X2=4.37 $Y2=1.905
r205 2 63 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.94
+ $Y=2.095 $X2=8.08 $Y2=2.24
r206 1 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.805
+ $Y=0.595 $X2=7.945 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%A2 1 3 7 9 10
r46 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.4
+ $Y=1.76 $X2=5.4 $Y2=1.76
r47 10 15 4.12815 $w=3.33e-07 $l=1.2e-07 $layer=LI1_cond $X=5.52 $Y=1.737
+ $X2=5.4 $Y2=1.737
r48 9 15 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=5.04 $Y=1.737 $X2=5.4
+ $Y2=1.737
r49 5 14 70.8721 $w=3.13e-07 $l=3.82426e-07 $layer=POLY_cond $X=5.31 $Y=1.385
+ $X2=5.325 $Y2=1.76
r50 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.31 $Y=1.385 $X2=5.31
+ $Y2=0.805
r51 1 14 38.5334 $w=3.13e-07 $l=2.33345e-07 $layer=POLY_cond $X=5.16 $Y=1.925
+ $X2=5.325 $Y2=1.76
r52 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=5.16 $Y=1.925 $X2=5.16
+ $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%A1 3 7 11 12 13 14 18 19
c45 3 0 1.8086e-19 $X=6.04 $Y=0.805
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.95
+ $Y=1.43 $X2=5.95 $Y2=1.43
r47 13 14 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=5.975 $Y=1.665
+ $X2=5.975 $Y2=2.035
r48 13 19 7.12695 $w=3.78e-07 $l=2.35e-07 $layer=LI1_cond $X=5.975 $Y=1.665
+ $X2=5.975 $Y2=1.43
r49 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.95 $Y=1.77
+ $X2=5.95 $Y2=1.43
r50 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.77
+ $X2=5.95 $Y2=1.935
r51 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.265
+ $X2=5.95 $Y2=1.43
r52 7 12 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.04 $Y=2.415
+ $X2=6.04 $Y2=1.935
r53 3 10 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=6.04 $Y=0.805
+ $X2=6.04 $Y2=1.265
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%A0 3 7 9 10 14
r36 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=1.77
+ $X2=7.39 $Y2=1.935
r37 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=1.77
+ $X2=7.39 $Y2=1.605
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.39
+ $Y=1.77 $X2=7.39 $Y2=1.77
r39 10 15 2.02183 $w=2.83e-07 $l=5e-08 $layer=LI1_cond $X=7.44 $Y=1.712 $X2=7.39
+ $Y2=1.712
r40 9 15 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=6.96 $Y=1.712
+ $X2=7.39 $Y2=1.712
r41 7 17 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.435 $Y=2.415
+ $X2=7.435 $Y2=1.935
r42 3 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=7.3 $Y=0.805 $X2=7.3
+ $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%S0 3 5 6 9 11 12 15 17 21 23 28 32 33 34 37
+ 39 40 43 44
c113 28 0 1.52601e-19 $X=7.73 $Y=0.805
r114 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.955
+ $Y=1.42 $X2=7.955 $Y2=1.42
r115 40 44 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=7.955 $Y=1.665
+ $X2=7.955 $Y2=1.42
r116 38 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.955 $Y=1.76
+ $X2=7.955 $Y2=1.42
r117 38 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.955 $Y=1.76
+ $X2=7.955 $Y2=1.925
r118 37 43 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=7.955 $Y=1.365
+ $X2=7.955 $Y2=1.42
r119 36 37 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=7.887 $Y=1.215
+ $X2=7.887 $Y2=1.365
r120 32 39 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=7.865 $Y=2.415
+ $X2=7.865 $Y2=1.925
r121 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.865 $Y=3.075
+ $X2=7.865 $Y2=2.415
r122 28 36 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.73 $Y=0.805
+ $X2=7.73 $Y2=1.215
r123 25 28 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.73 $Y=0.255
+ $X2=7.73 $Y2=0.805
r124 24 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7 $Y=3.15 $X2=6.925
+ $Y2=3.15
r125 23 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.79 $Y=3.15
+ $X2=7.865 $Y2=3.075
r126 23 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.79 $Y=3.15 $X2=7
+ $Y2=3.15
r127 19 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.925 $Y=3.075
+ $X2=6.925 $Y2=3.15
r128 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.925 $Y=3.075
+ $X2=6.925 $Y2=2.415
r129 18 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.475 $Y=0.18
+ $X2=6.4 $Y2=0.18
r130 17 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.655 $Y=0.18
+ $X2=7.73 $Y2=0.255
r131 17 18 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=7.655 $Y=0.18
+ $X2=6.475 $Y2=0.18
r132 13 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.4 $Y=0.255
+ $X2=6.4 $Y2=0.18
r133 13 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.4 $Y=0.255
+ $X2=6.4 $Y2=0.805
r134 11 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.85 $Y=3.15
+ $X2=6.925 $Y2=3.15
r135 11 12 1012.71 $w=1.5e-07 $l=1.975e-06 $layer=POLY_cond $X=6.85 $Y=3.15
+ $X2=4.875 $Y2=3.15
r136 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.8 $Y=3.075
+ $X2=4.875 $Y2=3.15
r137 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.8 $Y=3.075 $X2=4.8
+ $Y2=2.415
r138 5 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.325 $Y=0.18
+ $X2=6.4 $Y2=0.18
r139 5 6 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=6.325 $Y=0.18
+ $X2=4.485 $Y2=0.18
r140 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.41 $Y=0.255
+ $X2=4.485 $Y2=0.18
r141 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.41 $Y=0.255
+ $X2=4.41 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%A_27_125# 1 2 3 4 15 19 20 22 23 24 26 30 33
c98 30 0 3.60778e-20 $X=4.625 $Y=0.73
c99 26 0 1.49142e-19 $X=4.43 $Y=2.075
r100 33 34 8.78149 $w=3.89e-07 $l=2.8e-07 $layer=LI1_cond $X=4.547 $Y=2.24
+ $X2=4.547 $Y2=2.52
r101 27 30 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=4.43 $Y=0.695
+ $X2=4.625 $Y2=0.695
r102 26 33 9.10818 $w=3.89e-07 $l=2.15708e-07 $layer=LI1_cond $X=4.43 $Y=2.075
+ $X2=4.547 $Y2=2.24
r103 25 27 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.43 $Y=0.825
+ $X2=4.43 $Y2=0.695
r104 25 26 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.43 $Y=0.825
+ $X2=4.43 $Y2=2.075
r105 23 34 5.60925 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=4.345 $Y=2.52
+ $X2=4.547 $Y2=2.52
r106 23 24 176.802 $w=1.68e-07 $l=2.71e-06 $layer=LI1_cond $X=4.345 $Y=2.52
+ $X2=1.635 $Y2=2.52
r107 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.55 $Y=2.605
+ $X2=1.635 $Y2=2.52
r108 21 22 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.55 $Y=2.605
+ $X2=1.55 $Y2=2.815
r109 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.465 $Y=2.9
+ $X2=1.55 $Y2=2.815
r110 19 20 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=1.465 $Y=2.9
+ $X2=0.385 $Y2=2.9
r111 15 18 51.8599 $w=2.88e-07 $l=1.305e-06 $layer=LI1_cond $X=0.24 $Y=0.835
+ $X2=0.24 $Y2=2.14
r112 13 20 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=0.24 $Y=2.815
+ $X2=0.385 $Y2=2.9
r113 13 18 26.8241 $w=2.88e-07 $l=6.75e-07 $layer=LI1_cond $X=0.24 $Y=2.815
+ $X2=0.24 $Y2=2.14
r114 4 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.445
+ $Y=2.095 $X2=4.585 $Y2=2.24
r115 3 18 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.985 $X2=0.26 $Y2=2.14
r116 2 30 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=4.485
+ $Y=0.595 $X2=4.625 $Y2=0.73
r117 1 15 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.625 $X2=0.26 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%A_196_125# 1 2 3 4 20 24 25 29 31 32 35 38 44
+ 45
c105 32 0 4.91358e-20 $X=1.345 $Y=2.405
c106 29 0 3.51732e-20 $X=6.615 $Y=0.72
r107 44 45 9.08855 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=6.582 $Y=2.24
+ $X2=6.582 $Y2=2.075
r108 39 44 3.98693 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=6.582 $Y=2.405
+ $X2=6.582 $Y2=2.24
r109 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=2.405
+ $X2=6.48 $Y2=2.405
r110 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.405
+ $X2=1.2 $Y2=2.405
r111 32 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.405
+ $X2=1.2 $Y2=2.405
r112 31 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=2.405
+ $X2=6.48 $Y2=2.405
r113 31 32 6.17573 $w=1.4e-07 $l=4.99e-06 $layer=MET1_cond $X=6.335 $Y=2.405
+ $X2=1.345 $Y2=2.405
r114 26 29 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=6.425 $Y=0.71
+ $X2=6.615 $Y2=0.71
r115 24 25 7.45505 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.125 $Y=2.13
+ $X2=1.125 $Y2=1.995
r116 22 35 8.13489 $w=3.38e-07 $l=2.4e-07 $layer=LI1_cond $X=1.125 $Y=2.165
+ $X2=1.125 $Y2=2.405
r117 22 24 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=1.125 $Y=2.165
+ $X2=1.125 $Y2=2.13
r118 17 20 4.0085 $w=2.28e-07 $l=8e-08 $layer=LI1_cond $X=1.04 $Y=0.78 $X2=1.12
+ $Y2=0.78
r119 15 26 1.64051 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=6.425 $Y=0.815
+ $X2=6.425 $Y2=0.71
r120 15 45 77.6364 $w=1.78e-07 $l=1.26e-06 $layer=LI1_cond $X=6.425 $Y=0.815
+ $X2=6.425 $Y2=2.075
r121 13 17 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.04 $Y=0.895
+ $X2=1.04 $Y2=0.78
r122 13 25 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=1.04 $Y=0.895
+ $X2=1.04 $Y2=1.995
r123 4 44 300 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=2 $X=6.475
+ $Y=2.095 $X2=6.665 $Y2=2.24
r124 3 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.985 $X2=1.12 $Y2=2.13
r125 2 29 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=6.475
+ $Y=0.595 $X2=6.615 $Y2=0.72
r126 1 20 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.625 $X2=1.12 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%VPWR 1 2 3 4 15 19 21 22 25 32 33 34 36 44 49
+ 65 66 69 72 75
r97 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r98 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r99 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r101 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r102 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r103 60 63 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r104 60 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r105 59 62 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.44
+ $Y2=3.33
r106 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r107 57 75 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=5.99 $Y=3.33 $X2=5.6
+ $Y2=3.33
r108 57 59 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.99 $Y=3.33 $X2=6
+ $Y2=3.33
r109 56 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r111 53 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r112 52 55 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r113 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 50 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=3.55 $Y2=3.33
r115 50 52 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=4.08 $Y2=3.33
r116 49 75 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=5.21 $Y=3.33 $X2=5.6
+ $Y2=3.33
r117 49 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.04 $Y2=3.33
r118 48 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r119 48 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r121 45 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.69 $Y2=3.33
r122 45 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.12 $Y2=3.33
r123 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.55 $Y2=3.33
r124 44 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 43 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r126 42 43 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r127 39 43 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r128 38 42 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 38 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r130 36 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.69 $Y2=3.33
r131 36 42 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.16 $Y2=3.33
r132 34 56 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=5.04 $Y2=3.33
r133 34 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 32 62 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.44 $Y2=3.33
r135 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.65 $Y2=3.33
r136 31 65 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=7.815 $Y=3.33
+ $X2=8.4 $Y2=3.33
r137 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=3.33
+ $X2=7.65 $Y2=3.33
r138 28 30 6.69032 $w=6.2e-07 $l=4.38292e-07 $layer=LI1_cond $X=5.375 $Y=2.25
+ $X2=5.6 $Y2=2.59
r139 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.65 $Y=3.245
+ $X2=7.65 $Y2=3.33
r140 23 25 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=7.65 $Y=3.245
+ $X2=7.65 $Y2=2.25
r141 22 75 3.08259 $w=7.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.6 $Y=3.245 $X2=5.6
+ $Y2=3.33
r142 21 30 1.9557 $w=7.8e-07 $l=9e-08 $layer=LI1_cond $X=5.6 $Y=2.68 $X2=5.6
+ $Y2=2.59
r143 21 22 8.6639 $w=7.78e-07 $l=5.65e-07 $layer=LI1_cond $X=5.6 $Y=2.68 $X2=5.6
+ $Y2=3.245
r144 17 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.55 $Y2=3.33
r145 17 19 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.55 $Y2=2.89
r146 13 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=3.245
+ $X2=2.69 $Y2=3.33
r147 13 15 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.69 $Y=3.245
+ $X2=2.69 $Y2=2.89
r148 4 25 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=7.51
+ $Y=2.095 $X2=7.65 $Y2=2.25
r149 3 30 400 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=2.095 $X2=5.375 $Y2=2.59
r150 3 28 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=2.095 $X2=5.375 $Y2=2.25
r151 2 19 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.775 $X2=3.55 $Y2=2.89
r152 1 15 600 $w=1.7e-07 $l=1.37272e-06 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.775 $X2=2.69 $Y2=2.89
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%X 1 2 7 8 9 10 11 18
c17 18 0 8.02747e-20 $X=3.16 $Y=0.42
r18 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=1.665
+ $X2=3.14 $Y2=2.035
r19 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=1.295
+ $X2=3.14 $Y2=1.665
r20 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=0.925 $X2=3.14
+ $Y2=1.295
r21 7 8 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=0.555 $X2=3.14
+ $Y2=0.925
r22 7 18 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.14 $Y=0.555
+ $X2=3.14 $Y2=0.42
r23 2 11 600 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_PDIFF $count=1 $X=2.98
+ $Y=1.775 $X2=3.12 $Y2=2.1
r24 1 18 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.02
+ $Y=0.235 $X2=3.16 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_2%VGND 1 2 3 4 15 21 25 27 29 37 42 47 57 58 62
+ 68 71 74
c82 58 0 1.27692e-19 $X=8.4 $Y=0
r83 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r84 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r85 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r86 62 65 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.65 $Y=0 $X2=2.65
+ $Y2=0.26
r87 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r88 58 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r89 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r90 55 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.68 $Y=0 $X2=7.515
+ $Y2=0
r91 55 57 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.68 $Y=0 $X2=8.4
+ $Y2=0
r92 54 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r93 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r94 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r95 51 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r96 50 53 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=0 $X2=6.96 $Y2=0
r97 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r98 48 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=0 $X2=5.65
+ $Y2=0
r99 48 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.815 $Y=0 $X2=6
+ $Y2=0
r100 47 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.35 $Y=0 $X2=7.515
+ $Y2=0
r101 47 53 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.35 $Y=0 $X2=6.96
+ $Y2=0
r102 46 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r103 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r104 43 68 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.72
+ $Y2=0
r105 43 45 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.08
+ $Y2=0
r106 42 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.485 $Y=0 $X2=5.65
+ $Y2=0
r107 42 45 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=5.485 $Y=0
+ $X2=4.08 $Y2=0
r108 41 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r109 41 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r110 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r111 38 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.65
+ $Y2=0
r112 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.815 $Y=0
+ $X2=3.12 $Y2=0
r113 37 68 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.72
+ $Y2=0
r114 37 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=0
+ $X2=3.12 $Y2=0
r115 36 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r116 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r117 32 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=2.16 $Y2=0
r118 31 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r119 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r120 29 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.485 $Y=0 $X2=2.65
+ $Y2=0
r121 29 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.485 $Y=0
+ $X2=2.16 $Y2=0
r122 27 72 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=5.52
+ $Y2=0
r123 27 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r124 23 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.515 $Y=0.085
+ $X2=7.515 $Y2=0
r125 23 25 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=7.515 $Y=0.085
+ $X2=7.515 $Y2=0.72
r126 19 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.65 $Y=0.085
+ $X2=5.65 $Y2=0
r127 19 21 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.65 $Y=0.085
+ $X2=5.65 $Y2=0.72
r128 15 17 8.71718 $w=5.88e-07 $l=4.3e-07 $layer=LI1_cond $X=3.72 $Y=0.38
+ $X2=3.72 $Y2=0.81
r129 13 68 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0
r130 13 15 5.98039 $w=5.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0.38
r131 4 25 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=7.375
+ $Y=0.595 $X2=7.515 $Y2=0.72
r132 3 21 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=5.385
+ $Y=0.595 $X2=5.65 $Y2=0.72
r133 2 17 182 $w=1.7e-07 $l=7.42967e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.235 $X2=3.835 $Y2=0.81
r134 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.235 $X2=3.59 $Y2=0.38
r135 1 65 182 $w=1.7e-07 $l=5.06705e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.655 $X2=2.65 $Y2=0.26
.ends

