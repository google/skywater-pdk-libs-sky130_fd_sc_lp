* File: sky130_fd_sc_lp__dlxbp_1.pex.spice
* Created: Fri Aug 28 10:28:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXBP_1%D 3 6 9 10 11 12 13 17
c35 11 0 6.60299e-20 $X=0.55 $Y=1.51
c36 10 0 1.78633e-19 $X=0.55 $Y=1.345
c37 6 0 1.26821e-19 $X=0.64 $Y=2.415
r38 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.55
+ $Y=1.005 $X2=0.55 $Y2=1.005
r39 13 18 7.54049 $w=4.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.685 $Y=1.295
+ $X2=0.685 $Y2=1.005
r40 12 18 2.08014 $w=4.58e-07 $l=8e-08 $layer=LI1_cond $X=0.685 $Y=0.925
+ $X2=0.685 $Y2=1.005
r41 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.55 $Y=1.345
+ $X2=0.55 $Y2=1.005
r42 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.345
+ $X2=0.55 $Y2=1.51
r43 9 17 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=0.84
+ $X2=0.55 $Y2=1.005
r44 6 11 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=0.64 $Y=2.415
+ $X2=0.64 $Y2=1.51
r45 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.57 $Y=0.52 $X2=0.57
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%GATE 3 7 9 11 13 14 18
c46 9 0 2.01481e-20 $X=1.45 $Y=0.935
r47 13 14 19.7562 $w=2.43e-07 $l=4.2e-07 $layer=LI1_cond $X=1.652 $Y=0.505
+ $X2=1.652 $Y2=0.925
r48 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.615
+ $Y=0.505 $X2=1.615 $Y2=0.505
r49 12 18 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.615 $Y=0.86
+ $X2=1.615 $Y2=0.505
r50 10 11 5.30422 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.145 $Y=0.935
+ $X2=1.035 $Y2=0.935
r51 9 12 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.45 $Y=0.935
+ $X2=1.615 $Y2=0.86
r52 9 10 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.45 $Y=0.935
+ $X2=1.145 $Y2=0.935
r53 5 11 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.07 $Y=1.01
+ $X2=1.035 $Y2=0.935
r54 5 7 720.436 $w=1.5e-07 $l=1.405e-06 $layer=POLY_cond $X=1.07 $Y=1.01
+ $X2=1.07 $Y2=2.415
r55 1 11 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1 $Y=0.86
+ $X2=1.035 $Y2=0.935
r56 1 3 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1 $Y=0.86 $X2=1
+ $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%A_215_62# 1 2 8 9 11 14 18 20 24 28 32 36 37
+ 38 40 42 43 45 47 48 59
c128 47 0 1.66412e-19 $X=2.155 $Y=1.25
c129 42 0 9.58719e-20 $X=3.015 $Y=1.535
c130 37 0 3.05454e-19 $X=1.36 $Y=1.41
c131 24 0 1.79722e-19 $X=3.665 $Y=0.445
r132 55 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.53
+ $X2=3.055 $Y2=1.695
r133 55 59 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.055 $Y=1.53
+ $X2=3.055 $Y2=1.44
r134 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.055
+ $Y=1.53 $X2=3.055 $Y2=1.53
r135 50 51 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=2.155 $Y=1.41
+ $X2=2.155 $Y2=1.45
r136 48 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.25
+ $X2=2.155 $Y2=1.415
r137 48 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.25
+ $X2=2.155 $Y2=1.085
r138 47 50 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.155 $Y=1.25
+ $X2=2.155 $Y2=1.41
r139 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.155
+ $Y=1.25 $X2=2.155 $Y2=1.25
r140 42 54 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=1.535
+ $X2=3.015 $Y2=1.45
r141 42 43 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=3.015 $Y=1.535
+ $X2=3.015 $Y2=2.075
r142 41 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=1.45
+ $X2=2.155 $Y2=1.45
r143 40 54 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.89 $Y=1.45
+ $X2=3.015 $Y2=1.45
r144 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.89 $Y=1.45
+ $X2=2.32 $Y2=1.45
r145 39 45 4.57023 $w=1.8e-07 $l=1.48e-07 $layer=LI1_cond $X=1.45 $Y=2.165
+ $X2=1.302 $Y2=2.165
r146 38 43 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=2.89 $Y=2.165
+ $X2=3.015 $Y2=2.075
r147 38 39 88.7273 $w=1.78e-07 $l=1.44e-06 $layer=LI1_cond $X=2.89 $Y=2.165
+ $X2=1.45 $Y2=2.165
r148 36 50 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=1.41
+ $X2=2.155 $Y2=1.41
r149 36 37 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=1.99 $Y=1.41
+ $X2=1.36 $Y2=1.41
r150 30 37 6.83662 $w=2.5e-07 $l=1.9051e-07 $layer=LI1_cond $X=1.222 $Y=1.285
+ $X2=1.36 $Y2=1.41
r151 30 32 31.6398 $w=2.73e-07 $l=7.55e-07 $layer=LI1_cond $X=1.222 $Y=1.285
+ $X2=1.222 $Y2=0.53
r152 26 28 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=2.065 $Y=2.27
+ $X2=2.175 $Y2=2.27
r153 22 24 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=3.665 $Y=1.365
+ $X2=3.665 $Y2=0.445
r154 21 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.44
+ $X2=3.055 $Y2=1.44
r155 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.59 $Y=1.44
+ $X2=3.665 $Y2=1.365
r156 20 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.59 $Y=1.44
+ $X2=3.22 $Y2=1.44
r157 18 62 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=2.965 $Y=2.775
+ $X2=2.965 $Y2=1.695
r158 14 57 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.245 $Y=0.445
+ $X2=2.245 $Y2=1.085
r159 9 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.175 $Y=2.345
+ $X2=2.175 $Y2=2.27
r160 9 11 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.175 $Y=2.345
+ $X2=2.175 $Y2=2.775
r161 8 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.065 $Y=2.195
+ $X2=2.065 $Y2=2.27
r162 8 58 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.065 $Y=2.195
+ $X2=2.065 $Y2=1.415
r163 2 45 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=2.095 $X2=1.285 $Y2=2.24
r164 1 32 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.31 $X2=1.215 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%A_46_62# 1 2 11 15 19 22 25 29 30 35 37 39
c76 39 0 1.66412e-19 $X=2.515 $Y=1.655
c77 29 0 6.60299e-20 $X=2.515 $Y=1.82
r78 32 35 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.185 $Y=0.505
+ $X2=0.355 $Y2=0.505
r79 30 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.82
+ $X2=2.515 $Y2=1.985
r80 30 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.82
+ $X2=2.515 $Y2=1.655
r81 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.515
+ $Y=1.82 $X2=2.515 $Y2=1.82
r82 27 37 2.12 $w=2e-07 $l=2.35e-07 $layer=LI1_cond $X=0.555 $Y=1.805 $X2=0.32
+ $Y2=1.805
r83 27 29 108.691 $w=1.98e-07 $l=1.96e-06 $layer=LI1_cond $X=0.555 $Y=1.805
+ $X2=2.515 $Y2=1.805
r84 23 37 4.31155 $w=2.47e-07 $l=1.36748e-07 $layer=LI1_cond $X=0.407 $Y=1.905
+ $X2=0.32 $Y2=1.805
r85 23 25 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=0.407 $Y=1.905
+ $X2=0.407 $Y2=2.24
r86 22 37 4.31155 $w=2.47e-07 $l=1.78115e-07 $layer=LI1_cond $X=0.185 $Y=1.705
+ $X2=0.32 $Y2=1.805
r87 21 32 3.66692 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.185 $Y=0.67
+ $X2=0.185 $Y2=0.505
r88 21 22 57.3955 $w=1.98e-07 $l=1.035e-06 $layer=LI1_cond $X=0.185 $Y=0.67
+ $X2=0.185 $Y2=1.705
r89 17 19 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.605 $Y=1.05
+ $X2=2.765 $Y2=1.05
r90 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.765 $Y=0.975
+ $X2=2.765 $Y2=1.05
r91 13 15 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.765 $Y=0.975
+ $X2=2.765 $Y2=0.445
r92 11 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.605 $Y=2.775
+ $X2=2.605 $Y2=1.985
r93 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.605 $Y=1.125
+ $X2=2.605 $Y2=1.05
r94 7 39 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.605 $Y=1.125
+ $X2=2.605 $Y2=1.655
r95 2 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.3
+ $Y=2.095 $X2=0.425 $Y2=2.24
r96 1 35 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.23
+ $Y=0.31 $X2=0.355 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%A_367_491# 1 2 9 12 16 20 22 23 24 25 29 30
+ 32 33 36
c104 33 0 4.177e-19 $X=3.215 $Y=0.93
c105 22 0 1.59457e-19 $X=3.31 $Y=2.51
r106 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=0.93
+ $X2=3.215 $Y2=0.765
r107 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.215
+ $Y=0.93 $X2=3.215 $Y2=0.93
r108 30 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=2.13
+ $X2=3.415 $Y2=2.295
r109 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=2.13 $X2=3.415 $Y2=2.13
r110 27 29 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=3.41 $Y=2.425
+ $X2=3.41 $Y2=2.13
r111 26 32 7.3882 $w=3.22e-07 $l=3.02159e-07 $layer=LI1_cond $X=3.41 $Y=1.185
+ $X2=3.215 $Y2=0.965
r112 26 29 52.4045 $w=1.98e-07 $l=9.45e-07 $layer=LI1_cond $X=3.41 $Y=1.185
+ $X2=3.41 $Y2=2.13
r113 24 32 8.95589 $w=3.22e-07 $l=2.22486e-07 $layer=LI1_cond $X=3.05 $Y=0.83
+ $X2=3.215 $Y2=0.965
r114 24 25 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.05 $Y=0.83
+ $X2=2.135 $Y2=0.83
r115 22 27 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.31 $Y=2.51
+ $X2=3.41 $Y2=2.425
r116 22 23 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=3.31 $Y=2.51
+ $X2=2.125 $Y2=2.51
r117 18 25 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.04 $Y=0.745
+ $X2=2.135 $Y2=0.83
r118 18 20 17.512 $w=1.88e-07 $l=3e-07 $layer=LI1_cond $X=2.04 $Y=0.745 $X2=2.04
+ $Y2=0.445
r119 14 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.96 $Y=2.595
+ $X2=2.125 $Y2=2.51
r120 14 16 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.96 $Y=2.595
+ $X2=1.96 $Y2=2.6
r121 12 40 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.49 $Y=2.665
+ $X2=3.49 $Y2=2.295
r122 9 36 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.125 $Y=0.445
+ $X2=3.125 $Y2=0.765
r123 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.835
+ $Y=2.455 $X2=1.96 $Y2=2.6
r124 1 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.03 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%A_758_359# 1 2 9 13 15 17 19 22 24 26 28 31
+ 35 36 38 39 42 43 45 46 49 53 56 58 59 61 66 70
c129 42 0 3.5799e-19 $X=4.115 $Y=1.48
c130 9 0 1.59457e-19 $X=3.865 $Y=2.665
r131 67 70 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.23 $Y=1.43 $X2=5.23
+ $Y2=1.34
r132 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.23
+ $Y=1.43 $X2=5.23 $Y2=1.43
r133 64 66 6.39082 $w=3.28e-07 $l=1.83e-07 $layer=LI1_cond $X=5.047 $Y=1.43
+ $X2=5.23 $Y2=1.43
r134 62 64 0.942908 $w=3.28e-07 $l=2.7e-08 $layer=LI1_cond $X=5.02 $Y=1.43
+ $X2=5.047 $Y2=1.43
r135 58 61 3.80849 $w=2.42e-07 $l=9.31128e-08 $layer=LI1_cond $X=5.047 $Y=1.775
+ $X2=5.03 $Y2=1.86
r136 57 64 2.99809 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=5.047 $Y=1.595
+ $X2=5.047 $Y2=1.43
r137 57 58 9.21954 $w=2.23e-07 $l=1.8e-07 $layer=LI1_cond $X=5.047 $Y=1.595
+ $X2=5.047 $Y2=1.775
r138 56 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.02 $Y=1.265
+ $X2=5.02 $Y2=1.43
r139 56 59 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.02 $Y=1.265
+ $X2=5.02 $Y2=1.005
r140 51 61 3.80849 $w=2.42e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=1.945
+ $X2=5.03 $Y2=1.86
r141 51 53 41.8869 $w=2.58e-07 $l=9.45e-07 $layer=LI1_cond $X=5.03 $Y=1.945
+ $X2=5.03 $Y2=2.89
r142 47 59 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=4.912 $Y=0.813
+ $X2=4.912 $Y2=1.005
r143 47 49 11.7639 $w=3.83e-07 $l=3.93e-07 $layer=LI1_cond $X=4.912 $Y=0.813
+ $X2=4.912 $Y2=0.42
r144 45 61 2.64776 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.9 $Y=1.86 $X2=5.03
+ $Y2=1.86
r145 45 46 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.9 $Y=1.86 $X2=4.21
+ $Y2=1.86
r146 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.115
+ $Y=1.48 $X2=4.115 $Y2=1.48
r147 40 46 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.115 $Y=1.775
+ $X2=4.21 $Y2=1.86
r148 40 42 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=4.115 $Y=1.775
+ $X2=4.115 $Y2=1.48
r149 36 43 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.115 $Y=1.44
+ $X2=4.115 $Y2=1.48
r150 36 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.115 $Y=1.44
+ $X2=4.115 $Y2=1.275
r151 34 43 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=4.115 $Y=1.795
+ $X2=4.115 $Y2=1.48
r152 34 35 50.583 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.035 $Y=1.795
+ $X2=4.035 $Y2=1.985
r153 29 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.255 $Y=1.415
+ $X2=6.255 $Y2=1.34
r154 29 31 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.255 $Y=1.415
+ $X2=6.255 $Y2=2.155
r155 26 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.255 $Y=1.265
+ $X2=6.255 $Y2=1.34
r156 26 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.255 $Y=1.265
+ $X2=6.255 $Y2=0.945
r157 25 38 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.805 $Y=1.34 $X2=5.73
+ $Y2=1.34
r158 24 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.18 $Y=1.34
+ $X2=6.255 $Y2=1.34
r159 24 25 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=6.18 $Y=1.34
+ $X2=5.805 $Y2=1.34
r160 20 38 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.73 $Y=1.415 $X2=5.73
+ $Y2=1.34
r161 20 22 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=5.73 $Y=1.415
+ $X2=5.73 $Y2=2.465
r162 17 38 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.73 $Y=1.265 $X2=5.73
+ $Y2=1.34
r163 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.73 $Y=1.265
+ $X2=5.73 $Y2=0.735
r164 16 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.34
+ $X2=5.23 $Y2=1.34
r165 15 38 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.655 $Y=1.34 $X2=5.73
+ $Y2=1.34
r166 15 16 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.655 $Y=1.34
+ $X2=5.395 $Y2=1.34
r167 13 37 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.025 $Y=0.445
+ $X2=4.025 $Y2=1.275
r168 9 35 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.865 $Y=2.665
+ $X2=3.865 $Y2=1.985
r169 2 61 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.775 $X2=4.995 $Y2=1.94
r170 2 53 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.775 $X2=4.995 $Y2=2.89
r171 1 49 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=4.655
+ $Y=0.235 $X2=4.815 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%A_608_491# 1 2 7 9 12 14 19 21 22 25 27 35
c89 35 0 2.06947e-19 $X=4.78 $Y=1.35
c90 27 0 1.93528e-19 $X=3.765 $Y=1.06
r91 31 35 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.67 $Y=1.35
+ $X2=4.78 $Y2=1.35
r92 31 32 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.67 $Y=1.35 $X2=4.58
+ $Y2=1.35
r93 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.67
+ $Y=1.35 $X2=4.67 $Y2=1.35
r94 23 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=1.06
+ $X2=3.765 $Y2=1.06
r95 22 30 11.9932 $w=2.95e-07 $l=3.71927e-07 $layer=LI1_cond $X=4.38 $Y=1.06
+ $X2=4.567 $Y2=1.35
r96 22 23 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.38 $Y=1.06
+ $X2=3.85 $Y2=1.06
r97 20 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=1.145
+ $X2=3.765 $Y2=1.06
r98 20 21 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=3.765 $Y=1.145
+ $X2=3.765 $Y2=2.765
r99 19 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=0.975
+ $X2=3.765 $Y2=1.06
r100 18 25 13.9058 $w=3.29e-07 $l=4.95606e-07 $layer=LI1_cond $X=3.765 $Y=0.835
+ $X2=3.39 $Y2=0.555
r101 18 19 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.765 $Y=0.835
+ $X2=3.765 $Y2=0.975
r102 14 21 7.59919 $w=3.1e-07 $l=1.92873e-07 $layer=LI1_cond $X=3.68 $Y=2.92
+ $X2=3.765 $Y2=2.765
r103 14 16 18.5878 $w=3.08e-07 $l=5e-07 $layer=LI1_cond $X=3.68 $Y=2.92 $X2=3.18
+ $Y2=2.92
r104 10 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.78 $Y=1.515
+ $X2=4.78 $Y2=1.35
r105 10 12 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=4.78 $Y=1.515
+ $X2=4.78 $Y2=2.405
r106 7 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.58 $Y=1.185
+ $X2=4.58 $Y2=1.35
r107 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.58 $Y=1.185
+ $X2=4.58 $Y2=0.655
r108 2 16 600 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.455 $X2=3.18 $Y2=2.89
r109 1 25 182 $w=1.7e-07 $l=2.63344e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.235 $X2=3.39 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%A_1266_147# 1 2 9 12 16 20 24 25 27 29
c39 27 0 9.24665e-20 $X=6.47 $Y=1.51
r40 25 30 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.092 $Y=1.51
+ $X2=7.092 $Y2=1.675
r41 25 29 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.092 $Y=1.51
+ $X2=7.092 $Y2=1.345
r42 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.07
+ $Y=1.51 $X2=7.07 $Y2=1.51
r43 22 27 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.635 $Y=1.51
+ $X2=6.47 $Y2=1.51
r44 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.635 $Y=1.51
+ $X2=7.07 $Y2=1.51
r45 18 27 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.47 $Y=1.675
+ $X2=6.47 $Y2=1.51
r46 18 20 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.47 $Y=1.675
+ $X2=6.47 $Y2=1.98
r47 14 27 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.47 $Y=1.345
+ $X2=6.47 $Y2=1.51
r48 14 16 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.47 $Y=1.345
+ $X2=6.47 $Y2=0.955
r49 12 30 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.205 $Y=2.465
+ $X2=7.205 $Y2=1.675
r50 9 29 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.205 $Y=0.815
+ $X2=7.205 $Y2=1.345
r51 2 20 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.33
+ $Y=1.835 $X2=6.47 $Y2=1.98
r52 1 16 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.735 $X2=6.47 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%VPWR 1 2 3 4 5 18 22 24 27 30 36 41 42 44 45
+ 50 62 66 71 78 79 82 87 90
r98 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r99 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r100 83 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r101 82 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r102 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 79 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r104 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r105 76 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.155 $Y=3.33
+ $X2=6.99 $Y2=3.33
r106 76 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.155 $Y=3.33
+ $X2=7.44 $Y2=3.33
r107 75 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r108 75 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r109 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 72 87 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=5.985 $Y2=3.33
r111 72 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 71 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.99 $Y2=3.33
r113 71 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 70 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r115 70 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r117 67 82 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=4.375 $Y2=3.33
r118 67 69 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 66 87 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.985 $Y2=3.33
r120 66 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 62 82 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=4.375 $Y2=3.33
r123 62 64 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=2.64 $Y2=3.33
r124 61 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r125 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r127 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r128 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 54 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 50 85 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 50 65 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 47 49 7.46043 $w=5.56e-07 $l=4.245e-07 $layer=LI1_cond $X=4.565 $Y=2.21
+ $X2=4.375 $Y2=2.55
r134 44 60 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.16 $Y2=3.33
r135 44 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.425 $Y2=3.33
r136 43 64 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.64 $Y2=3.33
r137 43 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.425 $Y2=3.33
r138 41 53 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r139 41 42 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.855 $Y2=3.33
r140 40 57 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.2 $Y2=3.33
r141 40 42 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.855 $Y2=3.33
r142 36 39 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=6.99 $Y=1.98
+ $X2=6.99 $Y2=2.95
r143 34 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=3.245
+ $X2=6.99 $Y2=3.33
r144 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.99 $Y=3.245
+ $X2=6.99 $Y2=2.95
r145 30 33 18.0549 $w=2.98e-07 $l=4.7e-07 $layer=LI1_cond $X=5.985 $Y=1.98
+ $X2=5.985 $Y2=2.45
r146 28 87 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=3.33
r147 28 33 30.5397 $w=2.98e-07 $l=7.95e-07 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=2.45
r148 25 82 2.89202 $w=7.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=3.245
+ $X2=4.375 $Y2=3.33
r149 25 27 5.98039 $w=7.08e-07 $l=3.55e-07 $layer=LI1_cond $X=4.375 $Y=3.245
+ $X2=4.375 $Y2=2.89
r150 24 49 3.35657 $w=7.1e-07 $l=1.6e-07 $layer=LI1_cond $X=4.375 $Y=2.71
+ $X2=4.375 $Y2=2.55
r151 24 27 3.03231 $w=7.08e-07 $l=1.8e-07 $layer=LI1_cond $X=4.375 $Y=2.71
+ $X2=4.375 $Y2=2.89
r152 20 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=3.245
+ $X2=2.425 $Y2=3.33
r153 20 22 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.425 $Y=3.245
+ $X2=2.425 $Y2=2.93
r154 16 42 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=3.245
+ $X2=0.855 $Y2=3.33
r155 16 18 44.5464 $w=2.58e-07 $l=1.005e-06 $layer=LI1_cond $X=0.855 $Y=3.245
+ $X2=0.855 $Y2=2.24
r156 5 39 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=6.865
+ $Y=1.835 $X2=6.99 $Y2=2.95
r157 5 36 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.865
+ $Y=1.835 $X2=6.99 $Y2=1.98
r158 4 33 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=5.805
+ $Y=1.835 $X2=5.945 $Y2=2.45
r159 4 30 600 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.835 $X2=5.995 $Y2=1.98
r160 3 49 400 $w=1.7e-07 $l=6.7082e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=2.455 $X2=4.565 $Y2=2.55
r161 3 47 600 $w=1.7e-07 $l=7.37394e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=2.455 $X2=4.565 $Y2=2.21
r162 3 27 400 $w=1.7e-07 $l=8.13941e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=2.455 $X2=4.565 $Y2=2.89
r163 2 22 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=2.455 $X2=2.39 $Y2=2.93
r164 1 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.715
+ $Y=2.095 $X2=0.855 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%Q 1 2 7 9 15 16 17 28
c40 15 0 2.86787e-20 $X=5.507 $Y=1.815
r41 21 28 0.475611 $w=3.13e-07 $l=1.3e-08 $layer=LI1_cond $X=5.507 $Y=0.938
+ $X2=5.507 $Y2=0.925
r42 17 30 6.85281 $w=3.13e-07 $l=1.21e-07 $layer=LI1_cond $X=5.507 $Y=0.974
+ $X2=5.507 $Y2=1.095
r43 17 21 1.31708 $w=3.13e-07 $l=3.6e-08 $layer=LI1_cond $X=5.507 $Y=0.974
+ $X2=5.507 $Y2=0.938
r44 17 28 1.31708 $w=3.13e-07 $l=3.6e-08 $layer=LI1_cond $X=5.507 $Y=0.889
+ $X2=5.507 $Y2=0.925
r45 16 17 14.0488 $w=3.13e-07 $l=3.84e-07 $layer=LI1_cond $X=5.507 $Y=0.505
+ $X2=5.507 $Y2=0.889
r46 15 30 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.58 $Y=1.815
+ $X2=5.58 $Y2=1.095
r47 9 11 34.0245 $w=3.13e-07 $l=9.3e-07 $layer=LI1_cond $X=5.507 $Y=1.98
+ $X2=5.507 $Y2=2.91
r48 7 15 8.16989 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=5.507 $Y=1.972
+ $X2=5.507 $Y2=1.815
r49 7 9 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=5.507 $Y=1.972
+ $X2=5.507 $Y2=1.98
r50 2 11 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=1.835 $X2=5.515 $Y2=2.91
r51 2 9 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=1.835 $X2=5.515 $Y2=1.98
r52 1 16 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=5.39
+ $Y=0.315 $X2=5.515 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%Q_N 1 2 7 8 9 10 11 12 13
r10 13 39 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.46 $Y=2.775
+ $X2=7.46 $Y2=2.91
r11 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.46 $Y=2.405
+ $X2=7.46 $Y2=2.775
r12 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.46 $Y=1.98
+ $X2=7.46 $Y2=2.405
r13 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.46 $Y=1.665
+ $X2=7.46 $Y2=1.98
r14 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.46 $Y=1.295
+ $X2=7.46 $Y2=1.665
r15 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.46 $Y=0.925 $X2=7.46
+ $Y2=1.295
r16 7 8 16.433 $w=2.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.46 $Y=0.54 $X2=7.46
+ $Y2=0.925
r17 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.835 $X2=7.42 $Y2=2.91
r18 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.835 $X2=7.42 $Y2=1.98
r19 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.28
+ $Y=0.395 $X2=7.42 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_1%VGND 1 2 3 4 5 20 24 26 30 34 40 42 44 52 60
+ 67 68 71 74 77 80 83
c95 68 0 2.01481e-20 $X=7.44 $Y=0
c96 26 0 1.28299e-19 $X=4.075 $Y=0
r97 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r98 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r99 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r100 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r101 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r102 68 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r103 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r104 65 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.155 $Y=0 $X2=6.99
+ $Y2=0
r105 65 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.155 $Y=0
+ $X2=7.44 $Y2=0
r106 64 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r107 64 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r108 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r109 61 80 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.135 $Y=0 $X2=5.985
+ $Y2=0
r110 61 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.135 $Y=0 $X2=6.48
+ $Y2=0
r111 60 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=0 $X2=6.99
+ $Y2=0
r112 60 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.825 $Y=0 $X2=6.48
+ $Y2=0
r113 59 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r114 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r115 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r116 56 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r117 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r118 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r119 53 77 10.6558 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.302
+ $Y2=0
r120 53 55 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.56
+ $Y2=0
r121 52 80 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.985
+ $Y2=0
r122 52 58 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.835 $Y=0
+ $X2=5.52 $Y2=0
r123 51 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r124 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r125 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r126 48 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r127 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r128 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r129 45 71 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.915 $Y=0
+ $X2=0.787 $Y2=0
r130 45 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.2
+ $Y2=0
r131 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.505
+ $Y2=0
r132 44 50 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.16
+ $Y2=0
r133 42 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r134 42 75 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=2.64
+ $Y2=0
r135 38 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0
r136 38 40 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0.54
r137 34 36 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=5.985 $Y=0.46
+ $X2=5.985 $Y2=1.005
r138 32 80 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=0.085
+ $X2=5.985 $Y2=0
r139 32 34 14.4055 $w=2.98e-07 $l=3.75e-07 $layer=LI1_cond $X=5.985 $Y=0.085
+ $X2=5.985 $Y2=0.46
r140 28 77 1.82608 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.302 $Y=0.085
+ $X2=4.302 $Y2=0
r141 28 30 7.75479 $w=4.53e-07 $l=2.95e-07 $layer=LI1_cond $X=4.302 $Y=0.085
+ $X2=4.302 $Y2=0.38
r142 27 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.505
+ $Y2=0
r143 26 77 10.6558 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=4.075 $Y=0
+ $X2=4.302 $Y2=0
r144 26 27 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=4.075 $Y=0
+ $X2=2.67 $Y2=0
r145 22 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.085
+ $X2=2.505 $Y2=0
r146 22 24 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.505 $Y=0.085
+ $X2=2.505 $Y2=0.41
r147 18 71 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.787 $Y=0.085
+ $X2=0.787 $Y2=0
r148 18 20 18.9814 $w=2.53e-07 $l=4.2e-07 $layer=LI1_cond $X=0.787 $Y=0.085
+ $X2=0.787 $Y2=0.505
r149 5 40 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.865
+ $Y=0.395 $X2=6.99 $Y2=0.54
r150 4 36 182 $w=1.7e-07 $l=7.7479e-07 $layer=licon1_NDIFF $count=1 $X=5.805
+ $Y=0.315 $X2=5.985 $Y2=1.005
r151 4 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.805
+ $Y=0.315 $X2=5.945 $Y2=0.46
r152 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.1
+ $Y=0.235 $X2=4.24 $Y2=0.38
r153 2 24 182 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_NDIFF $count=1 $X=2.32
+ $Y=0.235 $X2=2.505 $Y2=0.41
r154 1 20 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.645
+ $Y=0.31 $X2=0.785 $Y2=0.505
.ends

