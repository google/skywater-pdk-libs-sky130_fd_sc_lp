* File: sky130_fd_sc_lp__dlrbp_2.pxi.spice
* Created: Fri Aug 28 10:26:09 2020
* 
x_PM_SKY130_FD_SC_LP__DLRBP_2%A_80_21# N_A_80_21#_M1009_s N_A_80_21#_M1021_s
+ N_A_80_21#_M1007_g N_A_80_21#_M1006_g N_A_80_21#_M1012_g N_A_80_21#_M1027_g
+ N_A_80_21#_c_176_n N_A_80_21#_c_177_n N_A_80_21#_c_178_n N_A_80_21#_c_179_n
+ N_A_80_21#_c_180_n N_A_80_21#_c_181_n PM_SKY130_FD_SC_LP__DLRBP_2%A_80_21#
x_PM_SKY130_FD_SC_LP__DLRBP_2%A_432_109# N_A_432_109#_M1005_d
+ N_A_432_109#_M1003_d N_A_432_109#_c_221_n N_A_432_109#_M1009_g
+ N_A_432_109#_M1021_g N_A_432_109#_c_222_n N_A_432_109#_M1011_g
+ N_A_432_109#_M1001_g N_A_432_109#_c_223_n N_A_432_109#_M1025_g
+ N_A_432_109#_M1014_g N_A_432_109#_M1015_g N_A_432_109#_M1019_g
+ N_A_432_109#_c_234_n N_A_432_109#_c_225_n N_A_432_109#_c_251_p
+ N_A_432_109#_c_333_p N_A_432_109#_c_235_n N_A_432_109#_c_253_p
+ N_A_432_109#_c_236_n N_A_432_109#_c_226_n N_A_432_109#_c_227_n
+ N_A_432_109#_c_237_n N_A_432_109#_c_228_n N_A_432_109#_c_229_n
+ PM_SKY130_FD_SC_LP__DLRBP_2%A_432_109#
x_PM_SKY130_FD_SC_LP__DLRBP_2%RESET_B N_RESET_B_M1002_g N_RESET_B_c_359_n
+ N_RESET_B_M1003_g RESET_B N_RESET_B_c_360_n
+ PM_SKY130_FD_SC_LP__DLRBP_2%RESET_B
x_PM_SKY130_FD_SC_LP__DLRBP_2%A_823_25# N_A_823_25#_M1013_d N_A_823_25#_M1000_d
+ N_A_823_25#_c_394_n N_A_823_25#_M1005_g N_A_823_25#_M1022_g
+ N_A_823_25#_c_396_n N_A_823_25#_c_397_n N_A_823_25#_c_398_n
+ N_A_823_25#_c_421_n N_A_823_25#_c_399_n N_A_823_25#_c_403_n
+ N_A_823_25#_c_400_n N_A_823_25#_c_401_n PM_SKY130_FD_SC_LP__DLRBP_2%A_823_25#
x_PM_SKY130_FD_SC_LP__DLRBP_2%A_1023_405# N_A_1023_405#_M1010_s
+ N_A_1023_405#_M1004_s N_A_1023_405#_M1000_g N_A_1023_405#_M1018_g
+ N_A_1023_405#_c_485_n N_A_1023_405#_c_486_n N_A_1023_405#_c_487_n
+ N_A_1023_405#_c_478_n N_A_1023_405#_c_521_p N_A_1023_405#_c_522_p
+ N_A_1023_405#_c_523_p N_A_1023_405#_c_489_n N_A_1023_405#_c_479_n
+ N_A_1023_405#_c_480_n N_A_1023_405#_c_481_n N_A_1023_405#_c_563_p
+ N_A_1023_405#_c_482_n N_A_1023_405#_c_491_n N_A_1023_405#_c_492_n
+ N_A_1023_405#_c_493_n N_A_1023_405#_c_483_n
+ PM_SKY130_FD_SC_LP__DLRBP_2%A_1023_405#
x_PM_SKY130_FD_SC_LP__DLRBP_2%A_1246_339# N_A_1246_339#_M1026_d
+ N_A_1246_339#_M1017_d N_A_1246_339#_M1023_g N_A_1246_339#_M1024_g
+ N_A_1246_339#_c_616_n N_A_1246_339#_c_617_n N_A_1246_339#_c_618_n
+ N_A_1246_339#_c_619_n N_A_1246_339#_c_620_n N_A_1246_339#_c_625_n
+ N_A_1246_339#_c_621_n N_A_1246_339#_c_627_n
+ PM_SKY130_FD_SC_LP__DLRBP_2%A_1246_339#
x_PM_SKY130_FD_SC_LP__DLRBP_2%D N_D_M1026_g N_D_M1017_g N_D_c_692_n N_D_c_697_n
+ D D N_D_c_694_n PM_SKY130_FD_SC_LP__DLRBP_2%D
x_PM_SKY130_FD_SC_LP__DLRBP_2%A_1109_21# N_A_1109_21#_M1020_d
+ N_A_1109_21#_M1008_d N_A_1109_21#_M1013_g N_A_1109_21#_c_740_n
+ N_A_1109_21#_c_741_n N_A_1109_21#_M1016_g N_A_1109_21#_c_742_n
+ N_A_1109_21#_c_743_n N_A_1109_21#_c_744_n N_A_1109_21#_c_745_n
+ N_A_1109_21#_M1010_g N_A_1109_21#_M1004_g N_A_1109_21#_c_755_n
+ N_A_1109_21#_c_746_n N_A_1109_21#_c_756_n N_A_1109_21#_c_757_n
+ N_A_1109_21#_c_747_n N_A_1109_21#_c_748_n N_A_1109_21#_c_749_n
+ N_A_1109_21#_c_760_n N_A_1109_21#_c_761_n N_A_1109_21#_c_762_n
+ N_A_1109_21#_c_750_n N_A_1109_21#_c_751_n N_A_1109_21#_c_764_n
+ PM_SKY130_FD_SC_LP__DLRBP_2%A_1109_21#
x_PM_SKY130_FD_SC_LP__DLRBP_2%GATE N_GATE_M1020_g N_GATE_M1008_g N_GATE_c_866_n
+ N_GATE_c_867_n GATE GATE GATE GATE N_GATE_c_869_n
+ PM_SKY130_FD_SC_LP__DLRBP_2%GATE
x_PM_SKY130_FD_SC_LP__DLRBP_2%VPWR N_VPWR_M1006_d N_VPWR_M1027_d N_VPWR_M1021_d
+ N_VPWR_M1014_s N_VPWR_M1022_d N_VPWR_M1023_d N_VPWR_M1004_d N_VPWR_c_900_n
+ N_VPWR_c_901_n N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_904_n N_VPWR_c_905_n
+ N_VPWR_c_906_n N_VPWR_c_907_n VPWR N_VPWR_c_908_n N_VPWR_c_909_n
+ N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_913_n N_VPWR_c_914_n
+ N_VPWR_c_899_n N_VPWR_c_916_n N_VPWR_c_917_n N_VPWR_c_918_n N_VPWR_c_919_n
+ N_VPWR_c_920_n N_VPWR_c_921_n PM_SKY130_FD_SC_LP__DLRBP_2%VPWR
x_PM_SKY130_FD_SC_LP__DLRBP_2%Q_N N_Q_N_M1007_d N_Q_N_M1006_s Q_N Q_N Q_N
+ N_Q_N_c_1017_n PM_SKY130_FD_SC_LP__DLRBP_2%Q_N
x_PM_SKY130_FD_SC_LP__DLRBP_2%Q N_Q_M1011_d N_Q_M1001_d N_Q_c_1035_n
+ N_Q_c_1053_n N_Q_c_1043_n N_Q_c_1036_n Q Q Q Q N_Q_c_1039_n N_Q_c_1065_n Q
+ N_Q_c_1067_n PM_SKY130_FD_SC_LP__DLRBP_2%Q
x_PM_SKY130_FD_SC_LP__DLRBP_2%VGND N_VGND_M1007_s N_VGND_M1012_s N_VGND_M1009_d
+ N_VGND_M1025_s N_VGND_M1019_s N_VGND_M1024_d N_VGND_M1010_d N_VGND_c_1096_n
+ N_VGND_c_1097_n N_VGND_c_1098_n N_VGND_c_1099_n N_VGND_c_1100_n
+ N_VGND_c_1101_n N_VGND_c_1102_n N_VGND_c_1103_n N_VGND_c_1104_n
+ N_VGND_c_1105_n N_VGND_c_1106_n N_VGND_c_1107_n VGND N_VGND_c_1108_n
+ N_VGND_c_1109_n N_VGND_c_1110_n N_VGND_c_1111_n N_VGND_c_1112_n
+ N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n N_VGND_c_1116_n
+ N_VGND_c_1117_n PM_SKY130_FD_SC_LP__DLRBP_2%VGND
cc_1 VNB N_A_80_21#_M1007_g 0.0307442f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A_80_21#_M1006_g 0.00192821f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_A_80_21#_M1012_g 0.030727f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_4 VNB N_A_80_21#_M1027_g 0.00192821f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_5 VNB N_A_80_21#_c_176_n 0.0448647f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.465
cc_6 VNB N_A_80_21#_c_177_n 0.0449641f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.465
cc_7 VNB N_A_80_21#_c_178_n 0.0413785f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=1.465
cc_8 VNB N_A_80_21#_c_179_n 0.015006f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=0.885
cc_9 VNB N_A_80_21#_c_180_n 0.00128353f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.985
cc_10 VNB N_A_80_21#_c_181_n 0.00569221f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.465
cc_11 VNB N_A_432_109#_c_221_n 0.023598f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.3
cc_12 VNB N_A_432_109#_c_222_n 0.0194203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_432_109#_c_223_n 0.0164903f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_14 VNB N_A_432_109#_M1019_g 0.0404542f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=0.885
cc_15 VNB N_A_432_109#_c_225_n 0.0131566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_432_109#_c_226_n 0.00815377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_432_109#_c_227_n 0.0010628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_432_109#_c_228_n 0.0338591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_432_109#_c_229_n 0.0908462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_RESET_B_M1002_g 0.0237154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_RESET_B_c_359_n 0.0272317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_RESET_B_c_360_n 0.00417485f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_23 VNB N_A_823_25#_c_394_n 0.0212176f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.3
cc_24 VNB N_A_823_25#_M1022_g 0.00703991f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_25 VNB N_A_823_25#_c_396_n 0.0323363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_823_25#_c_397_n 0.0013965f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_27 VNB N_A_823_25#_c_398_n 0.00418387f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_28 VNB N_A_823_25#_c_399_n 0.00101974f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=1.465
cc_29 VNB N_A_823_25#_c_400_n 0.00219351f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=0.885
cc_30 VNB N_A_823_25#_c_401_n 0.0434387f $X=-0.19 $Y=-0.245 $X2=2.062 $Y2=1.63
cc_31 VNB N_A_1023_405#_c_478_n 0.00279887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1023_405#_c_479_n 0.0169918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1023_405#_c_480_n 0.00199024f $X=-0.19 $Y=-0.245 $X2=2.04
+ $Y2=0.885
cc_34 VNB N_A_1023_405#_c_481_n 0.0382382f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=0.885
cc_35 VNB N_A_1023_405#_c_482_n 7.78343e-19 $X=-0.19 $Y=-0.245 $X2=1.165
+ $Y2=1.465
cc_36 VNB N_A_1023_405#_c_483_n 0.0158353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1246_339#_M1024_g 0.0411622f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=2.465
cc_38 VNB N_A_1246_339#_c_616_n 0.00274621f $X=-0.19 $Y=-0.245 $X2=0.905
+ $Y2=0.655
cc_39 VNB N_A_1246_339#_c_617_n 0.0110695f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_40 VNB N_A_1246_339#_c_618_n 0.00558666f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.465
cc_41 VNB N_A_1246_339#_c_619_n 0.00576393f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=1.465
cc_42 VNB N_A_1246_339#_c_620_n 0.0120106f $X=-0.19 $Y=-0.245 $X2=1.875
+ $Y2=1.465
cc_43 VNB N_A_1246_339#_c_621_n 0.00799261f $X=-0.19 $Y=-0.245 $X2=1.165
+ $Y2=1.465
cc_44 VNB N_D_M1026_g 0.0345111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_D_c_692_n 0.00300895f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.63
cc_46 VNB D 0.0029498f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_47 VNB N_D_c_694_n 0.0167375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1109_21#_M1013_g 0.0495584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1109_21#_c_740_n 0.146045f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.63
cc_50 VNB N_A_1109_21#_c_741_n 0.0125466f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_51 VNB N_A_1109_21#_c_742_n 0.0300612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1109_21#_c_743_n 0.0208548f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.63
cc_53 VNB N_A_1109_21#_c_744_n 0.0135695f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_54 VNB N_A_1109_21#_c_745_n 0.016975f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_55 VNB N_A_1109_21#_c_746_n 0.0386961f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.3
cc_56 VNB N_A_1109_21#_c_747_n 0.00534699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1109_21#_c_748_n 6.84479e-19 $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.985
cc_58 VNB N_A_1109_21#_c_749_n 0.0128524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1109_21#_c_750_n 0.050156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1109_21#_c_751_n 0.017037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_GATE_M1020_g 0.0241407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_GATE_M1008_g 0.00853481f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.3
cc_63 VNB N_GATE_c_866_n 0.0242144f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.63
cc_64 VNB N_GATE_c_867_n 0.0190903f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_65 VNB GATE 0.01178f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_66 VNB N_GATE_c_869_n 0.0168314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VPWR_c_899_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_Q_N_c_1017_n 0.00507155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_Q_c_1035_n 0.00173506f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_70 VNB N_Q_c_1036_n 0.00120514f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_71 VNB N_VGND_c_1096_n 0.0108094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1097_n 0.049388f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.465
cc_73 VNB N_VGND_c_1098_n 0.0315791f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.465
cc_74 VNB N_VGND_c_1099_n 0.015333f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1100_n 0.00626856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1101_n 0.0183093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1102_n 0.0115176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1103_n 0.00524934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1104_n 0.0405179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1105_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1106_n 0.0342111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1107_n 0.00507191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1108_n 0.0169258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1109_n 0.0341729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1110_n 0.0174868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1111_n 0.0330002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1112_n 0.0206396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1113_n 0.496923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1114_n 0.00548191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1115_n 0.00631443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1116_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1117_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VPB N_A_80_21#_M1006_g 0.0272796f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_94 VPB N_A_80_21#_M1027_g 0.0272796f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_95 VPB N_A_80_21#_c_180_n 0.0151221f $X=-0.19 $Y=1.655 $X2=2.1 $Y2=1.985
cc_96 VPB N_A_432_109#_M1021_g 0.0247645f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_97 VPB N_A_432_109#_M1001_g 0.020574f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.63
cc_98 VPB N_A_432_109#_M1014_g 0.0191184f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.465
cc_99 VPB N_A_432_109#_M1015_g 0.0577466f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=1.465
cc_100 VPB N_A_432_109#_c_234_n 0.00142203f $X=-0.19 $Y=1.655 $X2=2.1 $Y2=1.985
cc_101 VPB N_A_432_109#_c_235_n 0.00444711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_432_109#_c_236_n 0.0069408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_432_109#_c_237_n 0.00925285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_432_109#_c_228_n 0.0171849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_432_109#_c_229_n 0.0147324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_RESET_B_c_359_n 0.0289067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_RESET_B_c_360_n 0.00330621f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_108 VPB N_A_823_25#_M1022_g 0.0214399f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_109 VPB N_A_823_25#_c_403_n 7.50226e-19 $X=-0.19 $Y=1.655 $X2=2.04 $Y2=1.3
cc_110 VPB N_A_823_25#_c_400_n 0.0116596f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=0.885
cc_111 VPB N_A_1023_405#_M1000_g 0.0208632f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=0.655
cc_112 VPB N_A_1023_405#_c_485_n 0.00137967f $X=-0.19 $Y=1.655 $X2=0.905
+ $Y2=0.655
cc_113 VPB N_A_1023_405#_c_486_n 0.00469675f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.63
cc_114 VPB N_A_1023_405#_c_487_n 0.0022701f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_115 VPB N_A_1023_405#_c_478_n 0.0049121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_1023_405#_c_489_n 0.00139769f $X=-0.19 $Y=1.655 $X2=1.165
+ $Y2=1.465
cc_117 VPB N_A_1023_405#_c_479_n 0.0200456f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_1023_405#_c_491_n 0.0115812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_1023_405#_c_492_n 0.00663494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_1023_405#_c_493_n 0.0440083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_1246_339#_M1023_g 0.0271677f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=0.655
cc_122 VPB N_A_1246_339#_M1024_g 0.00220946f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=2.465
cc_123 VPB N_A_1246_339#_c_616_n 0.00291784f $X=-0.19 $Y=1.655 $X2=0.905
+ $Y2=0.655
cc_124 VPB N_A_1246_339#_c_625_n 0.0028323f $X=-0.19 $Y=1.655 $X2=1.165
+ $Y2=1.465
cc_125 VPB N_A_1246_339#_c_621_n 0.0127154f $X=-0.19 $Y=1.655 $X2=1.165
+ $Y2=1.465
cc_126 VPB N_A_1246_339#_c_627_n 0.0390412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_D_M1017_g 0.0263103f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.3
cc_128 VPB N_D_c_692_n 0.0230686f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.63
cc_129 VPB N_D_c_697_n 0.0187934f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_130 VPB D 0.00572469f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_131 VPB N_A_1109_21#_M1013_g 3.65257e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_1109_21#_M1016_g 0.0322763f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.3
cc_133 VPB N_A_1109_21#_M1004_g 0.0228829f $X=-0.19 $Y=1.655 $X2=1.875 $Y2=1.465
cc_134 VPB N_A_1109_21#_c_755_n 0.0377067f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=1.465
cc_135 VPB N_A_1109_21#_c_756_n 0.0286711f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=0.885
cc_136 VPB N_A_1109_21#_c_757_n 0.0183275f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=0.885
cc_137 VPB N_A_1109_21#_c_748_n 4.04609e-19 $X=-0.19 $Y=1.655 $X2=2.1 $Y2=1.985
cc_138 VPB N_A_1109_21#_c_749_n 0.00805843f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_1109_21#_c_760_n 0.00564023f $X=-0.19 $Y=1.655 $X2=1.165
+ $Y2=1.465
cc_140 VPB N_A_1109_21#_c_761_n 0.00107991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_1109_21#_c_762_n 0.0268487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_1109_21#_c_750_n 0.0310756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_1109_21#_c_764_n 0.0142804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_GATE_M1008_g 0.0571388f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.3
cc_145 VPB GATE 0.00927821f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_146 VPB N_VPWR_c_900_n 0.0107835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_901_n 0.0654008f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.465
cc_148 VPB N_VPWR_c_902_n 0.0442734f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=1.465
cc_149 VPB N_VPWR_c_903_n 0.0198296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_904_n 0.00442439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_905_n 0.00988942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_906_n 0.00839603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_907_n 0.00151893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_908_n 0.0169386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_909_n 0.0371681f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_910_n 0.0160372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_911_n 0.0157463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_912_n 0.0452663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_913_n 0.0377191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_914_n 0.0173809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_899_n 0.109231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_916_n 0.00555219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_917_n 0.00522677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_918_n 0.0063201f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_919_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_920_n 0.00651591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_921_n 0.00485691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_Q_N_c_1017_n 0.00353065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_Q_c_1035_n 0.00234053f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_170 VPB Q 8.78261e-19 $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.655
cc_171 VPB N_Q_c_1039_n 0.031946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 N_A_80_21#_c_179_n N_A_432_109#_c_221_n 0.00975599f $X=2.02 $Y=0.885
+ $X2=0 $Y2=0
cc_173 N_A_80_21#_c_179_n N_A_432_109#_c_229_n 0.00379584f $X=2.02 $Y=0.885
+ $X2=0 $Y2=0
cc_174 N_A_80_21#_c_180_n N_A_432_109#_c_229_n 0.00532908f $X=2.1 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_80_21#_c_181_n N_A_432_109#_c_229_n 0.0128515f $X=2.04 $Y=1.465 $X2=0
+ $Y2=0
cc_176 N_A_80_21#_M1006_g N_VPWR_c_901_n 0.00769005f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_80_21#_M1027_g N_VPWR_c_902_n 0.00769005f $X=0.91 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_80_21#_c_177_n N_VPWR_c_902_n 0.022791f $X=1.875 $Y=1.465 $X2=0 $Y2=0
cc_179 N_A_80_21#_c_178_n N_VPWR_c_902_n 0.00665919f $X=1.165 $Y=1.465 $X2=0
+ $Y2=0
cc_180 N_A_80_21#_c_180_n N_VPWR_c_902_n 0.0109699f $X=2.1 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_80_21#_M1006_g N_VPWR_c_908_n 0.00585385f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_80_21#_M1027_g N_VPWR_c_908_n 0.00585385f $X=0.91 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_80_21#_M1006_g N_VPWR_c_899_n 0.0114817f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_80_21#_M1027_g N_VPWR_c_899_n 0.0118488f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_80_21#_M1007_g N_Q_N_c_1017_n 0.0064542f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_186 N_A_80_21#_M1006_g N_Q_N_c_1017_n 0.00613418f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_80_21#_M1012_g N_Q_N_c_1017_n 0.00649413f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_188 N_A_80_21#_M1027_g N_Q_N_c_1017_n 0.00613418f $X=0.91 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_A_80_21#_c_176_n N_Q_N_c_1017_n 0.0315277f $X=0.985 $Y=1.465 $X2=0
+ $Y2=0
cc_190 N_A_80_21#_c_177_n N_Q_N_c_1017_n 0.0258419f $X=1.875 $Y=1.465 $X2=0
+ $Y2=0
cc_191 N_A_80_21#_c_179_n N_Q_c_1035_n 0.0270455f $X=2.02 $Y=0.885 $X2=0 $Y2=0
cc_192 N_A_80_21#_c_180_n N_Q_c_1035_n 0.0126828f $X=2.1 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_80_21#_c_181_n N_Q_c_1035_n 0.0209919f $X=2.04 $Y=1.465 $X2=0 $Y2=0
cc_194 N_A_80_21#_c_179_n N_Q_c_1043_n 0.00785117f $X=2.02 $Y=0.885 $X2=0 $Y2=0
cc_195 N_A_80_21#_M1021_s N_Q_c_1039_n 0.0033187f $X=1.955 $Y=1.835 $X2=0 $Y2=0
cc_196 N_A_80_21#_c_180_n N_Q_c_1039_n 0.0214214f $X=2.1 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_80_21#_M1007_g N_VGND_c_1097_n 0.00708945f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_198 N_A_80_21#_M1012_g N_VGND_c_1098_n 0.0070315f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_199 N_A_80_21#_c_177_n N_VGND_c_1098_n 0.0207405f $X=1.875 $Y=1.465 $X2=0
+ $Y2=0
cc_200 N_A_80_21#_c_178_n N_VGND_c_1098_n 0.00647511f $X=1.165 $Y=1.465 $X2=0
+ $Y2=0
cc_201 N_A_80_21#_c_179_n N_VGND_c_1098_n 0.0131827f $X=2.02 $Y=0.885 $X2=0
+ $Y2=0
cc_202 N_A_80_21#_M1007_g N_VGND_c_1108_n 0.00585385f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_203 N_A_80_21#_M1012_g N_VGND_c_1108_n 0.00585385f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_204 N_A_80_21#_c_179_n N_VGND_c_1109_n 0.00483641f $X=2.02 $Y=0.885 $X2=0
+ $Y2=0
cc_205 N_A_80_21#_M1007_g N_VGND_c_1113_n 0.0114687f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_206 N_A_80_21#_M1012_g N_VGND_c_1113_n 0.0118494f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_207 N_A_80_21#_c_179_n N_VGND_c_1113_n 0.009312f $X=2.02 $Y=0.885 $X2=0 $Y2=0
cc_208 N_A_432_109#_c_223_n N_RESET_B_M1002_g 0.0249889f $X=3.29 $Y=1.205 $X2=0
+ $Y2=0
cc_209 N_A_432_109#_c_225_n N_RESET_B_M1002_g 0.0171314f $X=3.91 $Y=1.09 $X2=0
+ $Y2=0
cc_210 N_A_432_109#_c_226_n N_RESET_B_M1002_g 0.00161331f $X=4.405 $Y=0.42 $X2=0
+ $Y2=0
cc_211 N_A_432_109#_c_227_n N_RESET_B_M1002_g 9.22877e-19 $X=3.2 $Y=1.37 $X2=0
+ $Y2=0
cc_212 N_A_432_109#_M1014_g N_RESET_B_c_359_n 0.0329166f $X=3.29 $Y=2.465 $X2=0
+ $Y2=0
cc_213 N_A_432_109#_c_234_n N_RESET_B_c_359_n 8.44003e-19 $X=3.25 $Y=1.92 $X2=0
+ $Y2=0
cc_214 N_A_432_109#_c_225_n N_RESET_B_c_359_n 0.00282936f $X=3.91 $Y=1.09 $X2=0
+ $Y2=0
cc_215 N_A_432_109#_c_251_p N_RESET_B_c_359_n 0.0161577f $X=3.925 $Y=2.005 $X2=0
+ $Y2=0
cc_216 N_A_432_109#_c_235_n N_RESET_B_c_359_n 0.00321692f $X=4.055 $Y=2.09 $X2=0
+ $Y2=0
cc_217 N_A_432_109#_c_253_p N_RESET_B_c_359_n 0.0137947f $X=4.09 $Y=2.91 $X2=0
+ $Y2=0
cc_218 N_A_432_109#_c_229_n N_RESET_B_c_359_n 0.0241805f $X=3.29 $Y=1.445 $X2=0
+ $Y2=0
cc_219 N_A_432_109#_c_234_n N_RESET_B_c_360_n 0.016124f $X=3.25 $Y=1.92 $X2=0
+ $Y2=0
cc_220 N_A_432_109#_c_225_n N_RESET_B_c_360_n 0.0244321f $X=3.91 $Y=1.09 $X2=0
+ $Y2=0
cc_221 N_A_432_109#_c_251_p N_RESET_B_c_360_n 0.0230841f $X=3.925 $Y=2.005 $X2=0
+ $Y2=0
cc_222 N_A_432_109#_c_235_n N_RESET_B_c_360_n 0.00290748f $X=4.055 $Y=2.09 $X2=0
+ $Y2=0
cc_223 N_A_432_109#_c_227_n N_RESET_B_c_360_n 0.0156746f $X=3.2 $Y=1.37 $X2=0
+ $Y2=0
cc_224 N_A_432_109#_c_229_n N_RESET_B_c_360_n 0.0026775f $X=3.29 $Y=1.445 $X2=0
+ $Y2=0
cc_225 N_A_432_109#_c_225_n N_A_823_25#_c_394_n 0.0154731f $X=3.91 $Y=1.09 $X2=0
+ $Y2=0
cc_226 N_A_432_109#_c_226_n N_A_823_25#_c_394_n 0.0106075f $X=4.405 $Y=0.42
+ $X2=0 $Y2=0
cc_227 N_A_432_109#_c_236_n N_A_823_25#_M1022_g 0.0145189f $X=4.805 $Y=1.8 $X2=0
+ $Y2=0
cc_228 N_A_432_109#_c_237_n N_A_823_25#_M1022_g 0.00108723f $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_229 N_A_432_109#_c_228_n N_A_823_25#_M1022_g 0.0268963f $X=4.97 $Y=1.62 $X2=0
+ $Y2=0
cc_230 N_A_432_109#_M1019_g N_A_823_25#_c_396_n 0.0161239f $X=5.26 $Y=0.805
+ $X2=0 $Y2=0
cc_231 N_A_432_109#_c_225_n N_A_823_25#_c_396_n 0.00210266f $X=3.91 $Y=1.09
+ $X2=0 $Y2=0
cc_232 N_A_432_109#_c_236_n N_A_823_25#_c_396_n 0.0114606f $X=4.805 $Y=1.8 $X2=0
+ $Y2=0
cc_233 N_A_432_109#_c_237_n N_A_823_25#_c_396_n 0.0249357f $X=4.97 $Y=1.62 $X2=0
+ $Y2=0
cc_234 N_A_432_109#_c_228_n N_A_823_25#_c_396_n 0.0115859f $X=4.97 $Y=1.62 $X2=0
+ $Y2=0
cc_235 N_A_432_109#_M1019_g N_A_823_25#_c_397_n 0.00123926f $X=5.26 $Y=0.805
+ $X2=0 $Y2=0
cc_236 N_A_432_109#_M1019_g N_A_823_25#_c_398_n 6.02135e-19 $X=5.26 $Y=0.805
+ $X2=0 $Y2=0
cc_237 N_A_432_109#_c_225_n N_A_823_25#_c_398_n 0.0229221f $X=3.91 $Y=1.09 $X2=0
+ $Y2=0
cc_238 N_A_432_109#_c_236_n N_A_823_25#_c_398_n 0.0207993f $X=4.805 $Y=1.8 $X2=0
+ $Y2=0
cc_239 N_A_432_109#_c_237_n N_A_823_25#_c_398_n 5.29882e-19 $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_240 N_A_432_109#_c_228_n N_A_823_25#_c_398_n 5.49534e-19 $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_241 N_A_432_109#_M1019_g N_A_823_25#_c_421_n 9.16434e-19 $X=5.26 $Y=0.805
+ $X2=0 $Y2=0
cc_242 N_A_432_109#_M1019_g N_A_823_25#_c_400_n 0.00129056f $X=5.26 $Y=0.805
+ $X2=0 $Y2=0
cc_243 N_A_432_109#_c_237_n N_A_823_25#_c_400_n 0.0115224f $X=4.97 $Y=1.62 $X2=0
+ $Y2=0
cc_244 N_A_432_109#_c_228_n N_A_823_25#_c_400_n 6.89982e-19 $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_245 N_A_432_109#_M1019_g N_A_823_25#_c_401_n 0.00382466f $X=5.26 $Y=0.805
+ $X2=0 $Y2=0
cc_246 N_A_432_109#_c_225_n N_A_823_25#_c_401_n 0.00191197f $X=3.91 $Y=1.09
+ $X2=0 $Y2=0
cc_247 N_A_432_109#_c_235_n N_A_823_25#_c_401_n 0.00276767f $X=4.055 $Y=2.09
+ $X2=0 $Y2=0
cc_248 N_A_432_109#_c_236_n N_A_823_25#_c_401_n 0.00276109f $X=4.805 $Y=1.8
+ $X2=0 $Y2=0
cc_249 N_A_432_109#_c_228_n N_A_823_25#_c_401_n 0.00439289f $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_250 N_A_432_109#_M1015_g N_A_1023_405#_M1000_g 0.0160219f $X=4.83 $Y=2.725
+ $X2=0 $Y2=0
cc_251 N_A_432_109#_M1015_g N_A_1023_405#_c_485_n 0.00535846f $X=4.83 $Y=2.725
+ $X2=0 $Y2=0
cc_252 N_A_432_109#_c_237_n N_A_1023_405#_c_485_n 0.00152785f $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_253 N_A_432_109#_c_228_n N_A_1023_405#_c_485_n 0.00126922f $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_254 N_A_432_109#_M1015_g N_A_1023_405#_c_487_n 0.0018782f $X=4.83 $Y=2.725
+ $X2=0 $Y2=0
cc_255 N_A_432_109#_M1015_g N_A_1023_405#_c_493_n 0.0203417f $X=4.83 $Y=2.725
+ $X2=0 $Y2=0
cc_256 N_A_432_109#_c_228_n N_A_1023_405#_c_493_n 0.00691002f $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_257 N_A_432_109#_M1019_g N_A_1109_21#_M1013_g 0.069253f $X=5.26 $Y=0.805
+ $X2=0 $Y2=0
cc_258 N_A_432_109#_c_237_n N_A_1109_21#_M1013_g 0.00105665f $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_259 N_A_432_109#_c_228_n N_A_1109_21#_M1013_g 0.00516921f $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_260 N_A_432_109#_M1015_g N_A_1109_21#_c_755_n 3.84066e-19 $X=4.83 $Y=2.725
+ $X2=0 $Y2=0
cc_261 N_A_432_109#_c_237_n N_A_1109_21#_c_755_n 4.48311e-19 $X=4.97 $Y=1.62
+ $X2=0 $Y2=0
cc_262 N_A_432_109#_c_251_p N_VPWR_M1014_s 0.00946867f $X=3.925 $Y=2.005 $X2=0
+ $Y2=0
cc_263 N_A_432_109#_c_236_n N_VPWR_M1022_d 0.00225176f $X=4.805 $Y=1.8 $X2=0
+ $Y2=0
cc_264 N_A_432_109#_M1001_g N_VPWR_c_903_n 0.0105471f $X=2.86 $Y=2.465 $X2=0
+ $Y2=0
cc_265 N_A_432_109#_M1014_g N_VPWR_c_903_n 5.99361e-19 $X=3.29 $Y=2.465 $X2=0
+ $Y2=0
cc_266 N_A_432_109#_M1014_g N_VPWR_c_904_n 0.00690677f $X=3.29 $Y=2.465 $X2=0
+ $Y2=0
cc_267 N_A_432_109#_c_251_p N_VPWR_c_904_n 0.0261161f $X=3.925 $Y=2.005 $X2=0
+ $Y2=0
cc_268 N_A_432_109#_M1015_g N_VPWR_c_905_n 0.014142f $X=4.83 $Y=2.725 $X2=0
+ $Y2=0
cc_269 N_A_432_109#_c_236_n N_VPWR_c_905_n 0.0220026f $X=4.805 $Y=1.8 $X2=0
+ $Y2=0
cc_270 N_A_432_109#_M1021_g N_VPWR_c_909_n 0.00312414f $X=2.315 $Y=2.155 $X2=0
+ $Y2=0
cc_271 N_A_432_109#_M1001_g N_VPWR_c_910_n 0.00564095f $X=2.86 $Y=2.465 $X2=0
+ $Y2=0
cc_272 N_A_432_109#_M1014_g N_VPWR_c_910_n 0.0054895f $X=3.29 $Y=2.465 $X2=0
+ $Y2=0
cc_273 N_A_432_109#_c_253_p N_VPWR_c_911_n 0.015688f $X=4.09 $Y=2.91 $X2=0 $Y2=0
cc_274 N_A_432_109#_M1015_g N_VPWR_c_912_n 0.00559701f $X=4.83 $Y=2.725 $X2=0
+ $Y2=0
cc_275 N_A_432_109#_M1003_d N_VPWR_c_899_n 0.00380103f $X=3.95 $Y=1.835 $X2=0
+ $Y2=0
cc_276 N_A_432_109#_M1021_g N_VPWR_c_899_n 0.00410284f $X=2.315 $Y=2.155 $X2=0
+ $Y2=0
cc_277 N_A_432_109#_M1001_g N_VPWR_c_899_n 0.00518386f $X=2.86 $Y=2.465 $X2=0
+ $Y2=0
cc_278 N_A_432_109#_M1014_g N_VPWR_c_899_n 0.0102673f $X=3.29 $Y=2.465 $X2=0
+ $Y2=0
cc_279 N_A_432_109#_M1015_g N_VPWR_c_899_n 0.00537853f $X=4.83 $Y=2.725 $X2=0
+ $Y2=0
cc_280 N_A_432_109#_c_253_p N_VPWR_c_899_n 0.00984745f $X=4.09 $Y=2.91 $X2=0
+ $Y2=0
cc_281 N_A_432_109#_c_221_n N_Q_c_1035_n 0.00328493f $X=2.235 $Y=1.205 $X2=0
+ $Y2=0
cc_282 N_A_432_109#_M1021_g N_Q_c_1035_n 0.00386906f $X=2.315 $Y=2.155 $X2=0
+ $Y2=0
cc_283 N_A_432_109#_c_222_n N_Q_c_1035_n 0.00602077f $X=2.86 $Y=1.205 $X2=0
+ $Y2=0
cc_284 N_A_432_109#_M1001_g N_Q_c_1035_n 0.00790116f $X=2.86 $Y=2.465 $X2=0
+ $Y2=0
cc_285 N_A_432_109#_c_234_n N_Q_c_1035_n 0.00994653f $X=3.25 $Y=1.92 $X2=0 $Y2=0
cc_286 N_A_432_109#_c_227_n N_Q_c_1035_n 0.029806f $X=3.2 $Y=1.37 $X2=0 $Y2=0
cc_287 N_A_432_109#_c_229_n N_Q_c_1035_n 0.0292119f $X=3.29 $Y=1.445 $X2=0 $Y2=0
cc_288 N_A_432_109#_c_222_n N_Q_c_1053_n 0.0111373f $X=2.86 $Y=1.205 $X2=0 $Y2=0
cc_289 N_A_432_109#_c_223_n N_Q_c_1053_n 0.00218767f $X=3.29 $Y=1.205 $X2=0
+ $Y2=0
cc_290 N_A_432_109#_c_227_n N_Q_c_1053_n 0.0167707f $X=3.2 $Y=1.37 $X2=0 $Y2=0
cc_291 N_A_432_109#_c_229_n N_Q_c_1053_n 0.00505525f $X=3.29 $Y=1.445 $X2=0
+ $Y2=0
cc_292 N_A_432_109#_c_221_n N_Q_c_1043_n 0.00308722f $X=2.235 $Y=1.205 $X2=0
+ $Y2=0
cc_293 N_A_432_109#_c_221_n N_Q_c_1036_n 4.85288e-19 $X=2.235 $Y=1.205 $X2=0
+ $Y2=0
cc_294 N_A_432_109#_c_222_n N_Q_c_1036_n 0.00825451f $X=2.86 $Y=1.205 $X2=0
+ $Y2=0
cc_295 N_A_432_109#_c_223_n N_Q_c_1036_n 0.00428601f $X=3.29 $Y=1.205 $X2=0
+ $Y2=0
cc_296 N_A_432_109#_M1014_g Q 0.00276097f $X=3.29 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A_432_109#_c_333_p Q 0.00207395f $X=3.335 $Y=2.005 $X2=0 $Y2=0
cc_298 N_A_432_109#_c_229_n Q 0.00303397f $X=3.29 $Y=1.445 $X2=0 $Y2=0
cc_299 N_A_432_109#_M1021_g N_Q_c_1039_n 0.0187697f $X=2.315 $Y=2.155 $X2=0
+ $Y2=0
cc_300 N_A_432_109#_M1001_g N_Q_c_1065_n 0.0170685f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A_432_109#_c_229_n N_Q_c_1065_n 0.00238641f $X=3.29 $Y=1.445 $X2=0
+ $Y2=0
cc_302 N_A_432_109#_M1014_g N_Q_c_1067_n 0.00761245f $X=3.29 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_432_109#_c_225_n N_VGND_M1025_s 0.00308172f $X=3.91 $Y=1.09 $X2=0
+ $Y2=0
cc_304 N_A_432_109#_c_222_n N_VGND_c_1099_n 0.00857457f $X=2.86 $Y=1.205 $X2=0
+ $Y2=0
cc_305 N_A_432_109#_c_223_n N_VGND_c_1100_n 0.00638719f $X=3.29 $Y=1.205 $X2=0
+ $Y2=0
cc_306 N_A_432_109#_c_225_n N_VGND_c_1100_n 0.022455f $X=3.91 $Y=1.09 $X2=0
+ $Y2=0
cc_307 N_A_432_109#_M1019_g N_VGND_c_1101_n 0.0118647f $X=5.26 $Y=0.805 $X2=0
+ $Y2=0
cc_308 N_A_432_109#_c_225_n N_VGND_c_1101_n 0.0078419f $X=3.91 $Y=1.09 $X2=0
+ $Y2=0
cc_309 N_A_432_109#_c_226_n N_VGND_c_1101_n 0.031824f $X=4.405 $Y=0.42 $X2=0
+ $Y2=0
cc_310 N_A_432_109#_M1019_g N_VGND_c_1104_n 0.0035863f $X=5.26 $Y=0.805 $X2=0
+ $Y2=0
cc_311 N_A_432_109#_c_221_n N_VGND_c_1109_n 0.00365453f $X=2.235 $Y=1.205 $X2=0
+ $Y2=0
cc_312 N_A_432_109#_c_222_n N_VGND_c_1110_n 0.0040172f $X=2.86 $Y=1.205 $X2=0
+ $Y2=0
cc_313 N_A_432_109#_c_223_n N_VGND_c_1110_n 0.00529818f $X=3.29 $Y=1.205 $X2=0
+ $Y2=0
cc_314 N_A_432_109#_c_226_n N_VGND_c_1111_n 0.0210192f $X=4.405 $Y=0.42 $X2=0
+ $Y2=0
cc_315 N_A_432_109#_c_221_n N_VGND_c_1113_n 0.00455831f $X=2.235 $Y=1.205 $X2=0
+ $Y2=0
cc_316 N_A_432_109#_c_222_n N_VGND_c_1113_n 0.00681483f $X=2.86 $Y=1.205 $X2=0
+ $Y2=0
cc_317 N_A_432_109#_c_223_n N_VGND_c_1113_n 0.00997058f $X=3.29 $Y=1.205 $X2=0
+ $Y2=0
cc_318 N_A_432_109#_M1019_g N_VGND_c_1113_n 0.00401353f $X=5.26 $Y=0.805 $X2=0
+ $Y2=0
cc_319 N_A_432_109#_c_225_n N_VGND_c_1113_n 0.0109859f $X=3.91 $Y=1.09 $X2=0
+ $Y2=0
cc_320 N_A_432_109#_c_226_n N_VGND_c_1113_n 0.0126321f $X=4.405 $Y=0.42 $X2=0
+ $Y2=0
cc_321 N_A_432_109#_c_225_n A_781_51# 0.00208937f $X=3.91 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_322 N_RESET_B_M1002_g N_A_823_25#_c_394_n 0.03684f $X=3.83 $Y=0.675 $X2=0
+ $Y2=0
cc_323 N_RESET_B_c_359_n N_A_823_25#_M1022_g 0.0267491f $X=3.875 $Y=1.715 $X2=0
+ $Y2=0
cc_324 N_RESET_B_c_360_n N_A_823_25#_M1022_g 9.12183e-19 $X=3.74 $Y=1.51 $X2=0
+ $Y2=0
cc_325 N_RESET_B_M1002_g N_A_823_25#_c_398_n 0.00151876f $X=3.83 $Y=0.675 $X2=0
+ $Y2=0
cc_326 N_RESET_B_c_360_n N_A_823_25#_c_398_n 0.00672639f $X=3.74 $Y=1.51 $X2=0
+ $Y2=0
cc_327 N_RESET_B_c_359_n N_A_823_25#_c_401_n 0.0438589f $X=3.875 $Y=1.715 $X2=0
+ $Y2=0
cc_328 N_RESET_B_c_360_n N_A_823_25#_c_401_n 6.80985e-19 $X=3.74 $Y=1.51 $X2=0
+ $Y2=0
cc_329 N_RESET_B_c_359_n N_VPWR_c_904_n 0.00681367f $X=3.875 $Y=1.715 $X2=0
+ $Y2=0
cc_330 N_RESET_B_c_359_n N_VPWR_c_905_n 8.47667e-19 $X=3.875 $Y=1.715 $X2=0
+ $Y2=0
cc_331 N_RESET_B_c_359_n N_VPWR_c_911_n 0.0054895f $X=3.875 $Y=1.715 $X2=0 $Y2=0
cc_332 N_RESET_B_c_359_n N_VPWR_c_899_n 0.0103063f $X=3.875 $Y=1.715 $X2=0 $Y2=0
cc_333 N_RESET_B_M1002_g N_VGND_c_1100_n 0.00325573f $X=3.83 $Y=0.675 $X2=0
+ $Y2=0
cc_334 N_RESET_B_M1002_g N_VGND_c_1111_n 0.00565115f $X=3.83 $Y=0.675 $X2=0
+ $Y2=0
cc_335 N_RESET_B_M1002_g N_VGND_c_1113_n 0.0106341f $X=3.83 $Y=0.675 $X2=0 $Y2=0
cc_336 N_A_823_25#_c_403_n N_A_1023_405#_M1000_g 0.00254358f $X=5.73 $Y=2.45
+ $X2=0 $Y2=0
cc_337 N_A_823_25#_c_400_n N_A_1023_405#_c_485_n 0.040103f $X=5.725 $Y=2.275
+ $X2=0 $Y2=0
cc_338 N_A_823_25#_M1000_d N_A_1023_405#_c_486_n 0.00493507f $X=5.495 $Y=2.515
+ $X2=0 $Y2=0
cc_339 N_A_823_25#_c_403_n N_A_1023_405#_c_486_n 0.0144872f $X=5.73 $Y=2.45
+ $X2=0 $Y2=0
cc_340 N_A_823_25#_c_403_n N_A_1023_405#_c_478_n 0.00341005f $X=5.73 $Y=2.45
+ $X2=0 $Y2=0
cc_341 N_A_823_25#_c_400_n N_A_1023_405#_c_478_n 0.0520623f $X=5.725 $Y=2.275
+ $X2=0 $Y2=0
cc_342 N_A_823_25#_c_397_n N_A_1023_405#_c_480_n 0.00430496f $X=5.71 $Y=1.185
+ $X2=0 $Y2=0
cc_343 N_A_823_25#_c_421_n N_A_1023_405#_c_480_n 0.00220334f $X=5.835 $Y=0.805
+ $X2=0 $Y2=0
cc_344 N_A_823_25#_c_399_n N_A_1023_405#_c_480_n 0.0138616f $X=5.71 $Y=1.27
+ $X2=0 $Y2=0
cc_345 N_A_823_25#_c_400_n N_A_1023_405#_c_480_n 0.00720002f $X=5.725 $Y=2.275
+ $X2=0 $Y2=0
cc_346 N_A_823_25#_c_397_n N_A_1023_405#_c_481_n 3.54593e-19 $X=5.71 $Y=1.185
+ $X2=0 $Y2=0
cc_347 N_A_823_25#_c_421_n N_A_1023_405#_c_481_n 0.00149362f $X=5.835 $Y=0.805
+ $X2=0 $Y2=0
cc_348 N_A_823_25#_c_399_n N_A_1023_405#_c_481_n 0.00117674f $X=5.71 $Y=1.27
+ $X2=0 $Y2=0
cc_349 N_A_823_25#_c_400_n N_A_1023_405#_c_481_n 5.92639e-19 $X=5.725 $Y=2.275
+ $X2=0 $Y2=0
cc_350 N_A_823_25#_c_396_n N_A_1023_405#_c_493_n 0.00456783f $X=5.625 $Y=1.27
+ $X2=0 $Y2=0
cc_351 N_A_823_25#_c_400_n N_A_1023_405#_c_493_n 0.00254358f $X=5.725 $Y=2.275
+ $X2=0 $Y2=0
cc_352 N_A_823_25#_c_397_n N_A_1023_405#_c_483_n 0.00304083f $X=5.71 $Y=1.185
+ $X2=0 $Y2=0
cc_353 N_A_823_25#_c_421_n N_A_1023_405#_c_483_n 0.00648177f $X=5.835 $Y=0.805
+ $X2=0 $Y2=0
cc_354 N_A_823_25#_c_421_n N_A_1246_339#_M1024_g 9.90281e-19 $X=5.835 $Y=0.805
+ $X2=0 $Y2=0
cc_355 N_A_823_25#_c_397_n N_A_1246_339#_c_618_n 9.37244e-19 $X=5.71 $Y=1.185
+ $X2=0 $Y2=0
cc_356 N_A_823_25#_c_396_n N_A_1109_21#_M1013_g 0.00952445f $X=5.625 $Y=1.27
+ $X2=0 $Y2=0
cc_357 N_A_823_25#_c_397_n N_A_1109_21#_M1013_g 0.00572356f $X=5.71 $Y=1.185
+ $X2=0 $Y2=0
cc_358 N_A_823_25#_c_421_n N_A_1109_21#_M1013_g 0.00749285f $X=5.835 $Y=0.805
+ $X2=0 $Y2=0
cc_359 N_A_823_25#_c_399_n N_A_1109_21#_M1013_g 0.00185925f $X=5.71 $Y=1.27
+ $X2=0 $Y2=0
cc_360 N_A_823_25#_c_400_n N_A_1109_21#_M1013_g 0.00847959f $X=5.725 $Y=2.275
+ $X2=0 $Y2=0
cc_361 N_A_823_25#_c_421_n N_A_1109_21#_c_740_n 0.00326233f $X=5.835 $Y=0.805
+ $X2=0 $Y2=0
cc_362 N_A_823_25#_c_400_n N_A_1109_21#_M1016_g 0.00597973f $X=5.725 $Y=2.275
+ $X2=0 $Y2=0
cc_363 N_A_823_25#_c_403_n N_A_1109_21#_c_755_n 8.37898e-19 $X=5.73 $Y=2.45
+ $X2=0 $Y2=0
cc_364 N_A_823_25#_c_400_n N_A_1109_21#_c_755_n 0.0139859f $X=5.725 $Y=2.275
+ $X2=0 $Y2=0
cc_365 N_A_823_25#_M1022_g N_VPWR_c_905_n 0.0162433f $X=4.305 $Y=2.465 $X2=0
+ $Y2=0
cc_366 N_A_823_25#_M1022_g N_VPWR_c_911_n 0.00486043f $X=4.305 $Y=2.465 $X2=0
+ $Y2=0
cc_367 N_A_823_25#_M1022_g N_VPWR_c_899_n 0.0082726f $X=4.305 $Y=2.465 $X2=0
+ $Y2=0
cc_368 N_A_823_25#_c_394_n N_VGND_c_1101_n 0.00327939f $X=4.19 $Y=1.205 $X2=0
+ $Y2=0
cc_369 N_A_823_25#_c_396_n N_VGND_c_1101_n 0.0206023f $X=5.625 $Y=1.27 $X2=0
+ $Y2=0
cc_370 N_A_823_25#_c_397_n N_VGND_c_1101_n 5.21178e-19 $X=5.71 $Y=1.185 $X2=0
+ $Y2=0
cc_371 N_A_823_25#_c_421_n N_VGND_c_1101_n 0.0115694f $X=5.835 $Y=0.805 $X2=0
+ $Y2=0
cc_372 N_A_823_25#_c_421_n N_VGND_c_1102_n 0.00810097f $X=5.835 $Y=0.805 $X2=0
+ $Y2=0
cc_373 N_A_823_25#_c_421_n N_VGND_c_1104_n 0.00566949f $X=5.835 $Y=0.805 $X2=0
+ $Y2=0
cc_374 N_A_823_25#_c_394_n N_VGND_c_1111_n 0.00529818f $X=4.19 $Y=1.205 $X2=0
+ $Y2=0
cc_375 N_A_823_25#_c_394_n N_VGND_c_1113_n 0.00716236f $X=4.19 $Y=1.205 $X2=0
+ $Y2=0
cc_376 N_A_823_25#_c_421_n N_VGND_c_1113_n 0.00931973f $X=5.835 $Y=0.805 $X2=0
+ $Y2=0
cc_377 N_A_1023_405#_c_491_n N_A_1246_339#_M1017_d 0.00339207f $X=7.615 $Y=2.81
+ $X2=0 $Y2=0
cc_378 N_A_1023_405#_c_486_n N_A_1246_339#_M1023_g 0.00125403f $X=5.995 $Y=2.87
+ $X2=0 $Y2=0
cc_379 N_A_1023_405#_c_521_p N_A_1246_339#_M1023_g 0.00438167f $X=6.08 $Y=2.785
+ $X2=0 $Y2=0
cc_380 N_A_1023_405#_c_522_p N_A_1246_339#_M1023_g 0.0156754f $X=6.865 $Y=2.44
+ $X2=0 $Y2=0
cc_381 N_A_1023_405#_c_523_p N_A_1246_339#_M1023_g 0.00244055f $X=6.95 $Y=2.81
+ $X2=0 $Y2=0
cc_382 N_A_1023_405#_c_489_n N_A_1246_339#_M1023_g 3.21961e-19 $X=7.035 $Y=2.895
+ $X2=0 $Y2=0
cc_383 N_A_1023_405#_c_478_n N_A_1246_339#_M1024_g 0.00122023f $X=6.08 $Y=2.355
+ $X2=0 $Y2=0
cc_384 N_A_1023_405#_c_480_n N_A_1246_339#_M1024_g 3.0392e-19 $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_385 N_A_1023_405#_c_481_n N_A_1246_339#_M1024_g 0.0203545f $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_386 N_A_1023_405#_c_483_n N_A_1246_339#_M1024_g 0.0248239f $X=6.07 $Y=1.125
+ $X2=0 $Y2=0
cc_387 N_A_1023_405#_c_522_p N_A_1246_339#_c_616_n 0.0107621f $X=6.865 $Y=2.44
+ $X2=0 $Y2=0
cc_388 N_A_1023_405#_c_480_n N_A_1246_339#_c_616_n 0.0568025f $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_389 N_A_1023_405#_c_481_n N_A_1246_339#_c_616_n 0.00116911f $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_390 N_A_1023_405#_c_480_n N_A_1246_339#_c_618_n 0.0118229f $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_391 N_A_1023_405#_c_481_n N_A_1246_339#_c_618_n 0.00102453f $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_392 N_A_1023_405#_c_483_n N_A_1246_339#_c_618_n 2.78513e-19 $X=6.07 $Y=1.125
+ $X2=0 $Y2=0
cc_393 N_A_1023_405#_c_479_n N_A_1246_339#_c_619_n 0.0238756f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_394 N_A_1023_405#_c_479_n N_A_1246_339#_c_620_n 0.0137878f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_395 N_A_1023_405#_c_522_p N_A_1246_339#_c_625_n 0.013649f $X=6.865 $Y=2.44
+ $X2=0 $Y2=0
cc_396 N_A_1023_405#_c_523_p N_A_1246_339#_c_625_n 0.00823307f $X=6.95 $Y=2.81
+ $X2=0 $Y2=0
cc_397 N_A_1023_405#_c_491_n N_A_1246_339#_c_625_n 0.0174686f $X=7.615 $Y=2.81
+ $X2=0 $Y2=0
cc_398 N_A_1023_405#_c_479_n N_A_1246_339#_c_621_n 0.099592f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_399 N_A_1023_405#_c_478_n N_A_1246_339#_c_627_n 0.00842476f $X=6.08 $Y=2.355
+ $X2=0 $Y2=0
cc_400 N_A_1023_405#_c_522_p N_A_1246_339#_c_627_n 0.00113211f $X=6.865 $Y=2.44
+ $X2=0 $Y2=0
cc_401 N_A_1023_405#_c_481_n N_A_1246_339#_c_627_n 3.49631e-19 $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_402 N_A_1023_405#_c_479_n N_D_M1026_g 0.00104176f $X=7.7 $Y=2.64 $X2=0 $Y2=0
cc_403 N_A_1023_405#_c_482_n N_D_M1026_g 6.51767e-19 $X=7.855 $Y=0.445 $X2=0
+ $Y2=0
cc_404 N_A_1023_405#_c_522_p N_D_M1017_g 0.00612719f $X=6.865 $Y=2.44 $X2=0
+ $Y2=0
cc_405 N_A_1023_405#_c_523_p N_D_M1017_g 0.00858822f $X=6.95 $Y=2.81 $X2=0 $Y2=0
cc_406 N_A_1023_405#_c_489_n N_D_M1017_g 0.00324565f $X=7.035 $Y=2.895 $X2=0
+ $Y2=0
cc_407 N_A_1023_405#_c_491_n N_D_M1017_g 0.0112559f $X=7.615 $Y=2.81 $X2=0 $Y2=0
cc_408 N_A_1023_405#_c_492_n N_D_M1017_g 0.00249111f $X=7.925 $Y=2.805 $X2=0
+ $Y2=0
cc_409 N_A_1023_405#_c_522_p N_D_c_697_n 9.08851e-19 $X=6.865 $Y=2.44 $X2=0
+ $Y2=0
cc_410 N_A_1023_405#_c_478_n D 0.00343001f $X=6.08 $Y=2.355 $X2=0 $Y2=0
cc_411 N_A_1023_405#_c_522_p D 0.0169726f $X=6.865 $Y=2.44 $X2=0 $Y2=0
cc_412 N_A_1023_405#_c_478_n N_A_1109_21#_M1013_g 6.51379e-19 $X=6.08 $Y=2.355
+ $X2=0 $Y2=0
cc_413 N_A_1023_405#_c_480_n N_A_1109_21#_M1013_g 3.15586e-19 $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_414 N_A_1023_405#_c_481_n N_A_1109_21#_M1013_g 0.0203711f $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_415 N_A_1023_405#_c_483_n N_A_1109_21#_M1013_g 0.0124302f $X=6.07 $Y=1.125
+ $X2=0 $Y2=0
cc_416 N_A_1023_405#_c_483_n N_A_1109_21#_c_740_n 0.0103123f $X=6.07 $Y=1.125
+ $X2=0 $Y2=0
cc_417 N_A_1023_405#_c_485_n N_A_1109_21#_M1016_g 6.67791e-19 $X=5.28 $Y=2.19
+ $X2=0 $Y2=0
cc_418 N_A_1023_405#_c_486_n N_A_1109_21#_M1016_g 0.0127992f $X=5.995 $Y=2.87
+ $X2=0 $Y2=0
cc_419 N_A_1023_405#_c_478_n N_A_1109_21#_M1016_g 0.00844455f $X=6.08 $Y=2.355
+ $X2=0 $Y2=0
cc_420 N_A_1023_405#_c_521_p N_A_1109_21#_M1016_g 0.00544109f $X=6.08 $Y=2.785
+ $X2=0 $Y2=0
cc_421 N_A_1023_405#_c_563_p N_A_1109_21#_M1016_g 0.00328964f $X=6.08 $Y=2.44
+ $X2=0 $Y2=0
cc_422 N_A_1023_405#_c_493_n N_A_1109_21#_M1016_g 0.0243036f $X=5.42 $Y=2.19
+ $X2=0 $Y2=0
cc_423 N_A_1023_405#_c_479_n N_A_1109_21#_c_742_n 0.00390444f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_424 N_A_1023_405#_c_482_n N_A_1109_21#_c_742_n 0.0160905f $X=7.855 $Y=0.445
+ $X2=0 $Y2=0
cc_425 N_A_1023_405#_c_479_n N_A_1109_21#_c_743_n 0.00867885f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_426 N_A_1023_405#_c_482_n N_A_1109_21#_c_743_n 0.00476686f $X=7.855 $Y=0.445
+ $X2=0 $Y2=0
cc_427 N_A_1023_405#_c_479_n N_A_1109_21#_c_744_n 0.00312057f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_428 N_A_1023_405#_c_479_n N_A_1109_21#_c_745_n 0.00302969f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_429 N_A_1023_405#_c_479_n N_A_1109_21#_M1004_g 0.0058906f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_430 N_A_1023_405#_c_478_n N_A_1109_21#_c_755_n 0.00398059f $X=6.08 $Y=2.355
+ $X2=0 $Y2=0
cc_431 N_A_1023_405#_c_480_n N_A_1109_21#_c_755_n 2.20068e-19 $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_432 N_A_1023_405#_c_481_n N_A_1109_21#_c_755_n 0.00730721f $X=6.07 $Y=1.29
+ $X2=0 $Y2=0
cc_433 N_A_1023_405#_c_479_n N_A_1109_21#_c_746_n 0.0144433f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_434 N_A_1023_405#_c_492_n N_A_1109_21#_c_757_n 0.00274508f $X=7.925 $Y=2.805
+ $X2=0 $Y2=0
cc_435 N_A_1023_405#_c_479_n N_A_1109_21#_c_748_n 0.0514141f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_436 N_A_1023_405#_c_479_n N_A_1109_21#_c_749_n 0.00993926f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_437 N_A_1023_405#_M1004_s N_A_1109_21#_c_761_n 0.00119091f $X=7.8 $Y=2.415
+ $X2=0 $Y2=0
cc_438 N_A_1023_405#_c_479_n N_A_1109_21#_c_761_n 0.0142597f $X=7.7 $Y=2.64
+ $X2=0 $Y2=0
cc_439 N_A_1023_405#_c_492_n N_A_1109_21#_c_761_n 0.00441513f $X=7.925 $Y=2.805
+ $X2=0 $Y2=0
cc_440 N_A_1023_405#_c_479_n GATE 0.0289697f $X=7.7 $Y=2.64 $X2=0 $Y2=0
cc_441 N_A_1023_405#_c_522_p N_VPWR_M1023_d 0.018514f $X=6.865 $Y=2.44 $X2=0
+ $Y2=0
cc_442 N_A_1023_405#_c_523_p N_VPWR_M1023_d 0.0036436f $X=6.95 $Y=2.81 $X2=0
+ $Y2=0
cc_443 N_A_1023_405#_c_489_n N_VPWR_M1023_d 0.00122627f $X=7.035 $Y=2.895 $X2=0
+ $Y2=0
cc_444 N_A_1023_405#_c_485_n N_VPWR_c_905_n 0.0297119f $X=5.28 $Y=2.19 $X2=0
+ $Y2=0
cc_445 N_A_1023_405#_c_487_n N_VPWR_c_905_n 0.00734033f $X=5.445 $Y=2.87 $X2=0
+ $Y2=0
cc_446 N_A_1023_405#_c_486_n N_VPWR_c_906_n 0.0129433f $X=5.995 $Y=2.87 $X2=0
+ $Y2=0
cc_447 N_A_1023_405#_c_521_p N_VPWR_c_906_n 0.00607901f $X=6.08 $Y=2.785 $X2=0
+ $Y2=0
cc_448 N_A_1023_405#_c_522_p N_VPWR_c_906_n 0.0222331f $X=6.865 $Y=2.44 $X2=0
+ $Y2=0
cc_449 N_A_1023_405#_c_523_p N_VPWR_c_906_n 0.00877273f $X=6.95 $Y=2.81 $X2=0
+ $Y2=0
cc_450 N_A_1023_405#_c_489_n N_VPWR_c_906_n 0.0146568f $X=7.035 $Y=2.895 $X2=0
+ $Y2=0
cc_451 N_A_1023_405#_M1000_g N_VPWR_c_912_n 0.0039943f $X=5.42 $Y=2.725 $X2=0
+ $Y2=0
cc_452 N_A_1023_405#_c_486_n N_VPWR_c_912_n 0.0265265f $X=5.995 $Y=2.87 $X2=0
+ $Y2=0
cc_453 N_A_1023_405#_c_487_n N_VPWR_c_912_n 0.0130756f $X=5.445 $Y=2.87 $X2=0
+ $Y2=0
cc_454 N_A_1023_405#_c_489_n N_VPWR_c_913_n 0.00740612f $X=7.035 $Y=2.895 $X2=0
+ $Y2=0
cc_455 N_A_1023_405#_c_491_n N_VPWR_c_913_n 0.0397642f $X=7.615 $Y=2.81 $X2=0
+ $Y2=0
cc_456 N_A_1023_405#_M1000_g N_VPWR_c_899_n 0.00537853f $X=5.42 $Y=2.725 $X2=0
+ $Y2=0
cc_457 N_A_1023_405#_c_486_n N_VPWR_c_899_n 0.0251132f $X=5.995 $Y=2.87 $X2=0
+ $Y2=0
cc_458 N_A_1023_405#_c_487_n N_VPWR_c_899_n 0.0119105f $X=5.445 $Y=2.87 $X2=0
+ $Y2=0
cc_459 N_A_1023_405#_c_522_p N_VPWR_c_899_n 0.0135731f $X=6.865 $Y=2.44 $X2=0
+ $Y2=0
cc_460 N_A_1023_405#_c_489_n N_VPWR_c_899_n 0.00622418f $X=7.035 $Y=2.895 $X2=0
+ $Y2=0
cc_461 N_A_1023_405#_c_491_n N_VPWR_c_899_n 0.0350291f $X=7.615 $Y=2.81 $X2=0
+ $Y2=0
cc_462 N_A_1023_405#_c_485_n A_981_503# 0.00411955f $X=5.28 $Y=2.19 $X2=-0.19
+ $Y2=-0.245
cc_463 N_A_1023_405#_c_487_n A_981_503# 0.00237995f $X=5.445 $Y=2.87 $X2=-0.19
+ $Y2=-0.245
cc_464 N_A_1023_405#_c_486_n A_1204_459# 0.00132782f $X=5.995 $Y=2.87 $X2=-0.19
+ $Y2=-0.245
cc_465 N_A_1023_405#_c_478_n A_1204_459# 6.49906e-19 $X=6.08 $Y=2.355 $X2=-0.19
+ $Y2=-0.245
cc_466 N_A_1023_405#_c_521_p A_1204_459# 0.00261797f $X=6.08 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_467 N_A_1023_405#_c_522_p A_1204_459# 4.03595e-19 $X=6.865 $Y=2.44 $X2=-0.19
+ $Y2=-0.245
cc_468 N_A_1023_405#_c_483_n N_VGND_c_1102_n 0.00171767f $X=6.07 $Y=1.125 $X2=0
+ $Y2=0
cc_469 N_A_1023_405#_c_482_n N_VGND_c_1106_n 0.0197797f $X=7.855 $Y=0.445 $X2=0
+ $Y2=0
cc_470 N_A_1023_405#_M1010_s N_VGND_c_1113_n 0.00266218f $X=7.73 $Y=0.235 $X2=0
+ $Y2=0
cc_471 N_A_1023_405#_c_482_n N_VGND_c_1113_n 0.0135505f $X=7.855 $Y=0.445 $X2=0
+ $Y2=0
cc_472 N_A_1023_405#_c_483_n N_VGND_c_1113_n 9.39239e-19 $X=6.07 $Y=1.125 $X2=0
+ $Y2=0
cc_473 N_A_1246_339#_M1024_g N_D_M1026_g 0.0262509f $X=6.52 $Y=0.805 $X2=0 $Y2=0
cc_474 N_A_1246_339#_c_616_n N_D_M1026_g 7.28012e-19 $X=6.43 $Y=1.86 $X2=0 $Y2=0
cc_475 N_A_1246_339#_c_617_n N_D_M1026_g 0.0157773f $X=7.07 $Y=1.185 $X2=0 $Y2=0
cc_476 N_A_1246_339#_c_619_n N_D_M1026_g 0.00375589f $X=7.165 $Y=0.805 $X2=0
+ $Y2=0
cc_477 N_A_1246_339#_c_621_n N_D_M1026_g 0.00392898f $X=7.32 $Y=2.3 $X2=0 $Y2=0
cc_478 N_A_1246_339#_M1023_g N_D_M1017_g 0.0128942f $X=6.305 $Y=2.615 $X2=0
+ $Y2=0
cc_479 N_A_1246_339#_c_621_n N_D_M1017_g 0.00618812f $X=7.32 $Y=2.3 $X2=0 $Y2=0
cc_480 N_A_1246_339#_c_627_n N_D_c_692_n 0.0148264f $X=6.52 $Y=1.86 $X2=0 $Y2=0
cc_481 N_A_1246_339#_M1023_g N_D_c_697_n 0.00202654f $X=6.305 $Y=2.615 $X2=0
+ $Y2=0
cc_482 N_A_1246_339#_M1023_g D 9.14515e-19 $X=6.305 $Y=2.615 $X2=0 $Y2=0
cc_483 N_A_1246_339#_M1024_g D 0.0033535f $X=6.52 $Y=0.805 $X2=0 $Y2=0
cc_484 N_A_1246_339#_c_616_n D 0.044695f $X=6.43 $Y=1.86 $X2=0 $Y2=0
cc_485 N_A_1246_339#_c_617_n D 0.0229751f $X=7.07 $Y=1.185 $X2=0 $Y2=0
cc_486 N_A_1246_339#_c_620_n D 0.0020369f $X=7.252 $Y=1.185 $X2=0 $Y2=0
cc_487 N_A_1246_339#_c_621_n D 0.0509893f $X=7.32 $Y=2.3 $X2=0 $Y2=0
cc_488 N_A_1246_339#_M1024_g N_D_c_694_n 0.0148264f $X=6.52 $Y=0.805 $X2=0 $Y2=0
cc_489 N_A_1246_339#_c_616_n N_D_c_694_n 6.36363e-19 $X=6.43 $Y=1.86 $X2=0 $Y2=0
cc_490 N_A_1246_339#_c_617_n N_D_c_694_n 5.82132e-19 $X=7.07 $Y=1.185 $X2=0
+ $Y2=0
cc_491 N_A_1246_339#_c_620_n N_D_c_694_n 0.00352194f $X=7.252 $Y=1.185 $X2=0
+ $Y2=0
cc_492 N_A_1246_339#_c_621_n N_D_c_694_n 0.00993926f $X=7.32 $Y=2.3 $X2=0 $Y2=0
cc_493 N_A_1246_339#_M1024_g N_A_1109_21#_c_740_n 0.0103107f $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_494 N_A_1246_339#_c_619_n N_A_1109_21#_c_740_n 0.00488616f $X=7.165 $Y=0.805
+ $X2=0 $Y2=0
cc_495 N_A_1246_339#_M1023_g N_A_1109_21#_M1016_g 0.0411796f $X=6.305 $Y=2.615
+ $X2=0 $Y2=0
cc_496 N_A_1246_339#_c_619_n N_A_1109_21#_c_742_n 0.00280408f $X=7.165 $Y=0.805
+ $X2=0 $Y2=0
cc_497 N_A_1246_339#_M1024_g N_A_1109_21#_c_755_n 4.3105e-19 $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_498 N_A_1246_339#_c_616_n N_A_1109_21#_c_755_n 2.6803e-19 $X=6.43 $Y=1.86
+ $X2=0 $Y2=0
cc_499 N_A_1246_339#_c_627_n N_A_1109_21#_c_755_n 0.0411796f $X=6.52 $Y=1.86
+ $X2=0 $Y2=0
cc_500 N_A_1246_339#_M1023_g N_VPWR_c_906_n 0.00754725f $X=6.305 $Y=2.615 $X2=0
+ $Y2=0
cc_501 N_A_1246_339#_M1023_g N_VPWR_c_912_n 0.00465077f $X=6.305 $Y=2.615 $X2=0
+ $Y2=0
cc_502 N_A_1246_339#_M1023_g N_VPWR_c_899_n 0.00451796f $X=6.305 $Y=2.615 $X2=0
+ $Y2=0
cc_503 N_A_1246_339#_M1024_g N_VGND_c_1102_n 0.0108613f $X=6.52 $Y=0.805 $X2=0
+ $Y2=0
cc_504 N_A_1246_339#_c_617_n N_VGND_c_1102_n 0.0197848f $X=7.07 $Y=1.185 $X2=0
+ $Y2=0
cc_505 N_A_1246_339#_c_618_n N_VGND_c_1102_n 0.0019893f $X=6.595 $Y=1.185 $X2=0
+ $Y2=0
cc_506 N_A_1246_339#_c_619_n N_VGND_c_1106_n 0.00483152f $X=7.165 $Y=0.805 $X2=0
+ $Y2=0
cc_507 N_A_1246_339#_M1024_g N_VGND_c_1113_n 7.88961e-19 $X=6.52 $Y=0.805 $X2=0
+ $Y2=0
cc_508 N_A_1246_339#_c_619_n N_VGND_c_1113_n 0.00676558f $X=7.165 $Y=0.805 $X2=0
+ $Y2=0
cc_509 N_D_M1026_g N_A_1109_21#_c_740_n 0.0103107f $X=6.95 $Y=0.805 $X2=0 $Y2=0
cc_510 N_D_M1026_g N_A_1109_21#_c_742_n 0.00591456f $X=6.95 $Y=0.805 $X2=0 $Y2=0
cc_511 N_D_c_692_n N_A_1109_21#_c_756_n 0.00156052f $X=7 $Y=1.955 $X2=0 $Y2=0
cc_512 N_D_c_697_n N_A_1109_21#_c_757_n 0.00156052f $X=7 $Y=2.12 $X2=0 $Y2=0
cc_513 N_D_c_694_n N_A_1109_21#_c_749_n 0.00156052f $X=7 $Y=1.615 $X2=0 $Y2=0
cc_514 N_D_M1017_g N_VPWR_c_906_n 0.00287474f $X=7.065 $Y=2.615 $X2=0 $Y2=0
cc_515 N_D_M1017_g N_VPWR_c_913_n 0.00396326f $X=7.065 $Y=2.615 $X2=0 $Y2=0
cc_516 N_D_M1017_g N_VPWR_c_899_n 0.00537853f $X=7.065 $Y=2.615 $X2=0 $Y2=0
cc_517 N_D_M1026_g N_VGND_c_1102_n 0.00899513f $X=6.95 $Y=0.805 $X2=0 $Y2=0
cc_518 N_D_M1026_g N_VGND_c_1113_n 7.88961e-19 $X=6.95 $Y=0.805 $X2=0 $Y2=0
cc_519 N_A_1109_21#_c_745_n N_GATE_M1020_g 0.0147193f $X=8.07 $Y=0.765 $X2=0
+ $Y2=0
cc_520 N_A_1109_21#_c_750_n N_GATE_M1020_g 0.00513797f $X=8.935 $Y=2.3 $X2=0
+ $Y2=0
cc_521 N_A_1109_21#_c_746_n N_GATE_M1008_g 0.00220447f $X=8.05 $Y=1.585 $X2=0
+ $Y2=0
cc_522 N_A_1109_21#_c_748_n N_GATE_M1008_g 0.00136212f $X=8.05 $Y=1.75 $X2=0
+ $Y2=0
cc_523 N_A_1109_21#_c_749_n N_GATE_M1008_g 0.052909f $X=8.05 $Y=1.75 $X2=0 $Y2=0
cc_524 N_A_1109_21#_c_760_n N_GATE_M1008_g 0.0121599f $X=8.69 $Y=2.385 $X2=0
+ $Y2=0
cc_525 N_A_1109_21#_c_762_n N_GATE_M1008_g 2.23531e-19 $X=8.79 $Y=2.56 $X2=0
+ $Y2=0
cc_526 N_A_1109_21#_c_750_n N_GATE_M1008_g 0.00974412f $X=8.935 $Y=2.3 $X2=0
+ $Y2=0
cc_527 N_A_1109_21#_c_746_n N_GATE_c_866_n 0.0147193f $X=8.05 $Y=1.585 $X2=0
+ $Y2=0
cc_528 N_A_1109_21#_c_747_n GATE 0.00869681f $X=8.07 $Y=0.84 $X2=0 $Y2=0
cc_529 N_A_1109_21#_c_748_n GATE 0.0416374f $X=8.05 $Y=1.75 $X2=0 $Y2=0
cc_530 N_A_1109_21#_c_749_n GATE 0.00422872f $X=8.05 $Y=1.75 $X2=0 $Y2=0
cc_531 N_A_1109_21#_c_760_n GATE 0.0298387f $X=8.69 $Y=2.385 $X2=0 $Y2=0
cc_532 N_A_1109_21#_c_750_n GATE 0.105561f $X=8.935 $Y=2.3 $X2=0 $Y2=0
cc_533 N_A_1109_21#_c_751_n GATE 0.00558853f $X=8.935 $Y=0.445 $X2=0 $Y2=0
cc_534 N_A_1109_21#_c_747_n N_GATE_c_869_n 0.0147193f $X=8.07 $Y=0.84 $X2=0
+ $Y2=0
cc_535 N_A_1109_21#_c_750_n N_GATE_c_869_n 0.0164925f $X=8.935 $Y=2.3 $X2=0
+ $Y2=0
cc_536 N_A_1109_21#_c_751_n N_GATE_c_869_n 0.00378778f $X=8.935 $Y=0.445 $X2=0
+ $Y2=0
cc_537 N_A_1109_21#_c_760_n N_VPWR_M1004_d 0.00174317f $X=8.69 $Y=2.385 $X2=0
+ $Y2=0
cc_538 N_A_1109_21#_M1016_g N_VPWR_c_906_n 7.62214e-19 $X=5.945 $Y=2.615 $X2=0
+ $Y2=0
cc_539 N_A_1109_21#_M1004_g N_VPWR_c_907_n 0.0137677f $X=8.14 $Y=2.735 $X2=0
+ $Y2=0
cc_540 N_A_1109_21#_c_760_n N_VPWR_c_907_n 0.0167297f $X=8.69 $Y=2.385 $X2=0
+ $Y2=0
cc_541 N_A_1109_21#_c_762_n N_VPWR_c_907_n 0.0163223f $X=8.79 $Y=2.56 $X2=0
+ $Y2=0
cc_542 N_A_1109_21#_M1016_g N_VPWR_c_912_n 0.00399493f $X=5.945 $Y=2.615 $X2=0
+ $Y2=0
cc_543 N_A_1109_21#_M1004_g N_VPWR_c_913_n 0.00452967f $X=8.14 $Y=2.735 $X2=0
+ $Y2=0
cc_544 N_A_1109_21#_c_762_n N_VPWR_c_914_n 0.0224523f $X=8.79 $Y=2.56 $X2=0
+ $Y2=0
cc_545 N_A_1109_21#_M1016_g N_VPWR_c_899_n 0.00537853f $X=5.945 $Y=2.615 $X2=0
+ $Y2=0
cc_546 N_A_1109_21#_M1004_g N_VPWR_c_899_n 0.00545486f $X=8.14 $Y=2.735 $X2=0
+ $Y2=0
cc_547 N_A_1109_21#_c_760_n N_VPWR_c_899_n 0.00736386f $X=8.69 $Y=2.385 $X2=0
+ $Y2=0
cc_548 N_A_1109_21#_c_761_n N_VPWR_c_899_n 0.00401925f $X=8.135 $Y=2.385 $X2=0
+ $Y2=0
cc_549 N_A_1109_21#_c_762_n N_VPWR_c_899_n 0.0128848f $X=8.79 $Y=2.56 $X2=0
+ $Y2=0
cc_550 N_A_1109_21#_M1013_g N_VGND_c_1101_n 0.00175674f $X=5.62 $Y=0.805 $X2=0
+ $Y2=0
cc_551 N_A_1109_21#_c_741_n N_VGND_c_1101_n 0.0106942f $X=5.695 $Y=0.18 $X2=0
+ $Y2=0
cc_552 N_A_1109_21#_c_740_n N_VGND_c_1102_n 0.0253184f $X=7.505 $Y=0.18 $X2=0
+ $Y2=0
cc_553 N_A_1109_21#_c_742_n N_VGND_c_1102_n 0.0057705f $X=7.58 $Y=0.765 $X2=0
+ $Y2=0
cc_554 N_A_1109_21#_c_745_n N_VGND_c_1103_n 0.00319852f $X=8.07 $Y=0.765 $X2=0
+ $Y2=0
cc_555 N_A_1109_21#_c_741_n N_VGND_c_1104_n 0.0330478f $X=5.695 $Y=0.18 $X2=0
+ $Y2=0
cc_556 N_A_1109_21#_c_740_n N_VGND_c_1106_n 0.0241663f $X=7.505 $Y=0.18 $X2=0
+ $Y2=0
cc_557 N_A_1109_21#_c_745_n N_VGND_c_1106_n 0.00585385f $X=8.07 $Y=0.765 $X2=0
+ $Y2=0
cc_558 N_A_1109_21#_c_751_n N_VGND_c_1112_n 0.0241407f $X=8.935 $Y=0.445 $X2=0
+ $Y2=0
cc_559 N_A_1109_21#_M1020_d N_VGND_c_1113_n 0.00222632f $X=8.575 $Y=0.235 $X2=0
+ $Y2=0
cc_560 N_A_1109_21#_c_740_n N_VGND_c_1113_n 0.0659465f $X=7.505 $Y=0.18 $X2=0
+ $Y2=0
cc_561 N_A_1109_21#_c_741_n N_VGND_c_1113_n 0.00929682f $X=5.695 $Y=0.18 $X2=0
+ $Y2=0
cc_562 N_A_1109_21#_c_745_n N_VGND_c_1113_n 0.0109106f $X=8.07 $Y=0.765 $X2=0
+ $Y2=0
cc_563 N_A_1109_21#_c_751_n N_VGND_c_1113_n 0.0165585f $X=8.935 $Y=0.445 $X2=0
+ $Y2=0
cc_564 N_GATE_M1008_g N_VPWR_c_907_n 0.0109737f $X=8.57 $Y=2.735 $X2=0 $Y2=0
cc_565 N_GATE_M1008_g N_VPWR_c_914_n 0.00452967f $X=8.57 $Y=2.735 $X2=0 $Y2=0
cc_566 N_GATE_M1008_g N_VPWR_c_899_n 0.00522258f $X=8.57 $Y=2.735 $X2=0 $Y2=0
cc_567 N_GATE_M1020_g N_VGND_c_1103_n 0.00316751f $X=8.5 $Y=0.445 $X2=0 $Y2=0
cc_568 GATE N_VGND_c_1103_n 0.00755763f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_569 N_GATE_M1020_g N_VGND_c_1112_n 0.00585385f $X=8.5 $Y=0.445 $X2=0 $Y2=0
cc_570 N_GATE_M1020_g N_VGND_c_1113_n 0.00728923f $X=8.5 $Y=0.445 $X2=0 $Y2=0
cc_571 GATE N_VGND_c_1113_n 0.00651156f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_572 N_VPWR_c_899_n N_Q_N_M1006_s 0.00262367f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_573 N_VPWR_c_901_n N_Q_N_c_1017_n 0.00154413f $X=0.26 $Y=1.98 $X2=0 $Y2=0
cc_574 N_VPWR_c_902_n N_Q_N_c_1017_n 0.00154413f $X=1.125 $Y=1.98 $X2=0 $Y2=0
cc_575 N_VPWR_c_908_n N_Q_N_c_1017_n 0.0156425f $X=1 $Y=3.33 $X2=0 $Y2=0
cc_576 N_VPWR_c_899_n N_Q_N_c_1017_n 0.0106136f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_577 N_VPWR_c_899_n N_Q_M1001_d 0.00238674f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_578 N_VPWR_M1021_d N_Q_c_1035_n 0.00811761f $X=2.39 $Y=1.835 $X2=0 $Y2=0
cc_579 N_VPWR_M1021_d Q 0.00158083f $X=2.39 $Y=1.835 $X2=0 $Y2=0
cc_580 N_VPWR_c_903_n Q 0.0127621f $X=2.625 $Y=2.79 $X2=0 $Y2=0
cc_581 N_VPWR_c_899_n Q 0.00154744f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_582 N_VPWR_c_902_n N_Q_c_1039_n 0.0122827f $X=1.125 $Y=1.98 $X2=0 $Y2=0
cc_583 N_VPWR_c_899_n N_Q_c_1039_n 0.0314425f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_584 N_VPWR_M1021_d N_Q_c_1065_n 0.00411357f $X=2.39 $Y=1.835 $X2=0 $Y2=0
cc_585 N_VPWR_c_903_n N_Q_c_1065_n 0.0102114f $X=2.625 $Y=2.79 $X2=0 $Y2=0
cc_586 N_VPWR_c_899_n N_Q_c_1065_n 0.00553076f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_587 N_VPWR_c_910_n N_Q_c_1067_n 0.0163977f $X=3.415 $Y=3.33 $X2=0 $Y2=0
cc_588 N_VPWR_c_899_n N_Q_c_1067_n 0.010625f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_589 N_Q_N_c_1017_n N_VGND_c_1097_n 0.00154413f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_590 N_Q_N_c_1017_n N_VGND_c_1098_n 0.0296698f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_591 N_Q_N_c_1017_n N_VGND_c_1108_n 0.0154684f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_592 N_Q_N_M1007_d N_VGND_c_1113_n 0.00240953f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_593 N_Q_N_c_1017_n N_VGND_c_1113_n 0.0106136f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_594 N_Q_c_1035_n N_VGND_M1009_d 0.00738081f $X=2.52 $Y=2.26 $X2=0 $Y2=0
cc_595 N_Q_c_1053_n N_VGND_M1009_d 0.00380679f $X=2.91 $Y=0.745 $X2=0 $Y2=0
cc_596 N_Q_c_1043_n N_VGND_M1009_d 0.00555592f $X=2.605 $Y=0.745 $X2=0 $Y2=0
cc_597 N_Q_c_1053_n N_VGND_c_1099_n 0.00854861f $X=2.91 $Y=0.745 $X2=0 $Y2=0
cc_598 N_Q_c_1043_n N_VGND_c_1099_n 0.0130251f $X=2.605 $Y=0.745 $X2=0 $Y2=0
cc_599 N_Q_c_1053_n N_VGND_c_1110_n 0.00245154f $X=2.91 $Y=0.745 $X2=0 $Y2=0
cc_600 N_Q_c_1036_n N_VGND_c_1110_n 0.0187529f $X=3.075 $Y=0.39 $X2=0 $Y2=0
cc_601 N_Q_c_1053_n N_VGND_c_1113_n 0.0050475f $X=2.91 $Y=0.745 $X2=0 $Y2=0
cc_602 N_Q_c_1043_n N_VGND_c_1113_n 8.80196e-19 $X=2.605 $Y=0.745 $X2=0 $Y2=0
cc_603 N_Q_c_1036_n N_VGND_c_1113_n 0.0124602f $X=3.075 $Y=0.39 $X2=0 $Y2=0
