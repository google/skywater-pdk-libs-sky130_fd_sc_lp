# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__nand2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.415000 3.770000 1.760000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.425000 2.245000 1.760000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.881600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.930000 3.770000 2.140000 ;
        RECT 0.635000 2.140000 0.965000 3.055000 ;
        RECT 1.635000 2.140000 1.825000 3.055000 ;
        RECT 2.425000 0.615000 2.755000 1.075000 ;
        RECT 2.425000 1.075000 3.775000 1.245000 ;
        RECT 2.425000 1.245000 2.755000 1.930000 ;
        RECT 2.495000 2.140000 2.750000 3.055000 ;
        RECT 3.420000 2.140000 3.770000 3.055000 ;
        RECT 3.435000 0.605000 3.775000 1.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.125000  1.805000 0.465000 3.245000 ;
      RECT 0.285000  0.305000 0.535000 1.085000 ;
      RECT 0.285000  1.085000 2.255000 1.255000 ;
      RECT 0.705000  0.085000 1.035000 0.915000 ;
      RECT 1.135000  2.310000 1.465000 3.245000 ;
      RECT 1.205000  0.305000 1.395000 1.085000 ;
      RECT 1.565000  0.085000 1.895000 0.915000 ;
      RECT 1.995000  2.310000 2.325000 3.245000 ;
      RECT 2.065000  0.265000 4.205000 0.435000 ;
      RECT 2.065000  0.435000 2.255000 1.085000 ;
      RECT 2.920000  2.310000 3.250000 3.245000 ;
      RECT 2.935000  0.435000 3.265000 0.905000 ;
      RECT 3.940000  1.815000 4.205000 3.245000 ;
      RECT 3.945000  0.435000 4.205000 1.185000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__nand2_4
END LIBRARY
