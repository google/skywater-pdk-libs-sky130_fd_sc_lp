* File: sky130_fd_sc_lp__a31o_1.spice
* Created: Wed Sep  2 09:26:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a31o_1.pex.spice"
.subckt sky130_fd_sc_lp__a31o_1  VNB VPB A3 A2 A1 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_80_21#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2709 AS=0.2226 PD=1.485 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1002 A_269_47# N_A3_M1002_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.2709 PD=1.08 PS=1.485 NRD=9.276 NRS=0 M=1 R=5.6 SA=75001 SB=75001.7
+ A=0.126 P=1.98 MULT=1
MM1003 A_347_47# N_A2_M1003_g A_269_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.1008 PD=1.23 PS=1.08 NRD=19.992 NRS=9.276 M=1 R=5.6 SA=75001.4 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1007 N_A_80_21#_M1007_d N_A1_M1007_g A_347_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=5.712 NRS=19.992 M=1 R=5.6 SA=75001.9
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_B1_M1008_g N_A_80_21#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_A_80_21#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.38115 AS=0.3339 PD=1.865 PS=3.05 NRD=12.4898 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1005 N_A_269_367#_M1005_d N_A3_M1005_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.21105 AS=0.38115 PD=1.595 PS=1.865 NRD=8.5892 NRS=38.2968 M=1
+ R=8.4 SA=75000.9 SB=75001.7 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A2_M1009_g N_A_269_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.25515 AS=0.21105 PD=1.665 PS=1.595 NRD=9.3772 NRS=0 M=1 R=8.4
+ SA=75001.4 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1000 N_A_269_367#_M1000_d N_A1_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.25515 PD=1.54 PS=1.665 NRD=0 NRS=10.1455 M=1 R=8.4
+ SA=75002 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_A_80_21#_M1006_d N_B1_M1006_g N_A_269_367#_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_30 VNB 0 1.17581e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__a31o_1.pxi.spice"
*
.ends
*
*
