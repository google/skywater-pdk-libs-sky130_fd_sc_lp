* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__einvn_8 A TE_B VGND VNB VPB VPWR Z
X0 a_305_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_305_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND a_110_57# a_305_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_305_47# a_110_57# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_305_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 Z A a_305_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR TE_B a_305_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VPWR TE_B a_305_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Z A a_305_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR TE_B a_110_57# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_305_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_305_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VPWR TE_B a_305_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_305_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_305_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Z A a_305_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 Z A a_305_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_305_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_305_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_305_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VPWR TE_B a_305_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_305_47# a_110_57# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 VGND a_110_57# a_305_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_305_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_305_47# a_110_57# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 Z A a_305_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 Z A a_305_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_305_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VGND a_110_57# a_305_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 Z A a_305_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_305_47# a_110_57# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 VGND TE_B a_110_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 VGND a_110_57# a_305_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 Z A a_305_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
