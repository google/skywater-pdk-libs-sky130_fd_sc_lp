* File: sky130_fd_sc_lp__dfrbp_lp.spice
* Created: Fri Aug 28 10:21:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfrbp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dfrbp_lp  VNB VPB D RESET_B CLK VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* D	D
* VPB	VPB
* VNB	VNB
MM1033 A_349_116# N_RESET_B_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.2184 PD=0.66 PS=1.88 NRD=18.564 NRS=67.14 M=1 R=2.8 SA=75000.4
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1023 N_A_111_457#_M1023_d N_D_M1023_g A_349_116# VNB NSHORT L=0.15 W=0.42
+ AD=0.13965 AS=0.0504 PD=1.085 PS=0.66 NRD=109.992 NRS=18.564 M=1 R=2.8
+ SA=75000.8 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1016 N_A_590_116#_M1016_d N_A_560_90#_M1016_g N_A_111_457#_M1023_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0756 AS=0.13965 PD=0.78 PS=1.085 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1045 A_692_116# N_A_662_90#_M1045_g N_A_590_116#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.13125 AS=0.0756 PD=1.045 PS=0.78 NRD=73.56 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1003 A_847_116# N_A_817_90#_M1003_g A_692_116# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.13125 PD=0.66 PS=1.045 NRD=18.564 NRS=73.56 M=1 R=2.8
+ SA=75002.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1040 N_VGND_M1040_d N_RESET_B_M1040_g A_847_116# VNB NSHORT L=0.15 W=0.42
+ AD=0.346 AS=0.0504 PD=2.48 PS=0.66 NRD=219.648 NRS=18.564 M=1 R=2.8 SA=75003.3
+ SB=75000.4 A=0.063 P=1.14 MULT=1
MM1004 A_1301_67# N_A_590_116#_M1004_g N_A_817_90#_M1004_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_A_590_116#_M1005_g A_1301_67# VNB NSHORT L=0.15 W=0.64
+ AD=0.165072 AS=0.0672 PD=1.33434 PS=0.85 NRD=13.116 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1006 A_1496_111# N_A_560_90#_M1006_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.108328 PD=0.63 PS=0.87566 NRD=14.28 NRS=33.564 M=1 R=2.8
+ SA=75001.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1041 N_A_662_90#_M1041_d N_A_560_90#_M1041_g A_1496_111# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 N_A_1799_379#_M1021_d N_A_662_90#_M1021_g N_A_817_90#_M1021_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.138023 AS=0.2336 PD=1.24981 PS=2.01 NRD=0 NRS=14.988 M=1
+ R=4.26667 SA=75000.3 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1036 A_2000_51# N_A_560_90#_M1036_g N_A_1799_379#_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1071 AS=0.0905774 PD=0.93 PS=0.820189 NRD=57.132 NRS=32.856 M=1
+ R=2.8 SA=75000.8 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_A_2102_25#_M1032_g A_2000_51# VNB NSHORT L=0.15 W=0.42
+ AD=0.34755 AS=0.1071 PD=2.075 PS=0.93 NRD=0 NRS=57.132 M=1 R=2.8 SA=75001.5
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1029 A_2493_51# N_RESET_B_M1029_g N_VGND_M1032_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.34755 PD=0.66 PS=2.075 NRD=18.564 NRS=392.856 M=1 R=2.8
+ SA=75003.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1030 N_A_2102_25#_M1030_d N_A_1799_379#_M1030_g A_2493_51# VNB NSHORT L=0.15
+ W=0.42 AD=0.2173 AS=0.0504 PD=1.98 PS=0.66 NRD=34.284 NRS=18.564 M=1 R=2.8
+ SA=75003.7 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1026 A_2825_48# N_CLK_M1026_g N_A_560_90#_M1026_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_CLK_M1027_g A_2825_48# VNB NSHORT L=0.15 W=0.42
+ AD=0.1071 AS=0.0504 PD=0.903333 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1050 A_3036_48# N_A_1799_379#_M1050_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2142 PD=1.05 PS=1.80667 NRD=7.14 NRS=33.564 M=1 R=5.6
+ SA=75000.7 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1035 N_Q_N_M1035_d N_A_1799_379#_M1035_g A_3036_48# VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1042 A_3309_137# N_A_1799_379#_M1042_g N_A_3222_137#_M1042_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1048 N_VGND_M1048_d N_A_1799_379#_M1048_g A_3309_137# VNB NSHORT L=0.15 W=0.42
+ AD=0.0952 AS=0.0441 PD=0.823333 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1015 A_3490_53# N_A_3222_137#_M1015_g N_VGND_M1048_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1904 PD=1.05 PS=1.64667 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1018 N_Q_M1018_d N_A_3222_137#_M1018_g A_3490_53# VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1043 N_A_111_457#_M1043_d N_D_M1043_g N_A_27_457#_M1043_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1134 PD=0.7 PS=1.38 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1014 A_197_457# N_RESET_B_M1014_g N_A_111_457#_M1043_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1022_d N_RESET_B_M1022_g A_197_457# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0938 AS=0.0441 PD=0.99 PS=0.63 NRD=51.5943 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.5 A=0.063 P=1.14 MULT=1
MM1012 N_A_27_457#_M1012_d N_D_M1012_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1134 AS=0.0938 PD=1.38 PS=0.99 NRD=0 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_A_590_116#_M1024_d N_A_560_90#_M1024_g N_A_484_411#_M1024_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.269575 PD=0.7 PS=2.21 NRD=0 NRS=128.976 M=1 R=2.8
+ SA=75000.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_111_457#_M1010_d N_A_662_90#_M1010_g N_A_590_116#_M1024_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1155 AS=0.0588 PD=1.39 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_817_90#_M1002_g N_A_484_411#_M1002_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.123975 AS=0.23115 PD=1.105 PS=2.13 NRD=112.645 NRS=232.342
+ M=1 R=2.8 SA=75000.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 A_1037_457# N_RESET_B_M1009_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.123975 PD=0.63 PS=1.105 NRD=23.443 NRS=112.645 M=1 R=2.8
+ SA=75000.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1038 N_A_590_116#_M1038_d N_RESET_B_M1038_g A_1037_457# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1134 AS=0.0441 PD=1.38 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75001.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_1301_373# N_A_590_116#_M1000_g N_A_817_90#_M1000_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.0882 AS=0.2268 PD=1.05 PS=2.22 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_A_590_116#_M1007_g A_1301_373# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.171065 AS=0.0882 PD=1.39054 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75001 A=0.126 P=1.98 MULT=1
MM1039 A_1480_413# N_A_560_90#_M1039_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.130335 PD=0.85 PS=1.05946 NRD=15.3857 NRS=32.308 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1047 N_A_662_90#_M1047_d N_A_560_90#_M1047_g A_1480_413# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.3924 AS=0.0672 PD=3.08 PS=0.85 NRD=171.784 NRS=15.3857 M=1
+ R=4.26667 SA=75001.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1019 N_A_1799_379#_M1019_d N_A_662_90#_M1019_g N_A_1712_379#_M1019_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0924 AS=0.1197 PD=0.816667 PS=1.41 NRD=77.3816
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1044 N_A_817_90#_M1044_d N_A_560_90#_M1044_g N_A_1799_379#_M1019_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2394 AS=0.1848 PD=2.25 PS=1.63333 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_A_2102_25#_M1013_g N_A_1712_379#_M1013_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_2102_25#_M1008_d N_A_1799_379#_M1008_g N_A_2185_397#_M1008_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1071 AS=0.2184 PD=0.93 PS=1.88 NRD=53.9386
+ NRS=110.222 M=1 R=2.8 SA=75000.4 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1017 A_2451_397# N_RESET_B_M1017_g N_A_2102_25#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1071 PD=0.63 PS=0.93 NRD=23.443 NRS=53.9386 M=1 R=2.8
+ SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_RESET_B_M1001_g A_2451_397# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.14625 AS=0.0441 PD=1.41 PS=0.63 NRD=137.526 NRS=23.443 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_A_2185_397#_M1020_d N_A_1799_379#_M1020_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1134 AS=0.14625 PD=1.38 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1049 A_2831_367# N_CLK_M1049_g N_A_560_90#_M1049_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.176 PD=0.85 PS=1.83 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1034 N_VPWR_M1034_d N_CLK_M1034_g A_2831_367# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.172632 AS=0.0672 PD=1.19579 PS=0.85 NRD=70.7821 NRS=15.3857 M=1 R=4.26667
+ SA=75000.6 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1031 A_3036_367# N_A_1799_379#_M1031_g N_VPWR_M1034_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.339868 PD=1.47 PS=2.35421 NRD=7.8012 NRS=1.5563 M=1
+ R=8.4 SA=75000.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1011 N_Q_N_M1011_d N_A_1799_379#_M1011_g A_3036_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1323 PD=3.09 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1028 A_3309_367# N_A_1799_379#_M1028_g N_A_3222_137#_M1028_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=15.3857 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1025 N_VPWR_M1025_d N_A_1799_379#_M1025_g A_3309_367# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.144674 AS=0.0672 PD=1.11495 PS=0.85 NRD=36.1495 NRS=15.3857 M=1
+ R=4.26667 SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1037 A_3490_367# N_A_3222_137#_M1037_g N_VPWR_M1025_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.284826 PD=1.47 PS=2.19505 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1046 N_Q_M1046_d N_A_3222_137#_M1046_g A_3490_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1323 PD=3.09 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX51_noxref VNB VPB NWDIODE A=35.0021 P=41.53
c_172 VNB 0 1.59406e-19 $X=0 $Y=0
c_327 VPB 0 2.15981e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dfrbp_lp.pxi.spice"
*
.ends
*
*
