* NGSPICE file created from sky130_fd_sc_lp__sdfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 a_1665_381# a_1517_63# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=2.4097e+12p ps=1.846e+07u
M1001 VPWR SCD a_414_487# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.048e+11p ps=1.92e+06u
M1002 VPWR a_1178_399# a_1136_451# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1003 Q a_1665_381# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=1.6005e+12p ps=1.41e+07u
M1004 a_328_119# D a_256_119# VNB nshort w=420000u l=150000u
+  ad=3.423e+11p pd=3.31e+06u as=8.82e+10p ps=1.26e+06u
M1005 a_414_487# a_55_119# a_328_119# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.905e+11p ps=3.21e+06u
M1006 a_831_47# a_610_487# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1007 a_256_119# a_55_119# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND SCE a_55_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1009 VGND SCD a_464_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 VGND a_1665_381# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1136_451# a_610_487# a_1047_125# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1012 a_1047_125# a_610_487# a_328_119# VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1013 Q a_1665_381# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1014 a_1178_399# a_1047_125# VPWR VPB phighvt w=840000u l=150000u
+  ad=4.62e+11p pd=2.78e+06u as=0p ps=0u
M1015 a_1178_399# a_1047_125# VGND VNB nshort w=640000u l=150000u
+  ad=2.158e+11p pd=2.03e+06u as=0p ps=0u
M1016 a_1623_493# a_831_47# a_1517_63# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.688e+11p ps=2.43e+06u
M1017 a_464_119# SCE a_328_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_328_119# D a_256_487# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1019 a_1517_63# a_610_487# a_1178_399# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1178_399# a_1149_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1021 a_1047_125# a_831_47# a_328_119# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_1665_381# a_1623_493# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_610_487# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1024 VPWR a_1665_381# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1665_381# a_1517_63# VGND VNB nshort w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1026 a_1670_63# a_610_487# a_1517_63# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.583e+11p ps=2.07e+06u
M1027 a_1149_125# a_831_47# a_1047_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_1665_381# a_1670_63# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR SCE a_55_119# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1030 a_256_487# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_610_487# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1032 a_831_47# a_610_487# VGND VNB nshort w=420000u l=150000u
+  ad=1.428e+11p pd=1.52e+06u as=0p ps=0u
M1033 a_1517_63# a_831_47# a_1178_399# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

