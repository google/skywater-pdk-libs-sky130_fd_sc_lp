* File: sky130_fd_sc_lp__and4bb_m.pex.spice
* Created: Fri Aug 28 10:09:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4BB_M%A_N 3 6 9 10 11 12 13 17
r34 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.56
+ $Y=0.97 $X2=0.56 $Y2=0.97
r35 13 18 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=0.97
r36 12 18 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.64 $Y=0.925
+ $X2=0.64 $Y2=0.97
r37 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.56 $Y=1.31
+ $X2=0.56 $Y2=0.97
r38 10 11 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=1.31
+ $X2=0.56 $Y2=1.475
r39 9 17 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=0.805
+ $X2=0.56 $Y2=0.97
r40 6 11 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.61 $Y=2.195
+ $X2=0.61 $Y2=1.475
r41 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.61 $Y=0.485 $X2=0.61
+ $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_M%B_N 3 6 9 10 11 12 13 17
r40 12 13 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.165 $Y=0.925
+ $X2=1.165 $Y2=1.295
r41 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.13
+ $Y=0.97 $X2=1.13 $Y2=0.97
r42 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.13 $Y=1.31
+ $X2=1.13 $Y2=0.97
r43 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.31
+ $X2=1.13 $Y2=1.475
r44 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=0.805
+ $X2=1.13 $Y2=0.97
r45 6 11 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.04 $Y=2.195
+ $X2=1.04 $Y2=1.475
r46 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.04 $Y=0.485 $X2=1.04
+ $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_M%A_54_55# 1 2 11 12 14 18 21 22 23 25 28 30
+ 34 35 40 42
c74 35 0 1.4009e-19 $X=1.7 $Y=1.32
r75 37 40 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.21 $Y=0.46
+ $X2=0.395 $Y2=0.46
r76 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.7 $Y=1.32
+ $X2=1.7 $Y2=1.32
r77 32 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.7 $Y=1.655
+ $X2=1.7 $Y2=1.32
r78 31 42 3.08518 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.5 $Y=1.74
+ $X2=0.312 $Y2=1.74
r79 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.615 $Y=1.74
+ $X2=1.7 $Y2=1.655
r80 30 31 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=1.615 $Y=1.74
+ $X2=0.5 $Y2=1.74
r81 26 42 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=0.312 $Y=1.825
+ $X2=0.312 $Y2=1.74
r82 26 28 9.3732 $w=3.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.312 $Y=1.825
+ $X2=0.312 $Y2=2.13
r83 25 42 3.43356 $w=2.72e-07 $l=1.38109e-07 $layer=LI1_cond $X=0.21 $Y=1.655
+ $X2=0.312 $Y2=1.74
r84 24 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.21 $Y=0.625
+ $X2=0.21 $Y2=0.46
r85 24 25 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.21 $Y=0.625
+ $X2=0.21 $Y2=1.655
r86 22 23 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.825 $Y=2.415
+ $X2=1.825 $Y2=2.565
r87 21 22 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.79 $Y=1.825
+ $X2=1.79 $Y2=2.415
r88 20 35 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.7 $Y=1.66 $X2=1.7
+ $Y2=1.32
r89 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.66 $X2=1.7
+ $Y2=1.825
r90 16 35 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.7 $Y=1.305 $X2=1.7
+ $Y2=1.32
r91 16 18 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.7 $Y=1.23 $X2=2
+ $Y2=1.23
r92 12 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2 $Y=1.155 $X2=2
+ $Y2=1.23
r93 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2 $Y=1.155 $X2=2
+ $Y2=0.835
r94 11 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.86 $Y=2.885
+ $X2=1.86 $Y2=2.565
r95 2 28 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.27
+ $Y=1.985 $X2=0.395 $Y2=2.13
r96 1 40 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.275 $X2=0.395 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_M%A_223_55# 1 2 9 14 17 18 21 22 24 28 29 31
+ 36
r73 36 39 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.255 $Y=2.09
+ $X2=1.255 $Y2=2.17
r74 31 34 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.255 $Y=0.35
+ $X2=1.255 $Y2=0.43
r75 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.27 $Y=1.7
+ $X2=2.27 $Y2=1.7
r76 26 28 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.27 $Y=2.005
+ $X2=2.27 $Y2=1.7
r77 25 36 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.36 $Y=2.09
+ $X2=1.255 $Y2=2.09
r78 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.105 $Y=2.09
+ $X2=2.27 $Y2=2.005
r79 24 25 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.105 $Y=2.09
+ $X2=1.36 $Y2=2.09
r80 22 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=0.35
+ $X2=2.45 $Y2=0.515
r81 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.45
+ $Y=0.35 $X2=2.45 $Y2=0.35
r82 19 31 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.36 $Y=0.35
+ $X2=1.255 $Y2=0.35
r83 19 21 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=1.36 $Y=0.35
+ $X2=2.45 $Y2=0.35
r84 17 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.27 $Y=2.04
+ $X2=2.27 $Y2=1.7
r85 17 18 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=2.04
+ $X2=2.27 $Y2=2.205
r86 16 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.535
+ $X2=2.27 $Y2=1.7
r87 14 16 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=2.36 $Y=0.835 $X2=2.36
+ $Y2=1.535
r88 14 44 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.36 $Y=0.835
+ $X2=2.36 $Y2=0.515
r89 9 18 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.29 $Y=2.885
+ $X2=2.29 $Y2=2.205
r90 2 39 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.985 $X2=1.255 $Y2=2.17
r91 1 34 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.275 $X2=1.255 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_M%C 3 7 8 9 13 14 15
r47 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.32
+ $X2=2.81 $Y2=1.485
r48 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.32
+ $X2=2.81 $Y2=1.155
r49 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=1.32 $X2=2.81 $Y2=1.32
r50 9 14 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=2.64 $Y=1.307 $X2=2.81
+ $Y2=1.307
r51 8 9 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.307 $X2=2.64
+ $Y2=1.307
r52 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.9 $Y=0.835 $X2=2.9
+ $Y2=1.155
r53 3 16 717.872 $w=1.5e-07 $l=1.4e-06 $layer=POLY_cond $X=2.72 $Y=2.885
+ $X2=2.72 $Y2=1.485
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_M%D 3 7 9 12
r44 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=2.035
+ $X2=3.17 $Y2=2.2
r45 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=2.035
+ $X2=3.17 $Y2=1.87
r46 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=2.035 $X2=3.17 $Y2=2.035
r47 7 14 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=3.26 $Y=0.835
+ $X2=3.26 $Y2=1.87
r48 3 15 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=3.15 $Y=2.885
+ $X2=3.15 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_M%A_332_125# 1 2 3 11 14 18 20 21 27 29 30 32
+ 33 34 35 37 40 41 48 50 51
c117 48 0 1.8805e-19 $X=3.24 $Y=1.67
c118 34 0 1.8253e-19 $X=2.825 $Y=1.67
r119 51 53 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.732 $Y=1.75
+ $X2=3.732 $Y2=1.585
r120 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.71
+ $Y=1.75 $X2=3.71 $Y2=1.75
r121 42 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=1.67
+ $X2=3.24 $Y2=1.67
r122 41 50 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=1.67
+ $X2=3.71 $Y2=1.67
r123 41 42 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.625 $Y=1.67
+ $X2=3.325 $Y2=1.67
r124 40 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=1.585
+ $X2=3.24 $Y2=1.67
r125 39 40 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.24 $Y=0.975
+ $X2=3.24 $Y2=1.585
r126 35 45 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.935 $Y=2.52
+ $X2=2.74 $Y2=2.52
r127 35 37 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.935 $Y=2.605
+ $X2=2.935 $Y2=2.82
r128 33 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=1.67
+ $X2=3.24 $Y2=1.67
r129 33 34 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.155 $Y=1.67
+ $X2=2.825 $Y2=1.67
r130 32 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=2.435
+ $X2=2.74 $Y2=2.52
r131 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.74 $Y=1.755
+ $X2=2.825 $Y2=1.67
r132 31 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.74 $Y=1.755
+ $X2=2.74 $Y2=2.435
r133 29 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.655 $Y=2.52
+ $X2=2.74 $Y2=2.52
r134 29 30 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.655 $Y=2.52
+ $X2=2.18 $Y2=2.52
r135 25 30 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.075 $Y=2.605
+ $X2=2.18 $Y2=2.52
r136 25 27 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.075 $Y=2.605
+ $X2=2.075 $Y2=2.82
r137 21 39 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.155 $Y=0.81
+ $X2=3.24 $Y2=0.975
r138 21 23 47.8438 $w=3.28e-07 $l=1.37e-06 $layer=LI1_cond $X=3.155 $Y=0.81
+ $X2=1.785 $Y2=0.81
r139 18 53 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=3.845 $Y=0.835
+ $X2=3.845 $Y2=1.585
r140 14 20 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.62 $Y=2.885
+ $X2=3.62 $Y2=2.255
r141 11 20 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=3.732 $Y=2.068
+ $X2=3.732 $Y2=2.255
r142 10 51 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=3.732 $Y=1.772
+ $X2=3.732 $Y2=1.75
r143 10 11 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=3.732 $Y=1.772
+ $X2=3.732 $Y2=2.068
r144 3 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=2.675 $X2=2.935 $Y2=2.82
r145 2 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=2.675 $X2=2.075 $Y2=2.82
r146 1 23 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.625 $X2=1.785 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_M%VPWR 1 2 3 4 17 21 25 29 32 33 35 36 38 39
+ 40 53 54 57
r50 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 42 57 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.93 $Y=3.33
+ $X2=0.825 $Y2=3.33
r57 42 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.93 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 40 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 40 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 40 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 38 50 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.22 $Y=3.33 $X2=3.12
+ $Y2=3.33
r62 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=3.33
+ $X2=3.385 $Y2=3.33
r63 37 53 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.55 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=3.33
+ $X2=3.385 $Y2=3.33
r65 35 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=3.33 $X2=2.16
+ $Y2=3.33
r66 35 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.505 $Y2=3.33
r67 34 50 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 34 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=2.505 $Y2=3.33
r69 32 44 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.54 $Y=3.33 $X2=1.2
+ $Y2=3.33
r70 32 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.645 $Y2=3.33
r71 31 47 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.75 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 31 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.75 $Y=3.33
+ $X2=1.645 $Y2=3.33
r73 27 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=3.245
+ $X2=3.385 $Y2=3.33
r74 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.385 $Y=3.245
+ $X2=3.385 $Y2=2.95
r75 23 36 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=3.245
+ $X2=2.505 $Y2=3.33
r76 23 25 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.505 $Y=3.245
+ $X2=2.505 $Y2=2.95
r77 19 33 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=3.245
+ $X2=1.645 $Y2=3.33
r78 19 21 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.645 $Y=3.245
+ $X2=1.645 $Y2=2.95
r79 15 57 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=3.33
r80 15 17 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=2.26
r81 4 29 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=2.675 $X2=3.385 $Y2=2.95
r82 3 25 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=2.675 $X2=2.505 $Y2=2.95
r83 2 21 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=2.675 $X2=1.645 $Y2=2.95
r84 1 17 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=1.985 $X2=0.825 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_M%X 1 2 10 13 14 15 16
r16 15 16 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=4.07 $Y=1.295
+ $X2=4.07 $Y2=1.665
r17 14 15 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=4.07 $Y=0.925
+ $X2=4.07 $Y2=1.295
r18 14 25 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=4.07 $Y=0.925
+ $X2=4.07 $Y2=0.77
r19 13 25 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=4.07 $Y=0.555
+ $X2=4.07 $Y2=0.77
r20 11 16 57.7895 $w=1.88e-07 $l=9.9e-07 $layer=LI1_cond $X=4.07 $Y=2.655
+ $X2=4.07 $Y2=1.665
r21 10 11 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=2.82
+ $X2=4.07 $Y2=2.655
r22 8 10 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=3.835 $Y=2.82
+ $X2=4.07 $Y2=2.82
r23 2 8 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.695
+ $Y=2.675 $X2=3.835 $Y2=2.82
r24 1 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.625 $X2=4.06 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_M%VGND 1 2 11 15 17 19 29 30 33 36
r42 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r43 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r45 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r46 27 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.61
+ $Y2=0
r47 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=4.08
+ $Y2=0
r48 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r49 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r52 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 20 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=0.825
+ $Y2=0
r54 20 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=1.2
+ $Y2=0
r55 19 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.61
+ $Y2=0
r56 19 25 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.12
+ $Y2=0
r57 17 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r58 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r59 13 36 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=0.085
+ $X2=3.61 $Y2=0
r60 13 15 36.1775 $w=2.08e-07 $l=6.85e-07 $layer=LI1_cond $X=3.61 $Y=0.085
+ $X2=3.61 $Y2=0.77
r61 9 33 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r62 9 11 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.42
r63 2 15 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.625 $X2=3.61 $Y2=0.77
r64 1 11 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.685
+ $Y=0.275 $X2=0.825 $Y2=0.42
.ends

