* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2i_0 A0 A1 S VGND VNB VPB VPWR Y
X0 a_465_491# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_47_48# S VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_47_48# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 Y A1 a_436_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_47_48# a_244_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_436_48# S VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_244_48# A0 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_47_48# a_292_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_292_491# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 Y A0 a_465_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
