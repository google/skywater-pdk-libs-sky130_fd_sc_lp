* File: sky130_fd_sc_lp__xor2_m.spice
* Created: Fri Aug 28 11:36:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xor2_m.pex.spice"
.subckt sky130_fd_sc_lp__xor2_m  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_A_41_535#_M1000_d N_B_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_41_535#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.12285 AS=0.0588 PD=1.005 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1007 A_357_156# N_A_M1007_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.12285 PD=0.63 PS=1.005 NRD=14.28 NRS=81.42 M=1 R=2.8 SA=75001.4
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_B_M1006_g A_357_156# VNB NSHORT L=0.15 W=0.42 AD=0.10605
+ AS=0.0441 PD=0.925 PS=0.63 NRD=64.284 NRS=14.28 M=1 R=2.8 SA=75001.7
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_41_535#_M1003_g N_X_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1512 AS=0.10605 PD=1.56 PS=0.925 NRD=27.132 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1004 A_124_535# N_B_M1004_g N_A_41_535#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_124_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_282_535#_M1008_d N_A_M1008_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_A_282_535#_M1008_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_41_535#_M1001_g N_A_282_535#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_29 VNB 0 1.46329e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__xor2_m.pxi.spice"
*
.ends
*
*
