* File: sky130_fd_sc_lp__nand4bb_4.pxi.spice
* Created: Fri Aug 28 10:52:36 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4BB_4%A_N N_A_N_M1032_g N_A_N_M1002_g A_N A_N
+ N_A_N_c_152_n N_A_N_c_153_n PM_SKY130_FD_SC_LP__NAND4BB_4%A_N
x_PM_SKY130_FD_SC_LP__NAND4BB_4%B_N N_B_N_c_180_n N_B_N_M1004_g N_B_N_M1011_g
+ B_N B_N N_B_N_c_183_n PM_SKY130_FD_SC_LP__NAND4BB_4%B_N
x_PM_SKY130_FD_SC_LP__NAND4BB_4%A_44_69# N_A_44_69#_M1032_s N_A_44_69#_M1002_s
+ N_A_44_69#_M1015_g N_A_44_69#_M1007_g N_A_44_69#_M1016_g N_A_44_69#_M1014_g
+ N_A_44_69#_M1025_g N_A_44_69#_M1028_g N_A_44_69#_M1035_g N_A_44_69#_M1029_g
+ N_A_44_69#_c_217_n N_A_44_69#_c_227_n N_A_44_69#_c_228_n N_A_44_69#_c_218_n
+ N_A_44_69#_c_219_n N_A_44_69#_c_263_p N_A_44_69#_c_220_n N_A_44_69#_c_230_n
+ N_A_44_69#_c_221_n N_A_44_69#_c_232_n N_A_44_69#_c_222_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%A_44_69#
x_PM_SKY130_FD_SC_LP__NAND4BB_4%A_217_69# N_A_217_69#_M1004_d
+ N_A_217_69#_M1011_d N_A_217_69#_M1005_g N_A_217_69#_M1000_g
+ N_A_217_69#_M1018_g N_A_217_69#_M1012_g N_A_217_69#_M1023_g
+ N_A_217_69#_M1022_g N_A_217_69#_M1031_g N_A_217_69#_M1030_g
+ N_A_217_69#_c_345_n N_A_217_69#_c_334_n N_A_217_69#_c_335_n
+ N_A_217_69#_c_370_n N_A_217_69#_c_336_n N_A_217_69#_c_337_n
+ N_A_217_69#_c_338_n N_A_217_69#_c_339_n N_A_217_69#_c_340_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%A_217_69#
x_PM_SKY130_FD_SC_LP__NAND4BB_4%C N_C_M1006_g N_C_c_473_n N_C_M1001_g
+ N_C_M1009_g N_C_c_475_n N_C_M1013_g N_C_M1020_g N_C_c_477_n N_C_M1017_g
+ N_C_M1033_g N_C_c_479_n N_C_M1019_g C C C C N_C_c_481_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%C
x_PM_SKY130_FD_SC_LP__NAND4BB_4%D N_D_M1003_g N_D_c_552_n N_D_M1008_g
+ N_D_M1021_g N_D_c_554_n N_D_M1010_g N_D_M1026_g N_D_c_556_n N_D_M1024_g
+ N_D_M1027_g N_D_c_558_n N_D_M1034_g D D D D N_D_c_560_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%D
x_PM_SKY130_FD_SC_LP__NAND4BB_4%VPWR N_VPWR_M1002_d N_VPWR_M1007_d
+ N_VPWR_M1014_d N_VPWR_M1035_d N_VPWR_M1018_s N_VPWR_M1031_s N_VPWR_M1009_d
+ N_VPWR_M1033_d N_VPWR_M1021_s N_VPWR_M1027_s N_VPWR_c_622_n N_VPWR_c_623_n
+ N_VPWR_c_624_n N_VPWR_c_625_n N_VPWR_c_626_n N_VPWR_c_627_n N_VPWR_c_628_n
+ N_VPWR_c_629_n N_VPWR_c_630_n N_VPWR_c_631_n N_VPWR_c_632_n N_VPWR_c_633_n
+ N_VPWR_c_634_n N_VPWR_c_635_n N_VPWR_c_636_n N_VPWR_c_637_n N_VPWR_c_638_n
+ N_VPWR_c_639_n VPWR N_VPWR_c_640_n N_VPWR_c_641_n N_VPWR_c_642_n
+ N_VPWR_c_643_n N_VPWR_c_644_n N_VPWR_c_645_n N_VPWR_c_646_n N_VPWR_c_647_n
+ N_VPWR_c_648_n N_VPWR_c_649_n N_VPWR_c_650_n N_VPWR_c_621_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%VPWR
x_PM_SKY130_FD_SC_LP__NAND4BB_4%Y N_Y_M1015_d N_Y_M1028_d N_Y_M1007_s
+ N_Y_M1025_s N_Y_M1005_d N_Y_M1023_d N_Y_M1006_s N_Y_M1020_s N_Y_M1003_d
+ N_Y_M1026_d N_Y_c_772_n N_Y_c_865_n N_Y_c_774_n N_Y_c_775_n N_Y_c_869_n
+ N_Y_c_773_n N_Y_c_777_n N_Y_c_778_n N_Y_c_874_n N_Y_c_876_n N_Y_c_779_n
+ N_Y_c_780_n N_Y_c_882_n N_Y_c_781_n N_Y_c_886_n N_Y_c_782_n N_Y_c_891_n
+ N_Y_c_783_n N_Y_c_784_n Y Y Y Y Y N_Y_c_787_n N_Y_c_788_n N_Y_c_835_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%Y
x_PM_SKY130_FD_SC_LP__NAND4BB_4%VGND N_VGND_M1032_d N_VGND_M1008_s
+ N_VGND_M1024_s N_VGND_c_905_n N_VGND_c_906_n N_VGND_c_907_n VGND
+ N_VGND_c_908_n N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n N_VGND_c_912_n
+ N_VGND_c_913_n N_VGND_c_914_n N_VGND_c_915_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%VGND
x_PM_SKY130_FD_SC_LP__NAND4BB_4%A_324_45# N_A_324_45#_M1015_s
+ N_A_324_45#_M1016_s N_A_324_45#_M1029_s N_A_324_45#_M1012_d
+ N_A_324_45#_M1030_d N_A_324_45#_c_1006_n N_A_324_45#_c_1025_n
+ N_A_324_45#_c_1007_n N_A_324_45#_c_1031_n N_A_324_45#_c_1008_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%A_324_45#
x_PM_SKY130_FD_SC_LP__NAND4BB_4%A_842_67# N_A_842_67#_M1000_s
+ N_A_842_67#_M1022_s N_A_842_67#_M1001_d N_A_842_67#_M1017_d
+ N_A_842_67#_c_1063_n N_A_842_67#_c_1064_n N_A_842_67#_c_1065_n
+ N_A_842_67#_c_1066_n N_A_842_67#_c_1067_n N_A_842_67#_c_1068_n
+ N_A_842_67#_c_1069_n N_A_842_67#_c_1091_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%A_842_67#
x_PM_SKY130_FD_SC_LP__NAND4BB_4%A_1251_47# N_A_1251_47#_M1001_s
+ N_A_1251_47#_M1013_s N_A_1251_47#_M1019_s N_A_1251_47#_M1010_d
+ N_A_1251_47#_M1034_d N_A_1251_47#_c_1125_n N_A_1251_47#_c_1129_n
+ N_A_1251_47#_c_1150_n N_A_1251_47#_c_1133_n N_A_1251_47#_c_1155_n
+ N_A_1251_47#_c_1137_n N_A_1251_47#_c_1160_n N_A_1251_47#_c_1132_n
+ N_A_1251_47#_c_1143_n N_A_1251_47#_c_1141_n
+ PM_SKY130_FD_SC_LP__NAND4BB_4%A_1251_47#
cc_1 VNB N_A_N_M1002_g 0.00167964f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_2 VNB A_N 0.00759102f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_N_c_152_n 0.0329407f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.46
cc_4 VNB N_A_N_c_153_n 0.0202539f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.295
cc_5 VNB N_B_N_c_180_n 0.0195161f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.295
cc_6 VNB N_B_N_M1011_g 0.00183824f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_7 VNB B_N 0.00437549f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_B_N_c_183_n 0.0470857f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.295
cc_9 VNB N_A_44_69#_M1015_g 0.0229488f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_10 VNB N_A_44_69#_M1016_g 0.0206128f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.295
cc_11 VNB N_A_44_69#_M1028_g 0.0205804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_44_69#_M1029_g 0.0199448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_44_69#_c_217_n 0.0259117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_44_69#_c_218_n 4.10739e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_44_69#_c_219_n 0.00389221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_44_69#_c_220_n 0.00800596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_44_69#_c_221_n 0.028412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_44_69#_c_222_n 0.0777913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_217_69#_M1000_g 0.0204831f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.46
cc_20 VNB N_A_217_69#_M1012_g 0.0181449f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.665
cc_21 VNB N_A_217_69#_M1022_g 0.0181498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_217_69#_M1030_g 0.024183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_217_69#_c_334_n 0.00206211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_217_69#_c_335_n 0.0151082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_217_69#_c_336_n 0.00750547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_217_69#_c_337_n 0.00347969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_217_69#_c_338_n 0.0023475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_217_69#_c_339_n 0.0298596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_217_69#_c_340_n 0.0737665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_M1006_g 0.00864269f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.765
cc_31 VNB N_C_c_473_n 0.019851f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_32 VNB N_C_M1009_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_C_c_475_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.46
cc_34 VNB N_C_M1020_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.295
cc_35 VNB N_C_c_477_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_C_M1033_g 0.00730538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_C_c_479_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB C 0.00895776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_C_c_481_n 0.0975121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_D_M1003_g 0.00730538f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.765
cc_41 VNB N_D_c_552_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_42 VNB N_D_M1021_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_D_c_554_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.46
cc_44 VNB N_D_M1026_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.295
cc_45 VNB N_D_c_556_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_D_M1027_g 0.0111859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_D_c_558_n 0.0218823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB D 0.0153863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_D_c_560_n 0.100731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VPWR_c_621_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_Y_c_772_n 0.00857568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_Y_c_773_n 0.00294896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_905_n 0.00332106f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.46
cc_54 VNB N_VGND_c_906_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.625
cc_55 VNB N_VGND_c_907_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.46
cc_56 VNB N_VGND_c_908_n 0.0188084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_909_n 0.173699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_910_n 0.0130339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_911_n 0.0159403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_912_n 0.505079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_913_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_914_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_915_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_324_45#_c_1006_n 0.0112634f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.625
cc_65 VNB N_A_324_45#_c_1007_n 0.00658237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_324_45#_c_1008_n 0.00203565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_842_67#_c_1063_n 0.0184784f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.295
cc_68 VNB N_A_842_67#_c_1064_n 0.0103733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_842_67#_c_1065_n 0.00782452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_842_67#_c_1066_n 0.00416423f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.46
cc_71 VNB N_A_842_67#_c_1067_n 0.00219381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_842_67#_c_1068_n 0.00319629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_842_67#_c_1069_n 0.0014302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VPB N_A_N_M1002_g 0.0235728f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.465
cc_75 VPB A_N 0.00571117f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_76 VPB N_B_N_M1011_g 0.0243795f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.465
cc_77 VPB B_N 0.00281621f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_78 VPB N_A_44_69#_M1007_g 0.0212049f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.46
cc_79 VPB N_A_44_69#_M1014_g 0.0180108f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.665
cc_80 VPB N_A_44_69#_M1025_g 0.0179863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_44_69#_M1035_g 0.0178455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_44_69#_c_227_n 0.00981458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A_44_69#_c_228_n 0.0208364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_44_69#_c_218_n 0.012511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A_44_69#_c_230_n 0.00790378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_44_69#_c_221_n 0.0130284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_44_69#_c_232_n 0.0279419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_44_69#_c_222_n 0.0195097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_217_69#_M1005_g 0.018914f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_90 VPB N_A_217_69#_M1018_g 0.0185025f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.295
cc_91 VPB N_A_217_69#_M1023_g 0.0185219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_217_69#_M1031_g 0.0246792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_217_69#_c_345_n 0.0128605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_217_69#_c_335_n 0.00631369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_217_69#_c_339_n 0.0100886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_217_69#_c_340_n 0.0143762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_C_M1006_g 0.0241614f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.765
cc_98 VPB N_C_M1009_g 0.0183287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_C_M1020_g 0.0183287f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.295
cc_100 VPB N_C_M1033_g 0.0184015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_D_M1003_g 0.0184015f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.765
cc_102 VPB N_D_M1021_g 0.0183287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_D_M1026_g 0.0183287f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.295
cc_104 VPB N_D_M1027_g 0.0272274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_622_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_623_n 0.0188957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_624_n 3.14366e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_625_n 0.0146078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_626_n 0.00375103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_627_n 3.20722e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_628_n 3.15883e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_629_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_630_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_631_n 3.14366e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_632_n 0.0119328f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_633_n 0.0572804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_634_n 0.027052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_635_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_636_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_637_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_638_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_639_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_640_n 0.0185059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_641_n 0.0154314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_642_n 0.0129339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_643_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_644_n 0.0146078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_645_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_646_n 0.00439477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_647_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_648_n 0.0285671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_649_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_650_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_621_n 0.0538593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_Y_c_774_n 0.00304705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_Y_c_775_n 0.00198153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_Y_c_773_n 0.00144235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_Y_c_777_n 0.00614929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_Y_c_778_n 0.00249758f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_Y_c_779_n 0.00308535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_Y_c_780_n 0.0170787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_Y_c_781_n 0.00484808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_Y_c_782_n 0.00677023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_Y_c_783_n 0.00145912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_Y_c_784_n 0.00145912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB Y 0.00186719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB Y 0.00144499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_Y_c_787_n 0.00308636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_Y_c_788_n 0.00463242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 A_N N_B_N_c_180_n 0.00413084f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_151 N_A_N_c_153_n N_B_N_c_180_n 0.0163566f $X=0.53 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_N_M1002_g N_B_N_M1011_g 0.0539128f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_153 A_N B_N 0.0426481f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A_N_c_152_n B_N 2.65922e-19 $X=0.53 $Y=1.46 $X2=0 $Y2=0
cc_155 N_A_N_c_152_n N_B_N_c_183_n 0.0174931f $X=0.53 $Y=1.46 $X2=0 $Y2=0
cc_156 N_A_N_c_153_n N_A_44_69#_c_217_n 4.52033e-19 $X=0.53 $Y=1.295 $X2=0 $Y2=0
cc_157 N_A_N_M1002_g N_A_44_69#_c_228_n 0.0116282f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_158 A_N N_A_44_69#_c_228_n 0.0111656f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_159 A_N N_A_44_69#_c_220_n 6.7912e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A_N_c_152_n N_A_44_69#_c_220_n 0.00333765f $X=0.53 $Y=1.46 $X2=0 $Y2=0
cc_161 N_A_N_c_152_n N_A_44_69#_c_230_n 0.00311636f $X=0.53 $Y=1.46 $X2=0 $Y2=0
cc_162 N_A_N_M1002_g N_A_44_69#_c_221_n 0.00498996f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_163 A_N N_A_44_69#_c_221_n 0.0425835f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A_N_c_152_n N_A_44_69#_c_221_n 0.00815572f $X=0.53 $Y=1.46 $X2=0 $Y2=0
cc_165 N_A_N_c_153_n N_A_44_69#_c_221_n 0.0044195f $X=0.53 $Y=1.295 $X2=0 $Y2=0
cc_166 N_A_N_M1002_g N_A_217_69#_c_345_n 7.68042e-19 $X=0.58 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_N_M1002_g N_VPWR_c_622_n 0.0150702f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A_N_M1002_g N_VPWR_c_640_n 0.00486043f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_N_M1002_g N_VPWR_c_621_n 0.0056736f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_170 A_N N_VGND_c_905_n 0.0182644f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A_N_c_153_n N_VGND_c_905_n 0.0151774f $X=0.53 $Y=1.295 $X2=0 $Y2=0
cc_172 N_A_N_c_153_n N_VGND_c_908_n 0.00400407f $X=0.53 $Y=1.295 $X2=0 $Y2=0
cc_173 N_A_N_c_153_n N_VGND_c_912_n 0.00797993f $X=0.53 $Y=1.295 $X2=0 $Y2=0
cc_174 N_B_N_c_183_n N_A_44_69#_M1015_g 5.39709e-19 $X=1.2 $Y=1.46 $X2=0 $Y2=0
cc_175 N_B_N_M1011_g N_A_44_69#_c_228_n 0.0171454f $X=1.01 $Y=2.465 $X2=0 $Y2=0
cc_176 B_N N_A_44_69#_c_228_n 6.39745e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_177 N_B_N_c_183_n N_A_44_69#_c_222_n 0.00347448f $X=1.2 $Y=1.46 $X2=0 $Y2=0
cc_178 N_B_N_M1011_g N_A_217_69#_c_345_n 0.00532463f $X=1.01 $Y=2.465 $X2=0
+ $Y2=0
cc_179 B_N N_A_217_69#_c_345_n 0.0163392f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_180 N_B_N_c_183_n N_A_217_69#_c_345_n 0.00372553f $X=1.2 $Y=1.46 $X2=0 $Y2=0
cc_181 N_B_N_c_180_n N_A_217_69#_c_334_n 4.43331e-19 $X=1.01 $Y=1.295 $X2=0
+ $Y2=0
cc_182 N_B_N_c_180_n N_A_217_69#_c_335_n 0.00486173f $X=1.01 $Y=1.295 $X2=0
+ $Y2=0
cc_183 N_B_N_M1011_g N_A_217_69#_c_335_n 0.00415075f $X=1.01 $Y=2.465 $X2=0
+ $Y2=0
cc_184 B_N N_A_217_69#_c_335_n 0.0343363f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_185 N_B_N_c_183_n N_A_217_69#_c_335_n 0.00392911f $X=1.2 $Y=1.46 $X2=0 $Y2=0
cc_186 B_N N_A_217_69#_c_336_n 0.0134181f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_187 N_B_N_c_183_n N_A_217_69#_c_336_n 0.00279125f $X=1.2 $Y=1.46 $X2=0 $Y2=0
cc_188 N_B_N_M1011_g N_VPWR_c_622_n 0.0235018f $X=1.01 $Y=2.465 $X2=0 $Y2=0
cc_189 N_B_N_M1011_g N_VPWR_c_634_n 0.00486043f $X=1.01 $Y=2.465 $X2=0 $Y2=0
cc_190 N_B_N_M1011_g N_VPWR_c_621_n 0.00597709f $X=1.01 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B_N_c_180_n N_VGND_c_905_n 0.0145378f $X=1.01 $Y=1.295 $X2=0 $Y2=0
cc_192 N_B_N_c_180_n N_VGND_c_909_n 0.00400407f $X=1.01 $Y=1.295 $X2=0 $Y2=0
cc_193 N_B_N_c_180_n N_VGND_c_912_n 0.00804497f $X=1.01 $Y=1.295 $X2=0 $Y2=0
cc_194 N_B_N_c_180_n N_A_324_45#_c_1006_n 0.00147458f $X=1.01 $Y=1.295 $X2=0
+ $Y2=0
cc_195 N_A_44_69#_c_228_n N_A_217_69#_M1011_d 0.00711717f $X=1.85 $Y=2.425 $X2=0
+ $Y2=0
cc_196 N_A_44_69#_M1035_g N_A_217_69#_M1005_g 0.0160692f $X=3.515 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_A_44_69#_M1029_g N_A_217_69#_M1000_g 0.026329f $X=3.545 $Y=0.755 $X2=0
+ $Y2=0
cc_198 N_A_44_69#_c_228_n N_A_217_69#_c_345_n 0.0439726f $X=1.85 $Y=2.425 $X2=0
+ $Y2=0
cc_199 N_A_44_69#_c_218_n N_A_217_69#_c_345_n 0.0209553f $X=1.935 $Y=2.34 $X2=0
+ $Y2=0
cc_200 N_A_44_69#_M1015_g N_A_217_69#_c_334_n 0.00385447f $X=2.095 $Y=0.755
+ $X2=0 $Y2=0
cc_201 N_A_44_69#_M1015_g N_A_217_69#_c_335_n 0.0128708f $X=2.095 $Y=0.755 $X2=0
+ $Y2=0
cc_202 N_A_44_69#_c_218_n N_A_217_69#_c_335_n 0.0237471f $X=1.935 $Y=2.34 $X2=0
+ $Y2=0
cc_203 N_A_44_69#_c_219_n N_A_217_69#_c_335_n 0.0186526f $X=2.02 $Y=1.495 $X2=0
+ $Y2=0
cc_204 N_A_44_69#_c_222_n N_A_217_69#_c_335_n 0.00183038f $X=3.515 $Y=1.51 $X2=0
+ $Y2=0
cc_205 N_A_44_69#_M1015_g N_A_217_69#_c_370_n 0.0142061f $X=2.095 $Y=0.755 $X2=0
+ $Y2=0
cc_206 N_A_44_69#_M1016_g N_A_217_69#_c_370_n 0.0112664f $X=2.525 $Y=0.755 $X2=0
+ $Y2=0
cc_207 N_A_44_69#_M1028_g N_A_217_69#_c_370_n 0.0112664f $X=3.115 $Y=0.755 $X2=0
+ $Y2=0
cc_208 N_A_44_69#_M1029_g N_A_217_69#_c_370_n 0.0110127f $X=3.545 $Y=0.755 $X2=0
+ $Y2=0
cc_209 N_A_44_69#_c_219_n N_A_217_69#_c_370_n 0.00475464f $X=2.02 $Y=1.495 $X2=0
+ $Y2=0
cc_210 N_A_44_69#_c_263_p N_A_217_69#_c_370_n 0.00303358f $X=3.175 $Y=1.51 $X2=0
+ $Y2=0
cc_211 N_A_44_69#_M1029_g N_A_217_69#_c_337_n 0.00466187f $X=3.545 $Y=0.755
+ $X2=0 $Y2=0
cc_212 N_A_44_69#_c_222_n N_A_217_69#_c_337_n 2.03617e-19 $X=3.515 $Y=1.51 $X2=0
+ $Y2=0
cc_213 N_A_44_69#_M1029_g N_A_217_69#_c_340_n 0.0084487f $X=3.545 $Y=0.755 $X2=0
+ $Y2=0
cc_214 N_A_44_69#_c_222_n N_A_217_69#_c_340_n 0.0160692f $X=3.515 $Y=1.51 $X2=0
+ $Y2=0
cc_215 N_A_44_69#_c_228_n N_VPWR_M1002_d 0.00526849f $X=1.85 $Y=2.425 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A_44_69#_c_228_n N_VPWR_M1007_d 0.00461511f $X=1.85 $Y=2.425 $X2=0
+ $Y2=0
cc_217 N_A_44_69#_c_218_n N_VPWR_M1007_d 0.00900444f $X=1.935 $Y=2.34 $X2=0
+ $Y2=0
cc_218 N_A_44_69#_c_228_n N_VPWR_c_622_n 0.0166722f $X=1.85 $Y=2.425 $X2=0 $Y2=0
cc_219 N_A_44_69#_M1007_g N_VPWR_c_623_n 0.0113675f $X=2.225 $Y=2.465 $X2=0
+ $Y2=0
cc_220 N_A_44_69#_M1014_g N_VPWR_c_623_n 5.6167e-19 $X=2.655 $Y=2.465 $X2=0
+ $Y2=0
cc_221 N_A_44_69#_c_228_n N_VPWR_c_623_n 0.0149622f $X=1.85 $Y=2.425 $X2=0 $Y2=0
cc_222 N_A_44_69#_M1007_g N_VPWR_c_624_n 7.21513e-19 $X=2.225 $Y=2.465 $X2=0
+ $Y2=0
cc_223 N_A_44_69#_M1014_g N_VPWR_c_624_n 0.014077f $X=2.655 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_44_69#_M1025_g N_VPWR_c_624_n 0.0141463f $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_225 N_A_44_69#_M1035_g N_VPWR_c_624_n 7.3372e-19 $X=3.515 $Y=2.465 $X2=0
+ $Y2=0
cc_226 N_A_44_69#_M1025_g N_VPWR_c_625_n 0.00486043f $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_227 N_A_44_69#_M1035_g N_VPWR_c_625_n 0.00585385f $X=3.515 $Y=2.465 $X2=0
+ $Y2=0
cc_228 N_A_44_69#_M1035_g N_VPWR_c_626_n 0.001584f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A_44_69#_M1007_g N_VPWR_c_636_n 0.00486043f $X=2.225 $Y=2.465 $X2=0
+ $Y2=0
cc_230 N_A_44_69#_M1014_g N_VPWR_c_636_n 0.00486043f $X=2.655 $Y=2.465 $X2=0
+ $Y2=0
cc_231 N_A_44_69#_c_232_n N_VPWR_c_640_n 0.0136951f $X=0.365 $Y=2.435 $X2=0
+ $Y2=0
cc_232 N_A_44_69#_M1002_s N_VPWR_c_621_n 0.0026298f $X=0.24 $Y=1.835 $X2=0 $Y2=0
cc_233 N_A_44_69#_M1007_g N_VPWR_c_621_n 0.00824727f $X=2.225 $Y=2.465 $X2=0
+ $Y2=0
cc_234 N_A_44_69#_M1014_g N_VPWR_c_621_n 0.00824727f $X=2.655 $Y=2.465 $X2=0
+ $Y2=0
cc_235 N_A_44_69#_M1025_g N_VPWR_c_621_n 0.00824727f $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_236 N_A_44_69#_M1035_g N_VPWR_c_621_n 0.0105341f $X=3.515 $Y=2.465 $X2=0
+ $Y2=0
cc_237 N_A_44_69#_c_228_n N_VPWR_c_621_n 0.0374031f $X=1.85 $Y=2.425 $X2=0 $Y2=0
cc_238 N_A_44_69#_c_232_n N_VPWR_c_621_n 0.0130717f $X=0.365 $Y=2.435 $X2=0
+ $Y2=0
cc_239 N_A_44_69#_M1015_g N_Y_c_772_n 0.00580551f $X=2.095 $Y=0.755 $X2=0 $Y2=0
cc_240 N_A_44_69#_M1016_g N_Y_c_772_n 0.0125591f $X=2.525 $Y=0.755 $X2=0 $Y2=0
cc_241 N_A_44_69#_M1028_g N_Y_c_772_n 0.0125486f $X=3.115 $Y=0.755 $X2=0 $Y2=0
cc_242 N_A_44_69#_M1029_g N_Y_c_772_n 0.00963327f $X=3.545 $Y=0.755 $X2=0 $Y2=0
cc_243 N_A_44_69#_c_263_p N_Y_c_772_n 0.0888233f $X=3.175 $Y=1.51 $X2=0 $Y2=0
cc_244 N_A_44_69#_c_222_n N_Y_c_772_n 0.0123057f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_245 N_A_44_69#_M1014_g N_Y_c_774_n 0.0128162f $X=2.655 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A_44_69#_M1025_g N_Y_c_774_n 0.0129249f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_247 N_A_44_69#_c_263_p N_Y_c_774_n 0.0574858f $X=3.175 $Y=1.51 $X2=0 $Y2=0
cc_248 N_A_44_69#_c_222_n N_Y_c_774_n 0.00243542f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_249 N_A_44_69#_M1007_g N_Y_c_775_n 6.73139e-19 $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A_44_69#_c_218_n N_Y_c_775_n 0.0056745f $X=1.935 $Y=2.34 $X2=0 $Y2=0
cc_251 N_A_44_69#_c_263_p N_Y_c_775_n 0.0155925f $X=3.175 $Y=1.51 $X2=0 $Y2=0
cc_252 N_A_44_69#_c_222_n N_Y_c_775_n 0.00296179f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_253 N_A_44_69#_M1025_g N_Y_c_773_n 5.31083e-19 $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_254 N_A_44_69#_M1028_g N_Y_c_773_n 7.31467e-19 $X=3.115 $Y=0.755 $X2=0 $Y2=0
cc_255 N_A_44_69#_M1035_g N_Y_c_773_n 0.00285752f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_256 N_A_44_69#_M1029_g N_Y_c_773_n 0.00396805f $X=3.545 $Y=0.755 $X2=0 $Y2=0
cc_257 N_A_44_69#_c_263_p N_Y_c_773_n 0.0158579f $X=3.175 $Y=1.51 $X2=0 $Y2=0
cc_258 N_A_44_69#_c_222_n N_Y_c_773_n 0.0129421f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_259 N_A_44_69#_M1035_g N_Y_c_778_n 0.013875f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A_44_69#_c_222_n N_Y_c_778_n 0.00271337f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_261 N_A_44_69#_M1035_g Y 4.43252e-19 $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A_44_69#_c_217_n N_VGND_c_905_n 0.0276344f $X=0.345 $Y=0.49 $X2=0 $Y2=0
cc_263 N_A_44_69#_c_217_n N_VGND_c_908_n 0.0185281f $X=0.345 $Y=0.49 $X2=0 $Y2=0
cc_264 N_A_44_69#_M1015_g N_VGND_c_909_n 0.00296932f $X=2.095 $Y=0.755 $X2=0
+ $Y2=0
cc_265 N_A_44_69#_M1016_g N_VGND_c_909_n 0.00296932f $X=2.525 $Y=0.755 $X2=0
+ $Y2=0
cc_266 N_A_44_69#_M1028_g N_VGND_c_909_n 0.00296932f $X=3.115 $Y=0.755 $X2=0
+ $Y2=0
cc_267 N_A_44_69#_M1029_g N_VGND_c_909_n 0.00296932f $X=3.545 $Y=0.755 $X2=0
+ $Y2=0
cc_268 N_A_44_69#_M1015_g N_VGND_c_912_n 0.00456657f $X=2.095 $Y=0.755 $X2=0
+ $Y2=0
cc_269 N_A_44_69#_M1016_g N_VGND_c_912_n 0.0042774f $X=2.525 $Y=0.755 $X2=0
+ $Y2=0
cc_270 N_A_44_69#_M1028_g N_VGND_c_912_n 0.0042774f $X=3.115 $Y=0.755 $X2=0
+ $Y2=0
cc_271 N_A_44_69#_M1029_g N_VGND_c_912_n 0.00427821f $X=3.545 $Y=0.755 $X2=0
+ $Y2=0
cc_272 N_A_44_69#_c_217_n N_VGND_c_912_n 0.013991f $X=0.345 $Y=0.49 $X2=0 $Y2=0
cc_273 N_A_44_69#_M1015_g N_A_324_45#_c_1006_n 0.0119541f $X=2.095 $Y=0.755
+ $X2=0 $Y2=0
cc_274 N_A_44_69#_M1016_g N_A_324_45#_c_1006_n 0.0110126f $X=2.525 $Y=0.755
+ $X2=0 $Y2=0
cc_275 N_A_44_69#_M1028_g N_A_324_45#_c_1006_n 0.0110126f $X=3.115 $Y=0.755
+ $X2=0 $Y2=0
cc_276 N_A_44_69#_M1029_g N_A_324_45#_c_1006_n 0.0109309f $X=3.545 $Y=0.755
+ $X2=0 $Y2=0
cc_277 N_A_217_69#_c_338_n N_C_M1006_g 4.41138e-19 $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_278 N_A_217_69#_c_339_n N_C_M1006_g 0.00308939f $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_279 N_A_217_69#_c_338_n C 0.00441862f $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_280 N_A_217_69#_c_339_n C 6.9573e-19 $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_281 N_A_217_69#_c_339_n N_C_c_481_n 0.00579295f $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_282 N_A_217_69#_M1005_g N_VPWR_c_626_n 0.00147373f $X=3.945 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_A_217_69#_M1005_g N_VPWR_c_627_n 7.34184e-19 $X=3.945 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_A_217_69#_M1018_g N_VPWR_c_627_n 0.0148745f $X=4.375 $Y=2.465 $X2=0
+ $Y2=0
cc_285 N_A_217_69#_M1023_g N_VPWR_c_627_n 0.014714f $X=4.805 $Y=2.465 $X2=0
+ $Y2=0
cc_286 N_A_217_69#_M1031_g N_VPWR_c_627_n 6.71593e-19 $X=5.235 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_A_217_69#_M1005_g N_VPWR_c_641_n 0.0054895f $X=3.945 $Y=2.465 $X2=0
+ $Y2=0
cc_288 N_A_217_69#_M1018_g N_VPWR_c_641_n 0.00486043f $X=4.375 $Y=2.465 $X2=0
+ $Y2=0
cc_289 N_A_217_69#_M1023_g N_VPWR_c_642_n 0.00486043f $X=4.805 $Y=2.465 $X2=0
+ $Y2=0
cc_290 N_A_217_69#_M1031_g N_VPWR_c_642_n 0.00486043f $X=5.235 $Y=2.465 $X2=0
+ $Y2=0
cc_291 N_A_217_69#_M1023_g N_VPWR_c_648_n 6.75557e-19 $X=4.805 $Y=2.465 $X2=0
+ $Y2=0
cc_292 N_A_217_69#_M1031_g N_VPWR_c_648_n 0.0174763f $X=5.235 $Y=2.465 $X2=0
+ $Y2=0
cc_293 N_A_217_69#_M1011_d N_VPWR_c_621_n 0.00383802f $X=1.085 $Y=1.835 $X2=0
+ $Y2=0
cc_294 N_A_217_69#_M1005_g N_VPWR_c_621_n 0.00979102f $X=3.945 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_217_69#_M1018_g N_VPWR_c_621_n 0.00824727f $X=4.375 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_217_69#_M1023_g N_VPWR_c_621_n 0.00824727f $X=4.805 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_A_217_69#_M1031_g N_VPWR_c_621_n 0.00819843f $X=5.235 $Y=2.465 $X2=0
+ $Y2=0
cc_298 N_A_217_69#_c_370_n N_Y_M1015_d 0.00336063f $X=3.87 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_299 N_A_217_69#_c_370_n N_Y_M1028_d 0.00336063f $X=3.87 $Y=0.7 $X2=0 $Y2=0
cc_300 N_A_217_69#_c_335_n N_Y_c_772_n 0.00934445f $X=1.59 $Y=1.92 $X2=0 $Y2=0
cc_301 N_A_217_69#_c_370_n N_Y_c_772_n 0.0841318f $X=3.87 $Y=0.7 $X2=0 $Y2=0
cc_302 N_A_217_69#_c_337_n N_Y_c_772_n 0.0203932f $X=3.955 $Y=1.415 $X2=0 $Y2=0
cc_303 N_A_217_69#_c_337_n N_Y_c_773_n 0.0286286f $X=3.955 $Y=1.415 $X2=0 $Y2=0
cc_304 N_A_217_69#_c_340_n N_Y_c_773_n 0.00466727f $X=5.5 $Y=1.5 $X2=0 $Y2=0
cc_305 N_A_217_69#_M1005_g N_Y_c_777_n 0.0110983f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_306 N_A_217_69#_c_337_n N_Y_c_777_n 0.00944573f $X=3.955 $Y=1.415 $X2=0 $Y2=0
cc_307 N_A_217_69#_c_338_n N_Y_c_780_n 5.42097e-19 $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_308 N_A_217_69#_M1005_g Y 0.00459077f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_309 N_A_217_69#_c_337_n Y 0.00385743f $X=3.955 $Y=1.415 $X2=0 $Y2=0
cc_310 N_A_217_69#_c_338_n Y 0.0174403f $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_311 N_A_217_69#_c_340_n Y 0.00292626f $X=5.5 $Y=1.5 $X2=0 $Y2=0
cc_312 N_A_217_69#_c_338_n Y 0.0154427f $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_313 N_A_217_69#_c_340_n Y 0.00292626f $X=5.5 $Y=1.5 $X2=0 $Y2=0
cc_314 N_A_217_69#_M1018_g N_Y_c_787_n 0.0180486f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_315 N_A_217_69#_M1023_g N_Y_c_787_n 0.0180627f $X=4.805 $Y=2.465 $X2=0 $Y2=0
cc_316 N_A_217_69#_c_338_n N_Y_c_787_n 0.0498546f $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_317 N_A_217_69#_c_340_n N_Y_c_787_n 0.00287088f $X=5.5 $Y=1.5 $X2=0 $Y2=0
cc_318 N_A_217_69#_M1031_g N_Y_c_788_n 0.0238562f $X=5.235 $Y=2.465 $X2=0 $Y2=0
cc_319 N_A_217_69#_c_338_n N_Y_c_788_n 0.0592135f $X=5.735 $Y=1.5 $X2=0 $Y2=0
cc_320 N_A_217_69#_c_340_n N_Y_c_788_n 0.0151033f $X=5.5 $Y=1.5 $X2=0 $Y2=0
cc_321 N_A_217_69#_M1005_g N_Y_c_835_n 0.0114253f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A_217_69#_c_334_n N_VGND_c_905_n 0.0116142f $X=1.225 $Y=0.49 $X2=0
+ $Y2=0
cc_323 N_A_217_69#_M1000_g N_VGND_c_909_n 0.00296932f $X=4.135 $Y=0.755 $X2=0
+ $Y2=0
cc_324 N_A_217_69#_M1012_g N_VGND_c_909_n 0.00296905f $X=4.565 $Y=0.755 $X2=0
+ $Y2=0
cc_325 N_A_217_69#_M1022_g N_VGND_c_909_n 0.00296905f $X=4.995 $Y=0.755 $X2=0
+ $Y2=0
cc_326 N_A_217_69#_M1030_g N_VGND_c_909_n 0.00296905f $X=5.425 $Y=0.755 $X2=0
+ $Y2=0
cc_327 N_A_217_69#_c_334_n N_VGND_c_909_n 0.00985379f $X=1.225 $Y=0.49 $X2=0
+ $Y2=0
cc_328 N_A_217_69#_c_336_n N_VGND_c_909_n 0.00553906f $X=1.68 $Y=0.7 $X2=0 $Y2=0
cc_329 N_A_217_69#_M1000_g N_VGND_c_912_n 0.00427821f $X=4.135 $Y=0.755 $X2=0
+ $Y2=0
cc_330 N_A_217_69#_M1012_g N_VGND_c_912_n 0.00416664f $X=4.565 $Y=0.755 $X2=0
+ $Y2=0
cc_331 N_A_217_69#_M1022_g N_VGND_c_912_n 0.00416664f $X=4.995 $Y=0.755 $X2=0
+ $Y2=0
cc_332 N_A_217_69#_M1030_g N_VGND_c_912_n 0.00456655f $X=5.425 $Y=0.755 $X2=0
+ $Y2=0
cc_333 N_A_217_69#_c_334_n N_VGND_c_912_n 0.00743302f $X=1.225 $Y=0.49 $X2=0
+ $Y2=0
cc_334 N_A_217_69#_c_336_n N_VGND_c_912_n 0.00840398f $X=1.68 $Y=0.7 $X2=0 $Y2=0
cc_335 N_A_217_69#_c_335_n N_A_324_45#_M1015_s 0.00656684f $X=1.59 $Y=1.92
+ $X2=-0.19 $Y2=-0.245
cc_336 N_A_217_69#_c_370_n N_A_324_45#_M1015_s 0.0130509f $X=3.87 $Y=0.7
+ $X2=-0.19 $Y2=-0.245
cc_337 N_A_217_69#_c_336_n N_A_324_45#_M1015_s 0.00120165f $X=1.68 $Y=0.7
+ $X2=-0.19 $Y2=-0.245
cc_338 N_A_217_69#_c_370_n N_A_324_45#_M1016_s 0.0072791f $X=3.87 $Y=0.7 $X2=0
+ $Y2=0
cc_339 N_A_217_69#_c_370_n N_A_324_45#_M1029_s 0.0121705f $X=3.87 $Y=0.7 $X2=0
+ $Y2=0
cc_340 N_A_217_69#_c_337_n N_A_324_45#_M1029_s 0.00670346f $X=3.955 $Y=1.415
+ $X2=0 $Y2=0
cc_341 N_A_217_69#_M1000_g N_A_324_45#_c_1006_n 0.0155882f $X=4.135 $Y=0.755
+ $X2=0 $Y2=0
cc_342 N_A_217_69#_M1012_g N_A_324_45#_c_1006_n 0.00862093f $X=4.565 $Y=0.755
+ $X2=0 $Y2=0
cc_343 N_A_217_69#_c_334_n N_A_324_45#_c_1006_n 0.00720715f $X=1.225 $Y=0.49
+ $X2=0 $Y2=0
cc_344 N_A_217_69#_c_370_n N_A_324_45#_c_1006_n 0.127452f $X=3.87 $Y=0.7 $X2=0
+ $Y2=0
cc_345 N_A_217_69#_c_336_n N_A_324_45#_c_1006_n 0.00622291f $X=1.68 $Y=0.7 $X2=0
+ $Y2=0
cc_346 N_A_217_69#_M1000_g N_A_324_45#_c_1025_n 0.00157086f $X=4.135 $Y=0.755
+ $X2=0 $Y2=0
cc_347 N_A_217_69#_M1012_g N_A_324_45#_c_1025_n 0.00832251f $X=4.565 $Y=0.755
+ $X2=0 $Y2=0
cc_348 N_A_217_69#_M1022_g N_A_324_45#_c_1025_n 0.0078735f $X=4.995 $Y=0.755
+ $X2=0 $Y2=0
cc_349 N_A_217_69#_M1030_g N_A_324_45#_c_1025_n 0.00130083f $X=5.425 $Y=0.755
+ $X2=0 $Y2=0
cc_350 N_A_217_69#_M1022_g N_A_324_45#_c_1007_n 0.00814149f $X=4.995 $Y=0.755
+ $X2=0 $Y2=0
cc_351 N_A_217_69#_M1030_g N_A_324_45#_c_1007_n 0.0117573f $X=5.425 $Y=0.755
+ $X2=0 $Y2=0
cc_352 N_A_217_69#_M1022_g N_A_324_45#_c_1031_n 0.00107475f $X=4.995 $Y=0.755
+ $X2=0 $Y2=0
cc_353 N_A_217_69#_M1030_g N_A_324_45#_c_1031_n 0.00668111f $X=5.425 $Y=0.755
+ $X2=0 $Y2=0
cc_354 N_A_217_69#_M1012_g N_A_324_45#_c_1008_n 0.00152423f $X=4.565 $Y=0.755
+ $X2=0 $Y2=0
cc_355 N_A_217_69#_M1022_g N_A_324_45#_c_1008_n 0.00182901f $X=4.995 $Y=0.755
+ $X2=0 $Y2=0
cc_356 N_A_217_69#_M1030_g N_A_842_67#_c_1063_n 0.0170713f $X=5.425 $Y=0.755
+ $X2=0 $Y2=0
cc_357 N_A_217_69#_c_339_n N_A_842_67#_c_1063_n 0.00996728f $X=5.735 $Y=1.5
+ $X2=0 $Y2=0
cc_358 N_A_217_69#_M1030_g N_A_842_67#_c_1064_n 0.00315269f $X=5.425 $Y=0.755
+ $X2=0 $Y2=0
cc_359 N_A_217_69#_M1030_g N_A_842_67#_c_1066_n 7.19256e-19 $X=5.425 $Y=0.755
+ $X2=0 $Y2=0
cc_360 N_A_217_69#_M1000_g N_A_842_67#_c_1067_n 5.53292e-19 $X=4.135 $Y=0.755
+ $X2=0 $Y2=0
cc_361 N_A_217_69#_c_337_n N_A_842_67#_c_1067_n 0.0046083f $X=3.955 $Y=1.415
+ $X2=0 $Y2=0
cc_362 N_A_217_69#_c_338_n N_A_842_67#_c_1067_n 0.0152507f $X=5.735 $Y=1.5 $X2=0
+ $Y2=0
cc_363 N_A_217_69#_c_340_n N_A_842_67#_c_1067_n 0.00294542f $X=5.5 $Y=1.5 $X2=0
+ $Y2=0
cc_364 N_A_217_69#_M1012_g N_A_842_67#_c_1068_n 0.0110129f $X=4.565 $Y=0.755
+ $X2=0 $Y2=0
cc_365 N_A_217_69#_M1022_g N_A_842_67#_c_1068_n 0.011531f $X=4.995 $Y=0.755
+ $X2=0 $Y2=0
cc_366 N_A_217_69#_c_338_n N_A_842_67#_c_1068_n 0.106265f $X=5.735 $Y=1.5 $X2=0
+ $Y2=0
cc_367 N_A_217_69#_c_340_n N_A_842_67#_c_1068_n 0.00290124f $X=5.5 $Y=1.5 $X2=0
+ $Y2=0
cc_368 N_A_217_69#_c_340_n N_A_842_67#_c_1069_n 0.00294793f $X=5.5 $Y=1.5 $X2=0
+ $Y2=0
cc_369 N_C_M1033_g N_D_M1003_g 0.0286582f $X=7.855 $Y=2.465 $X2=0 $Y2=0
cc_370 N_C_c_479_n N_D_c_552_n 0.0147597f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_371 C D 0.0242185f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_372 N_C_c_481_n D 3.61226e-19 $X=7.885 $Y=1.35 $X2=0 $Y2=0
cc_373 C N_D_c_560_n 0.00128571f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_374 N_C_c_481_n N_D_c_560_n 0.0177132f $X=7.885 $Y=1.35 $X2=0 $Y2=0
cc_375 N_C_M1006_g N_VPWR_c_628_n 7.37337e-19 $X=6.565 $Y=2.465 $X2=0 $Y2=0
cc_376 N_C_M1009_g N_VPWR_c_628_n 0.0141064f $X=6.995 $Y=2.465 $X2=0 $Y2=0
cc_377 N_C_M1020_g N_VPWR_c_628_n 0.0140168f $X=7.425 $Y=2.465 $X2=0 $Y2=0
cc_378 N_C_M1033_g N_VPWR_c_628_n 7.21513e-19 $X=7.855 $Y=2.465 $X2=0 $Y2=0
cc_379 N_C_M1020_g N_VPWR_c_629_n 0.00486043f $X=7.425 $Y=2.465 $X2=0 $Y2=0
cc_380 N_C_M1033_g N_VPWR_c_629_n 0.00486043f $X=7.855 $Y=2.465 $X2=0 $Y2=0
cc_381 N_C_M1020_g N_VPWR_c_630_n 7.21513e-19 $X=7.425 $Y=2.465 $X2=0 $Y2=0
cc_382 N_C_M1033_g N_VPWR_c_630_n 0.0139811f $X=7.855 $Y=2.465 $X2=0 $Y2=0
cc_383 N_C_M1006_g N_VPWR_c_638_n 0.00585385f $X=6.565 $Y=2.465 $X2=0 $Y2=0
cc_384 N_C_M1009_g N_VPWR_c_638_n 0.00486043f $X=6.995 $Y=2.465 $X2=0 $Y2=0
cc_385 N_C_M1006_g N_VPWR_c_648_n 0.00349091f $X=6.565 $Y=2.465 $X2=0 $Y2=0
cc_386 N_C_M1006_g N_VPWR_c_621_n 0.0118331f $X=6.565 $Y=2.465 $X2=0 $Y2=0
cc_387 N_C_M1009_g N_VPWR_c_621_n 0.00824727f $X=6.995 $Y=2.465 $X2=0 $Y2=0
cc_388 N_C_M1020_g N_VPWR_c_621_n 0.00824727f $X=7.425 $Y=2.465 $X2=0 $Y2=0
cc_389 N_C_M1033_g N_VPWR_c_621_n 0.00824727f $X=7.855 $Y=2.465 $X2=0 $Y2=0
cc_390 N_C_M1009_g N_Y_c_779_n 0.016691f $X=6.995 $Y=2.465 $X2=0 $Y2=0
cc_391 N_C_M1020_g N_Y_c_779_n 0.0167157f $X=7.425 $Y=2.465 $X2=0 $Y2=0
cc_392 C N_Y_c_779_n 0.0505913f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_393 N_C_c_481_n N_Y_c_779_n 0.00238281f $X=7.885 $Y=1.35 $X2=0 $Y2=0
cc_394 N_C_M1006_g N_Y_c_780_n 0.0213625f $X=6.565 $Y=2.465 $X2=0 $Y2=0
cc_395 C N_Y_c_780_n 0.0481976f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_396 N_C_c_481_n N_Y_c_780_n 0.00743395f $X=7.885 $Y=1.35 $X2=0 $Y2=0
cc_397 N_C_M1033_g N_Y_c_781_n 0.0166442f $X=7.855 $Y=2.465 $X2=0 $Y2=0
cc_398 C N_Y_c_781_n 0.0204479f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_399 N_C_c_481_n N_Y_c_781_n 7.97581e-19 $X=7.885 $Y=1.35 $X2=0 $Y2=0
cc_400 C N_Y_c_783_n 0.0159743f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_401 N_C_c_481_n N_Y_c_783_n 0.00244789f $X=7.885 $Y=1.35 $X2=0 $Y2=0
cc_402 N_C_c_479_n N_VGND_c_906_n 0.00121531f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_403 N_C_c_473_n N_VGND_c_909_n 0.00369121f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_404 N_C_c_475_n N_VGND_c_909_n 0.00369121f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_405 N_C_c_477_n N_VGND_c_909_n 0.00370545f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_406 N_C_c_479_n N_VGND_c_909_n 0.00585385f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_407 N_C_c_473_n N_VGND_c_912_n 0.00677279f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_408 N_C_c_475_n N_VGND_c_912_n 0.00537312f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_409 N_C_c_477_n N_VGND_c_912_n 0.0054347f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_410 N_C_c_479_n N_VGND_c_912_n 0.00653014f $X=7.885 $Y=1.185 $X2=0 $Y2=0
cc_411 N_C_c_473_n N_A_842_67#_c_1063_n 0.00450822f $X=6.595 $Y=1.185 $X2=0
+ $Y2=0
cc_412 C N_A_842_67#_c_1063_n 0.0039228f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_413 N_C_c_481_n N_A_842_67#_c_1063_n 0.00111826f $X=7.885 $Y=1.35 $X2=0 $Y2=0
cc_414 N_C_c_473_n N_A_842_67#_c_1064_n 0.00434268f $X=6.595 $Y=1.185 $X2=0
+ $Y2=0
cc_415 N_C_c_473_n N_A_842_67#_c_1065_n 0.0115125f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_416 N_C_c_475_n N_A_842_67#_c_1065_n 0.00917005f $X=7.025 $Y=1.185 $X2=0
+ $Y2=0
cc_417 N_C_c_477_n N_A_842_67#_c_1065_n 0.0105488f $X=7.455 $Y=1.185 $X2=0 $Y2=0
cc_418 N_C_c_481_n N_A_842_67#_c_1065_n 4.14624e-19 $X=7.885 $Y=1.35 $X2=0 $Y2=0
cc_419 N_C_c_475_n N_A_842_67#_c_1091_n 8.71093e-19 $X=7.025 $Y=1.185 $X2=0
+ $Y2=0
cc_420 N_C_c_477_n N_A_842_67#_c_1091_n 0.00433647f $X=7.455 $Y=1.185 $X2=0
+ $Y2=0
cc_421 N_C_c_473_n N_A_1251_47#_c_1125_n 0.0127195f $X=6.595 $Y=1.185 $X2=0
+ $Y2=0
cc_422 N_C_c_475_n N_A_1251_47#_c_1125_n 0.0126726f $X=7.025 $Y=1.185 $X2=0
+ $Y2=0
cc_423 C N_A_1251_47#_c_1125_n 0.11196f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_424 N_C_c_481_n N_A_1251_47#_c_1125_n 0.00797512f $X=7.885 $Y=1.35 $X2=0
+ $Y2=0
cc_425 N_C_c_477_n N_A_1251_47#_c_1129_n 0.0092537f $X=7.455 $Y=1.185 $X2=0
+ $Y2=0
cc_426 N_C_c_479_n N_A_1251_47#_c_1129_n 0.0100475f $X=7.885 $Y=1.185 $X2=0
+ $Y2=0
cc_427 N_C_c_481_n N_A_1251_47#_c_1129_n 0.00240196f $X=7.885 $Y=1.35 $X2=0
+ $Y2=0
cc_428 N_C_c_481_n N_A_1251_47#_c_1132_n 0.00243924f $X=7.885 $Y=1.35 $X2=0
+ $Y2=0
cc_429 N_D_M1003_g N_VPWR_c_630_n 0.0139811f $X=8.285 $Y=2.465 $X2=0 $Y2=0
cc_430 N_D_M1021_g N_VPWR_c_630_n 7.21513e-19 $X=8.715 $Y=2.465 $X2=0 $Y2=0
cc_431 N_D_M1003_g N_VPWR_c_631_n 7.21513e-19 $X=8.285 $Y=2.465 $X2=0 $Y2=0
cc_432 N_D_M1021_g N_VPWR_c_631_n 0.0140168f $X=8.715 $Y=2.465 $X2=0 $Y2=0
cc_433 N_D_M1026_g N_VPWR_c_631_n 0.0140861f $X=9.145 $Y=2.465 $X2=0 $Y2=0
cc_434 N_D_M1027_g N_VPWR_c_631_n 7.3372e-19 $X=9.575 $Y=2.465 $X2=0 $Y2=0
cc_435 N_D_M1027_g N_VPWR_c_633_n 0.00773581f $X=9.575 $Y=2.465 $X2=0 $Y2=0
cc_436 D N_VPWR_c_633_n 0.0149289f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_437 N_D_c_560_n N_VPWR_c_633_n 0.00535627f $X=9.735 $Y=1.35 $X2=0 $Y2=0
cc_438 N_D_M1003_g N_VPWR_c_643_n 0.00486043f $X=8.285 $Y=2.465 $X2=0 $Y2=0
cc_439 N_D_M1021_g N_VPWR_c_643_n 0.00486043f $X=8.715 $Y=2.465 $X2=0 $Y2=0
cc_440 N_D_M1026_g N_VPWR_c_644_n 0.00486043f $X=9.145 $Y=2.465 $X2=0 $Y2=0
cc_441 N_D_M1027_g N_VPWR_c_644_n 0.00585385f $X=9.575 $Y=2.465 $X2=0 $Y2=0
cc_442 N_D_M1003_g N_VPWR_c_621_n 0.00824727f $X=8.285 $Y=2.465 $X2=0 $Y2=0
cc_443 N_D_M1021_g N_VPWR_c_621_n 0.00824727f $X=8.715 $Y=2.465 $X2=0 $Y2=0
cc_444 N_D_M1026_g N_VPWR_c_621_n 0.00824727f $X=9.145 $Y=2.465 $X2=0 $Y2=0
cc_445 N_D_M1027_g N_VPWR_c_621_n 0.0114685f $X=9.575 $Y=2.465 $X2=0 $Y2=0
cc_446 N_D_M1003_g N_Y_c_781_n 0.0166442f $X=8.285 $Y=2.465 $X2=0 $Y2=0
cc_447 D N_Y_c_781_n 0.0144584f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_448 N_D_M1021_g N_Y_c_782_n 0.0166442f $X=8.715 $Y=2.465 $X2=0 $Y2=0
cc_449 N_D_M1026_g N_Y_c_782_n 0.0164008f $X=9.145 $Y=2.465 $X2=0 $Y2=0
cc_450 N_D_M1027_g N_Y_c_782_n 0.00449417f $X=9.575 $Y=2.465 $X2=0 $Y2=0
cc_451 D N_Y_c_782_n 0.0690881f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_452 N_D_c_560_n N_Y_c_782_n 0.0048307f $X=9.735 $Y=1.35 $X2=0 $Y2=0
cc_453 D N_Y_c_784_n 0.0159743f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_454 N_D_c_560_n N_Y_c_784_n 0.00244789f $X=9.735 $Y=1.35 $X2=0 $Y2=0
cc_455 N_D_c_552_n N_VGND_c_906_n 0.01106f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_456 N_D_c_554_n N_VGND_c_906_n 0.00986738f $X=8.745 $Y=1.185 $X2=0 $Y2=0
cc_457 N_D_c_556_n N_VGND_c_906_n 5.72987e-19 $X=9.175 $Y=1.185 $X2=0 $Y2=0
cc_458 N_D_c_554_n N_VGND_c_907_n 5.79734e-19 $X=8.745 $Y=1.185 $X2=0 $Y2=0
cc_459 N_D_c_556_n N_VGND_c_907_n 0.00996732f $X=9.175 $Y=1.185 $X2=0 $Y2=0
cc_460 N_D_c_558_n N_VGND_c_907_n 0.011549f $X=9.605 $Y=1.185 $X2=0 $Y2=0
cc_461 N_D_c_552_n N_VGND_c_909_n 0.00486043f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_462 N_D_c_554_n N_VGND_c_910_n 0.00486043f $X=8.745 $Y=1.185 $X2=0 $Y2=0
cc_463 N_D_c_556_n N_VGND_c_910_n 0.00486043f $X=9.175 $Y=1.185 $X2=0 $Y2=0
cc_464 N_D_c_558_n N_VGND_c_911_n 0.00486043f $X=9.605 $Y=1.185 $X2=0 $Y2=0
cc_465 N_D_c_552_n N_VGND_c_912_n 0.00460797f $X=8.315 $Y=1.185 $X2=0 $Y2=0
cc_466 N_D_c_554_n N_VGND_c_912_n 0.00458264f $X=8.745 $Y=1.185 $X2=0 $Y2=0
cc_467 N_D_c_556_n N_VGND_c_912_n 0.00458264f $X=9.175 $Y=1.185 $X2=0 $Y2=0
cc_468 N_D_c_558_n N_VGND_c_912_n 0.00551524f $X=9.605 $Y=1.185 $X2=0 $Y2=0
cc_469 N_D_c_552_n N_A_1251_47#_c_1133_n 0.00978727f $X=8.315 $Y=1.185 $X2=0
+ $Y2=0
cc_470 N_D_c_554_n N_A_1251_47#_c_1133_n 0.00978727f $X=8.745 $Y=1.185 $X2=0
+ $Y2=0
cc_471 D N_A_1251_47#_c_1133_n 0.0405304f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_472 N_D_c_560_n N_A_1251_47#_c_1133_n 0.00240196f $X=9.735 $Y=1.35 $X2=0
+ $Y2=0
cc_473 N_D_c_556_n N_A_1251_47#_c_1137_n 0.00974071f $X=9.175 $Y=1.185 $X2=0
+ $Y2=0
cc_474 N_D_c_558_n N_A_1251_47#_c_1137_n 0.00978727f $X=9.605 $Y=1.185 $X2=0
+ $Y2=0
cc_475 D N_A_1251_47#_c_1137_n 0.0574879f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_476 N_D_c_560_n N_A_1251_47#_c_1137_n 0.00651526f $X=9.735 $Y=1.35 $X2=0
+ $Y2=0
cc_477 D N_A_1251_47#_c_1141_n 0.0141881f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_478 N_D_c_560_n N_A_1251_47#_c_1141_n 0.00249225f $X=9.735 $Y=1.35 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_621_n N_Y_M1007_s 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_480 N_VPWR_c_621_n N_Y_M1025_s 0.00432284f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_481 N_VPWR_c_621_n N_Y_M1005_d 0.00380103f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_482 N_VPWR_c_621_n N_Y_M1023_d 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_483 N_VPWR_c_621_n N_Y_M1006_s 0.00397496f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_484 N_VPWR_c_621_n N_Y_M1020_s 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_485 N_VPWR_c_621_n N_Y_M1003_d 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_486 N_VPWR_c_621_n N_Y_M1026_d 0.00432284f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_487 N_VPWR_c_636_n N_Y_c_865_n 0.0124525f $X=2.705 $Y=3.33 $X2=0 $Y2=0
cc_488 N_VPWR_c_621_n N_Y_c_865_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_489 N_VPWR_M1014_d N_Y_c_774_n 0.00176461f $X=2.73 $Y=1.835 $X2=0 $Y2=0
cc_490 N_VPWR_c_624_n N_Y_c_774_n 0.0170777f $X=2.87 $Y=2.2 $X2=0 $Y2=0
cc_491 N_VPWR_c_625_n N_Y_c_869_n 0.0135169f $X=3.595 $Y=3.33 $X2=0 $Y2=0
cc_492 N_VPWR_c_621_n N_Y_c_869_n 0.00847534f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_493 N_VPWR_M1035_d N_Y_c_777_n 0.00129688f $X=3.59 $Y=1.835 $X2=0 $Y2=0
cc_494 N_VPWR_M1035_d N_Y_c_778_n 4.57098e-19 $X=3.59 $Y=1.835 $X2=0 $Y2=0
cc_495 N_VPWR_c_626_n N_Y_c_778_n 0.013469f $X=3.73 $Y=2.28 $X2=0 $Y2=0
cc_496 N_VPWR_c_642_n N_Y_c_874_n 0.0124525f $X=5.285 $Y=3.33 $X2=0 $Y2=0
cc_497 N_VPWR_c_621_n N_Y_c_874_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_498 N_VPWR_c_638_n N_Y_c_876_n 0.0138717f $X=7.045 $Y=3.33 $X2=0 $Y2=0
cc_499 N_VPWR_c_621_n N_Y_c_876_n 0.00886411f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_500 N_VPWR_M1009_d N_Y_c_779_n 0.00178786f $X=7.07 $Y=1.835 $X2=0 $Y2=0
cc_501 N_VPWR_c_628_n N_Y_c_779_n 0.0175857f $X=7.21 $Y=2.2 $X2=0 $Y2=0
cc_502 N_VPWR_M1031_s N_Y_c_780_n 0.0136665f $X=5.31 $Y=1.835 $X2=0 $Y2=0
cc_503 N_VPWR_c_648_n N_Y_c_780_n 0.0392272f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_504 N_VPWR_c_629_n N_Y_c_882_n 0.0124525f $X=7.905 $Y=3.33 $X2=0 $Y2=0
cc_505 N_VPWR_c_621_n N_Y_c_882_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_506 N_VPWR_M1033_d N_Y_c_781_n 0.00178786f $X=7.93 $Y=1.835 $X2=0 $Y2=0
cc_507 N_VPWR_c_630_n N_Y_c_781_n 0.0175857f $X=8.07 $Y=2.2 $X2=0 $Y2=0
cc_508 N_VPWR_c_643_n N_Y_c_886_n 0.0124525f $X=8.765 $Y=3.33 $X2=0 $Y2=0
cc_509 N_VPWR_c_621_n N_Y_c_886_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_510 N_VPWR_M1021_s N_Y_c_782_n 0.00178786f $X=8.79 $Y=1.835 $X2=0 $Y2=0
cc_511 N_VPWR_c_631_n N_Y_c_782_n 0.0175857f $X=8.93 $Y=2.2 $X2=0 $Y2=0
cc_512 N_VPWR_c_633_n N_Y_c_782_n 0.00166817f $X=9.79 $Y=1.98 $X2=0 $Y2=0
cc_513 N_VPWR_c_644_n N_Y_c_891_n 0.0135169f $X=9.655 $Y=3.33 $X2=0 $Y2=0
cc_514 N_VPWR_c_621_n N_Y_c_891_n 0.00847534f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_515 N_VPWR_M1018_s N_Y_c_787_n 0.00180346f $X=4.45 $Y=1.835 $X2=0 $Y2=0
cc_516 N_VPWR_c_627_n N_Y_c_787_n 0.0179414f $X=4.59 $Y=2.375 $X2=0 $Y2=0
cc_517 N_VPWR_M1031_s N_Y_c_788_n 0.0129322f $X=5.31 $Y=1.835 $X2=0 $Y2=0
cc_518 N_VPWR_c_648_n N_Y_c_788_n 0.0472237f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_519 N_VPWR_c_641_n N_Y_c_835_n 0.015688f $X=4.425 $Y=3.33 $X2=0 $Y2=0
cc_520 N_VPWR_c_621_n N_Y_c_835_n 0.00984745f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_521 N_Y_c_772_n N_A_324_45#_M1016_s 0.00448941f $X=3.52 $Y=1.085 $X2=0 $Y2=0
cc_522 N_Y_c_772_n N_A_324_45#_M1029_s 0.00226183f $X=3.52 $Y=1.085 $X2=0 $Y2=0
cc_523 N_Y_M1015_d N_A_324_45#_c_1006_n 0.001775f $X=2.17 $Y=0.335 $X2=0 $Y2=0
cc_524 N_Y_M1028_d N_A_324_45#_c_1006_n 0.001775f $X=3.19 $Y=0.335 $X2=0 $Y2=0
cc_525 N_Y_c_780_n N_A_842_67#_c_1063_n 0.00805696f $X=6.875 $Y=1.815 $X2=0
+ $Y2=0
cc_526 N_Y_c_781_n N_A_1251_47#_c_1143_n 0.00567402f $X=8.405 $Y=1.815 $X2=0
+ $Y2=0
cc_527 N_VGND_c_912_n N_A_324_45#_M1015_s 0.00248021f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_528 N_VGND_c_912_n N_A_324_45#_M1016_s 0.00238607f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_529 N_VGND_c_912_n N_A_324_45#_M1029_s 0.00238607f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_530 N_VGND_c_905_n N_A_324_45#_c_1006_n 0.00213148f $X=0.795 $Y=0.47 $X2=0
+ $Y2=0
cc_531 N_VGND_c_909_n N_A_324_45#_c_1006_n 0.192188f $X=8.365 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_912_n N_A_324_45#_c_1006_n 0.109638f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_c_909_n N_A_324_45#_c_1007_n 0.0533441f $X=8.365 $Y=0 $X2=0 $Y2=0
cc_534 N_VGND_c_912_n N_A_324_45#_c_1007_n 0.0296799f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_c_909_n N_A_324_45#_c_1008_n 0.023347f $X=8.365 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_912_n N_A_324_45#_c_1008_n 0.0125753f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_537 N_VGND_c_912_n N_A_842_67#_M1001_d 0.00227218f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_912_n N_A_842_67#_M1017_d 0.00253234f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_c_909_n N_A_842_67#_c_1065_n 0.0607734f $X=8.365 $Y=0 $X2=0 $Y2=0
cc_540 N_VGND_c_912_n N_A_842_67#_c_1065_n 0.0494948f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_c_909_n N_A_842_67#_c_1066_n 0.0090292f $X=8.365 $Y=0 $X2=0 $Y2=0
cc_542 N_VGND_c_912_n N_A_842_67#_c_1066_n 0.00642551f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_c_909_n N_A_842_67#_c_1091_n 0.011012f $X=8.365 $Y=0 $X2=0 $Y2=0
cc_544 N_VGND_c_912_n N_A_842_67#_c_1091_n 0.00950762f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_545 N_VGND_c_912_n N_A_1251_47#_M1001_s 0.0021945f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_546 N_VGND_c_912_n N_A_1251_47#_M1013_s 0.00228852f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_547 N_VGND_c_912_n N_A_1251_47#_M1019_s 0.00276017f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_548 N_VGND_c_912_n N_A_1251_47#_M1010_d 0.0028988f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_549 N_VGND_c_912_n N_A_1251_47#_M1034_d 0.00317907f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_550 N_VGND_c_912_n N_A_1251_47#_c_1129_n 0.00709098f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_551 N_VGND_c_909_n N_A_1251_47#_c_1150_n 0.0128073f $X=8.365 $Y=0 $X2=0 $Y2=0
cc_552 N_VGND_c_912_n N_A_1251_47#_c_1150_n 0.00769778f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_M1008_s N_A_1251_47#_c_1133_n 0.0032793f $X=8.39 $Y=0.235 $X2=0
+ $Y2=0
cc_554 N_VGND_c_906_n N_A_1251_47#_c_1133_n 0.0167297f $X=8.53 $Y=0.525 $X2=0
+ $Y2=0
cc_555 N_VGND_c_912_n N_A_1251_47#_c_1133_n 0.0106723f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_556 N_VGND_c_910_n N_A_1251_47#_c_1155_n 0.0120977f $X=9.225 $Y=0 $X2=0 $Y2=0
cc_557 N_VGND_c_912_n N_A_1251_47#_c_1155_n 0.00691495f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_558 N_VGND_M1024_s N_A_1251_47#_c_1137_n 0.0032793f $X=9.25 $Y=0.235 $X2=0
+ $Y2=0
cc_559 N_VGND_c_907_n N_A_1251_47#_c_1137_n 0.0167297f $X=9.39 $Y=0.525 $X2=0
+ $Y2=0
cc_560 N_VGND_c_912_n N_A_1251_47#_c_1137_n 0.0110118f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_561 N_VGND_c_911_n N_A_1251_47#_c_1160_n 0.0135387f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_562 N_VGND_c_912_n N_A_1251_47#_c_1160_n 0.00769778f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_563 N_A_324_45#_c_1006_n N_A_842_67#_M1000_s 0.00280802f $X=4.615 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_564 N_A_324_45#_c_1007_n N_A_842_67#_M1022_s 0.00278395f $X=5.475 $Y=0.34
+ $X2=0 $Y2=0
cc_565 N_A_324_45#_M1030_d N_A_842_67#_c_1063_n 0.00339163f $X=5.5 $Y=0.335
+ $X2=0 $Y2=0
cc_566 N_A_324_45#_c_1007_n N_A_842_67#_c_1063_n 0.00342117f $X=5.475 $Y=0.34
+ $X2=0 $Y2=0
cc_567 N_A_324_45#_c_1031_n N_A_842_67#_c_1063_n 0.018529f $X=5.64 $Y=0.625
+ $X2=0 $Y2=0
cc_568 N_A_324_45#_c_1031_n N_A_842_67#_c_1064_n 0.0207216f $X=5.64 $Y=0.625
+ $X2=0 $Y2=0
cc_569 N_A_324_45#_c_1007_n N_A_842_67#_c_1066_n 0.0106159f $X=5.475 $Y=0.34
+ $X2=0 $Y2=0
cc_570 N_A_324_45#_c_1031_n N_A_842_67#_c_1066_n 0.00813636f $X=5.64 $Y=0.625
+ $X2=0 $Y2=0
cc_571 N_A_324_45#_c_1006_n N_A_842_67#_c_1067_n 0.00639842f $X=4.615 $Y=0.35
+ $X2=0 $Y2=0
cc_572 N_A_324_45#_M1012_d N_A_842_67#_c_1068_n 0.00177068f $X=4.64 $Y=0.335
+ $X2=0 $Y2=0
cc_573 N_A_324_45#_c_1006_n N_A_842_67#_c_1068_n 0.00296726f $X=4.615 $Y=0.35
+ $X2=0 $Y2=0
cc_574 N_A_324_45#_c_1025_n N_A_842_67#_c_1068_n 0.0171014f $X=4.78 $Y=0.46
+ $X2=0 $Y2=0
cc_575 N_A_324_45#_c_1007_n N_A_842_67#_c_1068_n 0.0028551f $X=5.475 $Y=0.34
+ $X2=0 $Y2=0
cc_576 N_A_324_45#_c_1007_n N_A_842_67#_c_1069_n 0.00540831f $X=5.475 $Y=0.34
+ $X2=0 $Y2=0
cc_577 N_A_842_67#_c_1065_n N_A_1251_47#_M1001_s 0.0058172f $X=7.515 $Y=0.415
+ $X2=-0.19 $Y2=-0.245
cc_578 N_A_842_67#_c_1065_n N_A_1251_47#_M1013_s 0.00350443f $X=7.515 $Y=0.415
+ $X2=0 $Y2=0
cc_579 N_A_842_67#_M1001_d N_A_1251_47#_c_1125_n 0.00336306f $X=6.67 $Y=0.235
+ $X2=0 $Y2=0
cc_580 N_A_842_67#_c_1063_n N_A_1251_47#_c_1125_n 0.00608282f $X=5.93 $Y=1.102
+ $X2=0 $Y2=0
cc_581 N_A_842_67#_c_1064_n N_A_1251_47#_c_1125_n 0.0205044f $X=6.015 $Y=0.96
+ $X2=0 $Y2=0
cc_582 N_A_842_67#_c_1065_n N_A_1251_47#_c_1125_n 0.0560049f $X=7.515 $Y=0.415
+ $X2=0 $Y2=0
cc_583 N_A_842_67#_M1017_d N_A_1251_47#_c_1129_n 0.0032793f $X=7.53 $Y=0.235
+ $X2=0 $Y2=0
cc_584 N_A_842_67#_c_1065_n N_A_1251_47#_c_1129_n 0.00476298f $X=7.515 $Y=0.415
+ $X2=0 $Y2=0
cc_585 N_A_842_67#_c_1091_n N_A_1251_47#_c_1129_n 0.0136103f $X=7.645 $Y=0.415
+ $X2=0 $Y2=0
