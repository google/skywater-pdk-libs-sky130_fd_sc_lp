* File: sky130_fd_sc_lp__o21a_lp.pex.spice
* Created: Fri Aug 28 11:04:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21A_LP%A1 2 5 7 9 10 11 15
c34 10 0 2.37971e-20 $X=0.24 $Y=1.295
r35 15 17 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.425 $Y=1.34
+ $X2=0.425 $Y2=1.175
r36 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.34 $X2=0.385 $Y2=1.34
r37 11 16 8.8128 $w=4.23e-07 $l=3.25e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.34
r38 10 16 1.22023 $w=4.23e-07 $l=4.5e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.34
r39 7 9 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.605 $Y=1.97
+ $X2=0.605 $Y2=2.545
r40 5 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.495 $Y=0.495
+ $X2=0.495 $Y2=1.175
r41 2 7 45.5759 $w=3.49e-07 $l=4.10244e-07 $layer=POLY_cond $X=0.425 $Y=1.64
+ $X2=0.605 $Y2=1.97
r42 1 15 5.42589 $w=4.1e-07 $l=4e-08 $layer=POLY_cond $X=0.425 $Y=1.38 $X2=0.425
+ $Y2=1.34
r43 1 2 35.2683 $w=4.1e-07 $l=2.6e-07 $layer=POLY_cond $X=0.425 $Y=1.38
+ $X2=0.425 $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_LP%A2 3 7 9 11 12 13 14 15 16 23
c49 23 0 6.44844e-20 $X=1.035 $Y=1.345
c50 11 0 1.91533e-19 $X=1.095 $Y=1.745
c51 3 0 1.65657e-19 $X=1.005 $Y=0.495
r52 23 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.345
+ $X2=1.035 $Y2=1.51
r53 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.345
+ $X2=1.035 $Y2=1.18
r54 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.035
+ $Y=1.345 $X2=1.035 $Y2=1.345
r55 15 16 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.092 $Y=2.405
+ $X2=1.092 $Y2=2.775
r56 14 15 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.092 $Y=2.035
+ $X2=1.092 $Y2=2.405
r57 13 14 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.092 $Y=1.665
+ $X2=1.092 $Y2=2.035
r58 13 24 8.28723 $w=4.43e-07 $l=3.2e-07 $layer=LI1_cond $X=1.092 $Y=1.665
+ $X2=1.092 $Y2=1.345
r59 12 24 1.29488 $w=4.43e-07 $l=5e-08 $layer=LI1_cond $X=1.092 $Y=1.295
+ $X2=1.092 $Y2=1.345
r60 11 26 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=1.045 $Y=1.745
+ $X2=1.045 $Y2=1.51
r61 7 11 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.095 $Y=1.87
+ $X2=1.095 $Y2=1.745
r62 7 9 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.095 $Y=1.87
+ $X2=1.095 $Y2=2.545
r63 3 25 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=1.005 $Y=0.495
+ $X2=1.005 $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_LP%B1 3 7 9 16
c38 9 0 2.39711e-20 $X=1.68 $Y=1.295
c39 7 0 6.44844e-20 $X=1.925 $Y=2.545
r40 14 16 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.66 $Y=1.34
+ $X2=1.925 $Y2=1.34
r41 11 14 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.515 $Y=1.34
+ $X2=1.66 $Y2=1.34
r42 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=1.34 $X2=1.66 $Y2=1.34
r43 5 16 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.505
+ $X2=1.925 $Y2=1.34
r44 5 7 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.925 $Y=1.505
+ $X2=1.925 $Y2=2.545
r45 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.175
+ $X2=1.515 $Y2=1.34
r46 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.515 $Y=1.175
+ $X2=1.515 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_LP%A_244_409# 1 2 9 13 17 23 26 29 35 37 38 40
+ 41 42 49 50
c73 42 0 1.17889e-19 $X=2.175 $Y=0.91
c74 38 0 1.91533e-19 $X=1.825 $Y=1.77
r75 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=0.99 $X2=2.52 $Y2=0.99
r76 42 47 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.91
+ $X2=2.09 $Y2=0.91
r77 41 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=0.91
+ $X2=2.52 $Y2=0.91
r78 41 42 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.355 $Y=0.91
+ $X2=2.175 $Y2=0.91
r79 39 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=0.995
+ $X2=2.09 $Y2=0.91
r80 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.09 $Y=0.995
+ $X2=2.09 $Y2=1.685
r81 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.005 $Y=1.77
+ $X2=2.09 $Y2=1.685
r82 37 38 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.005 $Y=1.77
+ $X2=1.825 $Y2=1.77
r83 33 47 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.73 $Y=0.91
+ $X2=2.09 $Y2=0.91
r84 33 35 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.73 $Y=0.825
+ $X2=1.73 $Y2=0.495
r85 29 31 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.66 $Y=2.19 $X2=1.66
+ $Y2=2.9
r86 27 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.66 $Y=1.855
+ $X2=1.825 $Y2=1.77
r87 27 29 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.66 $Y=1.855
+ $X2=1.66 $Y2=2.19
r88 25 50 53.3155 $w=3.55e-07 $l=3.28e-07 $layer=POLY_cond $X=2.507 $Y=1.318
+ $X2=2.507 $Y2=0.99
r89 25 26 33.8903 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=2.507 $Y=1.318
+ $X2=2.507 $Y2=1.495
r90 22 50 2.43821 $w=3.55e-07 $l=1.5e-08 $layer=POLY_cond $X=2.507 $Y=0.975
+ $X2=2.507 $Y2=0.99
r91 22 23 183.57 $w=1.5e-07 $l=3.58e-07 $layer=POLY_cond $X=2.507 $Y=0.9
+ $X2=2.865 $Y2=0.9
r92 19 22 1.02553 $w=1.5e-07 $l=2e-09 $layer=POLY_cond $X=2.505 $Y=0.9 $X2=2.507
+ $Y2=0.9
r93 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=0.825
+ $X2=2.865 $Y2=0.9
r94 15 17 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.865 $Y=0.825
+ $X2=2.865 $Y2=0.445
r95 11 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=0.825
+ $X2=2.505 $Y2=0.9
r96 11 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.505 $Y=0.825
+ $X2=2.505 $Y2=0.445
r97 9 26 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.455 $Y=2.545
+ $X2=2.455 $Y2=1.495
r98 2 31 400 $w=1.7e-07 $l=1.05225e-06 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=2.045 $X2=1.66 $Y2=2.9
r99 2 29 400 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=2.045 $X2=1.66 $Y2=2.19
r100 1 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.285 $X2=1.73 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_LP%VPWR 1 2 7 9 15 19 21 31 32 38
r34 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 32 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.19 $Y2=3.33
r39 29 31 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 25 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r42 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 22 35 4.61231 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.252 $Y2=3.33
r44 22 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 21 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.19 $Y2=3.33
r46 21 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 19 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 19 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 19 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.19 $Y=2.2 $X2=2.19
+ $Y2=2.9
r51 13 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r52 13 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.9
r53 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.34 $Y=2.19 $X2=0.34
+ $Y2=2.9
r54 7 35 3.15387 $w=3.3e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.252 $Y2=3.33
r55 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.34 $Y2=2.9
r56 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=2.045 $X2=2.19 $Y2=2.9
r57 2 15 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=2.045 $X2=2.19 $Y2=2.2
r58 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=2.045 $X2=0.34 $Y2=2.9
r59 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=2.045 $X2=0.34 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_LP%X 1 2 9 15 17 18 19 20 26
r24 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.08 $Y=1.295
+ $X2=3.08 $Y2=1.665
r25 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.08 $Y=0.925
+ $X2=3.08 $Y2=1.295
r26 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.08 $Y=0.555
+ $X2=3.08 $Y2=0.925
r27 17 26 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.08 $Y=0.555
+ $X2=3.08 $Y2=0.445
r28 15 20 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.08 $Y=2.105
+ $X2=3.08 $Y2=1.665
r29 12 15 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.72 $Y=2.19
+ $X2=3.08 $Y2=2.19
r30 9 12 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=2.72 $Y=2.9 $X2=2.72
+ $Y2=2.275
r31 2 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=2.045 $X2=2.72 $Y2=2.19
r32 2 9 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=2.045 $X2=2.72 $Y2=2.9
r33 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_LP%A_27_57# 1 2 9 11 12 15
r29 13 15 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.22 $Y=0.825
+ $X2=1.22 $Y2=0.495
r30 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.055 $Y=0.91
+ $X2=1.22 $Y2=0.825
r31 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.055 $Y=0.91
+ $X2=0.445 $Y2=0.91
r32 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.825
+ $X2=0.445 $Y2=0.91
r33 7 9 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.28 $Y=0.825 $X2=0.28
+ $Y2=0.495
r34 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.285 $X2=1.22 $Y2=0.495
r35 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r45 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r46 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r48 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.29
+ $Y2=0
r50 27 29 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=3.12
+ $Y2=0
r51 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 23 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.75
+ $Y2=0
r54 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r55 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.29
+ $Y2=0
r56 22 25 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=1.2
+ $Y2=0
r57 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r58 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 17 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.75
+ $Y2=0
r60 17 19 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r61 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r62 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r63 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0
r64 11 13 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0.43
r65 7 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r66 7 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0.455
r67 2 13 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.235 $X2=2.29 $Y2=0.43
r68 1 9 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.285 $X2=0.71 $Y2=0.455
.ends

