* File: sky130_fd_sc_lp__einvp_2.pex.spice
* Created: Wed Sep  2 09:52:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVP_2%TE 3 8 9 11 13 15 17 18 20 22 23 24 26 32 33
r63 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=2.945
+ $X2=0.74 $Y2=2.945
r64 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=2.945 $X2=0.575 $Y2=2.945
r65 28 31 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=0.49 $Y=2.945
+ $X2=0.575 $Y2=2.945
r66 26 32 9.65171 $w=3.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=2.865
+ $X2=0.575 $Y2=2.865
r67 24 25 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.015 $Y=1.26
+ $X2=1.015 $Y2=1.41
r68 20 22 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.445 $Y=1.185
+ $X2=1.445 $Y2=0.655
r69 19 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.09 $Y=1.26
+ $X2=1.015 $Y2=1.26
r70 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.37 $Y=1.26
+ $X2=1.445 $Y2=1.185
r71 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.37 $Y=1.26
+ $X2=1.09 $Y2=1.26
r72 16 25 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.015 $Y=1.485
+ $X2=1.015 $Y2=1.41
r73 16 17 664.032 $w=1.5e-07 $l=1.295e-06 $layer=POLY_cond $X=1.015 $Y=1.485
+ $X2=1.015 $Y2=2.78
r74 13 24 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.015 $Y=1.185
+ $X2=1.015 $Y2=1.26
r75 13 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.015 $Y=1.185
+ $X2=1.015 $Y2=0.655
r76 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.94 $Y=2.855
+ $X2=1.015 $Y2=2.78
r77 11 33 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=0.94 $Y=2.855 $X2=0.74
+ $Y2=2.855
r78 10 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.565 $Y=1.41
+ $X2=0.49 $Y2=1.41
r79 9 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.94 $Y=1.41
+ $X2=1.015 $Y2=1.41
r80 9 10 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.94 $Y=1.41
+ $X2=0.565 $Y2=1.41
r81 6 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=2.78
+ $X2=0.49 $Y2=2.945
r82 6 8 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.49 $Y=2.78 $X2=0.49
+ $Y2=2.155
r83 5 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.49 $Y=1.485
+ $X2=0.49 $Y2=1.41
r84 5 8 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.49 $Y=1.485 $X2=0.49
+ $Y2=2.155
r85 1 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.49 $Y=1.335
+ $X2=0.49 $Y2=1.41
r86 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.49 $Y=1.335 $X2=0.49
+ $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_2%A_30_131# 1 2 7 9 10 12 15 19 23 24 26
c48 10 0 7.40582e-20 $X=2.015 $Y=1.725
r49 24 29 15.4929 $w=2.8e-07 $l=9e-08 $layer=POLY_cond $X=1.925 $Y=1.535
+ $X2=2.015 $Y2=1.535
r50 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.925
+ $Y=1.51 $X2=1.925 $Y2=1.51
r51 21 26 3.11956 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.4 $Y=1.51
+ $X2=0.255 $Y2=1.51
r52 21 23 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.4 $Y=1.51
+ $X2=1.925 $Y2=1.51
r53 17 26 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=1.595
+ $X2=0.255 $Y2=1.51
r54 17 19 15.2997 $w=2.88e-07 $l=3.85e-07 $layer=LI1_cond $X=0.255 $Y=1.595
+ $X2=0.255 $Y2=1.98
r55 13 26 3.40559 $w=2.75e-07 $l=9.21954e-08 $layer=LI1_cond $X=0.24 $Y=1.425
+ $X2=0.255 $Y2=1.51
r56 13 15 23.9354 $w=2.58e-07 $l=5.4e-07 $layer=LI1_cond $X=0.24 $Y=1.425
+ $X2=0.24 $Y2=0.885
r57 10 29 17.3521 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.015 $Y=1.725
+ $X2=2.015 $Y2=1.535
r58 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.015 $Y=1.725
+ $X2=2.015 $Y2=2.465
r59 7 24 58.5286 $w=2.8e-07 $l=4.245e-07 $layer=POLY_cond $X=1.585 $Y=1.725
+ $X2=1.925 $Y2=1.535
r60 7 9 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.585 $Y=1.725
+ $X2=1.585 $Y2=2.465
r61 2 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=1.98
r62 1 15 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.655 $X2=0.275 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_2%A 1 3 6 10 12 15 17 18 19 23 25
r42 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.46 $X2=3.09 $Y2=1.46
r43 22 25 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.875 $Y=1.46
+ $X2=3.09 $Y2=1.46
r44 22 23 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=1.46 $X2=2.8
+ $Y2=1.46
r45 19 26 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=3.125 $Y=1.665
+ $X2=3.125 $Y2=1.46
r46 18 26 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=1.295
+ $X2=3.125 $Y2=1.46
r47 13 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.625
+ $X2=2.875 $Y2=1.46
r48 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.875 $Y=1.625
+ $X2=2.875 $Y2=2.465
r49 10 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.295
+ $X2=2.875 $Y2=1.46
r50 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.875 $Y=1.295
+ $X2=2.875 $Y2=0.765
r51 9 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.52 $Y=1.37
+ $X2=2.445 $Y2=1.37
r52 9 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.52 $Y=1.37 $X2=2.8
+ $Y2=1.37
r53 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.445 $Y=1.445
+ $X2=2.445 $Y2=1.37
r54 4 6 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.445 $Y=1.445
+ $X2=2.445 $Y2=2.465
r55 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.445 $Y=1.295
+ $X2=2.445 $Y2=1.37
r56 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.445 $Y=1.295
+ $X2=2.445 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_2%VPWR 1 2 8 9 13 18 21 22 23 34 35 38
r57 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r60 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=1.8 $Y2=3.33
r62 29 31 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 23 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 23 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 23 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 21 26 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 21 22 5.53942 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=1.002 $Y2=3.33
r69 18 20 16.8252 $w=5.23e-07 $l=5.05e-07 $layer=LI1_cond $X=0.832 $Y=1.99
+ $X2=0.832 $Y2=2.495
r70 13 16 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.8 $Y=2.2 $X2=1.8
+ $Y2=2.97
r71 11 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.8 $Y=3.245 $X2=1.8
+ $Y2=3.33
r72 11 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.8 $Y=3.245
+ $X2=1.8 $Y2=2.97
r73 10 22 5.53942 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.002 $Y2=3.33
r74 9 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.635 $Y=3.33 $X2=1.8
+ $Y2=3.33
r75 9 10 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=1.095 $Y2=3.33
r76 8 22 1.03991 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.002 $Y=3.245
+ $X2=1.002 $Y2=3.33
r77 8 20 44.9631 $w=1.83e-07 $l=7.5e-07 $layer=LI1_cond $X=1.002 $Y=3.245
+ $X2=1.002 $Y2=2.495
r78 2 16 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=1.66
+ $Y=1.835 $X2=1.8 $Y2=2.97
r79 2 13 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.66
+ $Y=1.835 $X2=1.8 $Y2=2.2
r80 1 18 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_2%A_249_367# 1 2 3 12 16 17 19 22 24 26
r35 24 31 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=2.905
+ $X2=3.125 $Y2=2.99
r36 24 26 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=3.125 $Y=2.905
+ $X2=3.125 $Y2=2.085
r37 23 29 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.325 $Y=2.99
+ $X2=2.23 $Y2=2.99
r38 22 31 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.995 $Y=2.99
+ $X2=3.125 $Y2=2.99
r39 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.995 $Y=2.99
+ $X2=2.325 $Y2=2.99
r40 19 29 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.905
+ $X2=2.23 $Y2=2.99
r41 19 21 55.1627 $w=1.88e-07 $l=9.45e-07 $layer=LI1_cond $X=2.23 $Y=2.905
+ $X2=2.23 $Y2=1.96
r42 18 21 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=2.23 $Y=1.945
+ $X2=2.23 $Y2=1.96
r43 16 18 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.135 $Y=1.86
+ $X2=2.23 $Y2=1.945
r44 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.135 $Y=1.86
+ $X2=1.465 $Y2=1.86
r45 12 14 51.5727 $w=1.98e-07 $l=9.3e-07 $layer=LI1_cond $X=1.365 $Y=1.98
+ $X2=1.365 $Y2=2.91
r46 10 17 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.365 $Y=1.945
+ $X2=1.465 $Y2=1.86
r47 10 12 1.94091 $w=1.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.365 $Y=1.945
+ $X2=1.365 $Y2=1.98
r48 3 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.95
+ $Y=1.835 $X2=3.09 $Y2=2.91
r49 3 26 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=2.95
+ $Y=1.835 $X2=3.09 $Y2=2.085
r50 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.09
+ $Y=1.835 $X2=2.23 $Y2=2.91
r51 2 21 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.09
+ $Y=1.835 $X2=2.23 $Y2=1.96
r52 1 14 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.835 $X2=1.37 $Y2=2.91
r53 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.835 $X2=1.37 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_2%Z 1 2 7 8 9 10 11 18
c17 18 0 7.40582e-20 $X=2.66 $Y=0.68
r18 10 11 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.66 $Y=1.985
+ $X2=2.66 $Y2=2.405
r19 9 10 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.66 $Y=1.665
+ $X2=2.66 $Y2=1.985
r20 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=1.295 $X2=2.66
+ $Y2=1.665
r21 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=0.925 $X2=2.66
+ $Y2=1.295
r22 7 18 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.66 $Y=0.925
+ $X2=2.66 $Y2=0.68
r23 2 10 300 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=2 $X=2.52
+ $Y=1.835 $X2=2.66 $Y2=1.985
r24 1 18 91 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=2 $X=2.52
+ $Y=0.345 $X2=2.66 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_2%VGND 1 2 9 15 17 19 24 34 35 38 41
r40 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r43 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r44 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r45 29 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.66
+ $Y2=0
r46 29 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=2.16
+ $Y2=0
r47 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 25 38 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.732
+ $Y2=0
r50 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.2
+ $Y2=0
r51 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.66
+ $Y2=0
r52 24 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.2
+ $Y2=0
r53 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 19 38 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=0.732
+ $Y2=0
r56 19 21 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=0.24
+ $Y2=0
r57 17 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r58 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 17 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 13 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0
r61 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0.38
r62 9 11 16.4635 $w=3.83e-07 $l=5.5e-07 $layer=LI1_cond $X=0.732 $Y=0.38
+ $X2=0.732 $Y2=0.93
r63 7 38 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.732 $Y=0.085
+ $X2=0.732 $Y2=0
r64 7 9 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.732 $Y=0.085
+ $X2=0.732 $Y2=0.38
r65 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.52
+ $Y=0.235 $X2=1.66 $Y2=0.38
r66 1 11 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.655 $X2=0.705 $Y2=0.93
r67 1 9 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.655 $X2=0.8 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_2%A_218_47# 1 2 3 12 14 15 19 20 21 24
r36 22 24 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=3.125 $Y=0.425
+ $X2=3.125 $Y2=0.49
r37 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.995 $Y=0.34
+ $X2=3.125 $Y2=0.425
r38 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.995 $Y=0.34
+ $X2=2.325 $Y2=0.34
r39 17 19 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=2.195 $Y=1.065
+ $X2=2.195 $Y2=0.49
r40 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.195 $Y=0.425
+ $X2=2.325 $Y2=0.34
r41 16 19 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=2.195 $Y=0.425
+ $X2=2.195 $Y2=0.49
r42 14 17 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.065 $Y=1.15
+ $X2=2.195 $Y2=1.065
r43 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.065 $Y=1.15
+ $X2=1.325 $Y2=1.15
r44 10 15 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.21 $Y=1.065
+ $X2=1.325 $Y2=1.15
r45 10 12 32.3185 $w=2.28e-07 $l=6.45e-07 $layer=LI1_cond $X=1.21 $Y=1.065
+ $X2=1.21 $Y2=0.42
r46 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.95
+ $Y=0.345 $X2=3.09 $Y2=0.49
r47 2 19 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.105
+ $Y=0.345 $X2=2.23 $Y2=0.49
r48 1 12 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.42
.ends

