* File: sky130_fd_sc_lp__a41oi_lp.spice
* Created: Fri Aug 28 10:03:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41oi_lp.pex.spice"
.subckt sky130_fd_sc_lp__a41oi_lp  VNB VPB A4 A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* VPB	VPB
* VNB	VNB
MM1010 A_170_47# N_A4_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1001 A_248_47# N_A3_M1001_g A_170_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1009 A_326_47# N_A2_M1009_g A_248_47# VNB NSHORT L=0.15 W=0.42 AD=0.0756
+ AS=0.0504 PD=0.78 PS=0.66 NRD=35.712 NRS=18.564 M=1 R=2.8 SA=75001 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g A_326_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=35.712 M=1 R=2.8 SA=75001.5 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1005 A_514_47# N_B1_M1005_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.9 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_B1_M1006_g A_514_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.3 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A4_M1003_g N_A_27_409#_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1007 N_A_27_409#_M1007_d N_A3_M1007_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_27_409#_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.15 AS=0.14 PD=1.3 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1008 N_A_27_409#_M1008_d N_A1_M1008_g N_VPWR_M1002_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.15 PD=1.28 PS=1.3 NRD=0 NRS=3.9203 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_27_409#_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX11_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a41oi_lp.pxi.spice"
*
.ends
*
*
