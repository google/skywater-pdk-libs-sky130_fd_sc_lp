* File: sky130_fd_sc_lp__o21ai_0.pex.spice
* Created: Fri Aug 28 11:04:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21AI_0%A1 2 3 4 7 9 11 14 16 17 18 19 24 25
r43 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29 $Y=1.1
+ $X2=0.29 $Y2=1.1
r44 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=2.035
r45 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r46 17 25 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.1
r47 15 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.29 $Y=1.44
+ $X2=0.29 $Y2=1.1
r48 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.29 $Y=1.44
+ $X2=0.29 $Y2=1.605
r49 14 24 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.29 $Y=1.005
+ $X2=0.29 $Y2=1.1
r50 13 14 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.367 $Y=0.855
+ $X2=0.367 $Y2=1.005
r51 9 11 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.575 $Y=2.305
+ $X2=0.575 $Y2=2.735
r52 7 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.535 $Y=0.445
+ $X2=0.535 $Y2=0.855
r53 3 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.5 $Y=2.23
+ $X2=0.575 $Y2=2.305
r54 3 4 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=0.5 $Y=2.23 $X2=0.275
+ $Y2=2.23
r55 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.2 $Y=2.155
+ $X2=0.275 $Y2=2.23
r56 2 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.2 $Y=2.155 $X2=0.2
+ $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_0%A2 2 5 9 11 12 13 14 19
r46 19 21 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.855 $Y=1.41
+ $X2=0.855 $Y2=1.245
r47 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.835
+ $Y=1.41 $X2=0.835 $Y2=1.41
r48 13 14 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.772 $Y=1.665
+ $X2=0.772 $Y2=2.035
r49 13 20 9.9618 $w=2.93e-07 $l=2.55e-07 $layer=LI1_cond $X=0.772 $Y=1.665
+ $X2=0.772 $Y2=1.41
r50 12 20 4.49257 $w=2.93e-07 $l=1.15e-07 $layer=LI1_cond $X=0.772 $Y=1.295
+ $X2=0.772 $Y2=1.41
r51 9 11 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.965 $Y=2.735
+ $X2=0.965 $Y2=1.915
r52 5 21 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=0.965 $Y=0.445
+ $X2=0.965 $Y2=1.245
r53 2 11 49.8761 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=0.855 $Y=1.73
+ $X2=0.855 $Y2=1.915
r54 1 19 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=0.855 $Y=1.43 $X2=0.855
+ $Y2=1.41
r55 1 2 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=0.855 $Y=1.43 $X2=0.855
+ $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_0%B1 3 6 9 11 12 13 17 18
r32 17 19 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.51 $Y=1.635
+ $X2=1.51 $Y2=1.47
r33 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.535
+ $Y=1.635 $X2=1.535 $Y2=1.635
r34 12 13 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.642 $Y=1.665
+ $X2=1.642 $Y2=2.035
r35 12 18 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=1.642 $Y=1.665
+ $X2=1.642 $Y2=1.635
r36 9 11 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=1.395 $Y=2.735
+ $X2=1.395 $Y2=2.14
r37 6 11 48.9106 $w=3.8e-07 $l=1.9e-07 $layer=POLY_cond $X=1.51 $Y=1.95 $X2=1.51
+ $Y2=2.14
r38 5 17 3.65891 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.51 $Y=1.66 $X2=1.51
+ $Y2=1.635
r39 5 6 42.4433 $w=3.8e-07 $l=2.9e-07 $layer=POLY_cond $X=1.51 $Y=1.66 $X2=1.51
+ $Y2=1.95
r40 3 19 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=1.395 $Y=0.445
+ $X2=1.395 $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_0%VPWR 1 2 7 9 11 13 15 17 27
r26 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r30 18 23 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.262 $Y2=3.33
r31 18 20 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=1.2 $Y2=3.33
r32 17 26 4.14267 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.712 $Y2=3.33
r33 17 20 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.2 $Y2=3.33
r34 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r35 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 11 26 3.14202 $w=2.7e-07 $l=1.15521e-07 $layer=LI1_cond $X=1.64 $Y=3.245
+ $X2=1.712 $Y2=3.33
r37 11 13 29.2379 $w=2.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.64 $Y=3.245
+ $X2=1.64 $Y2=2.56
r38 7 23 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.262 $Y2=3.33
r39 7 9 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.36 $Y2=2.56
r40 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=2.415 $X2=1.61 $Y2=2.56
r41 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.235
+ $Y=2.415 $X2=0.36 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_0%Y 1 2 8 9 10 13 15 16 20 28
r37 20 28 2.90685 $w=3.2e-07 $l=7.5e-08 $layer=LI1_cond $X=1.175 $Y=2.48
+ $X2=1.175 $Y2=2.405
r38 15 28 0.20132 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=1.175 $Y=2.4 $X2=1.175
+ $Y2=2.405
r39 15 16 10.444 $w=3.18e-07 $l=2.9e-07 $layer=LI1_cond $X=1.175 $Y=2.485
+ $X2=1.175 $Y2=2.775
r40 15 20 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=1.175 $Y=2.485
+ $X2=1.175 $Y2=2.48
r41 11 13 27.2947 $w=2.83e-07 $l=6.75e-07 $layer=LI1_cond $X=1.632 $Y=1.12
+ $X2=1.632 $Y2=0.445
r42 9 11 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=1.49 $Y=1.205
+ $X2=1.632 $Y2=1.12
r43 9 10 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.49 $Y=1.205
+ $X2=1.27 $Y2=1.205
r44 8 15 7.16338 $w=3.03e-07 $l=1.249e-07 $layer=LI1_cond $X=1.185 $Y=2.28
+ $X2=1.175 $Y2=2.4
r45 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.185 $Y=1.29
+ $X2=1.27 $Y2=1.205
r46 7 8 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.185 $Y=1.29
+ $X2=1.185 $Y2=2.28
r47 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.415 $X2=1.18 $Y2=2.56
r48 1 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.47
+ $Y=0.235 $X2=1.61 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_0%A_39_47# 1 2 9 11 12 15
r30 13 15 11.2792 $w=2.33e-07 $l=2.3e-07 $layer=LI1_cond $X=1.202 $Y=0.675
+ $X2=1.202 $Y2=0.445
r31 11 13 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=1.085 $Y=0.76
+ $X2=1.202 $Y2=0.675
r32 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.085 $Y=0.76
+ $X2=0.415 $Y2=0.76
r33 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.285 $Y=0.675
+ $X2=0.415 $Y2=0.76
r34 7 9 10.1947 $w=2.58e-07 $l=2.3e-07 $layer=LI1_cond $X=0.285 $Y=0.675
+ $X2=0.285 $Y2=0.445
r35 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.235 $X2=1.18 $Y2=0.445
r36 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.195
+ $Y=0.235 $X2=0.32 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_0%VGND 1 6 8 10 17 18 21
r28 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r29 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r30 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r31 15 17 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.68
+ $Y2=0
r32 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r33 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r34 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r35 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r36 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r37 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r38 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0
r39 4 6 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.41
r40 1 6 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=0.61
+ $Y=0.235 $X2=0.75 $Y2=0.41
.ends

