* File: sky130_fd_sc_lp__dlrtn_4.pex.spice
* Created: Wed Sep  2 09:47:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRTN_4%D 2 5 9 10 11 12 13 18 20
r40 18 20 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.045
+ $X2=0.61 $Y2=0.88
r41 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.655
+ $Y=1.045 $X2=0.655 $Y2=1.045
r42 12 13 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.775 $Y=1.295
+ $X2=0.775 $Y2=1.665
r43 12 19 6.22958 $w=4.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.775 $Y=1.295
+ $X2=0.775 $Y2=1.045
r44 11 19 2.9902 $w=4.78e-07 $l=1.2e-07 $layer=LI1_cond $X=0.775 $Y=0.925
+ $X2=0.775 $Y2=1.045
r45 9 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.745 $Y=0.56
+ $X2=0.745 $Y2=0.88
r46 5 10 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.475 $Y=2.66
+ $X2=0.475 $Y2=1.55
r47 2 10 52.1105 $w=4.2e-07 $l=2.1e-07 $layer=POLY_cond $X=0.61 $Y=1.34 $X2=0.61
+ $Y2=1.55
r48 1 18 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=0.61 $Y=1.09 $X2=0.61
+ $Y2=1.045
r49 1 2 33.1044 $w=4.2e-07 $l=2.5e-07 $layer=POLY_cond $X=0.61 $Y=1.09 $X2=0.61
+ $Y2=1.34
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%GATE_N 3 7 9 13 15
r34 12 15 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.955 $Y=2.015
+ $X2=1.175 $Y2=2.015
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.955
+ $Y=2.015 $X2=0.955 $Y2=2.015
r36 9 13 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.955 $Y2=2.035
r37 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=2.18
+ $X2=1.175 $Y2=2.015
r38 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.175 $Y=2.18
+ $X2=1.175 $Y2=2.66
r39 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.85
+ $X2=1.175 $Y2=2.015
r40 1 3 661.468 $w=1.5e-07 $l=1.29e-06 $layer=POLY_cond $X=1.175 $Y=1.85
+ $X2=1.175 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%A_27_468# 1 2 9 13 17 18 20 23 26 27 28 30
+ 31 32 35 36 41 44
c110 31 0 9.02846e-20 $X=2.505 $Y=2.36
c111 13 0 2.83236e-20 $X=2.76 $Y=2.555
c112 9 0 3.16851e-19 $X=2.76 $Y=0.835
r113 38 41 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=0.23 $Y=0.5
+ $X2=0.51 $Y2=0.5
r114 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.67
+ $Y=1.57 $X2=2.67 $Y2=1.57
r115 33 35 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=2.67 $Y=2.275
+ $X2=2.67 $Y2=1.57
r116 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.505 $Y=2.36
+ $X2=2.67 $Y2=2.275
r117 31 32 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.505 $Y=2.36
+ $X2=2.01 $Y2=2.36
r118 29 32 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=1.842 $Y=2.445
+ $X2=2.01 $Y2=2.36
r119 29 30 13.2445 $w=3.33e-07 $l=3.85e-07 $layer=LI1_cond $X=1.842 $Y=2.445
+ $X2=1.842 $Y2=2.83
r120 27 30 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=1.675 $Y=2.915
+ $X2=1.842 $Y2=2.83
r121 27 28 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.675 $Y=2.915
+ $X2=1.125 $Y2=2.915
r122 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.04 $Y=2.83
+ $X2=1.125 $Y2=2.915
r123 25 26 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.04 $Y=2.49
+ $X2=1.04 $Y2=2.83
r124 24 44 3.05049 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.365 $Y=2.405
+ $X2=0.23 $Y2=2.405
r125 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.955 $Y=2.405
+ $X2=1.04 $Y2=2.49
r126 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.955 $Y=2.405
+ $X2=0.365 $Y2=2.405
r127 20 44 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=2.32
+ $X2=0.23 $Y2=2.405
r128 19 38 2.08978 $w=2.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.23 $Y=0.67
+ $X2=0.23 $Y2=0.5
r129 19 20 70.4271 $w=2.68e-07 $l=1.65e-06 $layer=LI1_cond $X=0.23 $Y=0.67
+ $X2=0.23 $Y2=2.32
r130 17 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.67 $Y=1.91
+ $X2=2.67 $Y2=1.57
r131 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.91
+ $X2=2.67 $Y2=2.075
r132 16 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.405
+ $X2=2.67 $Y2=1.57
r133 13 18 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.76 $Y=2.555
+ $X2=2.76 $Y2=2.075
r134 9 16 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.76 $Y=0.835
+ $X2=2.76 $Y2=1.405
r135 2 44 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.34 $X2=0.26 $Y2=2.485
r136 1 41 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.385
+ $Y=0.35 $X2=0.51 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%A_357_365# 1 2 9 13 14 20 23 24 25 27 28 30
+ 31 33 35 36 49
c114 35 0 1.5347e-19 $X=3.21 $Y=1.91
c115 31 0 1.65422e-19 $X=3.57 $Y=0.35
c116 28 0 1.46049e-19 $X=2.99 $Y=0.375
c117 23 0 7.94932e-20 $X=2.185 $Y=1.825
c118 14 0 2.83236e-20 $X=2.1 $Y=1.965
r119 36 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.91
+ $X2=3.21 $Y2=2.075
r120 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.21
+ $Y=1.91 $X2=3.21 $Y2=1.91
r121 33 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.21 $Y=1.14
+ $X2=2.905 $Y2=1.14
r122 33 35 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=3.21 $Y=1.225
+ $X2=3.21 $Y2=1.91
r123 31 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=0.35
+ $X2=3.57 $Y2=0.515
r124 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=0.35 $X2=3.57 $Y2=0.35
r125 28 30 27.8507 $w=2.38e-07 $l=5.8e-07 $layer=LI1_cond $X=2.99 $Y=0.375
+ $X2=3.57 $Y2=0.375
r126 27 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=1.055
+ $X2=2.905 $Y2=1.14
r127 26 28 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.905 $Y=0.495
+ $X2=2.99 $Y2=0.375
r128 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.905 $Y=0.495
+ $X2=2.905 $Y2=1.055
r129 25 40 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.27 $Y=1.14
+ $X2=2.185 $Y2=1.14
r130 24 41 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=1.14
+ $X2=2.905 $Y2=1.14
r131 24 25 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.82 $Y=1.14
+ $X2=2.27 $Y2=1.14
r132 22 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=1.225
+ $X2=2.185 $Y2=1.14
r133 22 23 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.185 $Y=1.225
+ $X2=2.185 $Y2=1.825
r134 18 40 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.005 $Y=1.14
+ $X2=2.185 $Y2=1.14
r135 18 20 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=2.005 $Y=1.055
+ $X2=2.005 $Y2=0.9
r136 14 23 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.1 $Y=1.965
+ $X2=2.185 $Y2=1.825
r137 14 16 7.82015 $w=2.78e-07 $l=1.9e-07 $layer=LI1_cond $X=2.1 $Y=1.965
+ $X2=1.91 $Y2=1.965
r138 13 49 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.55 $Y=0.835
+ $X2=3.55 $Y2=0.515
r139 9 46 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.12 $Y=2.555
+ $X2=3.12 $Y2=2.075
r140 2 16 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.785
+ $Y=1.825 $X2=1.91 $Y2=1.97
r141 1 20 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.625 $X2=2.005 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%A_250_70# 1 2 8 9 10 13 17 22 23 24 25 27 29
+ 30 31 35 39 43 46
c119 46 0 1.29453e-20 $X=1.4 $Y=1.525
c120 31 0 7.42903e-20 $X=2.22 $Y=1.49
c121 30 0 9.02846e-20 $X=2.145 $Y=1.49
c122 8 0 7.94932e-20 $X=1.665 $Y=1.325
r123 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.755
+ $Y=1.49 $X2=1.755 $Y2=1.49
r124 41 46 0.502427 $w=2.6e-07 $l=1.05e-07 $layer=LI1_cond $X=1.505 $Y=1.525
+ $X2=1.4 $Y2=1.525
r125 41 43 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=1.505 $Y=1.525
+ $X2=1.755 $Y2=1.525
r126 37 46 6.26566 $w=2.05e-07 $l=1.3e-07 $layer=LI1_cond $X=1.4 $Y=1.655
+ $X2=1.4 $Y2=1.525
r127 37 39 43.8355 $w=2.08e-07 $l=8.3e-07 $layer=LI1_cond $X=1.4 $Y=1.655
+ $X2=1.4 $Y2=2.485
r128 33 46 6.26566 $w=2.05e-07 $l=1.32476e-07 $layer=LI1_cond $X=1.395 $Y=1.395
+ $X2=1.4 $Y2=1.525
r129 33 35 49.9091 $w=1.98e-07 $l=9e-07 $layer=LI1_cond $X=1.395 $Y=1.395
+ $X2=1.395 $Y2=0.495
r130 30 44 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=2.145 $Y=1.49
+ $X2=1.755 $Y2=1.49
r131 30 31 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.145 $Y=1.49
+ $X2=2.22 $Y2=1.49
r132 29 44 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.74 $Y=1.49
+ $X2=1.755 $Y2=1.49
r133 25 32 71.3487 $w=1.52e-07 $l=2.26495e-07 $layer=POLY_cond $X=3.665 $Y=1.685
+ $X2=3.662 $Y2=1.46
r134 25 27 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.665 $Y=1.685
+ $X2=3.665 $Y2=2.445
r135 23 32 3.14937 $w=1.5e-07 $l=7.7e-08 $layer=POLY_cond $X=3.585 $Y=1.46
+ $X2=3.662 $Y2=1.46
r136 23 24 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.585 $Y=1.46
+ $X2=3.195 $Y2=1.46
r137 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.12 $Y=1.385
+ $X2=3.195 $Y2=1.46
r138 20 22 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.12 $Y=1.385
+ $X2=3.12 $Y2=0.835
r139 19 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.12 $Y=0.255
+ $X2=3.12 $Y2=0.835
r140 15 31 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.655
+ $X2=2.22 $Y2=1.49
r141 15 17 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.22 $Y=1.655
+ $X2=2.22 $Y2=2.555
r142 11 31 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.325
+ $X2=2.22 $Y2=1.49
r143 11 13 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.22 $Y=1.325
+ $X2=2.22 $Y2=0.835
r144 9 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.045 $Y=0.18
+ $X2=3.12 $Y2=0.255
r145 9 10 669.16 $w=1.5e-07 $l=1.305e-06 $layer=POLY_cond $X=3.045 $Y=0.18
+ $X2=1.74 $Y2=0.18
r146 8 29 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.665 $Y=1.325
+ $X2=1.74 $Y2=1.49
r147 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.665 $Y=0.255
+ $X2=1.74 $Y2=0.18
r148 7 8 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.665 $Y=0.255
+ $X2=1.665 $Y2=1.325
r149 2 39 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=2.34 $X2=1.39 $Y2=2.485
r150 1 35 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.25
+ $Y=0.35 $X2=1.39 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%A_789_99# 1 2 7 9 13 17 21 25 29 33 37 41 45
+ 48 49 52 55 56 59 63 64 65 68 70 76 81 82 91
c172 21 0 1.18362e-19 $X=5.905 $Y=0.655
c173 7 0 1.5347e-19 $X=4.02 $Y=1.175
r174 88 89 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.335 $Y=1.51
+ $X2=6.765 $Y2=1.51
r175 84 86 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.895 $Y=1.51
+ $X2=5.905 $Y2=1.51
r176 77 91 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=7.01 $Y=1.51
+ $X2=7.195 $Y2=1.51
r177 77 89 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=7.01 $Y=1.51
+ $X2=6.765 $Y2=1.51
r178 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.01
+ $Y=1.51 $X2=7.01 $Y2=1.51
r179 74 88 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=5.99 $Y=1.51
+ $X2=6.335 $Y2=1.51
r180 74 86 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.99 $Y=1.51
+ $X2=5.905 $Y2=1.51
r181 73 76 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=5.99 $Y=1.51
+ $X2=7.01 $Y2=1.51
r182 73 74 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.99
+ $Y=1.51 $X2=5.99 $Y2=1.51
r183 71 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.855 $Y=1.51
+ $X2=5.77 $Y2=1.51
r184 71 73 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.855 $Y=1.51
+ $X2=5.99 $Y2=1.51
r185 69 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.77 $Y=1.595
+ $X2=5.77 $Y2=1.51
r186 69 70 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=5.77 $Y=1.595
+ $X2=5.77 $Y2=2.3
r187 68 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.77 $Y=1.425
+ $X2=5.77 $Y2=1.51
r188 67 68 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.77 $Y=1.04
+ $X2=5.77 $Y2=1.425
r189 66 81 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=5.31 $Y=2.385
+ $X2=5.2 $Y2=2.385
r190 65 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.685 $Y=2.385
+ $X2=5.77 $Y2=2.3
r191 65 66 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.685 $Y=2.385
+ $X2=5.31 $Y2=2.385
r192 63 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.685 $Y=0.955
+ $X2=5.77 $Y2=1.04
r193 63 64 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.685 $Y=0.955
+ $X2=5.115 $Y2=0.955
r194 57 64 20.9205 $w=2.16e-07 $l=3.94816e-07 $layer=LI1_cond $X=4.755 $Y=0.882
+ $X2=5.115 $Y2=0.955
r195 57 59 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.755 $Y=0.725
+ $X2=4.755 $Y2=0.42
r196 55 81 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=5.09 $Y=2.385
+ $X2=5.2 $Y2=2.385
r197 55 56 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.09 $Y=2.385
+ $X2=4.28 $Y2=2.385
r198 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.115
+ $Y=1.57 $X2=4.115 $Y2=1.57
r199 50 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.115 $Y=2.3
+ $X2=4.28 $Y2=2.385
r200 50 52 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=4.115 $Y=2.3
+ $X2=4.115 $Y2=1.57
r201 48 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.115 $Y=1.91
+ $X2=4.115 $Y2=1.57
r202 48 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.115 $Y=1.91
+ $X2=4.115 $Y2=2.075
r203 43 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.195 $Y=1.675
+ $X2=7.195 $Y2=1.51
r204 43 45 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.195 $Y=1.675
+ $X2=7.195 $Y2=2.465
r205 39 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.195 $Y=1.345
+ $X2=7.195 $Y2=1.51
r206 39 41 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.195 $Y=1.345
+ $X2=7.195 $Y2=0.655
r207 35 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.765 $Y=1.675
+ $X2=6.765 $Y2=1.51
r208 35 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.765 $Y=1.675
+ $X2=6.765 $Y2=2.465
r209 31 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.765 $Y=1.345
+ $X2=6.765 $Y2=1.51
r210 31 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.765 $Y=1.345
+ $X2=6.765 $Y2=0.655
r211 27 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.675
+ $X2=6.335 $Y2=1.51
r212 27 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.335 $Y=1.675
+ $X2=6.335 $Y2=2.465
r213 23 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.345
+ $X2=6.335 $Y2=1.51
r214 23 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.335 $Y=1.345
+ $X2=6.335 $Y2=0.655
r215 19 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.905 $Y=1.345
+ $X2=5.905 $Y2=1.51
r216 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.905 $Y=1.345
+ $X2=5.905 $Y2=0.655
r217 15 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.895 $Y=1.675
+ $X2=5.895 $Y2=1.51
r218 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.895 $Y=1.675
+ $X2=5.895 $Y2=2.465
r219 13 49 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.025 $Y=2.445
+ $X2=4.025 $Y2=2.075
r220 7 53 79 $w=2.41e-07 $l=4.39943e-07 $layer=POLY_cond $X=4.02 $Y=1.175
+ $X2=4.115 $Y2=1.57
r221 7 9 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.02 $Y=1.175 $X2=4.02
+ $Y2=0.835
r222 2 81 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=5.045
+ $Y=1.835 $X2=5.185 $Y2=2.465
r223 1 59 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=4.63
+ $Y=0.235 $X2=4.755 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%A_639_125# 1 2 7 9 12 14 15 16 21 24 28 32
+ 33 35
c84 28 0 1.44123e-19 $X=4.69 $Y=1.35
c85 24 0 2.71061e-19 $X=4.525 $Y=1.15
c86 21 0 1.90545e-19 $X=3.635 $Y=1.065
c87 16 0 1.70802e-19 $X=3.545 $Y=0.775
r88 32 33 8.66191 $w=5.33e-07 $l=1.35e-07 $layer=LI1_cond $X=3.457 $Y=2.38
+ $X2=3.457 $Y2=2.245
r89 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.69
+ $Y=1.35 $X2=4.69 $Y2=1.35
r90 26 28 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.65 $Y=1.235
+ $X2=4.65 $Y2=1.35
r91 25 35 1.54918 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.725 $Y=1.15 $X2=3.635
+ $Y2=1.15
r92 24 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.525 $Y=1.15
+ $X2=4.65 $Y2=1.235
r93 24 25 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.525 $Y=1.15
+ $X2=3.725 $Y2=1.15
r94 22 35 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=1.235
+ $X2=3.635 $Y2=1.15
r95 22 33 62.2323 $w=1.78e-07 $l=1.01e-06 $layer=LI1_cond $X=3.635 $Y=1.235
+ $X2=3.635 $Y2=2.245
r96 21 35 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=1.065
+ $X2=3.635 $Y2=1.15
r97 20 21 11.0909 $w=1.78e-07 $l=1.8e-07 $layer=LI1_cond $X=3.635 $Y=0.885
+ $X2=3.635 $Y2=1.065
r98 16 20 6.90553 $w=2.2e-07 $l=1.48324e-07 $layer=LI1_cond $X=3.545 $Y=0.775
+ $X2=3.635 $Y2=0.885
r99 16 18 11.0006 $w=2.18e-07 $l=2.1e-07 $layer=LI1_cond $X=3.545 $Y=0.775
+ $X2=3.335 $Y2=0.775
r100 14 29 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.895 $Y=1.35
+ $X2=4.69 $Y2=1.35
r101 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.895 $Y=1.35
+ $X2=4.97 $Y2=1.35
r102 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.97 $Y=1.515
+ $X2=4.97 $Y2=1.35
r103 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.97 $Y=1.515
+ $X2=4.97 $Y2=2.465
r104 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.97 $Y=1.185
+ $X2=4.97 $Y2=1.35
r105 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.97 $Y=1.185
+ $X2=4.97 $Y2=0.655
r106 2 32 300 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=2 $X=3.195
+ $Y=2.235 $X2=3.4 $Y2=2.38
r107 1 18 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.625 $X2=3.335 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%RESET_B 3 7 9 10 11 16
c46 16 0 1.56858e-19 $X=5.42 $Y=1.375
c47 9 0 1.18362e-19 $X=5.04 $Y=1.295
c48 3 0 9.29041e-20 $X=5.33 $Y=0.655
r49 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.42 $Y=1.375
+ $X2=5.42 $Y2=1.54
r50 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.42 $Y=1.375
+ $X2=5.42 $Y2=1.21
r51 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.42
+ $Y=1.375 $X2=5.42 $Y2=1.375
r52 10 11 7.76402 $w=5.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.23 $Y=1.665
+ $X2=5.23 $Y2=2.035
r53 10 17 6.08531 $w=5.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.23 $Y=1.665
+ $X2=5.23 $Y2=1.375
r54 9 17 1.67871 $w=5.68e-07 $l=8e-08 $layer=LI1_cond $X=5.23 $Y=1.295 $X2=5.23
+ $Y2=1.375
r55 7 19 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=5.4 $Y=2.465 $X2=5.4
+ $Y2=1.54
r56 3 18 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.33 $Y=0.655
+ $X2=5.33 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%VPWR 1 2 3 4 5 6 21 25 29 31 35 39 43 45 49
+ 50 51 53 58 67 72 78 81 84 87 91
r106 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r107 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r108 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r109 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 76 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 76 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r113 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r114 73 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=3.33
+ $X2=6.55 $Y2=3.33
r115 73 75 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.715 $Y=3.33
+ $X2=6.96 $Y2=3.33
r116 72 90 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=7.245 $Y=3.33
+ $X2=7.462 $Y2=3.33
r117 72 75 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.245 $Y=3.33
+ $X2=6.96 $Y2=3.33
r118 71 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r119 71 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r120 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r121 68 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=3.33
+ $X2=5.645 $Y2=3.33
r122 68 70 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.81 $Y=3.33 $X2=6
+ $Y2=3.33
r123 67 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=3.33
+ $X2=6.55 $Y2=3.33
r124 67 70 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.385 $Y=3.33
+ $X2=6 $Y2=3.33
r125 66 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r126 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 63 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=3.33
+ $X2=2.49 $Y2=3.33
r128 63 65 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=2.655 $Y=3.33
+ $X2=4.56 $Y2=3.33
r129 62 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r130 62 79 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r132 59 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.66 $Y2=3.33
r133 59 61 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=2.16 $Y2=3.33
r134 58 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.49 $Y2=3.33
r135 58 61 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.16 $Y2=3.33
r136 56 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r137 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r138 53 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.66 $Y2=3.33
r139 53 55 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.24 $Y2=3.33
r140 51 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r141 51 82 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=2.64 $Y2=3.33
r142 49 65 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.59 $Y=3.33 $X2=4.56
+ $Y2=3.33
r143 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=3.33
+ $X2=4.755 $Y2=3.33
r144 45 48 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=7.41 $Y=2.19
+ $X2=7.41 $Y2=2.95
r145 43 90 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=7.41 $Y=3.245
+ $X2=7.462 $Y2=3.33
r146 43 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.41 $Y=3.245
+ $X2=7.41 $Y2=2.95
r147 39 42 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=6.55 $Y=2.19
+ $X2=6.55 $Y2=2.95
r148 37 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=3.245
+ $X2=6.55 $Y2=3.33
r149 37 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.55 $Y=3.245
+ $X2=6.55 $Y2=2.95
r150 33 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=3.33
r151 33 35 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=2.765
r152 32 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.92 $Y=3.33
+ $X2=4.755 $Y2=3.33
r153 31 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=5.645 $Y2=3.33
r154 31 32 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=4.92 $Y2=3.33
r155 27 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=3.245
+ $X2=4.755 $Y2=3.33
r156 27 29 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.755 $Y=3.245
+ $X2=4.755 $Y2=2.765
r157 23 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=3.245
+ $X2=2.49 $Y2=3.33
r158 23 25 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=2.49 $Y=3.245
+ $X2=2.49 $Y2=2.73
r159 19 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.66 $Y=3.245
+ $X2=0.66 $Y2=3.33
r160 19 21 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=0.66 $Y=3.245
+ $X2=0.66 $Y2=2.835
r161 6 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.27
+ $Y=1.835 $X2=7.41 $Y2=2.95
r162 6 45 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=7.27
+ $Y=1.835 $X2=7.41 $Y2=2.19
r163 5 42 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.41
+ $Y=1.835 $X2=6.55 $Y2=2.95
r164 5 39 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=6.41
+ $Y=1.835 $X2=6.55 $Y2=2.19
r165 4 35 600 $w=1.7e-07 $l=1.01143e-06 $layer=licon1_PDIFF $count=1 $X=5.475
+ $Y=1.835 $X2=5.645 $Y2=2.765
r166 3 29 600 $w=1.7e-07 $l=8.81008e-07 $layer=licon1_PDIFF $count=1 $X=4.1
+ $Y=2.235 $X2=4.755 $Y2=2.765
r167 2 25 600 $w=1.7e-07 $l=5.84423e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=2.235 $X2=2.49 $Y2=2.73
r168 1 21 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.34 $X2=0.69 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%Q 1 2 3 4 16 19 23 24 25 26 29 33 37 39 42
+ 45 46 48 51 53
c62 29 0 1.42181e-19 $X=6.98 $Y=0.42
c63 16 0 1.29923e-19 $X=6.12 $Y=0.93
r64 51 53 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=7.47 $Y=1.255 $X2=7.47
+ $Y2=1.295
r65 48 51 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.17 $X2=7.47
+ $Y2=1.255
r66 48 53 1.01415 $w=2.48e-07 $l=2.2e-08 $layer=LI1_cond $X=7.47 $Y=1.317
+ $X2=7.47 $Y2=1.295
r67 47 48 20.6518 $w=2.48e-07 $l=4.48e-07 $layer=LI1_cond $X=7.47 $Y=1.765
+ $X2=7.47 $Y2=1.317
r68 42 44 8.17035 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=0.42
+ $X2=6.085 $Y2=0.585
r69 40 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.075 $Y=1.85
+ $X2=6.98 $Y2=1.85
r70 39 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.345 $Y=1.85
+ $X2=7.47 $Y2=1.765
r71 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.345 $Y=1.85
+ $X2=7.075 $Y2=1.85
r72 38 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.075 $Y=1.17
+ $X2=6.98 $Y2=1.17
r73 37 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.345 $Y=1.17
+ $X2=7.47 $Y2=1.17
r74 37 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.345 $Y=1.17
+ $X2=7.075 $Y2=1.17
r75 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.98 $Y=1.98
+ $X2=6.98 $Y2=2.91
r76 31 46 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=1.935
+ $X2=6.98 $Y2=1.85
r77 31 33 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=6.98 $Y=1.935
+ $X2=6.98 $Y2=1.98
r78 27 45 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=1.085
+ $X2=6.98 $Y2=1.17
r79 27 29 38.8182 $w=1.88e-07 $l=6.65e-07 $layer=LI1_cond $X=6.98 $Y=1.085
+ $X2=6.98 $Y2=0.42
r80 25 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.885 $Y=1.85
+ $X2=6.98 $Y2=1.85
r81 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.885 $Y=1.85
+ $X2=6.215 $Y2=1.85
r82 23 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.885 $Y=1.17
+ $X2=6.98 $Y2=1.17
r83 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.885 $Y=1.17
+ $X2=6.215 $Y2=1.17
r84 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.12 $Y=1.98
+ $X2=6.12 $Y2=2.91
r85 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.12 $Y=1.935
+ $X2=6.215 $Y2=1.85
r86 17 19 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=6.12 $Y=1.935
+ $X2=6.12 $Y2=1.98
r87 16 44 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=6.12 $Y=0.93
+ $X2=6.12 $Y2=0.585
r88 14 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.12 $Y=1.085
+ $X2=6.215 $Y2=1.17
r89 14 16 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=6.12 $Y=1.085
+ $X2=6.12 $Y2=0.93
r90 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.835 $X2=6.98 $Y2=2.91
r91 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.835 $X2=6.98 $Y2=1.98
r92 3 21 400 $w=1.7e-07 $l=1.14755e-06 $layer=licon1_PDIFF $count=1 $X=5.97
+ $Y=1.835 $X2=6.12 $Y2=2.91
r93 3 19 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.97
+ $Y=1.835 $X2=6.12 $Y2=1.98
r94 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.84
+ $Y=0.235 $X2=6.98 $Y2=0.42
r95 1 42 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.98
+ $Y=0.235 $X2=6.12 $Y2=0.42
r96 1 16 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=5.98
+ $Y=0.235 $X2=6.12 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_4%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 47 48 49 61 65 70 75 81 84 87 91
r106 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r107 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r108 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r109 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r110 79 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r111 79 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r112 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r113 76 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=0 $X2=6.55
+ $Y2=0
r114 76 78 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.715 $Y=0 $X2=6.96
+ $Y2=0
r115 75 90 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=7.245 $Y=0
+ $X2=7.462 $Y2=0
r116 75 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.245 $Y=0
+ $X2=6.96 $Y2=0
r117 74 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r118 74 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r119 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r120 71 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=0 $X2=5.61
+ $Y2=0
r121 71 73 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.775 $Y=0 $X2=6
+ $Y2=0
r122 70 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=0 $X2=6.55
+ $Y2=0
r123 70 73 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.385 $Y=0 $X2=6
+ $Y2=0
r124 69 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r125 69 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r126 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r127 66 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=0 $X2=4.235
+ $Y2=0
r128 66 68 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.4 $Y=0 $X2=4.56
+ $Y2=0
r129 65 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.445 $Y=0 $X2=5.61
+ $Y2=0
r130 65 68 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=5.445 $Y=0 $X2=4.56
+ $Y2=0
r131 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r132 61 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.235
+ $Y2=0
r133 61 63 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=4.07 $Y=0 $X2=2.64
+ $Y2=0
r134 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r135 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r136 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r137 56 59 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r138 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r139 53 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r140 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r141 49 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r142 49 64 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=2.64
+ $Y2=0
r143 47 59 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.29 $Y=0 $X2=2.16
+ $Y2=0
r144 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=0 $X2=2.455
+ $Y2=0
r145 46 63 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.62 $Y=0 $X2=2.64
+ $Y2=0
r146 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=0 $X2=2.455
+ $Y2=0
r147 44 52 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.72
+ $Y2=0
r148 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.96
+ $Y2=0
r149 43 56 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.2
+ $Y2=0
r150 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=0.96
+ $Y2=0
r151 39 90 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.462 $Y2=0
r152 39 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0.38
r153 35 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=0.085
+ $X2=6.55 $Y2=0
r154 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.55 $Y=0.085
+ $X2=6.55 $Y2=0.38
r155 31 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.61 $Y=0.085
+ $X2=5.61 $Y2=0
r156 31 33 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.61 $Y=0.085
+ $X2=5.61 $Y2=0.58
r157 27 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.235 $Y=0.085
+ $X2=4.235 $Y2=0
r158 27 29 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=4.235 $Y=0.085
+ $X2=4.235 $Y2=0.79
r159 23 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=0.085
+ $X2=2.455 $Y2=0
r160 23 25 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.455 $Y=0.085
+ $X2=2.455 $Y2=0.77
r161 19 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=0.085
+ $X2=0.96 $Y2=0
r162 19 21 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.96 $Y=0.085
+ $X2=0.96 $Y2=0.495
r163 6 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.27
+ $Y=0.235 $X2=7.41 $Y2=0.38
r164 5 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.41
+ $Y=0.235 $X2=6.55 $Y2=0.38
r165 4 33 182 $w=1.7e-07 $l=4.35603e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.235 $X2=5.61 $Y2=0.58
r166 3 29 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.625 $X2=4.235 $Y2=0.79
r167 2 25 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.625 $X2=2.455 $Y2=0.77
r168 1 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.82
+ $Y=0.35 $X2=0.96 $Y2=0.495
.ends

