* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fa_lp A B CIN VGND VNB VPB VPWR COUT SUM
M1000 a_1049_419# B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.6e+11p pd=5.12e+06u as=2.64e+12p ps=1.528e+07u
M1001 SUM a_1574_141# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1002 a_355_141# CIN a_84_209# VNB nshort w=420000u l=150000u
+  ad=4.4395e+11p pd=4.02e+06u as=1.764e+11p ps=1.68e+06u
M1003 a_1049_419# A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND CIN a_1005_141# VNB nshort w=420000u l=150000u
+  ad=1.44145e+12p pd=1.129e+07u as=4.0825e+11p ps=3.85e+06u
M1005 VGND a_84_209# a_134_85# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_1956_66# a_1574_141# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 a_84_209# B a_577_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 a_1005_141# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1720_419# CIN a_1574_141# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=2.8e+11p ps=2.56e+06u
M1010 a_1574_141# a_84_209# a_1005_141# VNB nshort w=420000u l=150000u
+  ad=1.722e+11p pd=1.66e+06u as=0p ps=0u
M1011 a_84_209# B a_245_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.8e+11p pd=2.56e+06u as=7.45e+11p ps=5.49e+06u
M1012 a_1764_141# B a_1686_141# VNB nshort w=420000u l=150000u
+  ad=2.02125e+11p pd=2.24e+06u as=1.008e+11p ps=1.32e+06u
M1013 VGND A a_1764_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_84_209# COUT VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1015 VGND B a_355_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B a_458_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=6.65e+11p ps=5.33e+06u
M1017 VPWR A a_1818_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1018 a_134_85# a_84_209# COUT VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1019 VGND A a_355_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_577_141# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_458_409# A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1686_141# CIN a_1574_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1574_141# a_84_209# a_1049_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1005_141# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1818_419# B a_1720_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1026 SUM a_1574_141# a_1956_66# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1027 a_458_409# CIN a_84_209# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR CIN a_1049_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A a_245_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends
