* File: sky130_fd_sc_lp__o2111a_4.pex.spice
* Created: Fri Aug 28 11:00:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111A_4%D1 3 5 7 10 12 14 15 22
c42 12 0 5.72713e-20 $X=0.94 $Y=1.275
r43 22 23 1.47401 $w=3.27e-07 $l=1e-08 $layer=POLY_cond $X=0.93 $Y=1.44 $X2=0.94
+ $Y2=1.44
r44 21 22 61.9083 $w=3.27e-07 $l=4.2e-07 $layer=POLY_cond $X=0.51 $Y=1.44
+ $X2=0.93 $Y2=1.44
r45 20 21 1.47401 $w=3.27e-07 $l=1e-08 $layer=POLY_cond $X=0.5 $Y=1.44 $X2=0.51
+ $Y2=1.44
r46 18 20 31.6911 $w=3.27e-07 $l=2.15e-07 $layer=POLY_cond $X=0.285 $Y=1.44
+ $X2=0.5 $Y2=1.44
r47 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.285
+ $Y=1.44 $X2=0.285 $Y2=1.44
r48 15 19 5.47883 $w=3.03e-07 $l=1.45e-07 $layer=LI1_cond $X=0.237 $Y=1.295
+ $X2=0.237 $Y2=1.44
r49 12 23 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.275
+ $X2=0.94 $Y2=1.44
r50 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.94 $Y=1.275
+ $X2=0.94 $Y2=0.745
r51 8 22 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.605
+ $X2=0.93 $Y2=1.44
r52 8 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.93 $Y=1.605
+ $X2=0.93 $Y2=2.465
r53 5 21 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.275
+ $X2=0.51 $Y2=1.44
r54 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.51 $Y=1.275 $X2=0.51
+ $Y2=0.745
r55 1 20 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.605 $X2=0.5
+ $Y2=1.44
r56 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.5 $Y=1.605 $X2=0.5
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%C1 3 7 11 15 18 21 23 25 30 31 33
c97 30 0 1.58704e-19 $X=2.82 $Y=1.51
c98 18 0 1.86413e-19 $X=1.515 $Y=1.95
c99 7 0 1.76405e-19 $X=1.37 $Y=0.745
c100 3 0 1.59948e-19 $X=1.36 $Y=2.465
r101 31 42 46.2775 $w=4.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.867 $Y=1.51
+ $X2=2.867 $Y2=1.675
r102 31 41 46.2775 $w=4.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.867 $Y=1.51
+ $X2=2.867 $Y2=1.345
r103 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.51 $X2=2.82 $Y2=1.51
r104 27 33 13.0851 $w=3.48e-07 $l=3.55e-07 $layer=LI1_cond $X=2.645 $Y=1.595
+ $X2=2.645 $Y2=1.95
r105 26 30 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.645 $Y=1.51
+ $X2=2.82 $Y2=1.51
r106 26 27 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=1.51
+ $X2=2.645 $Y2=1.595
r107 25 33 33.8097 $w=3.38e-07 $l=9.55e-07 $layer=LI1_cond $X=1.6 $Y=2.035
+ $X2=2.555 $Y2=2.035
r108 21 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.51
+ $X2=1.39 $Y2=1.675
r109 21 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.51
+ $X2=1.39 $Y2=1.345
r110 20 23 6.54797 $w=2.18e-07 $l=1.25e-07 $layer=LI1_cond $X=1.39 $Y=1.535
+ $X2=1.515 $Y2=1.535
r111 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.39
+ $Y=1.51 $X2=1.39 $Y2=1.51
r112 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=1.95
+ $X2=1.6 $Y2=2.035
r113 17 23 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.515 $Y=1.645
+ $X2=1.515 $Y2=1.535
r114 17 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.515 $Y=1.645
+ $X2=1.515 $Y2=1.95
r115 15 42 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.73 $Y=2.465
+ $X2=2.73 $Y2=1.675
r116 11 41 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.73 $Y=0.745 $X2=2.73
+ $Y2=1.345
r117 7 38 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.37 $Y=0.745 $X2=1.37
+ $Y2=1.345
r118 3 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.36 $Y=2.465
+ $X2=1.36 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%B1 3 7 11 15 17 23 24
c51 3 0 4.22428e-20 $X=1.87 $Y=0.745
r52 22 24 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.08 $Y=1.51 $X2=2.3
+ $Y2=1.51
r53 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.51 $X2=2.08 $Y2=1.51
r54 19 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.87 $Y=1.51
+ $X2=2.08 $Y2=1.51
r55 17 23 3.06433 $w=6.03e-07 $l=1.55e-07 $layer=LI1_cond $X=2.072 $Y=1.665
+ $X2=2.072 $Y2=1.51
r56 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.675
+ $X2=2.3 $Y2=1.51
r57 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.3 $Y=1.675 $X2=2.3
+ $Y2=2.465
r58 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.345 $X2=2.3
+ $Y2=1.51
r59 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.3 $Y=1.345 $X2=2.3
+ $Y2=0.745
r60 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.675
+ $X2=1.87 $Y2=1.51
r61 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.87 $Y=1.675 $X2=1.87
+ $Y2=2.465
r62 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.345
+ $X2=1.87 $Y2=1.51
r63 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.87 $Y=1.345 $X2=1.87
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%A2 3 5 7 9 10 12 13 14 17 19 21 24 25 26 30
+ 40 42
c117 42 0 1.97215e-19 $X=3.6 $Y=1.295
c118 30 0 8.94706e-20 $X=3.61 $Y=1.26
c119 21 0 6.80566e-21 $X=5.33 $Y=1.16
c120 3 0 6.92333e-20 $X=3.63 $Y=2.465
r121 40 42 1.42277 $w=4.03e-07 $l=5e-08 $layer=LI1_cond $X=3.572 $Y=1.245
+ $X2=3.572 $Y2=1.295
r122 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.61 $Y=1.35
+ $X2=3.61 $Y2=1.515
r123 30 33 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.61 $Y=1.26 $X2=3.61
+ $Y2=1.35
r124 25 40 2.48344 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.572 $Y=1.16
+ $X2=3.572 $Y2=1.245
r125 25 26 10.0448 $w=4.03e-07 $l=3.53e-07 $layer=LI1_cond $X=3.572 $Y=1.312
+ $X2=3.572 $Y2=1.665
r126 25 42 0.483741 $w=4.03e-07 $l=1.7e-08 $layer=LI1_cond $X=3.572 $Y=1.312
+ $X2=3.572 $Y2=1.295
r127 25 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.61
+ $Y=1.35 $X2=3.61 $Y2=1.35
r128 24 38 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.33 $Y=1.49
+ $X2=5.33 $Y2=1.65
r129 24 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.33 $Y=1.49
+ $X2=5.33 $Y2=1.325
r130 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.33
+ $Y=1.49 $X2=5.33 $Y2=1.49
r131 21 23 16.0398 $w=2.51e-07 $l=3.3e-07 $layer=LI1_cond $X=5.33 $Y=1.16
+ $X2=5.33 $Y2=1.49
r132 20 25 5.93104 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=3.775 $Y=1.16
+ $X2=3.572 $Y2=1.16
r133 19 21 3.01842 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=1.16
+ $X2=5.33 $Y2=1.16
r134 19 20 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=5.165 $Y=1.16
+ $X2=3.775 $Y2=1.16
r135 17 37 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.31 $Y=0.655
+ $X2=5.31 $Y2=1.325
r136 13 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.165 $Y=1.65
+ $X2=5.33 $Y2=1.65
r137 13 14 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.165 $Y=1.65
+ $X2=4.995 $Y2=1.65
r138 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.92 $Y=1.725
+ $X2=4.995 $Y2=1.65
r139 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.92 $Y=1.725
+ $X2=4.92 $Y2=2.465
r140 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.02 $Y=1.185
+ $X2=4.02 $Y2=0.655
r141 6 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.775 $Y=1.26
+ $X2=3.61 $Y2=1.26
r142 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.945 $Y=1.26
+ $X2=4.02 $Y2=1.185
r143 5 6 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.945 $Y=1.26
+ $X2=3.775 $Y2=1.26
r144 3 35 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.63 $Y=2.465
+ $X2=3.63 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%A1 1 3 4 5 6 8 9 11 12 14 16 18 20 21 22 26
c68 26 0 1.97215e-19 $X=4.47 $Y=1.51
c69 20 0 6.80566e-21 $X=4.47 $Y=1.65
c70 18 0 1.19211e-19 $X=4.47 $Y=1.26
r71 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.47
+ $Y=1.51 $X2=4.47 $Y2=1.51
r72 22 27 3.00637 $w=3.43e-07 $l=9e-08 $layer=LI1_cond $X=4.56 $Y=1.587 $X2=4.47
+ $Y2=1.587
r73 21 27 13.0276 $w=3.43e-07 $l=3.9e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.47 $Y2=1.587
r74 19 26 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=4.47 $Y=1.575
+ $X2=4.47 $Y2=1.51
r75 19 20 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.47 $Y=1.575
+ $X2=4.47 $Y2=1.65
r76 17 26 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=4.47 $Y=1.335
+ $X2=4.47 $Y2=1.51
r77 17 18 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.47 $Y=1.335
+ $X2=4.47 $Y2=1.26
r78 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.88 $Y=1.185
+ $X2=4.88 $Y2=0.655
r79 13 18 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=1.26
+ $X2=4.47 $Y2=1.26
r80 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.805 $Y=1.26
+ $X2=4.88 $Y2=1.185
r81 12 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.805 $Y=1.26
+ $X2=4.635 $Y2=1.26
r82 9 20 13.5877 $w=2.4e-07 $l=8.44097e-08 $layer=POLY_cond $X=4.49 $Y=1.725
+ $X2=4.47 $Y2=1.65
r83 9 11 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.49 $Y=1.725
+ $X2=4.49 $Y2=2.465
r84 6 18 13.5877 $w=2.4e-07 $l=8.44097e-08 $layer=POLY_cond $X=4.45 $Y=1.185
+ $X2=4.47 $Y2=1.26
r85 6 8 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.45 $Y=1.185 $X2=4.45
+ $Y2=0.655
r86 4 20 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.65
+ $X2=4.47 $Y2=1.65
r87 4 5 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.305 $Y=1.65
+ $X2=4.135 $Y2=1.65
r88 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.06 $Y=1.725
+ $X2=4.135 $Y2=1.65
r89 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.06 $Y=1.725 $X2=4.06
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%A_32_367# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 51 53 55 59 65 67 71 73 75 79 81 84 85 90 97 101 105 108 124
c182 124 0 1.87664e-19 $X=7.185 $Y=1.49
c183 97 0 1.59948e-19 $X=1.145 $Y=1.98
r184 123 124 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.07 $Y=1.49
+ $X2=7.185 $Y2=1.49
r185 120 121 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=6.64 $Y=1.49
+ $X2=6.755 $Y2=1.49
r186 119 120 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=6.325 $Y=1.49
+ $X2=6.64 $Y2=1.49
r187 118 119 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=6.21 $Y=1.49
+ $X2=6.325 $Y2=1.49
r188 117 118 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=5.895 $Y=1.49
+ $X2=6.21 $Y2=1.49
r189 112 113 3.16711 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.135 $Y=2.015
+ $X2=5.135 $Y2=2.1
r190 111 112 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=5.135 $Y=1.98
+ $X2=5.135 $Y2=2.015
r191 108 111 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=5.135 $Y=1.84
+ $X2=5.135 $Y2=1.98
r192 105 107 9.55096 $w=6.77e-07 $l=5.3e-07 $layer=LI1_cond $X=3.197 $Y=2.38
+ $X2=3.197 $Y2=2.91
r193 104 105 5.13589 $w=6.77e-07 $l=2.85e-07 $layer=LI1_cond $X=3.197 $Y=2.095
+ $X2=3.197 $Y2=2.38
r194 102 104 1.44165 $w=6.77e-07 $l=8e-08 $layer=LI1_cond $X=3.197 $Y=2.015
+ $X2=3.197 $Y2=2.095
r195 91 123 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=6.89 $Y=1.49
+ $X2=7.07 $Y2=1.49
r196 91 121 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.89 $Y=1.49
+ $X2=6.755 $Y2=1.49
r197 90 91 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.89
+ $Y=1.49 $X2=6.89 $Y2=1.49
r198 88 117 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=5.87 $Y=1.49
+ $X2=5.895 $Y2=1.49
r199 88 114 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.87 $Y=1.49
+ $X2=5.78 $Y2=1.49
r200 87 90 62.8485 $w=1.78e-07 $l=1.02e-06 $layer=LI1_cond $X=5.87 $Y=1.495
+ $X2=6.89 $Y2=1.495
r201 87 88 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.87
+ $Y=1.49 $X2=5.87 $Y2=1.49
r202 85 87 1.5404 $w=1.78e-07 $l=2.5e-08 $layer=LI1_cond $X=5.845 $Y=1.495
+ $X2=5.87 $Y2=1.495
r203 83 85 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.76 $Y=1.585
+ $X2=5.845 $Y2=1.495
r204 83 84 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.76 $Y=1.585
+ $X2=5.76 $Y2=1.755
r205 82 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=1.84
+ $X2=5.135 $Y2=1.84
r206 81 84 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.675 $Y=1.84
+ $X2=5.76 $Y2=1.755
r207 81 82 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.675 $Y=1.84
+ $X2=5.3 $Y2=1.84
r208 79 113 14.1075 $w=2.88e-07 $l=3.55e-07 $layer=LI1_cond $X=5.155 $Y=2.455
+ $X2=5.155 $Y2=2.1
r209 76 102 9.10194 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=3.545 $Y=2.015
+ $X2=3.197 $Y2=2.015
r210 75 112 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.97 $Y=2.015
+ $X2=5.135 $Y2=2.015
r211 75 76 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=4.97 $Y=2.015
+ $X2=3.545 $Y2=2.015
r212 74 101 6.55305 $w=1.75e-07 $l=1.18e-07 $layer=LI1_cond $X=2.18 $Y=2.38
+ $X2=2.062 $Y2=2.38
r213 73 105 8.7286 $w=1.8e-07 $l=3.47e-07 $layer=LI1_cond $X=2.85 $Y=2.38
+ $X2=3.197 $Y2=2.38
r214 73 74 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.85 $Y=2.38
+ $X2=2.18 $Y2=2.38
r215 69 101 0.305871 $w=2.35e-07 $l=9e-08 $layer=LI1_cond $X=2.062 $Y=2.47
+ $X2=2.062 $Y2=2.38
r216 69 71 21.5777 $w=2.33e-07 $l=4.4e-07 $layer=LI1_cond $X=2.062 $Y=2.47
+ $X2=2.062 $Y2=2.91
r217 68 99 2.15711 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.275 $Y=2.375
+ $X2=1.162 $Y2=2.375
r218 67 101 6.55305 $w=1.75e-07 $l=1.19474e-07 $layer=LI1_cond $X=1.945 $Y=2.375
+ $X2=2.062 $Y2=2.38
r219 67 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.945 $Y=2.375
+ $X2=1.275 $Y2=2.375
r220 63 99 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=1.162 $Y=2.46
+ $X2=1.162 $Y2=2.375
r221 63 65 0.256098 $w=2.23e-07 $l=5e-09 $layer=LI1_cond $X=1.162 $Y=2.46
+ $X2=1.162 $Y2=2.465
r222 62 99 4.27425 $w=2.12e-07 $l=9.0802e-08 $layer=LI1_cond $X=1.15 $Y=2.29
+ $X2=1.162 $Y2=2.375
r223 62 97 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=1.15 $Y=2.29
+ $X2=1.15 $Y2=1.985
r224 57 97 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.725 $Y=1.9
+ $X2=1.145 $Y2=1.9
r225 57 59 39.6371 $w=3.28e-07 $l=1.135e-06 $layer=LI1_cond $X=0.725 $Y=1.815
+ $X2=0.725 $Y2=0.68
r226 56 94 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.38 $Y=1.9 $X2=0.25
+ $Y2=1.9
r227 55 57 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=1.9
+ $X2=0.725 $Y2=1.9
r228 55 56 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.56 $Y=1.9
+ $X2=0.38 $Y2=1.9
r229 51 94 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.25 $Y=1.985
+ $X2=0.25 $Y2=1.9
r230 51 53 41.0004 $w=2.58e-07 $l=9.25e-07 $layer=LI1_cond $X=0.25 $Y=1.985
+ $X2=0.25 $Y2=2.91
r231 47 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.185 $Y=1.655
+ $X2=7.185 $Y2=1.49
r232 47 49 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.185 $Y=1.655
+ $X2=7.185 $Y2=2.465
r233 43 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.07 $Y=1.325
+ $X2=7.07 $Y2=1.49
r234 43 45 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.07 $Y=1.325
+ $X2=7.07 $Y2=0.655
r235 39 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.755 $Y=1.655
+ $X2=6.755 $Y2=1.49
r236 39 41 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.755 $Y=1.655
+ $X2=6.755 $Y2=2.465
r237 35 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.64 $Y=1.325
+ $X2=6.64 $Y2=1.49
r238 35 37 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.64 $Y=1.325
+ $X2=6.64 $Y2=0.655
r239 31 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.325 $Y=1.655
+ $X2=6.325 $Y2=1.49
r240 31 33 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.325 $Y=1.655
+ $X2=6.325 $Y2=2.465
r241 27 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.21 $Y=1.325
+ $X2=6.21 $Y2=1.49
r242 27 29 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.21 $Y=1.325
+ $X2=6.21 $Y2=0.655
r243 23 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.895 $Y=1.655
+ $X2=5.895 $Y2=1.49
r244 23 25 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.895 $Y=1.655
+ $X2=5.895 $Y2=2.465
r245 19 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.78 $Y=1.325
+ $X2=5.78 $Y2=1.49
r246 19 21 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.78 $Y=1.325
+ $X2=5.78 $Y2=0.655
r247 6 111 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.995
+ $Y=1.835 $X2=5.135 $Y2=1.98
r248 6 79 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=4.995
+ $Y=1.835 $X2=5.135 $Y2=2.455
r249 5 107 200 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=3 $X=2.805
+ $Y=1.835 $X2=2.945 $Y2=2.91
r250 5 104 200 $w=1.7e-07 $l=3.40147e-07 $layer=licon1_PDIFF $count=3 $X=2.805
+ $Y=1.835 $X2=2.99 $Y2=2.095
r251 4 101 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.835 $X2=2.085 $Y2=2.375
r252 4 71 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.835 $X2=2.085 $Y2=2.91
r253 3 97 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.835 $X2=1.145 $Y2=1.98
r254 3 65 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=1.005
+ $Y=1.835 $X2=1.145 $Y2=2.465
r255 2 94 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=1.98
r256 2 53 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=2.91
r257 1 59 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.325 $X2=0.725 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%VPWR 1 2 3 4 5 6 7 24 30 34 38 42 48 52 54
+ 59 60 61 63 68 73 82 86 91 97 100 103 106 109 113
r121 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r122 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r124 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r125 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r126 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 95 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r128 95 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r129 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r130 92 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.54 $Y2=3.33
r131 92 94 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.96 $Y2=3.33
r132 91 112 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.235 $Y=3.33
+ $X2=7.457 $Y2=3.33
r133 91 94 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.235 $Y=3.33
+ $X2=6.96 $Y2=3.33
r134 90 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r135 90 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r136 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r137 87 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.68 $Y2=3.33
r138 87 89 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6 $Y2=3.33
r139 86 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=3.33
+ $X2=6.54 $Y2=3.33
r140 86 89 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.375 $Y=3.33
+ $X2=6 $Y2=3.33
r141 85 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r142 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 82 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.515 $Y=3.33
+ $X2=5.68 $Y2=3.33
r144 82 84 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=5.515 $Y=3.33
+ $X2=4.56 $Y2=3.33
r145 81 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r146 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r147 78 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=3.33
+ $X2=2.515 $Y2=3.33
r148 78 80 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.68 $Y=3.33
+ $X2=4.08 $Y2=3.33
r149 77 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r150 77 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r151 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r152 74 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=3.33
+ $X2=1.61 $Y2=3.33
r153 74 76 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.775 $Y=3.33
+ $X2=2.16 $Y2=3.33
r154 73 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.515 $Y2=3.33
r155 73 76 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.16 $Y2=3.33
r156 72 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r157 72 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r158 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r159 69 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=3.33
+ $X2=0.715 $Y2=3.33
r160 69 71 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=3.33 $X2=1.2
+ $Y2=3.33
r161 68 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.61 $Y2=3.33
r162 68 71 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r163 66 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r164 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r165 63 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.715 $Y2=3.33
r166 63 65 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.24 $Y2=3.33
r167 61 81 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r168 61 104 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=2.64 $Y2=3.33
r169 59 80 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.11 $Y=3.33 $X2=4.08
+ $Y2=3.33
r170 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.11 $Y=3.33
+ $X2=4.275 $Y2=3.33
r171 58 84 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.56 $Y2=3.33
r172 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.275 $Y2=3.33
r173 54 57 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=7.4 $Y=2.18 $X2=7.4
+ $Y2=2.95
r174 52 112 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.457 $Y2=3.33
r175 52 57 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.4 $Y2=2.95
r176 48 51 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.54 $Y=2.18
+ $X2=6.54 $Y2=2.95
r177 46 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.54 $Y=3.245
+ $X2=6.54 $Y2=3.33
r178 46 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.54 $Y=3.245
+ $X2=6.54 $Y2=2.95
r179 42 45 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.68 $Y=2.19
+ $X2=5.68 $Y2=2.95
r180 40 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=3.245
+ $X2=5.68 $Y2=3.33
r181 40 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.68 $Y=3.245
+ $X2=5.68 $Y2=2.95
r182 36 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.275 $Y=3.245
+ $X2=4.275 $Y2=3.33
r183 36 38 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.275 $Y=3.245
+ $X2=4.275 $Y2=2.745
r184 32 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=3.245
+ $X2=2.515 $Y2=3.33
r185 32 34 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.515 $Y=3.245
+ $X2=2.515 $Y2=2.775
r186 28 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=3.245
+ $X2=1.61 $Y2=3.33
r187 28 30 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=1.61 $Y=3.245
+ $X2=1.61 $Y2=2.745
r188 24 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.715 $Y=2.24
+ $X2=0.715 $Y2=2.95
r189 22 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=3.33
r190 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=2.95
r191 7 57 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.835 $X2=7.4 $Y2=2.95
r192 7 54 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.835 $X2=7.4 $Y2=2.18
r193 6 51 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.4
+ $Y=1.835 $X2=6.54 $Y2=2.95
r194 6 48 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=6.4
+ $Y=1.835 $X2=6.54 $Y2=2.18
r195 5 45 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=5.555
+ $Y=1.835 $X2=5.68 $Y2=2.95
r196 5 42 400 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_PDIFF $count=1 $X=5.555
+ $Y=1.835 $X2=5.68 $Y2=2.19
r197 4 38 600 $w=1.7e-07 $l=9.77497e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.835 $X2=4.275 $Y2=2.745
r198 3 34 600 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.835 $X2=2.515 $Y2=2.775
r199 2 30 600 $w=1.7e-07 $l=9.93655e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.835 $X2=1.61 $Y2=2.745
r200 1 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.715 $Y2=2.95
r201 1 24 400 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.715 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%A_741_367# 1 2 9 14 16
r15 10 14 3.98913 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.94 $Y=2.365
+ $X2=3.827 $Y2=2.365
r16 9 16 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.61 $Y=2.365
+ $X2=4.725 $Y2=2.365
r17 9 10 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.61 $Y=2.365
+ $X2=3.94 $Y2=2.365
r18 2 16 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=4.565
+ $Y=1.835 $X2=4.705 $Y2=2.445
r19 1 14 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=3.705
+ $Y=1.835 $X2=3.845 $Y2=2.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 42
+ 44 45 49 51
r60 49 51 1.92074 $w=3.58e-07 $l=6e-08 $layer=LI1_cond $X=7.415 $Y=1.235
+ $X2=7.415 $Y2=1.295
r61 44 49 2.57345 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=1.15
+ $X2=7.415 $Y2=1.235
r62 44 45 11.4604 $w=3.58e-07 $l=3.58e-07 $layer=LI1_cond $X=7.415 $Y=1.307
+ $X2=7.415 $Y2=1.665
r63 44 51 0.384148 $w=3.58e-07 $l=1.2e-08 $layer=LI1_cond $X=7.415 $Y=1.307
+ $X2=7.415 $Y2=1.295
r64 42 45 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=7.415 $Y=1.755
+ $X2=7.415 $Y2=1.665
r65 40 42 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.97 $Y=1.84
+ $X2=7.415 $Y2=1.84
r66 38 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.95 $Y=1.15
+ $X2=6.855 $Y2=1.15
r67 37 44 5.44966 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=7.235 $Y=1.15
+ $X2=7.415 $Y2=1.15
r68 37 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.235 $Y=1.15
+ $X2=6.95 $Y2=1.15
r69 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.97 $Y=1.98
+ $X2=6.97 $Y2=2.91
r70 31 40 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=1.925
+ $X2=6.97 $Y2=1.84
r71 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.97 $Y=1.925
+ $X2=6.97 $Y2=1.98
r72 27 39 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.855 $Y=1.065
+ $X2=6.855 $Y2=1.15
r73 27 29 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=6.855 $Y=1.065
+ $X2=6.855 $Y2=0.42
r74 25 40 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.875 $Y=1.84
+ $X2=6.97 $Y2=1.84
r75 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.875 $Y=1.84
+ $X2=6.205 $Y2=1.84
r76 23 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.76 $Y=1.15
+ $X2=6.855 $Y2=1.15
r77 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.76 $Y=1.15
+ $X2=6.09 $Y2=1.15
r78 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.11 $Y=1.98
+ $X2=6.11 $Y2=2.91
r79 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.11 $Y=1.925
+ $X2=6.205 $Y2=1.84
r80 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.11 $Y=1.925
+ $X2=6.11 $Y2=1.98
r81 13 24 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=5.977 $Y=1.065
+ $X2=6.09 $Y2=1.15
r82 13 15 33.0367 $w=2.23e-07 $l=6.45e-07 $layer=LI1_cond $X=5.977 $Y=1.065
+ $X2=5.977 $Y2=0.42
r83 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.83
+ $Y=1.835 $X2=6.97 $Y2=2.91
r84 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.83
+ $Y=1.835 $X2=6.97 $Y2=1.98
r85 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.97
+ $Y=1.835 $X2=6.11 $Y2=2.91
r86 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.97
+ $Y=1.835 $X2=6.11 $Y2=1.98
r87 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.715
+ $Y=0.235 $X2=6.855 $Y2=0.42
r88 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.855
+ $Y=0.235 $X2=5.995 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%A_32_65# 1 2 3 12 14 15 20 21 24
r49 22 24 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.015 $Y=1.085
+ $X2=3.015 $Y2=0.7
r50 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.85 $Y=1.17
+ $X2=3.015 $Y2=1.085
r51 20 21 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=2.85 $Y=1.17
+ $X2=1.25 $Y2=1.17
r52 17 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.155 $Y=1.085
+ $X2=1.25 $Y2=1.17
r53 17 19 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=1.155 $Y=1.085
+ $X2=1.155 $Y2=0.47
r54 16 19 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=1.155 $Y=0.425
+ $X2=1.155 $Y2=0.47
r55 14 16 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.06 $Y=0.34
+ $X2=1.155 $Y2=0.425
r56 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.06 $Y=0.34
+ $X2=0.39 $Y2=0.34
r57 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.26 $Y=0.425
+ $X2=0.39 $Y2=0.34
r58 10 12 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=0.26 $Y=0.425
+ $X2=0.26 $Y2=0.47
r59 3 24 91 $w=1.7e-07 $l=4.68375e-07 $layer=licon1_NDIFF $count=2 $X=2.805
+ $Y=0.325 $X2=3.015 $Y2=0.7
r60 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.325 $X2=1.155 $Y2=0.47
r61 1 12 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.325 $X2=0.295 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%A_289_65# 1 2 9 12 14 15
c22 9 0 5.72713e-20 $X=1.585 $Y=0.45
r23 14 15 7.3219 $w=2.33e-07 $l=1.4e-07 $layer=LI1_cond $X=2.515 $Y=0.797
+ $X2=2.375 $Y2=0.797
r24 12 15 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=1.75 $Y=0.82
+ $X2=2.375 $Y2=0.82
r25 7 12 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=1.585 $Y=0.725
+ $X2=1.75 $Y2=0.82
r26 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.585 $Y=0.725
+ $X2=1.585 $Y2=0.45
r27 2 14 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.325 $X2=2.515 $Y2=0.81
r28 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.445
+ $Y=0.325 $X2=1.585 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%A_389_65# 1 2 3 10 13 14 15 18 20 22 24 26
+ 32
c64 32 0 1.19211e-19 $X=4.235 $Y=0.82
c65 26 0 1.76405e-19 $X=2.085 $Y=0.34
c66 10 0 4.22428e-20 $X=3.35 $Y=0.34
r67 26 29 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.085 $Y=0.34
+ $X2=2.085 $Y2=0.45
r68 22 34 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.13 $Y=0.735
+ $X2=5.13 $Y2=0.82
r69 22 24 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=5.13 $Y=0.735
+ $X2=5.13 $Y2=0.42
r70 21 32 6.33349 $w=1.75e-07 $l=1.15473e-07 $layer=LI1_cond $X=4.33 $Y=0.82
+ $X2=4.217 $Y2=0.815
r71 20 34 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5 $Y=0.82 $X2=5.13
+ $Y2=0.82
r72 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5 $Y=0.82 $X2=4.33
+ $Y2=0.82
r73 16 32 0.455276 $w=2.25e-07 $l=9e-08 $layer=LI1_cond $X=4.217 $Y=0.725
+ $X2=4.217 $Y2=0.815
r74 16 18 15.622 $w=2.23e-07 $l=3.05e-07 $layer=LI1_cond $X=4.217 $Y=0.725
+ $X2=4.217 $Y2=0.42
r75 14 32 6.33349 $w=1.75e-07 $l=1.12e-07 $layer=LI1_cond $X=4.105 $Y=0.815
+ $X2=4.217 $Y2=0.815
r76 14 15 36.0455 $w=1.78e-07 $l=5.85e-07 $layer=LI1_cond $X=4.105 $Y=0.815
+ $X2=3.52 $Y2=0.815
r77 13 15 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.435 $Y=0.725
+ $X2=3.52 $Y2=0.815
r78 12 13 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.435 $Y=0.425
+ $X2=3.435 $Y2=0.725
r79 11 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=0.34
+ $X2=2.085 $Y2=0.34
r80 10 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.35 $Y=0.34
+ $X2=3.435 $Y2=0.425
r81 10 11 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=3.35 $Y=0.34
+ $X2=2.25 $Y2=0.34
r82 3 34 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.095 $Y2=0.82
r83 3 24 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.095 $Y2=0.42
r84 2 32 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.235 $X2=4.235 $Y2=0.82
r85 2 18 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.235 $X2=4.235 $Y2=0.42
r86 1 29 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.325 $X2=2.085 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_4%VGND 1 2 3 4 5 18 20 24 28 32 34 36 38 39
+ 40 49 54 59 65 68 71 75
c102 36 0 1.87664e-19 $X=7.285 $Y=0.36
r103 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r104 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r105 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r106 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r107 63 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r108 63 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r109 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r110 60 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.59 $Y=0 $X2=6.425
+ $Y2=0
r111 60 62 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.59 $Y=0 $X2=6.96
+ $Y2=0
r112 59 74 4.53027 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=7.12 $Y=0 $X2=7.4
+ $Y2=0
r113 59 62 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.12 $Y=0 $X2=6.96
+ $Y2=0
r114 58 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r115 58 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r116 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r117 55 68 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.695 $Y=0
+ $X2=5.562 $Y2=0
r118 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.695 $Y=0 $X2=6
+ $Y2=0
r119 54 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.26 $Y=0 $X2=6.425
+ $Y2=0
r120 54 57 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.26 $Y=0 $X2=6
+ $Y2=0
r121 53 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r122 53 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r123 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r124 50 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.665
+ $Y2=0
r125 50 52 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.04
+ $Y2=0
r126 49 68 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=5.43 $Y=0 $X2=5.562
+ $Y2=0
r127 49 52 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.43 $Y=0 $X2=5.04
+ $Y2=0
r128 47 48 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r129 44 48 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r130 43 47 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r131 43 44 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r132 40 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=4.56
+ $Y2=0
r133 40 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r134 38 47 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.69 $Y=0 $X2=3.6
+ $Y2=0
r135 38 39 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=3.812
+ $Y2=0
r136 34 74 3.23591 $w=3.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.285 $Y=0.085
+ $X2=7.4 $Y2=0
r137 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.285 $Y=0.085
+ $X2=7.285 $Y2=0.36
r138 30 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=0.085
+ $X2=6.425 $Y2=0
r139 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.425 $Y=0.085
+ $X2=6.425 $Y2=0.36
r140 26 68 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.562 $Y=0.085
+ $X2=5.562 $Y2=0
r141 26 28 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=5.562 $Y=0.085
+ $X2=5.562 $Y2=0.38
r142 22 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=0.085
+ $X2=4.665 $Y2=0
r143 22 24 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.665 $Y=0.085
+ $X2=4.665 $Y2=0.445
r144 21 39 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=3.935 $Y=0
+ $X2=3.812 $Y2=0
r145 20 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=4.665
+ $Y2=0
r146 20 21 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=3.935
+ $Y2=0
r147 16 39 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.812 $Y=0.085
+ $X2=3.812 $Y2=0
r148 16 18 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=3.812 $Y=0.085
+ $X2=3.812 $Y2=0.38
r149 5 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.145
+ $Y=0.235 $X2=7.285 $Y2=0.36
r150 4 32 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.285
+ $Y=0.235 $X2=6.425 $Y2=0.36
r151 3 28 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=5.385
+ $Y=0.235 $X2=5.545 $Y2=0.38
r152 2 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.235 $X2=4.665 $Y2=0.445
r153 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.68
+ $Y=0.235 $X2=3.805 $Y2=0.38
.ends

