* File: sky130_fd_sc_lp__nor4bb_m.spice
* Created: Wed Sep  2 10:12:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4bb_m.pex.spice"
.subckt sky130_fd_sc_lp__nor4bb_m  VNB VPB D_N B A C_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C_N	C_N
* A	A
* B	B
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_D_N_M1002_g N_A_27_507#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A_27_507#_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.7
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_284_99#_M1008_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.0588 PD=0.97 PS=0.7 NRD=9.996 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 N_Y_M1011_d N_B_M1011_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1155 PD=0.7 PS=0.97 NRD=0 NRS=67.14 M=1 R=2.8 SA=75001.8 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1011_d VNB NSHORT L=0.15 W=0.42 AD=0.0903
+ AS=0.0588 PD=0.85 PS=0.7 NRD=42.852 NRS=0 M=1 R=2.8 SA=75002.2 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_284_99#_M1005_d N_C_N_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0903 PD=1.37 PS=0.85 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_D_N_M1010_g N_A_27_507#_M1010_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_310_397# N_A_27_507#_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1006 A_382_397# N_A_284_99#_M1006_g A_310_397# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1009 A_454_397# N_B_M1009_g A_382_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.9
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g A_454_397# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.12915 AS=0.0441 PD=1.035 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1007 N_A_284_99#_M1007_d N_C_N_M1007_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.12915 PD=1.37 PS=1.035 NRD=0 NRS=157.127 M=1 R=2.8
+ SA=75002 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_80 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__nor4bb_m.pxi.spice"
*
.ends
*
*
