* File: sky130_fd_sc_lp__a32oi_1.pex.spice
* Created: Fri Aug 28 10:01:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32OI_1%B2 1 3 6 8 9 16
r26 13 16 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.425 $Y=1.46
+ $X2=0.63 $Y2=1.46
r27 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.425
+ $Y=1.46 $X2=0.425 $Y2=1.46
r28 9 14 6.65495 $w=3.53e-07 $l=2.05e-07 $layer=LI1_cond $X=0.332 $Y=1.665
+ $X2=0.332 $Y2=1.46
r29 8 14 5.35643 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.332 $Y=1.295
+ $X2=0.332 $Y2=1.46
r30 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.625
+ $X2=0.63 $Y2=1.46
r31 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.63 $Y=1.625 $X2=0.63
+ $Y2=2.465
r32 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.46
r33 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.63 $Y=1.295 $X2=0.63
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_1%B1 3 6 8 9 13 15
c34 6 0 1.02479e-19 $X=1.06 $Y=2.465
r35 13 16 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.46 $X2=1.1
+ $Y2=1.625
r36 13 15 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.46 $X2=1.1
+ $Y2=1.295
r37 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=1.46 $X2=1.105 $Y2=1.46
r38 9 14 6.84785 $w=3.43e-07 $l=2.05e-07 $layer=LI1_cond $X=1.192 $Y=1.665
+ $X2=1.192 $Y2=1.46
r39 8 14 5.51168 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.192 $Y=1.295
+ $X2=1.192 $Y2=1.46
r40 6 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.06 $Y=2.465
+ $X2=1.06 $Y2=1.625
r41 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.005 $Y=0.765
+ $X2=1.005 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_1%A1 3 6 8 9 10 11 17 19
c39 8 0 1.02479e-19 $X=1.68 $Y=0.555
r40 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.645 $Y=1.46
+ $X2=1.645 $Y2=1.625
r41 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.645 $Y=1.46
+ $X2=1.645 $Y2=1.295
r42 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.645
+ $Y=1.46 $X2=1.645 $Y2=1.46
r43 11 18 8.59094 $w=2.73e-07 $l=2.05e-07 $layer=LI1_cond $X=1.697 $Y=1.665
+ $X2=1.697 $Y2=1.46
r44 10 18 6.91466 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.697 $Y=1.295
+ $X2=1.697 $Y2=1.46
r45 9 10 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.697 $Y=0.925
+ $X2=1.697 $Y2=1.295
r46 8 9 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.697 $Y=0.555
+ $X2=1.697 $Y2=0.925
r47 6 20 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.555 $Y=2.465
+ $X2=1.555 $Y2=1.625
r48 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.555 $Y=0.765
+ $X2=1.555 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_1%A2 1 3 6 8 9 10 11 21
c39 8 0 1.11746e-19 $X=2.16 $Y=0.555
r40 19 21 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.185 $Y=1.46
+ $X2=2.325 $Y2=1.46
r41 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.185
+ $Y=1.46 $X2=2.185 $Y2=1.46
r42 16 19 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.095 $Y=1.46
+ $X2=2.185 $Y2=1.46
r43 11 20 6.84785 $w=3.43e-07 $l=2.05e-07 $layer=LI1_cond $X=2.177 $Y=1.665
+ $X2=2.177 $Y2=1.46
r44 10 20 5.51168 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.177 $Y=1.295
+ $X2=2.177 $Y2=1.46
r45 9 10 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.177 $Y=0.925
+ $X2=2.177 $Y2=1.295
r46 8 9 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.177 $Y=0.555
+ $X2=2.177 $Y2=0.925
r47 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.625
+ $X2=2.325 $Y2=1.46
r48 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.325 $Y=1.625
+ $X2=2.325 $Y2=2.465
r49 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.295
+ $X2=2.095 $Y2=1.46
r50 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.095 $Y=1.295
+ $X2=2.095 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_1%A3 3 6 8 10 17 19
c26 17 0 1.1209e-19 $X=2.775 $Y=1.46
c27 6 0 1.11746e-19 $X=2.755 $Y=2.465
r28 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.46
+ $X2=2.775 $Y2=1.625
r29 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.46
+ $X2=2.775 $Y2=1.295
r30 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.775
+ $Y=1.46 $X2=2.775 $Y2=1.46
r31 10 18 7.64161 $w=5.38e-07 $l=3.45e-07 $layer=LI1_cond $X=3.12 $Y=1.48
+ $X2=2.775 $Y2=1.48
r32 8 18 2.9902 $w=5.38e-07 $l=1.35e-07 $layer=LI1_cond $X=2.64 $Y=1.48
+ $X2=2.775 $Y2=1.48
r33 6 20 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.755 $Y=2.465
+ $X2=2.755 $Y2=1.625
r34 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.685 $Y=0.765
+ $X2=2.685 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_1%A_58_367# 1 2 3 10 12 14 16 18 22 26
c26 22 0 1.1209e-19 $X=2.54 $Y=2.085
r27 24 32 4.50329 $w=2e-07 $l=8.9861e-08 $layer=LI1_cond $X=2.54 $Y=2.46
+ $X2=2.53 $Y2=2.375
r28 24 26 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=2.54 $Y=2.46
+ $X2=2.54 $Y2=2.495
r29 20 32 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=2.29 $X2=2.53
+ $Y2=2.375
r30 20 22 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=2.53 $Y=2.29
+ $X2=2.53 $Y2=2.085
r31 19 31 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.435 $Y=2.375
+ $X2=1.307 $Y2=2.375
r32 18 32 1.93381 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.425 $Y=2.375
+ $X2=2.53 $Y2=2.375
r33 18 19 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=2.425 $Y=2.375
+ $X2=1.435 $Y2=2.375
r34 16 31 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.307 $Y=2.46
+ $X2=1.307 $Y2=2.375
r35 16 17 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=1.307 $Y=2.46
+ $X2=1.307 $Y2=2.905
r36 15 29 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.51 $Y=2.99 $X2=0.38
+ $Y2=2.99
r37 14 17 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.18 $Y=2.99
+ $X2=1.307 $Y2=2.905
r38 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.18 $Y=2.99
+ $X2=0.51 $Y2=2.99
r39 10 29 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.38 $Y=2.905
+ $X2=0.38 $Y2=2.99
r40 10 12 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=0.38 $Y=2.905
+ $X2=0.38 $Y2=2.085
r41 3 26 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=2.4
+ $Y=1.835 $X2=2.54 $Y2=2.495
r42 3 22 600 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.835 $X2=2.54 $Y2=2.085
r43 2 31 300 $w=1.7e-07 $l=7.04273e-07 $layer=licon1_PDIFF $count=2 $X=1.135
+ $Y=1.835 $X2=1.315 $Y2=2.455
r44 1 29 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.29
+ $Y=1.835 $X2=0.415 $Y2=2.91
r45 1 12 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.29
+ $Y=1.835 $X2=0.415 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_1%Y 1 2 8 11 12 15 19 20 21 22
r46 21 22 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.02
+ $X2=2.16 $Y2=2.02
r47 20 21 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.02 $X2=1.68
+ $Y2=2.02
r48 17 20 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=1.01 $Y=2.02 $X2=1.2
+ $Y2=2.02
r49 17 19 2.15711 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=2.02 $X2=0.845
+ $Y2=2.02
r50 13 15 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.245 $Y=0.86
+ $X2=1.245 $Y2=0.49
r51 11 13 7.31368 $w=1.8e-07 $l=1.84594e-07 $layer=LI1_cond $X=1.1 $Y=0.95
+ $X2=1.245 $Y2=0.86
r52 11 12 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=1.1 $Y=0.95 $X2=0.85
+ $Y2=0.95
r53 8 19 4.27425 $w=2.5e-07 $l=1.34164e-07 $layer=LI1_cond $X=0.765 $Y=1.92
+ $X2=0.845 $Y2=2.02
r54 7 12 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.765 $Y=1.04
+ $X2=0.85 $Y2=0.95
r55 7 8 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.765 $Y=1.04
+ $X2=0.765 $Y2=1.92
r56 2 19 300 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=2 $X=0.705
+ $Y=1.835 $X2=0.845 $Y2=2.035
r57 1 15 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.08
+ $Y=0.345 $X2=1.265 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_1%VPWR 1 2 7 9 13 15 20 26 36
r38 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 29 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 26 29 10.2649 $w=6.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.94 $Y=2.755
+ $X2=1.94 $Y2=3.33
r41 24 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 21 29 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=1.94 $Y2=3.33
r45 21 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 20 35 4.53846 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=3.082 $Y2=3.33
r47 20 23 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 15 29 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.605 $Y=3.33
+ $X2=1.94 $Y2=3.33
r50 15 17 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=1.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 13 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 13 18 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 13 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 9 12 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=2.97 $Y=2.01 $X2=2.97
+ $Y2=2.95
r55 7 35 3.22771 $w=3.3e-07 $l=1.4854e-07 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=3.082 $Y2=3.33
r56 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=2.95
r57 2 12 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.835 $X2=2.97 $Y2=2.95
r58 2 9 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.835 $X2=2.97 $Y2=2.01
r59 1 26 300 $w=1.7e-07 $l=1.1349e-06 $layer=licon1_PDIFF $count=2 $X=1.63
+ $Y=1.835 $X2=2.11 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_1%VGND 1 2 7 9 13 15 16 17 18 29
r34 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r36 26 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r37 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 23 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r39 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r40 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 20 31 3.95509 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.255
+ $Y2=0
r42 20 22 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.72
+ $Y2=0
r43 18 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r44 18 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r45 16 25 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.64
+ $Y2=0
r46 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.9
+ $Y2=0
r47 15 28 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=3.065 $Y=0 $X2=3.12
+ $Y2=0
r48 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=2.9
+ $Y2=0
r49 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=0.085 $X2=2.9
+ $Y2=0
r50 11 13 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=2.9 $Y=0.085
+ $X2=2.9 $Y2=0.49
r51 7 31 3.25713 $w=2.6e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.38 $Y=0.085
+ $X2=0.255 $Y2=0
r52 7 9 17.9515 $w=2.58e-07 $l=4.05e-07 $layer=LI1_cond $X=0.38 $Y=0.085
+ $X2=0.38 $Y2=0.49
r53 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.76
+ $Y=0.345 $X2=2.9 $Y2=0.49
r54 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.29
+ $Y=0.345 $X2=0.415 $Y2=0.49
.ends

