* File: sky130_fd_sc_lp__xnor2_1.pxi.spice
* Created: Fri Aug 28 11:34:58 2020
* 
x_PM_SKY130_FD_SC_LP__XNOR2_1%B N_B_M1004_g N_B_M1002_g N_B_M1000_g N_B_M1001_g
+ N_B_c_77_p N_B_c_71_n N_B_c_64_n N_B_c_65_n B B N_B_c_67_n N_B_c_68_n
+ PM_SKY130_FD_SC_LP__XNOR2_1%B
x_PM_SKY130_FD_SC_LP__XNOR2_1%A N_A_c_143_n N_A_M1007_g N_A_M1006_g N_A_c_144_n
+ N_A_M1009_g N_A_M1008_g N_A_c_145_n N_A_c_146_n N_A_c_147_n A A N_A_c_148_n
+ PM_SKY130_FD_SC_LP__XNOR2_1%A
x_PM_SKY130_FD_SC_LP__XNOR2_1%A_33_47# N_A_33_47#_M1004_s N_A_33_47#_M1002_d
+ N_A_33_47#_M1003_g N_A_33_47#_M1005_g N_A_33_47#_c_205_n N_A_33_47#_c_217_n
+ N_A_33_47#_c_219_n N_A_33_47#_c_206_n N_A_33_47#_c_207_n N_A_33_47#_c_227_n
+ N_A_33_47#_c_230_n N_A_33_47#_c_208_n N_A_33_47#_c_211_n N_A_33_47#_c_237_n
+ N_A_33_47#_c_209_n PM_SKY130_FD_SC_LP__XNOR2_1%A_33_47#
x_PM_SKY130_FD_SC_LP__XNOR2_1%VPWR N_VPWR_M1002_s N_VPWR_M1006_d N_VPWR_M1005_d
+ N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_297_n VPWR
+ N_VPWR_c_298_n N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_293_n VPWR
+ PM_SKY130_FD_SC_LP__XNOR2_1%VPWR
x_PM_SKY130_FD_SC_LP__XNOR2_1%Y N_Y_M1003_d N_Y_M1001_d N_Y_c_352_n N_Y_c_364_n
+ N_Y_c_354_n N_Y_c_343_n Y Y Y Y N_Y_c_344_n N_Y_c_347_n Y N_Y_c_345_n
+ PM_SKY130_FD_SC_LP__XNOR2_1%Y
x_PM_SKY130_FD_SC_LP__XNOR2_1%VGND N_VGND_M1007_d N_VGND_M1009_d N_VGND_c_378_n
+ N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n VGND N_VGND_c_382_n
+ N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n VGND
+ PM_SKY130_FD_SC_LP__XNOR2_1%VGND
x_PM_SKY130_FD_SC_LP__XNOR2_1%A_302_47# N_A_302_47#_M1009_s N_A_302_47#_M1000_d
+ N_A_302_47#_c_425_n N_A_302_47#_c_428_n N_A_302_47#_c_426_n
+ N_A_302_47#_c_436_n N_A_302_47#_c_440_n PM_SKY130_FD_SC_LP__XNOR2_1%A_302_47#
cc_1 VNB N_B_M1002_g 0.00843998f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_2 VNB N_B_M1000_g 0.0258974f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.655
cc_3 VNB N_B_c_64_n 0.00349564f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.51
cc_4 VNB N_B_c_65_n 0.0223855f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.51
cc_5 VNB B 0.0221204f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_B_c_67_n 0.0423263f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.35
cc_7 VNB N_B_c_68_n 0.0219524f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.185
cc_8 VNB N_A_c_143_n 0.0187051f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.185
cc_9 VNB N_A_c_144_n 0.0208843f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=1.345
cc_10 VNB N_A_c_145_n 0.0179297f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=2.005
cc_11 VNB N_A_c_146_n 0.0557674f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=2.005
cc_12 VNB N_A_c_147_n 0.0145743f $X=-0.19 $Y=-0.245 $X2=0.262 $Y2=1.92
cc_13 VNB N_A_c_148_n 0.0028508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_33_47#_M1003_g 0.0281005f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.655
cc_15 VNB N_A_33_47#_c_205_n 0.0227027f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=2.005
cc_16 VNB N_A_33_47#_c_206_n 0.0295692f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A_33_47#_c_207_n 0.0109276f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_A_33_47#_c_208_n 0.00449354f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.35
cc_19 VNB N_A_33_47#_c_209_n 0.0273863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_293_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_343_n 0.00745412f $X=-0.19 $Y=-0.245 $X2=0.262 $Y2=1.92
cc_22 VNB N_Y_c_344_n 0.0303447f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.185
cc_23 VNB N_Y_c_345_n 0.0225054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_378_n 0.00928581f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.655
cc_25 VNB N_VGND_c_379_n 0.0055721f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=2.465
cc_26 VNB N_VGND_c_380_n 0.0283014f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=2.005
cc_27 VNB N_VGND_c_381_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=2.005
cc_28 VNB N_VGND_c_382_n 0.018068f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_VGND_c_383_n 0.0294937f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.185
cc_30 VNB N_VGND_c_384_n 0.197645f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_31 VNB N_VGND_c_385_n 0.00631724f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.675
cc_32 VNB N_A_302_47#_c_425_n 0.00465065f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.655
cc_33 VNB N_A_302_47#_c_426_n 0.00178967f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=1.675
cc_34 VPB N_B_M1002_g 0.0247181f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_35 VPB N_B_M1001_g 0.0193441f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.465
cc_36 VPB N_B_c_71_n 0.00942129f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=2.005
cc_37 VPB N_B_c_64_n 0.00127155f $X=-0.19 $Y=1.655 $X2=2.3 $Y2=1.51
cc_38 VPB N_B_c_65_n 0.00622484f $X=-0.19 $Y=1.655 $X2=2.3 $Y2=1.51
cc_39 VPB B 0.0110219f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_40 VPB N_A_M1006_g 0.0238138f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_41 VPB N_A_M1008_g 0.0237863f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.465
cc_42 VPB N_A_c_145_n 0.00266858f $X=-0.19 $Y=1.655 $X2=1.825 $Y2=2.005
cc_43 VPB N_A_c_146_n 0.0182643f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=2.005
cc_44 VPB N_A_c_147_n 5.21411e-19 $X=-0.19 $Y=1.655 $X2=0.262 $Y2=1.92
cc_45 VPB N_A_c_148_n 0.00910704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_33_47#_M1005_g 0.0213198f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.465
cc_47 VPB N_A_33_47#_c_211_n 0.00103837f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.185
cc_48 VPB N_A_33_47#_c_209_n 0.00674542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_294_n 0.0111601f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=0.655
cc_50 VPB N_VPWR_c_295_n 0.036146f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=1.675
cc_51 VPB N_VPWR_c_296_n 0.0103403f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.465
cc_52 VPB N_VPWR_c_297_n 0.0172906f $X=-0.19 $Y=1.655 $X2=1.825 $Y2=2.005
cc_53 VPB N_VPWR_c_298_n 0.0307321f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_299_n 0.0154255f $X=-0.19 $Y=1.655 $X2=0.262 $Y2=1.295
cc_55 VPB N_VPWR_c_300_n 0.0162327f $X=-0.19 $Y=1.655 $X2=0.262 $Y2=1.665
cc_56 VPB N_VPWR_c_293_n 0.0446846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB Y 0.00494099f $X=-0.19 $Y=1.655 $X2=2.3 $Y2=1.51
cc_58 VPB N_Y_c_347_n 0.00905019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB Y 0.0143669f $X=-0.19 $Y=1.655 $X2=0.262 $Y2=1.665
cc_60 VPB N_Y_c_345_n 0.00887046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 N_B_c_68_n N_A_c_143_n 0.0524063f $X=0.385 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_62 N_B_M1002_g N_A_M1006_g 0.0350083f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_63 N_B_c_77_p N_A_M1006_g 0.0124865f $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_64 B N_A_M1006_g 8.62061e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_B_M1000_g N_A_c_144_n 0.0322384f $X=2.39 $Y=0.655 $X2=0 $Y2=0
cc_66 N_B_M1001_g N_A_M1008_g 0.0446796f $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_67 N_B_c_77_p N_A_M1008_g 0.00690275f $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_68 N_B_c_64_n N_A_M1008_g 0.0171373f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_69 N_B_c_77_p N_A_c_145_n 2.92856e-19 $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_70 B N_A_c_145_n 0.00120753f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 N_B_c_67_n N_A_c_145_n 0.0320257f $X=0.355 $Y=1.35 $X2=0 $Y2=0
cc_72 N_B_c_77_p N_A_c_146_n 0.00398658f $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_73 N_B_c_64_n N_A_c_147_n 0.00968613f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_74 N_B_c_65_n N_A_c_147_n 0.0226036f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_75 N_B_c_77_p N_A_c_148_n 0.0742199f $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_76 N_B_c_64_n N_A_c_148_n 0.0275076f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_77 B N_A_c_148_n 0.024655f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_B_c_67_n N_A_c_148_n 0.00260468f $X=0.355 $Y=1.35 $X2=0 $Y2=0
cc_79 N_B_c_77_p N_A_33_47#_M1002_d 0.00350685f $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_80 N_B_M1000_g N_A_33_47#_M1003_g 0.0284187f $X=2.39 $Y=0.655 $X2=0 $Y2=0
cc_81 N_B_M1001_g N_A_33_47#_M1005_g 0.0364649f $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_82 N_B_c_68_n N_A_33_47#_c_205_n 0.0114925f $X=0.385 $Y=1.185 $X2=0 $Y2=0
cc_83 N_B_M1002_g N_A_33_47#_c_217_n 0.00216614f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_84 N_B_c_77_p N_A_33_47#_c_217_n 0.0153678f $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_85 N_B_M1002_g N_A_33_47#_c_219_n 0.00869234f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_86 N_B_M1000_g N_A_33_47#_c_206_n 0.0113142f $X=2.39 $Y=0.655 $X2=0 $Y2=0
cc_87 N_B_c_77_p N_A_33_47#_c_206_n 0.00318133f $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_88 N_B_c_64_n N_A_33_47#_c_206_n 0.0496995f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_89 N_B_c_65_n N_A_33_47#_c_206_n 0.00443399f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_90 B N_A_33_47#_c_207_n 0.0311053f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B_c_67_n N_A_33_47#_c_207_n 0.0017268f $X=0.355 $Y=1.35 $X2=0 $Y2=0
cc_92 N_B_c_68_n N_A_33_47#_c_207_n 0.0174528f $X=0.385 $Y=1.185 $X2=0 $Y2=0
cc_93 N_B_M1001_g N_A_33_47#_c_227_n 2.45189e-19 $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_94 N_B_c_77_p N_A_33_47#_c_227_n 0.0607726f $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_95 N_B_c_64_n N_A_33_47#_c_227_n 0.0155362f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_96 N_B_M1001_g N_A_33_47#_c_230_n 0.0124023f $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_97 N_B_c_64_n N_A_33_47#_c_230_n 0.00951562f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_98 N_B_M1000_g N_A_33_47#_c_208_n 0.00183209f $X=2.39 $Y=0.655 $X2=0 $Y2=0
cc_99 N_B_c_64_n N_A_33_47#_c_208_n 0.0164964f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_100 N_B_c_65_n N_A_33_47#_c_208_n 8.92009e-19 $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_101 N_B_M1001_g N_A_33_47#_c_211_n 0.00402332f $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_102 N_B_c_64_n N_A_33_47#_c_211_n 0.0114396f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_103 N_B_M1001_g N_A_33_47#_c_237_n 0.00977301f $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_104 N_B_c_64_n N_A_33_47#_c_237_n 0.015311f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B_c_65_n N_A_33_47#_c_237_n 6.40793e-19 $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_106 N_B_c_64_n N_A_33_47#_c_209_n 3.13661e-19 $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_107 N_B_c_65_n N_A_33_47#_c_209_n 0.0212538f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_108 N_B_c_71_n N_VPWR_M1002_s 0.00310159f $X=0.44 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_109 B N_VPWR_M1002_s 3.95201e-19 $X=0.155 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_110 N_B_c_77_p N_VPWR_M1006_d 0.0169813f $X=1.825 $Y=2.005 $X2=0 $Y2=0
cc_111 N_B_M1002_g N_VPWR_c_295_n 0.00579872f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_112 N_B_c_71_n N_VPWR_c_295_n 0.0224079f $X=0.44 $Y=2.005 $X2=0 $Y2=0
cc_113 N_B_M1001_g N_VPWR_c_297_n 0.00112063f $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_114 N_B_M1001_g N_VPWR_c_298_n 0.00585385f $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_115 N_B_M1002_g N_VPWR_c_299_n 0.0054895f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B_M1002_g N_VPWR_c_300_n 6.82747e-19 $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B_M1001_g N_VPWR_c_300_n 0.00335725f $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_118 N_B_M1002_g N_VPWR_c_293_n 0.0107508f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B_M1001_g N_VPWR_c_293_n 0.0114566f $X=2.39 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B_c_64_n A_385_367# 0.00714446f $X=2.3 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_121 N_B_c_68_n N_VGND_c_378_n 0.00293265f $X=0.385 $Y=1.185 $X2=0 $Y2=0
cc_122 N_B_M1000_g N_VGND_c_379_n 0.00346025f $X=2.39 $Y=0.655 $X2=0 $Y2=0
cc_123 N_B_c_68_n N_VGND_c_380_n 0.00549284f $X=0.385 $Y=1.185 $X2=0 $Y2=0
cc_124 N_B_M1000_g N_VGND_c_383_n 0.00440547f $X=2.39 $Y=0.655 $X2=0 $Y2=0
cc_125 N_B_M1000_g N_VGND_c_384_n 0.00654212f $X=2.39 $Y=0.655 $X2=0 $Y2=0
cc_126 N_B_c_68_n N_VGND_c_384_n 0.00716953f $X=0.385 $Y=1.185 $X2=0 $Y2=0
cc_127 N_B_M1000_g N_A_302_47#_c_425_n 6.72946e-19 $X=2.39 $Y=0.655 $X2=0 $Y2=0
cc_128 N_B_M1000_g N_A_302_47#_c_428_n 0.0131412f $X=2.39 $Y=0.655 $X2=0 $Y2=0
cc_129 N_A_c_143_n N_A_33_47#_c_205_n 0.0016502f $X=0.9 $Y=1.185 $X2=0 $Y2=0
cc_130 N_A_c_143_n N_A_33_47#_c_206_n 0.0104312f $X=0.9 $Y=1.185 $X2=0 $Y2=0
cc_131 N_A_c_144_n N_A_33_47#_c_206_n 0.00727111f $X=1.85 $Y=1.185 $X2=0 $Y2=0
cc_132 N_A_c_145_n N_A_33_47#_c_206_n 0.00544694f $X=0.9 $Y=1.43 $X2=0 $Y2=0
cc_133 N_A_c_146_n N_A_33_47#_c_206_n 0.0271397f $X=1.775 $Y=1.43 $X2=0 $Y2=0
cc_134 N_A_c_147_n N_A_33_47#_c_206_n 0.00484188f $X=1.85 $Y=1.43 $X2=0 $Y2=0
cc_135 N_A_c_148_n N_A_33_47#_c_206_n 0.062379f $X=1.49 $Y=1.51 $X2=0 $Y2=0
cc_136 N_A_c_143_n N_A_33_47#_c_207_n 0.00109753f $X=0.9 $Y=1.185 $X2=0 $Y2=0
cc_137 N_A_c_148_n N_A_33_47#_c_207_n 0.0123174f $X=1.49 $Y=1.51 $X2=0 $Y2=0
cc_138 N_A_M1006_g N_A_33_47#_c_227_n 0.0142704f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_M1008_g N_A_33_47#_c_227_n 0.0155369f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A_M1008_g N_A_33_47#_c_237_n 0.00380756f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_M1008_g N_VPWR_c_298_n 0.00388479f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_M1006_g N_VPWR_c_299_n 0.00486043f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_M1006_g N_VPWR_c_300_n 0.0151507f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_M1008_g N_VPWR_c_300_n 0.0235783f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1006_g N_VPWR_c_293_n 0.00822376f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_M1008_g N_VPWR_c_293_n 0.00704974f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_c_143_n N_VGND_c_378_n 0.0183425f $X=0.9 $Y=1.185 $X2=0 $Y2=0
cc_148 N_A_c_144_n N_VGND_c_378_n 0.00346595f $X=1.85 $Y=1.185 $X2=0 $Y2=0
cc_149 N_A_c_146_n N_VGND_c_378_n 0.00131022f $X=1.775 $Y=1.43 $X2=0 $Y2=0
cc_150 N_A_c_144_n N_VGND_c_379_n 0.00506054f $X=1.85 $Y=1.185 $X2=0 $Y2=0
cc_151 N_A_c_143_n N_VGND_c_380_n 0.00486043f $X=0.9 $Y=1.185 $X2=0 $Y2=0
cc_152 N_A_c_144_n N_VGND_c_382_n 0.00428252f $X=1.85 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A_c_143_n N_VGND_c_384_n 0.00828783f $X=0.9 $Y=1.185 $X2=0 $Y2=0
cc_154 N_A_c_144_n N_VGND_c_384_n 0.00751064f $X=1.85 $Y=1.185 $X2=0 $Y2=0
cc_155 N_A_c_143_n N_A_302_47#_c_425_n 9.01218e-19 $X=0.9 $Y=1.185 $X2=0 $Y2=0
cc_156 N_A_c_144_n N_A_302_47#_c_425_n 0.00806553f $X=1.85 $Y=1.185 $X2=0 $Y2=0
cc_157 N_A_c_144_n N_A_302_47#_c_428_n 0.00938814f $X=1.85 $Y=1.185 $X2=0 $Y2=0
cc_158 N_A_c_144_n N_A_302_47#_c_426_n 7.17169e-19 $X=1.85 $Y=1.185 $X2=0 $Y2=0
cc_159 N_A_c_146_n N_A_302_47#_c_426_n 0.00130701f $X=1.775 $Y=1.43 $X2=0 $Y2=0
cc_160 N_A_33_47#_c_227_n N_VPWR_M1006_d 0.0170845f $X=2.165 $Y=2.345 $X2=0
+ $Y2=0
cc_161 N_A_33_47#_M1005_g N_VPWR_c_297_n 0.0111902f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_33_47#_M1005_g N_VPWR_c_298_n 0.00486043f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_33_47#_c_219_n N_VPWR_c_299_n 0.015688f $X=0.72 $Y=2.91 $X2=0 $Y2=0
cc_164 N_A_33_47#_c_227_n N_VPWR_c_300_n 0.0583344f $X=2.165 $Y=2.345 $X2=0
+ $Y2=0
cc_165 N_A_33_47#_M1002_d N_VPWR_c_293_n 0.00380103f $X=0.58 $Y=1.835 $X2=0
+ $Y2=0
cc_166 N_A_33_47#_M1005_g N_VPWR_c_293_n 0.00458005f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_33_47#_c_219_n N_VPWR_c_293_n 0.00984745f $X=0.72 $Y=2.91 $X2=0 $Y2=0
cc_168 N_A_33_47#_c_227_n A_385_367# 0.0105198f $X=2.165 $Y=2.345 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_33_47#_c_237_n A_385_367# 0.00790073f $X=2.25 $Y=2.1 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A_33_47#_c_230_n N_Y_M1001_d 0.00826753f $X=2.675 $Y=2.1 $X2=0 $Y2=0
cc_171 N_A_33_47#_c_211_n N_Y_M1001_d 0.00210879f $X=2.76 $Y=2.015 $X2=0 $Y2=0
cc_172 N_A_33_47#_c_230_n N_Y_c_352_n 0.0194873f $X=2.675 $Y=2.1 $X2=0 $Y2=0
cc_173 N_A_33_47#_c_209_n N_Y_c_352_n 2.458e-19 $X=2.84 $Y=1.51 $X2=0 $Y2=0
cc_174 N_A_33_47#_M1005_g N_Y_c_354_n 0.015592f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A_33_47#_c_230_n N_Y_c_354_n 0.00266139f $X=2.675 $Y=2.1 $X2=0 $Y2=0
cc_176 N_A_33_47#_M1003_g N_Y_c_343_n 0.00468351f $X=2.885 $Y=0.655 $X2=0 $Y2=0
cc_177 N_A_33_47#_c_208_n N_Y_c_343_n 0.00741808f $X=2.76 $Y=1.675 $X2=0 $Y2=0
cc_178 N_A_33_47#_M1003_g N_Y_c_345_n 0.00353612f $X=2.885 $Y=0.655 $X2=0 $Y2=0
cc_179 N_A_33_47#_M1005_g N_Y_c_345_n 0.00353817f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_33_47#_c_208_n N_Y_c_345_n 0.0341285f $X=2.76 $Y=1.675 $X2=0 $Y2=0
cc_181 N_A_33_47#_c_211_n N_Y_c_345_n 0.0090955f $X=2.76 $Y=2.015 $X2=0 $Y2=0
cc_182 N_A_33_47#_c_209_n N_Y_c_345_n 0.00814023f $X=2.84 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A_33_47#_c_207_n A_116_47# 0.00296772f $X=0.78 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_33_47#_c_205_n N_VGND_c_378_n 0.0181973f $X=0.29 $Y=0.38 $X2=0 $Y2=0
cc_185 N_A_33_47#_c_206_n N_VGND_c_378_n 0.0244341f $X=2.675 $Y=1.17 $X2=0 $Y2=0
cc_186 N_A_33_47#_c_205_n N_VGND_c_380_n 0.0197852f $X=0.29 $Y=0.38 $X2=0 $Y2=0
cc_187 N_A_33_47#_M1003_g N_VGND_c_383_n 0.0054895f $X=2.885 $Y=0.655 $X2=0
+ $Y2=0
cc_188 N_A_33_47#_M1004_s N_VGND_c_384_n 0.00215406f $X=0.165 $Y=0.235 $X2=0
+ $Y2=0
cc_189 N_A_33_47#_M1003_g N_VGND_c_384_n 0.0110197f $X=2.885 $Y=0.655 $X2=0
+ $Y2=0
cc_190 N_A_33_47#_c_205_n N_VGND_c_384_n 0.012508f $X=0.29 $Y=0.38 $X2=0 $Y2=0
cc_191 N_A_33_47#_c_207_n N_VGND_c_384_n 0.0107989f $X=0.78 $Y=1.17 $X2=0 $Y2=0
cc_192 N_A_33_47#_c_206_n N_A_302_47#_c_428_n 0.0448188f $X=2.675 $Y=1.17 $X2=0
+ $Y2=0
cc_193 N_A_33_47#_c_206_n N_A_302_47#_c_426_n 0.0245409f $X=2.675 $Y=1.17 $X2=0
+ $Y2=0
cc_194 N_A_33_47#_M1003_g N_A_302_47#_c_436_n 0.00219412f $X=2.885 $Y=0.655
+ $X2=0 $Y2=0
cc_195 N_A_33_47#_c_206_n N_A_302_47#_c_436_n 0.0132261f $X=2.675 $Y=1.17 $X2=0
+ $Y2=0
cc_196 N_A_33_47#_c_208_n N_A_302_47#_c_436_n 0.0118949f $X=2.76 $Y=1.675 $X2=0
+ $Y2=0
cc_197 N_A_33_47#_c_209_n N_A_302_47#_c_436_n 4.92304e-19 $X=2.84 $Y=1.51 $X2=0
+ $Y2=0
cc_198 N_A_33_47#_M1003_g N_A_302_47#_c_440_n 0.00625231f $X=2.885 $Y=0.655
+ $X2=0 $Y2=0
cc_199 N_VPWR_c_293_n A_385_367# 0.016774f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_200 N_VPWR_c_293_n N_Y_M1001_d 0.00443357f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_298_n N_Y_c_364_n 0.0172687f $X=2.935 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_c_293_n N_Y_c_364_n 0.0100457f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_203 N_VPWR_c_297_n N_Y_c_354_n 0.00175662f $X=3.1 $Y=2.85 $X2=0 $Y2=0
cc_204 N_VPWR_c_293_n N_Y_c_354_n 0.00561519f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_M1005_d Y 0.00295493f $X=2.96 $Y=1.835 $X2=0 $Y2=0
cc_206 N_VPWR_M1005_d N_Y_c_347_n 0.00318869f $X=2.96 $Y=1.835 $X2=0 $Y2=0
cc_207 N_VPWR_c_297_n N_Y_c_347_n 0.0217628f $X=3.1 $Y=2.85 $X2=0 $Y2=0
cc_208 N_VPWR_c_293_n N_Y_c_347_n 0.00143554f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_209 N_VPWR_M1005_d Y 0.00305146f $X=2.96 $Y=1.835 $X2=0 $Y2=0
cc_210 N_Y_c_344_n N_VGND_c_383_n 0.0181731f $X=3.1 $Y=0.42 $X2=0 $Y2=0
cc_211 N_Y_M1003_d N_VGND_c_384_n 0.0040649f $X=2.96 $Y=0.235 $X2=0 $Y2=0
cc_212 N_Y_c_344_n N_VGND_c_384_n 0.0100252f $X=3.1 $Y=0.42 $X2=0 $Y2=0
cc_213 A_116_47# N_VGND_c_384_n 0.00487419f $X=0.58 $Y=0.235 $X2=0.29 $Y2=1.015
cc_214 N_VGND_c_384_n N_A_302_47#_M1009_s 0.00215158f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_215 N_VGND_c_384_n N_A_302_47#_M1000_d 0.00296667f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_378_n N_A_302_47#_c_425_n 0.0376927f $X=1.115 $Y=0.38 $X2=0
+ $Y2=0
cc_217 N_VGND_c_382_n N_A_302_47#_c_425_n 0.0210049f $X=1.97 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_384_n N_A_302_47#_c_425_n 0.0125589f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_M1009_d N_A_302_47#_c_428_n 0.005915f $X=1.925 $Y=0.235 $X2=0
+ $Y2=0
cc_220 N_VGND_c_379_n N_A_302_47#_c_428_n 0.0216986f $X=2.135 $Y=0.455 $X2=0
+ $Y2=0
cc_221 N_VGND_c_382_n N_A_302_47#_c_428_n 0.00191958f $X=1.97 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_383_n N_A_302_47#_c_428_n 0.00231886f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_384_n N_A_302_47#_c_428_n 0.00966551f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_224 N_VGND_c_378_n N_A_302_47#_c_426_n 0.0139f $X=1.115 $Y=0.38 $X2=0 $Y2=0
cc_225 N_VGND_c_383_n N_A_302_47#_c_440_n 0.0203968f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_226 N_VGND_c_384_n N_A_302_47#_c_440_n 0.0125589f $X=3.12 $Y=0 $X2=0 $Y2=0
