* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21bo_0 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VGND B1_N a_216_526# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR A2 a_467_458# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_467_458# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 VPWR B1_N a_216_526# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 X a_72_212# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_533_52# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_216_526# a_72_212# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_72_212# A1 a_533_52# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_72_212# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_72_212# a_216_526# a_467_458# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
