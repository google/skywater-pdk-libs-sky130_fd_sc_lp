* File: sky130_fd_sc_lp__o21bai_1.pex.spice
* Created: Wed Sep  2 10:17:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BAI_1%B1_N 3 5 6 7 9 12 13 14 18
c38 18 0 5.38984e-20 $X=0.385 $Y=1.35
r39 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.35 $X2=0.385 $Y2=1.35
r40 14 19 8.44232 $w=4.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.3 $Y=1.665
+ $X2=0.3 $Y2=1.35
r41 13 19 1.47406 $w=4.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.3 $Y=1.295 $X2=0.3
+ $Y2=1.35
r42 12 18 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=0.385 $Y=1.755
+ $X2=0.385 $Y2=1.35
r43 11 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.185
+ $X2=0.385 $Y2=1.35
r44 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.95 $Y=1.905 $X2=0.95
+ $Y2=2.225
r45 6 12 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.55 $Y=1.83
+ $X2=0.385 $Y2=1.755
r46 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.875 $Y=1.83
+ $X2=0.95 $Y2=1.905
r47 5 6 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.875 $Y=1.83
+ $X2=0.55 $Y2=1.83
r48 3 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.475 $Y=0.555
+ $X2=0.475 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_1%A_27_69# 1 2 7 9 12 14 15 18 20 21 23 27 28
+ 34
r64 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.955
+ $Y=1.35 $X2=0.955 $Y2=1.35
r65 32 34 5.51776 $w=3.28e-07 $l=1.58e-07 $layer=LI1_cond $X=0.797 $Y=1.35
+ $X2=0.955 $Y2=1.35
r66 30 32 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.792 $Y=1.35
+ $X2=0.797 $Y2=1.35
r67 27 28 7.16023 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=2.225
+ $X2=0.735 $Y2=2.06
r68 24 30 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=0.792 $Y=1.515
+ $X2=0.792 $Y2=1.35
r69 24 28 29.2131 $w=2.13e-07 $l=5.45e-07 $layer=LI1_cond $X=0.792 $Y=1.515
+ $X2=0.792 $Y2=2.06
r70 23 32 2.99809 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=0.797 $Y=1.185
+ $X2=0.797 $Y2=1.35
r71 22 23 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=0.797 $Y=1.015
+ $X2=0.797 $Y2=1.185
r72 20 22 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=0.685 $Y=0.93
+ $X2=0.797 $Y2=1.015
r73 20 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.685 $Y=0.93
+ $X2=0.355 $Y2=0.93
r74 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=0.845
+ $X2=0.355 $Y2=0.93
r75 16 18 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=0.845
+ $X2=0.225 $Y2=0.55
r76 14 35 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=1.4 $Y=1.35
+ $X2=0.955 $Y2=1.35
r77 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.4 $Y=1.35
+ $X2=1.475 $Y2=1.35
r78 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.515
+ $X2=1.475 $Y2=1.35
r79 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.475 $Y=1.515
+ $X2=1.475 $Y2=2.465
r80 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.185
+ $X2=1.475 $Y2=1.35
r81 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.475 $Y=1.185
+ $X2=1.475 $Y2=0.655
r82 2 27 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=2.015 $X2=0.735 $Y2=2.225
r83 1 18 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.345 $X2=0.26 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_1%A2 3 7 9 10 14
r34 14 17 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.94 $Y=1.51
+ $X2=1.94 $Y2=1.675
r35 14 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.94 $Y=1.51
+ $X2=1.94 $Y2=1.345
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.925
+ $Y=1.51 $X2=1.925 $Y2=1.51
r37 10 15 7.22198 $w=3.73e-07 $l=2.35e-07 $layer=LI1_cond $X=2.16 $Y=1.562
+ $X2=1.925 $Y2=1.562
r38 9 15 7.52929 $w=3.73e-07 $l=2.45e-07 $layer=LI1_cond $X=1.68 $Y=1.562
+ $X2=1.925 $Y2=1.562
r39 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.045 $Y=2.465
+ $X2=2.045 $Y2=1.675
r40 3 16 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.91 $Y=0.655
+ $X2=1.91 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_1%A1 3 7 9 14 15
r23 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.46 $X2=2.59 $Y2=1.46
r24 11 14 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.405 $Y=1.46
+ $X2=2.59 $Y2=1.46
r25 9 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.46
r26 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.625
+ $X2=2.405 $Y2=1.46
r27 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.405 $Y=1.625
+ $X2=2.405 $Y2=2.465
r28 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.295
+ $X2=2.405 $Y2=1.46
r29 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.405 $Y=1.295
+ $X2=2.405 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_1%VPWR 1 2 9 11 13 17 19 24 30 34
r31 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 25 30 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.247 $Y2=3.33
r36 25 27 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 24 33 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.455 $Y=3.33
+ $X2=2.667 $Y2=3.33
r38 24 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.455 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 19 30 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.07 $Y=3.33
+ $X2=1.247 $Y2=3.33
r42 19 21 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 17 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 17 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 13 16 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=2.62 $Y=2.005
+ $X2=2.62 $Y2=2.95
r46 11 33 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.62 $Y=3.245
+ $X2=2.667 $Y2=3.33
r47 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.62 $Y=3.245
+ $X2=2.62 $Y2=2.95
r48 7 30 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.247 $Y=3.245
+ $X2=1.247 $Y2=3.33
r49 7 9 28.0807 $w=3.53e-07 $l=8.65e-07 $layer=LI1_cond $X=1.247 $Y=3.245
+ $X2=1.247 $Y2=2.38
r50 2 16 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2.95
r51 2 13 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2.005
r52 1 9 300 $w=1.7e-07 $l=4.67974e-07 $layer=licon1_PDIFF $count=2 $X=1.025
+ $Y=2.015 $X2=1.26 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_1%Y 1 2 9 12 13 14 15 16 17 23
c39 12 0 5.38984e-20 $X=1.325 $Y=1.93
r40 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.76 $Y=2.405
+ $X2=1.76 $Y2=2.775
r41 15 23 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=2.015 $X2=1.76
+ $Y2=2.1
r42 15 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.76 $Y=2.11
+ $X2=1.76 $Y2=2.405
r43 15 23 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.76 $Y=2.11 $X2=1.76
+ $Y2=2.1
r44 14 15 8.01147 $w=3.18e-07 $l=1.85e-07 $layer=LI1_cond $X=1.41 $Y=2.015
+ $X2=1.595 $Y2=2.015
r45 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.325 $Y=1.93
+ $X2=1.41 $Y2=2.015
r46 12 13 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.325 $Y=1.93
+ $X2=1.325 $Y2=1.015
r47 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=0.85
+ $X2=1.245 $Y2=1.015
r48 7 9 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.245 $Y=0.85
+ $X2=1.245 $Y2=0.38
r49 2 15 600 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.835 $X2=1.76 $Y2=2.015
r50 2 16 300 $w=1.7e-07 $l=7.27461e-07 $layer=licon1_PDIFF $count=2 $X=1.55
+ $Y=1.835 $X2=1.76 $Y2=2.465
r51 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.12
+ $Y=0.235 $X2=1.245 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r38 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r41 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.145
+ $Y2=0
r43 27 29 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.64
+ $Y2=0
r44 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r45 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r46 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r47 23 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.68
+ $Y2=0
r48 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=0 $X2=2.145
+ $Y2=0
r49 22 25 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.98 $Y=0 $X2=1.68
+ $Y2=0
r50 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r51 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r53 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r54 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r55 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r56 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=0.085
+ $X2=2.145 $Y2=0
r57 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.145 $Y=0.085
+ $X2=2.145 $Y2=0.38
r58 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r59 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0.55
r60 2 13 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.985
+ $Y=0.235 $X2=2.145 $Y2=0.38
r61 1 9 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.345 $X2=0.69 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_1%A_310_47# 1 2 9 11 12 15
r21 13 15 23.2378 $w=3.03e-07 $l=6.15e-07 $layer=LI1_cond $X=2.632 $Y=1.035
+ $X2=2.632 $Y2=0.42
r22 11 13 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=2.48 $Y=1.12
+ $X2=2.632 $Y2=1.035
r23 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.48 $Y=1.12
+ $X2=1.81 $Y2=1.12
r24 7 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.695 $Y=1.035
+ $X2=1.81 $Y2=1.12
r25 7 9 30.8153 $w=2.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.695 $Y=1.035
+ $X2=1.695 $Y2=0.42
r26 2 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.48
+ $Y=0.235 $X2=2.62 $Y2=0.42
r27 1 9 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.55
+ $Y=0.235 $X2=1.695 $Y2=0.42
.ends

