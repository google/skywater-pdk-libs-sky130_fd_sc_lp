* File: sky130_fd_sc_lp__o21ba_lp.spice
* Created: Wed Sep  2 10:17:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ba_lp.pex.spice"
.subckt sky130_fd_sc_lp__o21ba_lp  VNB VPB A1 A2 B1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1_N	B1_N
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A1_M1001_g N_A_34_55#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.1197 PD=0.86 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1002 N_A_34_55#_M1002_d N_A2_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0924 PD=0.81 PS=0.86 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_253_389#_M1005_d N_A_317_29#_M1005_g N_A_34_55#_M1002_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0819 PD=1.41 PS=0.81 NRD=0 NRS=31.428 M=1 R=2.8
+ SA=75001.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_550_75# N_B1_N_M1007_g N_A_317_29#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B1_N_M1003_g A_550_75# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1011 A_708_75# N_A_253_389#_M1011_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_253_389#_M1009_g A_708_75# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_155_389# N_A1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1010 N_A_253_389#_M1010_d N_A2_M1010_g A_155_389# VPB PHIGHVT L=0.25 W=1
+ AD=0.16 AS=0.12 PD=1.32 PS=1.24 NRD=7.8603 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_A_317_29#_M1008_g N_A_253_389#_M1010_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.24175 AS=0.16 PD=1.59 PS=1.32 NRD=16.7253 NRS=0 M=1 R=4
+ SA=125001 SB=125001 A=0.25 P=2.5 MULT=1
MM1000 N_A_317_29#_M1000_d N_B1_N_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.24175 PD=2.57 PS=1.59 NRD=0 NRS=16.7253 M=1 R=4 SA=125002
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1006 N_X_M1006_d N_A_253_389#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__o21ba_lp.pxi.spice"
*
.ends
*
*
