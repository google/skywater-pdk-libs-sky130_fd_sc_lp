# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a2111o_m
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a2111o_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.700000 2.665000 3.205000 2.995000 ;
        RECT 2.890000 2.320000 3.205000 2.665000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 0.840000 3.205000 1.380000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 2.320000 1.765000 2.735000 ;
        RECT 1.500000 2.735000 2.170000 3.065000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 2.320000 1.330000 2.965000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.095000 1.295000 1.750000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 0.345000 0.390000 0.675000 ;
        RECT 0.155000 0.675000 0.325000 2.530000 ;
        RECT 0.155000 2.530000 0.390000 2.860000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
        RECT 0.570000  0.085000 0.900000 0.485000 ;
        RECT 1.690000  0.085000 1.900000 0.545000 ;
        RECT 2.850000  0.085000 3.180000 0.485000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 3.360000 3.415000 ;
        RECT 0.610000 2.645000 0.820000 3.245000 ;
        RECT 2.340000 2.305000 2.710000 2.495000 ;
        RECT 2.340000 2.495000 2.530000 3.245000 ;
        RECT 2.520000 1.955000 2.710000 2.305000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.505000 1.470000 0.675000 1.930000 ;
      RECT 0.505000 1.930000 1.645000 2.140000 ;
      RECT 1.260000 0.345000 1.470000 0.725000 ;
      RECT 1.260000 0.725000 2.330000 0.895000 ;
      RECT 1.475000 0.895000 1.645000 1.930000 ;
      RECT 2.090000 1.605000 3.260000 1.775000 ;
      RECT 2.090000 1.775000 2.300000 2.135000 ;
      RECT 2.120000 0.345000 2.330000 0.725000 ;
      RECT 2.930000 1.775000 3.260000 2.095000 ;
  END
END sky130_fd_sc_lp__a2111o_m
