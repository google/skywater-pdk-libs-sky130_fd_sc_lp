# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__ha_0
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__ha_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.055000 2.800000 1.385000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.915000 3.270000 2.295000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.255000 2.435000 4.715000 3.075000 ;
        RECT 4.355000 0.375000 4.715000 1.425000 ;
        RECT 4.435000 1.425000 4.715000 2.435000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.293700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.385000 0.425000 1.425000 ;
        RECT 0.095000 1.425000 0.325000 2.495000 ;
        RECT 0.095000 2.495000 0.500000 3.075000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.800000 0.085000 ;
        RECT 0.595000  0.085000 0.805000 0.805000 ;
        RECT 1.940000  0.085000 2.270000 0.545000 ;
        RECT 3.855000  0.085000 4.185000 1.050000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.800000 3.415000 ;
        RECT 0.670000 2.435000 1.000000 3.245000 ;
        RECT 2.330000 2.500000 3.180000 3.245000 ;
        RECT 3.780000 2.435000 4.085000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.505000 1.595000 1.145000 2.095000 ;
      RECT 0.505000 2.095000 1.415000 2.265000 ;
      RECT 0.975000 0.280000 1.390000 0.610000 ;
      RECT 0.975000 0.610000 1.145000 1.595000 ;
      RECT 1.170000 2.265000 1.415000 2.500000 ;
      RECT 1.170000 2.500000 1.840000 2.830000 ;
      RECT 1.315000 1.055000 1.575000 1.565000 ;
      RECT 1.315000 1.565000 3.610000 1.595000 ;
      RECT 1.315000 1.595000 4.265000 1.735000 ;
      RECT 1.560000 0.280000 1.770000 0.715000 ;
      RECT 1.560000 0.715000 2.700000 0.885000 ;
      RECT 2.440000 0.280000 2.700000 0.715000 ;
      RECT 3.010000 0.720000 3.610000 1.565000 ;
      RECT 3.350000 2.500000 3.610000 2.830000 ;
      RECT 3.440000 1.735000 4.265000 2.265000 ;
      RECT 3.440000 2.265000 3.610000 2.500000 ;
  END
END sky130_fd_sc_lp__ha_0
