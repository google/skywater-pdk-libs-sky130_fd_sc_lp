* NGSPICE file created from sky130_fd_sc_lp__nor4bb_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor4bb_m A B C_N D_N VGND VNB VPB VPWR Y
M1000 VGND A Y VNB nshort w=420000u l=150000u
+  ad=5.46e+11p pd=5.12e+06u as=2.352e+11p ps=2.8e+06u
M1001 VPWR A a_454_397# VPB phighvt w=420000u l=150000u
+  ad=3.696e+11p pd=3.44e+06u as=8.82e+10p ps=1.26e+06u
M1002 VGND D_N a_27_507# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 a_310_397# a_27_507# Y VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1004 Y a_27_507# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_284_99# C_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 a_382_397# a_284_99# a_310_397# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 a_284_99# C_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 VGND a_284_99# Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_454_397# B a_382_397# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR D_N a_27_507# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 Y B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

