* File: sky130_fd_sc_lp__clkdlybuf4s25_1.pxi.spice
* Created: Fri Aug 28 10:16:50 2020
* 
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%A N_A_M1003_g N_A_M1007_g A A N_A_c_62_n
+ PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%A
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%A_27_52# N_A_27_52#_M1003_s
+ N_A_27_52#_M1007_s N_A_27_52#_c_95_n N_A_27_52#_M1004_g N_A_27_52#_c_96_n
+ N_A_27_52#_M1002_g N_A_27_52#_c_97_n N_A_27_52#_c_104_n N_A_27_52#_c_105_n
+ N_A_27_52#_c_98_n N_A_27_52#_c_99_n N_A_27_52#_c_106_n N_A_27_52#_c_100_n
+ N_A_27_52#_c_101_n PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%A_27_52#
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%A_282_52# N_A_282_52#_M1004_d
+ N_A_282_52#_M1002_d N_A_282_52#_c_162_n N_A_282_52#_M1006_g
+ N_A_282_52#_M1001_g N_A_282_52#_c_163_n N_A_282_52#_c_164_n
+ N_A_282_52#_c_168_n N_A_282_52#_c_165_n N_A_282_52#_c_166_n
+ N_A_282_52#_c_170_n PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%A_282_52#
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%A_394_52# N_A_394_52#_M1006_s
+ N_A_394_52#_M1001_s N_A_394_52#_M1005_g N_A_394_52#_M1000_g
+ N_A_394_52#_c_234_n N_A_394_52#_c_236_n N_A_394_52#_c_239_n
+ N_A_394_52#_c_229_n N_A_394_52#_c_230_n N_A_394_52#_c_225_n
+ N_A_394_52#_c_226_n N_A_394_52#_c_257_n N_A_394_52#_c_227_n
+ PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%A_394_52#
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%VPWR N_VPWR_M1007_d N_VPWR_M1001_d
+ N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n VPWR
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_294_n N_VPWR_c_302_n
+ PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%VPWR
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%X N_X_M1005_d N_X_M1000_d X X X X X X X
+ N_X_c_337_n N_X_c_340_n X PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%X
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%VGND N_VGND_M1003_d N_VGND_M1006_d
+ N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n VGND
+ N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n
+ PM_SKY130_FD_SC_LP__CLKDLYBUF4S25_1%VGND
cc_1 VNB N_A_M1003_g 0.0647104f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.47
cc_2 VNB A 0.0208018f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A_c_62_n 0.0329141f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_4 VNB N_A_27_52#_c_95_n 0.0276919f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_5 VNB N_A_27_52#_c_96_n 0.0421651f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_27_52#_c_97_n 0.0205357f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.335
cc_7 VNB N_A_27_52#_c_98_n 0.0050785f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.665
cc_8 VNB N_A_27_52#_c_99_n 0.0115829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_52#_c_100_n 0.00219081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_52#_c_101_n 9.66126e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_282_52#_c_162_n 0.0288054f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_12 VNB N_A_282_52#_c_163_n 0.011676f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.335
cc_13 VNB N_A_282_52#_c_164_n 0.0150178f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.295
cc_14 VNB N_A_282_52#_c_165_n 0.0124045f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.665
cc_15 VNB N_A_282_52#_c_166_n 0.0456811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_394_52#_M1005_g 0.0568356f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A_394_52#_M1000_g 0.00175473f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_18 VNB N_A_394_52#_c_225_n 0.014306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_394_52#_c_226_n 4.63484e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_394_52#_c_227_n 0.0354556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_294_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB X 0.0542411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_337_n 0.0186904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_360_n 0.00646702f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_25 VNB N_VGND_c_361_n 0.00646199f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_26 VNB N_VGND_c_362_n 0.0512685f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.335
cc_27 VNB N_VGND_c_363_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.665
cc_28 VNB N_VGND_c_364_n 0.0179296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_365_n 0.0230432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_366_n 0.241616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_367_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_A_M1007_g 0.0257865f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_33 VPB A 0.00827303f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_34 VPB N_A_c_62_n 0.00600603f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_35 VPB N_A_27_52#_c_96_n 0.043701f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_36 VPB N_A_27_52#_M1002_g 0.0314916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_27_52#_c_104_n 0.00794922f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.295
cc_38 VPB N_A_27_52#_c_105_n 0.0339238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_52#_c_106_n 0.00375793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_27_52#_c_100_n 0.00497175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_282_52#_M1001_g 0.0509536f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_282_52#_c_168_n 0.0102217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_282_52#_c_166_n 0.017645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_282_52#_c_170_n 0.0138541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_394_52#_M1000_g 0.0265621f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_46 VPB N_A_394_52#_c_229_n 0.0112289f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_394_52#_c_230_n 0.0040145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_394_52#_c_226_n 0.00362728f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_295_n 0.00558649f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_50 VPB N_VPWR_c_296_n 0.00563065f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_51 VPB N_VPWR_c_297_n 0.0498697f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.295
cc_52 VPB N_VPWR_c_298_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_299_n 0.0178675f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.665
cc_54 VPB N_VPWR_c_300_n 0.0226035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_294_n 0.0532965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_302_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB X 0.00848832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB X 0.0499319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_X_c_340_n 0.0178335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 A N_A_27_52#_M1007_s 0.00237131f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_A_M1003_g N_A_27_52#_c_95_n 0.0161521f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_62 A N_A_27_52#_c_96_n 0.00135678f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A_c_62_n N_A_27_52#_c_96_n 0.0175907f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_64 N_A_M1007_g N_A_27_52#_M1002_g 0.0186474f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_65 N_A_M1003_g N_A_27_52#_c_97_n 0.013604f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_66 N_A_M1007_g N_A_27_52#_c_104_n 7.4234e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_67 A N_A_27_52#_c_104_n 0.0239868f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A_c_62_n N_A_27_52#_c_104_n 7.87914e-19 $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_69 N_A_M1007_g N_A_27_52#_c_105_n 0.0151418f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_M1003_g N_A_27_52#_c_98_n 0.0116934f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_71 A N_A_27_52#_c_98_n 0.0106601f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_M1003_g N_A_27_52#_c_99_n 0.00435937f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_73 A N_A_27_52#_c_99_n 0.0289379f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_c_62_n N_A_27_52#_c_99_n 0.00100334f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_75 N_A_M1007_g N_A_27_52#_c_106_n 0.0125269f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_76 A N_A_27_52#_c_106_n 0.00941865f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_M1007_g N_A_27_52#_c_100_n 0.00214268f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_78 A N_A_27_52#_c_100_n 0.0114464f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A_c_62_n N_A_27_52#_c_100_n 0.0013726f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_80 N_A_M1003_g N_A_27_52#_c_101_n 0.00511688f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_81 A N_A_27_52#_c_101_n 0.0179575f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_c_62_n N_A_27_52#_c_101_n 9.52655e-19 $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_83 N_A_M1007_g N_VPWR_c_295_n 0.00922071f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_84 N_A_M1007_g N_VPWR_c_299_n 0.0054895f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_M1007_g N_VPWR_c_294_n 0.0114819f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A_M1003_g N_VGND_c_360_n 0.00360601f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_87 N_A_M1003_g N_VGND_c_364_n 0.00547602f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_VGND_c_366_n 0.00732141f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_89 N_A_27_52#_c_96_n N_A_282_52#_M1001_g 0.00272427f $X=1.285 $Y=1.93 $X2=0
+ $Y2=0
cc_90 N_A_27_52#_c_95_n N_A_282_52#_c_164_n 0.00532265f $X=1.285 $Y=1.37 $X2=0
+ $Y2=0
cc_91 N_A_27_52#_c_96_n N_A_282_52#_c_164_n 0.00414437f $X=1.285 $Y=1.93 $X2=0
+ $Y2=0
cc_92 N_A_27_52#_c_100_n N_A_282_52#_c_164_n 0.00828764f $X=1.087 $Y=1.6 $X2=0
+ $Y2=0
cc_93 N_A_27_52#_c_101_n N_A_282_52#_c_164_n 0.022177f $X=1.085 $Y=1.535 $X2=0
+ $Y2=0
cc_94 N_A_27_52#_c_96_n N_A_282_52#_c_168_n 0.00361912f $X=1.285 $Y=1.93 $X2=0
+ $Y2=0
cc_95 N_A_27_52#_M1002_g N_A_282_52#_c_168_n 0.00350396f $X=1.285 $Y=2.595 $X2=0
+ $Y2=0
cc_96 N_A_27_52#_c_100_n N_A_282_52#_c_168_n 0.0285056f $X=1.087 $Y=1.6 $X2=0
+ $Y2=0
cc_97 N_A_27_52#_c_96_n N_A_282_52#_c_166_n 0.00552637f $X=1.285 $Y=1.93 $X2=0
+ $Y2=0
cc_98 N_A_27_52#_c_96_n N_A_282_52#_c_170_n 0.00392394f $X=1.285 $Y=1.93 $X2=0
+ $Y2=0
cc_99 N_A_27_52#_M1002_g N_A_282_52#_c_170_n 0.0145229f $X=1.285 $Y=2.595 $X2=0
+ $Y2=0
cc_100 N_A_27_52#_c_100_n N_A_282_52#_c_170_n 0.00501863f $X=1.087 $Y=1.6 $X2=0
+ $Y2=0
cc_101 N_A_27_52#_c_106_n N_VPWR_M1007_d 0.0115736f $X=0.91 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_27_52#_c_100_n N_VPWR_M1007_d 0.00859969f $X=1.087 $Y=1.6 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_27_52#_M1002_g N_VPWR_c_295_n 0.0110096f $X=1.285 $Y=2.595 $X2=0
+ $Y2=0
cc_104 N_A_27_52#_c_106_n N_VPWR_c_295_n 0.0241337f $X=0.91 $Y=2.117 $X2=0 $Y2=0
cc_105 N_A_27_52#_c_100_n N_VPWR_c_295_n 0.00123499f $X=1.087 $Y=1.6 $X2=0 $Y2=0
cc_106 N_A_27_52#_M1002_g N_VPWR_c_297_n 0.00937688f $X=1.285 $Y=2.595 $X2=0
+ $Y2=0
cc_107 N_A_27_52#_c_105_n N_VPWR_c_299_n 0.0210467f $X=0.26 $Y=2.915 $X2=0 $Y2=0
cc_108 N_A_27_52#_M1007_s N_VPWR_c_294_n 0.00215158f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_109 N_A_27_52#_M1002_g N_VPWR_c_294_n 0.0181716f $X=1.285 $Y=2.595 $X2=0
+ $Y2=0
cc_110 N_A_27_52#_c_105_n N_VPWR_c_294_n 0.0125689f $X=0.26 $Y=2.915 $X2=0 $Y2=0
cc_111 N_A_27_52#_c_98_n N_VGND_M1003_d 0.0195513f $X=0.91 $Y=0.92 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_27_52#_c_101_n N_VGND_M1003_d 0.00404045f $X=1.085 $Y=1.535 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_27_52#_c_95_n N_VGND_c_360_n 0.00723954f $X=1.285 $Y=1.37 $X2=0 $Y2=0
cc_114 N_A_27_52#_c_98_n N_VGND_c_360_n 0.0252704f $X=0.91 $Y=0.92 $X2=0 $Y2=0
cc_115 N_A_27_52#_c_95_n N_VGND_c_362_n 0.00933598f $X=1.285 $Y=1.37 $X2=0 $Y2=0
cc_116 N_A_27_52#_c_97_n N_VGND_c_364_n 0.0152237f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_117 N_A_27_52#_c_95_n N_VGND_c_366_n 0.0154889f $X=1.285 $Y=1.37 $X2=0 $Y2=0
cc_118 N_A_27_52#_c_97_n N_VGND_c_366_n 0.0118277f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_119 N_A_27_52#_c_98_n N_VGND_c_366_n 0.0196037f $X=0.91 $Y=0.92 $X2=0 $Y2=0
cc_120 N_A_282_52#_c_162_n N_A_394_52#_M1005_g 0.0196394f $X=2.36 $Y=1.37 $X2=0
+ $Y2=0
cc_121 N_A_282_52#_M1001_g N_A_394_52#_M1000_g 0.0187947f $X=2.36 $Y=2.595 $X2=0
+ $Y2=0
cc_122 N_A_282_52#_c_162_n N_A_394_52#_c_234_n 0.0257681f $X=2.36 $Y=1.37 $X2=0
+ $Y2=0
cc_123 N_A_282_52#_c_163_n N_A_394_52#_c_234_n 0.0577683f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_124 N_A_282_52#_c_162_n N_A_394_52#_c_236_n 0.0226716f $X=2.36 $Y=1.37 $X2=0
+ $Y2=0
cc_125 N_A_282_52#_c_165_n N_A_394_52#_c_236_n 0.0288942f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_126 N_A_282_52#_c_166_n N_A_394_52#_c_236_n 0.00585462f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_127 N_A_282_52#_c_162_n N_A_394_52#_c_239_n 8.78991e-19 $X=2.36 $Y=1.37 $X2=0
+ $Y2=0
cc_128 N_A_282_52#_c_163_n N_A_394_52#_c_239_n 0.00858119f $X=1.55 $Y=0.435
+ $X2=0 $Y2=0
cc_129 N_A_282_52#_c_164_n N_A_394_52#_c_239_n 0.0121129f $X=1.755 $Y=1.655
+ $X2=0 $Y2=0
cc_130 N_A_282_52#_c_165_n N_A_394_52#_c_239_n 0.0177106f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_131 N_A_282_52#_c_166_n N_A_394_52#_c_239_n 0.00503939f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_132 N_A_282_52#_c_165_n N_A_394_52#_c_229_n 0.0106947f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_133 N_A_282_52#_c_166_n N_A_394_52#_c_229_n 0.0048475f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_134 N_A_282_52#_M1001_g N_A_394_52#_c_230_n 0.0325688f $X=2.36 $Y=2.595 $X2=0
+ $Y2=0
cc_135 N_A_282_52#_c_168_n N_A_394_52#_c_230_n 0.00990869f $X=1.755 $Y=2.1 $X2=0
+ $Y2=0
cc_136 N_A_282_52#_c_165_n N_A_394_52#_c_230_n 0.0272343f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_137 N_A_282_52#_c_166_n N_A_394_52#_c_230_n 0.00593164f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_138 N_A_282_52#_c_170_n N_A_394_52#_c_230_n 0.0129926f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_139 N_A_282_52#_c_162_n N_A_394_52#_c_225_n 0.0032529f $X=2.36 $Y=1.37 $X2=0
+ $Y2=0
cc_140 N_A_282_52#_c_165_n N_A_394_52#_c_225_n 0.0207685f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_141 N_A_282_52#_c_166_n N_A_394_52#_c_225_n 0.0027866f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_142 N_A_282_52#_M1001_g N_A_394_52#_c_226_n 0.00236812f $X=2.36 $Y=2.595
+ $X2=0 $Y2=0
cc_143 N_A_282_52#_c_165_n N_A_394_52#_c_226_n 0.00227963f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_144 N_A_282_52#_c_166_n N_A_394_52#_c_226_n 0.00140233f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_145 N_A_282_52#_M1001_g N_A_394_52#_c_257_n 0.021788f $X=2.36 $Y=2.595 $X2=0
+ $Y2=0
cc_146 N_A_282_52#_c_170_n N_A_394_52#_c_257_n 0.0679402f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_147 N_A_282_52#_c_166_n N_A_394_52#_c_227_n 0.0101747f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_148 N_A_282_52#_c_170_n N_VPWR_c_295_n 0.0250587f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_149 N_A_282_52#_M1001_g N_VPWR_c_296_n 0.0130235f $X=2.36 $Y=2.595 $X2=0
+ $Y2=0
cc_150 N_A_282_52#_M1001_g N_VPWR_c_297_n 0.00939206f $X=2.36 $Y=2.595 $X2=0
+ $Y2=0
cc_151 N_A_282_52#_c_170_n N_VPWR_c_297_n 0.0301474f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_152 N_A_282_52#_M1002_d N_VPWR_c_294_n 0.00215158f $X=1.41 $Y=2.095 $X2=0
+ $Y2=0
cc_153 N_A_282_52#_M1001_g N_VPWR_c_294_n 0.0182087f $X=2.36 $Y=2.595 $X2=0
+ $Y2=0
cc_154 N_A_282_52#_c_170_n N_VPWR_c_294_n 0.0175018f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_155 N_A_282_52#_c_162_n N_VGND_c_361_n 0.00753134f $X=2.36 $Y=1.37 $X2=0
+ $Y2=0
cc_156 N_A_282_52#_c_162_n N_VGND_c_362_n 0.00899047f $X=2.36 $Y=1.37 $X2=0
+ $Y2=0
cc_157 N_A_282_52#_c_163_n N_VGND_c_362_n 0.0250858f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_158 N_A_282_52#_c_162_n N_VGND_c_366_n 0.0177497f $X=2.36 $Y=1.37 $X2=0 $Y2=0
cc_159 N_A_282_52#_c_163_n N_VGND_c_366_n 0.0155553f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_160 N_A_394_52#_c_229_n N_VPWR_M1001_d 0.00502062f $X=2.855 $Y=1.91 $X2=0
+ $Y2=0
cc_161 N_A_394_52#_M1000_g N_VPWR_c_296_n 0.0107614f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_394_52#_c_229_n N_VPWR_c_296_n 0.027185f $X=2.855 $Y=1.91 $X2=0 $Y2=0
cc_163 N_A_394_52#_c_225_n N_VPWR_c_296_n 5.09408e-19 $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_164 N_A_394_52#_c_257_n N_VPWR_c_296_n 0.0295704f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_165 N_A_394_52#_c_257_n N_VPWR_c_297_n 0.0153681f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_166 N_A_394_52#_M1000_g N_VPWR_c_300_n 0.00564131f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_394_52#_M1001_s N_VPWR_c_294_n 0.00357787f $X=1.97 $Y=2.095 $X2=0
+ $Y2=0
cc_168 N_A_394_52#_M1000_g N_VPWR_c_294_n 0.0120194f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_394_52#_c_257_n N_VPWR_c_294_n 0.00945867f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_170 N_A_394_52#_M1005_g X 0.0163897f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_171 N_A_394_52#_M1000_g X 0.00381153f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A_394_52#_c_225_n X 0.0389414f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_173 N_A_394_52#_c_226_n X 0.00696747f $X=2.94 $Y=1.825 $X2=0 $Y2=0
cc_174 N_A_394_52#_c_227_n X 0.00819462f $X=3.26 $Y=1.46 $X2=0 $Y2=0
cc_175 N_A_394_52#_M1000_g X 0.0170331f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_394_52#_M1005_g N_X_c_337_n 0.00509113f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_177 N_A_394_52#_c_225_n N_X_c_337_n 0.00268942f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_178 N_A_394_52#_c_227_n N_X_c_337_n 0.00229273f $X=3.26 $Y=1.46 $X2=0 $Y2=0
cc_179 N_A_394_52#_M1000_g N_X_c_340_n 0.00618036f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_394_52#_c_229_n N_X_c_340_n 0.012527f $X=2.855 $Y=1.91 $X2=0 $Y2=0
cc_181 N_A_394_52#_c_225_n N_X_c_340_n 0.00881742f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_182 N_A_394_52#_c_226_n N_X_c_340_n 6.43138e-19 $X=2.94 $Y=1.825 $X2=0 $Y2=0
cc_183 N_A_394_52#_c_227_n N_X_c_340_n 0.00425967f $X=3.26 $Y=1.46 $X2=0 $Y2=0
cc_184 N_A_394_52#_c_236_n N_VGND_M1006_d 0.0152079f $X=2.855 $Y=1.097 $X2=0
+ $Y2=0
cc_185 N_A_394_52#_c_225_n N_VGND_M1006_d 0.00394571f $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_186 N_A_394_52#_M1005_g N_VGND_c_361_n 0.00659723f $X=3.17 $Y=0.47 $X2=0
+ $Y2=0
cc_187 N_A_394_52#_c_234_n N_VGND_c_361_n 0.0143451f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_188 N_A_394_52#_c_236_n N_VGND_c_361_n 0.0076609f $X=2.855 $Y=1.097 $X2=0
+ $Y2=0
cc_189 N_A_394_52#_c_225_n N_VGND_c_361_n 0.0103475f $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_190 N_A_394_52#_c_234_n N_VGND_c_362_n 0.0140261f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_191 N_A_394_52#_M1005_g N_VGND_c_365_n 0.0051159f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_192 N_A_394_52#_M1005_g N_VGND_c_366_n 0.0107972f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_193 N_A_394_52#_c_234_n N_VGND_c_366_n 0.00945114f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_294_n N_X_M1000_d 0.00215158f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_300_n X 0.0347023f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_294_n X 0.0200014f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_197 N_X_c_337_n N_VGND_c_365_n 0.0254f $X=3.632 $Y=0.475 $X2=0 $Y2=0
cc_198 N_X_c_337_n N_VGND_c_366_n 0.0197894f $X=3.632 $Y=0.475 $X2=0 $Y2=0
