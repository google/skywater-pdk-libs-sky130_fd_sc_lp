* File: sky130_fd_sc_lp__and4_4.pex.spice
* Created: Fri Aug 28 10:07:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4_4%A 1 3 4 6 7 8
c21 7 0 1.68603e-19 $X=0.24 $Y=1.295
r22 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.375 $X2=0.37 $Y2=1.375
r23 8 13 9.41432 $w=3.53e-07 $l=2.9e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.375
r24 7 13 2.59705 $w=3.53e-07 $l=8e-08 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.375
r25 4 12 60.9298 $w=4.31e-07 $l=4.28661e-07 $layer=POLY_cond $X=0.63 $Y=1.725
+ $X2=0.455 $Y2=1.375
r26 4 6 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.63 $Y=1.725 $X2=0.63
+ $Y2=2.465
r27 1 12 43.0365 $w=4.31e-07 $l=2.63344e-07 $layer=POLY_cond $X=0.63 $Y=1.185
+ $X2=0.455 $Y2=1.375
r28 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.63 $Y=1.185 $X2=0.63
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_4%B 3 6 8 9 13 15
c35 13 0 1.68603e-19 $X=1.08 $Y=1.35
c36 6 0 1.35108e-19 $X=1.06 $Y=2.465
r37 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.08 $Y=1.35
+ $X2=1.08 $Y2=1.515
r38 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.08 $Y=1.35
+ $X2=1.08 $Y2=1.185
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.35 $X2=1.08 $Y2=1.35
r40 9 14 4.39026 $w=3.13e-07 $l=1.2e-07 $layer=LI1_cond $X=1.2 $Y=1.357 $X2=1.08
+ $Y2=1.357
r41 8 14 13.1708 $w=3.13e-07 $l=3.6e-07 $layer=LI1_cond $X=0.72 $Y=1.357
+ $X2=1.08 $Y2=1.357
r42 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.06 $Y=2.465
+ $X2=1.06 $Y2=1.515
r43 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.99 $Y=0.655
+ $X2=0.99 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_4%C 3 7 9 12
c34 9 0 1.35108e-19 $X=1.68 $Y=1.295
c35 3 0 8.28477e-21 $X=1.53 $Y=0.655
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.375
+ $X2=1.62 $Y2=1.54
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.375
+ $X2=1.62 $Y2=1.21
r38 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.375 $X2=1.62 $Y2=1.375
r39 7 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.64 $Y=2.465
+ $X2=1.64 $Y2=1.54
r40 3 14 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.53 $Y=0.655
+ $X2=1.53 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_4%D 3 7 9 12
c37 9 0 8.28477e-21 $X=2.16 $Y=1.295
r38 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.375
+ $X2=2.16 $Y2=1.54
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.375
+ $X2=2.16 $Y2=1.21
r40 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.375 $X2=2.16 $Y2=1.375
r41 7 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.07 $Y=2.465
+ $X2=2.07 $Y2=1.54
r42 3 14 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.07 $Y=0.655
+ $X2=2.07 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_4%A_58_47# 1 2 3 12 16 20 24 28 32 36 40 44 46
+ 47 50 54 55 58 62 65 67 73 74 76 77
r147 82 83 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.505 $Y=1.5
+ $X2=3.935 $Y2=1.5
r148 81 82 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.075 $Y=1.5
+ $X2=3.505 $Y2=1.5
r149 74 83 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=4.095 $Y=1.5
+ $X2=3.935 $Y2=1.5
r150 73 74 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.095
+ $Y=1.5 $X2=4.095 $Y2=1.5
r151 71 81 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.735 $Y=1.5
+ $X2=3.075 $Y2=1.5
r152 71 78 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.735 $Y=1.5
+ $X2=2.645 $Y2=1.5
r153 70 73 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.735 $Y=1.5
+ $X2=4.095 $Y2=1.5
r154 70 71 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.735
+ $Y=1.5 $X2=2.735 $Y2=1.5
r155 68 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.5
+ $X2=2.51 $Y2=1.5
r156 68 70 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.595 $Y=1.5
+ $X2=2.735 $Y2=1.5
r157 66 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.585
+ $X2=2.51 $Y2=1.5
r158 66 67 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.51 $Y=1.585
+ $X2=2.51 $Y2=1.755
r159 65 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.415
+ $X2=2.51 $Y2=1.5
r160 64 65 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.51 $Y=1.03
+ $X2=2.51 $Y2=1.415
r161 63 76 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=2.01 $Y=1.84
+ $X2=1.847 $Y2=1.84
r162 62 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.425 $Y=1.84
+ $X2=2.51 $Y2=1.755
r163 62 63 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.425 $Y=1.84
+ $X2=2.01 $Y2=1.84
r164 58 60 32.9776 $w=3.23e-07 $l=9.3e-07 $layer=LI1_cond $X=1.847 $Y=1.98
+ $X2=1.847 $Y2=2.91
r165 56 76 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.847 $Y=1.925
+ $X2=1.847 $Y2=1.84
r166 56 58 1.95029 $w=3.23e-07 $l=5.5e-08 $layer=LI1_cond $X=1.847 $Y=1.925
+ $X2=1.847 $Y2=1.98
r167 54 76 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=1.685 $Y=1.84
+ $X2=1.847 $Y2=1.84
r168 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.685 $Y=1.84
+ $X2=1.015 $Y2=1.84
r169 50 52 40.4442 $w=2.63e-07 $l=9.3e-07 $layer=LI1_cond $X=0.882 $Y=1.98
+ $X2=0.882 $Y2=2.91
r170 48 55 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.882 $Y=1.925
+ $X2=1.015 $Y2=1.84
r171 48 50 2.39186 $w=2.63e-07 $l=5.5e-08 $layer=LI1_cond $X=0.882 $Y=1.925
+ $X2=0.882 $Y2=1.98
r172 46 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.425 $Y=0.945
+ $X2=2.51 $Y2=1.03
r173 46 47 125.588 $w=1.68e-07 $l=1.925e-06 $layer=LI1_cond $X=2.425 $Y=0.945
+ $X2=0.5 $Y2=0.945
r174 42 47 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.405 $Y=0.86
+ $X2=0.5 $Y2=0.945
r175 42 44 19.555 $w=1.88e-07 $l=3.35e-07 $layer=LI1_cond $X=0.405 $Y=0.86
+ $X2=0.405 $Y2=0.525
r176 38 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.935 $Y=1.665
+ $X2=3.935 $Y2=1.5
r177 38 40 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.935 $Y=1.665
+ $X2=3.935 $Y2=2.465
r178 34 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.935 $Y=1.335
+ $X2=3.935 $Y2=1.5
r179 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.935 $Y=1.335
+ $X2=3.935 $Y2=0.655
r180 30 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.665
+ $X2=3.505 $Y2=1.5
r181 30 32 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.505 $Y=1.665
+ $X2=3.505 $Y2=2.465
r182 26 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.335
+ $X2=3.505 $Y2=1.5
r183 26 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.505 $Y=1.335
+ $X2=3.505 $Y2=0.655
r184 22 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.665
+ $X2=3.075 $Y2=1.5
r185 22 24 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.075 $Y=1.665
+ $X2=3.075 $Y2=2.465
r186 18 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.335
+ $X2=3.075 $Y2=1.5
r187 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.075 $Y=1.335
+ $X2=3.075 $Y2=0.655
r188 14 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.665
+ $X2=2.645 $Y2=1.5
r189 14 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.645 $Y=1.665
+ $X2=2.645 $Y2=2.465
r190 10 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.335
+ $X2=2.645 $Y2=1.5
r191 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.645 $Y=1.335
+ $X2=2.645 $Y2=0.655
r192 3 60 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=1.835 $X2=1.855 $Y2=2.91
r193 3 58 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=1.835 $X2=1.855 $Y2=1.98
r194 2 52 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.705
+ $Y=1.835 $X2=0.845 $Y2=2.91
r195 2 50 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.705
+ $Y=1.835 $X2=0.845 $Y2=1.98
r196 1 44 91 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=2 $X=0.29
+ $Y=0.235 $X2=0.415 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_4%VPWR 1 2 3 4 5 16 18 22 26 32 38 44 49 50 52
+ 53 54 63 69 70 76 79
r66 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r68 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r70 70 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r71 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r72 67 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.15 $Y2=3.33
r73 67 69 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.56 $Y2=3.33
r74 66 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r75 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r76 63 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=4.15 $Y2=3.33
r77 63 65 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r78 62 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r79 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r80 59 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r81 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 56 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.35 $Y2=3.33
r83 56 58 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 54 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 54 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r86 52 61 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=3.12 $Y2=3.33
r87 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=3.29 $Y2=3.33
r88 51 65 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.455 $Y=3.33
+ $X2=3.6 $Y2=3.33
r89 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=3.33
+ $X2=3.29 $Y2=3.33
r90 49 58 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.18 $Y=3.33 $X2=2.16
+ $Y2=3.33
r91 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=3.33
+ $X2=2.345 $Y2=3.33
r92 48 61 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.51 $Y=3.33
+ $X2=3.12 $Y2=3.33
r93 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=3.33
+ $X2=2.345 $Y2=3.33
r94 44 47 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=4.15 $Y=2.2 $X2=4.15
+ $Y2=2.95
r95 42 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.15 $Y=3.245
+ $X2=4.15 $Y2=3.33
r96 42 47 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.15 $Y=3.245
+ $X2=4.15 $Y2=2.95
r97 38 41 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.29 $Y=2.2 $X2=3.29
+ $Y2=2.97
r98 36 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=3.245
+ $X2=3.29 $Y2=3.33
r99 36 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.29 $Y=3.245
+ $X2=3.29 $Y2=2.97
r100 32 35 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.345 $Y=2.19
+ $X2=2.345 $Y2=2.95
r101 30 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=3.245
+ $X2=2.345 $Y2=3.33
r102 30 35 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.245
+ $X2=2.345 $Y2=2.95
r103 26 29 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.35 $Y=2.19
+ $X2=1.35 $Y2=2.95
r104 24 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=3.245
+ $X2=1.35 $Y2=3.33
r105 24 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.35 $Y=3.245
+ $X2=1.35 $Y2=2.95
r106 23 73 4.50438 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.29 $Y2=3.33
r107 22 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=3.33
+ $X2=1.35 $Y2=3.33
r108 22 23 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.185 $Y=3.33
+ $X2=0.58 $Y2=3.33
r109 18 21 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.415 $Y=2.005
+ $X2=0.415 $Y2=2.95
r110 16 73 3.26179 $w=3.3e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.415 $Y=3.245
+ $X2=0.29 $Y2=3.33
r111 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.415 $Y=3.245
+ $X2=0.415 $Y2=2.95
r112 5 47 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.01
+ $Y=1.835 $X2=4.15 $Y2=2.95
r113 5 44 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=4.01
+ $Y=1.835 $X2=4.15 $Y2=2.2
r114 4 41 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.835 $X2=3.29 $Y2=2.97
r115 4 38 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.835 $X2=3.29 $Y2=2.2
r116 3 35 400 $w=1.7e-07 $l=1.21088e-06 $layer=licon1_PDIFF $count=1 $X=2.145
+ $Y=1.835 $X2=2.345 $Y2=2.95
r117 3 32 400 $w=1.7e-07 $l=4.43875e-07 $layer=licon1_PDIFF $count=1 $X=2.145
+ $Y=1.835 $X2=2.345 $Y2=2.19
r118 2 29 400 $w=1.7e-07 $l=1.21776e-06 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.835 $X2=1.35 $Y2=2.95
r119 2 26 400 $w=1.7e-07 $l=4.49833e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.835 $X2=1.35 $Y2=2.19
r120 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.29
+ $Y=1.835 $X2=0.415 $Y2=2.95
r121 1 18 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.29
+ $Y=1.835 $X2=0.415 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_4%X 1 2 3 4 15 21 23 24 25 26 29 33 37 39 41 42
+ 44 45 46 47 61
r68 59 61 2.56098 $w=2.68e-07 $l=6e-08 $layer=LI1_cond $X=4.565 $Y=1.235
+ $X2=4.565 $Y2=1.295
r69 46 53 3.49088 $w=2.67e-07 $l=8.59942e-08 $layer=LI1_cond $X=4.565 $Y=1.15
+ $X2=4.567 $Y2=1.065
r70 46 59 3.49088 $w=2.67e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=1.15
+ $X2=4.565 $Y2=1.235
r71 46 47 15.2805 $w=2.68e-07 $l=3.58e-07 $layer=LI1_cond $X=4.565 $Y=1.307
+ $X2=4.565 $Y2=1.665
r72 46 61 0.512197 $w=2.68e-07 $l=1.2e-08 $layer=LI1_cond $X=4.565 $Y=1.307
+ $X2=4.565 $Y2=1.295
r73 45 53 6.08838 $w=2.63e-07 $l=1.4e-07 $layer=LI1_cond $X=4.567 $Y=0.925
+ $X2=4.567 $Y2=1.065
r74 44 45 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=4.567 $Y=0.555
+ $X2=4.567 $Y2=0.925
r75 43 47 4.69514 $w=2.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.565 $Y=1.775
+ $X2=4.565 $Y2=1.665
r76 40 41 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.865 $Y=1.15
+ $X2=3.745 $Y2=1.15
r77 39 46 3.01551 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.43 $Y=1.15
+ $X2=4.565 $Y2=1.15
r78 39 40 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.43 $Y=1.15
+ $X2=3.865 $Y2=1.15
r79 38 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.815 $Y=1.86
+ $X2=3.72 $Y2=1.86
r80 37 43 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.43 $Y=1.86
+ $X2=4.565 $Y2=1.775
r81 37 38 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.43 $Y=1.86
+ $X2=3.815 $Y2=1.86
r82 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.72 $Y=1.98
+ $X2=3.72 $Y2=2.91
r83 31 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=1.945
+ $X2=3.72 $Y2=1.86
r84 31 33 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=3.72 $Y=1.945
+ $X2=3.72 $Y2=1.98
r85 27 41 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.745 $Y=1.065
+ $X2=3.745 $Y2=1.15
r86 27 29 30.9719 $w=2.38e-07 $l=6.45e-07 $layer=LI1_cond $X=3.745 $Y=1.065
+ $X2=3.745 $Y2=0.42
r87 25 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.625 $Y=1.86
+ $X2=3.72 $Y2=1.86
r88 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.625 $Y=1.86
+ $X2=2.955 $Y2=1.86
r89 23 41 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.625 $Y=1.15
+ $X2=3.745 $Y2=1.15
r90 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.625 $Y=1.15
+ $X2=2.955 $Y2=1.15
r91 19 24 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.865 $Y=1.065
+ $X2=2.955 $Y2=1.15
r92 19 21 39.7424 $w=1.78e-07 $l=6.45e-07 $layer=LI1_cond $X=2.865 $Y=1.065
+ $X2=2.865 $Y2=0.42
r93 15 17 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.86 $Y=1.98
+ $X2=2.86 $Y2=2.91
r94 13 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.86 $Y=1.945
+ $X2=2.955 $Y2=1.86
r95 13 15 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=2.86 $Y=1.945
+ $X2=2.86 $Y2=1.98
r96 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.835 $X2=3.72 $Y2=2.91
r97 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.835 $X2=3.72 $Y2=1.98
r98 3 17 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=2.91
r99 3 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=1.98
r100 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.58
+ $Y=0.235 $X2=3.72 $Y2=0.42
r101 1 21 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.72
+ $Y=0.235 $X2=2.86 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_4%VGND 1 2 3 12 16 18 22 25 26 27 28 29 43 44
+ 47
r57 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r58 44 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r59 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r60 41 47 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4.15
+ $Y2=0
r61 41 43 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4.56
+ $Y2=0
r62 40 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r63 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r64 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r65 33 37 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r66 32 36 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r67 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r68 29 40 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r69 29 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r70 27 39 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.12
+ $Y2=0
r71 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.29
+ $Y2=0
r72 25 36 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.16
+ $Y2=0
r73 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.345
+ $Y2=0
r74 24 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=3.12
+ $Y2=0
r75 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.345
+ $Y2=0
r76 20 47 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.15 $Y=0.085
+ $X2=4.15 $Y2=0
r77 20 22 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.15 $Y=0.085
+ $X2=4.15 $Y2=0.38
r78 19 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.29
+ $Y2=0
r79 18 47 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.035 $Y=0 $X2=4.15
+ $Y2=0
r80 18 19 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.035 $Y=0 $X2=3.455
+ $Y2=0
r81 14 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=0.085
+ $X2=3.29 $Y2=0
r82 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.29 $Y=0.085
+ $X2=3.29 $Y2=0.38
r83 10 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=0.085
+ $X2=2.345 $Y2=0
r84 10 12 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.345 $Y=0.085
+ $X2=2.345 $Y2=0.525
r85 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.01
+ $Y=0.235 $X2=4.15 $Y2=0.38
r86 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.15
+ $Y=0.235 $X2=3.29 $Y2=0.38
r87 1 12 182 $w=1.7e-07 $l=3.76962e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.235 $X2=2.345 $Y2=0.525
.ends

