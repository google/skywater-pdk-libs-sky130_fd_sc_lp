* File: sky130_fd_sc_lp__sdfrtp_2.pxi.spice
* Created: Fri Aug 28 11:28:28 2020
* 
x_PM_SKY130_FD_SC_LP__SDFRTP_2%A_35_74# N_A_35_74#_M1023_s N_A_35_74#_M1022_s
+ N_A_35_74#_c_283_n N_A_35_74#_M1003_g N_A_35_74#_M1018_g N_A_35_74#_c_284_n
+ N_A_35_74#_c_285_n N_A_35_74#_c_290_n N_A_35_74#_c_291_n N_A_35_74#_c_286_n
+ N_A_35_74#_c_292_n N_A_35_74#_c_287_n N_A_35_74#_c_288_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%A_35_74#
x_PM_SKY130_FD_SC_LP__SDFRTP_2%SCE N_SCE_M1023_g N_SCE_c_353_n N_SCE_c_359_n
+ N_SCE_c_360_n N_SCE_M1022_g N_SCE_c_362_n N_SCE_M1007_g N_SCE_M1039_g
+ N_SCE_c_364_n SCE SCE SCE SCE SCE N_SCE_c_356_n N_SCE_c_357_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%SCE
x_PM_SKY130_FD_SC_LP__SDFRTP_2%D N_D_M1033_g N_D_c_420_n N_D_M1032_g D D D D D
+ PM_SKY130_FD_SC_LP__SDFRTP_2%D
x_PM_SKY130_FD_SC_LP__SDFRTP_2%SCD N_SCD_c_455_n N_SCD_M1000_g N_SCD_M1012_g
+ N_SCD_c_460_n SCD SCD SCD N_SCD_c_458_n PM_SKY130_FD_SC_LP__SDFRTP_2%SCD
x_PM_SKY130_FD_SC_LP__SDFRTP_2%A_756_265# N_A_756_265#_M1006_s
+ N_A_756_265#_M1002_s N_A_756_265#_M1016_g N_A_756_265#_M1036_g
+ N_A_756_265#_c_501_n N_A_756_265#_M1015_g N_A_756_265#_c_502_n
+ N_A_756_265#_c_503_n N_A_756_265#_M1021_g N_A_756_265#_c_521_n
+ N_A_756_265#_c_504_n N_A_756_265#_c_505_n N_A_756_265#_c_506_n
+ N_A_756_265#_c_507_n N_A_756_265#_c_524_n N_A_756_265#_c_525_n
+ N_A_756_265#_c_508_n N_A_756_265#_c_509_n N_A_756_265#_c_510_n
+ N_A_756_265#_c_537_p N_A_756_265#_c_511_n N_A_756_265#_c_637_p
+ N_A_756_265#_c_512_n N_A_756_265#_c_513_n N_A_756_265#_c_514_n
+ N_A_756_265#_c_515_n N_A_756_265#_c_516_n N_A_756_265#_c_517_n
+ N_A_756_265#_c_518_n PM_SKY130_FD_SC_LP__SDFRTP_2%A_756_265#
x_PM_SKY130_FD_SC_LP__SDFRTP_2%A_936_333# N_A_936_333#_M1030_d
+ N_A_936_333#_M1025_d N_A_936_333#_M1004_g N_A_936_333#_c_711_n
+ N_A_936_333#_M1005_g N_A_936_333#_c_704_n N_A_936_333#_c_705_n
+ N_A_936_333#_c_706_n N_A_936_333#_c_707_n N_A_936_333#_c_714_n
+ N_A_936_333#_c_708_n N_A_936_333#_c_709_n N_A_936_333#_c_736_n
+ N_A_936_333#_c_717_n PM_SKY130_FD_SC_LP__SDFRTP_2%A_936_333#
x_PM_SKY130_FD_SC_LP__SDFRTP_2%RESET_B N_RESET_B_M1019_g N_RESET_B_c_803_n
+ N_RESET_B_c_804_n N_RESET_B_M1026_g N_RESET_B_c_806_n N_RESET_B_c_807_n
+ N_RESET_B_c_808_n N_RESET_B_c_809_n N_RESET_B_c_818_n N_RESET_B_M1013_g
+ N_RESET_B_c_819_n N_RESET_B_c_820_n N_RESET_B_M1037_g N_RESET_B_M1034_g
+ N_RESET_B_c_812_n N_RESET_B_c_813_n N_RESET_B_M1014_g N_RESET_B_c_814_n
+ N_RESET_B_c_815_n N_RESET_B_c_824_n N_RESET_B_c_881_p N_RESET_B_c_825_n
+ N_RESET_B_c_862_n N_RESET_B_c_826_n N_RESET_B_c_827_n RESET_B
+ N_RESET_B_c_828_n N_RESET_B_c_816_n N_RESET_B_c_830_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%RESET_B
x_PM_SKY130_FD_SC_LP__SDFRTP_2%A_808_463# N_A_808_463#_M1031_d
+ N_A_808_463#_M1016_d N_A_808_463#_M1013_d N_A_808_463#_c_1005_n
+ N_A_808_463#_M1030_g N_A_808_463#_M1025_g N_A_808_463#_c_1043_n
+ N_A_808_463#_c_1007_n N_A_808_463#_c_1013_n N_A_808_463#_c_1008_n
+ N_A_808_463#_c_1054_n N_A_808_463#_c_1009_n N_A_808_463#_c_1014_n
+ N_A_808_463#_c_1033_n N_A_808_463#_c_1010_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%A_808_463#
x_PM_SKY130_FD_SC_LP__SDFRTP_2%A_864_255# N_A_864_255#_M1008_d
+ N_A_864_255#_M1020_d N_A_864_255#_M1001_g N_A_864_255#_M1031_g
+ N_A_864_255#_c_1138_n N_A_864_255#_c_1139_n N_A_864_255#_M1009_g
+ N_A_864_255#_c_1126_n N_A_864_255#_c_1127_n N_A_864_255#_M1027_g
+ N_A_864_255#_M1006_g N_A_864_255#_M1002_g N_A_864_255#_c_1130_n
+ N_A_864_255#_c_1131_n N_A_864_255#_c_1132_n N_A_864_255#_c_1133_n
+ N_A_864_255#_c_1147_n N_A_864_255#_c_1148_n N_A_864_255#_c_1149_n
+ N_A_864_255#_c_1134_n N_A_864_255#_c_1150_n N_A_864_255#_c_1277_p
+ N_A_864_255#_c_1135_n N_A_864_255#_c_1136_n N_A_864_255#_c_1278_p
+ N_A_864_255#_c_1153_n PM_SKY130_FD_SC_LP__SDFRTP_2%A_864_255#
x_PM_SKY130_FD_SC_LP__SDFRTP_2%A_1406_69# N_A_1406_69#_M1015_d
+ N_A_1406_69#_M1009_d N_A_1406_69#_c_1322_n N_A_1406_69#_M1040_g
+ N_A_1406_69#_c_1323_n N_A_1406_69#_c_1324_n N_A_1406_69#_M1038_g
+ N_A_1406_69#_M1011_g N_A_1406_69#_M1028_g N_A_1406_69#_c_1328_n
+ N_A_1406_69#_c_1329_n N_A_1406_69#_c_1330_n N_A_1406_69#_c_1331_n
+ N_A_1406_69#_c_1332_n N_A_1406_69#_c_1333_n N_A_1406_69#_c_1346_n
+ N_A_1406_69#_c_1334_n N_A_1406_69#_c_1335_n N_A_1406_69#_c_1336_n
+ N_A_1406_69#_c_1337_n N_A_1406_69#_c_1338_n N_A_1406_69#_c_1339_n
+ N_A_1406_69#_c_1340_n N_A_1406_69#_c_1341_n N_A_1406_69#_c_1342_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%A_1406_69#
x_PM_SKY130_FD_SC_LP__SDFRTP_2%A_1635_21# N_A_1635_21#_M1040_d
+ N_A_1635_21#_M1014_d N_A_1635_21#_M1017_g N_A_1635_21#_M1035_g
+ N_A_1635_21#_c_1520_n N_A_1635_21#_c_1521_n N_A_1635_21#_c_1522_n
+ N_A_1635_21#_c_1523_n N_A_1635_21#_c_1524_n N_A_1635_21#_c_1531_n
+ N_A_1635_21#_c_1558_n N_A_1635_21#_c_1525_n N_A_1635_21#_c_1532_n
+ N_A_1635_21#_c_1526_n N_A_1635_21#_c_1527_n N_A_1635_21#_c_1533_n
+ N_A_1635_21#_c_1534_n N_A_1635_21#_c_1528_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%A_1635_21#
x_PM_SKY130_FD_SC_LP__SDFRTP_2%CLK N_CLK_M1008_g N_CLK_M1020_g N_CLK_c_1638_n
+ N_CLK_c_1639_n CLK CLK CLK N_CLK_c_1640_n N_CLK_c_1641_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%CLK
x_PM_SKY130_FD_SC_LP__SDFRTP_2%A_2431_47# N_A_2431_47#_M1011_s
+ N_A_2431_47#_M1028_s N_A_2431_47#_M1024_g N_A_2431_47#_M1010_g
+ N_A_2431_47#_M1041_g N_A_2431_47#_M1029_g N_A_2431_47#_c_1694_n
+ N_A_2431_47#_c_1702_n N_A_2431_47#_c_1695_n N_A_2431_47#_c_1696_n
+ N_A_2431_47#_c_1686_n N_A_2431_47#_c_1687_n N_A_2431_47#_c_1688_n
+ N_A_2431_47#_c_1689_n N_A_2431_47#_c_1690_n N_A_2431_47#_c_1691_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%A_2431_47#
x_PM_SKY130_FD_SC_LP__SDFRTP_2%VPWR N_VPWR_M1022_d N_VPWR_M1012_d N_VPWR_M1004_d
+ N_VPWR_M1025_s N_VPWR_M1035_d N_VPWR_M1038_d N_VPWR_M1002_d N_VPWR_M1028_d
+ N_VPWR_M1029_d N_VPWR_c_1771_n N_VPWR_c_1772_n N_VPWR_c_1773_n N_VPWR_c_1774_n
+ N_VPWR_c_1775_n N_VPWR_c_1776_n N_VPWR_c_1777_n N_VPWR_c_1778_n
+ N_VPWR_c_1779_n N_VPWR_c_1780_n N_VPWR_c_1781_n N_VPWR_c_1782_n
+ N_VPWR_c_1783_n N_VPWR_c_1784_n N_VPWR_c_1785_n VPWR N_VPWR_c_1786_n
+ N_VPWR_c_1787_n N_VPWR_c_1788_n N_VPWR_c_1789_n N_VPWR_c_1790_n
+ N_VPWR_c_1791_n N_VPWR_c_1792_n N_VPWR_c_1793_n N_VPWR_c_1794_n
+ N_VPWR_c_1795_n N_VPWR_c_1796_n N_VPWR_c_1770_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%VPWR
x_PM_SKY130_FD_SC_LP__SDFRTP_2%A_380_50# N_A_380_50#_M1033_d N_A_380_50#_M1031_s
+ N_A_380_50#_M1032_d N_A_380_50#_M1026_d N_A_380_50#_c_1931_n
+ N_A_380_50#_c_1937_n N_A_380_50#_c_1932_n N_A_380_50#_c_1933_n
+ N_A_380_50#_c_1934_n N_A_380_50#_c_1939_n N_A_380_50#_c_1935_n
+ N_A_380_50#_c_1940_n N_A_380_50#_c_1936_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%A_380_50#
x_PM_SKY130_FD_SC_LP__SDFRTP_2%Q N_Q_M1024_d N_Q_M1010_s N_Q_c_2038_n
+ N_Q_c_2039_n N_Q_c_2036_n N_Q_c_2035_n Q Q Q PM_SKY130_FD_SC_LP__SDFRTP_2%Q
x_PM_SKY130_FD_SC_LP__SDFRTP_2%VGND N_VGND_M1023_d N_VGND_M1019_d N_VGND_M1037_d
+ N_VGND_M1017_d N_VGND_M1006_d N_VGND_M1011_d N_VGND_M1041_s N_VGND_c_2061_n
+ N_VGND_c_2062_n N_VGND_c_2063_n N_VGND_c_2064_n N_VGND_c_2065_n
+ N_VGND_c_2066_n N_VGND_c_2067_n N_VGND_c_2068_n N_VGND_c_2069_n
+ N_VGND_c_2070_n N_VGND_c_2071_n N_VGND_c_2072_n N_VGND_c_2073_n
+ N_VGND_c_2074_n VGND N_VGND_c_2075_n N_VGND_c_2076_n N_VGND_c_2077_n
+ N_VGND_c_2078_n N_VGND_c_2079_n N_VGND_c_2080_n N_VGND_c_2081_n
+ N_VGND_c_2082_n PM_SKY130_FD_SC_LP__SDFRTP_2%VGND
x_PM_SKY130_FD_SC_LP__SDFRTP_2%noxref_24 N_noxref_24_M1003_s N_noxref_24_M1000_d
+ N_noxref_24_c_2204_n N_noxref_24_c_2205_n N_noxref_24_c_2206_n
+ PM_SKY130_FD_SC_LP__SDFRTP_2%noxref_24
cc_1 VNB N_A_35_74#_c_283_n 0.0212422f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.78
cc_2 VNB N_A_35_74#_c_284_n 0.0179504f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.58
cc_3 VNB N_A_35_74#_c_285_n 0.014408f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_4 VNB N_A_35_74#_c_286_n 0.00791735f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.945
cc_5 VNB N_A_35_74#_c_287_n 0.0326912f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.93
cc_6 VNB N_A_35_74#_c_288_n 0.0403563f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.945
cc_7 VNB N_SCE_M1023_g 0.0395444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_353_n 0.0337086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCE_M1039_g 0.0261313f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_10 VNB SCE 0.0336513f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.015
cc_11 VNB N_SCE_c_356_n 0.034328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_SCE_c_357_n 0.034075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D_M1033_g 0.0670496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_D_c_420_n 0.0223501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB D 0.0157732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCD_c_455_n 0.0165707f $X=-0.19 $Y=-0.245 $X2=0.175 $Y2=0.37
cc_17 VNB N_SCD_M1000_g 0.0265639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB SCD 0.00547455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_SCD_c_458_n 0.023828f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=0.945
cc_20 VNB N_A_756_265#_c_501_n 0.0216893f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.86
cc_21 VNB N_A_756_265#_c_502_n 0.0149208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_756_265#_c_503_n 0.0101942f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.03
cc_23 VNB N_A_756_265#_c_504_n 0.00298648f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.03
cc_24 VNB N_A_756_265#_c_505_n 0.0172381f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.015
cc_25 VNB N_A_756_265#_c_506_n 0.00611513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_756_265#_c_507_n 0.0032265f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.03
cc_27 VNB N_A_756_265#_c_508_n 0.0151454f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.945
cc_28 VNB N_A_756_265#_c_509_n 0.00147433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_756_265#_c_510_n 0.0153033f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.015
cc_30 VNB N_A_756_265#_c_511_n 0.00703168f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.18
cc_31 VNB N_A_756_265#_c_512_n 0.00642786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_756_265#_c_513_n 0.00256014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_756_265#_c_514_n 0.0285812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_756_265#_c_515_n 0.0289815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_756_265#_c_516_n 0.00636165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_756_265#_c_517_n 0.0158609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_756_265#_c_518_n 0.0330939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_936_333#_M1005_g 0.024004f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_39 VNB N_A_936_333#_c_704_n 0.0167487f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.03
cc_40 VNB N_A_936_333#_c_705_n 0.00885581f $X=-0.19 $Y=-0.245 $X2=0.405
+ $Y2=0.945
cc_41 VNB N_A_936_333#_c_706_n 0.0108991f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_42 VNB N_A_936_333#_c_707_n 0.0104872f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.03
cc_43 VNB N_A_936_333#_c_708_n 0.00193935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_936_333#_c_709_n 4.45643e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_M1019_g 0.00993309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_RESET_B_c_803_n 0.0235722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_804_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_RESET_B_M1026_g 0.0310576f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.46
cc_49 VNB N_RESET_B_c_806_n 0.0263834f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.66
cc_50 VNB N_RESET_B_c_807_n 0.0150584f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.66
cc_51 VNB N_RESET_B_c_808_n 0.0432014f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.86
cc_52 VNB N_RESET_B_c_809_n 0.149307f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_53 VNB N_RESET_B_M1037_g 0.0318232f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.015
cc_54 VNB N_RESET_B_M1034_g 0.0364663f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.945
cc_55 VNB N_RESET_B_c_812_n 0.0143436f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.93
cc_56 VNB N_RESET_B_c_813_n 0.00394614f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.485
cc_57 VNB N_RESET_B_c_814_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_c_815_n 0.00973448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_RESET_B_c_816_n 0.0224138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_808_463#_c_1005_n 0.0179652f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.18
cc_61 VNB N_A_808_463#_M1025_g 0.00110046f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_62 VNB N_A_808_463#_c_1007_n 0.00842474f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_63 VNB N_A_808_463#_c_1008_n 0.00375229f $X=-0.19 $Y=-0.245 $X2=1.035
+ $Y2=2.03
cc_64 VNB N_A_808_463#_c_1009_n 0.00396822f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=2.485
cc_65 VNB N_A_808_463#_c_1010_n 0.0747433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_864_255#_M1001_g 0.013419f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.18
cc_67 VNB N_A_864_255#_M1031_g 0.0248611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_864_255#_c_1126_n 0.0110246f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_69 VNB N_A_864_255#_c_1127_n 0.00316727f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_70 VNB N_A_864_255#_M1027_g 0.0440125f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.03
cc_71 VNB N_A_864_255#_M1006_g 0.02239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_864_255#_c_1130_n 0.0113368f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_73 VNB N_A_864_255#_c_1131_n 0.00384825f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=0.945
cc_74 VNB N_A_864_255#_c_1132_n 0.00800365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_864_255#_c_1133_n 0.0012281f $X=-0.19 $Y=-0.245 $X2=2.395
+ $Y2=2.015
cc_76 VNB N_A_864_255#_c_1134_n 0.0157205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_864_255#_c_1135_n 0.0139559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_864_255#_c_1136_n 0.0294614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1406_69#_c_1322_n 0.0160964f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.78
cc_80 VNB N_A_1406_69#_c_1323_n 0.0138651f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.18
cc_81 VNB N_A_1406_69#_c_1324_n 0.00620811f $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.66
cc_82 VNB N_A_1406_69#_M1038_g 0.0094489f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.86
cc_83 VNB N_A_1406_69#_M1011_g 0.0258606f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.03
cc_84 VNB N_A_1406_69#_M1028_g 0.00429678f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_85 VNB N_A_1406_69#_c_1328_n 0.0209677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1406_69#_c_1329_n 0.0178053f $X=-0.19 $Y=-0.245 $X2=2.395
+ $Y2=2.015
cc_87 VNB N_A_1406_69#_c_1330_n 0.00119189f $X=-0.19 $Y=-0.245 $X2=2.395
+ $Y2=2.015
cc_88 VNB N_A_1406_69#_c_1331_n 0.00696254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1406_69#_c_1332_n 0.0112643f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.945
cc_90 VNB N_A_1406_69#_c_1333_n 0.00247664f $X=-0.19 $Y=-0.245 $X2=0.94
+ $Y2=2.485
cc_91 VNB N_A_1406_69#_c_1334_n 0.00163504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1406_69#_c_1335_n 0.0213833f $X=-0.19 $Y=-0.245 $X2=2.395
+ $Y2=2.015
cc_93 VNB N_A_1406_69#_c_1336_n 0.00170636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1406_69#_c_1337_n 0.00800408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1406_69#_c_1338_n 0.0216293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1406_69#_c_1339_n 0.00313421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1406_69#_c_1340_n 0.023598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1406_69#_c_1341_n 0.0308494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1406_69#_c_1342_n 0.0428435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1635_21#_M1017_g 0.0219387f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.18
cc_101 VNB N_A_1635_21#_c_1520_n 0.109613f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_102 VNB N_A_1635_21#_c_1521_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.58
cc_103 VNB N_A_1635_21#_c_1522_n 0.0260034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1635_21#_c_1523_n 0.00606018f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.03
cc_105 VNB N_A_1635_21#_c_1524_n 0.0188331f $X=-0.19 $Y=-0.245 $X2=0.405
+ $Y2=0.945
cc_106 VNB N_A_1635_21#_c_1525_n 0.00337432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1635_21#_c_1526_n 0.00372955f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=2.485
cc_108 VNB N_A_1635_21#_c_1527_n 0.00607331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1635_21#_c_1528_n 0.0522379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_CLK_M1008_g 0.0244479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_CLK_M1020_g 0.00586985f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.78
cc_112 VNB N_CLK_c_1638_n 0.0182093f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.46
cc_113 VNB N_CLK_c_1639_n 0.00391068f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.66
cc_114 VNB N_CLK_c_1640_n 0.0262869f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.03
cc_115 VNB N_CLK_c_1641_n 0.00368549f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_116 VNB N_A_2431_47#_M1024_g 0.0192472f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.46
cc_117 VNB N_A_2431_47#_M1010_g 0.00431392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2431_47#_M1041_g 0.0256705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2431_47#_M1029_g 0.00602717f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_120 VNB N_A_2431_47#_c_1686_n 0.00377889f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=2.03
cc_121 VNB N_A_2431_47#_c_1687_n 0.00245565f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.93
cc_122 VNB N_A_2431_47#_c_1688_n 0.00102726f $X=-0.19 $Y=-0.245 $X2=0.94
+ $Y2=2.485
cc_123 VNB N_A_2431_47#_c_1689_n 0.00426398f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_124 VNB N_A_2431_47#_c_1690_n 0.00418217f $X=-0.19 $Y=-0.245 $X2=2.395
+ $Y2=2.015
cc_125 VNB N_A_2431_47#_c_1691_n 0.0611355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VPWR_c_1770_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_380_50#_c_1931_n 0.013305f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_128 VNB N_A_380_50#_c_1932_n 0.00426068f $X=-0.19 $Y=-0.245 $X2=0.405
+ $Y2=0.945
cc_129 VNB N_A_380_50#_c_1933_n 0.00225068f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_130 VNB N_A_380_50#_c_1934_n 0.00810127f $X=-0.19 $Y=-0.245 $X2=2.395
+ $Y2=2.03
cc_131 VNB N_A_380_50#_c_1935_n 0.00162082f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.93
cc_132 VNB N_A_380_50#_c_1936_n 0.00284405f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_133 VNB N_Q_c_2035_n 0.00171756f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_134 VNB N_VGND_c_2061_n 0.00993588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2062_n 0.00889572f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.015
cc_136 VNB N_VGND_c_2063_n 0.00864254f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.93
cc_137 VNB N_VGND_c_2064_n 0.0109665f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_138 VNB N_VGND_c_2065_n 0.00864305f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.015
cc_139 VNB N_VGND_c_2066_n 0.00276358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2067_n 0.0107404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2068_n 0.0481093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2069_n 0.0726178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2070_n 0.00594344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2071_n 0.0504328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2072_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2073_n 0.0546665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2074_n 0.00631504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2075_n 0.0181906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2076_n 0.0590578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2077_n 0.0371839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2078_n 0.0154348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2079_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2080_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2081_n 0.00516105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2082_n 0.682965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_noxref_24_c_2204_n 0.00432969f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=0.78
cc_157 VNB N_noxref_24_c_2205_n 0.00390834f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=0.46
cc_158 VNB N_noxref_24_c_2206_n 0.00236766f $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=0.86
cc_159 VPB N_A_35_74#_M1018_g 0.0203099f $X=-0.19 $Y=1.655 $X2=2.375 $Y2=2.66
cc_160 VPB N_A_35_74#_c_290_n 0.0200503f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=2.015
cc_161 VPB N_A_35_74#_c_291_n 0.0319044f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=2.015
cc_162 VPB N_A_35_74#_c_292_n 0.0729262f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.03
cc_163 VPB N_A_35_74#_c_287_n 0.0139259f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.93
cc_164 VPB N_SCE_c_353_n 0.0462946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_SCE_c_359_n 0.0127327f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.78
cc_166 VPB N_SCE_c_360_n 0.0253985f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.46
cc_167 VPB N_SCE_M1022_g 0.0209361f $X=-0.19 $Y=1.655 $X2=2.375 $Y2=2.66
cc_168 VPB N_SCE_c_362_n 0.0232878f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_SCE_M1007_g 0.0177003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_SCE_c_364_n 0.00666874f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_171 VPB N_D_c_420_n 0.0244722f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_D_M1032_g 0.0410389f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.78
cc_173 VPB D 0.0152853f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_SCD_M1012_g 0.0320543f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.78
cc_175 VPB N_SCD_c_460_n 0.018347f $X=-0.19 $Y=1.655 $X2=2.375 $Y2=2.66
cc_176 VPB SCD 0.00622066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_SCD_c_458_n 0.0153015f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=0.945
cc_178 VPB N_A_756_265#_M1016_g 0.0301572f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.46
cc_179 VPB N_A_756_265#_M1021_g 0.0266706f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_180 VPB N_A_756_265#_c_521_n 0.0156771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_756_265#_c_504_n 0.00516087f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=2.03
cc_182 VPB N_A_756_265#_c_506_n 0.00794753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_756_265#_c_524_n 0.00259066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_756_265#_c_525_n 0.0372553f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_185 VPB N_A_756_265#_c_512_n 0.00475318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_756_265#_c_514_n 0.0111211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_936_333#_M1004_g 0.0269928f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.46
cc_188 VPB N_A_936_333#_c_711_n 0.025819f $X=-0.19 $Y=1.655 $X2=2.375 $Y2=2.66
cc_189 VPB N_A_936_333#_c_704_n 0.00186275f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.03
cc_190 VPB N_A_936_333#_c_706_n 0.0127244f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_191 VPB N_A_936_333#_c_714_n 0.00103499f $X=-0.19 $Y=1.655 $X2=2.395
+ $Y2=2.015
cc_192 VPB N_A_936_333#_c_708_n 0.00178195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_936_333#_c_709_n 7.29702e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_936_333#_c_717_n 0.0350077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_RESET_B_M1026_g 0.0495042f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.46
cc_196 VPB N_RESET_B_c_818_n 0.019097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_RESET_B_c_819_n 0.0216981f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=0.945
cc_198 VPB N_RESET_B_c_820_n 0.0083369f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_199 VPB N_RESET_B_c_812_n 0.00497343f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.93
cc_200 VPB N_RESET_B_c_813_n 0.00454165f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.485
cc_201 VPB N_RESET_B_M1014_g 0.0225139f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_202 VPB N_RESET_B_c_824_n 0.00351546f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_RESET_B_c_825_n 0.0161988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_RESET_B_c_826_n 0.0016088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_RESET_B_c_827_n 0.0354135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_RESET_B_c_828_n 0.0764971f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_816_n 0.0156389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_RESET_B_c_830_n 0.026967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_808_463#_M1025_g 0.0255057f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=0.58
cc_210 VPB N_A_808_463#_c_1007_n 0.00371024f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_211 VPB N_A_808_463#_c_1013_n 0.00804597f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_212 VPB N_A_808_463#_c_1014_n 0.00699661f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_213 VPB N_A_864_255#_M1001_g 0.0513431f $X=-0.19 $Y=1.655 $X2=2.375 $Y2=2.18
cc_214 VPB N_A_864_255#_c_1138_n 0.204793f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=0.58
cc_215 VPB N_A_864_255#_c_1139_n 0.012806f $X=-0.19 $Y=1.655 $X2=0.3 $Y2=0.58
cc_216 VPB N_A_864_255#_M1009_g 0.0291f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=0.945
cc_217 VPB N_A_864_255#_c_1126_n 0.0268847f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_218 VPB N_A_864_255#_c_1127_n 0.00381747f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_219 VPB N_A_864_255#_M1002_g 0.0226368f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.485
cc_220 VPB N_A_864_255#_c_1131_n 0.00787526f $X=-0.19 $Y=1.655 $X2=1.465
+ $Y2=0.945
cc_221 VPB N_A_864_255#_c_1132_n 0.0156721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_864_255#_c_1133_n 0.00558761f $X=-0.19 $Y=1.655 $X2=2.395
+ $Y2=2.015
cc_223 VPB N_A_864_255#_c_1147_n 0.01386f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=2.18
cc_224 VPB N_A_864_255#_c_1148_n 0.0163242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_864_255#_c_1149_n 0.00375656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_864_255#_c_1150_n 0.00151381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_864_255#_c_1135_n 0.0193117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_864_255#_c_1136_n 0.00806119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_864_255#_c_1153_n 0.0118506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_1406_69#_M1038_g 0.06887f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=0.86
cc_231 VPB N_A_1406_69#_M1028_g 0.0258827f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_232 VPB N_A_1406_69#_c_1333_n 0.00135887f $X=-0.19 $Y=1.655 $X2=0.94
+ $Y2=2.485
cc_233 VPB N_A_1406_69#_c_1346_n 0.00161251f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_234 VPB N_A_1635_21#_M1035_g 0.0386939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_1635_21#_c_1524_n 0.0170452f $X=-0.19 $Y=1.655 $X2=0.405
+ $Y2=0.945
cc_236 VPB N_A_1635_21#_c_1531_n 0.0142536f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_237 VPB N_A_1635_21#_c_1532_n 0.00424123f $X=-0.19 $Y=1.655 $X2=0.585
+ $Y2=1.93
cc_238 VPB N_A_1635_21#_c_1533_n 0.00518188f $X=-0.19 $Y=1.655 $X2=1.465
+ $Y2=0.945
cc_239 VPB N_A_1635_21#_c_1534_n 0.0509975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_CLK_M1020_g 0.024773f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.78
cc_241 VPB N_CLK_c_1640_n 0.0106975f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.03
cc_242 VPB N_CLK_c_1641_n 0.0207771f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_243 VPB N_A_2431_47#_M1010_g 0.022325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_2431_47#_M1029_g 0.0264965f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_245 VPB N_A_2431_47#_c_1694_n 0.00458841f $X=-0.19 $Y=1.655 $X2=1.035
+ $Y2=2.03
cc_246 VPB N_A_2431_47#_c_1695_n 0.00537492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_2431_47#_c_1696_n 0.00333047f $X=-0.19 $Y=1.655 $X2=0.27
+ $Y2=0.945
cc_248 VPB N_A_2431_47#_c_1690_n 0.00183434f $X=-0.19 $Y=1.655 $X2=2.395
+ $Y2=2.015
cc_249 VPB N_VPWR_c_1771_n 0.00760603f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.945
cc_250 VPB N_VPWR_c_1772_n 0.00964855f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.485
cc_251 VPB N_VPWR_c_1773_n 0.0153711f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.945
cc_252 VPB N_VPWR_c_1774_n 0.0207158f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=2.18
cc_253 VPB N_VPWR_c_1775_n 0.00950882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1776_n 0.00268089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1777_n 0.02302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1778_n 0.0107145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1779_n 0.0639877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1780_n 0.0329037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1781_n 0.00482629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1782_n 0.0197332f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1783_n 0.0047802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1784_n 0.0189374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1785_n 0.00481989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1786_n 0.0448455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1787_n 0.0440347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1788_n 0.030381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1789_n 0.042172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1790_n 0.0154348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1791_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1792_n 0.00435574f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1793_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1794_n 0.0489093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1795_n 0.0180895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1796_n 0.00651403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1770_n 0.107685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_380_50#_c_1937_n 0.0100215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_A_380_50#_c_1932_n 0.00484411f $X=-0.19 $Y=1.655 $X2=0.405
+ $Y2=0.945
cc_278 VPB N_A_380_50#_c_1939_n 0.00471706f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.03
cc_279 VPB N_A_380_50#_c_1940_n 0.0122559f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.485
cc_280 VPB N_Q_c_2036_n 0.00323231f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=0.86
cc_281 VPB N_Q_c_2035_n 7.12541e-19 $X=-0.19 $Y=1.655 $X2=0.265 $Y2=0.58
cc_282 N_A_35_74#_c_284_n N_SCE_M1023_g 0.00313661f $X=0.3 $Y=0.58 $X2=0 $Y2=0
cc_283 N_A_35_74#_c_285_n N_SCE_M1023_g 0.0184567f $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_284 N_A_35_74#_c_287_n N_SCE_M1023_g 0.0349739f $X=0.585 $Y=1.93 $X2=0 $Y2=0
cc_285 N_A_35_74#_c_288_n N_SCE_M1023_g 0.00681185f $X=1.465 $Y=0.945 $X2=0
+ $Y2=0
cc_286 N_A_35_74#_c_290_n N_SCE_c_353_n 7.56281e-19 $X=2.395 $Y=2.015 $X2=0
+ $Y2=0
cc_287 N_A_35_74#_c_292_n N_SCE_c_353_n 0.0224464f $X=0.585 $Y=2.03 $X2=0 $Y2=0
cc_288 N_A_35_74#_c_290_n N_SCE_c_359_n 0.00293037f $X=2.395 $Y=2.015 $X2=0
+ $Y2=0
cc_289 N_A_35_74#_c_292_n N_SCE_c_359_n 0.0107508f $X=0.585 $Y=2.03 $X2=0 $Y2=0
cc_290 N_A_35_74#_c_292_n N_SCE_c_360_n 0.0216778f $X=0.585 $Y=2.03 $X2=0 $Y2=0
cc_291 N_A_35_74#_c_292_n N_SCE_M1022_g 0.00608296f $X=0.585 $Y=2.03 $X2=0 $Y2=0
cc_292 N_A_35_74#_c_290_n N_SCE_c_362_n 0.0218464f $X=2.395 $Y=2.015 $X2=0 $Y2=0
cc_293 N_A_35_74#_c_290_n N_SCE_c_364_n 0.00953865f $X=2.395 $Y=2.015 $X2=0
+ $Y2=0
cc_294 N_A_35_74#_c_285_n SCE 0.0681126f $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_295 N_A_35_74#_c_287_n SCE 0.0146701f $X=0.585 $Y=1.93 $X2=0 $Y2=0
cc_296 N_A_35_74#_c_288_n SCE 0.0100266f $X=1.465 $Y=0.945 $X2=0 $Y2=0
cc_297 N_A_35_74#_c_285_n N_SCE_c_356_n 0.0092968f $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_298 N_A_35_74#_c_291_n N_SCE_c_357_n 0.00845332f $X=2.395 $Y=2.015 $X2=0
+ $Y2=0
cc_299 N_A_35_74#_c_283_n N_D_M1033_g 0.0635766f $X=1.465 $Y=0.78 $X2=0 $Y2=0
cc_300 N_A_35_74#_c_285_n N_D_M1033_g 6.37375e-19 $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_301 N_A_35_74#_c_290_n N_D_c_420_n 0.00557826f $X=2.395 $Y=2.015 $X2=0 $Y2=0
cc_302 N_A_35_74#_M1018_g N_D_M1032_g 0.0143482f $X=2.375 $Y=2.66 $X2=0 $Y2=0
cc_303 N_A_35_74#_c_290_n N_D_M1032_g 0.0163411f $X=2.395 $Y=2.015 $X2=0 $Y2=0
cc_304 N_A_35_74#_c_291_n N_D_M1032_g 0.0220528f $X=2.395 $Y=2.015 $X2=0 $Y2=0
cc_305 N_A_35_74#_c_290_n D 0.114889f $X=2.395 $Y=2.015 $X2=0 $Y2=0
cc_306 N_A_35_74#_c_291_n D 0.00313801f $X=2.395 $Y=2.015 $X2=0 $Y2=0
cc_307 N_A_35_74#_c_292_n D 0.036479f $X=0.585 $Y=2.03 $X2=0 $Y2=0
cc_308 N_A_35_74#_c_287_n D 0.0171918f $X=0.585 $Y=1.93 $X2=0 $Y2=0
cc_309 N_A_35_74#_M1018_g N_SCD_M1012_g 0.035782f $X=2.375 $Y=2.66 $X2=0 $Y2=0
cc_310 N_A_35_74#_c_290_n N_SCD_c_460_n 6.98602e-19 $X=2.395 $Y=2.015 $X2=0
+ $Y2=0
cc_311 N_A_35_74#_c_291_n N_SCD_c_460_n 0.0212646f $X=2.395 $Y=2.015 $X2=0 $Y2=0
cc_312 N_A_35_74#_c_290_n SCD 0.00900903f $X=2.395 $Y=2.015 $X2=0 $Y2=0
cc_313 N_A_35_74#_c_291_n SCD 6.31533e-19 $X=2.395 $Y=2.015 $X2=0 $Y2=0
cc_314 N_A_35_74#_c_290_n N_VPWR_c_1771_n 0.0199655f $X=2.395 $Y=2.015 $X2=0
+ $Y2=0
cc_315 N_A_35_74#_c_292_n N_VPWR_c_1771_n 0.0265069f $X=0.585 $Y=2.03 $X2=0
+ $Y2=0
cc_316 N_A_35_74#_c_292_n N_VPWR_c_1780_n 0.0435581f $X=0.585 $Y=2.03 $X2=0
+ $Y2=0
cc_317 N_A_35_74#_M1018_g N_VPWR_c_1786_n 0.00449508f $X=2.375 $Y=2.66 $X2=0
+ $Y2=0
cc_318 N_A_35_74#_M1018_g N_VPWR_c_1770_n 0.00488839f $X=2.375 $Y=2.66 $X2=0
+ $Y2=0
cc_319 N_A_35_74#_c_292_n N_VPWR_c_1770_n 0.0335596f $X=0.585 $Y=2.03 $X2=0
+ $Y2=0
cc_320 N_A_35_74#_M1018_g N_A_380_50#_c_1937_n 0.00877292f $X=2.375 $Y=2.66
+ $X2=0 $Y2=0
cc_321 N_A_35_74#_c_290_n N_A_380_50#_c_1937_n 0.0165074f $X=2.395 $Y=2.015
+ $X2=0 $Y2=0
cc_322 N_A_35_74#_c_291_n N_A_380_50#_c_1937_n 0.00261593f $X=2.395 $Y=2.015
+ $X2=0 $Y2=0
cc_323 N_A_35_74#_c_285_n N_A_380_50#_c_1934_n 0.00550184f $X=1.345 $Y=0.945
+ $X2=0 $Y2=0
cc_324 N_A_35_74#_M1018_g N_A_380_50#_c_1939_n 0.0118252f $X=2.375 $Y=2.66 $X2=0
+ $Y2=0
cc_325 N_A_35_74#_c_290_n N_A_380_50#_c_1939_n 0.0275609f $X=2.395 $Y=2.015
+ $X2=0 $Y2=0
cc_326 N_A_35_74#_c_291_n N_A_380_50#_c_1939_n 0.00173089f $X=2.395 $Y=2.015
+ $X2=0 $Y2=0
cc_327 N_A_35_74#_c_283_n N_VGND_c_2061_n 0.00386287f $X=1.465 $Y=0.78 $X2=0
+ $Y2=0
cc_328 N_A_35_74#_c_285_n N_VGND_c_2061_n 0.0238773f $X=1.345 $Y=0.945 $X2=0
+ $Y2=0
cc_329 N_A_35_74#_c_284_n N_VGND_c_2075_n 0.00870147f $X=0.3 $Y=0.58 $X2=0 $Y2=0
cc_330 N_A_35_74#_c_283_n N_VGND_c_2076_n 0.00351389f $X=1.465 $Y=0.78 $X2=0
+ $Y2=0
cc_331 N_A_35_74#_c_283_n N_VGND_c_2082_n 0.0063493f $X=1.465 $Y=0.78 $X2=0
+ $Y2=0
cc_332 N_A_35_74#_c_284_n N_VGND_c_2082_n 0.00914631f $X=0.3 $Y=0.58 $X2=0 $Y2=0
cc_333 N_A_35_74#_c_285_n N_VGND_c_2082_n 0.0128604f $X=1.345 $Y=0.945 $X2=0
+ $Y2=0
cc_334 N_A_35_74#_c_286_n N_VGND_c_2082_n 3.87486e-19 $X=0.27 $Y=0.945 $X2=0
+ $Y2=0
cc_335 N_A_35_74#_c_283_n N_noxref_24_c_2204_n 0.00854136f $X=1.465 $Y=0.78
+ $X2=0 $Y2=0
cc_336 N_A_35_74#_c_285_n N_noxref_24_c_2204_n 0.00262689f $X=1.345 $Y=0.945
+ $X2=0 $Y2=0
cc_337 N_A_35_74#_c_283_n N_noxref_24_c_2205_n 0.00476417f $X=1.465 $Y=0.78
+ $X2=0 $Y2=0
cc_338 N_A_35_74#_c_285_n N_noxref_24_c_2205_n 0.0166978f $X=1.345 $Y=0.945
+ $X2=0 $Y2=0
cc_339 N_A_35_74#_c_288_n N_noxref_24_c_2205_n 0.00487372f $X=1.465 $Y=0.945
+ $X2=0 $Y2=0
cc_340 N_SCE_M1039_g N_D_M1033_g 0.0176354f $X=2.485 $Y=0.615 $X2=0 $Y2=0
cc_341 SCE N_D_M1033_g 0.0179101f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_342 N_SCE_c_357_n N_D_M1033_g 0.013574f $X=2.395 $Y=1.295 $X2=0 $Y2=0
cc_343 SCE N_D_c_420_n 0.00487125f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_344 N_SCE_c_362_n N_D_M1032_g 0.063563f $X=1.51 $Y=2.135 $X2=0 $Y2=0
cc_345 N_SCE_c_353_n D 0.0230165f $X=0.677 $Y=2.06 $X2=0 $Y2=0
cc_346 N_SCE_c_359_n D 0.00382924f $X=1.08 $Y=2.135 $X2=0 $Y2=0
cc_347 SCE D 0.160301f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_348 N_SCE_c_357_n D 0.00313801f $X=2.395 $Y=1.295 $X2=0 $Y2=0
cc_349 SCE N_SCD_c_455_n 0.00125075f $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_350 N_SCE_c_357_n N_SCD_c_455_n 0.0334662f $X=2.395 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_351 N_SCE_M1039_g N_SCD_M1000_g 0.0334662f $X=2.485 $Y=0.615 $X2=0 $Y2=0
cc_352 SCE SCD 0.0143507f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_353 N_SCE_c_357_n SCD 5.97719e-19 $X=2.395 $Y=1.295 $X2=0 $Y2=0
cc_354 SCE N_SCD_c_458_n 3.50187e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_355 N_SCE_c_357_n N_SCD_c_458_n 0.00635576f $X=2.395 $Y=1.295 $X2=0 $Y2=0
cc_356 N_SCE_M1022_g N_VPWR_c_1771_n 0.0136472f $X=1.155 $Y=2.66 $X2=0 $Y2=0
cc_357 N_SCE_c_362_n N_VPWR_c_1771_n 0.00218665f $X=1.51 $Y=2.135 $X2=0 $Y2=0
cc_358 N_SCE_M1007_g N_VPWR_c_1771_n 0.00332228f $X=1.585 $Y=2.66 $X2=0 $Y2=0
cc_359 N_SCE_M1022_g N_VPWR_c_1780_n 0.00396895f $X=1.155 $Y=2.66 $X2=0 $Y2=0
cc_360 N_SCE_M1007_g N_VPWR_c_1786_n 0.00478016f $X=1.585 $Y=2.66 $X2=0 $Y2=0
cc_361 N_SCE_M1022_g N_VPWR_c_1770_n 0.00796233f $X=1.155 $Y=2.66 $X2=0 $Y2=0
cc_362 N_SCE_M1007_g N_VPWR_c_1770_n 0.00935327f $X=1.585 $Y=2.66 $X2=0 $Y2=0
cc_363 N_SCE_M1039_g N_A_380_50#_c_1931_n 0.011034f $X=2.485 $Y=0.615 $X2=0
+ $Y2=0
cc_364 SCE N_A_380_50#_c_1931_n 0.0270001f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_365 N_SCE_c_357_n N_A_380_50#_c_1931_n 0.00215661f $X=2.395 $Y=1.295 $X2=0
+ $Y2=0
cc_366 N_SCE_M1039_g N_A_380_50#_c_1934_n 0.00620309f $X=2.485 $Y=0.615 $X2=0
+ $Y2=0
cc_367 SCE N_A_380_50#_c_1934_n 0.0238303f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_368 N_SCE_c_357_n N_A_380_50#_c_1934_n 0.00218697f $X=2.395 $Y=1.295 $X2=0
+ $Y2=0
cc_369 N_SCE_M1007_g N_A_380_50#_c_1939_n 0.00200928f $X=1.585 $Y=2.66 $X2=0
+ $Y2=0
cc_370 N_SCE_M1023_g N_VGND_c_2061_n 0.0138465f $X=0.515 $Y=0.58 $X2=0 $Y2=0
cc_371 N_SCE_M1023_g N_VGND_c_2075_n 0.00383152f $X=0.515 $Y=0.58 $X2=0 $Y2=0
cc_372 N_SCE_M1039_g N_VGND_c_2076_n 9.29198e-19 $X=2.485 $Y=0.615 $X2=0 $Y2=0
cc_373 N_SCE_M1023_g N_VGND_c_2082_n 0.0039187f $X=0.515 $Y=0.58 $X2=0 $Y2=0
cc_374 N_SCE_M1039_g N_noxref_24_c_2204_n 0.0118723f $X=2.485 $Y=0.615 $X2=0
+ $Y2=0
cc_375 N_SCE_M1023_g N_noxref_24_c_2205_n 8.06104e-19 $X=0.515 $Y=0.58 $X2=0
+ $Y2=0
cc_376 N_SCE_M1039_g N_noxref_24_c_2206_n 0.00109906f $X=2.485 $Y=0.615 $X2=0
+ $Y2=0
cc_377 D SCD 0.0177105f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_378 D N_SCD_c_458_n 0.00534059f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_379 N_D_M1032_g N_VPWR_c_1786_n 0.00449508f $X=1.945 $Y=2.66 $X2=0 $Y2=0
cc_380 N_D_M1032_g N_VPWR_c_1770_n 0.00854629f $X=1.945 $Y=2.66 $X2=0 $Y2=0
cc_381 D N_A_380_50#_c_1937_n 0.00601221f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_382 N_D_M1033_g N_A_380_50#_c_1934_n 0.00904098f $X=1.825 $Y=0.46 $X2=0 $Y2=0
cc_383 N_D_M1032_g N_A_380_50#_c_1939_n 0.0131282f $X=1.945 $Y=2.66 $X2=0 $Y2=0
cc_384 N_D_M1033_g N_VGND_c_2076_n 0.00349953f $X=1.825 $Y=0.46 $X2=0 $Y2=0
cc_385 N_D_M1033_g N_VGND_c_2082_n 0.00635843f $X=1.825 $Y=0.46 $X2=0 $Y2=0
cc_386 N_D_M1033_g N_noxref_24_c_2204_n 0.0148629f $X=1.825 $Y=0.46 $X2=0 $Y2=0
cc_387 N_D_M1033_g N_noxref_24_c_2205_n 9.87143e-19 $X=1.825 $Y=0.46 $X2=0 $Y2=0
cc_388 N_SCD_M1000_g N_RESET_B_M1019_g 0.0211242f $X=2.845 $Y=0.615 $X2=0 $Y2=0
cc_389 N_SCD_c_455_n N_RESET_B_M1026_g 0.0428382f $X=2.845 $Y=1.185 $X2=0 $Y2=0
cc_390 N_SCD_M1000_g N_RESET_B_M1026_g 0.00278588f $X=2.845 $Y=0.615 $X2=0 $Y2=0
cc_391 N_SCD_M1012_g N_RESET_B_M1026_g 0.0240943f $X=2.845 $Y=2.66 $X2=0 $Y2=0
cc_392 SCD N_RESET_B_M1026_g 0.00640013f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_393 SCD N_RESET_B_c_807_n 0.00202629f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_394 N_SCD_M1012_g N_VPWR_c_1772_n 0.00582729f $X=2.845 $Y=2.66 $X2=0 $Y2=0
cc_395 N_SCD_M1012_g N_VPWR_c_1786_n 0.00478016f $X=2.845 $Y=2.66 $X2=0 $Y2=0
cc_396 N_SCD_M1012_g N_VPWR_c_1770_n 0.00527534f $X=2.845 $Y=2.66 $X2=0 $Y2=0
cc_397 N_SCD_c_455_n N_A_380_50#_c_1931_n 0.00237845f $X=2.845 $Y=1.185 $X2=0
+ $Y2=0
cc_398 N_SCD_M1000_g N_A_380_50#_c_1931_n 0.014929f $X=2.845 $Y=0.615 $X2=0
+ $Y2=0
cc_399 SCD N_A_380_50#_c_1931_n 0.0273322f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_400 N_SCD_M1012_g N_A_380_50#_c_1937_n 0.0169075f $X=2.845 $Y=2.66 $X2=0
+ $Y2=0
cc_401 N_SCD_c_460_n N_A_380_50#_c_1937_n 0.00116918f $X=2.962 $Y=1.995 $X2=0
+ $Y2=0
cc_402 SCD N_A_380_50#_c_1937_n 0.0318088f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_403 N_SCD_c_455_n N_A_380_50#_c_1932_n 7.81287e-19 $X=2.845 $Y=1.185 $X2=0
+ $Y2=0
cc_404 N_SCD_M1000_g N_A_380_50#_c_1932_n 7.90567e-19 $X=2.845 $Y=0.615 $X2=0
+ $Y2=0
cc_405 N_SCD_M1012_g N_A_380_50#_c_1932_n 9.06689e-19 $X=2.845 $Y=2.66 $X2=0
+ $Y2=0
cc_406 SCD N_A_380_50#_c_1932_n 0.0716565f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_407 N_SCD_M1012_g N_A_380_50#_c_1939_n 0.00193047f $X=2.845 $Y=2.66 $X2=0
+ $Y2=0
cc_408 N_SCD_M1012_g N_A_380_50#_c_1940_n 8.09944e-19 $X=2.845 $Y=2.66 $X2=0
+ $Y2=0
cc_409 N_SCD_M1000_g N_VGND_c_2076_n 9.22791e-19 $X=2.845 $Y=0.615 $X2=0 $Y2=0
cc_410 N_SCD_M1000_g N_noxref_24_c_2204_n 0.00824966f $X=2.845 $Y=0.615 $X2=0
+ $Y2=0
cc_411 N_SCD_M1000_g N_noxref_24_c_2206_n 0.00708705f $X=2.845 $Y=0.615 $X2=0
+ $Y2=0
cc_412 N_A_756_265#_c_515_n N_A_936_333#_c_711_n 0.00284672f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_413 N_A_756_265#_c_516_n N_A_936_333#_c_711_n 8.37161e-19 $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_414 N_A_756_265#_c_510_n N_A_936_333#_M1005_g 0.00230372f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_415 N_A_756_265#_c_515_n N_A_936_333#_M1005_g 0.0192524f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_416 N_A_756_265#_c_516_n N_A_936_333#_M1005_g 0.00620794f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_417 N_A_756_265#_c_517_n N_A_936_333#_M1005_g 0.027489f $X=4.9 $Y=1.125 $X2=0
+ $Y2=0
cc_418 N_A_756_265#_c_515_n N_A_936_333#_c_704_n 0.00181244f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_419 N_A_756_265#_c_510_n N_A_936_333#_c_705_n 0.00349273f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_420 N_A_756_265#_c_510_n N_A_936_333#_c_706_n 0.0339737f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_421 N_A_756_265#_c_537_p N_A_936_333#_c_706_n 0.00126513f $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_422 N_A_756_265#_c_515_n N_A_936_333#_c_706_n 3.27937e-19 $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_423 N_A_756_265#_c_516_n N_A_936_333#_c_706_n 0.013295f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_424 N_A_756_265#_c_501_n N_A_936_333#_c_707_n 0.00224374f $X=6.955 $Y=1.095
+ $X2=0 $Y2=0
cc_425 N_A_756_265#_c_510_n N_A_936_333#_c_707_n 0.0198631f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_426 N_A_756_265#_c_508_n N_A_936_333#_c_708_n 0.00139051f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_427 N_A_756_265#_c_537_p N_A_936_333#_c_708_n 8.82602e-19 $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_428 N_A_756_265#_c_515_n N_A_936_333#_c_708_n 0.00174887f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_429 N_A_756_265#_c_516_n N_A_936_333#_c_708_n 0.0197641f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_430 N_A_756_265#_c_510_n N_A_936_333#_c_736_n 0.00569077f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_431 N_A_756_265#_c_508_n N_A_936_333#_c_717_n 0.00118695f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_432 N_A_756_265#_c_515_n N_A_936_333#_c_717_n 0.0177235f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_433 N_A_756_265#_c_516_n N_A_936_333#_c_717_n 2.87131e-19 $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_434 N_A_756_265#_M1016_g N_RESET_B_M1026_g 0.015492f $X=3.965 $Y=2.525 $X2=0
+ $Y2=0
cc_435 N_A_756_265#_c_512_n N_RESET_B_M1026_g 0.00134802f $X=4.08 $Y=1.295 $X2=0
+ $Y2=0
cc_436 N_A_756_265#_c_514_n N_RESET_B_M1026_g 0.0305402f $X=3.945 $Y=1.49 $X2=0
+ $Y2=0
cc_437 N_A_756_265#_c_512_n N_RESET_B_c_806_n 5.84967e-19 $X=4.08 $Y=1.295 $X2=0
+ $Y2=0
cc_438 N_A_756_265#_c_514_n N_RESET_B_c_806_n 0.00856697f $X=3.945 $Y=1.49 $X2=0
+ $Y2=0
cc_439 N_A_756_265#_c_517_n N_RESET_B_c_809_n 0.0099884f $X=4.9 $Y=1.125 $X2=0
+ $Y2=0
cc_440 N_A_756_265#_c_510_n N_RESET_B_c_815_n 0.00223631f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_441 N_A_756_265#_c_516_n N_RESET_B_c_815_n 4.47828e-19 $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_442 N_A_756_265#_M1021_g N_RESET_B_c_825_n 0.0142324f $X=7.77 $Y=2.88 $X2=0
+ $Y2=0
cc_443 N_A_756_265#_c_524_n N_RESET_B_c_825_n 0.0253467f $X=7.91 $Y=2.26 $X2=0
+ $Y2=0
cc_444 N_A_756_265#_c_525_n N_RESET_B_c_825_n 0.00560147f $X=7.91 $Y=2.26 $X2=0
+ $Y2=0
cc_445 N_A_756_265#_c_510_n N_RESET_B_c_816_n 0.00371297f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_446 N_A_756_265#_c_501_n N_A_808_463#_c_1005_n 0.0081345f $X=6.955 $Y=1.095
+ $X2=0 $Y2=0
cc_447 N_A_756_265#_M1016_g N_A_808_463#_c_1007_n 9.89135e-19 $X=3.965 $Y=2.525
+ $X2=0 $Y2=0
cc_448 N_A_756_265#_c_508_n N_A_808_463#_c_1007_n 0.0164278f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_449 N_A_756_265#_c_509_n N_A_808_463#_c_1007_n 0.00256146f $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_450 N_A_756_265#_c_537_p N_A_808_463#_c_1007_n 4.63228e-19 $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_451 N_A_756_265#_c_512_n N_A_808_463#_c_1007_n 0.0602052f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_452 N_A_756_265#_c_514_n N_A_808_463#_c_1007_n 6.35916e-19 $X=3.945 $Y=1.49
+ $X2=0 $Y2=0
cc_453 N_A_756_265#_c_515_n N_A_808_463#_c_1007_n 0.00208175f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_454 N_A_756_265#_c_516_n N_A_808_463#_c_1007_n 0.01744f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_455 N_A_756_265#_c_517_n N_A_808_463#_c_1007_n 0.00208975f $X=4.9 $Y=1.125
+ $X2=0 $Y2=0
cc_456 N_A_756_265#_c_510_n N_A_808_463#_c_1008_n 0.0261117f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_457 N_A_756_265#_c_537_p N_A_808_463#_c_1008_n 0.00213368f $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_458 N_A_756_265#_c_515_n N_A_808_463#_c_1008_n 0.00245586f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_459 N_A_756_265#_c_517_n N_A_808_463#_c_1008_n 0.00895602f $X=4.9 $Y=1.125
+ $X2=0 $Y2=0
cc_460 N_A_756_265#_c_510_n N_A_808_463#_c_1009_n 0.0205864f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_461 N_A_756_265#_M1016_g N_A_808_463#_c_1014_n 0.00184766f $X=3.965 $Y=2.525
+ $X2=0 $Y2=0
cc_462 N_A_756_265#_c_521_n N_A_808_463#_c_1014_n 4.15402e-19 $X=3.945 $Y=1.995
+ $X2=0 $Y2=0
cc_463 N_A_756_265#_c_512_n N_A_808_463#_c_1014_n 0.0137691f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_464 N_A_756_265#_c_508_n N_A_808_463#_c_1033_n 0.00993354f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_465 N_A_756_265#_c_515_n N_A_808_463#_c_1033_n 0.00151523f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_466 N_A_756_265#_c_516_n N_A_808_463#_c_1033_n 0.0279281f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_467 N_A_756_265#_c_503_n N_A_808_463#_c_1010_n 0.0081345f $X=7.03 $Y=1.17
+ $X2=0 $Y2=0
cc_468 N_A_756_265#_c_510_n N_A_808_463#_c_1010_n 0.00957152f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_469 N_A_756_265#_c_518_n N_A_808_463#_c_1010_n 0.00256292f $X=7.44 $Y=1.17
+ $X2=0 $Y2=0
cc_470 N_A_756_265#_M1016_g N_A_864_255#_M1001_g 0.020324f $X=3.965 $Y=2.525
+ $X2=0 $Y2=0
cc_471 N_A_756_265#_c_521_n N_A_864_255#_M1001_g 0.0198374f $X=3.945 $Y=1.995
+ $X2=0 $Y2=0
cc_472 N_A_756_265#_c_515_n N_A_864_255#_M1001_g 0.00137082f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_473 N_A_756_265#_c_508_n N_A_864_255#_M1031_g 0.00111681f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_474 N_A_756_265#_c_509_n N_A_864_255#_M1031_g 0.001085f $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_475 N_A_756_265#_c_512_n N_A_864_255#_M1031_g 0.00172363f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_476 N_A_756_265#_c_515_n N_A_864_255#_M1031_g 0.0192773f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_477 N_A_756_265#_c_516_n N_A_864_255#_M1031_g 3.98441e-19 $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_478 N_A_756_265#_c_517_n N_A_864_255#_M1031_g 0.0125029f $X=4.9 $Y=1.125
+ $X2=0 $Y2=0
cc_479 N_A_756_265#_M1021_g N_A_864_255#_c_1138_n 0.0136739f $X=7.77 $Y=2.88
+ $X2=0 $Y2=0
cc_480 N_A_756_265#_c_525_n N_A_864_255#_M1009_g 0.0136739f $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_481 N_A_756_265#_c_504_n N_A_864_255#_c_1126_n 0.00640393f $X=7.81 $Y=2.095
+ $X2=0 $Y2=0
cc_482 N_A_756_265#_c_507_n N_A_864_255#_c_1126_n 0.00482866f $X=7.725 $Y=1.26
+ $X2=0 $Y2=0
cc_483 N_A_756_265#_c_525_n N_A_864_255#_c_1126_n 0.00502506f $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_484 N_A_756_265#_c_518_n N_A_864_255#_c_1126_n 0.0206671f $X=7.44 $Y=1.17
+ $X2=0 $Y2=0
cc_485 N_A_756_265#_c_502_n N_A_864_255#_c_1127_n 0.00604095f $X=7.275 $Y=1.17
+ $X2=0 $Y2=0
cc_486 N_A_756_265#_c_504_n N_A_864_255#_M1027_g 0.00527992f $X=7.81 $Y=2.095
+ $X2=0 $Y2=0
cc_487 N_A_756_265#_c_507_n N_A_864_255#_M1027_g 0.00886932f $X=7.725 $Y=1.26
+ $X2=0 $Y2=0
cc_488 N_A_756_265#_c_511_n N_A_864_255#_M1027_g 0.00521164f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_489 N_A_756_265#_c_518_n N_A_864_255#_M1027_g 0.021379f $X=7.44 $Y=1.17 $X2=0
+ $Y2=0
cc_490 N_A_756_265#_c_505_n N_A_864_255#_M1006_g 0.0111347f $X=10.505 $Y=1.425
+ $X2=0 $Y2=0
cc_491 N_A_756_265#_c_506_n N_A_864_255#_M1002_g 0.00357707f $X=10.54 $Y=1.98
+ $X2=0 $Y2=0
cc_492 N_A_756_265#_c_508_n N_A_864_255#_c_1130_n 0.00405164f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_493 N_A_756_265#_c_509_n N_A_864_255#_c_1130_n 7.07929e-19 $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_494 N_A_756_265#_c_512_n N_A_864_255#_c_1130_n 0.00479343f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_495 N_A_756_265#_c_514_n N_A_864_255#_c_1130_n 0.0198374f $X=3.945 $Y=1.49
+ $X2=0 $Y2=0
cc_496 N_A_756_265#_c_504_n N_A_864_255#_c_1131_n 0.00992611f $X=7.81 $Y=2.095
+ $X2=0 $Y2=0
cc_497 N_A_756_265#_c_524_n N_A_864_255#_c_1131_n 0.0013102f $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_498 N_A_756_265#_c_525_n N_A_864_255#_c_1131_n 0.0175875f $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_499 N_A_756_265#_c_506_n N_A_864_255#_c_1132_n 0.0107027f $X=10.54 $Y=1.98
+ $X2=0 $Y2=0
cc_500 N_A_756_265#_c_511_n N_A_864_255#_c_1132_n 0.0176112f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_501 N_A_756_265#_c_504_n N_A_864_255#_c_1133_n 0.0242106f $X=7.81 $Y=2.095
+ $X2=0 $Y2=0
cc_502 N_A_756_265#_c_524_n N_A_864_255#_c_1133_n 6.25038e-19 $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_503 N_A_756_265#_c_511_n N_A_864_255#_c_1133_n 0.00192646f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_504 N_A_756_265#_c_506_n N_A_864_255#_c_1147_n 0.0239473f $X=10.54 $Y=1.98
+ $X2=0 $Y2=0
cc_505 N_A_756_265#_M1002_s N_A_864_255#_c_1148_n 0.00716549f $X=10.415 $Y=1.835
+ $X2=0 $Y2=0
cc_506 N_A_756_265#_c_506_n N_A_864_255#_c_1148_n 0.0202165f $X=10.54 $Y=1.98
+ $X2=0 $Y2=0
cc_507 N_A_756_265#_c_505_n N_A_864_255#_c_1134_n 0.0160491f $X=10.505 $Y=1.425
+ $X2=0 $Y2=0
cc_508 N_A_756_265#_c_506_n N_A_864_255#_c_1134_n 0.0202589f $X=10.54 $Y=1.98
+ $X2=0 $Y2=0
cc_509 N_A_756_265#_c_513_n N_A_864_255#_c_1134_n 3.36705e-19 $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_510 N_A_756_265#_c_506_n N_A_864_255#_c_1150_n 0.0264598f $X=10.54 $Y=1.98
+ $X2=0 $Y2=0
cc_511 N_A_756_265#_c_511_n N_A_864_255#_c_1135_n 0.0023718f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_512 N_A_756_265#_c_506_n N_A_864_255#_c_1136_n 0.00680211f $X=10.54 $Y=1.98
+ $X2=0 $Y2=0
cc_513 N_A_756_265#_c_506_n N_A_1406_69#_M1038_g 0.00282009f $X=10.54 $Y=1.98
+ $X2=0 $Y2=0
cc_514 N_A_756_265#_c_501_n N_A_1406_69#_c_1330_n 0.0067812f $X=6.955 $Y=1.095
+ $X2=0 $Y2=0
cc_515 N_A_756_265#_c_501_n N_A_1406_69#_c_1331_n 0.0035691f $X=6.955 $Y=1.095
+ $X2=0 $Y2=0
cc_516 N_A_756_265#_c_502_n N_A_1406_69#_c_1331_n 0.0095692f $X=7.275 $Y=1.17
+ $X2=0 $Y2=0
cc_517 N_A_756_265#_c_503_n N_A_1406_69#_c_1331_n 0.00196911f $X=7.03 $Y=1.17
+ $X2=0 $Y2=0
cc_518 N_A_756_265#_c_504_n N_A_1406_69#_c_1331_n 0.00598746f $X=7.81 $Y=2.095
+ $X2=0 $Y2=0
cc_519 N_A_756_265#_c_507_n N_A_1406_69#_c_1331_n 0.0224549f $X=7.725 $Y=1.26
+ $X2=0 $Y2=0
cc_520 N_A_756_265#_c_510_n N_A_1406_69#_c_1331_n 0.0164876f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_521 N_A_756_265#_c_637_p N_A_1406_69#_c_1331_n 0.00234811f $X=7.585 $Y=1.295
+ $X2=0 $Y2=0
cc_522 N_A_756_265#_c_518_n N_A_1406_69#_c_1331_n 0.00185918f $X=7.44 $Y=1.17
+ $X2=0 $Y2=0
cc_523 N_A_756_265#_c_502_n N_A_1406_69#_c_1332_n 0.0130244f $X=7.275 $Y=1.17
+ $X2=0 $Y2=0
cc_524 N_A_756_265#_c_507_n N_A_1406_69#_c_1332_n 0.0405372f $X=7.725 $Y=1.26
+ $X2=0 $Y2=0
cc_525 N_A_756_265#_c_510_n N_A_1406_69#_c_1332_n 0.00498772f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_526 N_A_756_265#_c_511_n N_A_1406_69#_c_1332_n 0.00909529f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_527 N_A_756_265#_c_637_p N_A_1406_69#_c_1332_n 0.00393315f $X=7.585 $Y=1.295
+ $X2=0 $Y2=0
cc_528 N_A_756_265#_c_502_n N_A_1406_69#_c_1333_n 0.00165058f $X=7.275 $Y=1.17
+ $X2=0 $Y2=0
cc_529 N_A_756_265#_c_503_n N_A_1406_69#_c_1333_n 2.73427e-19 $X=7.03 $Y=1.17
+ $X2=0 $Y2=0
cc_530 N_A_756_265#_c_504_n N_A_1406_69#_c_1333_n 0.0128089f $X=7.81 $Y=2.095
+ $X2=0 $Y2=0
cc_531 N_A_756_265#_c_507_n N_A_1406_69#_c_1333_n 0.0136185f $X=7.725 $Y=1.26
+ $X2=0 $Y2=0
cc_532 N_A_756_265#_c_510_n N_A_1406_69#_c_1333_n 0.00569361f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_533 N_A_756_265#_c_637_p N_A_1406_69#_c_1333_n 0.00366248f $X=7.585 $Y=1.295
+ $X2=0 $Y2=0
cc_534 N_A_756_265#_c_518_n N_A_1406_69#_c_1333_n 0.00252219f $X=7.44 $Y=1.17
+ $X2=0 $Y2=0
cc_535 N_A_756_265#_c_504_n N_A_1406_69#_c_1346_n 0.0247031f $X=7.81 $Y=2.095
+ $X2=0 $Y2=0
cc_536 N_A_756_265#_c_524_n N_A_1406_69#_c_1346_n 0.0199905f $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_537 N_A_756_265#_c_525_n N_A_1406_69#_c_1346_n 0.00249054f $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_538 N_A_756_265#_c_507_n N_A_1406_69#_c_1334_n 0.00853839f $X=7.725 $Y=1.26
+ $X2=0 $Y2=0
cc_539 N_A_756_265#_c_505_n N_A_1406_69#_c_1335_n 0.0101909f $X=10.505 $Y=1.425
+ $X2=0 $Y2=0
cc_540 N_A_756_265#_c_511_n N_A_1406_69#_c_1335_n 0.106559f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_541 N_A_756_265#_c_513_n N_A_1406_69#_c_1335_n 9.05304e-19 $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_542 N_A_756_265#_c_507_n N_A_1406_69#_c_1336_n 0.0123982f $X=7.725 $Y=1.26
+ $X2=0 $Y2=0
cc_543 N_A_756_265#_c_511_n N_A_1406_69#_c_1336_n 0.0150173f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_544 N_A_756_265#_c_505_n N_A_1406_69#_c_1337_n 0.0151241f $X=10.505 $Y=1.425
+ $X2=0 $Y2=0
cc_545 N_A_756_265#_c_513_n N_A_1406_69#_c_1337_n 7.23216e-19 $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_546 N_A_756_265#_M1006_s N_A_1406_69#_c_1338_n 0.00738119f $X=10.39 $Y=0.365
+ $X2=0 $Y2=0
cc_547 N_A_756_265#_c_505_n N_A_1406_69#_c_1338_n 0.0338824f $X=10.505 $Y=1.425
+ $X2=0 $Y2=0
cc_548 N_A_756_265#_c_511_n N_A_1406_69#_c_1338_n 0.00625944f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_549 N_A_756_265#_c_513_n N_A_1406_69#_c_1338_n 0.00261237f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_550 N_A_756_265#_c_505_n N_A_1406_69#_c_1342_n 0.00310076f $X=10.505 $Y=1.425
+ $X2=0 $Y2=0
cc_551 N_A_756_265#_c_506_n N_A_1406_69#_c_1342_n 0.00207875f $X=10.54 $Y=1.98
+ $X2=0 $Y2=0
cc_552 N_A_756_265#_c_513_n N_A_1406_69#_c_1342_n 9.04676e-19 $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_553 N_A_756_265#_M1021_g N_A_1635_21#_M1035_g 0.0234947f $X=7.77 $Y=2.88
+ $X2=0 $Y2=0
cc_554 N_A_756_265#_c_504_n N_A_1635_21#_c_1524_n 0.0030717f $X=7.81 $Y=2.095
+ $X2=0 $Y2=0
cc_555 N_A_756_265#_c_507_n N_A_1635_21#_c_1524_n 2.61975e-19 $X=7.725 $Y=1.26
+ $X2=0 $Y2=0
cc_556 N_A_756_265#_c_511_n N_A_1635_21#_c_1525_n 0.00225503f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_557 N_A_756_265#_c_504_n N_A_1635_21#_c_1533_n 0.00505417f $X=7.81 $Y=2.095
+ $X2=0 $Y2=0
cc_558 N_A_756_265#_c_524_n N_A_1635_21#_c_1533_n 0.00602931f $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_559 N_A_756_265#_c_525_n N_A_1635_21#_c_1533_n 2.22756e-19 $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_560 N_A_756_265#_c_524_n N_A_1635_21#_c_1534_n 0.00120163f $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_561 N_A_756_265#_c_525_n N_A_1635_21#_c_1534_n 0.0195609f $X=7.91 $Y=2.26
+ $X2=0 $Y2=0
cc_562 N_A_756_265#_c_505_n N_CLK_M1008_g 5.49749e-19 $X=10.505 $Y=1.425 $X2=0
+ $Y2=0
cc_563 N_A_756_265#_M1016_g N_VPWR_c_1787_n 0.00431487f $X=3.965 $Y=2.525 $X2=0
+ $Y2=0
cc_564 N_A_756_265#_M1021_g N_VPWR_c_1794_n 0.00420905f $X=7.77 $Y=2.88 $X2=0
+ $Y2=0
cc_565 N_A_756_265#_M1021_g N_VPWR_c_1795_n 0.00186772f $X=7.77 $Y=2.88 $X2=0
+ $Y2=0
cc_566 N_A_756_265#_M1002_s N_VPWR_c_1770_n 0.00389753f $X=10.415 $Y=1.835 $X2=0
+ $Y2=0
cc_567 N_A_756_265#_M1016_g N_VPWR_c_1770_n 0.00477801f $X=3.965 $Y=2.525 $X2=0
+ $Y2=0
cc_568 N_A_756_265#_M1021_g N_VPWR_c_1770_n 0.0067778f $X=7.77 $Y=2.88 $X2=0
+ $Y2=0
cc_569 N_A_756_265#_M1016_g N_A_380_50#_c_1932_n 0.00494899f $X=3.965 $Y=2.525
+ $X2=0 $Y2=0
cc_570 N_A_756_265#_c_509_n N_A_380_50#_c_1932_n 0.00139523f $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_571 N_A_756_265#_c_512_n N_A_380_50#_c_1932_n 0.0626292f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_572 N_A_756_265#_c_514_n N_A_380_50#_c_1932_n 0.00473435f $X=3.945 $Y=1.49
+ $X2=0 $Y2=0
cc_573 N_A_756_265#_c_512_n N_A_380_50#_c_1933_n 0.00838218f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_574 N_A_756_265#_c_514_n N_A_380_50#_c_1933_n 6.79402e-19 $X=3.945 $Y=1.49
+ $X2=0 $Y2=0
cc_575 N_A_756_265#_M1016_g N_A_380_50#_c_1940_n 0.0044447f $X=3.965 $Y=2.525
+ $X2=0 $Y2=0
cc_576 N_A_756_265#_c_521_n N_A_380_50#_c_1940_n 0.00317185f $X=3.945 $Y=1.995
+ $X2=0 $Y2=0
cc_577 N_A_756_265#_c_512_n N_A_380_50#_c_1940_n 0.00195293f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_578 N_A_756_265#_c_509_n N_A_380_50#_c_1936_n 0.00206819f $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_579 N_A_756_265#_c_512_n N_A_380_50#_c_1936_n 0.0207892f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_580 N_A_756_265#_c_514_n N_A_380_50#_c_1936_n 7.9056e-19 $X=3.945 $Y=1.49
+ $X2=0 $Y2=0
cc_581 N_A_756_265#_c_501_n N_VGND_c_2063_n 7.03502e-19 $X=6.955 $Y=1.095 $X2=0
+ $Y2=0
cc_582 N_A_756_265#_c_510_n N_VGND_c_2063_n 0.00121302f $X=7.295 $Y=1.295 $X2=0
+ $Y2=0
cc_583 N_A_756_265#_c_511_n N_VGND_c_2064_n 0.00266917f $X=10.175 $Y=1.295 $X2=0
+ $Y2=0
cc_584 N_A_756_265#_c_501_n N_VGND_c_2071_n 0.00452196f $X=6.955 $Y=1.095 $X2=0
+ $Y2=0
cc_585 N_A_756_265#_c_501_n N_VGND_c_2082_n 0.00892994f $X=6.955 $Y=1.095 $X2=0
+ $Y2=0
cc_586 N_A_756_265#_c_517_n N_VGND_c_2082_n 9.39239e-19 $X=4.9 $Y=1.125 $X2=0
+ $Y2=0
cc_587 N_A_936_333#_M1005_g N_RESET_B_c_809_n 0.0099884f $X=5.35 $Y=0.805 $X2=0
+ $Y2=0
cc_588 N_A_936_333#_c_706_n N_RESET_B_c_819_n 0.00771516f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_589 N_A_936_333#_M1004_g N_RESET_B_c_820_n 0.0186613f $X=4.755 $Y=2.525 $X2=0
+ $Y2=0
cc_590 N_A_936_333#_c_711_n N_RESET_B_c_820_n 0.0159515f $X=5.305 $Y=1.77 $X2=0
+ $Y2=0
cc_591 N_A_936_333#_c_706_n N_RESET_B_c_820_n 8.98955e-19 $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_592 N_A_936_333#_M1005_g N_RESET_B_M1037_g 0.0237671f $X=5.35 $Y=0.805 $X2=0
+ $Y2=0
cc_593 N_A_936_333#_M1005_g N_RESET_B_c_815_n 0.00756074f $X=5.35 $Y=0.805 $X2=0
+ $Y2=0
cc_594 N_A_936_333#_c_706_n N_RESET_B_c_815_n 2.62424e-19 $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_595 N_A_936_333#_c_706_n N_RESET_B_c_824_n 0.0162313f $X=6.645 $Y=1.685 $X2=0
+ $Y2=0
cc_596 N_A_936_333#_c_709_n N_RESET_B_c_824_n 2.96862e-19 $X=6.74 $Y=1.685 $X2=0
+ $Y2=0
cc_597 N_A_936_333#_c_736_n N_RESET_B_c_824_n 0.00683654f $X=6.935 $Y=2.04 $X2=0
+ $Y2=0
cc_598 N_A_936_333#_M1025_d N_RESET_B_c_825_n 0.0032773f $X=6.795 $Y=1.895 $X2=0
+ $Y2=0
cc_599 N_A_936_333#_c_736_n N_RESET_B_c_825_n 0.00455612f $X=6.935 $Y=2.04 $X2=0
+ $Y2=0
cc_600 N_A_936_333#_M1025_d N_RESET_B_c_862_n 0.00472583f $X=6.795 $Y=1.895
+ $X2=0 $Y2=0
cc_601 N_A_936_333#_c_736_n N_RESET_B_c_862_n 0.00847209f $X=6.935 $Y=2.04 $X2=0
+ $Y2=0
cc_602 N_A_936_333#_c_706_n RESET_B 0.0234126f $X=6.645 $Y=1.685 $X2=0 $Y2=0
cc_603 N_A_936_333#_c_736_n RESET_B 0.00558095f $X=6.935 $Y=2.04 $X2=0 $Y2=0
cc_604 N_A_936_333#_c_706_n N_RESET_B_c_828_n 0.00578877f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_605 N_A_936_333#_c_714_n N_RESET_B_c_828_n 4.43831e-19 $X=6.745 $Y=1.945
+ $X2=0 $Y2=0
cc_606 N_A_936_333#_c_736_n N_RESET_B_c_828_n 8.62668e-19 $X=6.935 $Y=2.04 $X2=0
+ $Y2=0
cc_607 N_A_936_333#_c_705_n N_RESET_B_c_816_n 0.0260645f $X=5.365 $Y=1.425 $X2=0
+ $Y2=0
cc_608 N_A_936_333#_c_706_n N_RESET_B_c_816_n 0.0153102f $X=6.645 $Y=1.685 $X2=0
+ $Y2=0
cc_609 N_A_936_333#_c_707_n N_A_808_463#_c_1005_n 0.00665378f $X=6.74 $Y=0.49
+ $X2=0 $Y2=0
cc_610 N_A_936_333#_c_714_n N_A_808_463#_M1025_g 0.0080555f $X=6.745 $Y=1.945
+ $X2=0 $Y2=0
cc_611 N_A_936_333#_c_709_n N_A_808_463#_M1025_g 0.00596229f $X=6.74 $Y=1.685
+ $X2=0 $Y2=0
cc_612 N_A_936_333#_c_736_n N_A_808_463#_M1025_g 0.00716141f $X=6.935 $Y=2.04
+ $X2=0 $Y2=0
cc_613 N_A_936_333#_M1004_g N_A_808_463#_c_1043_n 0.00146248f $X=4.755 $Y=2.525
+ $X2=0 $Y2=0
cc_614 N_A_936_333#_c_708_n N_A_808_463#_c_1007_n 0.0296188f $X=4.867 $Y=1.685
+ $X2=0 $Y2=0
cc_615 N_A_936_333#_c_717_n N_A_808_463#_c_1007_n 0.00576607f $X=5.01 $Y=1.83
+ $X2=0 $Y2=0
cc_616 N_A_936_333#_M1004_g N_A_808_463#_c_1013_n 0.0160791f $X=4.755 $Y=2.525
+ $X2=0 $Y2=0
cc_617 N_A_936_333#_c_711_n N_A_808_463#_c_1013_n 0.00446241f $X=5.305 $Y=1.77
+ $X2=0 $Y2=0
cc_618 N_A_936_333#_c_706_n N_A_808_463#_c_1013_n 0.0229505f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_619 N_A_936_333#_c_708_n N_A_808_463#_c_1013_n 0.0203583f $X=4.867 $Y=1.685
+ $X2=0 $Y2=0
cc_620 N_A_936_333#_c_717_n N_A_808_463#_c_1013_n 0.00124625f $X=5.01 $Y=1.83
+ $X2=0 $Y2=0
cc_621 N_A_936_333#_M1005_g N_A_808_463#_c_1008_n 0.013664f $X=5.35 $Y=0.805
+ $X2=0 $Y2=0
cc_622 N_A_936_333#_c_706_n N_A_808_463#_c_1008_n 0.0101864f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_623 N_A_936_333#_c_707_n N_A_808_463#_c_1008_n 0.0091919f $X=6.74 $Y=0.49
+ $X2=0 $Y2=0
cc_624 N_A_936_333#_M1004_g N_A_808_463#_c_1054_n 5.74677e-19 $X=4.755 $Y=2.525
+ $X2=0 $Y2=0
cc_625 N_A_936_333#_c_706_n N_A_808_463#_c_1009_n 0.0253868f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_626 N_A_936_333#_c_707_n N_A_808_463#_c_1009_n 0.0318053f $X=6.74 $Y=0.49
+ $X2=0 $Y2=0
cc_627 N_A_936_333#_c_717_n N_A_808_463#_c_1033_n 0.00127399f $X=5.01 $Y=1.83
+ $X2=0 $Y2=0
cc_628 N_A_936_333#_c_706_n N_A_808_463#_c_1010_n 0.00971916f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_629 N_A_936_333#_c_707_n N_A_808_463#_c_1010_n 0.0115221f $X=6.74 $Y=0.49
+ $X2=0 $Y2=0
cc_630 N_A_936_333#_c_709_n N_A_808_463#_c_1010_n 9.96648e-19 $X=6.74 $Y=1.685
+ $X2=0 $Y2=0
cc_631 N_A_936_333#_c_708_n N_A_864_255#_M1001_g 7.14877e-19 $X=4.867 $Y=1.685
+ $X2=0 $Y2=0
cc_632 N_A_936_333#_c_717_n N_A_864_255#_M1001_g 0.0734882f $X=5.01 $Y=1.83
+ $X2=0 $Y2=0
cc_633 N_A_936_333#_M1004_g N_A_864_255#_c_1138_n 0.0104164f $X=4.755 $Y=2.525
+ $X2=0 $Y2=0
cc_634 N_A_936_333#_c_736_n N_A_864_255#_M1009_g 0.00284124f $X=6.935 $Y=2.04
+ $X2=0 $Y2=0
cc_635 N_A_936_333#_c_714_n N_A_864_255#_c_1127_n 9.13899e-19 $X=6.745 $Y=1.945
+ $X2=0 $Y2=0
cc_636 N_A_936_333#_c_709_n N_A_864_255#_c_1127_n 4.54168e-19 $X=6.74 $Y=1.685
+ $X2=0 $Y2=0
cc_637 N_A_936_333#_c_707_n N_A_1406_69#_c_1330_n 0.0260046f $X=6.74 $Y=0.49
+ $X2=0 $Y2=0
cc_638 N_A_936_333#_c_707_n N_A_1406_69#_c_1331_n 0.0466069f $X=6.74 $Y=0.49
+ $X2=0 $Y2=0
cc_639 N_A_936_333#_c_709_n N_A_1406_69#_c_1331_n 4.22241e-19 $X=6.74 $Y=1.685
+ $X2=0 $Y2=0
cc_640 N_A_936_333#_c_709_n N_A_1406_69#_c_1333_n 0.0151212f $X=6.74 $Y=1.685
+ $X2=0 $Y2=0
cc_641 N_A_936_333#_c_736_n N_A_1406_69#_c_1333_n 0.00472143f $X=6.935 $Y=2.04
+ $X2=0 $Y2=0
cc_642 N_A_936_333#_c_714_n N_A_1406_69#_c_1346_n 0.00482692f $X=6.745 $Y=1.945
+ $X2=0 $Y2=0
cc_643 N_A_936_333#_M1004_g N_VPWR_c_1773_n 0.00382662f $X=4.755 $Y=2.525 $X2=0
+ $Y2=0
cc_644 N_A_936_333#_M1004_g N_VPWR_c_1770_n 9.39239e-19 $X=4.755 $Y=2.525 $X2=0
+ $Y2=0
cc_645 N_A_936_333#_c_707_n N_VGND_c_2063_n 0.0116085f $X=6.74 $Y=0.49 $X2=0
+ $Y2=0
cc_646 N_A_936_333#_c_707_n N_VGND_c_2071_n 0.00932149f $X=6.74 $Y=0.49 $X2=0
+ $Y2=0
cc_647 N_A_936_333#_M1005_g N_VGND_c_2082_n 9.39239e-19 $X=5.35 $Y=0.805 $X2=0
+ $Y2=0
cc_648 N_A_936_333#_c_707_n N_VGND_c_2082_n 0.00704609f $X=6.74 $Y=0.49 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_809_n N_A_808_463#_c_1005_n 0.0134019f $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_650 N_RESET_B_c_824_n N_A_808_463#_M1025_g 0.00801229f $X=6.755 $Y=2.39 $X2=0
+ $Y2=0
cc_651 N_RESET_B_c_825_n N_A_808_463#_M1025_g 2.03236e-19 $X=9.075 $Y=2.61 $X2=0
+ $Y2=0
cc_652 N_RESET_B_c_862_n N_A_808_463#_M1025_g 0.0113586f $X=6.84 $Y=2.39 $X2=0
+ $Y2=0
cc_653 RESET_B N_A_808_463#_M1025_g 0.00157507f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_654 N_RESET_B_c_828_n N_A_808_463#_M1025_g 0.0148666f $X=5.96 $Y=2.035 $X2=0
+ $Y2=0
cc_655 N_RESET_B_c_806_n N_A_808_463#_c_1007_n 5.43998e-19 $X=3.77 $Y=1.01 $X2=0
+ $Y2=0
cc_656 N_RESET_B_c_818_n N_A_808_463#_c_1013_n 0.0111585f $X=5.295 $Y=2.205
+ $X2=0 $Y2=0
cc_657 N_RESET_B_c_819_n N_A_808_463#_c_1013_n 0.00830323f $X=5.755 $Y=2.13
+ $X2=0 $Y2=0
cc_658 N_RESET_B_c_820_n N_A_808_463#_c_1013_n 0.00272396f $X=5.37 $Y=2.13 $X2=0
+ $Y2=0
cc_659 N_RESET_B_c_881_p N_A_808_463#_c_1013_n 0.00351361f $X=6.125 $Y=2.39
+ $X2=0 $Y2=0
cc_660 RESET_B N_A_808_463#_c_1013_n 0.0107899f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_661 N_RESET_B_c_828_n N_A_808_463#_c_1013_n 0.00128374f $X=5.96 $Y=2.035
+ $X2=0 $Y2=0
cc_662 N_RESET_B_c_809_n N_A_808_463#_c_1008_n 0.0131328f $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_663 N_RESET_B_M1037_g N_A_808_463#_c_1008_n 0.0167315f $X=5.86 $Y=0.775 $X2=0
+ $Y2=0
cc_664 N_RESET_B_c_815_n N_A_808_463#_c_1008_n 0.00101861f $X=5.845 $Y=1.245
+ $X2=0 $Y2=0
cc_665 N_RESET_B_c_818_n N_A_808_463#_c_1054_n 0.005098f $X=5.295 $Y=2.205 $X2=0
+ $Y2=0
cc_666 N_RESET_B_c_881_p N_A_808_463#_c_1054_n 0.0105188f $X=6.125 $Y=2.39 $X2=0
+ $Y2=0
cc_667 N_RESET_B_c_828_n N_A_808_463#_c_1054_n 0.0027915f $X=5.96 $Y=2.035 $X2=0
+ $Y2=0
cc_668 N_RESET_B_M1037_g N_A_808_463#_c_1009_n 0.00243259f $X=5.86 $Y=0.775
+ $X2=0 $Y2=0
cc_669 N_RESET_B_c_815_n N_A_808_463#_c_1009_n 0.00109845f $X=5.845 $Y=1.245
+ $X2=0 $Y2=0
cc_670 N_RESET_B_c_816_n N_A_808_463#_c_1009_n 0.00175977f $X=5.94 $Y=1.87 $X2=0
+ $Y2=0
cc_671 N_RESET_B_c_809_n N_A_808_463#_c_1033_n 0.00488344f $X=5.785 $Y=0.18
+ $X2=0 $Y2=0
cc_672 N_RESET_B_c_815_n N_A_808_463#_c_1010_n 0.0100968f $X=5.845 $Y=1.245
+ $X2=0 $Y2=0
cc_673 N_RESET_B_c_824_n N_A_808_463#_c_1010_n 6.9488e-19 $X=6.755 $Y=2.39 $X2=0
+ $Y2=0
cc_674 N_RESET_B_c_816_n N_A_808_463#_c_1010_n 0.0162747f $X=5.94 $Y=1.87 $X2=0
+ $Y2=0
cc_675 N_RESET_B_c_808_n N_A_864_255#_M1031_g 0.0136977f $X=3.845 $Y=0.935 $X2=0
+ $Y2=0
cc_676 N_RESET_B_c_809_n N_A_864_255#_M1031_g 0.0098336f $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_677 N_RESET_B_c_818_n N_A_864_255#_c_1138_n 0.0103572f $X=5.295 $Y=2.205
+ $X2=0 $Y2=0
cc_678 N_RESET_B_c_824_n N_A_864_255#_c_1138_n 0.00488319f $X=6.755 $Y=2.39
+ $X2=0 $Y2=0
cc_679 N_RESET_B_c_881_p N_A_864_255#_c_1138_n 0.00154627f $X=6.125 $Y=2.39
+ $X2=0 $Y2=0
cc_680 N_RESET_B_c_825_n N_A_864_255#_c_1138_n 0.00106324f $X=9.075 $Y=2.61
+ $X2=0 $Y2=0
cc_681 N_RESET_B_c_862_n N_A_864_255#_c_1138_n 0.00221383f $X=6.84 $Y=2.39 $X2=0
+ $Y2=0
cc_682 N_RESET_B_c_828_n N_A_864_255#_c_1138_n 0.00856175f $X=5.96 $Y=2.035
+ $X2=0 $Y2=0
cc_683 N_RESET_B_c_825_n N_A_864_255#_M1009_g 0.0159644f $X=9.075 $Y=2.61 $X2=0
+ $Y2=0
cc_684 N_RESET_B_c_862_n N_A_864_255#_M1009_g 0.00419552f $X=6.84 $Y=2.39 $X2=0
+ $Y2=0
cc_685 N_RESET_B_c_812_n N_A_864_255#_c_1132_n 0.00877029f $X=9.255 $Y=1.59
+ $X2=0 $Y2=0
cc_686 N_RESET_B_c_813_n N_A_864_255#_c_1132_n 0.00679121f $X=9.045 $Y=1.59
+ $X2=0 $Y2=0
cc_687 N_RESET_B_c_830_n N_A_864_255#_c_1132_n 0.00474148f $X=9.24 $Y=2.18 $X2=0
+ $Y2=0
cc_688 N_RESET_B_c_825_n N_A_864_255#_c_1133_n 0.00670596f $X=9.075 $Y=2.61
+ $X2=0 $Y2=0
cc_689 N_RESET_B_c_825_n N_A_864_255#_c_1135_n 0.00106466f $X=9.075 $Y=2.61
+ $X2=0 $Y2=0
cc_690 N_RESET_B_c_825_n N_A_1406_69#_M1009_d 0.0112959f $X=9.075 $Y=2.61 $X2=0
+ $Y2=0
cc_691 N_RESET_B_M1034_g N_A_1406_69#_c_1322_n 0.0499387f $X=8.97 $Y=0.805 $X2=0
+ $Y2=0
cc_692 N_RESET_B_c_812_n N_A_1406_69#_c_1324_n 0.00836713f $X=9.255 $Y=1.59
+ $X2=0 $Y2=0
cc_693 N_RESET_B_c_812_n N_A_1406_69#_M1038_g 0.0629713f $X=9.255 $Y=1.59 $X2=0
+ $Y2=0
cc_694 N_RESET_B_M1014_g N_A_1406_69#_M1038_g 0.0177344f $X=9.26 $Y=2.88 $X2=0
+ $Y2=0
cc_695 N_RESET_B_c_826_n N_A_1406_69#_M1038_g 9.25684e-19 $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_696 N_RESET_B_c_825_n N_A_1406_69#_c_1346_n 0.0218449f $X=9.075 $Y=2.61 $X2=0
+ $Y2=0
cc_697 N_RESET_B_M1034_g N_A_1406_69#_c_1334_n 0.00161777f $X=8.97 $Y=0.805
+ $X2=0 $Y2=0
cc_698 N_RESET_B_M1034_g N_A_1406_69#_c_1335_n 0.0151403f $X=8.97 $Y=0.805 $X2=0
+ $Y2=0
cc_699 N_RESET_B_c_812_n N_A_1406_69#_c_1335_n 0.00519904f $X=9.255 $Y=1.59
+ $X2=0 $Y2=0
cc_700 N_RESET_B_M1034_g N_A_1406_69#_c_1342_n 0.00540417f $X=8.97 $Y=0.805
+ $X2=0 $Y2=0
cc_701 N_RESET_B_c_826_n N_A_1635_21#_M1014_d 3.47647e-19 $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_702 N_RESET_B_M1034_g N_A_1635_21#_M1017_g 0.00687393f $X=8.97 $Y=0.805 $X2=0
+ $Y2=0
cc_703 N_RESET_B_c_825_n N_A_1635_21#_M1035_g 0.0176553f $X=9.075 $Y=2.61 $X2=0
+ $Y2=0
cc_704 N_RESET_B_c_826_n N_A_1635_21#_M1035_g 0.00181127f $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_705 N_RESET_B_c_827_n N_A_1635_21#_M1035_g 0.00478863f $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_706 N_RESET_B_M1034_g N_A_1635_21#_c_1520_n 0.0104164f $X=8.97 $Y=0.805 $X2=0
+ $Y2=0
cc_707 N_RESET_B_M1034_g N_A_1635_21#_c_1522_n 0.0190129f $X=8.97 $Y=0.805 $X2=0
+ $Y2=0
cc_708 N_RESET_B_c_813_n N_A_1635_21#_c_1524_n 0.0190129f $X=9.045 $Y=1.59 $X2=0
+ $Y2=0
cc_709 N_RESET_B_c_830_n N_A_1635_21#_c_1524_n 0.00627154f $X=9.24 $Y=2.18 $X2=0
+ $Y2=0
cc_710 N_RESET_B_c_813_n N_A_1635_21#_c_1531_n 0.00162926f $X=9.045 $Y=1.59
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_825_n N_A_1635_21#_c_1531_n 0.00813358f $X=9.075 $Y=2.61
+ $X2=0 $Y2=0
cc_712 N_RESET_B_c_826_n N_A_1635_21#_c_1531_n 0.0247905f $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_713 N_RESET_B_c_827_n N_A_1635_21#_c_1531_n 0.00195903f $X=9.24 $Y=2.345
+ $X2=0 $Y2=0
cc_714 N_RESET_B_c_830_n N_A_1635_21#_c_1531_n 0.0105392f $X=9.24 $Y=2.18 $X2=0
+ $Y2=0
cc_715 N_RESET_B_M1014_g N_A_1635_21#_c_1558_n 0.0027538f $X=9.26 $Y=2.88 $X2=0
+ $Y2=0
cc_716 N_RESET_B_c_826_n N_A_1635_21#_c_1558_n 0.00263578f $X=9.24 $Y=2.345
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_827_n N_A_1635_21#_c_1558_n 2.22629e-19 $X=9.24 $Y=2.345
+ $X2=0 $Y2=0
cc_718 N_RESET_B_M1034_g N_A_1635_21#_c_1525_n 0.00146886f $X=8.97 $Y=0.805
+ $X2=0 $Y2=0
cc_719 N_RESET_B_M1014_g N_A_1635_21#_c_1532_n 4.47615e-19 $X=9.26 $Y=2.88 $X2=0
+ $Y2=0
cc_720 N_RESET_B_c_826_n N_A_1635_21#_c_1532_n 0.0318225f $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_721 N_RESET_B_c_830_n N_A_1635_21#_c_1532_n 0.00473438f $X=9.24 $Y=2.18 $X2=0
+ $Y2=0
cc_722 N_RESET_B_c_825_n N_A_1635_21#_c_1533_n 0.0186812f $X=9.075 $Y=2.61 $X2=0
+ $Y2=0
cc_723 N_RESET_B_c_826_n N_A_1635_21#_c_1533_n 0.00158434f $X=9.24 $Y=2.345
+ $X2=0 $Y2=0
cc_724 N_RESET_B_c_827_n N_A_1635_21#_c_1533_n 5.86558e-19 $X=9.24 $Y=2.345
+ $X2=0 $Y2=0
cc_725 N_RESET_B_c_830_n N_A_1635_21#_c_1533_n 6.9692e-19 $X=9.24 $Y=2.18 $X2=0
+ $Y2=0
cc_726 N_RESET_B_c_825_n N_A_1635_21#_c_1534_n 0.00530107f $X=9.075 $Y=2.61
+ $X2=0 $Y2=0
cc_727 N_RESET_B_c_827_n N_A_1635_21#_c_1534_n 0.00655646f $X=9.24 $Y=2.345
+ $X2=0 $Y2=0
cc_728 N_RESET_B_c_830_n N_A_1635_21#_c_1534_n 0.00750546f $X=9.24 $Y=2.18 $X2=0
+ $Y2=0
cc_729 N_RESET_B_c_824_n N_VPWR_M1025_s 0.0097762f $X=6.755 $Y=2.39 $X2=0 $Y2=0
cc_730 N_RESET_B_c_825_n N_VPWR_M1035_d 0.00642498f $X=9.075 $Y=2.61 $X2=0 $Y2=0
cc_731 N_RESET_B_c_826_n N_VPWR_M1035_d 6.14024e-19 $X=9.24 $Y=2.345 $X2=0 $Y2=0
cc_732 N_RESET_B_M1026_g N_VPWR_c_1772_n 0.00659433f $X=3.44 $Y=2.635 $X2=0
+ $Y2=0
cc_733 N_RESET_B_c_818_n N_VPWR_c_1773_n 0.00505974f $X=5.295 $Y=2.205 $X2=0
+ $Y2=0
cc_734 N_RESET_B_c_824_n N_VPWR_c_1774_n 0.0262522f $X=6.755 $Y=2.39 $X2=0 $Y2=0
cc_735 N_RESET_B_c_862_n N_VPWR_c_1774_n 0.00354025f $X=6.84 $Y=2.39 $X2=0 $Y2=0
cc_736 N_RESET_B_M1014_g N_VPWR_c_1782_n 0.00409721f $X=9.26 $Y=2.88 $X2=0 $Y2=0
cc_737 N_RESET_B_c_826_n N_VPWR_c_1782_n 0.00260876f $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_738 N_RESET_B_M1026_g N_VPWR_c_1787_n 0.00452955f $X=3.44 $Y=2.635 $X2=0
+ $Y2=0
cc_739 N_RESET_B_c_825_n N_VPWR_c_1794_n 0.0232542f $X=9.075 $Y=2.61 $X2=0 $Y2=0
cc_740 N_RESET_B_c_862_n N_VPWR_c_1794_n 0.00256552f $X=6.84 $Y=2.39 $X2=0 $Y2=0
cc_741 N_RESET_B_M1014_g N_VPWR_c_1795_n 0.00920347f $X=9.26 $Y=2.88 $X2=0 $Y2=0
cc_742 N_RESET_B_c_825_n N_VPWR_c_1795_n 0.0459408f $X=9.075 $Y=2.61 $X2=0 $Y2=0
cc_743 N_RESET_B_c_826_n N_VPWR_c_1795_n 0.00422691f $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_744 N_RESET_B_c_827_n N_VPWR_c_1795_n 2.96715e-19 $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_745 N_RESET_B_M1026_g N_VPWR_c_1770_n 0.00544287f $X=3.44 $Y=2.635 $X2=0
+ $Y2=0
cc_746 N_RESET_B_c_818_n N_VPWR_c_1770_n 9.39239e-19 $X=5.295 $Y=2.205 $X2=0
+ $Y2=0
cc_747 N_RESET_B_M1014_g N_VPWR_c_1770_n 0.00705209f $X=9.26 $Y=2.88 $X2=0 $Y2=0
cc_748 N_RESET_B_c_824_n N_VPWR_c_1770_n 0.00980357f $X=6.755 $Y=2.39 $X2=0
+ $Y2=0
cc_749 N_RESET_B_c_881_p N_VPWR_c_1770_n 0.0100179f $X=6.125 $Y=2.39 $X2=0 $Y2=0
cc_750 N_RESET_B_c_825_n N_VPWR_c_1770_n 0.0426704f $X=9.075 $Y=2.61 $X2=0 $Y2=0
cc_751 N_RESET_B_c_862_n N_VPWR_c_1770_n 0.00426564f $X=6.84 $Y=2.39 $X2=0 $Y2=0
cc_752 N_RESET_B_c_826_n N_VPWR_c_1770_n 0.00492433f $X=9.24 $Y=2.345 $X2=0
+ $Y2=0
cc_753 N_RESET_B_c_828_n N_VPWR_c_1770_n 0.00235298f $X=5.96 $Y=2.035 $X2=0
+ $Y2=0
cc_754 N_RESET_B_M1019_g N_A_380_50#_c_1931_n 0.00624478f $X=3.29 $Y=0.615 $X2=0
+ $Y2=0
cc_755 N_RESET_B_c_807_n N_A_380_50#_c_1931_n 0.00995357f $X=3.515 $Y=1.01 $X2=0
+ $Y2=0
cc_756 N_RESET_B_M1026_g N_A_380_50#_c_1937_n 0.0101934f $X=3.44 $Y=2.635 $X2=0
+ $Y2=0
cc_757 N_RESET_B_M1026_g N_A_380_50#_c_1932_n 0.0302853f $X=3.44 $Y=2.635 $X2=0
+ $Y2=0
cc_758 N_RESET_B_c_806_n N_A_380_50#_c_1932_n 0.00673681f $X=3.77 $Y=1.01 $X2=0
+ $Y2=0
cc_759 N_RESET_B_c_807_n N_A_380_50#_c_1932_n 0.00184838f $X=3.515 $Y=1.01 $X2=0
+ $Y2=0
cc_760 N_RESET_B_c_806_n N_A_380_50#_c_1933_n 0.00716031f $X=3.77 $Y=1.01 $X2=0
+ $Y2=0
cc_761 N_RESET_B_c_808_n N_A_380_50#_c_1933_n 0.00585807f $X=3.845 $Y=0.935
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_803_n N_A_380_50#_c_1935_n 4.69055e-19 $X=3.77 $Y=0.18 $X2=0
+ $Y2=0
cc_763 N_RESET_B_c_806_n N_A_380_50#_c_1935_n 0.00313934f $X=3.77 $Y=1.01 $X2=0
+ $Y2=0
cc_764 N_RESET_B_c_807_n N_A_380_50#_c_1935_n 0.00114854f $X=3.515 $Y=1.01 $X2=0
+ $Y2=0
cc_765 N_RESET_B_M1026_g N_A_380_50#_c_1940_n 0.013489f $X=3.44 $Y=2.635 $X2=0
+ $Y2=0
cc_766 N_RESET_B_c_808_n N_A_380_50#_c_1936_n 0.00579032f $X=3.845 $Y=0.935
+ $X2=0 $Y2=0
cc_767 N_RESET_B_c_809_n N_A_380_50#_c_1936_n 0.0037685f $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_768 N_RESET_B_c_825_n A_1569_534# 0.00578273f $X=9.075 $Y=2.61 $X2=-0.19
+ $Y2=-0.245
cc_769 N_RESET_B_M1019_g N_VGND_c_2062_n 0.00211288f $X=3.29 $Y=0.615 $X2=0
+ $Y2=0
cc_770 N_RESET_B_c_803_n N_VGND_c_2062_n 0.0217783f $X=3.77 $Y=0.18 $X2=0 $Y2=0
cc_771 N_RESET_B_c_807_n N_VGND_c_2062_n 8.80271e-19 $X=3.515 $Y=1.01 $X2=0
+ $Y2=0
cc_772 N_RESET_B_c_808_n N_VGND_c_2062_n 0.00893666f $X=3.845 $Y=0.935 $X2=0
+ $Y2=0
cc_773 N_RESET_B_c_809_n N_VGND_c_2063_n 0.0128616f $X=5.785 $Y=0.18 $X2=0 $Y2=0
cc_774 N_RESET_B_M1034_g N_VGND_c_2064_n 0.00763063f $X=8.97 $Y=0.805 $X2=0
+ $Y2=0
cc_775 N_RESET_B_c_803_n N_VGND_c_2069_n 0.0723339f $X=3.77 $Y=0.18 $X2=0 $Y2=0
cc_776 N_RESET_B_c_804_n N_VGND_c_2076_n 0.00724047f $X=3.365 $Y=0.18 $X2=0
+ $Y2=0
cc_777 N_RESET_B_c_803_n N_VGND_c_2082_n 0.00217301f $X=3.77 $Y=0.18 $X2=0 $Y2=0
cc_778 N_RESET_B_c_804_n N_VGND_c_2082_n 0.00691715f $X=3.365 $Y=0.18 $X2=0
+ $Y2=0
cc_779 N_RESET_B_c_809_n N_VGND_c_2082_n 0.0636944f $X=5.785 $Y=0.18 $X2=0 $Y2=0
cc_780 N_RESET_B_M1034_g N_VGND_c_2082_n 9.39239e-19 $X=8.97 $Y=0.805 $X2=0
+ $Y2=0
cc_781 N_RESET_B_c_814_n N_VGND_c_2082_n 0.00463263f $X=3.845 $Y=0.18 $X2=0
+ $Y2=0
cc_782 N_RESET_B_M1019_g N_noxref_24_c_2206_n 0.00624612f $X=3.29 $Y=0.615 $X2=0
+ $Y2=0
cc_783 N_A_808_463#_c_1043_n N_A_864_255#_M1001_g 0.00825723f $X=4.18 $Y=2.53
+ $X2=0 $Y2=0
cc_784 N_A_808_463#_c_1007_n N_A_864_255#_M1001_g 0.0173643f $X=4.47 $Y=2.175
+ $X2=0 $Y2=0
cc_785 N_A_808_463#_c_1014_n N_A_864_255#_M1001_g 0.0130765f $X=4.305 $Y=2.26
+ $X2=0 $Y2=0
cc_786 N_A_808_463#_c_1007_n N_A_864_255#_M1031_g 0.0101271f $X=4.47 $Y=2.175
+ $X2=0 $Y2=0
cc_787 N_A_808_463#_c_1033_n N_A_864_255#_M1031_g 0.00893971f $X=4.8 $Y=0.817
+ $X2=0 $Y2=0
cc_788 N_A_808_463#_M1025_g N_A_864_255#_c_1138_n 0.00999463f $X=6.72 $Y=2.315
+ $X2=0 $Y2=0
cc_789 N_A_808_463#_c_1054_n N_A_864_255#_c_1138_n 0.00454409f $X=5.51 $Y=2.53
+ $X2=0 $Y2=0
cc_790 N_A_808_463#_M1025_g N_A_864_255#_c_1127_n 0.0389841f $X=6.72 $Y=2.315
+ $X2=0 $Y2=0
cc_791 N_A_808_463#_c_1007_n N_A_864_255#_c_1130_n 0.00426747f $X=4.47 $Y=2.175
+ $X2=0 $Y2=0
cc_792 N_A_808_463#_c_1010_n N_A_1406_69#_c_1331_n 7.72467e-19 $X=6.525 $Y=1.365
+ $X2=0 $Y2=0
cc_793 N_A_808_463#_c_1010_n N_A_1406_69#_c_1333_n 7.61567e-19 $X=6.525 $Y=1.365
+ $X2=0 $Y2=0
cc_794 N_A_808_463#_c_1013_n N_VPWR_M1004_d 0.00298209f $X=5.355 $Y=2.26 $X2=0
+ $Y2=0
cc_795 N_A_808_463#_c_1013_n N_VPWR_c_1773_n 0.022455f $X=5.355 $Y=2.26 $X2=0
+ $Y2=0
cc_796 N_A_808_463#_M1025_g N_VPWR_c_1774_n 0.00813936f $X=6.72 $Y=2.315 $X2=0
+ $Y2=0
cc_797 N_A_808_463#_c_1054_n N_VPWR_c_1774_n 0.00158406f $X=5.51 $Y=2.53 $X2=0
+ $Y2=0
cc_798 N_A_808_463#_c_1043_n N_VPWR_c_1787_n 0.00521857f $X=4.18 $Y=2.53 $X2=0
+ $Y2=0
cc_799 N_A_808_463#_c_1054_n N_VPWR_c_1788_n 0.00452011f $X=5.51 $Y=2.53 $X2=0
+ $Y2=0
cc_800 N_A_808_463#_M1025_g N_VPWR_c_1770_n 9.39239e-19 $X=6.72 $Y=2.315 $X2=0
+ $Y2=0
cc_801 N_A_808_463#_c_1043_n N_VPWR_c_1770_n 0.00949055f $X=4.18 $Y=2.53 $X2=0
+ $Y2=0
cc_802 N_A_808_463#_c_1054_n N_VPWR_c_1770_n 0.00694919f $X=5.51 $Y=2.53 $X2=0
+ $Y2=0
cc_803 N_A_808_463#_c_1014_n N_A_380_50#_c_1932_n 0.00616821f $X=4.305 $Y=2.26
+ $X2=0 $Y2=0
cc_804 N_A_808_463#_c_1014_n N_A_380_50#_c_1940_n 0.00131082f $X=4.305 $Y=2.26
+ $X2=0 $Y2=0
cc_805 N_A_808_463#_c_1007_n N_A_380_50#_c_1936_n 7.25909e-19 $X=4.47 $Y=2.175
+ $X2=0 $Y2=0
cc_806 N_A_808_463#_c_1033_n N_A_380_50#_c_1936_n 0.0281522f $X=4.8 $Y=0.817
+ $X2=0 $Y2=0
cc_807 N_A_808_463#_c_1013_n A_894_463# 0.00255642f $X=5.355 $Y=2.26 $X2=-0.19
+ $Y2=-0.245
cc_808 N_A_808_463#_c_1014_n A_894_463# 0.00126309f $X=4.305 $Y=2.26 $X2=-0.19
+ $Y2=-0.245
cc_809 N_A_808_463#_c_1008_n N_VGND_M1037_d 0.00677207f $X=6.145 $Y=0.89 $X2=0
+ $Y2=0
cc_810 N_A_808_463#_c_1005_n N_VGND_c_2063_n 0.00777284f $X=6.525 $Y=1.095 $X2=0
+ $Y2=0
cc_811 N_A_808_463#_c_1008_n N_VGND_c_2063_n 0.0229474f $X=6.145 $Y=0.89 $X2=0
+ $Y2=0
cc_812 N_A_808_463#_c_1010_n N_VGND_c_2063_n 0.00113735f $X=6.525 $Y=1.365 $X2=0
+ $Y2=0
cc_813 N_A_808_463#_c_1033_n N_VGND_c_2069_n 0.00642607f $X=4.8 $Y=0.817 $X2=0
+ $Y2=0
cc_814 N_A_808_463#_c_1005_n N_VGND_c_2071_n 0.00400407f $X=6.525 $Y=1.095 $X2=0
+ $Y2=0
cc_815 N_A_808_463#_c_1005_n N_VGND_c_2082_n 0.00775088f $X=6.525 $Y=1.095 $X2=0
+ $Y2=0
cc_816 N_A_808_463#_c_1008_n N_VGND_c_2082_n 0.0449925f $X=6.145 $Y=0.89 $X2=0
+ $Y2=0
cc_817 N_A_808_463#_c_1033_n N_VGND_c_2082_n 0.0103691f $X=4.8 $Y=0.817 $X2=0
+ $Y2=0
cc_818 N_A_808_463#_c_1008_n A_991_119# 0.00370984f $X=6.145 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_819 N_A_808_463#_c_1008_n A_1085_119# 0.00569011f $X=6.145 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_820 N_A_864_255#_c_1132_n N_A_1406_69#_c_1323_n 0.00114455f $X=9.935 $Y=1.645
+ $X2=0 $Y2=0
cc_821 N_A_864_255#_c_1132_n N_A_1406_69#_M1038_g 0.0118345f $X=9.935 $Y=1.645
+ $X2=0 $Y2=0
cc_822 N_A_864_255#_c_1147_n N_A_1406_69#_M1038_g 0.0141129f $X=10.02 $Y=2.325
+ $X2=0 $Y2=0
cc_823 N_A_864_255#_c_1149_n N_A_1406_69#_M1038_g 0.0034218f $X=10.105 $Y=2.41
+ $X2=0 $Y2=0
cc_824 N_A_864_255#_c_1134_n N_A_1406_69#_c_1328_n 9.70421e-19 $X=11.132
+ $Y=1.672 $X2=0 $Y2=0
cc_825 N_A_864_255#_c_1127_n N_A_1406_69#_c_1331_n 3.44645e-19 $X=7.225 $Y=1.71
+ $X2=0 $Y2=0
cc_826 N_A_864_255#_M1027_g N_A_1406_69#_c_1331_n 0.00418298f $X=7.89 $Y=0.775
+ $X2=0 $Y2=0
cc_827 N_A_864_255#_M1027_g N_A_1406_69#_c_1332_n 0.0193956f $X=7.89 $Y=0.775
+ $X2=0 $Y2=0
cc_828 N_A_864_255#_c_1135_n N_A_1406_69#_c_1332_n 0.00184846f $X=8.16 $Y=1.72
+ $X2=0 $Y2=0
cc_829 N_A_864_255#_c_1126_n N_A_1406_69#_c_1333_n 0.00973464f $X=7.815 $Y=1.71
+ $X2=0 $Y2=0
cc_830 N_A_864_255#_c_1127_n N_A_1406_69#_c_1333_n 0.00946274f $X=7.225 $Y=1.71
+ $X2=0 $Y2=0
cc_831 N_A_864_255#_M1009_g N_A_1406_69#_c_1346_n 0.00370806f $X=7.15 $Y=2.315
+ $X2=0 $Y2=0
cc_832 N_A_864_255#_c_1126_n N_A_1406_69#_c_1346_n 0.00791899f $X=7.815 $Y=1.71
+ $X2=0 $Y2=0
cc_833 N_A_864_255#_c_1131_n N_A_1406_69#_c_1346_n 3.35785e-19 $X=7.89 $Y=1.72
+ $X2=0 $Y2=0
cc_834 N_A_864_255#_M1027_g N_A_1406_69#_c_1334_n 0.00426555f $X=7.89 $Y=0.775
+ $X2=0 $Y2=0
cc_835 N_A_864_255#_c_1132_n N_A_1406_69#_c_1335_n 0.103381f $X=9.935 $Y=1.645
+ $X2=0 $Y2=0
cc_836 N_A_864_255#_c_1133_n N_A_1406_69#_c_1335_n 0.00569984f $X=8.325 $Y=1.645
+ $X2=0 $Y2=0
cc_837 N_A_864_255#_c_1135_n N_A_1406_69#_c_1335_n 5.58847e-19 $X=8.16 $Y=1.72
+ $X2=0 $Y2=0
cc_838 N_A_864_255#_M1027_g N_A_1406_69#_c_1336_n 0.00217729f $X=7.89 $Y=0.775
+ $X2=0 $Y2=0
cc_839 N_A_864_255#_c_1133_n N_A_1406_69#_c_1336_n 0.0125877f $X=8.325 $Y=1.645
+ $X2=0 $Y2=0
cc_840 N_A_864_255#_c_1135_n N_A_1406_69#_c_1336_n 0.00111299f $X=8.16 $Y=1.72
+ $X2=0 $Y2=0
cc_841 N_A_864_255#_M1006_g N_A_1406_69#_c_1337_n 0.00244513f $X=10.75 $Y=0.785
+ $X2=0 $Y2=0
cc_842 N_A_864_255#_M1008_d N_A_1406_69#_c_1338_n 0.00716655f $X=11.415 $Y=0.365
+ $X2=0 $Y2=0
cc_843 N_A_864_255#_M1006_g N_A_1406_69#_c_1338_n 0.0179382f $X=10.75 $Y=0.785
+ $X2=0 $Y2=0
cc_844 N_A_864_255#_c_1134_n N_A_1406_69#_c_1338_n 0.0429283f $X=11.132 $Y=1.672
+ $X2=0 $Y2=0
cc_845 N_A_864_255#_c_1136_n N_A_1406_69#_c_1338_n 0.00104471f $X=10.89 $Y=1.51
+ $X2=0 $Y2=0
cc_846 N_A_864_255#_c_1134_n N_A_1406_69#_c_1340_n 0.0223818f $X=11.132 $Y=1.672
+ $X2=0 $Y2=0
cc_847 N_A_864_255#_c_1132_n N_A_1406_69#_c_1342_n 0.00472619f $X=9.935 $Y=1.645
+ $X2=0 $Y2=0
cc_848 N_A_864_255#_M1027_g N_A_1635_21#_M1017_g 0.0504619f $X=7.89 $Y=0.775
+ $X2=0 $Y2=0
cc_849 N_A_864_255#_c_1132_n N_A_1635_21#_c_1522_n 0.0010707f $X=9.935 $Y=1.645
+ $X2=0 $Y2=0
cc_850 N_A_864_255#_c_1135_n N_A_1635_21#_c_1523_n 0.00581981f $X=8.16 $Y=1.72
+ $X2=0 $Y2=0
cc_851 N_A_864_255#_M1027_g N_A_1635_21#_c_1524_n 0.00456443f $X=7.89 $Y=0.775
+ $X2=0 $Y2=0
cc_852 N_A_864_255#_c_1132_n N_A_1635_21#_c_1524_n 0.0101757f $X=9.935 $Y=1.645
+ $X2=0 $Y2=0
cc_853 N_A_864_255#_c_1133_n N_A_1635_21#_c_1524_n 0.00106783f $X=8.325 $Y=1.645
+ $X2=0 $Y2=0
cc_854 N_A_864_255#_c_1135_n N_A_1635_21#_c_1524_n 0.0206052f $X=8.16 $Y=1.72
+ $X2=0 $Y2=0
cc_855 N_A_864_255#_c_1132_n N_A_1635_21#_c_1531_n 0.061251f $X=9.935 $Y=1.645
+ $X2=0 $Y2=0
cc_856 N_A_864_255#_c_1147_n N_A_1635_21#_c_1531_n 0.0130074f $X=10.02 $Y=2.325
+ $X2=0 $Y2=0
cc_857 N_A_864_255#_c_1147_n N_A_1635_21#_c_1532_n 0.0167184f $X=10.02 $Y=2.325
+ $X2=0 $Y2=0
cc_858 N_A_864_255#_c_1149_n N_A_1635_21#_c_1532_n 0.01314f $X=10.105 $Y=2.41
+ $X2=0 $Y2=0
cc_859 N_A_864_255#_M1006_g N_A_1635_21#_c_1527_n 0.00110762f $X=10.75 $Y=0.785
+ $X2=0 $Y2=0
cc_860 N_A_864_255#_c_1132_n N_A_1635_21#_c_1533_n 0.023213f $X=9.935 $Y=1.645
+ $X2=0 $Y2=0
cc_861 N_A_864_255#_c_1132_n N_A_1635_21#_c_1534_n 0.00741488f $X=9.935 $Y=1.645
+ $X2=0 $Y2=0
cc_862 N_A_864_255#_c_1133_n N_A_1635_21#_c_1534_n 2.05003e-19 $X=8.325 $Y=1.645
+ $X2=0 $Y2=0
cc_863 N_A_864_255#_c_1135_n N_A_1635_21#_c_1534_n 0.00226456f $X=8.16 $Y=1.72
+ $X2=0 $Y2=0
cc_864 N_A_864_255#_M1006_g N_A_1635_21#_c_1528_n 0.00517184f $X=10.75 $Y=0.785
+ $X2=0 $Y2=0
cc_865 N_A_864_255#_M1006_g N_CLK_M1008_g 0.0282234f $X=10.75 $Y=0.785 $X2=0
+ $Y2=0
cc_866 N_A_864_255#_c_1134_n N_CLK_M1008_g 0.0135117f $X=11.132 $Y=1.672 $X2=0
+ $Y2=0
cc_867 N_A_864_255#_M1002_g N_CLK_M1020_g 0.0328257f $X=10.755 $Y=2.465 $X2=0
+ $Y2=0
cc_868 N_A_864_255#_c_1134_n N_CLK_M1020_g 0.00459986f $X=11.132 $Y=1.672 $X2=0
+ $Y2=0
cc_869 N_A_864_255#_c_1150_n N_CLK_M1020_g 0.029339f $X=11.132 $Y=2.325 $X2=0
+ $Y2=0
cc_870 N_A_864_255#_c_1277_p N_CLK_M1020_g 0.00624229f $X=11.375 $Y=2.66 $X2=0
+ $Y2=0
cc_871 N_A_864_255#_c_1278_p N_CLK_M1020_g 0.00838452f $X=11.132 $Y=2.41 $X2=0
+ $Y2=0
cc_872 N_A_864_255#_c_1153_n N_CLK_M1020_g 0.00685311f $X=11.555 $Y=2.765 $X2=0
+ $Y2=0
cc_873 N_A_864_255#_c_1134_n N_CLK_c_1638_n 0.0159706f $X=11.132 $Y=1.672 $X2=0
+ $Y2=0
cc_874 N_A_864_255#_c_1134_n N_CLK_c_1639_n 0.00417528f $X=11.132 $Y=1.672 $X2=0
+ $Y2=0
cc_875 N_A_864_255#_c_1136_n N_CLK_c_1639_n 0.0213932f $X=10.89 $Y=1.51 $X2=0
+ $Y2=0
cc_876 N_A_864_255#_c_1134_n N_CLK_c_1640_n 6.51906e-19 $X=11.132 $Y=1.672 $X2=0
+ $Y2=0
cc_877 N_A_864_255#_M1020_d N_CLK_c_1641_n 0.00796345f $X=11.415 $Y=1.835 $X2=0
+ $Y2=0
cc_878 N_A_864_255#_c_1134_n N_CLK_c_1641_n 0.0295074f $X=11.132 $Y=1.672 $X2=0
+ $Y2=0
cc_879 N_A_864_255#_c_1150_n N_CLK_c_1641_n 0.0343805f $X=11.132 $Y=2.325 $X2=0
+ $Y2=0
cc_880 N_A_864_255#_c_1153_n N_CLK_c_1641_n 0.00742316f $X=11.555 $Y=2.765 $X2=0
+ $Y2=0
cc_881 N_A_864_255#_c_1150_n N_VPWR_M1002_d 0.00194695f $X=11.132 $Y=2.325 $X2=0
+ $Y2=0
cc_882 N_A_864_255#_c_1278_p N_VPWR_M1002_d 0.00534194f $X=11.132 $Y=2.41 $X2=0
+ $Y2=0
cc_883 N_A_864_255#_M1001_g N_VPWR_c_1773_n 0.00678956f $X=4.395 $Y=2.525 $X2=0
+ $Y2=0
cc_884 N_A_864_255#_c_1138_n N_VPWR_c_1773_n 0.0256572f $X=7.075 $Y=3.15 $X2=0
+ $Y2=0
cc_885 N_A_864_255#_c_1138_n N_VPWR_c_1774_n 0.0253374f $X=7.075 $Y=3.15 $X2=0
+ $Y2=0
cc_886 N_A_864_255#_M1009_g N_VPWR_c_1774_n 0.00581309f $X=7.15 $Y=2.315 $X2=0
+ $Y2=0
cc_887 N_A_864_255#_M1002_g N_VPWR_c_1775_n 0.00749395f $X=10.755 $Y=2.465 $X2=0
+ $Y2=0
cc_888 N_A_864_255#_c_1148_n N_VPWR_c_1775_n 0.00473761f $X=10.805 $Y=2.41 $X2=0
+ $Y2=0
cc_889 N_A_864_255#_c_1149_n N_VPWR_c_1775_n 0.0128433f $X=10.105 $Y=2.41 $X2=0
+ $Y2=0
cc_890 N_A_864_255#_M1002_g N_VPWR_c_1776_n 0.0153983f $X=10.755 $Y=2.465 $X2=0
+ $Y2=0
cc_891 N_A_864_255#_c_1278_p N_VPWR_c_1776_n 0.0223431f $X=11.132 $Y=2.41 $X2=0
+ $Y2=0
cc_892 N_A_864_255#_c_1153_n N_VPWR_c_1776_n 0.0217248f $X=11.555 $Y=2.765 $X2=0
+ $Y2=0
cc_893 N_A_864_255#_M1002_g N_VPWR_c_1784_n 0.00486043f $X=10.755 $Y=2.465 $X2=0
+ $Y2=0
cc_894 N_A_864_255#_c_1139_n N_VPWR_c_1787_n 0.0190557f $X=4.47 $Y=3.15 $X2=0
+ $Y2=0
cc_895 N_A_864_255#_c_1138_n N_VPWR_c_1788_n 0.0345146f $X=7.075 $Y=3.15 $X2=0
+ $Y2=0
cc_896 N_A_864_255#_c_1153_n N_VPWR_c_1789_n 0.0140235f $X=11.555 $Y=2.765 $X2=0
+ $Y2=0
cc_897 N_A_864_255#_c_1138_n N_VPWR_c_1794_n 0.0187969f $X=7.075 $Y=3.15 $X2=0
+ $Y2=0
cc_898 N_A_864_255#_M1020_d N_VPWR_c_1770_n 0.00232647f $X=11.415 $Y=1.835 $X2=0
+ $Y2=0
cc_899 N_A_864_255#_c_1138_n N_VPWR_c_1770_n 0.0724812f $X=7.075 $Y=3.15 $X2=0
+ $Y2=0
cc_900 N_A_864_255#_c_1139_n N_VPWR_c_1770_n 0.0094884f $X=4.47 $Y=3.15 $X2=0
+ $Y2=0
cc_901 N_A_864_255#_M1002_g N_VPWR_c_1770_n 0.00599211f $X=10.755 $Y=2.465 $X2=0
+ $Y2=0
cc_902 N_A_864_255#_c_1148_n N_VPWR_c_1770_n 0.0212343f $X=10.805 $Y=2.41 $X2=0
+ $Y2=0
cc_903 N_A_864_255#_c_1149_n N_VPWR_c_1770_n 6.93057e-19 $X=10.105 $Y=2.41 $X2=0
+ $Y2=0
cc_904 N_A_864_255#_c_1278_p N_VPWR_c_1770_n 0.00771847f $X=11.132 $Y=2.41 $X2=0
+ $Y2=0
cc_905 N_A_864_255#_c_1153_n N_VPWR_c_1770_n 0.0143844f $X=11.555 $Y=2.765 $X2=0
+ $Y2=0
cc_906 N_A_864_255#_M1001_g N_A_380_50#_c_1932_n 3.12444e-19 $X=4.395 $Y=2.525
+ $X2=0 $Y2=0
cc_907 N_A_864_255#_M1031_g N_A_380_50#_c_1932_n 0.0022481f $X=4.45 $Y=0.805
+ $X2=0 $Y2=0
cc_908 N_A_864_255#_M1001_g N_A_380_50#_c_1940_n 0.00327967f $X=4.395 $Y=2.525
+ $X2=0 $Y2=0
cc_909 N_A_864_255#_M1031_g N_A_380_50#_c_1936_n 0.00282073f $X=4.45 $Y=0.805
+ $X2=0 $Y2=0
cc_910 N_A_864_255#_M1006_g N_VGND_c_2065_n 0.00438183f $X=10.75 $Y=0.785 $X2=0
+ $Y2=0
cc_911 N_A_864_255#_M1027_g N_VGND_c_2071_n 6.694e-19 $X=7.89 $Y=0.775 $X2=0
+ $Y2=0
cc_912 N_A_864_255#_M1006_g N_VGND_c_2073_n 0.00330473f $X=10.75 $Y=0.785 $X2=0
+ $Y2=0
cc_913 N_A_864_255#_M1031_g N_VGND_c_2082_n 9.39239e-19 $X=4.45 $Y=0.805 $X2=0
+ $Y2=0
cc_914 N_A_864_255#_M1006_g N_VGND_c_2082_n 0.00430341f $X=10.75 $Y=0.785 $X2=0
+ $Y2=0
cc_915 N_A_1406_69#_c_1332_n N_A_1635_21#_M1017_g 0.0166968f $X=8.065 $Y=0.625
+ $X2=0 $Y2=0
cc_916 N_A_1406_69#_c_1334_n N_A_1635_21#_M1017_g 0.00478174f $X=8.15 $Y=1.205
+ $X2=0 $Y2=0
cc_917 N_A_1406_69#_c_1322_n N_A_1635_21#_c_1520_n 0.0103024f $X=9.33 $Y=1.125
+ $X2=0 $Y2=0
cc_918 N_A_1406_69#_c_1335_n N_A_1635_21#_c_1522_n 0.012848f $X=9.83 $Y=1.29
+ $X2=0 $Y2=0
cc_919 N_A_1406_69#_c_1334_n N_A_1635_21#_c_1523_n 0.00328963f $X=8.15 $Y=1.205
+ $X2=0 $Y2=0
cc_920 N_A_1406_69#_c_1335_n N_A_1635_21#_c_1523_n 0.00493696f $X=9.83 $Y=1.29
+ $X2=0 $Y2=0
cc_921 N_A_1406_69#_c_1336_n N_A_1635_21#_c_1523_n 8.66673e-19 $X=8.235 $Y=1.29
+ $X2=0 $Y2=0
cc_922 N_A_1406_69#_c_1335_n N_A_1635_21#_c_1524_n 0.00579209f $X=9.83 $Y=1.29
+ $X2=0 $Y2=0
cc_923 N_A_1406_69#_M1038_g N_A_1635_21#_c_1531_n 0.00674732f $X=9.69 $Y=2.88
+ $X2=0 $Y2=0
cc_924 N_A_1406_69#_M1038_g N_A_1635_21#_c_1558_n 0.00497329f $X=9.69 $Y=2.88
+ $X2=0 $Y2=0
cc_925 N_A_1406_69#_c_1322_n N_A_1635_21#_c_1525_n 0.011476f $X=9.33 $Y=1.125
+ $X2=0 $Y2=0
cc_926 N_A_1406_69#_c_1323_n N_A_1635_21#_c_1525_n 0.00548896f $X=9.615 $Y=1.2
+ $X2=0 $Y2=0
cc_927 N_A_1406_69#_c_1335_n N_A_1635_21#_c_1525_n 0.0130016f $X=9.83 $Y=1.29
+ $X2=0 $Y2=0
cc_928 N_A_1406_69#_c_1337_n N_A_1635_21#_c_1525_n 0.0118636f $X=9.915 $Y=1.205
+ $X2=0 $Y2=0
cc_929 N_A_1406_69#_c_1339_n N_A_1635_21#_c_1525_n 0.0146126f $X=10 $Y=0.73
+ $X2=0 $Y2=0
cc_930 N_A_1406_69#_M1038_g N_A_1635_21#_c_1532_n 0.0228357f $X=9.69 $Y=2.88
+ $X2=0 $Y2=0
cc_931 N_A_1406_69#_c_1322_n N_A_1635_21#_c_1526_n 5.55733e-19 $X=9.33 $Y=1.125
+ $X2=0 $Y2=0
cc_932 N_A_1406_69#_c_1338_n N_A_1635_21#_c_1527_n 0.00756892f $X=11.9 $Y=0.73
+ $X2=0 $Y2=0
cc_933 N_A_1406_69#_c_1339_n N_A_1635_21#_c_1527_n 0.0131623f $X=10 $Y=0.73
+ $X2=0 $Y2=0
cc_934 N_A_1406_69#_c_1342_n N_A_1635_21#_c_1527_n 0.00341365f $X=9.78 $Y=1.2
+ $X2=0 $Y2=0
cc_935 N_A_1406_69#_c_1322_n N_A_1635_21#_c_1528_n 0.00144479f $X=9.33 $Y=1.125
+ $X2=0 $Y2=0
cc_936 N_A_1406_69#_c_1335_n N_A_1635_21#_c_1528_n 2.53161e-19 $X=9.83 $Y=1.29
+ $X2=0 $Y2=0
cc_937 N_A_1406_69#_c_1338_n N_A_1635_21#_c_1528_n 0.00270068f $X=11.9 $Y=0.73
+ $X2=0 $Y2=0
cc_938 N_A_1406_69#_c_1339_n N_A_1635_21#_c_1528_n 0.00278863f $X=10 $Y=0.73
+ $X2=0 $Y2=0
cc_939 N_A_1406_69#_c_1342_n N_A_1635_21#_c_1528_n 0.0023655f $X=9.78 $Y=1.2
+ $X2=0 $Y2=0
cc_940 N_A_1406_69#_c_1338_n N_CLK_M1008_g 0.0147012f $X=11.9 $Y=0.73 $X2=0
+ $Y2=0
cc_941 N_A_1406_69#_c_1340_n N_CLK_M1008_g 0.00348461f $X=11.985 $Y=0.995 $X2=0
+ $Y2=0
cc_942 N_A_1406_69#_M1028_g N_CLK_c_1640_n 0.00197204f $X=12.495 $Y=2.155 $X2=0
+ $Y2=0
cc_943 N_A_1406_69#_c_1338_n N_CLK_c_1640_n 0.003407f $X=11.9 $Y=0.73 $X2=0
+ $Y2=0
cc_944 N_A_1406_69#_c_1340_n N_CLK_c_1640_n 0.00239682f $X=11.985 $Y=0.995 $X2=0
+ $Y2=0
cc_945 N_A_1406_69#_c_1341_n N_CLK_c_1640_n 0.0131692f $X=12.375 $Y=1.08 $X2=0
+ $Y2=0
cc_946 N_A_1406_69#_M1028_g N_CLK_c_1641_n 0.00245703f $X=12.495 $Y=2.155 $X2=0
+ $Y2=0
cc_947 N_A_1406_69#_c_1329_n N_CLK_c_1641_n 0.00219417f $X=12.39 $Y=1.585 $X2=0
+ $Y2=0
cc_948 N_A_1406_69#_c_1338_n N_CLK_c_1641_n 0.00546696f $X=11.9 $Y=0.73 $X2=0
+ $Y2=0
cc_949 N_A_1406_69#_c_1340_n N_CLK_c_1641_n 0.0156163f $X=11.985 $Y=0.995 $X2=0
+ $Y2=0
cc_950 N_A_1406_69#_M1011_g N_A_2431_47#_M1024_g 0.029911f $X=12.495 $Y=0.445
+ $X2=0 $Y2=0
cc_951 N_A_1406_69#_c_1340_n N_A_2431_47#_M1024_g 2.23991e-19 $X=11.985 $Y=0.995
+ $X2=0 $Y2=0
cc_952 N_A_1406_69#_c_1329_n N_A_2431_47#_M1010_g 0.0208771f $X=12.39 $Y=1.585
+ $X2=0 $Y2=0
cc_953 N_A_1406_69#_M1028_g N_A_2431_47#_c_1694_n 4.43331e-19 $X=12.495 $Y=2.155
+ $X2=0 $Y2=0
cc_954 N_A_1406_69#_M1011_g N_A_2431_47#_c_1702_n 0.00481975f $X=12.495 $Y=0.445
+ $X2=0 $Y2=0
cc_955 N_A_1406_69#_M1028_g N_A_2431_47#_c_1695_n 0.016321f $X=12.495 $Y=2.155
+ $X2=0 $Y2=0
cc_956 N_A_1406_69#_c_1329_n N_A_2431_47#_c_1695_n 0.00129934f $X=12.39 $Y=1.585
+ $X2=0 $Y2=0
cc_957 N_A_1406_69#_c_1340_n N_A_2431_47#_c_1695_n 0.0124014f $X=11.985 $Y=0.995
+ $X2=0 $Y2=0
cc_958 N_A_1406_69#_c_1329_n N_A_2431_47#_c_1696_n 0.00494327f $X=12.39 $Y=1.585
+ $X2=0 $Y2=0
cc_959 N_A_1406_69#_c_1340_n N_A_2431_47#_c_1696_n 0.0160084f $X=11.985 $Y=0.995
+ $X2=0 $Y2=0
cc_960 N_A_1406_69#_M1011_g N_A_2431_47#_c_1686_n 0.00986832f $X=12.495 $Y=0.445
+ $X2=0 $Y2=0
cc_961 N_A_1406_69#_c_1340_n N_A_2431_47#_c_1686_n 0.00671434f $X=11.985
+ $Y=0.995 $X2=0 $Y2=0
cc_962 N_A_1406_69#_M1011_g N_A_2431_47#_c_1687_n 0.00368082f $X=12.495 $Y=0.445
+ $X2=0 $Y2=0
cc_963 N_A_1406_69#_c_1328_n N_A_2431_47#_c_1687_n 0.00455766f $X=12.39 $Y=1.035
+ $X2=0 $Y2=0
cc_964 N_A_1406_69#_c_1338_n N_A_2431_47#_c_1687_n 0.0139124f $X=11.9 $Y=0.73
+ $X2=0 $Y2=0
cc_965 N_A_1406_69#_c_1340_n N_A_2431_47#_c_1687_n 0.0133932f $X=11.985 $Y=0.995
+ $X2=0 $Y2=0
cc_966 N_A_1406_69#_M1011_g N_A_2431_47#_c_1688_n 0.00423999f $X=12.495 $Y=0.445
+ $X2=0 $Y2=0
cc_967 N_A_1406_69#_c_1340_n N_A_2431_47#_c_1688_n 0.0242821f $X=11.985 $Y=0.995
+ $X2=0 $Y2=0
cc_968 N_A_1406_69#_M1011_g N_A_2431_47#_c_1689_n 0.00223315f $X=12.495 $Y=0.445
+ $X2=0 $Y2=0
cc_969 N_A_1406_69#_c_1328_n N_A_2431_47#_c_1689_n 0.00151548f $X=12.39 $Y=1.035
+ $X2=0 $Y2=0
cc_970 N_A_1406_69#_c_1340_n N_A_2431_47#_c_1689_n 0.0053936f $X=11.985 $Y=0.995
+ $X2=0 $Y2=0
cc_971 N_A_1406_69#_c_1340_n N_A_2431_47#_c_1690_n 0.0197606f $X=11.985 $Y=0.995
+ $X2=0 $Y2=0
cc_972 N_A_1406_69#_c_1341_n N_A_2431_47#_c_1690_n 0.00543695f $X=12.375 $Y=1.08
+ $X2=0 $Y2=0
cc_973 N_A_1406_69#_c_1340_n N_A_2431_47#_c_1691_n 2.71544e-19 $X=11.985
+ $Y=0.995 $X2=0 $Y2=0
cc_974 N_A_1406_69#_c_1341_n N_A_2431_47#_c_1691_n 0.0207537f $X=12.375 $Y=1.08
+ $X2=0 $Y2=0
cc_975 N_A_1406_69#_M1038_g N_VPWR_c_1775_n 0.0114001f $X=9.69 $Y=2.88 $X2=0
+ $Y2=0
cc_976 N_A_1406_69#_M1028_g N_VPWR_c_1777_n 0.0153559f $X=12.495 $Y=2.155 $X2=0
+ $Y2=0
cc_977 N_A_1406_69#_M1038_g N_VPWR_c_1782_n 0.00369389f $X=9.69 $Y=2.88 $X2=0
+ $Y2=0
cc_978 N_A_1406_69#_M1028_g N_VPWR_c_1789_n 0.00259749f $X=12.495 $Y=2.155 $X2=0
+ $Y2=0
cc_979 N_A_1406_69#_M1009_d N_VPWR_c_1770_n 0.00420488f $X=7.225 $Y=1.895 $X2=0
+ $Y2=0
cc_980 N_A_1406_69#_M1038_g N_VPWR_c_1770_n 0.00707264f $X=9.69 $Y=2.88 $X2=0
+ $Y2=0
cc_981 N_A_1406_69#_M1028_g N_VPWR_c_1770_n 0.00344639f $X=12.495 $Y=2.155 $X2=0
+ $Y2=0
cc_982 N_A_1406_69#_c_1338_n N_VGND_M1006_d 0.00966466f $X=11.9 $Y=0.73 $X2=0
+ $Y2=0
cc_983 N_A_1406_69#_c_1332_n N_VGND_c_2064_n 0.038876f $X=8.065 $Y=0.625 $X2=0
+ $Y2=0
cc_984 N_A_1406_69#_c_1334_n N_VGND_c_2064_n 0.00170602f $X=8.15 $Y=1.205 $X2=0
+ $Y2=0
cc_985 N_A_1406_69#_c_1335_n N_VGND_c_2064_n 0.0166618f $X=9.83 $Y=1.29 $X2=0
+ $Y2=0
cc_986 N_A_1406_69#_c_1338_n N_VGND_c_2065_n 0.0249306f $X=11.9 $Y=0.73 $X2=0
+ $Y2=0
cc_987 N_A_1406_69#_M1011_g N_VGND_c_2066_n 0.00435875f $X=12.495 $Y=0.445 $X2=0
+ $Y2=0
cc_988 N_A_1406_69#_c_1330_n N_VGND_c_2071_n 0.00835105f $X=7.09 $Y=0.925 $X2=0
+ $Y2=0
cc_989 N_A_1406_69#_c_1332_n N_VGND_c_2071_n 0.0517156f $X=8.065 $Y=0.625 $X2=0
+ $Y2=0
cc_990 N_A_1406_69#_c_1338_n N_VGND_c_2073_n 0.0123458f $X=11.9 $Y=0.73 $X2=0
+ $Y2=0
cc_991 N_A_1406_69#_M1011_g N_VGND_c_2077_n 0.00415809f $X=12.495 $Y=0.445 $X2=0
+ $Y2=0
cc_992 N_A_1406_69#_c_1338_n N_VGND_c_2077_n 0.0142494f $X=11.9 $Y=0.73 $X2=0
+ $Y2=0
cc_993 N_A_1406_69#_c_1322_n N_VGND_c_2082_n 7.82699e-19 $X=9.33 $Y=1.125 $X2=0
+ $Y2=0
cc_994 N_A_1406_69#_M1011_g N_VGND_c_2082_n 0.00723931f $X=12.495 $Y=0.445 $X2=0
+ $Y2=0
cc_995 N_A_1406_69#_c_1330_n N_VGND_c_2082_n 0.00625229f $X=7.09 $Y=0.925 $X2=0
+ $Y2=0
cc_996 N_A_1406_69#_c_1332_n N_VGND_c_2082_n 0.039273f $X=8.065 $Y=0.625 $X2=0
+ $Y2=0
cc_997 N_A_1406_69#_c_1338_n N_VGND_c_2082_n 0.0467133f $X=11.9 $Y=0.73 $X2=0
+ $Y2=0
cc_998 N_A_1406_69#_c_1332_n A_1593_113# 3.28039e-19 $X=8.065 $Y=0.625 $X2=-0.19
+ $Y2=-0.245
cc_999 N_A_1406_69#_c_1334_n A_1593_113# 6.58248e-19 $X=8.15 $Y=1.205 $X2=-0.19
+ $Y2=-0.245
cc_1000 N_A_1635_21#_c_1558_n N_VPWR_c_1775_n 0.0164138f $X=9.585 $Y=2.97 $X2=0
+ $Y2=0
cc_1001 N_A_1635_21#_c_1532_n N_VPWR_c_1775_n 0.0115444f $X=9.67 $Y=2.865 $X2=0
+ $Y2=0
cc_1002 N_A_1635_21#_c_1558_n N_VPWR_c_1782_n 0.0257432f $X=9.585 $Y=2.97 $X2=0
+ $Y2=0
cc_1003 N_A_1635_21#_M1035_g N_VPWR_c_1794_n 0.00350055f $X=8.36 $Y=2.88 $X2=0
+ $Y2=0
cc_1004 N_A_1635_21#_M1035_g N_VPWR_c_1795_n 0.0116953f $X=8.36 $Y=2.88 $X2=0
+ $Y2=0
cc_1005 N_A_1635_21#_M1014_d N_VPWR_c_1770_n 0.00222771f $X=9.335 $Y=2.67 $X2=0
+ $Y2=0
cc_1006 N_A_1635_21#_M1035_g N_VPWR_c_1770_n 0.00452722f $X=8.36 $Y=2.88 $X2=0
+ $Y2=0
cc_1007 N_A_1635_21#_c_1558_n N_VPWR_c_1770_n 0.0160875f $X=9.585 $Y=2.97 $X2=0
+ $Y2=0
cc_1008 N_A_1635_21#_M1017_g N_VGND_c_2064_n 0.00741095f $X=8.25 $Y=0.775 $X2=0
+ $Y2=0
cc_1009 N_A_1635_21#_c_1520_n N_VGND_c_2064_n 0.0256773f $X=9.78 $Y=0.18 $X2=0
+ $Y2=0
cc_1010 N_A_1635_21#_c_1522_n N_VGND_c_2064_n 0.00583476f $X=8.535 $Y=1.17 $X2=0
+ $Y2=0
cc_1011 N_A_1635_21#_c_1525_n N_VGND_c_2064_n 0.0142015f $X=9.545 $Y=0.805 $X2=0
+ $Y2=0
cc_1012 N_A_1635_21#_c_1526_n N_VGND_c_2064_n 0.00822729f $X=9.66 $Y=0.365 $X2=0
+ $Y2=0
cc_1013 N_A_1635_21#_c_1521_n N_VGND_c_2071_n 0.0104146f $X=8.325 $Y=0.18 $X2=0
+ $Y2=0
cc_1014 N_A_1635_21#_c_1520_n N_VGND_c_2073_n 0.0362227f $X=9.78 $Y=0.18 $X2=0
+ $Y2=0
cc_1015 N_A_1635_21#_c_1526_n N_VGND_c_2073_n 0.0191579f $X=9.66 $Y=0.365 $X2=0
+ $Y2=0
cc_1016 N_A_1635_21#_c_1527_n N_VGND_c_2073_n 0.0284865f $X=9.945 $Y=0.35 $X2=0
+ $Y2=0
cc_1017 N_A_1635_21#_c_1520_n N_VGND_c_2082_n 0.043107f $X=9.78 $Y=0.18 $X2=0
+ $Y2=0
cc_1018 N_A_1635_21#_c_1521_n N_VGND_c_2082_n 0.00939353f $X=8.325 $Y=0.18 $X2=0
+ $Y2=0
cc_1019 N_A_1635_21#_c_1526_n N_VGND_c_2082_n 0.00961889f $X=9.66 $Y=0.365 $X2=0
+ $Y2=0
cc_1020 N_A_1635_21#_c_1527_n N_VGND_c_2082_n 0.0149973f $X=9.945 $Y=0.35 $X2=0
+ $Y2=0
cc_1021 N_A_1635_21#_c_1528_n N_VGND_c_2082_n 0.0100496f $X=9.945 $Y=0.18 $X2=0
+ $Y2=0
cc_1022 N_CLK_c_1641_n N_A_2431_47#_c_1694_n 0.0513631f $X=11.805 $Y=1.51 $X2=0
+ $Y2=0
cc_1023 N_CLK_c_1641_n N_A_2431_47#_c_1696_n 0.0152191f $X=11.805 $Y=1.51 $X2=0
+ $Y2=0
cc_1024 N_CLK_M1008_g N_A_2431_47#_c_1689_n 0.00405327f $X=11.34 $Y=0.785 $X2=0
+ $Y2=0
cc_1025 N_CLK_M1020_g N_VPWR_c_1776_n 0.00861626f $X=11.34 $Y=2.465 $X2=0 $Y2=0
cc_1026 N_CLK_M1020_g N_VPWR_c_1789_n 0.00417974f $X=11.34 $Y=2.465 $X2=0 $Y2=0
cc_1027 N_CLK_M1020_g N_VPWR_c_1770_n 0.00746349f $X=11.34 $Y=2.465 $X2=0 $Y2=0
cc_1028 N_CLK_c_1641_n N_VPWR_c_1770_n 0.0113624f $X=11.805 $Y=1.51 $X2=0 $Y2=0
cc_1029 N_CLK_M1008_g N_VGND_c_2065_n 0.00438183f $X=11.34 $Y=0.785 $X2=0 $Y2=0
cc_1030 N_CLK_M1008_g N_VGND_c_2077_n 0.00330473f $X=11.34 $Y=0.785 $X2=0 $Y2=0
cc_1031 N_CLK_M1008_g N_VGND_c_2082_n 0.00435988f $X=11.34 $Y=0.785 $X2=0 $Y2=0
cc_1032 N_A_2431_47#_c_1695_n N_VPWR_M1028_d 9.77978e-19 $X=12.72 $Y=1.76 $X2=0
+ $Y2=0
cc_1033 N_A_2431_47#_c_1690_n N_VPWR_M1028_d 0.00169314f $X=12.945 $Y=1.41 $X2=0
+ $Y2=0
cc_1034 N_A_2431_47#_M1010_g N_VPWR_c_1777_n 0.0206387f $X=13.005 $Y=2.465 $X2=0
+ $Y2=0
cc_1035 N_A_2431_47#_M1029_g N_VPWR_c_1777_n 8.36898e-19 $X=13.435 $Y=2.465
+ $X2=0 $Y2=0
cc_1036 N_A_2431_47#_c_1694_n N_VPWR_c_1777_n 0.0192815f $X=12.28 $Y=1.98 $X2=0
+ $Y2=0
cc_1037 N_A_2431_47#_c_1695_n N_VPWR_c_1777_n 0.00931595f $X=12.72 $Y=1.76 $X2=0
+ $Y2=0
cc_1038 N_A_2431_47#_c_1690_n N_VPWR_c_1777_n 0.0151204f $X=12.945 $Y=1.41 $X2=0
+ $Y2=0
cc_1039 N_A_2431_47#_c_1691_n N_VPWR_c_1777_n 4.499e-19 $X=13.435 $Y=1.41 $X2=0
+ $Y2=0
cc_1040 N_A_2431_47#_M1029_g N_VPWR_c_1779_n 0.00742903f $X=13.435 $Y=2.465
+ $X2=0 $Y2=0
cc_1041 N_A_2431_47#_M1010_g N_VPWR_c_1790_n 0.00525069f $X=13.005 $Y=2.465
+ $X2=0 $Y2=0
cc_1042 N_A_2431_47#_M1029_g N_VPWR_c_1790_n 0.00564131f $X=13.435 $Y=2.465
+ $X2=0 $Y2=0
cc_1043 N_A_2431_47#_M1010_g N_VPWR_c_1770_n 0.00886509f $X=13.005 $Y=2.465
+ $X2=0 $Y2=0
cc_1044 N_A_2431_47#_M1029_g N_VPWR_c_1770_n 0.0110509f $X=13.435 $Y=2.465 $X2=0
+ $Y2=0
cc_1045 N_A_2431_47#_c_1694_n N_VPWR_c_1770_n 0.00784141f $X=12.28 $Y=1.98 $X2=0
+ $Y2=0
cc_1046 N_A_2431_47#_M1041_g N_Q_c_2038_n 0.00773436f $X=13.435 $Y=0.655 $X2=0
+ $Y2=0
cc_1047 N_A_2431_47#_M1041_g N_Q_c_2039_n 0.00129524f $X=13.435 $Y=0.655 $X2=0
+ $Y2=0
cc_1048 N_A_2431_47#_c_1691_n N_Q_c_2039_n 0.00131892f $X=13.435 $Y=1.41 $X2=0
+ $Y2=0
cc_1049 N_A_2431_47#_M1010_g N_Q_c_2036_n 0.00142104f $X=13.005 $Y=2.465 $X2=0
+ $Y2=0
cc_1050 N_A_2431_47#_M1029_g N_Q_c_2036_n 0.00393417f $X=13.435 $Y=2.465 $X2=0
+ $Y2=0
cc_1051 N_A_2431_47#_c_1690_n N_Q_c_2036_n 0.00565781f $X=12.945 $Y=1.41 $X2=0
+ $Y2=0
cc_1052 N_A_2431_47#_c_1691_n N_Q_c_2036_n 0.00131892f $X=13.435 $Y=1.41 $X2=0
+ $Y2=0
cc_1053 N_A_2431_47#_M1024_g N_Q_c_2035_n 0.00125464f $X=13.005 $Y=0.655 $X2=0
+ $Y2=0
cc_1054 N_A_2431_47#_M1010_g N_Q_c_2035_n 0.00140799f $X=13.005 $Y=2.465 $X2=0
+ $Y2=0
cc_1055 N_A_2431_47#_M1041_g N_Q_c_2035_n 0.0074857f $X=13.435 $Y=0.655 $X2=0
+ $Y2=0
cc_1056 N_A_2431_47#_M1029_g N_Q_c_2035_n 0.00842182f $X=13.435 $Y=2.465 $X2=0
+ $Y2=0
cc_1057 N_A_2431_47#_c_1688_n N_Q_c_2035_n 0.00966485f $X=12.832 $Y=1.245 $X2=0
+ $Y2=0
cc_1058 N_A_2431_47#_c_1690_n N_Q_c_2035_n 0.0330383f $X=12.945 $Y=1.41 $X2=0
+ $Y2=0
cc_1059 N_A_2431_47#_c_1691_n N_Q_c_2035_n 0.025808f $X=13.435 $Y=1.41 $X2=0
+ $Y2=0
cc_1060 N_A_2431_47#_M1029_g Q 0.0135782f $X=13.435 $Y=2.465 $X2=0 $Y2=0
cc_1061 N_A_2431_47#_c_1686_n N_VGND_M1011_d 0.00406008f $X=12.72 $Y=0.73 $X2=0
+ $Y2=0
cc_1062 N_A_2431_47#_c_1688_n N_VGND_M1011_d 0.00341772f $X=12.832 $Y=1.245
+ $X2=0 $Y2=0
cc_1063 N_A_2431_47#_M1024_g N_VGND_c_2066_n 0.00616302f $X=13.005 $Y=0.655
+ $X2=0 $Y2=0
cc_1064 N_A_2431_47#_M1041_g N_VGND_c_2066_n 4.66399e-19 $X=13.435 $Y=0.655
+ $X2=0 $Y2=0
cc_1065 N_A_2431_47#_c_1686_n N_VGND_c_2066_n 0.0210712f $X=12.72 $Y=0.73 $X2=0
+ $Y2=0
cc_1066 N_A_2431_47#_M1041_g N_VGND_c_2068_n 0.00684158f $X=13.435 $Y=0.655
+ $X2=0 $Y2=0
cc_1067 N_A_2431_47#_c_1686_n N_VGND_c_2077_n 0.00240763f $X=12.72 $Y=0.73 $X2=0
+ $Y2=0
cc_1068 N_A_2431_47#_c_1689_n N_VGND_c_2077_n 0.0172428f $X=12.28 $Y=0.38 $X2=0
+ $Y2=0
cc_1069 N_A_2431_47#_M1024_g N_VGND_c_2078_n 0.00525069f $X=13.005 $Y=0.655
+ $X2=0 $Y2=0
cc_1070 N_A_2431_47#_M1041_g N_VGND_c_2078_n 0.00564131f $X=13.435 $Y=0.655
+ $X2=0 $Y2=0
cc_1071 N_A_2431_47#_M1011_s N_VGND_c_2082_n 0.00215867f $X=12.155 $Y=0.235
+ $X2=0 $Y2=0
cc_1072 N_A_2431_47#_M1024_g N_VGND_c_2082_n 0.00886509f $X=13.005 $Y=0.655
+ $X2=0 $Y2=0
cc_1073 N_A_2431_47#_M1041_g N_VGND_c_2082_n 0.0110509f $X=13.435 $Y=0.655 $X2=0
+ $Y2=0
cc_1074 N_A_2431_47#_c_1686_n N_VGND_c_2082_n 0.00575328f $X=12.72 $Y=0.73 $X2=0
+ $Y2=0
cc_1075 N_A_2431_47#_c_1689_n N_VGND_c_2082_n 0.0121041f $X=12.28 $Y=0.38 $X2=0
+ $Y2=0
cc_1076 N_VPWR_M1012_d N_A_380_50#_c_1937_n 0.00426912f $X=2.92 $Y=2.34 $X2=0
+ $Y2=0
cc_1077 N_VPWR_c_1772_n N_A_380_50#_c_1937_n 0.0256659f $X=3.135 $Y=2.765 $X2=0
+ $Y2=0
cc_1078 N_VPWR_c_1770_n N_A_380_50#_c_1937_n 0.0256306f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1079 N_VPWR_c_1771_n N_A_380_50#_c_1939_n 0.0111757f $X=1.37 $Y=2.485 $X2=0
+ $Y2=0
cc_1080 N_VPWR_c_1772_n N_A_380_50#_c_1939_n 0.00475219f $X=3.135 $Y=2.765 $X2=0
+ $Y2=0
cc_1081 N_VPWR_c_1786_n N_A_380_50#_c_1939_n 0.0157949f $X=2.97 $Y=3.33 $X2=0
+ $Y2=0
cc_1082 N_VPWR_c_1770_n N_A_380_50#_c_1939_n 0.0120401f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1083 N_VPWR_c_1772_n N_A_380_50#_c_1940_n 0.0220038f $X=3.135 $Y=2.765 $X2=0
+ $Y2=0
cc_1084 N_VPWR_c_1787_n N_A_380_50#_c_1940_n 0.0159799f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_1085 N_VPWR_c_1770_n N_A_380_50#_c_1940_n 0.0153628f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1086 N_VPWR_c_1770_n A_1569_534# 0.00513015f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1087 N_VPWR_c_1770_n N_Q_M1010_s 0.00345315f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1088 N_VPWR_c_1779_n N_Q_c_2036_n 0.0463129f $X=13.65 $Y=1.98 $X2=0 $Y2=0
cc_1089 N_VPWR_c_1790_n Q 0.0153611f $X=13.545 $Y=3.33 $X2=0 $Y2=0
cc_1090 N_VPWR_c_1770_n Q 0.00989321f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1091 N_A_380_50#_c_1937_n A_490_468# 0.00421169f $X=3.455 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_1092 N_A_380_50#_c_1931_n N_VGND_c_2062_n 0.00320548f $X=3.455 $Y=0.92 $X2=0
+ $Y2=0
cc_1093 N_A_380_50#_c_1933_n N_VGND_c_2062_n 0.00439668f $X=3.955 $Y=0.92 $X2=0
+ $Y2=0
cc_1094 N_A_380_50#_c_1935_n N_VGND_c_2062_n 0.0201661f $X=3.567 $Y=0.92 $X2=0
+ $Y2=0
cc_1095 N_A_380_50#_c_1936_n N_VGND_c_2062_n 0.00170514f $X=4.13 $Y=0.805 $X2=0
+ $Y2=0
cc_1096 N_A_380_50#_c_1936_n N_VGND_c_2069_n 0.00473837f $X=4.13 $Y=0.805 $X2=0
+ $Y2=0
cc_1097 N_A_380_50#_c_1931_n N_VGND_c_2082_n 0.00737337f $X=3.455 $Y=0.92 $X2=0
+ $Y2=0
cc_1098 N_A_380_50#_c_1933_n N_VGND_c_2082_n 0.00646725f $X=3.955 $Y=0.92 $X2=0
+ $Y2=0
cc_1099 N_A_380_50#_c_1935_n N_VGND_c_2082_n 8.24991e-19 $X=3.567 $Y=0.92 $X2=0
+ $Y2=0
cc_1100 N_A_380_50#_c_1936_n N_VGND_c_2082_n 0.00657042f $X=4.13 $Y=0.805 $X2=0
+ $Y2=0
cc_1101 N_A_380_50#_M1033_d N_noxref_24_c_2204_n 0.00989114f $X=1.9 $Y=0.25
+ $X2=0 $Y2=0
cc_1102 N_A_380_50#_c_1931_n N_noxref_24_c_2204_n 0.0150529f $X=3.455 $Y=0.92
+ $X2=0 $Y2=0
cc_1103 N_A_380_50#_c_1934_n N_noxref_24_c_2204_n 0.0240309f $X=2.155 $Y=0.7
+ $X2=0 $Y2=0
cc_1104 N_A_380_50#_c_1934_n N_noxref_24_c_2205_n 5.95629e-19 $X=2.155 $Y=0.7
+ $X2=0 $Y2=0
cc_1105 N_A_380_50#_c_1931_n N_noxref_24_c_2206_n 0.0203788f $X=3.455 $Y=0.92
+ $X2=0 $Y2=0
cc_1106 N_A_380_50#_c_1934_n N_noxref_24_c_2206_n 0.00178689f $X=2.155 $Y=0.7
+ $X2=0 $Y2=0
cc_1107 N_Q_c_2038_n N_VGND_c_2068_n 0.0310208f $X=13.22 $Y=0.42 $X2=0 $Y2=0
cc_1108 N_Q_c_2038_n N_VGND_c_2078_n 0.0153611f $X=13.22 $Y=0.42 $X2=0 $Y2=0
cc_1109 N_Q_M1024_d N_VGND_c_2082_n 0.00345315f $X=13.08 $Y=0.235 $X2=0 $Y2=0
cc_1110 N_Q_c_2038_n N_VGND_c_2082_n 0.00989321f $X=13.22 $Y=0.42 $X2=0 $Y2=0
cc_1111 N_VGND_c_2076_n N_noxref_24_c_2204_n 0.0838299f $X=3.405 $Y=0 $X2=0
+ $Y2=0
cc_1112 N_VGND_c_2082_n N_noxref_24_c_2204_n 0.0540533f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1113 N_VGND_c_2061_n N_noxref_24_c_2205_n 0.0277209f $X=0.73 $Y=0.565 $X2=0
+ $Y2=0
cc_1114 N_VGND_c_2076_n N_noxref_24_c_2205_n 0.0189903f $X=3.405 $Y=0 $X2=0
+ $Y2=0
cc_1115 N_VGND_c_2082_n N_noxref_24_c_2205_n 0.0123641f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1116 N_VGND_c_2062_n N_noxref_24_c_2206_n 0.0198933f $X=3.57 $Y=0.55 $X2=0
+ $Y2=0
cc_1117 N_VGND_c_2076_n N_noxref_24_c_2206_n 0.021233f $X=3.405 $Y=0 $X2=0 $Y2=0
cc_1118 N_VGND_c_2082_n N_noxref_24_c_2206_n 0.0124747f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1119 N_noxref_24_c_2204_n noxref_25 0.00458445f $X=2.895 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_1120 N_noxref_24_c_2204_n noxref_26 0.00154019f $X=2.895 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
