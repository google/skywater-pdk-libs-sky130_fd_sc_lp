* File: sky130_fd_sc_lp__invlp_0.pex.spice
* Created: Fri Aug 28 10:39:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INVLP_0%A 3 7 9 13 17 20 22 23 24 25 26 37
r36 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.455
+ $Y=1.345 $X2=0.455 $Y2=1.345
r37 25 26 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=2.035
r38 25 38 5.39078 $w=7.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=1.345
r39 24 38 0.842309 $w=7.08e-07 $l=5e-08 $layer=LI1_cond $X=0.48 $Y=1.295
+ $X2=0.48 $Y2=1.345
r40 21 37 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.455 $Y=1.685
+ $X2=0.455 $Y2=1.345
r41 21 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.455 $Y=1.685
+ $X2=0.455 $Y2=1.85
r42 19 37 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.455 $Y=1.33
+ $X2=0.455 $Y2=1.345
r43 19 20 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=0.455 $Y=1.33
+ $X2=0.455 $Y2=1.255
r44 15 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.935 $Y=1.33
+ $X2=0.935 $Y2=1.255
r45 15 17 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.935 $Y=1.33
+ $X2=0.935 $Y2=2.66
r46 11 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.935 $Y=1.18
+ $X2=0.935 $Y2=1.255
r47 11 13 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.935 $Y=1.18
+ $X2=0.935 $Y2=0.67
r48 10 20 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.62 $Y=1.255
+ $X2=0.455 $Y2=1.255
r49 9 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.86 $Y=1.255
+ $X2=0.935 $Y2=1.255
r50 9 10 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.86 $Y=1.255
+ $X2=0.62 $Y2=1.255
r51 7 22 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.545 $Y=2.66
+ $X2=0.545 $Y2=1.85
r52 1 20 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.545 $Y=1.18
+ $X2=0.455 $Y2=1.255
r53 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.545 $Y=1.18
+ $X2=0.545 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_0%VPWR 1 4 6 8 12 13
r16 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r17 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r18 10 16 4.62984 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=0.495 $Y=3.33
+ $X2=0.247 $Y2=3.33
r19 10 12 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.495 $Y=3.33
+ $X2=1.2 $Y2=3.33
r20 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33 $X2=1.2
+ $Y2=3.33
r21 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r22 4 16 3.13634 $w=3.3e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.247 $Y2=3.33
r23 4 6 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.33 $Y=3.245 $X2=0.33
+ $Y2=2.485
r24 1 6 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=2.34 $X2=0.33 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_0%Y 1 2 7 8 9 10 11 12 13 27 51
r18 27 47 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.2 $Y=0.925 $X2=1.2
+ $Y2=0.9
r19 12 51 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.15 $Y=2.485 $X2=1.15
+ $Y2=2.405
r20 12 51 0.104768 $w=3.28e-07 $l=3e-09 $layer=LI1_cond $X=1.15 $Y=2.402
+ $X2=1.15 $Y2=2.405
r21 12 13 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.15 $Y=2.485
+ $X2=1.15 $Y2=2.775
r22 11 12 10.2753 $w=3.98e-07 $l=2.85e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.32
r23 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.2
+ $Y2=2.035
r24 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.665
r25 8 47 2.11807 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.15 $Y=0.87 $X2=1.15
+ $Y2=0.9
r26 8 45 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.15 $Y=0.87 $X2=1.15
+ $Y2=0.67
r27 8 9 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.2 $Y=0.955 $X2=1.2
+ $Y2=1.295
r28 8 27 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=1.2 $Y=0.955 $X2=1.2
+ $Y2=0.925
r29 7 45 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.15 $Y=0.555
+ $X2=1.15 $Y2=0.67
r30 2 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.34 $X2=1.15 $Y2=2.485
r31 1 45 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.46 $X2=1.15 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_0%VGND 1 4 6 8 12 13
r15 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r16 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r17 10 16 4.62984 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=0.495 $Y=0 $X2=0.247
+ $Y2=0
r18 10 12 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.495 $Y=0 $X2=1.2
+ $Y2=0
r19 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r20 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r21 4 16 3.13634 $w=3.3e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.247 $Y2=0
r22 4 6 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.33 $Y2=0.67
r23 1 6 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.46 $X2=0.33 $Y2=0.67
.ends

