* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 X a_102_53# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_753_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VGND a_102_53# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_645_367# A2 a_753_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR B1 a_102_53# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR a_102_53# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND A3 a_465_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_102_53# A4 a_573_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_573_367# A3 a_645_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_465_49# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VGND A1 a_465_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_102_53# B1 a_465_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_465_49# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 X a_102_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
