* NGSPICE file created from sky130_fd_sc_lp__dlxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlxtp_1 D GATE VGND VNB VPB VPWR Q
M1000 VPWR a_196_425# a_317_461# VPB phighvt w=640000u l=150000u
+  ad=1.2717e+12p pd=1.084e+07u as=1.696e+11p ps=1.81e+06u
M1001 VGND a_196_425# a_317_461# VNB nshort w=420000u l=150000u
+  ad=7.329e+11p pd=7.47e+06u as=1.113e+11p ps=1.37e+06u
M1002 VGND a_733_99# a_691_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1003 a_530_125# a_27_425# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_701_419# a_317_461# a_596_419# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.158e+11p ps=2.03e+06u
M1005 a_691_125# a_196_425# a_596_419# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.239e+11p ps=1.43e+06u
M1006 VPWR a_733_99# a_701_419# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR D a_27_425# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1008 VGND D a_27_425# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 a_196_425# GATE VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1010 a_524_419# a_27_425# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1011 Q a_733_99# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1012 a_596_419# a_196_425# a_524_419# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_733_99# a_596_419# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1014 Q a_733_99# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1015 a_196_425# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1016 a_733_99# a_596_419# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1017 a_596_419# a_317_461# a_530_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

