* File: sky130_fd_sc_lp__o221ai_2.pxi.spice
* Created: Wed Sep  2 10:19:11 2020
* 
x_PM_SKY130_FD_SC_LP__O221AI_2%C1 N_C1_c_90_n N_C1_M1002_g N_C1_M1004_g
+ N_C1_c_92_n N_C1_M1005_g N_C1_M1015_g C1 C1 N_C1_c_95_n
+ PM_SKY130_FD_SC_LP__O221AI_2%C1
x_PM_SKY130_FD_SC_LP__O221AI_2%B1 N_B1_M1003_g N_B1_M1001_g N_B1_M1013_g
+ N_B1_M1010_g N_B1_c_138_n N_B1_c_132_n N_B1_c_133_n N_B1_c_134_n B1 B1
+ N_B1_c_135_n PM_SKY130_FD_SC_LP__O221AI_2%B1
x_PM_SKY130_FD_SC_LP__O221AI_2%B2 N_B2_c_226_n N_B2_M1006_g N_B2_M1007_g
+ N_B2_c_228_n N_B2_M1014_g N_B2_M1019_g B2 N_B2_c_231_n
+ PM_SKY130_FD_SC_LP__O221AI_2%B2
x_PM_SKY130_FD_SC_LP__O221AI_2%A1 N_A1_M1011_g N_A1_M1000_g N_A1_c_283_n
+ N_A1_M1012_g N_A1_M1016_g N_A1_c_285_n N_A1_c_286_n N_A1_c_293_n N_A1_c_294_n
+ A1 A1 N_A1_c_288_n N_A1_c_296_n A1 PM_SKY130_FD_SC_LP__O221AI_2%A1
x_PM_SKY130_FD_SC_LP__O221AI_2%A2 N_A2_c_367_n N_A2_M1009_g N_A2_M1008_g
+ N_A2_c_369_n N_A2_M1017_g N_A2_M1018_g A2 A2 N_A2_c_372_n
+ PM_SKY130_FD_SC_LP__O221AI_2%A2
x_PM_SKY130_FD_SC_LP__O221AI_2%VPWR N_VPWR_M1004_d N_VPWR_M1015_d N_VPWR_M1013_d
+ N_VPWR_M1016_d N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n
+ N_VPWR_c_427_n N_VPWR_c_428_n VPWR N_VPWR_c_429_n N_VPWR_c_430_n
+ N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_422_n
+ PM_SKY130_FD_SC_LP__O221AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O221AI_2%Y N_Y_M1002_d N_Y_M1004_s N_Y_M1007_s N_Y_M1008_s
+ N_Y_c_501_n N_Y_c_511_n N_Y_c_500_n N_Y_c_517_n N_Y_c_520_n N_Y_c_534_n Y Y Y
+ Y Y N_Y_c_504_n PM_SKY130_FD_SC_LP__O221AI_2%Y
x_PM_SKY130_FD_SC_LP__O221AI_2%A_388_367# N_A_388_367#_M1001_s
+ N_A_388_367#_M1019_d N_A_388_367#_c_581_n N_A_388_367#_c_567_n
+ N_A_388_367#_c_576_n N_A_388_367#_c_568_n
+ PM_SKY130_FD_SC_LP__O221AI_2%A_388_367#
x_PM_SKY130_FD_SC_LP__O221AI_2%A_794_367# N_A_794_367#_M1000_s
+ N_A_794_367#_M1018_d N_A_794_367#_c_599_n N_A_794_367#_c_588_n
+ N_A_794_367#_c_594_n N_A_794_367#_c_596_n N_A_794_367#_c_587_n
+ PM_SKY130_FD_SC_LP__O221AI_2%A_794_367#
x_PM_SKY130_FD_SC_LP__O221AI_2%A_29_69# N_A_29_69#_M1002_s N_A_29_69#_M1005_s
+ N_A_29_69#_M1003_s N_A_29_69#_M1014_s N_A_29_69#_c_602_n N_A_29_69#_c_603_n
+ N_A_29_69#_c_604_n N_A_29_69#_c_614_n N_A_29_69#_c_605_n N_A_29_69#_c_606_n
+ N_A_29_69#_c_618_n N_A_29_69#_c_607_n N_A_29_69#_c_622_n
+ PM_SKY130_FD_SC_LP__O221AI_2%A_29_69#
x_PM_SKY130_FD_SC_LP__O221AI_2%A_305_65# N_A_305_65#_M1003_d N_A_305_65#_M1006_d
+ N_A_305_65#_M1010_d N_A_305_65#_M1009_d N_A_305_65#_M1012_s
+ N_A_305_65#_c_658_n N_A_305_65#_c_659_n N_A_305_65#_c_660_n
+ N_A_305_65#_c_704_n N_A_305_65#_c_661_n N_A_305_65#_c_675_n
+ N_A_305_65#_c_679_n N_A_305_65#_c_662_n N_A_305_65#_c_680_n
+ N_A_305_65#_c_663_n N_A_305_65#_c_664_n N_A_305_65#_c_665_n
+ N_A_305_65#_c_693_n PM_SKY130_FD_SC_LP__O221AI_2%A_305_65#
x_PM_SKY130_FD_SC_LP__O221AI_2%VGND N_VGND_M1011_d N_VGND_M1017_s N_VGND_c_728_n
+ N_VGND_c_729_n VGND N_VGND_c_730_n N_VGND_c_731_n N_VGND_c_732_n
+ N_VGND_c_733_n N_VGND_c_734_n N_VGND_c_735_n PM_SKY130_FD_SC_LP__O221AI_2%VGND
cc_1 VNB N_C1_c_90_n 0.0191041f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.295
cc_2 VNB N_C1_M1004_g 0.00146396f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_3 VNB N_C1_c_92_n 0.0194651f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.295
cc_4 VNB N_C1_M1015_g 0.00148155f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_5 VNB C1 0.019736f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_C1_c_95_n 0.074719f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.46
cc_7 VNB N_B1_M1003_g 0.0263901f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_8 VNB N_B1_M1010_g 0.0222466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_132_n 0.00481956f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_10 VNB N_B1_c_133_n 0.00176867f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.46
cc_11 VNB N_B1_c_134_n 0.0298017f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.46
cc_12 VNB N_B1_c_135_n 0.0441794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B2_c_226_n 0.0165074f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.295
cc_14 VNB N_B2_M1007_g 0.00227023f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_15 VNB N_B2_c_228_n 0.0175636f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.295
cc_16 VNB N_B2_M1019_g 0.00242959f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_17 VNB B2 0.00262528f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_B2_c_231_n 0.0371913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1011_g 0.0210814f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.765
cc_20 VNB N_A1_c_283_n 0.0209775f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.765
cc_21 VNB N_A1_M1016_g 0.00275546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_c_285_n 0.00472528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_286_n 0.024507f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_24 VNB A1 0.0233806f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.46
cc_25 VNB N_A1_c_288_n 0.0536738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_c_367_n 0.0162509f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.295
cc_27 VNB N_A2_M1008_g 0.00263923f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_28 VNB N_A2_c_369_n 0.0162509f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.295
cc_29 VNB N_A2_M1018_g 0.00257203f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_30 VNB A2 0.0104154f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB N_A2_c_372_n 0.0435939f $X=-0.19 $Y=-0.245 $X2=0.222 $Y2=1.46
cc_32 VNB N_VPWR_c_422_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_29_69#_c_602_n 0.023359f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_A_29_69#_c_603_n 0.00506087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_29_69#_c_604_n 0.00935084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_29_69#_c_605_n 0.0152544f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.46
cc_37 VNB N_A_29_69#_c_606_n 0.0039075f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.46
cc_38 VNB N_A_29_69#_c_607_n 0.00289575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_305_65#_c_658_n 0.00500387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_305_65#_c_659_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_41 VNB N_A_305_65#_c_660_n 0.00407928f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_42 VNB N_A_305_65#_c_661_n 0.00595553f $X=-0.19 $Y=-0.245 $X2=0.222 $Y2=1.295
cc_43 VNB N_A_305_65#_c_662_n 0.00218621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_305_65#_c_663_n 0.00742831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_305_65#_c_664_n 0.0239025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_305_65#_c_665_n 0.00150323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_728_n 0.00232955f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.765
cc_48 VNB N_VGND_c_729_n 0.00232955f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_49 VNB N_VGND_c_730_n 0.0931964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_731_n 0.0152212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_732_n 0.0195242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_733_n 0.328125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_734_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_735_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VPB N_C1_M1004_g 0.024561f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_56 VPB N_C1_M1015_g 0.0226316f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_57 VPB C1 0.00691937f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_58 VPB N_B1_M1001_g 0.0224024f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.765
cc_59 VPB N_B1_M1013_g 0.0196206f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_60 VPB N_B1_c_138_n 0.00744879f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_61 VPB N_B1_c_132_n 0.00407099f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_62 VPB N_B1_c_133_n 5.34044e-19 $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.46
cc_63 VPB N_B1_c_134_n 0.00795669f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.46
cc_64 VPB N_B1_c_135_n 0.0168406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_B2_M1007_g 0.019297f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_66 VPB N_B2_M1019_g 0.0187406f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_67 VPB N_A1_M1000_g 0.0204706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A1_M1016_g 0.0227736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A1_c_285_n 5.96505e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A1_c_286_n 0.00644416f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_71 VPB N_A1_c_293_n 0.00866827f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_72 VPB N_A1_c_294_n 0.00102826f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB A1 0.00183157f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.46
cc_74 VPB N_A1_c_296_n 0.0090853f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A2_M1008_g 0.019598f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_76 VPB N_A2_M1018_g 0.0187224f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_77 VPB N_VPWR_c_423_n 0.0105221f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_78 VPB N_VPWR_c_424_n 0.0488337f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_79 VPB N_VPWR_c_425_n 0.00283718f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_80 VPB N_VPWR_c_426_n 0.00564356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_427_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_428_n 0.043525f $X=-0.19 $Y=1.655 $X2=0.222 $Y2=1.46
cc_83 VPB N_VPWR_c_429_n 0.0154314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_430_n 0.0376032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_431_n 0.0386847f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_432_n 0.0138973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_433_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_422_n 0.0450415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_Y_c_500_n 0.00440089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 N_C1_M1015_g N_B1_c_132_n 0.00266411f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_91 N_C1_c_95_n N_B1_c_132_n 0.00118591f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_92 N_C1_c_95_n N_B1_c_135_n 0.011878f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_93 N_C1_M1004_g N_VPWR_c_424_n 0.00483162f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_94 C1 N_VPWR_c_424_n 0.0224262f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_95 N_C1_c_95_n N_VPWR_c_424_n 0.00144108f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_96 N_C1_M1004_g N_VPWR_c_425_n 7.28915e-19 $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_97 N_C1_M1015_g N_VPWR_c_425_n 0.0147054f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_98 N_C1_M1004_g N_VPWR_c_429_n 0.0054895f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_99 N_C1_M1015_g N_VPWR_c_429_n 0.00486043f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_100 N_C1_M1004_g N_VPWR_c_422_n 0.0107076f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_101 N_C1_M1015_g N_VPWR_c_422_n 0.00824727f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_102 N_C1_M1004_g N_Y_c_501_n 0.010366f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_103 N_C1_M1004_g N_Y_c_500_n 0.00879487f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_104 N_C1_M1015_g N_Y_c_500_n 0.0277462f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_105 N_C1_c_90_n N_Y_c_504_n 0.0146534f $X=0.485 $Y=1.295 $X2=0 $Y2=0
cc_106 N_C1_M1004_g N_Y_c_504_n 0.00638994f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_107 N_C1_c_92_n N_Y_c_504_n 0.0105158f $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_108 N_C1_M1015_g N_Y_c_504_n 0.00611876f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_109 C1 N_Y_c_504_n 0.0388367f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_110 N_C1_c_95_n N_Y_c_504_n 0.0262323f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_111 C1 N_A_29_69#_c_602_n 0.022426f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_112 N_C1_c_95_n N_A_29_69#_c_602_n 0.0015759f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_113 N_C1_c_90_n N_A_29_69#_c_603_n 0.0128219f $X=0.485 $Y=1.295 $X2=0 $Y2=0
cc_114 N_C1_c_92_n N_A_29_69#_c_603_n 0.0127816f $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_115 N_C1_c_92_n N_A_29_69#_c_606_n 0.00162302f $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_116 N_C1_c_92_n N_A_305_65#_c_660_n 6.09955e-19 $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_117 N_C1_c_90_n N_VGND_c_730_n 0.0029147f $X=0.485 $Y=1.295 $X2=0 $Y2=0
cc_118 N_C1_c_92_n N_VGND_c_730_n 0.0029147f $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_119 N_C1_c_90_n N_VGND_c_733_n 0.00420369f $X=0.485 $Y=1.295 $X2=0 $Y2=0
cc_120 N_C1_c_92_n N_VGND_c_733_n 0.00428625f $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_121 N_B1_M1003_g N_B2_c_226_n 0.0258829f $X=1.865 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_122 N_B1_M1001_g N_B2_M1007_g 0.0296432f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B1_c_138_n N_B2_M1007_g 0.00923201f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_124 N_B1_c_132_n N_B2_M1007_g 0.00628799f $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_125 N_B1_M1010_g N_B2_c_228_n 0.0198867f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_126 N_B1_M1013_g N_B2_M1019_g 0.0381109f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B1_c_138_n N_B2_M1019_g 0.0109831f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_128 N_B1_c_132_n N_B2_M1019_g 4.78402e-19 $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_129 N_B1_c_133_n N_B2_M1019_g 6.09034e-19 $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_130 N_B1_M1003_g B2 2.9131e-19 $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_131 N_B1_M1010_g B2 6.98768e-19 $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_132 N_B1_c_138_n B2 0.025828f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_133 N_B1_c_132_n B2 0.00881824f $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_134 N_B1_c_133_n B2 0.00897351f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_135 N_B1_c_134_n B2 6.74005e-19 $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_136 N_B1_c_135_n B2 4.71921e-19 $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_137 N_B1_c_138_n N_B2_c_231_n 0.00243405f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_138 N_B1_c_132_n N_B2_c_231_n 0.00788422f $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_139 N_B1_c_133_n N_B2_c_231_n 0.00154435f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_140 N_B1_c_134_n N_B2_c_231_n 0.0220693f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_141 N_B1_c_135_n N_B2_c_231_n 0.0166692f $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_142 N_B1_M1010_g N_A1_M1011_g 0.019821f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_143 N_B1_M1013_g N_A1_M1000_g 0.0293007f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_144 N_B1_c_138_n N_A1_M1000_g 6.00451e-19 $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_145 N_B1_c_133_n N_A1_c_285_n 0.022339f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_146 N_B1_c_134_n N_A1_c_285_n 0.00118578f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_147 N_B1_c_133_n N_A1_c_286_n 0.00114936f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_148 N_B1_c_134_n N_A1_c_286_n 0.0203676f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_149 N_B1_M1013_g N_A1_c_294_n 6.00967e-19 $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_150 N_B1_c_138_n N_A1_c_294_n 0.0135638f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_151 N_B1_c_133_n N_A1_c_294_n 7.26095e-19 $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_152 N_B1_c_132_n N_VPWR_M1015_d 0.00304131f $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_153 N_B1_c_138_n N_VPWR_M1013_d 0.00163876f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_154 N_B1_M1001_g N_VPWR_c_425_n 0.0158272f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_155 N_B1_M1013_g N_VPWR_c_426_n 0.0105261f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_156 N_B1_M1001_g N_VPWR_c_430_n 0.00486043f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_157 N_B1_M1013_g N_VPWR_c_430_n 0.00547432f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B1_M1001_g N_VPWR_c_422_n 0.00843225f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B1_M1013_g N_VPWR_c_422_n 0.010534f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_160 N_B1_c_138_n N_Y_M1007_s 0.00176461f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_161 N_B1_M1001_g N_Y_c_511_n 0.0167067f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_162 N_B1_c_138_n N_Y_c_511_n 0.00671026f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_163 N_B1_c_132_n N_Y_c_511_n 0.0555727f $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_164 N_B1_c_135_n N_Y_c_511_n 0.00235675f $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_165 N_B1_M1001_g N_Y_c_500_n 0.00543679f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_166 N_B1_c_132_n N_Y_c_500_n 0.00444706f $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_167 N_B1_M1013_g N_Y_c_517_n 0.0152971f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_168 N_B1_c_138_n N_Y_c_517_n 0.040698f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_169 N_B1_c_134_n N_Y_c_517_n 6.86769e-19 $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_170 N_B1_M1001_g N_Y_c_520_n 8.13212e-19 $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_171 N_B1_M1013_g N_Y_c_520_n 7.61432e-19 $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_172 N_B1_c_138_n N_Y_c_520_n 0.0172505f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_173 N_B1_c_132_n N_Y_c_504_n 0.0127724f $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_174 N_B1_c_135_n N_Y_c_504_n 7.12728e-19 $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_175 N_B1_c_132_n N_A_388_367#_M1001_s 0.00258529f $X=2.315 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_176 N_B1_c_138_n N_A_388_367#_M1019_d 0.00176891f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_177 N_B1_M1013_g N_A_388_367#_c_567_n 0.00218451f $X=3.225 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_B1_M1013_g N_A_388_367#_c_568_n 0.00637863f $X=3.225 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_B1_M1003_g N_A_29_69#_c_603_n 5.15082e-19 $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_180 N_B1_M1003_g N_A_29_69#_c_614_n 0.00269095f $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_181 N_B1_M1003_g N_A_29_69#_c_605_n 0.0133735f $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_182 N_B1_c_132_n N_A_29_69#_c_605_n 0.0479888f $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_183 N_B1_c_135_n N_A_29_69#_c_605_n 0.0119251f $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_184 N_B1_c_138_n N_A_29_69#_c_618_n 0.00403051f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_185 N_B1_M1003_g N_A_29_69#_c_607_n 4.46099e-19 $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_186 N_B1_c_132_n N_A_29_69#_c_607_n 0.0293817f $X=2.315 $Y=1.79 $X2=0 $Y2=0
cc_187 N_B1_c_135_n N_A_29_69#_c_607_n 8.69935e-19 $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_188 N_B1_M1010_g N_A_29_69#_c_622_n 0.0113094f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_189 N_B1_c_138_n N_A_29_69#_c_622_n 0.00785499f $X=3.14 $Y=1.79 $X2=0 $Y2=0
cc_190 N_B1_c_133_n N_A_29_69#_c_622_n 0.0128684f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_191 N_B1_c_134_n N_A_29_69#_c_622_n 0.00284053f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_192 N_B1_M1003_g N_A_305_65#_c_658_n 0.00697855f $X=1.865 $Y=0.745 $X2=0
+ $Y2=0
cc_193 N_B1_M1003_g N_A_305_65#_c_659_n 0.00863921f $X=1.865 $Y=0.745 $X2=0
+ $Y2=0
cc_194 N_B1_M1003_g N_A_305_65#_c_660_n 0.00193542f $X=1.865 $Y=0.745 $X2=0
+ $Y2=0
cc_195 N_B1_M1010_g N_A_305_65#_c_661_n 0.0125548f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_196 N_B1_M1010_g N_VGND_c_728_n 4.97374e-19 $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_197 N_B1_M1003_g N_VGND_c_730_n 0.00302473f $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_198 N_B1_M1010_g N_VGND_c_730_n 0.00302501f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_199 N_B1_M1003_g N_VGND_c_733_n 0.00491773f $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_200 N_B1_M1010_g N_VGND_c_733_n 0.00450282f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_201 N_B2_M1007_g N_VPWR_c_425_n 0.00104976f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B2_M1007_g N_VPWR_c_430_n 0.00357877f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B2_M1019_g N_VPWR_c_430_n 0.00357877f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B2_M1007_g N_VPWR_c_422_n 0.00553619f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B2_M1019_g N_VPWR_c_422_n 0.00537654f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_206 N_B2_M1007_g N_Y_c_511_n 0.0114816f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B2_M1019_g N_Y_c_517_n 0.0111034f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B2_M1007_g N_Y_c_520_n 0.00944955f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_209 N_B2_M1019_g N_Y_c_520_n 0.00923548f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_210 N_B2_M1007_g N_A_388_367#_c_567_n 0.0115031f $X=2.365 $Y=2.465 $X2=0
+ $Y2=0
cc_211 N_B2_M1019_g N_A_388_367#_c_567_n 0.0115031f $X=2.795 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_B2_c_226_n N_A_29_69#_c_618_n 0.0109883f $X=2.365 $Y=1.275 $X2=0 $Y2=0
cc_213 N_B2_c_228_n N_A_29_69#_c_618_n 0.0100482f $X=2.795 $Y=1.275 $X2=0 $Y2=0
cc_214 B2 N_A_29_69#_c_618_n 0.0239985f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_215 N_B2_c_231_n N_A_29_69#_c_618_n 5.91533e-19 $X=2.795 $Y=1.44 $X2=0 $Y2=0
cc_216 N_B2_c_226_n N_A_29_69#_c_607_n 0.0102547f $X=2.365 $Y=1.275 $X2=0 $Y2=0
cc_217 N_B2_c_228_n N_A_29_69#_c_607_n 0.00141777f $X=2.795 $Y=1.275 $X2=0 $Y2=0
cc_218 B2 N_A_29_69#_c_607_n 0.00357748f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_219 N_B2_c_226_n N_A_29_69#_c_622_n 4.49684e-19 $X=2.365 $Y=1.275 $X2=0 $Y2=0
cc_220 N_B2_c_228_n N_A_29_69#_c_622_n 0.00946355f $X=2.795 $Y=1.275 $X2=0 $Y2=0
cc_221 N_B2_c_226_n N_A_305_65#_c_658_n 2.75259e-19 $X=2.365 $Y=1.275 $X2=0
+ $Y2=0
cc_222 N_B2_c_226_n N_A_305_65#_c_659_n 0.0098642f $X=2.365 $Y=1.275 $X2=0 $Y2=0
cc_223 N_B2_c_228_n N_A_305_65#_c_661_n 0.0105038f $X=2.795 $Y=1.275 $X2=0 $Y2=0
cc_224 N_B2_c_226_n N_VGND_c_730_n 0.00302501f $X=2.365 $Y=1.275 $X2=0 $Y2=0
cc_225 N_B2_c_228_n N_VGND_c_730_n 0.00302501f $X=2.795 $Y=1.275 $X2=0 $Y2=0
cc_226 N_B2_c_226_n N_VGND_c_733_n 0.00441786f $X=2.365 $Y=1.275 $X2=0 $Y2=0
cc_227 N_B2_c_228_n N_VGND_c_733_n 0.00449308f $X=2.795 $Y=1.275 $X2=0 $Y2=0
cc_228 N_A1_M1011_g N_A2_c_367_n 0.0293926f $X=3.825 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_229 N_A1_M1000_g N_A2_M1008_g 0.0378042f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A1_c_285_n N_A2_M1008_g 0.0018065f $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_231 N_A1_c_286_n N_A2_M1008_g 0.00244667f $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_232 N_A1_c_293_n N_A2_M1008_g 0.0112859f $X=5.345 $Y=1.785 $X2=0 $Y2=0
cc_233 N_A1_c_283_n N_A2_c_369_n 0.0270857f $X=5.195 $Y=1.275 $X2=0 $Y2=0
cc_234 N_A1_M1016_g N_A2_M1018_g 0.0258539f $X=5.265 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A1_c_293_n N_A2_M1018_g 0.0146827f $X=5.345 $Y=1.785 $X2=0 $Y2=0
cc_236 N_A1_M1011_g A2 8.01844e-19 $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_237 N_A1_c_283_n A2 0.00234406f $X=5.195 $Y=1.275 $X2=0 $Y2=0
cc_238 N_A1_c_285_n A2 0.0130552f $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_239 N_A1_c_286_n A2 2.223e-19 $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_240 N_A1_c_293_n A2 0.0715647f $X=5.345 $Y=1.785 $X2=0 $Y2=0
cc_241 A1 A2 0.0251761f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_242 N_A1_c_288_n A2 0.00757403f $X=5.49 $Y=1.44 $X2=0 $Y2=0
cc_243 N_A1_c_285_n N_A2_c_372_n 0.00247602f $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_244 N_A1_c_286_n N_A2_c_372_n 0.0170413f $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_245 N_A1_c_293_n N_A2_c_372_n 0.00608571f $X=5.345 $Y=1.785 $X2=0 $Y2=0
cc_246 A1 N_A2_c_372_n 5.29727e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_247 N_A1_c_288_n N_A2_c_372_n 0.0224852f $X=5.49 $Y=1.44 $X2=0 $Y2=0
cc_248 N_A1_c_294_n N_VPWR_M1013_d 0.00131337f $X=4.015 $Y=1.785 $X2=0 $Y2=0
cc_249 N_A1_c_296_n N_VPWR_M1016_d 0.0024884f $X=5.507 $Y=1.695 $X2=0 $Y2=0
cc_250 N_A1_M1000_g N_VPWR_c_426_n 0.0113483f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A1_M1016_g N_VPWR_c_428_n 0.017873f $X=5.265 $Y=2.465 $X2=0 $Y2=0
cc_252 N_A1_c_293_n N_VPWR_c_428_n 0.0017933f $X=5.345 $Y=1.785 $X2=0 $Y2=0
cc_253 N_A1_c_288_n N_VPWR_c_428_n 0.00120978f $X=5.49 $Y=1.44 $X2=0 $Y2=0
cc_254 N_A1_c_296_n N_VPWR_c_428_n 0.0223707f $X=5.507 $Y=1.695 $X2=0 $Y2=0
cc_255 N_A1_M1000_g N_VPWR_c_431_n 0.00585385f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_256 N_A1_M1016_g N_VPWR_c_431_n 0.00486043f $X=5.265 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A1_M1000_g N_VPWR_c_422_n 0.0117279f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A1_M1016_g N_VPWR_c_422_n 0.0082726f $X=5.265 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A1_c_293_n N_Y_M1008_s 0.00176773f $X=5.345 $Y=1.785 $X2=0 $Y2=0
cc_260 N_A1_M1000_g N_Y_c_517_n 0.016459f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A1_c_286_n N_Y_c_517_n 5.23226e-19 $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_262 N_A1_c_293_n N_Y_c_517_n 0.0264208f $X=5.345 $Y=1.785 $X2=0 $Y2=0
cc_263 N_A1_c_294_n N_Y_c_517_n 0.0178103f $X=4.015 $Y=1.785 $X2=0 $Y2=0
cc_264 N_A1_M1000_g N_Y_c_534_n 8.75385e-19 $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A1_c_293_n N_Y_c_534_n 0.0172972f $X=5.345 $Y=1.785 $X2=0 $Y2=0
cc_266 N_A1_c_293_n N_A_794_367#_M1000_s 0.00262603f $X=5.345 $Y=1.785 $X2=-0.19
+ $Y2=-0.245
cc_267 N_A1_c_293_n N_A_794_367#_M1018_d 0.00176773f $X=5.345 $Y=1.785 $X2=0
+ $Y2=0
cc_268 N_A1_c_293_n N_A_794_367#_c_587_n 0.0135577f $X=5.345 $Y=1.785 $X2=0
+ $Y2=0
cc_269 N_A1_M1011_g N_A_29_69#_c_622_n 4.48052e-19 $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_270 N_A1_M1011_g N_A_305_65#_c_661_n 6.00676e-19 $X=3.825 $Y=0.745 $X2=0
+ $Y2=0
cc_271 N_A1_M1011_g N_A_305_65#_c_675_n 0.013485f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_272 N_A1_c_285_n N_A_305_65#_c_675_n 0.0121224f $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_273 N_A1_c_286_n N_A_305_65#_c_675_n 5.1677e-19 $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_274 N_A1_c_293_n N_A_305_65#_c_675_n 0.00497222f $X=5.345 $Y=1.785 $X2=0
+ $Y2=0
cc_275 N_A1_c_285_n N_A_305_65#_c_679_n 0.00121501f $X=3.845 $Y=1.51 $X2=0 $Y2=0
cc_276 N_A1_c_283_n N_A_305_65#_c_680_n 0.0141116f $X=5.195 $Y=1.275 $X2=0 $Y2=0
cc_277 N_A1_c_293_n N_A_305_65#_c_680_n 0.00241788f $X=5.345 $Y=1.785 $X2=0
+ $Y2=0
cc_278 N_A1_c_293_n N_A_305_65#_c_663_n 8.48612e-19 $X=5.345 $Y=1.785 $X2=0
+ $Y2=0
cc_279 A1 N_A_305_65#_c_663_n 0.021086f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_280 N_A1_c_288_n N_A_305_65#_c_663_n 0.00283538f $X=5.49 $Y=1.44 $X2=0 $Y2=0
cc_281 N_A1_c_283_n N_A_305_65#_c_664_n 0.00234009f $X=5.195 $Y=1.275 $X2=0
+ $Y2=0
cc_282 N_A1_M1011_g N_VGND_c_728_n 0.00755047f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_283 N_A1_c_283_n N_VGND_c_729_n 0.00958261f $X=5.195 $Y=1.275 $X2=0 $Y2=0
cc_284 N_A1_M1011_g N_VGND_c_730_n 0.00481374f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_285 N_A1_c_283_n N_VGND_c_732_n 0.00481374f $X=5.195 $Y=1.275 $X2=0 $Y2=0
cc_286 N_A1_M1011_g N_VGND_c_733_n 0.00912395f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_287 N_A1_c_283_n N_VGND_c_733_n 0.00950163f $X=5.195 $Y=1.275 $X2=0 $Y2=0
cc_288 N_A2_M1018_g N_VPWR_c_428_n 0.00109252f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_289 N_A2_M1008_g N_VPWR_c_431_n 0.00357877f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_290 N_A2_M1018_g N_VPWR_c_431_n 0.00357877f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A2_M1008_g N_VPWR_c_422_n 0.00555738f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A2_M1018_g N_VPWR_c_422_n 0.00537654f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A2_M1008_g N_Y_c_517_n 0.0115313f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A2_M1008_g N_Y_c_534_n 0.00925722f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_295 N_A2_M1018_g N_Y_c_534_n 0.00897551f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_296 N_A2_M1008_g N_A_794_367#_c_588_n 0.011751f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A2_M1018_g N_A_794_367#_c_588_n 0.0118004f $X=4.835 $Y=2.465 $X2=0
+ $Y2=0
cc_298 N_A2_c_367_n N_A_305_65#_c_675_n 0.0127501f $X=4.295 $Y=1.275 $X2=0 $Y2=0
cc_299 A2 N_A_305_65#_c_675_n 0.0116716f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_300 N_A2_c_367_n N_A_305_65#_c_662_n 5.75621e-19 $X=4.295 $Y=1.275 $X2=0
+ $Y2=0
cc_301 N_A2_c_369_n N_A_305_65#_c_662_n 5.75621e-19 $X=4.725 $Y=1.275 $X2=0
+ $Y2=0
cc_302 N_A2_c_369_n N_A_305_65#_c_680_n 0.0127501f $X=4.725 $Y=1.275 $X2=0 $Y2=0
cc_303 A2 N_A_305_65#_c_680_n 0.0362956f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_304 N_A2_c_372_n N_A_305_65#_c_680_n 5.33262e-19 $X=4.835 $Y=1.44 $X2=0 $Y2=0
cc_305 A2 N_A_305_65#_c_693_n 0.0169989f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_306 N_A2_c_372_n N_A_305_65#_c_693_n 6.61019e-19 $X=4.835 $Y=1.44 $X2=0 $Y2=0
cc_307 N_A2_c_367_n N_VGND_c_728_n 0.00748198f $X=4.295 $Y=1.275 $X2=0 $Y2=0
cc_308 N_A2_c_369_n N_VGND_c_728_n 4.3911e-19 $X=4.725 $Y=1.275 $X2=0 $Y2=0
cc_309 N_A2_c_367_n N_VGND_c_729_n 4.3911e-19 $X=4.295 $Y=1.275 $X2=0 $Y2=0
cc_310 N_A2_c_369_n N_VGND_c_729_n 0.00748198f $X=4.725 $Y=1.275 $X2=0 $Y2=0
cc_311 N_A2_c_367_n N_VGND_c_731_n 0.00481374f $X=4.295 $Y=1.275 $X2=0 $Y2=0
cc_312 N_A2_c_369_n N_VGND_c_731_n 0.00481374f $X=4.725 $Y=1.275 $X2=0 $Y2=0
cc_313 N_A2_c_367_n N_VGND_c_733_n 0.00911421f $X=4.295 $Y=1.275 $X2=0 $Y2=0
cc_314 N_A2_c_369_n N_VGND_c_733_n 0.00911421f $X=4.725 $Y=1.275 $X2=0 $Y2=0
cc_315 N_VPWR_c_422_n N_Y_M1004_s 0.00380103f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_316 N_VPWR_c_422_n N_Y_M1007_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_317 N_VPWR_c_422_n N_Y_M1008_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_318 N_VPWR_c_429_n N_Y_c_501_n 0.015688f $X=0.965 $Y=3.33 $X2=0 $Y2=0
cc_319 N_VPWR_c_422_n N_Y_c_501_n 0.00984745f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_M1015_d N_Y_c_511_n 0.0113083f $X=0.99 $Y=1.835 $X2=0 $Y2=0
cc_321 N_VPWR_c_425_n N_Y_c_511_n 0.0341303f $X=1.65 $Y=2.49 $X2=0 $Y2=0
cc_322 N_VPWR_M1015_d N_Y_c_500_n 0.012957f $X=0.99 $Y=1.835 $X2=0 $Y2=0
cc_323 N_VPWR_c_425_n N_Y_c_500_n 0.0268202f $X=1.65 $Y=2.49 $X2=0 $Y2=0
cc_324 N_VPWR_M1013_d N_Y_c_517_n 0.017714f $X=3.3 $Y=1.835 $X2=0 $Y2=0
cc_325 N_VPWR_c_426_n N_Y_c_517_n 0.0266856f $X=3.56 $Y=2.51 $X2=0 $Y2=0
cc_326 N_VPWR_c_422_n N_A_388_367#_M1001_s 0.00432919f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_327 N_VPWR_c_422_n N_A_388_367#_M1019_d 0.00223562f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_426_n N_A_388_367#_c_567_n 0.0114735f $X=3.56 $Y=2.51 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_430_n N_A_388_367#_c_567_n 0.0519231f $X=3.395 $Y=3.33 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_422_n N_A_388_367#_c_567_n 0.0336005f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_430_n N_A_388_367#_c_576_n 0.0174631f $X=3.395 $Y=3.33 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_422_n N_A_388_367#_c_576_n 0.0101068f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_426_n N_A_388_367#_c_568_n 0.0325112f $X=3.56 $Y=2.51 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_422_n N_A_794_367#_M1000_s 0.00480031f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_335 N_VPWR_c_422_n N_A_794_367#_M1018_d 0.00376627f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_336 N_VPWR_c_431_n N_A_794_367#_c_588_n 0.0362264f $X=5.315 $Y=3.33 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_422_n N_A_794_367#_c_588_n 0.0237058f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_431_n N_A_794_367#_c_594_n 0.0178122f $X=5.315 $Y=3.33 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_422_n N_A_794_367#_c_594_n 0.0101015f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_431_n N_A_794_367#_c_596_n 0.0125234f $X=5.315 $Y=3.33 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_422_n N_A_794_367#_c_596_n 0.00738676f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_342 N_Y_c_511_n N_A_388_367#_M1001_s 0.00498051f $X=2.415 $Y=2.13 $X2=-0.19
+ $Y2=1.655
cc_343 N_Y_c_517_n N_A_388_367#_M1019_d 0.00351257f $X=4.455 $Y=2.13 $X2=0 $Y2=0
cc_344 N_Y_c_511_n N_A_388_367#_c_581_n 0.0192236f $X=2.415 $Y=2.13 $X2=0 $Y2=0
cc_345 N_Y_M1007_s N_A_388_367#_c_567_n 0.00332344f $X=2.44 $Y=1.835 $X2=0 $Y2=0
cc_346 N_Y_c_520_n N_A_388_367#_c_567_n 0.0159985f $X=2.58 $Y=2.13 $X2=0 $Y2=0
cc_347 N_Y_c_517_n N_A_388_367#_c_568_n 0.0153099f $X=4.455 $Y=2.13 $X2=0 $Y2=0
cc_348 N_Y_c_517_n N_A_794_367#_M1000_s 0.00516361f $X=4.455 $Y=2.13 $X2=-0.19
+ $Y2=1.655
cc_349 N_Y_c_517_n N_A_794_367#_c_599_n 0.0200381f $X=4.455 $Y=2.13 $X2=0 $Y2=0
cc_350 N_Y_M1008_s N_A_794_367#_c_588_n 0.00332931f $X=4.48 $Y=1.835 $X2=0 $Y2=0
cc_351 N_Y_c_534_n N_A_794_367#_c_588_n 0.0160814f $X=4.62 $Y=2.13 $X2=0 $Y2=0
cc_352 N_Y_M1002_d N_A_29_69#_c_603_n 0.00176461f $X=0.56 $Y=0.345 $X2=0 $Y2=0
cc_353 N_Y_c_504_n N_A_29_69#_c_603_n 0.0159805f $X=0.7 $Y=0.68 $X2=0 $Y2=0
cc_354 N_Y_c_500_n N_A_29_69#_c_605_n 0.00318646f $X=1.335 $Y=2.13 $X2=0 $Y2=0
cc_355 N_Y_c_500_n N_A_29_69#_c_606_n 0.00725788f $X=1.335 $Y=2.13 $X2=0 $Y2=0
cc_356 N_Y_c_504_n N_A_29_69#_c_606_n 0.009209f $X=0.7 $Y=0.68 $X2=0 $Y2=0
cc_357 N_A_29_69#_c_605_n N_A_305_65#_M1003_d 0.00258276f $X=1.985 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_358 N_A_29_69#_c_618_n N_A_305_65#_M1006_d 0.00332139f $X=2.865 $Y=0.955
+ $X2=0 $Y2=0
cc_359 N_A_29_69#_c_614_n N_A_305_65#_c_658_n 0.0291516f $X=1.13 $Y=0.49 $X2=0
+ $Y2=0
cc_360 N_A_29_69#_c_605_n N_A_305_65#_c_658_n 0.0219488f $X=1.985 $Y=1.17 $X2=0
+ $Y2=0
cc_361 N_A_29_69#_M1003_s N_A_305_65#_c_659_n 0.00250873f $X=1.94 $Y=0.325 $X2=0
+ $Y2=0
cc_362 N_A_29_69#_c_605_n N_A_305_65#_c_659_n 0.00272017f $X=1.985 $Y=1.17 $X2=0
+ $Y2=0
cc_363 N_A_29_69#_c_618_n N_A_305_65#_c_659_n 0.00387154f $X=2.865 $Y=0.955
+ $X2=0 $Y2=0
cc_364 N_A_29_69#_c_607_n N_A_305_65#_c_659_n 0.0195903f $X=2.15 $Y=0.68 $X2=0
+ $Y2=0
cc_365 N_A_29_69#_c_603_n N_A_305_65#_c_660_n 0.0119903f $X=1.045 $Y=0.34 $X2=0
+ $Y2=0
cc_366 N_A_29_69#_c_618_n N_A_305_65#_c_704_n 0.0130514f $X=2.865 $Y=0.955 $X2=0
+ $Y2=0
cc_367 N_A_29_69#_M1014_s N_A_305_65#_c_661_n 0.00406492f $X=2.87 $Y=0.325 $X2=0
+ $Y2=0
cc_368 N_A_29_69#_c_618_n N_A_305_65#_c_661_n 0.00447792f $X=2.865 $Y=0.955
+ $X2=0 $Y2=0
cc_369 N_A_29_69#_c_622_n N_A_305_65#_c_661_n 0.0271302f $X=3.03 $Y=0.68 $X2=0
+ $Y2=0
cc_370 N_A_29_69#_c_603_n N_VGND_c_730_n 0.0564933f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_371 N_A_29_69#_c_604_n N_VGND_c_730_n 0.0186386f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_372 N_A_29_69#_c_603_n N_VGND_c_733_n 0.03158f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_373 N_A_29_69#_c_604_n N_VGND_c_733_n 0.0101082f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_374 N_A_305_65#_c_675_n N_VGND_M1011_d 0.0058703f $X=4.395 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_375 N_A_305_65#_c_680_n N_VGND_M1017_s 0.00427446f $X=5.295 $Y=0.955 $X2=0
+ $Y2=0
cc_376 N_A_305_65#_c_661_n N_VGND_c_728_n 0.00920891f $X=3.515 $Y=0.34 $X2=0
+ $Y2=0
cc_377 N_A_305_65#_c_675_n N_VGND_c_728_n 0.017285f $X=4.395 $Y=0.955 $X2=0
+ $Y2=0
cc_378 N_A_305_65#_c_662_n N_VGND_c_728_n 0.0155698f $X=4.51 $Y=0.47 $X2=0 $Y2=0
cc_379 N_A_305_65#_c_662_n N_VGND_c_729_n 0.0155698f $X=4.51 $Y=0.47 $X2=0 $Y2=0
cc_380 N_A_305_65#_c_680_n N_VGND_c_729_n 0.017285f $X=5.295 $Y=0.955 $X2=0
+ $Y2=0
cc_381 N_A_305_65#_c_664_n N_VGND_c_729_n 0.0155924f $X=5.41 $Y=0.47 $X2=0 $Y2=0
cc_382 N_A_305_65#_c_659_n N_VGND_c_730_n 0.0423044f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_383 N_A_305_65#_c_660_n N_VGND_c_730_n 0.0235159f $X=1.815 $Y=0.34 $X2=0
+ $Y2=0
cc_384 N_A_305_65#_c_661_n N_VGND_c_730_n 0.0662288f $X=3.515 $Y=0.34 $X2=0
+ $Y2=0
cc_385 N_A_305_65#_c_665_n N_VGND_c_730_n 0.0145891f $X=2.59 $Y=0.34 $X2=0 $Y2=0
cc_386 N_A_305_65#_c_662_n N_VGND_c_731_n 0.0124036f $X=4.51 $Y=0.47 $X2=0 $Y2=0
cc_387 N_A_305_65#_c_664_n N_VGND_c_732_n 0.0151237f $X=5.41 $Y=0.47 $X2=0 $Y2=0
cc_388 N_A_305_65#_c_659_n N_VGND_c_733_n 0.0239316f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_389 N_A_305_65#_c_660_n N_VGND_c_733_n 0.0127052f $X=1.815 $Y=0.34 $X2=0
+ $Y2=0
cc_390 N_A_305_65#_c_661_n N_VGND_c_733_n 0.0372325f $X=3.515 $Y=0.34 $X2=0
+ $Y2=0
cc_391 N_A_305_65#_c_662_n N_VGND_c_733_n 0.00864148f $X=4.51 $Y=0.47 $X2=0
+ $Y2=0
cc_392 N_A_305_65#_c_664_n N_VGND_c_733_n 0.0105365f $X=5.41 $Y=0.47 $X2=0 $Y2=0
cc_393 N_A_305_65#_c_665_n N_VGND_c_733_n 0.00807735f $X=2.59 $Y=0.34 $X2=0
+ $Y2=0
