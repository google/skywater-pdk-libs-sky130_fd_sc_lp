* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfxtp_lp CLK D SCD SCE VGND VNB VPB VPWR Q
X0 VGND a_733_66# a_978_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND a_1957_347# a_2359_69# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_733_66# CLK a_820_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_457_417# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_1576_99# a_733_66# a_1957_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_531_125# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_1263_155# a_1722_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_351_417# D a_457_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_1263_155# a_733_66# a_351_417# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_733_66# a_998_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VPWR a_1263_155# a_1576_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_1160_155# a_998_347# a_1263_155# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1957_347# a_998_347# a_1576_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_27_409# a_351_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 Q a_2148_185# a_2628_69# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_27_409# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_1263_155# a_733_66# a_1528_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_27_409# SCE a_159_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_351_417# SCE a_531_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_2359_69# a_1957_347# a_2148_185# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1528_347# a_1576_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 Q a_2148_185# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_351_125# D a_351_417# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_1957_347# a_998_347# a_2095_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X24 VPWR SCD a_244_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 a_159_125# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_244_417# a_27_409# a_351_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 a_733_66# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X28 a_820_66# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1910_155# a_2148_185# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_2628_69# a_2148_185# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_1910_155# a_733_66# a_1957_347# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VPWR a_1957_347# a_2148_185# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X33 a_1160_155# a_1576_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_351_417# a_998_347# a_1263_155# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X35 a_1722_125# a_1263_155# a_1576_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_2095_361# a_2148_185# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X37 a_978_66# a_733_66# a_998_347# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
