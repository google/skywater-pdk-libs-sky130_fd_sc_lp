* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a41o_lp A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_314_47# A1 a_428_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR A3 a_27_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VPWR A1 a_27_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_27_409# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_700_47# a_428_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_27_409# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_128_47# A3 a_206_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_428_47# B1 a_542_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND A4 a_128_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_206_47# A2 a_314_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_542_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_428_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 VGND a_428_47# a_700_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_409# B1 a_428_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
