# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__o2111a_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o2111a_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.035000 3.755000 2.200000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715000 1.140000 3.215000 1.825000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 1.140000 2.510000 1.865000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 0.375000 1.855000 1.865000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.080000 1.360000 1.865000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.265000 0.355000 2.385000 ;
        RECT 0.085000 2.385000 0.670000 3.065000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.840000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 4.030000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.525000  0.085000 0.855000 0.570000 ;
      RECT 0.525000  0.740000 1.375000 0.910000 ;
      RECT 0.525000  0.910000 0.795000 2.035000 ;
      RECT 0.525000  2.035000 2.800000 2.215000 ;
      RECT 0.840000  2.385000 1.135000 3.245000 ;
      RECT 1.120000  0.280000 1.375000 0.740000 ;
      RECT 1.305000  2.215000 1.570000 3.075000 ;
      RECT 1.740000  2.385000 2.340000 3.245000 ;
      RECT 2.270000  0.280000 2.565000 0.695000 ;
      RECT 2.270000  0.695000 3.530000 0.865000 ;
      RECT 2.510000  2.215000 2.800000 3.075000 ;
      RECT 2.735000  0.085000 3.065000 0.525000 ;
      RECT 3.250000  0.280000 3.530000 0.695000 ;
      RECT 3.260000  2.385000 3.590000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__o2111a_0
END LIBRARY
