* NGSPICE file created from sky130_fd_sc_lp__buf_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__buf_2 A VGND VNB VPB VPWR X
M1000 X a_90_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=6.405e+11p ps=5.35e+06u
M1001 X a_90_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=9.832e+11p ps=6.95e+06u
M1002 a_90_21# A VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1003 VGND a_90_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_90_21# A VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 VPWR a_90_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

