* File: sky130_fd_sc_lp__or3b_lp.pex.spice
* Created: Fri Aug 28 11:24:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3B_LP%C_N 1 3 7 10 12 14 16 17 18 19 20 24 26
r48 24 26 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.34
+ $X2=0.597 $Y2=1.175
r49 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.34 $X2=0.61 $Y2=1.34
r50 20 25 9.60369 $w=3.88e-07 $l=3.25e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.34
r51 19 25 1.32974 $w=3.88e-07 $l=4.5e-08 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.34
r52 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.855 $Y=0.73
+ $X2=0.855 $Y2=0.445
r53 13 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.57 $Y=0.805
+ $X2=0.495 $Y2=0.805
r54 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.855 $Y2=0.73
r55 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.57 $Y2=0.805
r56 10 18 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.545 $Y=2.545
+ $X2=0.545 $Y2=1.845
r57 7 18 33.8903 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.597 $Y=1.668
+ $X2=0.597 $Y2=1.845
r58 6 24 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.597 $Y=1.352
+ $X2=0.597 $Y2=1.34
r59 6 7 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.597 $Y=1.352
+ $X2=0.597 $Y2=1.668
r60 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=0.805
r61 4 26 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=1.175
r62 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.73
+ $X2=0.495 $Y2=0.805
r63 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.73 $X2=0.495
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_LP%A_27_47# 1 2 9 11 15 19 21 23 24 27 33 35 39
+ 42 44 45 49
r87 48 49 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.285 $Y=1.285
+ $X2=1.36 $Y2=1.285
r88 44 45 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=2.19
+ $X2=0.27 $Y2=2.025
r89 40 48 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=1.18 $Y=1.285
+ $X2=1.285 $Y2=1.285
r90 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.285 $X2=1.18 $Y2=1.285
r91 37 39 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.18 $Y=0.995
+ $X2=1.18 $Y2=1.285
r92 36 42 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.445 $Y=0.91
+ $X2=0.27 $Y2=0.91
r93 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.015 $Y=0.91
+ $X2=1.18 $Y2=0.995
r94 35 36 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.015 $Y=0.91
+ $X2=0.445 $Y2=0.91
r95 31 44 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.27 $Y=2.2 $X2=0.27
+ $Y2=2.19
r96 31 33 23.0489 $w=3.48e-07 $l=7e-07 $layer=LI1_cond $X=0.27 $Y=2.2 $X2=0.27
+ $Y2=2.9
r97 29 42 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.18 $Y=0.995
+ $X2=0.27 $Y2=0.91
r98 29 45 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.18 $Y=0.995
+ $X2=0.18 $Y2=2.025
r99 25 42 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=0.825
+ $X2=0.27 $Y2=0.91
r100 25 27 11.6891 $w=3.48e-07 $l=3.55e-07 $layer=LI1_cond $X=0.27 $Y=0.825
+ $X2=0.27 $Y2=0.47
r101 19 24 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.725 $Y=1.545
+ $X2=1.725 $Y2=1.42
r102 19 21 203.732 $w=2.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.725 $Y=1.545
+ $X2=1.725 $Y2=2.365
r103 17 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.675 $Y=1.27
+ $X2=1.675 $Y2=1.195
r104 17 24 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.675 $Y=1.27
+ $X2=1.675 $Y2=1.42
r105 13 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.675 $Y=1.12
+ $X2=1.675 $Y2=1.195
r106 13 15 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.675 $Y=1.12
+ $X2=1.675 $Y2=0.445
r107 11 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.6 $Y=1.195
+ $X2=1.675 $Y2=1.195
r108 11 49 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.6 $Y=1.195
+ $X2=1.36 $Y2=1.195
r109 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.12
+ $X2=1.285 $Y2=1.285
r110 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.285 $Y=1.12
+ $X2=1.285 $Y2=0.445
r111 2 44 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r112 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r113 1 27 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_LP%B 3 6 9 13 15 16 20 24
c60 3 0 7.0949e-20 $X=2.255 $Y=1.135
r61 22 24 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=2.975 $Y=1.77
+ $X2=3.015 $Y2=1.77
r62 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.77 $X2=2.975 $Y2=1.77
r63 19 22 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.615 $Y=1.77
+ $X2=2.975 $Y2=1.77
r64 19 20 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.615 $Y=1.77
+ $X2=2.54 $Y2=1.77
r65 15 16 12.0867 $w=4.73e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.912
+ $X2=3.6 $Y2=1.912
r66 15 23 3.65119 $w=4.73e-07 $l=1.45e-07 $layer=LI1_cond $X=3.12 $Y=1.912
+ $X2=2.975 $Y2=1.912
r67 11 24 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.015 $Y=1.935
+ $X2=3.015 $Y2=1.77
r68 11 13 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.015 $Y=1.935
+ $X2=3.015 $Y2=2.595
r69 7 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=1.605
+ $X2=2.615 $Y2=1.77
r70 7 9 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.615 $Y=1.605 $X2=2.615
+ $Y2=1.135
r71 6 20 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.33 $Y=1.68 $X2=2.54
+ $Y2=1.68
r72 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.255 $Y=1.605
+ $X2=2.33 $Y2=1.68
r73 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.255 $Y=1.605 $X2=2.255
+ $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_LP%A 1 3 6 8 10 11 12 19
c46 12 0 1.53875e-20 $X=3.6 $Y=1.295
c47 6 0 1.96911e-19 $X=3.505 $Y=2.595
r48 19 20 1.33518 $w=3.61e-07 $l=1e-08 $layer=POLY_cond $X=3.505 $Y=1.262
+ $X2=3.515 $Y2=1.262
r49 17 19 23.3657 $w=3.61e-07 $l=1.75e-07 $layer=POLY_cond $X=3.33 $Y=1.262
+ $X2=3.505 $Y2=1.262
r50 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.33
+ $Y=1.2 $X2=3.33 $Y2=1.2
r51 15 17 27.3712 $w=3.61e-07 $l=2.05e-07 $layer=POLY_cond $X=3.125 $Y=1.262
+ $X2=3.33 $Y2=1.262
r52 12 18 8.29759 $w=3.73e-07 $l=2.7e-07 $layer=LI1_cond $X=3.6 $Y=1.222
+ $X2=3.33 $Y2=1.222
r53 11 18 6.45368 $w=3.73e-07 $l=2.1e-07 $layer=LI1_cond $X=3.12 $Y=1.222
+ $X2=3.33 $Y2=1.222
r54 8 20 23.3725 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=3.515 $Y=1.035
+ $X2=3.515 $Y2=1.262
r55 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.515 $Y=1.035
+ $X2=3.515 $Y2=0.715
r56 4 19 11.4134 $w=2.5e-07 $l=2.28e-07 $layer=POLY_cond $X=3.505 $Y=1.49
+ $X2=3.505 $Y2=1.262
r57 4 6 274.541 $w=2.5e-07 $l=1.105e-06 $layer=POLY_cond $X=3.505 $Y=1.49
+ $X2=3.505 $Y2=2.595
r58 1 15 23.3725 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=3.125 $Y=1.035
+ $X2=3.125 $Y2=1.262
r59 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.125 $Y=1.035
+ $X2=3.125 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_LP%A_350_47# 1 2 3 12 16 20 24 26 28 31 33 34
+ 36 37 38 40 43 44 47 51 57 62
c138 62 0 5.55614e-20 $X=2.91 $Y=0.67
r139 59 62 5.29501 $w=3.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.74 $Y=0.67
+ $X2=2.91 $Y2=0.67
r140 56 57 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.545 $Y=1.41
+ $X2=2.74 $Y2=1.41
r141 48 51 7.87034 $w=4.08e-07 $l=2.8e-07 $layer=LI1_cond $X=1.61 $Y=0.47
+ $X2=1.89 $Y2=0.47
r142 47 64 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.98 $Y=2.33
+ $X2=3.98 $Y2=1.895
r143 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.06
+ $Y=1.39 $X2=4.06 $Y2=1.39
r144 41 64 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=1.73
+ $X2=4.06 $Y2=1.895
r145 41 43 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=4.06 $Y=1.73
+ $X2=4.06 $Y2=1.39
r146 40 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=1.325
+ $X2=2.74 $Y2=1.41
r147 39 59 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.74 $Y=0.855
+ $X2=2.74 $Y2=0.67
r148 39 40 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.74 $Y=0.855
+ $X2=2.74 $Y2=1.325
r149 37 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.895 $Y=2.415
+ $X2=3.98 $Y2=2.33
r150 37 38 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=3.895 $Y=2.415
+ $X2=2.63 $Y2=2.415
r151 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.545 $Y=2.33
+ $X2=2.63 $Y2=2.415
r152 35 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=1.495
+ $X2=2.545 $Y2=1.41
r153 35 36 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.545 $Y=1.495
+ $X2=2.545 $Y2=2.33
r154 33 56 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=1.41
+ $X2=2.545 $Y2=1.41
r155 33 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.46 $Y=1.41
+ $X2=2.155 $Y2=1.41
r156 29 34 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=1.41
+ $X2=2.155 $Y2=1.41
r157 29 53 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.99 $Y=1.41
+ $X2=1.61 $Y2=1.41
r158 29 31 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=1.99 $Y=1.495
+ $X2=1.99 $Y2=2.01
r159 28 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=1.325
+ $X2=1.61 $Y2=1.41
r160 27 48 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.61 $Y=0.675
+ $X2=1.61 $Y2=0.47
r161 27 28 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.61 $Y=0.675
+ $X2=1.61 $Y2=1.325
r162 25 44 42.4067 $w=4e-07 $l=3.05e-07 $layer=POLY_cond $X=4.07 $Y=1.695
+ $X2=4.07 $Y2=1.39
r163 25 26 35.5859 $w=4e-07 $l=2e-07 $layer=POLY_cond $X=4.07 $Y=1.695 $X2=4.07
+ $Y2=1.895
r164 24 44 2.08558 $w=4e-07 $l=1.5e-08 $layer=POLY_cond $X=4.07 $Y=1.375
+ $X2=4.07 $Y2=1.39
r165 16 26 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=4.145 $Y=2.595
+ $X2=4.145 $Y2=1.895
r166 10 24 24.4565 $w=4e-07 $l=1.5e-07 $layer=POLY_cond $X=4.125 $Y=1.225
+ $X2=4.125 $Y2=1.375
r167 10 20 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.305 $Y=1.225
+ $X2=4.305 $Y2=0.715
r168 10 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.945 $Y=1.225
+ $X2=3.945 $Y2=0.715
r169 3 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.85
+ $Y=1.865 $X2=1.99 $Y2=2.01
r170 2 62 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=2.69
+ $Y=0.925 $X2=2.91 $Y2=0.67
r171 1 51 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.235 $X2=1.89 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_LP%VPWR 1 2 11 17 20 21 22 32 33 36
r47 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r49 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r50 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r51 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 26 29 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r55 24 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 22 30 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 22 27 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 20 29 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.605 $Y=3.33 $X2=3.6
+ $Y2=3.33
r59 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.77 $Y2=3.33
r60 19 32 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=3.77 $Y2=3.33
r62 15 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=3.245
+ $X2=3.77 $Y2=3.33
r63 15 17 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=3.77 $Y=3.245
+ $X2=3.77 $Y2=2.895
r64 11 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.19 $X2=0.81
+ $Y2=2.9
r65 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245 $X2=0.81
+ $Y2=3.33
r66 9 14 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.9
r67 2 17 600 $w=1.7e-07 $l=8.67179e-07 $layer=licon1_PDIFF $count=1 $X=3.63
+ $Y=2.095 $X2=3.77 $Y2=2.895
r68 1 14 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.9
r69 1 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_LP%A_263_373# 1 2 9 13 14 16
r34 16 18 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=2.87
+ $X2=2.75 $Y2=2.98
r35 13 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=2.98
+ $X2=2.75 $Y2=2.98
r36 13 14 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.585 $Y=2.98
+ $X2=1.625 $Y2=2.98
r37 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.46 $Y=2.01 $X2=1.46
+ $Y2=2.72
r38 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.46 $Y=2.895
+ $X2=1.625 $Y2=2.98
r39 7 12 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.46 $Y=2.895
+ $X2=1.46 $Y2=2.72
r40 2 16 600 $w=1.7e-07 $l=8.44393e-07 $layer=licon1_PDIFF $count=1 $X=2.605
+ $Y=2.095 $X2=2.75 $Y2=2.87
r41 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.865 $X2=1.46 $Y2=2.72
r42 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.865 $X2=1.46 $Y2=2.01
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_LP%X 1 2 7 8 9 10 11 12 13 38 45
c26 13 0 1.62489e-19 $X=4.56 $Y=2.775
c27 11 0 3.44213e-20 $X=4.475 $Y=1.95
r28 45 46 1.57618 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=4.52 $Y=0.925 $X2=4.52
+ $Y2=0.945
r29 39 50 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=4.465 $Y=2.295
+ $X2=4.465 $Y2=2.24
r30 38 48 1.92074 $w=2.38e-07 $l=4e-08 $layer=LI1_cond $X=4.565 $Y=2.035
+ $X2=4.565 $Y2=2.075
r31 23 28 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=4.52 $Y=0.78
+ $X2=4.52 $Y2=0.715
r32 13 40 3.09184 $w=4.4e-07 $l=1.05e-07 $layer=LI1_cond $X=4.465 $Y=2.775
+ $X2=4.465 $Y2=2.67
r33 12 40 6.94085 $w=4.38e-07 $l=2.65e-07 $layer=LI1_cond $X=4.465 $Y=2.405
+ $X2=4.465 $Y2=2.67
r34 12 39 2.88111 $w=4.38e-07 $l=1.1e-07 $layer=LI1_cond $X=4.465 $Y=2.405
+ $X2=4.465 $Y2=2.295
r35 11 50 3.74544 $w=4.38e-07 $l=1.43e-07 $layer=LI1_cond $X=4.465 $Y=2.097
+ $X2=4.465 $Y2=2.24
r36 11 48 2.94049 $w=4.38e-07 $l=2.2e-08 $layer=LI1_cond $X=4.465 $Y=2.097
+ $X2=4.465 $Y2=2.075
r37 11 38 1.10442 $w=2.38e-07 $l=2.3e-08 $layer=LI1_cond $X=4.565 $Y=2.012
+ $X2=4.565 $Y2=2.035
r38 10 11 16.6624 $w=2.38e-07 $l=3.47e-07 $layer=LI1_cond $X=4.565 $Y=1.665
+ $X2=4.565 $Y2=2.012
r39 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.565 $Y=1.295
+ $X2=4.565 $Y2=1.665
r40 8 45 1.15244 $w=3.28e-07 $l=3.3e-08 $layer=LI1_cond $X=4.52 $Y=0.892
+ $X2=4.52 $Y2=0.925
r41 8 23 3.91132 $w=3.28e-07 $l=1.12e-07 $layer=LI1_cond $X=4.52 $Y=0.892
+ $X2=4.52 $Y2=0.78
r42 8 9 15.2699 $w=2.38e-07 $l=3.18e-07 $layer=LI1_cond $X=4.565 $Y=0.977
+ $X2=4.565 $Y2=1.295
r43 8 46 1.53659 $w=2.38e-07 $l=3.2e-08 $layer=LI1_cond $X=4.565 $Y=0.977
+ $X2=4.565 $Y2=0.945
r44 7 28 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.52 $Y=0.555 $X2=4.52
+ $Y2=0.715
r45 2 50 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.27
+ $Y=2.095 $X2=4.41 $Y2=2.24
r46 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.505 $X2=4.52 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_LP%VGND 1 2 3 12 14 19 22 25 26 27 29 38 44 45
+ 48 51
r78 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r79 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r80 45 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r81 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r82 42 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=3.73
+ $Y2=0
r83 42 44 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=4.56
+ $Y2=0
r84 41 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r85 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r86 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.565 $Y=0 $X2=3.73
+ $Y2=0
r87 38 40 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=3.565 $Y=0 $X2=2.64
+ $Y2=0
r88 37 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r89 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r90 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r91 34 36 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=2.16
+ $Y2=0
r92 32 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r93 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r94 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r95 29 31 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r96 27 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r97 27 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r98 25 36 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.16
+ $Y2=0
r99 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.32
+ $Y2=0
r100 24 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.405 $Y=0
+ $X2=2.64 $Y2=0
r101 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.32
+ $Y2=0
r102 20 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=0.085
+ $X2=3.73 $Y2=0
r103 20 22 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=3.73 $Y=0.085
+ $X2=3.73 $Y2=0.67
r104 18 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.32 $Y=0.085
+ $X2=2.32 $Y2=0
r105 18 19 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.32 $Y=0.085
+ $X2=2.32 $Y2=0.895
r106 14 19 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.235 $Y=1.02
+ $X2=2.32 $Y2=0.895
r107 14 16 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=2.235 $Y=1.02
+ $X2=2.04 $Y2=1.02
r108 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r109 10 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.43
r110 3 22 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.505 $X2=3.73 $Y2=0.67
r111 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.925 $X2=2.04 $Y2=1.06
r112 1 12 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.235 $X2=1.07 $Y2=0.43
.ends

