* File: sky130_fd_sc_lp__isobufsrc_2.pex.spice
* Created: Fri Aug 28 10:41:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_2%A 1 3 6 8 15
r25 13 15 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.72 $Y=1.35
+ $X2=0.815 $Y2=1.35
r26 10 13 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.54 $Y=1.35 $X2=0.72
+ $Y2=1.35
r27 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.35 $X2=0.72 $Y2=1.35
r28 4 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.815 $Y=1.515
+ $X2=0.815 $Y2=1.35
r29 4 6 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.815 $Y=1.515
+ $X2=0.815 $Y2=2.045
r30 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.185
+ $X2=0.54 $Y2=1.35
r31 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=1.185 $X2=0.54
+ $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_2%SLEEP 3 7 10 14 15 17 21 23 24 29 31 34
+ 43
c80 17 0 8.67399e-20 $X=2.685 $Y=1.16
r81 29 32 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.292 $Y=1.35
+ $X2=1.292 $Y2=1.515
r82 29 31 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.292 $Y=1.35
+ $X2=1.292 $Y2=1.185
r83 24 43 6.27016 $w=3.58e-07 $l=9.5e-08 $layer=LI1_cond $X=1.68 $Y=1.255
+ $X2=1.775 $Y2=1.255
r84 23 24 10.1518 $w=5.28e-07 $l=3.95e-07 $layer=LI1_cond $X=1.2 $Y=1.255
+ $X2=1.595 $Y2=1.255
r85 23 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.35 $X2=1.265 $Y2=1.35
r86 21 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.72 $Y=1.35
+ $X2=2.72 $Y2=1.515
r87 21 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.72 $Y=1.35
+ $X2=2.72 $Y2=1.185
r88 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.72
+ $Y=1.35 $X2=2.72 $Y2=1.35
r89 17 20 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=2.685 $Y=1.16
+ $X2=2.685 $Y2=1.35
r90 15 17 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.555 $Y=1.16
+ $X2=2.685 $Y2=1.16
r91 15 43 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.555 $Y=1.16
+ $X2=1.775 $Y2=1.16
r92 14 34 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.675 $Y=0.655
+ $X2=2.675 $Y2=1.185
r93 10 35 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.63 $Y=2.465
+ $X2=2.63 $Y2=1.515
r94 7 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.385 $Y=0.655
+ $X2=1.385 $Y2=1.185
r95 3 32 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.34 $Y=2.465
+ $X2=1.34 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_2%A_40_131# 1 2 9 13 17 21 25 27 33 35 43
c75 43 0 8.67399e-20 $X=2.2 $Y=1.505
r76 43 44 6.77812 $w=3.2e-07 $l=4.5e-08 $layer=POLY_cond $X=2.2 $Y=1.505
+ $X2=2.245 $Y2=1.505
r77 40 41 6.77812 $w=3.2e-07 $l=4.5e-08 $layer=POLY_cond $X=1.77 $Y=1.505
+ $X2=1.815 $Y2=1.505
r78 36 43 13.5562 $w=3.2e-07 $l=9e-08 $layer=POLY_cond $X=2.11 $Y=1.505 $X2=2.2
+ $Y2=1.505
r79 36 41 44.4344 $w=3.2e-07 $l=2.95e-07 $layer=POLY_cond $X=2.11 $Y=1.505
+ $X2=1.815 $Y2=1.505
r80 35 38 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.11 $Y=1.51
+ $X2=2.11 $Y2=1.77
r81 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.51 $X2=2.11 $Y2=1.51
r82 32 33 8.07799 $w=5.23e-07 $l=9.5e-08 $layer=LI1_cond $X=0.6 $Y=1.947
+ $X2=0.695 $Y2=1.947
r83 27 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=1.77
+ $X2=2.11 $Y2=1.77
r84 27 33 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.945 $Y=1.77
+ $X2=0.695 $Y2=1.77
r85 23 32 6.94865 $w=5.23e-07 $l=3.05e-07 $layer=LI1_cond $X=0.295 $Y=1.947
+ $X2=0.6 $Y2=1.947
r86 23 25 35.0001 $w=2.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.295 $Y=1.685
+ $X2=0.295 $Y2=0.865
r87 19 44 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.245 $Y=1.345
+ $X2=2.245 $Y2=1.505
r88 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.245 $Y=1.345
+ $X2=2.245 $Y2=0.655
r89 15 43 20.4921 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.2 $Y=1.675 $X2=2.2
+ $Y2=1.505
r90 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.2 $Y=1.675 $X2=2.2
+ $Y2=2.465
r91 11 41 20.4921 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.815 $Y=1.335
+ $X2=1.815 $Y2=1.505
r92 11 13 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.815 $Y=1.335
+ $X2=1.815 $Y2=0.655
r93 7 40 20.4921 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.77 $Y=1.675
+ $X2=1.77 $Y2=1.505
r94 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.77 $Y=1.675 $X2=1.77
+ $Y2=2.465
r95 2 32 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.475
+ $Y=1.835 $X2=0.6 $Y2=2.045
r96 1 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.655 $X2=0.325 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_2%VPWR 1 2 9 15 18 19 20 22 32 33 36
r33 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r34 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 27 36 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.057 $Y2=3.33
r38 27 29 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 25 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 22 36 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.865 $Y=3.33
+ $X2=1.057 $Y2=3.33
r42 22 24 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.865 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 20 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 18 29 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r46 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=3.33
+ $X2=2.845 $Y2=3.33
r47 17 32 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.01 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=3.33
+ $X2=2.845 $Y2=3.33
r49 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=3.245
+ $X2=2.845 $Y2=3.33
r50 13 15 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=2.845 $Y=3.245
+ $X2=2.845 $Y2=2.47
r51 9 12 13.0211 $w=3.83e-07 $l=4.35e-07 $layer=LI1_cond $X=1.057 $Y=2.11
+ $X2=1.057 $Y2=2.545
r52 7 36 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.057 $Y=3.245
+ $X2=1.057 $Y2=3.33
r53 7 12 20.9535 $w=3.83e-07 $l=7e-07 $layer=LI1_cond $X=1.057 $Y=3.245
+ $X2=1.057 $Y2=2.545
r54 2 15 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=2.705
+ $Y=1.835 $X2=2.845 $Y2=2.47
r55 1 12 300 $w=1.7e-07 $l=8.19115e-07 $layer=licon1_PDIFF $count=2 $X=0.89
+ $Y=1.835 $X2=1.125 $Y2=2.545
r56 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.89
+ $Y=1.835 $X2=1.03 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_2%A_283_367# 1 2 7 9 11 15
r14 13 15 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=2.415 $Y=2.895
+ $X2=2.415 $Y2=2.53
r15 12 18 3.89832 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=1.65 $Y=2.985
+ $X2=1.535 $Y2=2.985
r16 11 13 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=2.32 $Y=2.985
+ $X2=2.415 $Y2=2.895
r17 11 12 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.32 $Y=2.985
+ $X2=1.65 $Y2=2.985
r18 7 18 3.05086 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=1.535 $Y=2.895 $X2=1.535
+ $Y2=2.985
r19 7 9 35.3249 $w=2.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.535 $Y=2.895
+ $X2=1.535 $Y2=2.19
r20 2 15 300 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=1.835 $X2=2.415 $Y2=2.53
r21 1 18 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.415
+ $Y=1.835 $X2=1.555 $Y2=2.91
r22 1 9 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.415
+ $Y=1.835 $X2=1.555 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_2%X 1 2 3 10 12 14 18 22 24 29 31 32 33 34
+ 35 42 43 45
r62 42 45 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=3.13 $Y=0.905
+ $X2=3.13 $Y2=0.925
r63 35 43 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=2.11 $X2=3.13
+ $Y2=2.025
r64 35 43 1.5101 $w=2.88e-07 $l=3.8e-08 $layer=LI1_cond $X=3.13 $Y=1.987
+ $X2=3.13 $Y2=2.025
r65 34 35 12.7961 $w=2.88e-07 $l=3.22e-07 $layer=LI1_cond $X=3.13 $Y=1.665
+ $X2=3.13 $Y2=1.987
r66 33 34 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=1.295
+ $X2=3.13 $Y2=1.665
r67 32 42 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.82 $X2=3.13
+ $Y2=0.905
r68 32 33 13.4319 $w=2.88e-07 $l=3.38e-07 $layer=LI1_cond $X=3.13 $Y=0.957
+ $X2=3.13 $Y2=1.295
r69 32 45 1.27166 $w=2.88e-07 $l=3.2e-08 $layer=LI1_cond $X=3.13 $Y=0.957
+ $X2=3.13 $Y2=0.925
r70 25 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.555 $Y=0.82
+ $X2=2.46 $Y2=0.82
r71 24 32 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.985 $Y=0.82
+ $X2=3.13 $Y2=0.82
r72 24 25 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.985 $Y=0.82
+ $X2=2.555 $Y2=0.82
r73 20 31 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.735
+ $X2=2.46 $Y2=0.82
r74 20 22 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=2.46 $Y=0.735
+ $X2=2.46 $Y2=0.42
r75 19 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=2.11
+ $X2=1.985 $Y2=2.11
r76 18 35 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.985 $Y=2.11
+ $X2=3.13 $Y2=2.11
r77 18 19 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.985 $Y=2.11
+ $X2=2.15 $Y2=2.11
r78 15 27 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.695 $Y=0.82
+ $X2=1.565 $Y2=0.82
r79 14 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.365 $Y=0.82
+ $X2=2.46 $Y2=0.82
r80 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.365 $Y=0.82
+ $X2=1.695 $Y2=0.82
r81 10 27 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=0.735
+ $X2=1.565 $Y2=0.82
r82 10 12 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.565 $Y=0.735
+ $X2=1.565 $Y2=0.42
r83 3 29 300 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=2 $X=1.845
+ $Y=1.835 $X2=1.985 $Y2=2.11
r84 2 31 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=2.32
+ $Y=0.235 $X2=2.46 $Y2=0.82
r85 2 22 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.32
+ $Y=0.235 $X2=2.46 $Y2=0.42
r86 1 27 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=1.46
+ $Y=0.235 $X2=1.6 $Y2=0.82
r87 1 12 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.46
+ $Y=0.235 $X2=1.6 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_2%VGND 1 2 3 11 13 16 20 25 26 27 28 29 30
+ 32 46 48
r61 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r62 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r63 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r64 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r65 37 48 13.073 $w=1.7e-07 $l=3.23e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=0.942
+ $Y2=0
r66 37 39 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.68
+ $Y2=0
r67 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r68 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r69 32 48 13.073 $w=1.7e-07 $l=3.22e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.942
+ $Y2=0
r70 32 34 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r71 30 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r72 30 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r73 30 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 28 42 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.64
+ $Y2=0
r75 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.89
+ $Y2=0
r76 27 45 4.66471 $w=1.7e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=0 $X2=3.12
+ $Y2=0
r77 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=2.89
+ $Y2=0
r78 25 39 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.68
+ $Y2=0
r79 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.03
+ $Y2=0
r80 24 42 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.64
+ $Y2=0
r81 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.03
+ $Y2=0
r82 18 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=0.085
+ $X2=2.89 $Y2=0
r83 18 20 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.89 $Y=0.085
+ $X2=2.89 $Y2=0.44
r84 14 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0
r85 14 16 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0.44
r86 11 23 5.80021 $w=6.45e-07 $l=2.87e-07 $layer=LI1_cond $X=0.942 $Y=0.563
+ $X2=0.942 $Y2=0.85
r87 11 13 3.39352 $w=6.43e-07 $l=1.83e-07 $layer=LI1_cond $X=0.942 $Y=0.563
+ $X2=0.942 $Y2=0.38
r88 10 48 2.68498 $w=6.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.942 $Y=0.085
+ $X2=0.942 $Y2=0
r89 10 13 5.47044 $w=6.43e-07 $l=2.95e-07 $layer=LI1_cond $X=0.942 $Y=0.085
+ $X2=0.942 $Y2=0.38
r90 3 20 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.75
+ $Y=0.235 $X2=2.89 $Y2=0.44
r91 2 16 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.235 $X2=2.03 $Y2=0.44
r92 1 23 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=0.655 $X2=0.755 $Y2=0.85
r93 1 13 91 $w=1.7e-07 $l=3.67083e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=0.655 $X2=0.83 $Y2=0.38
.ends

