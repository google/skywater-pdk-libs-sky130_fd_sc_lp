* File: sky130_fd_sc_lp__buflp_8.spice
* Created: Wed Sep  2 09:36:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__buflp_8.pex.spice"
.subckt sky130_fd_sc_lp__buflp_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_A_114_47#_M1003_d N_A_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75009.8 A=0.126 P=1.98 MULT=1
MM1006 N_A_114_47#_M1003_d N_A_M1006_g N_A_27_47#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.6
+ SB=75009.3 A=0.126 P=1.98 MULT=1
MM1008 N_A_114_47#_M1008_d N_A_M1008_g N_A_27_47#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75008.9 A=0.126 P=1.98 MULT=1
MM1000 N_A_114_47#_M1008_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75008.4 A=0.126 P=1.98 MULT=1
MM1024 N_A_114_47#_M1024_d N_A_M1024_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75008
+ A=0.126 P=1.98 MULT=1
MM1027 N_A_114_47#_M1024_d N_A_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75007.6 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1027_s N_A_27_47#_M1001_g N_A_644_47#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75007.1 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A_27_47#_M1012_g N_A_644_47#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75006.7 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1012_d N_A_27_47#_M1013_g N_A_644_47#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.7
+ SB=75006.3 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1019_d N_A_27_47#_M1019_g N_A_644_47#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.168 AS=0.1176 PD=1.24 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.1
+ SB=75005.8 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1019_d N_A_27_47#_M1022_g N_A_644_47#_M1022_s VNB NSHORT L=0.15
+ W=0.84 AD=0.168 AS=0.1176 PD=1.24 PS=1.12 NRD=17.136 NRS=0 M=1 R=5.6
+ SA=75004.7 SB=75005.3 A=0.126 P=1.98 MULT=1
MM1029 N_VGND_M1029_d N_A_27_47#_M1029_g N_A_644_47#_M1022_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.1
+ SB=75004.9 A=0.126 P=1.98 MULT=1
MM1040 N_VGND_M1029_d N_A_27_47#_M1040_g N_A_644_47#_M1040_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.6
+ SB=75004.4 A=0.126 P=1.98 MULT=1
MM1010 N_A_644_47#_M1040_s N_A_27_47#_M1010_g N_X_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006
+ SB=75004 A=0.126 P=1.98 MULT=1
MM1017 N_A_644_47#_M1017_d N_A_27_47#_M1017_g N_X_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.4
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1025 N_A_644_47#_M1017_d N_A_27_47#_M1025_g N_X_M1025_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.9
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1028 N_A_644_47#_M1028_d N_A_27_47#_M1028_g N_X_M1025_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75007.3
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1031 N_A_644_47#_M1028_d N_A_27_47#_M1031_g N_X_M1031_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75007.8
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1033 N_A_644_47#_M1033_d N_A_27_47#_M1033_g N_X_M1031_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=9.996 NRS=0 M=1 R=5.6 SA=75008.3
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1036 N_A_644_47#_M1033_d N_A_27_47#_M1036_g N_X_M1036_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75008.8
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1039 N_A_644_47#_M1039_d N_A_27_47#_M1039_g N_X_M1036_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1386 AS=0.147 PD=1.17 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75009.3
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1043 N_VGND_M1043_d N_A_27_47#_M1043_g N_A_644_47#_M1039_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2562 AS=0.1386 PD=2.29 PS=1.17 NRD=2.856 NRS=7.14 M=1 R=5.6
+ SA=75009.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1020 N_A_114_367#_M1020_d N_A_M1020_g N_A_27_47#_M1020_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75009.8 A=0.189 P=2.82 MULT=1
MM1026 N_A_114_367#_M1020_d N_A_M1026_g N_A_27_47#_M1026_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75009.3 A=0.189 P=2.82 MULT=1
MM1041 N_A_114_367#_M1041_d N_A_M1041_g N_A_27_47#_M1026_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75008.9 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_A_114_367#_M1041_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75008.5 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1009_d N_A_M1018_g N_A_114_367#_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9 SB=75008
+ A=0.189 P=2.82 MULT=1
MM1042 N_VPWR_M1042_d N_A_M1042_g N_A_114_367#_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1953 AS=0.1764 PD=1.57 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75007.6 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1042_d N_A_27_47#_M1002_g N_A_636_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1953 AS=0.1764 PD=1.57 PS=1.54 NRD=4.6886 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75007.2 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_27_47#_M1005_g N_A_636_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75006.7 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1005_d N_A_27_47#_M1007_g N_A_636_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75006.3 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A_27_47#_M1014_g N_A_636_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75005.9 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1014_d N_A_27_47#_M1021_g N_A_636_367#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75005.4 A=0.189 P=2.82 MULT=1
MM1023 N_VPWR_M1023_d N_A_27_47#_M1023_g N_A_636_367#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005
+ SB=75005 A=0.189 P=2.82 MULT=1
MM1034 N_VPWR_M1023_d N_A_27_47#_M1034_g N_A_636_367#_M1034_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.4
+ SB=75004.6 A=0.189 P=2.82 MULT=1
MM1004 N_A_636_367#_M1034_s N_A_27_47#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2205 PD=1.54 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75005.8 SB=75004.1 A=0.189 P=2.82 MULT=1
MM1011 N_A_636_367#_M1011_d N_A_27_47#_M1011_g N_X_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75006.3 SB=75003.6 A=0.189 P=2.82 MULT=1
MM1015 N_A_636_367#_M1011_d N_A_27_47#_M1015_g N_X_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75006.8 SB=75003.1 A=0.189 P=2.82 MULT=1
MM1016 N_A_636_367#_M1016_d N_A_27_47#_M1016_g N_X_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75007.3 SB=75002.6 A=0.189 P=2.82 MULT=1
MM1030 N_A_636_367#_M1016_d N_A_27_47#_M1030_g N_X_M1030_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75007.8 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1032 N_A_636_367#_M1032_d N_A_27_47#_M1032_g N_X_M1030_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75008.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1037 N_A_636_367#_M1032_d N_A_27_47#_M1037_g N_X_M1037_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75008.8 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1038 N_A_636_367#_M1038_d N_A_27_47#_M1038_g N_X_M1037_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2205 PD=1.54 PS=1.61 NRD=0 NRS=0 M=1 R=8.4 SA=75009.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1035 N_VPWR_M1035_d N_A_27_47#_M1035_g N_A_636_367#_M1038_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75009.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX44_noxref VNB VPB NWDIODE A=20.4031 P=25.61
*
.include "sky130_fd_sc_lp__buflp_8.pxi.spice"
*
.ends
*
*
