* File: sky130_fd_sc_lp__or3_2.spice
* Created: Wed Sep  2 10:30:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or3_2.pex.spice"
.subckt sky130_fd_sc_lp__or3_2  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_C_M1006_g N_A_35_60#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.1113 PD=1.04 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1008 N_A_35_60#_M1008_d N_B_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1302 PD=0.7 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_35_60#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.123333 AS=0.0588 PD=0.926667 PS=0.7 NRD=24.276 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_35_60#_M1005_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.246667 PD=1.12 PS=1.85333 NRD=0 NRS=12.132 M=1 R=5.6 SA=75001.1
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1005_d N_A_35_60#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3679 PD=1.12 PS=2.7 NRD=0 NRS=17.136 M=1 R=5.6 SA=75001.6
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1009 A_132_367# N_C_M1009_g N_A_35_60#_M1009_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.04725 AS=0.1113 PD=0.645 PS=1.37 NRD=26.9693 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1001 A_207_367# N_B_M1001_g A_132_367# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.04725 PD=0.63 PS=0.645 NRD=23.443 NRS=26.9693 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_207_367# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.164325 AS=0.0441 PD=1.0625 PS=0.63 NRD=30.4759 NRS=23.443 M=1 R=2.8
+ SA=75000.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1002_d N_A_35_60#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.492975 AS=0.1764 PD=3.1875 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A_35_60#_M1004_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__or3_2.pxi.spice"
*
.ends
*
*
