* File: sky130_fd_sc_lp__o31ai_1.pex.spice
* Created: Wed Sep  2 10:25:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31AI_1%A1 3 7 9 10 17
c25 9 0 1.35027e-19 $X=0.24 $Y=1.295
r26 14 17 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.375
+ $X2=0.475 $Y2=1.375
r27 9 10 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295 $X2=0.24
+ $Y2=1.665
r28 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.375 $X2=0.27 $Y2=1.375
r29 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=1.375
r30 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=2.465
r31 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.21
+ $X2=0.475 $Y2=1.375
r32 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.475 $Y=1.21
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_1%A2 3 7 9 10 11 12 19 20
c42 19 0 1.35027e-19 $X=0.925 $Y=1.51
r43 20 35 5.49189 $w=4.03e-07 $l=1.93e-07 $layer=LI1_cond $X=0.925 $Y=1.547
+ $X2=0.732 $Y2=1.547
r44 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.675
r45 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.345
r46 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.51 $X2=0.925 $Y2=1.51
r47 11 12 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.732 $Y=2.405
+ $X2=0.732 $Y2=2.775
r48 10 11 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.732 $Y=2.035
+ $X2=0.732 $Y2=2.405
r49 9 35 0.341465 $w=4.03e-07 $l=1.2e-08 $layer=LI1_cond $X=0.72 $Y=1.547
+ $X2=0.732 $Y2=1.547
r50 9 35 3.01869 $w=2.75e-07 $l=2.03e-07 $layer=LI1_cond $X=0.732 $Y=1.75
+ $X2=0.732 $Y2=1.547
r51 9 10 9.05215 $w=4.43e-07 $l=2.85e-07 $layer=LI1_cond $X=0.732 $Y=1.75
+ $X2=0.732 $Y2=2.035
r52 7 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.905 $Y=0.655
+ $X2=0.905 $Y2=1.345
r53 3 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.835 $Y=2.465
+ $X2=0.835 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_1%A3 3 7 9 10 17
c34 17 0 1.06993e-19 $X=1.69 $Y=1.51
r35 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.51 $X2=1.69 $Y2=1.51
r36 15 17 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.675 $Y=1.51
+ $X2=1.69 $Y2=1.51
r37 13 15 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=1.375 $Y=1.51
+ $X2=1.675 $Y2=1.51
r38 10 18 14.444 $w=3.73e-07 $l=4.7e-07 $layer=LI1_cond $X=2.16 $Y=1.562
+ $X2=1.69 $Y2=1.562
r39 9 18 0.307318 $w=3.73e-07 $l=1e-08 $layer=LI1_cond $X=1.68 $Y=1.562 $X2=1.69
+ $Y2=1.562
r40 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.345
+ $X2=1.675 $Y2=1.51
r41 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.675 $Y=1.345
+ $X2=1.675 $Y2=0.655
r42 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.675
+ $X2=1.375 $Y2=1.51
r43 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.375 $Y=1.675
+ $X2=1.375 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_1%B1 3 7 10 11 14 15
c30 15 0 1.06993e-19 $X=2.59 $Y=1.46
r31 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.46 $X2=2.59 $Y2=1.46
r32 11 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.46
r33 9 14 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.25 $Y=1.46 $X2=2.59
+ $Y2=1.46
r34 9 10 5.03009 $w=3.3e-07 $l=8.3e-08 $layer=POLY_cond $X=2.25 $Y=1.46
+ $X2=2.167 $Y2=1.46
r35 5 10 37.0704 $w=1.5e-07 $l=1.68953e-07 $layer=POLY_cond $X=2.175 $Y=1.295
+ $X2=2.167 $Y2=1.46
r36 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.175 $Y=1.295
+ $X2=2.175 $Y2=0.655
r37 1 10 37.0704 $w=1.5e-07 $l=1.68464e-07 $layer=POLY_cond $X=2.16 $Y=1.625
+ $X2=2.167 $Y2=1.46
r38 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.16 $Y=1.625 $X2=2.16
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_1%VPWR 1 2 7 9 15 20 21 22 32 33
r31 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 24 36 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r39 24 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 22 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 22 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 20 29 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 20 21 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=3.33 $X2=2.41
+ $Y2=3.33
r44 19 32 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.54 $Y=3.33 $X2=2.64
+ $Y2=3.33
r45 19 21 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=3.33 $X2=2.41
+ $Y2=3.33
r46 15 18 38.3409 $w=2.58e-07 $l=8.65e-07 $layer=LI1_cond $X=2.41 $Y=2.085
+ $X2=2.41 $Y2=2.95
r47 13 21 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=3.245
+ $X2=2.41 $Y2=3.33
r48 13 18 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.41 $Y=3.245
+ $X2=2.41 $Y2=2.95
r49 9 12 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.26 $Y=2.005
+ $X2=0.26 $Y2=2.95
r50 7 36 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r51 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r52 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.835 $X2=2.375 $Y2=2.95
r53 2 15 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.835 $X2=2.375 $Y2=2.085
r54 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r55 1 9 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_1%Y 1 2 7 8 11 14 15 16
r37 16 32 1.99533 $w=1.068e-06 $l=1.75e-07 $layer=LI1_cond $X=1.575 $Y=2.775
+ $X2=1.575 $Y2=2.95
r38 15 16 4.21869 $w=1.068e-06 $l=3.7e-07 $layer=LI1_cond $X=1.575 $Y=2.405
+ $X2=1.575 $Y2=2.775
r39 14 15 4.21869 $w=1.068e-06 $l=3.7e-07 $layer=LI1_cond $X=1.575 $Y=2.035
+ $X2=1.575 $Y2=2.405
r40 13 14 32.4466 $w=2.73e-07 $l=7.45e-07 $layer=LI1_cond $X=1.265 $Y=1.205
+ $X2=1.265 $Y2=1.95
r41 9 11 27.2597 $w=2.58e-07 $l=6.15e-07 $layer=LI1_cond $X=2.425 $Y=1.035
+ $X2=2.425 $Y2=0.42
r42 8 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.35 $Y=1.12
+ $X2=1.265 $Y2=1.205
r43 7 9 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.295 $Y=1.12
+ $X2=2.425 $Y2=1.035
r44 7 8 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=2.295 $Y=1.12
+ $X2=1.35 $Y2=1.12
r45 2 32 200 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=3 $X=1.45
+ $Y=1.835 $X2=1.59 $Y2=2.95
r46 2 14 200 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=3 $X=1.45
+ $Y=1.835 $X2=1.59 $Y2=2.035
r47 1 11 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.25
+ $Y=0.235 $X2=2.39 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_1%VGND 1 2 7 9 11 23 24 32 35
r40 34 35 10.2213 $w=6.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=0.22
+ $X2=1.625 $Y2=0.22
r41 30 34 5.09804 $w=6.08e-07 $l=2.6e-07 $layer=LI1_cond $X=1.2 $Y=0.22 $X2=1.46
+ $Y2=0.22
r42 30 32 11.986 $w=6.08e-07 $l=2.55e-07 $layer=LI1_cond $X=1.2 $Y=0.22
+ $X2=0.945 $Y2=0.22
r43 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r45 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 21 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r47 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r48 20 35 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.625
+ $Y2=0
r49 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r50 17 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r51 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r52 16 32 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.945
+ $Y2=0
r53 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r54 14 27 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r55 14 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r56 11 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r57 11 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r58 7 27 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r59 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r60 2 34 91 $w=1.7e-07 $l=5.5857e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.235 $X2=1.46 $Y2=0.405
r61 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_1%A_110_47# 1 2 9 11 15 17
r29 17 20 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=0.725 $Y=0.78
+ $X2=0.725 $Y2=0.93
r30 17 18 4.86943 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.78
+ $X2=0.725 $Y2=0.695
r31 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.96 $Y=0.695
+ $X2=1.96 $Y2=0.36
r32 12 17 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.855 $Y=0.78
+ $X2=0.725 $Y2=0.78
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.795 $Y=0.78
+ $X2=1.96 $Y2=0.695
r34 11 12 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.795 $Y=0.78
+ $X2=0.855 $Y2=0.78
r35 9 18 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=0.685 $Y=0.42
+ $X2=0.685 $Y2=0.695
r36 2 15 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=1.75
+ $Y=0.235 $X2=1.96 $Y2=0.36
r37 1 20 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.93
r38 1 9 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

