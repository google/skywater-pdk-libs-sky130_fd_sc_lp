# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__and4bb_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__and4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.425000 0.550000 1.750000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.945000 0.255000 4.645000 0.650000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.335000 2.690000 3.735000 3.020000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.410000 1.180000 4.185000 1.415000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.080000 0.255000 1.310000 1.935000 ;
        RECT 1.080000 1.935000 1.445000 2.215000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.800000 0.085000 ;
        RECT 0.525000  0.085000 0.910000 0.905000 ;
        RECT 1.480000  0.085000 1.810000 0.825000 ;
        RECT 3.435000  0.085000 3.775000 0.820000 ;
        RECT 3.435000  0.820000 4.145000 1.010000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.800000 3.415000 ;
        RECT 0.685000 2.725000 1.015000 3.245000 ;
        RECT 1.545000 2.725000 2.220000 3.245000 ;
        RECT 1.955000 2.135000 2.220000 2.725000 ;
        RECT 2.985000 2.275000 3.315000 2.520000 ;
        RECT 2.985000 2.520000 3.155000 3.245000 ;
        RECT 3.905000 2.120000 4.185000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.710000 0.355000 1.075000 ;
      RECT 0.095000 1.075000 0.900000 1.245000 ;
      RECT 0.160000 1.920000 0.900000 2.385000 ;
      RECT 0.730000 1.245000 0.900000 1.920000 ;
      RECT 0.730000 2.385000 1.785000 2.555000 ;
      RECT 1.480000 0.995000 2.560000 1.175000 ;
      RECT 1.480000 1.175000 1.750000 1.615000 ;
      RECT 1.615000 1.795000 2.220000 1.965000 ;
      RECT 1.615000 1.965000 1.785000 2.385000 ;
      RECT 1.960000 1.345000 2.220000 1.795000 ;
      RECT 2.125000 0.670000 2.560000 0.995000 ;
      RECT 2.390000 1.175000 2.560000 1.935000 ;
      RECT 2.390000 1.935000 3.735000 2.105000 ;
      RECT 2.390000 2.105000 2.815000 2.450000 ;
      RECT 2.790000 1.245000 3.120000 1.585000 ;
      RECT 2.790000 1.585000 4.685000 1.765000 ;
      RECT 3.485000 2.105000 3.735000 2.450000 ;
      RECT 4.355000 0.820000 4.685000 1.585000 ;
      RECT 4.355000 1.765000 4.685000 2.450000 ;
  END
END sky130_fd_sc_lp__and4bb_2
