# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__mux2i_m
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__mux2i_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.030000 1.580000 2.360000 1.795000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 0.265000 2.150000 0.435000 ;
        RECT 1.355000 0.435000 1.525000 1.210000 ;
        RECT 1.355000 1.210000 1.765000 2.120000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.520000 1.995000 0.690000 2.300000 ;
        RECT 0.520000 2.300000 1.505000 2.470000 ;
        RECT 1.335000 2.470000 1.505000 2.895000 ;
        RECT 1.335000 2.895000 2.465000 3.065000 ;
        RECT 2.295000 2.325000 3.205000 2.495000 ;
        RECT 2.295000 2.495000 2.465000 2.895000 ;
        RECT 2.890000 1.155000 3.205000 2.325000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  0.331800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705000 0.700000 2.245000 1.030000 ;
        RECT 1.710000 2.525000 2.115000 2.715000 ;
        RECT 1.945000 1.975000 2.710000 2.145000 ;
        RECT 1.945000 2.145000 2.115000 2.525000 ;
        RECT 2.075000 1.030000 2.245000 1.055000 ;
        RECT 2.075000 1.055000 2.710000 1.225000 ;
        RECT 2.540000 1.225000 2.710000 1.975000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.360000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 3.550000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.170000  0.795000 0.565000 1.005000 ;
      RECT 0.170000  1.005000 0.340000 1.425000 ;
      RECT 0.170000  1.425000 1.170000 1.755000 ;
      RECT 0.170000  1.755000 0.340000 2.650000 ;
      RECT 0.170000  2.650000 0.645000 2.860000 ;
      RECT 0.745000  0.085000 1.075000 0.875000 ;
      RECT 0.825000  2.655000 1.155000 3.245000 ;
      RECT 2.600000  0.085000 2.930000 0.875000 ;
      RECT 2.790000  2.675000 3.120000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__mux2i_m
END LIBRARY
