* File: sky130_fd_sc_lp__dfbbp_1.pxi.spice
* Created: Wed Sep  2 09:43:07 2020
* 
x_PM_SKY130_FD_SC_LP__DFBBP_1%CLK N_CLK_c_259_n N_CLK_M1018_g N_CLK_c_266_n
+ N_CLK_M1033_g N_CLK_c_261_n N_CLK_c_262_n N_CLK_c_267_n CLK CLK CLK
+ N_CLK_c_263_n N_CLK_c_264_n PM_SKY130_FD_SC_LP__DFBBP_1%CLK
x_PM_SKY130_FD_SC_LP__DFBBP_1%D N_D_c_296_n N_D_c_300_n N_D_c_297_n N_D_M1002_g
+ N_D_c_301_n N_D_M1006_g D D D N_D_c_299_n N_D_c_303_n
+ PM_SKY130_FD_SC_LP__DFBBP_1%D
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_225_47# N_A_225_47#_M1008_s N_A_225_47#_M1011_s
+ N_A_225_47#_M1032_g N_A_225_47#_M1031_g N_A_225_47#_M1013_g
+ N_A_225_47#_M1007_g N_A_225_47#_c_360_n N_A_225_47#_c_361_n
+ N_A_225_47#_c_362_n N_A_225_47#_c_375_n N_A_225_47#_c_376_n
+ N_A_225_47#_c_377_n N_A_225_47#_c_363_n N_A_225_47#_c_378_n
+ N_A_225_47#_c_364_n N_A_225_47#_c_380_n N_A_225_47#_c_381_n
+ N_A_225_47#_c_365_n N_A_225_47#_c_366_n N_A_225_47#_c_367_n
+ N_A_225_47#_c_422_p N_A_225_47#_c_368_n N_A_225_47#_c_369_n
+ PM_SKY130_FD_SC_LP__DFBBP_1%A_225_47#
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_767_21# N_A_767_21#_M1023_d N_A_767_21#_M1030_d
+ N_A_767_21#_M1028_g N_A_767_21#_M1009_g N_A_767_21#_M1026_g
+ N_A_767_21#_c_556_n N_A_767_21#_c_557_n N_A_767_21#_M1012_g
+ N_A_767_21#_c_559_n N_A_767_21#_c_560_n N_A_767_21#_c_601_p
+ N_A_767_21#_c_633_p N_A_767_21#_c_584_n N_A_767_21#_c_612_p
+ N_A_767_21#_c_585_n N_A_767_21#_c_586_n N_A_767_21#_c_561_n
+ N_A_767_21#_c_571_n N_A_767_21#_c_562_n N_A_767_21#_c_563_n
+ N_A_767_21#_c_574_n N_A_767_21#_c_608_p PM_SKY130_FD_SC_LP__DFBBP_1%A_767_21#
x_PM_SKY130_FD_SC_LP__DFBBP_1%SET_B N_SET_B_M1003_g N_SET_B_c_715_n
+ N_SET_B_M1030_g N_SET_B_M1020_g N_SET_B_M1010_g SET_B N_SET_B_c_722_n
+ N_SET_B_c_733_n N_SET_B_c_723_n N_SET_B_c_724_n N_SET_B_c_717_n
+ N_SET_B_c_718_n N_SET_B_c_719_n PM_SKY130_FD_SC_LP__DFBBP_1%SET_B
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_617_47# N_A_617_47#_M1021_d N_A_617_47#_M1032_d
+ N_A_617_47#_M1023_g N_A_617_47#_c_834_n N_A_617_47#_M1015_g
+ N_A_617_47#_c_836_n N_A_617_47#_c_837_n N_A_617_47#_c_838_n
+ N_A_617_47#_c_848_n N_A_617_47#_c_850_n PM_SKY130_FD_SC_LP__DFBBP_1%A_617_47#
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_1091_21# N_A_1091_21#_M1035_s
+ N_A_1091_21#_M1025_s N_A_1091_21#_c_922_n N_A_1091_21#_M1019_g
+ N_A_1091_21#_M1016_g N_A_1091_21#_M1001_g N_A_1091_21#_M1014_g
+ N_A_1091_21#_c_926_n N_A_1091_21#_c_927_n N_A_1091_21#_c_928_n
+ N_A_1091_21#_c_929_n N_A_1091_21#_c_930_n N_A_1091_21#_c_952_n
+ N_A_1091_21#_c_931_n N_A_1091_21#_c_932_n N_A_1091_21#_c_933_n
+ N_A_1091_21#_c_934_n N_A_1091_21#_c_935_n N_A_1091_21#_c_936_n
+ N_A_1091_21#_c_937_n N_A_1091_21#_c_938_n N_A_1091_21#_c_939_n
+ N_A_1091_21#_c_945_n N_A_1091_21#_c_946_n N_A_1091_21#_c_940_n
+ PM_SKY130_FD_SC_LP__DFBBP_1%A_1091_21#
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_114_57# N_A_114_57#_M1018_d N_A_114_57#_M1033_d
+ N_A_114_57#_c_1100_n N_A_114_57#_M1008_g N_A_114_57#_M1011_g
+ N_A_114_57#_c_1103_n N_A_114_57#_c_1104_n N_A_114_57#_c_1114_n
+ N_A_114_57#_c_1115_n N_A_114_57#_c_1105_n N_A_114_57#_M1021_g
+ N_A_114_57#_M1034_g N_A_114_57#_c_1117_n N_A_114_57#_c_1118_n
+ N_A_114_57#_M1017_g N_A_114_57#_c_1120_n N_A_114_57#_M1004_g
+ N_A_114_57#_c_1108_n N_A_114_57#_c_1122_n N_A_114_57#_c_1109_n
+ N_A_114_57#_c_1110_n N_A_114_57#_c_1124_n N_A_114_57#_c_1111_n
+ N_A_114_57#_c_1112_n PM_SKY130_FD_SC_LP__DFBBP_1%A_114_57#
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_1545_332# N_A_1545_332#_M1029_d
+ N_A_1545_332#_M1010_d N_A_1545_332#_M1005_g N_A_1545_332#_M1036_g
+ N_A_1545_332#_M1027_g N_A_1545_332#_M1037_g N_A_1545_332#_c_1259_n
+ N_A_1545_332#_c_1260_n N_A_1545_332#_M1000_g N_A_1545_332#_M1022_g
+ N_A_1545_332#_c_1262_n N_A_1545_332#_c_1272_n N_A_1545_332#_c_1273_n
+ N_A_1545_332#_c_1274_n N_A_1545_332#_c_1275_n N_A_1545_332#_c_1276_n
+ N_A_1545_332#_c_1277_n N_A_1545_332#_c_1263_n N_A_1545_332#_c_1279_n
+ N_A_1545_332#_c_1264_n N_A_1545_332#_c_1281_n N_A_1545_332#_c_1265_n
+ N_A_1545_332#_c_1328_n N_A_1545_332#_c_1266_n N_A_1545_332#_c_1267_n
+ N_A_1545_332#_c_1268_n PM_SKY130_FD_SC_LP__DFBBP_1%A_1545_332#
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_1307_428# N_A_1307_428#_M1013_d
+ N_A_1307_428#_M1017_d N_A_1307_428#_M1029_g N_A_1307_428#_M1038_g
+ N_A_1307_428#_c_1438_n N_A_1307_428#_c_1453_n N_A_1307_428#_c_1439_n
+ N_A_1307_428#_c_1440_n N_A_1307_428#_c_1441_n N_A_1307_428#_c_1442_n
+ N_A_1307_428#_c_1448_n N_A_1307_428#_c_1443_n N_A_1307_428#_c_1444_n
+ N_A_1307_428#_c_1445_n PM_SKY130_FD_SC_LP__DFBBP_1%A_1307_428#
x_PM_SKY130_FD_SC_LP__DFBBP_1%RESET_B N_RESET_B_M1025_g N_RESET_B_M1035_g
+ RESET_B N_RESET_B_c_1560_n N_RESET_B_c_1561_n
+ PM_SKY130_FD_SC_LP__DFBBP_1%RESET_B
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_2317_367# N_A_2317_367#_M1000_s
+ N_A_2317_367#_M1022_s N_A_2317_367#_M1039_g N_A_2317_367#_M1024_g
+ N_A_2317_367#_c_1592_n N_A_2317_367#_c_1600_n N_A_2317_367#_c_1593_n
+ N_A_2317_367#_c_1594_n N_A_2317_367#_c_1595_n N_A_2317_367#_c_1596_n
+ N_A_2317_367#_c_1597_n N_A_2317_367#_c_1598_n
+ PM_SKY130_FD_SC_LP__DFBBP_1%A_2317_367#
x_PM_SKY130_FD_SC_LP__DFBBP_1%VPWR N_VPWR_M1033_s N_VPWR_M1011_d N_VPWR_M1009_d
+ N_VPWR_M1016_d N_VPWR_M1036_d N_VPWR_M1001_d N_VPWR_M1025_d N_VPWR_M1022_d
+ N_VPWR_c_1652_n N_VPWR_c_1653_n N_VPWR_c_1654_n N_VPWR_c_1655_n
+ N_VPWR_c_1656_n N_VPWR_c_1657_n N_VPWR_c_1658_n N_VPWR_c_1659_n
+ N_VPWR_c_1660_n N_VPWR_c_1661_n N_VPWR_c_1662_n N_VPWR_c_1663_n
+ N_VPWR_c_1664_n N_VPWR_c_1665_n N_VPWR_c_1666_n VPWR N_VPWR_c_1667_n
+ N_VPWR_c_1668_n N_VPWR_c_1669_n N_VPWR_c_1670_n N_VPWR_c_1671_n
+ N_VPWR_c_1651_n N_VPWR_c_1673_n N_VPWR_c_1674_n N_VPWR_c_1675_n
+ N_VPWR_c_1676_n PM_SKY130_FD_SC_LP__DFBBP_1%VPWR
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_531_47# N_A_531_47#_M1002_d N_A_531_47#_M1006_d
+ N_A_531_47#_c_1799_n N_A_531_47#_c_1796_n N_A_531_47#_c_1793_n
+ N_A_531_47#_c_1794_n N_A_531_47#_c_1795_n N_A_531_47#_c_1798_n
+ PM_SKY130_FD_SC_LP__DFBBP_1%A_531_47#
x_PM_SKY130_FD_SC_LP__DFBBP_1%Q_N N_Q_N_M1037_d N_Q_N_M1027_d N_Q_N_c_1865_n
+ N_Q_N_c_1866_n N_Q_N_c_1868_n N_Q_N_c_1867_n Q_N Q_N Q_N
+ PM_SKY130_FD_SC_LP__DFBBP_1%Q_N
x_PM_SKY130_FD_SC_LP__DFBBP_1%Q N_Q_M1039_d N_Q_M1024_d N_Q_c_1904_n
+ N_Q_c_1905_n N_Q_c_1901_n Q Q N_Q_c_1902_n Q PM_SKY130_FD_SC_LP__DFBBP_1%Q
x_PM_SKY130_FD_SC_LP__DFBBP_1%VGND N_VGND_M1018_s N_VGND_M1008_d N_VGND_M1028_d
+ N_VGND_M1012_s N_VGND_M1005_d N_VGND_M1035_d N_VGND_M1000_d N_VGND_c_1928_n
+ N_VGND_c_1929_n N_VGND_c_1930_n N_VGND_c_1931_n N_VGND_c_1932_n
+ N_VGND_c_1933_n N_VGND_c_1934_n N_VGND_c_1935_n N_VGND_c_1936_n
+ N_VGND_c_1937_n N_VGND_c_1938_n N_VGND_c_1939_n N_VGND_c_1940_n
+ N_VGND_c_1941_n VGND N_VGND_c_1942_n N_VGND_c_1943_n N_VGND_c_1944_n
+ N_VGND_c_1945_n N_VGND_c_1946_n N_VGND_c_1947_n N_VGND_c_1948_n
+ N_VGND_c_1949_n PM_SKY130_FD_SC_LP__DFBBP_1%VGND
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_917_47# N_A_917_47#_M1003_d N_A_917_47#_M1019_d
+ N_A_917_47#_c_2075_n N_A_917_47#_c_2080_n N_A_917_47#_c_2076_n
+ N_A_917_47#_c_2077_n PM_SKY130_FD_SC_LP__DFBBP_1%A_917_47#
x_PM_SKY130_FD_SC_LP__DFBBP_1%A_1705_54# N_A_1705_54#_M1020_d
+ N_A_1705_54#_M1014_d N_A_1705_54#_c_2105_n
+ PM_SKY130_FD_SC_LP__DFBBP_1%A_1705_54#
cc_1 VNB N_CLK_c_259_n 0.00489886f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=2.18
cc_2 VNB N_CLK_M1018_g 0.0299316f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_3 VNB N_CLK_c_261_n 0.0335688f $X=-0.19 $Y=-0.245 $X2=0.347 $Y2=1.03
cc_4 VNB N_CLK_c_262_n 0.0222535f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.575
cc_5 VNB N_CLK_c_263_n 0.0410503f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_6 VNB N_CLK_c_264_n 0.00298149f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_7 VNB N_D_c_296_n 0.0329536f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.575
cc_8 VNB N_D_c_297_n 0.0216705f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_9 VNB D 0.0151111f $X=-0.19 $Y=-0.245 $X2=0.347 $Y2=0.88
cc_10 VNB N_D_c_299_n 0.0354251f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.255
cc_11 VNB N_A_225_47#_M1031_g 0.055205f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.41
cc_12 VNB N_A_225_47#_M1013_g 0.0242067f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.255
cc_13 VNB N_A_225_47#_c_360_n 0.0158456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_225_47#_c_361_n 0.0170642f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_15 VNB N_A_225_47#_c_362_n 0.0161321f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_16 VNB N_A_225_47#_c_363_n 0.00704797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_225_47#_c_364_n 0.0013649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_225_47#_c_365_n 0.0496142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_225_47#_c_366_n 6.558e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_225_47#_c_367_n 0.00463802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_225_47#_c_368_n 0.0305926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_225_47#_c_369_n 0.00516627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_767_21#_M1028_g 0.0512547f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.725
cc_24 VNB N_A_767_21#_c_556_n 0.00715355f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_25 VNB N_A_767_21#_c_557_n 0.0080337f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_A_767_21#_M1012_g 0.0242948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_767_21#_c_559_n 0.00132918f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_28 VNB N_A_767_21#_c_560_n 0.0224588f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_29 VNB N_A_767_21#_c_561_n 0.00623319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_767_21#_c_562_n 0.00440047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_767_21#_c_563_n 0.046867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_SET_B_M1003_g 0.0403016f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_33 VNB N_SET_B_c_715_n 0.0268952f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_34 VNB N_SET_B_M1020_g 0.0546996f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.03
cc_35 VNB N_SET_B_c_717_n 0.00131955f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_36 VNB N_SET_B_c_718_n 0.0139766f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_37 VNB N_SET_B_c_719_n 3.23736e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_617_47#_M1023_g 0.019726f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.725
cc_39 VNB N_A_617_47#_c_834_n 0.037785f $X=-0.19 $Y=-0.245 $X2=0.347 $Y2=0.88
cc_40 VNB N_A_617_47#_M1015_g 0.0149584f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.41
cc_41 VNB N_A_617_47#_c_836_n 0.00334864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_617_47#_c_837_n 0.00366115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_617_47#_c_838_n 0.0240244f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_44 VNB N_A_1091_21#_c_922_n 0.0201976f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.33
cc_45 VNB N_A_1091_21#_M1016_g 0.017631f $X=-0.19 $Y=-0.245 $X2=0.347 $Y2=1.03
cc_46 VNB N_A_1091_21#_M1001_g 0.0153336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1091_21#_M1014_g 0.0332683f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_48 VNB N_A_1091_21#_c_926_n 0.0159086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1091_21#_c_927_n 0.00361822f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_50 VNB N_A_1091_21#_c_928_n 0.0515332f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_51 VNB N_A_1091_21#_c_929_n 0.00679306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1091_21#_c_930_n 0.00232304f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_53 VNB N_A_1091_21#_c_931_n 0.0141496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1091_21#_c_932_n 0.0010739f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=2.035
cc_55 VNB N_A_1091_21#_c_933_n 7.19767e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1091_21#_c_934_n 0.0204823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1091_21#_c_935_n 0.00173127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1091_21#_c_936_n 0.00324996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1091_21#_c_937_n 0.0166604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1091_21#_c_938_n 0.00483494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1091_21#_c_939_n 0.0390063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1091_21#_c_940_n 0.00131128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_114_57#_c_1100_n 0.0306328f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.725
cc_64 VNB N_A_114_57#_M1008_g 0.0587055f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.41
cc_65 VNB N_A_114_57#_M1011_g 0.00794326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_114_57#_c_1103_n 0.0327238f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_67 VNB N_A_114_57#_c_1104_n 0.0141373f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_68 VNB N_A_114_57#_c_1105_n 0.0334632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_114_57#_M1021_g 0.0397064f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_70 VNB N_A_114_57#_M1004_g 0.0451628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_114_57#_c_1108_n 0.0211809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_114_57#_c_1109_n 0.00606839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_114_57#_c_1110_n 0.0354215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_114_57#_c_1111_n 0.0114121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_114_57#_c_1112_n 0.0115074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1545_332#_M1005_g 0.0511432f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=2.725
cc_77 VNB N_A_1545_332#_M1027_g 0.00105714f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=2.255
cc_78 VNB N_A_1545_332#_c_1259_n 0.0579671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1545_332#_c_1260_n 0.01992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1545_332#_M1022_g 0.0182088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1545_332#_c_1262_n 0.00497842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1545_332#_c_1263_n 0.00390291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1545_332#_c_1264_n 2.81183e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1545_332#_c_1265_n 0.00812166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1545_332#_c_1266_n 0.00411923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1545_332#_c_1267_n 0.0311474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1545_332#_c_1268_n 0.0226398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1307_428#_M1029_g 0.0509833f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=2.725
cc_89 VNB N_A_1307_428#_c_1438_n 0.00747573f $X=-0.19 $Y=-0.245 $X2=0.38
+ $Y2=2.255
cc_90 VNB N_A_1307_428#_c_1439_n 0.00304526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1307_428#_c_1440_n 0.00164857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1307_428#_c_1441_n 0.0241465f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_93 VNB N_A_1307_428#_c_1442_n 0.00171028f $X=-0.19 $Y=-0.245 $X2=0.29
+ $Y2=1.07
cc_94 VNB N_A_1307_428#_c_1443_n 0.00491209f $X=-0.19 $Y=-0.245 $X2=0.29
+ $Y2=2.035
cc_95 VNB N_A_1307_428#_c_1444_n 0.00497605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1307_428#_c_1445_n 0.0296136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_RESET_B_M1025_g 0.00113044f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_98 VNB RESET_B 0.00697606f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.725
cc_99 VNB N_RESET_B_c_1560_n 0.0286972f $X=-0.19 $Y=-0.245 $X2=0.347 $Y2=0.88
cc_100 VNB N_RESET_B_c_1561_n 0.0208713f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.41
cc_101 VNB N_A_2317_367#_M1039_g 0.0309878f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=2.725
cc_102 VNB N_A_2317_367#_M1024_g 0.00114377f $X=-0.19 $Y=-0.245 $X2=0.29
+ $Y2=1.41
cc_103 VNB N_A_2317_367#_c_1592_n 0.00346631f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=2.255
cc_104 VNB N_A_2317_367#_c_1593_n 0.00356065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2317_367#_c_1594_n 5.67915e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2317_367#_c_1595_n 0.00356065f $X=-0.19 $Y=-0.245 $X2=0.29
+ $Y2=1.07
cc_107 VNB N_A_2317_367#_c_1596_n 0.0026183f $X=-0.19 $Y=-0.245 $X2=0.29
+ $Y2=1.07
cc_108 VNB N_A_2317_367#_c_1597_n 0.0097818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2317_367#_c_1598_n 0.0327828f $X=-0.19 $Y=-0.245 $X2=0.29
+ $Y2=1.295
cc_110 VNB N_VPWR_c_1651_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_531_47#_c_1793_n 0.00482125f $X=-0.19 $Y=-0.245 $X2=0.38
+ $Y2=2.255
cc_112 VNB N_A_531_47#_c_1794_n 0.00275587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_531_47#_c_1795_n 0.0100127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_Q_N_c_1865_n 0.0100281f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.725
cc_115 VNB N_Q_N_c_1866_n 0.00259606f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.41
cc_116 VNB N_Q_N_c_1867_n 0.00586888f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.255
cc_117 VNB N_Q_c_1901_n 0.0263603f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=2.255
cc_118 VNB N_Q_c_1902_n 0.0261045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB Q 0.0133613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1928_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1929_n 0.0259355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1930_n 0.00564356f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_123 VNB N_VGND_c_1931_n 0.00999718f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_124 VNB N_VGND_c_1932_n 0.00951844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1933_n 0.00674438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1934_n 0.0168508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1935_n 0.0117393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1936_n 0.0370513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1937_n 0.00632108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1938_n 0.0427133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1939_n 0.00478223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1940_n 0.0411239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1941_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1942_n 0.0546863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1943_n 0.0580007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1944_n 0.034456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1945_n 0.0190013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1946_n 0.660643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1947_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1948_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1949_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_A_917_47#_c_2075_n 0.00128814f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=2.725
cc_143 VNB N_A_917_47#_c_2076_n 0.00260912f $X=-0.19 $Y=-0.245 $X2=0.29
+ $Y2=1.575
cc_144 VNB N_A_1705_54#_c_2105_n 0.0196256f $X=-0.19 $Y=-0.245 $X2=0.347
+ $Y2=0.88
cc_145 VPB N_CLK_c_259_n 0.0344292f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=2.18
cc_146 VPB N_CLK_c_266_n 0.0218224f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.33
cc_147 VPB N_CLK_c_267_n 0.0389681f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.255
cc_148 VPB N_CLK_c_264_n 0.0221476f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_149 VPB N_D_c_300_n 0.0368901f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.88
cc_150 VPB N_D_c_301_n 0.0145975f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.725
cc_151 VPB D 0.00635081f $X=-0.19 $Y=1.655 $X2=0.347 $Y2=0.88
cc_152 VPB N_D_c_303_n 0.0446498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_225_47#_M1032_g 0.0368587f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.725
cc_154 VPB N_A_225_47#_M1007_g 0.0247098f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_155 VPB N_A_225_47#_c_360_n 0.0247742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_225_47#_c_361_n 0.0251508f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_157 VPB N_A_225_47#_c_362_n 0.00750216f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_158 VPB N_A_225_47#_c_375_n 0.00774175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_225_47#_c_376_n 0.00549286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_225_47#_c_377_n 0.00402215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_225_47#_c_378_n 0.00183635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_225_47#_c_364_n 0.0026483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_225_47#_c_380_n 0.0074129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_225_47#_c_381_n 0.0343615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_225_47#_c_369_n 0.00352882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_767_21#_M1009_g 0.0465823f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.41
cc_167 VPB N_A_767_21#_M1026_g 0.0223642f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.255
cc_168 VPB N_A_767_21#_c_556_n 0.00427013f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_169 VPB N_A_767_21#_c_557_n 7.19928e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_170 VPB N_A_767_21#_c_559_n 0.00408757f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_171 VPB N_A_767_21#_c_560_n 0.0119198f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_172 VPB N_A_767_21#_c_561_n 0.00231882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_767_21#_c_571_n 0.0042165f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_767_21#_c_562_n 0.00379487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_767_21#_c_563_n 0.00514433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_767_21#_c_574_n 0.00198183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_SET_B_c_715_n 0.03439f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.495
cc_178 VPB N_SET_B_M1010_g 0.0220795f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.575
cc_179 VPB N_SET_B_c_722_n 0.020858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_SET_B_c_723_n 7.53232e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_SET_B_c_724_n 7.85201e-19 $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_182 VPB N_SET_B_c_718_n 0.0184111f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.665
cc_183 VPB N_SET_B_c_719_n 0.00169882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_617_47#_M1015_g 0.0218333f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.41
cc_185 VPB N_A_617_47#_c_837_n 0.00940689f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_1091_21#_M1016_g 0.0197811f $X=-0.19 $Y=1.655 $X2=0.347 $Y2=1.03
cc_187 VPB N_A_1091_21#_M1001_g 0.0250327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_1091_21#_c_938_n 6.29763e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1091_21#_c_939_n 0.0178038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_1091_21#_c_945_n 0.00750098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_1091_21#_c_946_n 0.00950855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_114_57#_M1011_g 0.0474235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_114_57#_c_1114_n 0.140972f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_194 VPB N_A_114_57#_c_1115_n 0.012806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_114_57#_M1034_g 0.0388379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_114_57#_c_1117_n 0.20692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_114_57#_c_1118_n 0.0404248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_114_57#_M1017_g 0.00995358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_114_57#_c_1120_n 0.0472906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_114_57#_M1004_g 0.00120062f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_114_57#_c_1122_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_114_57#_c_1110_n 0.0313142f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_114_57#_c_1124_n 0.0156273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1545_332#_M1036_g 0.0512038f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.41
cc_205 VPB N_A_1545_332#_M1027_g 0.0263449f $X=-0.19 $Y=1.655 $X2=0.645
+ $Y2=2.255
cc_206 VPB N_A_1545_332#_M1022_g 0.0257447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_1545_332#_c_1272_n 0.00457671f $X=-0.19 $Y=1.655 $X2=0.29
+ $Y2=2.035
cc_208 VPB N_A_1545_332#_c_1273_n 0.034132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_1545_332#_c_1274_n 0.00342301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_1545_332#_c_1275_n 0.00344006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_1545_332#_c_1276_n 0.0019974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_1545_332#_c_1277_n 0.00650563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_1545_332#_c_1263_n 0.00170618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_1545_332#_c_1279_n 0.0248295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_1545_332#_c_1264_n 0.00174475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_1545_332#_c_1281_n 0.00164229f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_1307_428#_M1038_g 0.021883f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.41
cc_218 VPB N_A_1307_428#_c_1440_n 0.0142048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1307_428#_c_1448_n 0.00279081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_RESET_B_M1025_g 0.0278194f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.88
cc_221 VPB N_A_2317_367#_M1024_g 0.0281185f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.41
cc_222 VPB N_A_2317_367#_c_1600_n 0.00647927f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_223 VPB N_VPWR_c_1652_n 0.0144238f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_224 VPB N_VPWR_c_1653_n 0.0365901f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_225 VPB N_VPWR_c_1654_n 0.0139513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1655_n 0.0139329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1656_n 0.0111336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1657_n 0.00598237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1658_n 0.0250478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1659_n 0.0252991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1660_n 0.0190075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1661_n 0.0331037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1662_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1663_n 0.0284211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1664_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1665_n 0.0299474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1666_n 0.00590455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1667_n 0.063342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1668_n 0.0636406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1669_n 0.0236438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1670_n 0.0340313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1671_n 0.0190013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1651_n 0.149692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1673_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1674_n 0.00590455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1675_n 0.00601829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1676_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_531_47#_c_1796_n 0.00285974f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.41
cc_249 VPB N_A_531_47#_c_1795_n 0.0016501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_531_47#_c_1798_n 0.00690786f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_251 VPB N_Q_N_c_1868_n 0.00492403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_Q_N_c_1867_n 0.00304868f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.255
cc_253 VPB Q_N 0.0208894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_Q_c_1904_n 0.0427906f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.725
cc_255 VPB N_Q_c_1905_n 0.0133536f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.575
cc_256 VPB N_Q_c_1901_n 0.00776535f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=2.255
cc_257 N_CLK_c_267_n N_A_225_47#_c_362_n 2.11074e-19 $X=0.645 $Y=2.255 $X2=0
+ $Y2=0
cc_258 N_CLK_M1018_g N_A_225_47#_c_363_n 8.52124e-19 $X=0.495 $Y=0.495 $X2=0
+ $Y2=0
cc_259 N_CLK_c_267_n N_A_225_47#_c_378_n 7.17472e-19 $X=0.645 $Y=2.255 $X2=0
+ $Y2=0
cc_260 N_CLK_c_263_n N_A_114_57#_c_1109_n 0.00113859f $X=0.29 $Y=1.07 $X2=0
+ $Y2=0
cc_261 N_CLK_c_262_n N_A_114_57#_c_1110_n 0.0170166f $X=0.29 $Y=1.575 $X2=0
+ $Y2=0
cc_262 N_CLK_c_267_n N_A_114_57#_c_1110_n 0.00140388f $X=0.645 $Y=2.255 $X2=0
+ $Y2=0
cc_263 N_CLK_c_263_n N_A_114_57#_c_1110_n 0.0170166f $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_264 N_CLK_c_264_n N_A_114_57#_c_1110_n 0.00255104f $X=0.29 $Y=1.07 $X2=0
+ $Y2=0
cc_265 N_CLK_c_259_n N_A_114_57#_c_1124_n 0.00494999f $X=0.38 $Y=2.18 $X2=0
+ $Y2=0
cc_266 N_CLK_c_266_n N_A_114_57#_c_1124_n 0.0118143f $X=0.645 $Y=2.33 $X2=0
+ $Y2=0
cc_267 N_CLK_c_262_n N_A_114_57#_c_1124_n 0.00113859f $X=0.29 $Y=1.575 $X2=0
+ $Y2=0
cc_268 N_CLK_c_267_n N_A_114_57#_c_1124_n 0.0102281f $X=0.645 $Y=2.255 $X2=0
+ $Y2=0
cc_269 N_CLK_M1018_g N_A_114_57#_c_1111_n 0.00770576f $X=0.495 $Y=0.495 $X2=0
+ $Y2=0
cc_270 N_CLK_M1018_g N_A_114_57#_c_1112_n 0.00986148f $X=0.495 $Y=0.495 $X2=0
+ $Y2=0
cc_271 N_CLK_c_263_n N_A_114_57#_c_1112_n 0.00511962f $X=0.29 $Y=1.07 $X2=0
+ $Y2=0
cc_272 N_CLK_c_264_n N_A_114_57#_c_1112_n 0.0721364f $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_273 N_CLK_c_266_n N_VPWR_c_1653_n 0.0171119f $X=0.645 $Y=2.33 $X2=0 $Y2=0
cc_274 N_CLK_c_267_n N_VPWR_c_1653_n 0.0076598f $X=0.645 $Y=2.255 $X2=0 $Y2=0
cc_275 N_CLK_c_264_n N_VPWR_c_1653_n 0.0192751f $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_276 N_CLK_c_266_n N_VPWR_c_1661_n 0.00502664f $X=0.645 $Y=2.33 $X2=0 $Y2=0
cc_277 N_CLK_c_266_n N_VPWR_c_1651_n 0.011051f $X=0.645 $Y=2.33 $X2=0 $Y2=0
cc_278 N_CLK_M1018_g N_VGND_c_1929_n 0.00533583f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_279 N_CLK_c_261_n N_VGND_c_1929_n 0.00664962f $X=0.347 $Y=1.03 $X2=0 $Y2=0
cc_280 N_CLK_c_264_n N_VGND_c_1929_n 0.0203156f $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_281 N_CLK_M1018_g N_VGND_c_1936_n 0.00502664f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_282 N_CLK_M1018_g N_VGND_c_1946_n 0.0109766f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_283 N_CLK_c_261_n N_VGND_c_1946_n 0.00140006f $X=0.347 $Y=1.03 $X2=0 $Y2=0
cc_284 N_D_c_300_n N_A_225_47#_M1032_g 0.0180119f $X=2.685 $Y=2.165 $X2=0 $Y2=0
cc_285 N_D_c_300_n N_A_225_47#_c_360_n 0.0114375f $X=2.685 $Y=2.165 $X2=0 $Y2=0
cc_286 D N_A_225_47#_c_360_n 9.58754e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_287 N_D_c_303_n N_A_225_47#_c_360_n 0.00422899f $X=2.115 $Y=1.89 $X2=0 $Y2=0
cc_288 D N_A_225_47#_c_362_n 0.0994686f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_289 N_D_c_299_n N_A_225_47#_c_362_n 0.00195887f $X=1.935 $Y=0.84 $X2=0 $Y2=0
cc_290 N_D_c_303_n N_A_225_47#_c_362_n 0.0012251f $X=2.115 $Y=1.89 $X2=0 $Y2=0
cc_291 N_D_c_300_n N_A_225_47#_c_376_n 0.0131926f $X=2.685 $Y=2.165 $X2=0 $Y2=0
cc_292 N_D_c_301_n N_A_225_47#_c_376_n 0.00344592f $X=2.76 $Y=2.24 $X2=0 $Y2=0
cc_293 D N_A_225_47#_c_376_n 0.0391292f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_294 N_D_c_303_n N_A_225_47#_c_376_n 0.0060529f $X=2.115 $Y=1.89 $X2=0 $Y2=0
cc_295 N_D_c_300_n N_A_225_47#_c_377_n 0.0130624f $X=2.685 $Y=2.165 $X2=0 $Y2=0
cc_296 D N_A_225_47#_c_377_n 0.0130297f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_297 N_D_c_303_n N_A_225_47#_c_377_n 0.00508382f $X=2.115 $Y=1.89 $X2=0 $Y2=0
cc_298 N_D_c_300_n N_A_225_47#_c_364_n 0.00327696f $X=2.685 $Y=2.165 $X2=0 $Y2=0
cc_299 D N_A_225_47#_c_364_n 0.0267152f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_300 N_D_c_303_n N_A_225_47#_c_364_n 0.00126301f $X=2.115 $Y=1.89 $X2=0 $Y2=0
cc_301 D N_A_225_47#_c_366_n 0.00165575f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_302 N_D_c_296_n N_A_225_47#_c_367_n 0.00181458f $X=2.505 $Y=0.84 $X2=0 $Y2=0
cc_303 D N_A_225_47#_c_367_n 0.0281931f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_304 D N_A_114_57#_M1008_g 0.00211913f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_305 N_D_c_299_n N_A_114_57#_M1008_g 0.0211581f $X=1.935 $Y=0.84 $X2=0 $Y2=0
cc_306 D N_A_114_57#_M1011_g 0.00589074f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_307 N_D_c_303_n N_A_114_57#_M1011_g 0.0222844f $X=2.115 $Y=1.89 $X2=0 $Y2=0
cc_308 N_D_c_296_n N_A_114_57#_c_1103_n 0.0056548f $X=2.505 $Y=0.84 $X2=0 $Y2=0
cc_309 N_D_c_300_n N_A_114_57#_c_1103_n 0.0047146f $X=2.685 $Y=2.165 $X2=0 $Y2=0
cc_310 D N_A_114_57#_c_1103_n 0.0245662f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_311 N_D_c_299_n N_A_114_57#_c_1103_n 0.0180853f $X=1.935 $Y=0.84 $X2=0 $Y2=0
cc_312 N_D_c_303_n N_A_114_57#_c_1103_n 0.0181064f $X=2.115 $Y=1.89 $X2=0 $Y2=0
cc_313 N_D_c_301_n N_A_114_57#_c_1114_n 0.0103003f $X=2.76 $Y=2.24 $X2=0 $Y2=0
cc_314 N_D_c_297_n N_A_114_57#_M1021_g 0.0202573f $X=2.58 $Y=0.765 $X2=0 $Y2=0
cc_315 D N_A_114_57#_M1021_g 0.00410768f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_316 N_D_c_296_n N_A_114_57#_c_1108_n 0.0202029f $X=2.505 $Y=0.84 $X2=0 $Y2=0
cc_317 D N_A_114_57#_c_1108_n 0.00608116f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_318 N_D_c_301_n N_VPWR_c_1654_n 0.00671345f $X=2.76 $Y=2.24 $X2=0 $Y2=0
cc_319 N_D_c_301_n N_VPWR_c_1651_n 9.39239e-19 $X=2.76 $Y=2.24 $X2=0 $Y2=0
cc_320 N_D_c_296_n N_A_531_47#_c_1799_n 0.0022486f $X=2.505 $Y=0.84 $X2=0 $Y2=0
cc_321 N_D_c_297_n N_A_531_47#_c_1799_n 0.0156311f $X=2.58 $Y=0.765 $X2=0 $Y2=0
cc_322 D N_A_531_47#_c_1799_n 0.00280632f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_323 N_D_c_300_n N_A_531_47#_c_1796_n 3.3619e-19 $X=2.685 $Y=2.165 $X2=0 $Y2=0
cc_324 N_D_c_301_n N_A_531_47#_c_1796_n 0.0187162f $X=2.76 $Y=2.24 $X2=0 $Y2=0
cc_325 N_D_c_296_n N_A_531_47#_c_1794_n 0.0031719f $X=2.505 $Y=0.84 $X2=0 $Y2=0
cc_326 D N_A_531_47#_c_1794_n 0.00865372f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_327 N_D_c_299_n N_A_531_47#_c_1794_n 4.45107e-19 $X=1.935 $Y=0.84 $X2=0 $Y2=0
cc_328 N_D_c_300_n N_A_531_47#_c_1798_n 0.00423644f $X=2.685 $Y=2.165 $X2=0
+ $Y2=0
cc_329 N_D_c_297_n N_VGND_c_1930_n 0.0088163f $X=2.58 $Y=0.765 $X2=0 $Y2=0
cc_330 D N_VGND_c_1930_n 0.0259955f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_331 N_D_c_299_n N_VGND_c_1930_n 0.00252096f $X=1.935 $Y=0.84 $X2=0 $Y2=0
cc_332 N_D_c_296_n N_VGND_c_1942_n 0.00350456f $X=2.505 $Y=0.84 $X2=0 $Y2=0
cc_333 N_D_c_297_n N_VGND_c_1942_n 0.00549284f $X=2.58 $Y=0.765 $X2=0 $Y2=0
cc_334 N_D_c_299_n N_VGND_c_1942_n 0.00133406f $X=1.935 $Y=0.84 $X2=0 $Y2=0
cc_335 N_D_c_297_n N_VGND_c_1946_n 0.0115186f $X=2.58 $Y=0.765 $X2=0 $Y2=0
cc_336 D N_VGND_c_1946_n 0.0082716f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_337 N_D_c_299_n N_VGND_c_1946_n 0.00481363f $X=1.935 $Y=0.84 $X2=0 $Y2=0
cc_338 N_A_225_47#_M1031_g N_A_767_21#_M1028_g 0.0424617f $X=3.52 $Y=0.445 $X2=0
+ $Y2=0
cc_339 N_A_225_47#_c_365_n N_A_767_21#_M1028_g 0.00664788f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_340 N_A_225_47#_c_361_n N_A_767_21#_M1009_g 0.00373941f $X=3.52 $Y=1.715
+ $X2=0 $Y2=0
cc_341 N_A_225_47#_c_365_n N_A_767_21#_c_557_n 0.00614479f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_342 N_A_225_47#_M1013_g N_A_767_21#_M1012_g 0.051395f $X=6.91 $Y=0.59 $X2=0
+ $Y2=0
cc_343 N_A_225_47#_M1031_g N_A_767_21#_c_559_n 3.20736e-19 $X=3.52 $Y=0.445
+ $X2=0 $Y2=0
cc_344 N_A_225_47#_c_361_n N_A_767_21#_c_559_n 4.30772e-19 $X=3.52 $Y=1.715
+ $X2=0 $Y2=0
cc_345 N_A_225_47#_c_365_n N_A_767_21#_c_559_n 0.00813614f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_346 N_A_225_47#_c_361_n N_A_767_21#_c_560_n 0.0424617f $X=3.52 $Y=1.715 $X2=0
+ $Y2=0
cc_347 N_A_225_47#_c_365_n N_A_767_21#_c_584_n 0.00348578f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_348 N_A_225_47#_c_365_n N_A_767_21#_c_585_n 0.00770185f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_349 N_A_225_47#_c_365_n N_A_767_21#_c_586_n 0.00572941f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_350 N_A_225_47#_c_365_n N_A_767_21#_c_561_n 0.0234933f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_351 N_A_225_47#_c_365_n N_A_767_21#_c_571_n 0.0167243f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_352 N_A_225_47#_c_369_n N_A_767_21#_c_571_n 0.00863979f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_353 N_A_225_47#_c_365_n N_A_767_21#_c_562_n 0.0267614f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_354 N_A_225_47#_c_422_p N_A_767_21#_c_562_n 6.18576e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_355 N_A_225_47#_c_368_n N_A_767_21#_c_562_n 0.00107576f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_356 N_A_225_47#_c_369_n N_A_767_21#_c_562_n 0.0479339f $X=6.97 $Y=1.275 $X2=0
+ $Y2=0
cc_357 N_A_225_47#_c_365_n N_A_767_21#_c_563_n 0.00281319f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_358 N_A_225_47#_c_368_n N_A_767_21#_c_563_n 0.0217086f $X=6.97 $Y=1.275 $X2=0
+ $Y2=0
cc_359 N_A_225_47#_c_369_n N_A_767_21#_c_563_n 0.00234154f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_360 N_A_225_47#_c_365_n N_SET_B_M1003_g 0.00545234f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_361 N_A_225_47#_c_365_n N_SET_B_c_715_n 0.00255946f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_362 N_A_225_47#_c_380_n N_SET_B_c_722_n 0.0111487f $X=7.11 $Y=2.235 $X2=0
+ $Y2=0
cc_363 N_A_225_47#_c_381_n N_SET_B_c_722_n 8.97701e-19 $X=7.11 $Y=2.235 $X2=0
+ $Y2=0
cc_364 N_A_225_47#_c_422_p N_SET_B_c_722_n 0.0110708f $X=6.96 $Y=1.295 $X2=0
+ $Y2=0
cc_365 N_A_225_47#_c_369_n N_SET_B_c_722_n 0.0159225f $X=6.97 $Y=1.275 $X2=0
+ $Y2=0
cc_366 N_A_225_47#_c_365_n N_SET_B_c_733_n 0.012286f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_367 N_A_225_47#_c_365_n N_SET_B_c_717_n 0.00517532f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_368 N_A_225_47#_c_365_n N_A_617_47#_c_834_n 0.00282295f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_369 N_A_225_47#_M1031_g N_A_617_47#_c_836_n 0.0088702f $X=3.52 $Y=0.445 $X2=0
+ $Y2=0
cc_370 N_A_225_47#_M1032_g N_A_617_47#_c_837_n 0.00504683f $X=3.19 $Y=2.525
+ $X2=0 $Y2=0
cc_371 N_A_225_47#_M1031_g N_A_617_47#_c_837_n 0.00554466f $X=3.52 $Y=0.445
+ $X2=0 $Y2=0
cc_372 N_A_225_47#_c_361_n N_A_617_47#_c_837_n 0.015799f $X=3.52 $Y=1.715 $X2=0
+ $Y2=0
cc_373 N_A_225_47#_c_365_n N_A_617_47#_c_837_n 0.0176827f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_374 N_A_225_47#_c_365_n N_A_617_47#_c_838_n 0.0732074f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_375 N_A_225_47#_M1031_g N_A_617_47#_c_848_n 0.0116458f $X=3.52 $Y=0.445 $X2=0
+ $Y2=0
cc_376 N_A_225_47#_c_365_n N_A_617_47#_c_848_n 0.00604375f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_377 N_A_225_47#_M1031_g N_A_617_47#_c_850_n 0.00399103f $X=3.52 $Y=0.445
+ $X2=0 $Y2=0
cc_378 N_A_225_47#_c_365_n N_A_617_47#_c_850_n 0.00908224f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_379 N_A_225_47#_c_365_n N_A_1091_21#_M1016_g 0.00156241f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_380 N_A_225_47#_c_365_n N_A_1091_21#_c_927_n 0.0218603f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_381 N_A_225_47#_c_365_n N_A_1091_21#_c_928_n 0.00987012f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_382 N_A_225_47#_M1013_g N_A_1091_21#_c_929_n 0.00135798f $X=6.91 $Y=0.59
+ $X2=0 $Y2=0
cc_383 N_A_225_47#_c_365_n N_A_1091_21#_c_929_n 0.018502f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_384 N_A_225_47#_M1013_g N_A_1091_21#_c_952_n 0.00494431f $X=6.91 $Y=0.59
+ $X2=0 $Y2=0
cc_385 N_A_225_47#_M1013_g N_A_1091_21#_c_931_n 0.0125081f $X=6.91 $Y=0.59 $X2=0
+ $Y2=0
cc_386 N_A_225_47#_c_369_n N_A_1091_21#_c_931_n 0.00337848f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_387 N_A_225_47#_c_362_n N_A_114_57#_c_1100_n 0.0120137f $X=1.42 $Y=2.235
+ $X2=0 $Y2=0
cc_388 N_A_225_47#_c_363_n N_A_114_57#_c_1100_n 0.00347188f $X=1.27 $Y=0.47
+ $X2=0 $Y2=0
cc_389 N_A_225_47#_c_362_n N_A_114_57#_M1008_g 0.0256296f $X=1.42 $Y=2.235 $X2=0
+ $Y2=0
cc_390 N_A_225_47#_c_363_n N_A_114_57#_M1008_g 0.0135811f $X=1.27 $Y=0.47 $X2=0
+ $Y2=0
cc_391 N_A_225_47#_c_362_n N_A_114_57#_M1011_g 0.0230791f $X=1.42 $Y=2.235 $X2=0
+ $Y2=0
cc_392 N_A_225_47#_c_375_n N_A_114_57#_M1011_g 0.0127087f $X=1.42 $Y=2.46 $X2=0
+ $Y2=0
cc_393 N_A_225_47#_c_376_n N_A_114_57#_M1011_g 0.0168813f $X=2.46 $Y=2.32 $X2=0
+ $Y2=0
cc_394 N_A_225_47#_c_378_n N_A_114_57#_M1011_g 0.0019878f $X=1.42 $Y=2.32 $X2=0
+ $Y2=0
cc_395 N_A_225_47#_c_362_n N_A_114_57#_c_1104_n 0.00677719f $X=1.42 $Y=2.235
+ $X2=0 $Y2=0
cc_396 N_A_225_47#_M1032_g N_A_114_57#_c_1114_n 0.0103003f $X=3.19 $Y=2.525
+ $X2=0 $Y2=0
cc_397 N_A_225_47#_c_376_n N_A_114_57#_c_1114_n 0.0122483f $X=2.46 $Y=2.32 $X2=0
+ $Y2=0
cc_398 N_A_225_47#_c_360_n N_A_114_57#_c_1105_n 0.023749f $X=3.115 $Y=1.715
+ $X2=0 $Y2=0
cc_399 N_A_225_47#_c_364_n N_A_114_57#_c_1105_n 0.00166488f $X=2.835 $Y=1.715
+ $X2=0 $Y2=0
cc_400 N_A_225_47#_c_365_n N_A_114_57#_c_1105_n 0.00415482f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_401 N_A_225_47#_c_366_n N_A_114_57#_c_1105_n 0.00397741f $X=2.785 $Y=1.295
+ $X2=0 $Y2=0
cc_402 N_A_225_47#_c_367_n N_A_114_57#_c_1105_n 0.0142624f $X=2.64 $Y=1.295
+ $X2=0 $Y2=0
cc_403 N_A_225_47#_M1031_g N_A_114_57#_M1021_g 0.0296078f $X=3.52 $Y=0.445 $X2=0
+ $Y2=0
cc_404 N_A_225_47#_M1032_g N_A_114_57#_M1034_g 0.0152735f $X=3.19 $Y=2.525 $X2=0
+ $Y2=0
cc_405 N_A_225_47#_M1007_g N_A_114_57#_c_1117_n 0.0116078f $X=7.02 $Y=2.77 $X2=0
+ $Y2=0
cc_406 N_A_225_47#_c_365_n N_A_114_57#_c_1118_n 0.00473279f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_407 N_A_225_47#_c_369_n N_A_114_57#_c_1118_n 0.00547227f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_408 N_A_225_47#_c_380_n N_A_114_57#_M1017_g 0.00624953f $X=7.11 $Y=2.235
+ $X2=0 $Y2=0
cc_409 N_A_225_47#_c_381_n N_A_114_57#_M1017_g 0.0116078f $X=7.11 $Y=2.235 $X2=0
+ $Y2=0
cc_410 N_A_225_47#_c_369_n N_A_114_57#_M1017_g 2.33135e-19 $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_411 N_A_225_47#_c_380_n N_A_114_57#_c_1120_n 0.0010972f $X=7.11 $Y=2.235
+ $X2=0 $Y2=0
cc_412 N_A_225_47#_c_381_n N_A_114_57#_c_1120_n 0.0178119f $X=7.11 $Y=2.235
+ $X2=0 $Y2=0
cc_413 N_A_225_47#_c_368_n N_A_114_57#_c_1120_n 0.0181215f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_414 N_A_225_47#_c_369_n N_A_114_57#_c_1120_n 0.0176575f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_415 N_A_225_47#_M1013_g N_A_114_57#_M1004_g 0.0177094f $X=6.91 $Y=0.59 $X2=0
+ $Y2=0
cc_416 N_A_225_47#_c_368_n N_A_114_57#_M1004_g 0.0205681f $X=6.97 $Y=1.275 $X2=0
+ $Y2=0
cc_417 N_A_225_47#_c_369_n N_A_114_57#_M1004_g 0.00463403f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_418 N_A_225_47#_c_367_n N_A_114_57#_c_1108_n 0.00565087f $X=2.64 $Y=1.295
+ $X2=0 $Y2=0
cc_419 N_A_225_47#_c_362_n N_A_114_57#_c_1109_n 0.0614794f $X=1.42 $Y=2.235
+ $X2=0 $Y2=0
cc_420 N_A_225_47#_c_362_n N_A_114_57#_c_1110_n 0.00468928f $X=1.42 $Y=2.235
+ $X2=0 $Y2=0
cc_421 N_A_225_47#_c_375_n N_A_114_57#_c_1124_n 0.0383948f $X=1.42 $Y=2.46 $X2=0
+ $Y2=0
cc_422 N_A_225_47#_c_378_n N_A_114_57#_c_1124_n 0.0121616f $X=1.42 $Y=2.32 $X2=0
+ $Y2=0
cc_423 N_A_225_47#_c_362_n N_A_114_57#_c_1111_n 0.027207f $X=1.42 $Y=2.235 $X2=0
+ $Y2=0
cc_424 N_A_225_47#_c_363_n N_A_114_57#_c_1111_n 0.0284467f $X=1.27 $Y=0.47 $X2=0
+ $Y2=0
cc_425 N_A_225_47#_M1007_g N_A_1545_332#_M1036_g 0.0120961f $X=7.02 $Y=2.77
+ $X2=0 $Y2=0
cc_426 N_A_225_47#_c_381_n N_A_1545_332#_M1036_g 0.0063142f $X=7.11 $Y=2.235
+ $X2=0 $Y2=0
cc_427 N_A_225_47#_M1013_g N_A_1307_428#_c_1438_n 0.00445671f $X=6.91 $Y=0.59
+ $X2=0 $Y2=0
cc_428 N_A_225_47#_c_422_p N_A_1307_428#_c_1438_n 9.5169e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_429 N_A_225_47#_c_368_n N_A_1307_428#_c_1438_n 0.00108863f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_430 N_A_225_47#_c_369_n N_A_1307_428#_c_1438_n 0.0128505f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_431 N_A_225_47#_M1007_g N_A_1307_428#_c_1453_n 0.00984282f $X=7.02 $Y=2.77
+ $X2=0 $Y2=0
cc_432 N_A_225_47#_c_380_n N_A_1307_428#_c_1453_n 0.0165257f $X=7.11 $Y=2.235
+ $X2=0 $Y2=0
cc_433 N_A_225_47#_c_381_n N_A_1307_428#_c_1453_n 0.00236287f $X=7.11 $Y=2.235
+ $X2=0 $Y2=0
cc_434 N_A_225_47#_M1013_g N_A_1307_428#_c_1439_n 0.00317119f $X=6.91 $Y=0.59
+ $X2=0 $Y2=0
cc_435 N_A_225_47#_c_422_p N_A_1307_428#_c_1439_n 8.76507e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_436 N_A_225_47#_c_368_n N_A_1307_428#_c_1439_n 0.00105498f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_437 N_A_225_47#_c_369_n N_A_1307_428#_c_1439_n 0.0134695f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_438 N_A_225_47#_M1007_g N_A_1307_428#_c_1440_n 0.00356074f $X=7.02 $Y=2.77
+ $X2=0 $Y2=0
cc_439 N_A_225_47#_c_380_n N_A_1307_428#_c_1440_n 0.0239123f $X=7.11 $Y=2.235
+ $X2=0 $Y2=0
cc_440 N_A_225_47#_c_381_n N_A_1307_428#_c_1440_n 0.00288152f $X=7.11 $Y=2.235
+ $X2=0 $Y2=0
cc_441 N_A_225_47#_c_369_n N_A_1307_428#_c_1440_n 0.0297083f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_442 N_A_225_47#_M1007_g N_A_1307_428#_c_1448_n 0.0127968f $X=7.02 $Y=2.77
+ $X2=0 $Y2=0
cc_443 N_A_225_47#_c_380_n N_A_1307_428#_c_1448_n 0.011054f $X=7.11 $Y=2.235
+ $X2=0 $Y2=0
cc_444 N_A_225_47#_c_422_p N_A_1307_428#_c_1443_n 7.6822e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_445 N_A_225_47#_c_368_n N_A_1307_428#_c_1443_n 8.02731e-19 $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_446 N_A_225_47#_c_369_n N_A_1307_428#_c_1443_n 0.0130481f $X=6.97 $Y=1.275
+ $X2=0 $Y2=0
cc_447 N_A_225_47#_c_376_n N_VPWR_M1011_d 0.0134815f $X=2.46 $Y=2.32 $X2=0 $Y2=0
cc_448 N_A_225_47#_c_375_n N_VPWR_c_1654_n 0.0147373f $X=1.42 $Y=2.46 $X2=0
+ $Y2=0
cc_449 N_A_225_47#_c_376_n N_VPWR_c_1654_n 0.0254908f $X=2.46 $Y=2.32 $X2=0
+ $Y2=0
cc_450 N_A_225_47#_c_375_n N_VPWR_c_1661_n 0.0142766f $X=1.42 $Y=2.46 $X2=0
+ $Y2=0
cc_451 N_A_225_47#_M1007_g N_VPWR_c_1668_n 0.0032848f $X=7.02 $Y=2.77 $X2=0
+ $Y2=0
cc_452 N_A_225_47#_M1032_g N_VPWR_c_1651_n 9.39239e-19 $X=3.19 $Y=2.525 $X2=0
+ $Y2=0
cc_453 N_A_225_47#_M1007_g N_VPWR_c_1651_n 0.004474f $X=7.02 $Y=2.77 $X2=0 $Y2=0
cc_454 N_A_225_47#_c_375_n N_VPWR_c_1651_n 0.0119616f $X=1.42 $Y=2.46 $X2=0
+ $Y2=0
cc_455 N_A_225_47#_M1031_g N_A_531_47#_c_1799_n 5.44874e-19 $X=3.52 $Y=0.445
+ $X2=0 $Y2=0
cc_456 N_A_225_47#_M1032_g N_A_531_47#_c_1796_n 0.00829939f $X=3.19 $Y=2.525
+ $X2=0 $Y2=0
cc_457 N_A_225_47#_c_376_n N_A_531_47#_c_1796_n 0.00959795f $X=2.46 $Y=2.32
+ $X2=0 $Y2=0
cc_458 N_A_225_47#_c_377_n N_A_531_47#_c_1796_n 3.08694e-19 $X=2.545 $Y=2.235
+ $X2=0 $Y2=0
cc_459 N_A_225_47#_M1031_g N_A_531_47#_c_1793_n 0.00145813f $X=3.52 $Y=0.445
+ $X2=0 $Y2=0
cc_460 N_A_225_47#_c_360_n N_A_531_47#_c_1793_n 0.00297439f $X=3.115 $Y=1.715
+ $X2=0 $Y2=0
cc_461 N_A_225_47#_c_364_n N_A_531_47#_c_1793_n 4.37441e-19 $X=2.835 $Y=1.715
+ $X2=0 $Y2=0
cc_462 N_A_225_47#_c_365_n N_A_531_47#_c_1793_n 0.00803236f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_463 N_A_225_47#_c_364_n N_A_531_47#_c_1794_n 0.00286266f $X=2.835 $Y=1.715
+ $X2=0 $Y2=0
cc_464 N_A_225_47#_c_365_n N_A_531_47#_c_1794_n 0.0047119f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_465 N_A_225_47#_c_366_n N_A_531_47#_c_1794_n 0.00202377f $X=2.785 $Y=1.295
+ $X2=0 $Y2=0
cc_466 N_A_225_47#_c_367_n N_A_531_47#_c_1794_n 0.00830591f $X=2.64 $Y=1.295
+ $X2=0 $Y2=0
cc_467 N_A_225_47#_M1032_g N_A_531_47#_c_1795_n 0.00741878f $X=3.19 $Y=2.525
+ $X2=0 $Y2=0
cc_468 N_A_225_47#_M1031_g N_A_531_47#_c_1795_n 0.00711489f $X=3.52 $Y=0.445
+ $X2=0 $Y2=0
cc_469 N_A_225_47#_c_361_n N_A_531_47#_c_1795_n 0.0200733f $X=3.52 $Y=1.715
+ $X2=0 $Y2=0
cc_470 N_A_225_47#_c_377_n N_A_531_47#_c_1795_n 0.00531167f $X=2.545 $Y=2.235
+ $X2=0 $Y2=0
cc_471 N_A_225_47#_c_364_n N_A_531_47#_c_1795_n 0.0226912f $X=2.835 $Y=1.715
+ $X2=0 $Y2=0
cc_472 N_A_225_47#_c_365_n N_A_531_47#_c_1795_n 0.0145154f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_473 N_A_225_47#_c_366_n N_A_531_47#_c_1795_n 0.00209117f $X=2.785 $Y=1.295
+ $X2=0 $Y2=0
cc_474 N_A_225_47#_c_367_n N_A_531_47#_c_1795_n 0.011938f $X=2.64 $Y=1.295 $X2=0
+ $Y2=0
cc_475 N_A_225_47#_M1032_g N_A_531_47#_c_1798_n 0.0154202f $X=3.19 $Y=2.525
+ $X2=0 $Y2=0
cc_476 N_A_225_47#_c_360_n N_A_531_47#_c_1798_n 0.00806151f $X=3.115 $Y=1.715
+ $X2=0 $Y2=0
cc_477 N_A_225_47#_c_361_n N_A_531_47#_c_1798_n 3.96493e-19 $X=3.52 $Y=1.715
+ $X2=0 $Y2=0
cc_478 N_A_225_47#_c_377_n N_A_531_47#_c_1798_n 0.0122262f $X=2.545 $Y=2.235
+ $X2=0 $Y2=0
cc_479 N_A_225_47#_c_364_n N_A_531_47#_c_1798_n 0.0136458f $X=2.835 $Y=1.715
+ $X2=0 $Y2=0
cc_480 N_A_225_47#_c_363_n N_VGND_c_1936_n 0.0282984f $X=1.27 $Y=0.47 $X2=0
+ $Y2=0
cc_481 N_A_225_47#_M1013_g N_VGND_c_1940_n 0.00337062f $X=6.91 $Y=0.59 $X2=0
+ $Y2=0
cc_482 N_A_225_47#_M1031_g N_VGND_c_1942_n 0.00393552f $X=3.52 $Y=0.445 $X2=0
+ $Y2=0
cc_483 N_A_225_47#_M1008_s N_VGND_c_1946_n 0.00232985f $X=1.125 $Y=0.235 $X2=0
+ $Y2=0
cc_484 N_A_225_47#_M1031_g N_VGND_c_1946_n 0.00577637f $X=3.52 $Y=0.445 $X2=0
+ $Y2=0
cc_485 N_A_225_47#_M1013_g N_VGND_c_1946_n 0.00602632f $X=6.91 $Y=0.59 $X2=0
+ $Y2=0
cc_486 N_A_225_47#_c_363_n N_VGND_c_1946_n 0.0177283f $X=1.27 $Y=0.47 $X2=0
+ $Y2=0
cc_487 N_A_767_21#_M1028_g N_SET_B_M1003_g 0.0299917f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_488 N_A_767_21#_M1009_g N_SET_B_c_715_n 0.0215931f $X=4.09 $Y=2.525 $X2=0
+ $Y2=0
cc_489 N_A_767_21#_c_559_n N_SET_B_c_715_n 0.00262119f $X=4 $Y=1.57 $X2=0 $Y2=0
cc_490 N_A_767_21#_c_560_n N_SET_B_c_715_n 0.0225622f $X=4 $Y=1.57 $X2=0 $Y2=0
cc_491 N_A_767_21#_c_601_p N_SET_B_c_715_n 0.0104299f $X=4.855 $Y=2.415 $X2=0
+ $Y2=0
cc_492 N_A_767_21#_M1030_d N_SET_B_c_722_n 0.00246114f $X=4.8 $Y=1.895 $X2=0
+ $Y2=0
cc_493 N_A_767_21#_c_601_p N_SET_B_c_722_n 0.00565077f $X=4.855 $Y=2.415 $X2=0
+ $Y2=0
cc_494 N_A_767_21#_c_584_n N_SET_B_c_722_n 0.0244889f $X=4.98 $Y=2.13 $X2=0
+ $Y2=0
cc_495 N_A_767_21#_c_586_n N_SET_B_c_722_n 0.0246749f $X=5.38 $Y=2.045 $X2=0
+ $Y2=0
cc_496 N_A_767_21#_c_571_n N_SET_B_c_722_n 0.0838384f $X=6.225 $Y=2.045 $X2=0
+ $Y2=0
cc_497 N_A_767_21#_c_563_n N_SET_B_c_722_n 2.27217e-19 $X=6.39 $Y=1.275 $X2=0
+ $Y2=0
cc_498 N_A_767_21#_c_608_p N_SET_B_c_722_n 0.0189773f $X=5.465 $Y=2.045 $X2=0
+ $Y2=0
cc_499 N_A_767_21#_c_559_n N_SET_B_c_733_n 0.00145194f $X=4 $Y=1.57 $X2=0 $Y2=0
cc_500 N_A_767_21#_c_601_p N_SET_B_c_733_n 0.00281995f $X=4.855 $Y=2.415 $X2=0
+ $Y2=0
cc_501 N_A_767_21#_c_584_n N_SET_B_c_733_n 7.96392e-19 $X=4.98 $Y=2.13 $X2=0
+ $Y2=0
cc_502 N_A_767_21#_c_612_p N_SET_B_c_733_n 5.12238e-19 $X=4.98 $Y=2.33 $X2=0
+ $Y2=0
cc_503 N_A_767_21#_c_601_p N_SET_B_c_723_n 0.0163278f $X=4.855 $Y=2.415 $X2=0
+ $Y2=0
cc_504 N_A_767_21#_c_584_n N_SET_B_c_723_n 0.0076826f $X=4.98 $Y=2.13 $X2=0
+ $Y2=0
cc_505 N_A_767_21#_M1009_g N_SET_B_c_717_n 0.0029146f $X=4.09 $Y=2.525 $X2=0
+ $Y2=0
cc_506 N_A_767_21#_c_559_n N_SET_B_c_717_n 0.046019f $X=4 $Y=1.57 $X2=0 $Y2=0
cc_507 N_A_767_21#_c_560_n N_SET_B_c_717_n 0.00126755f $X=4 $Y=1.57 $X2=0 $Y2=0
cc_508 N_A_767_21#_c_601_p N_SET_B_c_717_n 3.20975e-19 $X=4.855 $Y=2.415 $X2=0
+ $Y2=0
cc_509 N_A_767_21#_c_561_n N_SET_B_c_717_n 0.00970892f $X=5.465 $Y=1.96 $X2=0
+ $Y2=0
cc_510 N_A_767_21#_c_561_n N_A_617_47#_M1023_g 0.0024409f $X=5.465 $Y=1.96 $X2=0
+ $Y2=0
cc_511 N_A_767_21#_c_584_n N_A_617_47#_c_834_n 7.95803e-19 $X=4.98 $Y=2.13 $X2=0
+ $Y2=0
cc_512 N_A_767_21#_c_585_n N_A_617_47#_c_834_n 0.00553179f $X=5.38 $Y=0.745
+ $X2=0 $Y2=0
cc_513 N_A_767_21#_c_561_n N_A_617_47#_c_834_n 0.00260671f $X=5.465 $Y=1.96
+ $X2=0 $Y2=0
cc_514 N_A_767_21#_c_584_n N_A_617_47#_M1015_g 0.00105405f $X=4.98 $Y=2.13 $X2=0
+ $Y2=0
cc_515 N_A_767_21#_c_612_p N_A_617_47#_M1015_g 0.003477f $X=4.98 $Y=2.33 $X2=0
+ $Y2=0
cc_516 N_A_767_21#_c_586_n N_A_617_47#_M1015_g 0.012339f $X=5.38 $Y=2.045 $X2=0
+ $Y2=0
cc_517 N_A_767_21#_c_561_n N_A_617_47#_M1015_g 0.00804604f $X=5.465 $Y=1.96
+ $X2=0 $Y2=0
cc_518 N_A_767_21#_c_574_n N_A_617_47#_M1015_g 0.00812069f $X=4.98 $Y=2.415
+ $X2=0 $Y2=0
cc_519 N_A_767_21#_M1028_g N_A_617_47#_c_836_n 0.00549101f $X=3.91 $Y=0.445
+ $X2=0 $Y2=0
cc_520 N_A_767_21#_M1028_g N_A_617_47#_c_837_n 0.00526429f $X=3.91 $Y=0.445
+ $X2=0 $Y2=0
cc_521 N_A_767_21#_M1009_g N_A_617_47#_c_837_n 0.00344136f $X=4.09 $Y=2.525
+ $X2=0 $Y2=0
cc_522 N_A_767_21#_c_559_n N_A_617_47#_c_837_n 0.0676646f $X=4 $Y=1.57 $X2=0
+ $Y2=0
cc_523 N_A_767_21#_c_633_p N_A_617_47#_c_837_n 0.0131757f $X=4.165 $Y=2.415
+ $X2=0 $Y2=0
cc_524 N_A_767_21#_M1028_g N_A_617_47#_c_838_n 0.0154915f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_525 N_A_767_21#_c_559_n N_A_617_47#_c_838_n 0.0161137f $X=4 $Y=1.57 $X2=0
+ $Y2=0
cc_526 N_A_767_21#_c_560_n N_A_617_47#_c_838_n 0.00123268f $X=4 $Y=1.57 $X2=0
+ $Y2=0
cc_527 N_A_767_21#_c_584_n N_A_617_47#_c_838_n 0.00288911f $X=4.98 $Y=2.13 $X2=0
+ $Y2=0
cc_528 N_A_767_21#_c_585_n N_A_617_47#_c_838_n 0.00875788f $X=5.38 $Y=0.745
+ $X2=0 $Y2=0
cc_529 N_A_767_21#_c_586_n N_A_617_47#_c_838_n 0.00144162f $X=5.38 $Y=2.045
+ $X2=0 $Y2=0
cc_530 N_A_767_21#_c_561_n N_A_617_47#_c_838_n 0.0224711f $X=5.465 $Y=1.96 $X2=0
+ $Y2=0
cc_531 N_A_767_21#_M1028_g N_A_617_47#_c_848_n 0.0021704f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_532 N_A_767_21#_c_585_n N_A_1091_21#_c_922_n 0.00884894f $X=5.38 $Y=0.745
+ $X2=0 $Y2=0
cc_533 N_A_767_21#_c_561_n N_A_1091_21#_c_922_n 0.00260986f $X=5.465 $Y=1.96
+ $X2=0 $Y2=0
cc_534 N_A_767_21#_c_557_n N_A_1091_21#_M1016_g 0.0411592f $X=6.06 $Y=1.6 $X2=0
+ $Y2=0
cc_535 N_A_767_21#_c_612_p N_A_1091_21#_M1016_g 0.00215432f $X=4.98 $Y=2.33
+ $X2=0 $Y2=0
cc_536 N_A_767_21#_c_561_n N_A_1091_21#_M1016_g 0.0181806f $X=5.465 $Y=1.96
+ $X2=0 $Y2=0
cc_537 N_A_767_21#_c_571_n N_A_1091_21#_M1016_g 0.00709788f $X=6.225 $Y=2.045
+ $X2=0 $Y2=0
cc_538 N_A_767_21#_c_562_n N_A_1091_21#_M1016_g 0.00106779f $X=6.39 $Y=1.275
+ $X2=0 $Y2=0
cc_539 N_A_767_21#_c_563_n N_A_1091_21#_M1016_g 0.00350914f $X=6.39 $Y=1.275
+ $X2=0 $Y2=0
cc_540 N_A_767_21#_c_608_p N_A_1091_21#_M1016_g 0.00711245f $X=5.465 $Y=2.045
+ $X2=0 $Y2=0
cc_541 N_A_767_21#_c_557_n N_A_1091_21#_c_927_n 7.36814e-19 $X=6.06 $Y=1.6 $X2=0
+ $Y2=0
cc_542 N_A_767_21#_M1012_g N_A_1091_21#_c_927_n 0.00220886f $X=6.52 $Y=0.59
+ $X2=0 $Y2=0
cc_543 N_A_767_21#_c_561_n N_A_1091_21#_c_927_n 0.0255314f $X=5.465 $Y=1.96
+ $X2=0 $Y2=0
cc_544 N_A_767_21#_c_571_n N_A_1091_21#_c_927_n 0.00284012f $X=6.225 $Y=2.045
+ $X2=0 $Y2=0
cc_545 N_A_767_21#_c_562_n N_A_1091_21#_c_927_n 0.0118491f $X=6.39 $Y=1.275
+ $X2=0 $Y2=0
cc_546 N_A_767_21#_c_563_n N_A_1091_21#_c_927_n 7.13951e-19 $X=6.39 $Y=1.275
+ $X2=0 $Y2=0
cc_547 N_A_767_21#_c_557_n N_A_1091_21#_c_928_n 0.00701575f $X=6.06 $Y=1.6 $X2=0
+ $Y2=0
cc_548 N_A_767_21#_M1012_g N_A_1091_21#_c_928_n 0.00402472f $X=6.52 $Y=0.59
+ $X2=0 $Y2=0
cc_549 N_A_767_21#_c_561_n N_A_1091_21#_c_928_n 0.00868941f $X=5.465 $Y=1.96
+ $X2=0 $Y2=0
cc_550 N_A_767_21#_c_571_n N_A_1091_21#_c_928_n 0.00206251f $X=6.225 $Y=2.045
+ $X2=0 $Y2=0
cc_551 N_A_767_21#_c_562_n N_A_1091_21#_c_928_n 7.58238e-19 $X=6.39 $Y=1.275
+ $X2=0 $Y2=0
cc_552 N_A_767_21#_c_563_n N_A_1091_21#_c_928_n 0.0138069f $X=6.39 $Y=1.275
+ $X2=0 $Y2=0
cc_553 N_A_767_21#_c_557_n N_A_1091_21#_c_929_n 0.0048015f $X=6.06 $Y=1.6 $X2=0
+ $Y2=0
cc_554 N_A_767_21#_M1012_g N_A_1091_21#_c_929_n 0.0129042f $X=6.52 $Y=0.59 $X2=0
+ $Y2=0
cc_555 N_A_767_21#_c_562_n N_A_1091_21#_c_929_n 0.022921f $X=6.39 $Y=1.275 $X2=0
+ $Y2=0
cc_556 N_A_767_21#_c_563_n N_A_1091_21#_c_929_n 0.00151536f $X=6.39 $Y=1.275
+ $X2=0 $Y2=0
cc_557 N_A_767_21#_c_585_n N_A_1091_21#_c_930_n 0.00937466f $X=5.38 $Y=0.745
+ $X2=0 $Y2=0
cc_558 N_A_767_21#_c_561_n N_A_1091_21#_c_930_n 0.00421833f $X=5.465 $Y=1.96
+ $X2=0 $Y2=0
cc_559 N_A_767_21#_M1012_g N_A_1091_21#_c_952_n 0.0108439f $X=6.52 $Y=0.59 $X2=0
+ $Y2=0
cc_560 N_A_767_21#_M1012_g N_A_1091_21#_c_932_n 0.00376448f $X=6.52 $Y=0.59
+ $X2=0 $Y2=0
cc_561 N_A_767_21#_M1009_g N_A_114_57#_M1034_g 0.0347175f $X=4.09 $Y=2.525 $X2=0
+ $Y2=0
cc_562 N_A_767_21#_c_559_n N_A_114_57#_M1034_g 9.07749e-19 $X=4 $Y=1.57 $X2=0
+ $Y2=0
cc_563 N_A_767_21#_c_633_p N_A_114_57#_M1034_g 0.00120751f $X=4.165 $Y=2.415
+ $X2=0 $Y2=0
cc_564 N_A_767_21#_M1009_g N_A_114_57#_c_1117_n 0.0100385f $X=4.09 $Y=2.525
+ $X2=0 $Y2=0
cc_565 N_A_767_21#_M1026_g N_A_114_57#_c_1117_n 0.0103562f $X=5.985 $Y=2.315
+ $X2=0 $Y2=0
cc_566 N_A_767_21#_c_601_p N_A_114_57#_c_1117_n 0.0031423f $X=4.855 $Y=2.415
+ $X2=0 $Y2=0
cc_567 N_A_767_21#_c_633_p N_A_114_57#_c_1117_n 0.00319983f $X=4.165 $Y=2.415
+ $X2=0 $Y2=0
cc_568 N_A_767_21#_c_574_n N_A_114_57#_c_1117_n 0.00461852f $X=4.98 $Y=2.415
+ $X2=0 $Y2=0
cc_569 N_A_767_21#_M1026_g N_A_114_57#_c_1118_n 0.039839f $X=5.985 $Y=2.315
+ $X2=0 $Y2=0
cc_570 N_A_767_21#_c_571_n N_A_114_57#_c_1118_n 0.00421626f $X=6.225 $Y=2.045
+ $X2=0 $Y2=0
cc_571 N_A_767_21#_c_562_n N_A_114_57#_c_1118_n 0.00792902f $X=6.39 $Y=1.275
+ $X2=0 $Y2=0
cc_572 N_A_767_21#_c_563_n N_A_114_57#_c_1118_n 0.00515849f $X=6.39 $Y=1.275
+ $X2=0 $Y2=0
cc_573 N_A_767_21#_c_571_n N_A_114_57#_M1017_g 0.00990695f $X=6.225 $Y=2.045
+ $X2=0 $Y2=0
cc_574 N_A_767_21#_M1012_g N_A_1307_428#_c_1438_n 2.63425e-19 $X=6.52 $Y=0.59
+ $X2=0 $Y2=0
cc_575 N_A_767_21#_c_601_p N_VPWR_M1009_d 0.0125711f $X=4.855 $Y=2.415 $X2=0
+ $Y2=0
cc_576 N_A_767_21#_c_571_n N_VPWR_M1016_d 0.0045064f $X=6.225 $Y=2.045 $X2=0
+ $Y2=0
cc_577 N_A_767_21#_M1009_g N_VPWR_c_1655_n 0.00416523f $X=4.09 $Y=2.525 $X2=0
+ $Y2=0
cc_578 N_A_767_21#_c_601_p N_VPWR_c_1655_n 0.0242478f $X=4.855 $Y=2.415 $X2=0
+ $Y2=0
cc_579 N_A_767_21#_c_574_n N_VPWR_c_1655_n 0.00115075f $X=4.98 $Y=2.415 $X2=0
+ $Y2=0
cc_580 N_A_767_21#_M1026_g N_VPWR_c_1656_n 0.0124229f $X=5.985 $Y=2.315 $X2=0
+ $Y2=0
cc_581 N_A_767_21#_c_612_p N_VPWR_c_1656_n 0.0137891f $X=4.98 $Y=2.33 $X2=0
+ $Y2=0
cc_582 N_A_767_21#_c_571_n N_VPWR_c_1656_n 0.0147371f $X=6.225 $Y=2.045 $X2=0
+ $Y2=0
cc_583 N_A_767_21#_c_574_n N_VPWR_c_1663_n 0.00565285f $X=4.98 $Y=2.415 $X2=0
+ $Y2=0
cc_584 N_A_767_21#_M1009_g N_VPWR_c_1651_n 9.39239e-19 $X=4.09 $Y=2.525 $X2=0
+ $Y2=0
cc_585 N_A_767_21#_M1026_g N_VPWR_c_1651_n 8.51577e-19 $X=5.985 $Y=2.315 $X2=0
+ $Y2=0
cc_586 N_A_767_21#_c_601_p N_VPWR_c_1651_n 0.0117711f $X=4.855 $Y=2.415 $X2=0
+ $Y2=0
cc_587 N_A_767_21#_c_633_p N_VPWR_c_1651_n 0.00962881f $X=4.165 $Y=2.415 $X2=0
+ $Y2=0
cc_588 N_A_767_21#_c_574_n N_VPWR_c_1651_n 0.00685297f $X=4.98 $Y=2.415 $X2=0
+ $Y2=0
cc_589 N_A_767_21#_c_633_p A_755_463# 0.00225479f $X=4.165 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_590 N_A_767_21#_c_586_n A_1046_379# 0.00535996f $X=5.38 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_591 N_A_767_21#_c_561_n A_1046_379# 7.32932e-19 $X=5.465 $Y=1.96 $X2=-0.19
+ $Y2=-0.245
cc_592 N_A_767_21#_c_608_p A_1046_379# 0.00144354f $X=5.465 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_593 N_A_767_21#_c_571_n A_1212_379# 0.0085875f $X=6.225 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_594 N_A_767_21#_c_562_n A_1212_379# 8.9883e-19 $X=6.39 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_595 N_A_767_21#_M1028_g N_VGND_c_1931_n 0.0118921f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_596 N_A_767_21#_M1012_g N_VGND_c_1932_n 0.00449201f $X=6.52 $Y=0.59 $X2=0
+ $Y2=0
cc_597 N_A_767_21#_M1012_g N_VGND_c_1940_n 0.00400146f $X=6.52 $Y=0.59 $X2=0
+ $Y2=0
cc_598 N_A_767_21#_M1028_g N_VGND_c_1942_n 0.00585385f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_599 N_A_767_21#_M1023_d N_VGND_c_1946_n 0.00356992f $X=5.015 $Y=0.235 $X2=0
+ $Y2=0
cc_600 N_A_767_21#_M1028_g N_VGND_c_1946_n 0.0112164f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_601 N_A_767_21#_M1012_g N_VGND_c_1946_n 0.00666425f $X=6.52 $Y=0.59 $X2=0
+ $Y2=0
cc_602 N_A_767_21#_M1023_d N_A_917_47#_c_2077_n 0.00725784f $X=5.015 $Y=0.235
+ $X2=0 $Y2=0
cc_603 N_A_767_21#_c_585_n N_A_917_47#_c_2077_n 0.0264198f $X=5.38 $Y=0.745
+ $X2=0 $Y2=0
cc_604 N_SET_B_M1003_g N_A_617_47#_M1023_g 0.0321335f $X=4.51 $Y=0.555 $X2=0
+ $Y2=0
cc_605 N_SET_B_M1003_g N_A_617_47#_c_834_n 0.00893733f $X=4.51 $Y=0.555 $X2=0
+ $Y2=0
cc_606 N_SET_B_M1003_g N_A_617_47#_M1015_g 5.74421e-19 $X=4.51 $Y=0.555 $X2=0
+ $Y2=0
cc_607 N_SET_B_c_715_n N_A_617_47#_M1015_g 0.0293055f $X=4.725 $Y=1.775 $X2=0
+ $Y2=0
cc_608 N_SET_B_c_723_n N_A_617_47#_M1015_g 9.50455e-19 $X=4.56 $Y=2.035 $X2=0
+ $Y2=0
cc_609 N_SET_B_c_717_n N_A_617_47#_M1015_g 0.00139099f $X=4.54 $Y=1.57 $X2=0
+ $Y2=0
cc_610 N_SET_B_M1003_g N_A_617_47#_c_838_n 0.0166082f $X=4.51 $Y=0.555 $X2=0
+ $Y2=0
cc_611 N_SET_B_c_715_n N_A_617_47#_c_838_n 0.00432362f $X=4.725 $Y=1.775 $X2=0
+ $Y2=0
cc_612 N_SET_B_c_722_n N_A_617_47#_c_838_n 0.00168272f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_613 N_SET_B_c_717_n N_A_617_47#_c_838_n 0.0185151f $X=4.54 $Y=1.57 $X2=0
+ $Y2=0
cc_614 N_SET_B_M1020_g N_A_1091_21#_c_933_n 9.87872e-19 $X=8.45 $Y=0.59 $X2=0
+ $Y2=0
cc_615 N_SET_B_M1020_g N_A_1091_21#_c_934_n 0.0150231f $X=8.45 $Y=0.59 $X2=0
+ $Y2=0
cc_616 N_SET_B_M1020_g N_A_1091_21#_c_940_n 0.00348817f $X=8.45 $Y=0.59 $X2=0
+ $Y2=0
cc_617 N_SET_B_c_715_n N_A_114_57#_c_1117_n 0.0100396f $X=4.725 $Y=1.775 $X2=0
+ $Y2=0
cc_618 N_SET_B_c_722_n N_A_114_57#_c_1118_n 0.00920743f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_619 N_SET_B_c_722_n N_A_114_57#_c_1120_n 0.0068292f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_620 N_SET_B_M1020_g N_A_1545_332#_M1005_g 0.0289429f $X=8.45 $Y=0.59 $X2=0
+ $Y2=0
cc_621 N_SET_B_M1010_g N_A_1545_332#_M1036_g 0.0161649f $X=8.52 $Y=2.57 $X2=0
+ $Y2=0
cc_622 N_SET_B_c_722_n N_A_1545_332#_M1036_g 0.00286838f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_623 N_SET_B_c_719_n N_A_1545_332#_M1036_g 3.50268e-19 $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_624 N_SET_B_M1010_g N_A_1545_332#_c_1272_n 0.00388593f $X=8.52 $Y=2.57 $X2=0
+ $Y2=0
cc_625 N_SET_B_c_722_n N_A_1545_332#_c_1272_n 0.0262812f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_626 N_SET_B_c_724_n N_A_1545_332#_c_1272_n 0.00255335f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_627 N_SET_B_c_718_n N_A_1545_332#_c_1272_n 0.00111008f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_628 N_SET_B_c_719_n N_A_1545_332#_c_1272_n 0.0288863f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_629 N_SET_B_c_722_n N_A_1545_332#_c_1273_n 0.0011552f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_630 N_SET_B_c_724_n N_A_1545_332#_c_1273_n 6.6973e-19 $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_631 N_SET_B_c_718_n N_A_1545_332#_c_1273_n 0.0205842f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_632 N_SET_B_c_719_n N_A_1545_332#_c_1273_n 0.00117787f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_633 N_SET_B_M1010_g N_A_1545_332#_c_1274_n 0.0142689f $X=8.52 $Y=2.57 $X2=0
+ $Y2=0
cc_634 N_SET_B_c_722_n N_A_1545_332#_c_1274_n 0.00855392f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_635 N_SET_B_c_724_n N_A_1545_332#_c_1274_n 0.00258598f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_636 N_SET_B_c_718_n N_A_1545_332#_c_1274_n 7.53951e-19 $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_637 N_SET_B_c_719_n N_A_1545_332#_c_1274_n 0.016037f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_638 N_SET_B_M1010_g N_A_1545_332#_c_1276_n 0.00703392f $X=8.52 $Y=2.57 $X2=0
+ $Y2=0
cc_639 N_SET_B_M1010_g N_A_1545_332#_c_1281_n 0.00532104f $X=8.52 $Y=2.57 $X2=0
+ $Y2=0
cc_640 N_SET_B_c_719_n N_A_1545_332#_c_1281_n 3.56909e-19 $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_641 N_SET_B_M1020_g N_A_1307_428#_M1029_g 0.0522619f $X=8.45 $Y=0.59 $X2=0
+ $Y2=0
cc_642 N_SET_B_c_718_n N_A_1307_428#_M1038_g 0.0234742f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_643 N_SET_B_c_719_n N_A_1307_428#_M1038_g 9.88939e-19 $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_644 N_SET_B_c_722_n N_A_1307_428#_c_1453_n 0.00702661f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_645 N_SET_B_c_722_n N_A_1307_428#_c_1440_n 0.0218471f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_646 N_SET_B_M1020_g N_A_1307_428#_c_1441_n 0.0115456f $X=8.45 $Y=0.59 $X2=0
+ $Y2=0
cc_647 N_SET_B_c_722_n N_A_1307_428#_c_1441_n 0.0136612f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_648 N_SET_B_c_724_n N_A_1307_428#_c_1441_n 0.00153502f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_649 N_SET_B_c_718_n N_A_1307_428#_c_1441_n 0.00247069f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_650 N_SET_B_c_719_n N_A_1307_428#_c_1441_n 0.0203351f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_651 N_SET_B_M1020_g N_A_1307_428#_c_1442_n 0.00301856f $X=8.45 $Y=0.59 $X2=0
+ $Y2=0
cc_652 N_SET_B_c_722_n N_A_1307_428#_c_1448_n 0.006875f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_653 N_SET_B_c_722_n N_A_1307_428#_c_1443_n 0.00361522f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_654 N_SET_B_M1020_g N_A_1307_428#_c_1444_n 5.52915e-19 $X=8.45 $Y=0.59 $X2=0
+ $Y2=0
cc_655 N_SET_B_c_724_n N_A_1307_428#_c_1444_n 3.40683e-19 $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_656 N_SET_B_c_718_n N_A_1307_428#_c_1444_n 0.00188136f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_657 N_SET_B_c_719_n N_A_1307_428#_c_1444_n 0.0229459f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_658 N_SET_B_c_718_n N_A_1307_428#_c_1445_n 0.0190067f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_659 N_SET_B_c_719_n N_A_1307_428#_c_1445_n 3.15876e-19 $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_660 N_SET_B_c_733_n N_VPWR_M1009_d 0.00148894f $X=4.705 $Y=2.035 $X2=0 $Y2=0
cc_661 N_SET_B_c_723_n N_VPWR_M1009_d 0.00474174f $X=4.56 $Y=2.035 $X2=0 $Y2=0
cc_662 N_SET_B_c_724_n N_VPWR_M1036_d 0.00158932f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_663 N_SET_B_c_719_n N_VPWR_M1036_d 8.96001e-19 $X=8.43 $Y=1.825 $X2=0 $Y2=0
cc_664 N_SET_B_c_715_n N_VPWR_c_1655_n 0.00384677f $X=4.725 $Y=1.775 $X2=0 $Y2=0
cc_665 N_SET_B_c_722_n N_VPWR_c_1656_n 0.00264794f $X=8.255 $Y=2.035 $X2=0 $Y2=0
cc_666 N_SET_B_M1010_g N_VPWR_c_1657_n 0.00924924f $X=8.52 $Y=2.57 $X2=0 $Y2=0
cc_667 N_SET_B_M1010_g N_VPWR_c_1665_n 0.0040395f $X=8.52 $Y=2.57 $X2=0 $Y2=0
cc_668 N_SET_B_c_715_n N_VPWR_c_1651_n 9.39239e-19 $X=4.725 $Y=1.775 $X2=0 $Y2=0
cc_669 N_SET_B_M1010_g N_VPWR_c_1651_n 0.00408208f $X=8.52 $Y=2.57 $X2=0 $Y2=0
cc_670 N_SET_B_M1003_g N_VGND_c_1931_n 0.00716677f $X=4.51 $Y=0.555 $X2=0 $Y2=0
cc_671 N_SET_B_M1020_g N_VGND_c_1933_n 0.00896652f $X=8.45 $Y=0.59 $X2=0 $Y2=0
cc_672 N_SET_B_M1003_g N_VGND_c_1938_n 0.0054778f $X=4.51 $Y=0.555 $X2=0 $Y2=0
cc_673 N_SET_B_M1020_g N_VGND_c_1943_n 0.00514823f $X=8.45 $Y=0.59 $X2=0 $Y2=0
cc_674 N_SET_B_M1003_g N_VGND_c_1946_n 0.0103714f $X=4.51 $Y=0.555 $X2=0 $Y2=0
cc_675 N_SET_B_M1020_g N_VGND_c_1946_n 0.0106184f $X=8.45 $Y=0.59 $X2=0 $Y2=0
cc_676 N_SET_B_M1003_g N_A_917_47#_c_2075_n 0.00628215f $X=4.51 $Y=0.555 $X2=0
+ $Y2=0
cc_677 N_SET_B_M1003_g N_A_917_47#_c_2080_n 0.00331806f $X=4.51 $Y=0.555 $X2=0
+ $Y2=0
cc_678 N_SET_B_M1020_g N_A_1705_54#_c_2105_n 0.00423725f $X=8.45 $Y=0.59 $X2=0
+ $Y2=0
cc_679 N_A_617_47#_M1023_g N_A_1091_21#_c_922_n 0.0218838f $X=4.94 $Y=0.555
+ $X2=0 $Y2=0
cc_680 N_A_617_47#_c_834_n N_A_1091_21#_M1016_g 0.00422241f $X=5.155 $Y=1.385
+ $X2=0 $Y2=0
cc_681 N_A_617_47#_M1015_g N_A_1091_21#_M1016_g 0.0747717f $X=5.155 $Y=2.315
+ $X2=0 $Y2=0
cc_682 N_A_617_47#_c_834_n N_A_1091_21#_c_928_n 0.0193242f $X=5.155 $Y=1.385
+ $X2=0 $Y2=0
cc_683 N_A_617_47#_c_838_n N_A_1091_21#_c_928_n 3.08461e-19 $X=4.915 $Y=1.14
+ $X2=0 $Y2=0
cc_684 N_A_617_47#_c_837_n N_A_114_57#_c_1114_n 0.00416667f $X=3.615 $Y=2.41
+ $X2=0 $Y2=0
cc_685 N_A_617_47#_c_836_n N_A_114_57#_M1021_g 7.44203e-19 $X=3.615 $Y=1.055
+ $X2=0 $Y2=0
cc_686 N_A_617_47#_c_837_n N_A_114_57#_M1034_g 0.0154131f $X=3.615 $Y=2.41 $X2=0
+ $Y2=0
cc_687 N_A_617_47#_M1015_g N_A_114_57#_c_1117_n 0.0103003f $X=5.155 $Y=2.315
+ $X2=0 $Y2=0
cc_688 N_A_617_47#_c_837_n N_VPWR_c_1655_n 0.00229416f $X=3.615 $Y=2.41 $X2=0
+ $Y2=0
cc_689 N_A_617_47#_M1015_g N_VPWR_c_1656_n 0.00180485f $X=5.155 $Y=2.315 $X2=0
+ $Y2=0
cc_690 N_A_617_47#_c_837_n N_VPWR_c_1667_n 0.00813654f $X=3.615 $Y=2.41 $X2=0
+ $Y2=0
cc_691 N_A_617_47#_M1015_g N_VPWR_c_1651_n 9.39239e-19 $X=5.155 $Y=2.315 $X2=0
+ $Y2=0
cc_692 N_A_617_47#_c_837_n N_VPWR_c_1651_n 0.0100775f $X=3.615 $Y=2.41 $X2=0
+ $Y2=0
cc_693 N_A_617_47#_c_836_n N_A_531_47#_c_1799_n 0.00471886f $X=3.615 $Y=1.055
+ $X2=0 $Y2=0
cc_694 N_A_617_47#_c_837_n N_A_531_47#_c_1796_n 0.0202193f $X=3.615 $Y=2.41
+ $X2=0 $Y2=0
cc_695 N_A_617_47#_c_836_n N_A_531_47#_c_1793_n 0.0132041f $X=3.615 $Y=1.055
+ $X2=0 $Y2=0
cc_696 N_A_617_47#_c_848_n N_A_531_47#_c_1793_n 0.0162668f $X=3.305 $Y=0.455
+ $X2=0 $Y2=0
cc_697 N_A_617_47#_c_836_n N_A_531_47#_c_1795_n 0.00369954f $X=3.615 $Y=1.055
+ $X2=0 $Y2=0
cc_698 N_A_617_47#_c_837_n N_A_531_47#_c_1795_n 0.0559215f $X=3.615 $Y=2.41
+ $X2=0 $Y2=0
cc_699 N_A_617_47#_c_850_n N_A_531_47#_c_1795_n 0.0130061f $X=3.615 $Y=1.14
+ $X2=0 $Y2=0
cc_700 N_A_617_47#_c_837_n N_A_531_47#_c_1798_n 0.0155357f $X=3.615 $Y=2.41
+ $X2=0 $Y2=0
cc_701 N_A_617_47#_c_836_n N_VGND_c_1931_n 0.0107508f $X=3.615 $Y=1.055 $X2=0
+ $Y2=0
cc_702 N_A_617_47#_c_838_n N_VGND_c_1931_n 0.0241496f $X=4.915 $Y=1.14 $X2=0
+ $Y2=0
cc_703 N_A_617_47#_c_848_n N_VGND_c_1931_n 0.0147262f $X=3.305 $Y=0.455 $X2=0
+ $Y2=0
cc_704 N_A_617_47#_M1023_g N_VGND_c_1938_n 0.0035993f $X=4.94 $Y=0.555 $X2=0
+ $Y2=0
cc_705 N_A_617_47#_c_848_n N_VGND_c_1942_n 0.0244899f $X=3.305 $Y=0.455 $X2=0
+ $Y2=0
cc_706 N_A_617_47#_M1021_d N_VGND_c_1946_n 0.00325445f $X=3.085 $Y=0.235 $X2=0
+ $Y2=0
cc_707 N_A_617_47#_M1023_g N_VGND_c_1946_n 0.0058413f $X=4.94 $Y=0.555 $X2=0
+ $Y2=0
cc_708 N_A_617_47#_c_848_n N_VGND_c_1946_n 0.0195235f $X=3.305 $Y=0.455 $X2=0
+ $Y2=0
cc_709 N_A_617_47#_c_848_n A_719_47# 0.00267563f $X=3.305 $Y=0.455 $X2=-0.19
+ $Y2=-0.245
cc_710 N_A_617_47#_M1023_g N_A_917_47#_c_2075_n 0.00808861f $X=4.94 $Y=0.555
+ $X2=0 $Y2=0
cc_711 N_A_617_47#_c_838_n N_A_917_47#_c_2075_n 0.0194758f $X=4.915 $Y=1.14
+ $X2=0 $Y2=0
cc_712 N_A_617_47#_M1023_g N_A_917_47#_c_2080_n 0.0018944f $X=4.94 $Y=0.555
+ $X2=0 $Y2=0
cc_713 N_A_617_47#_M1023_g N_A_917_47#_c_2076_n 4.02471e-19 $X=4.94 $Y=0.555
+ $X2=0 $Y2=0
cc_714 N_A_617_47#_M1023_g N_A_917_47#_c_2077_n 0.00923314f $X=4.94 $Y=0.555
+ $X2=0 $Y2=0
cc_715 N_A_617_47#_c_834_n N_A_917_47#_c_2077_n 9.35671e-19 $X=5.155 $Y=1.385
+ $X2=0 $Y2=0
cc_716 N_A_617_47#_c_838_n N_A_917_47#_c_2077_n 0.00369659f $X=4.915 $Y=1.14
+ $X2=0 $Y2=0
cc_717 N_A_1091_21#_M1016_g N_A_114_57#_c_1117_n 0.0103107f $X=5.545 $Y=2.315
+ $X2=0 $Y2=0
cc_718 N_A_1091_21#_c_931_n N_A_114_57#_M1004_g 0.00767583f $X=7.665 $Y=0.35
+ $X2=0 $Y2=0
cc_719 N_A_1091_21#_c_933_n N_A_114_57#_M1004_g 0.00534318f $X=7.75 $Y=0.945
+ $X2=0 $Y2=0
cc_720 N_A_1091_21#_c_935_n N_A_114_57#_M1004_g 0.00104127f $X=7.835 $Y=1.03
+ $X2=0 $Y2=0
cc_721 N_A_1091_21#_c_936_n N_A_1545_332#_M1029_d 0.00763252f $X=9.68 $Y=0.86
+ $X2=-0.19 $Y2=-0.245
cc_722 N_A_1091_21#_c_931_n N_A_1545_332#_M1005_g 0.00365588f $X=7.665 $Y=0.35
+ $X2=0 $Y2=0
cc_723 N_A_1091_21#_c_933_n N_A_1545_332#_M1005_g 0.0123324f $X=7.75 $Y=0.945
+ $X2=0 $Y2=0
cc_724 N_A_1091_21#_c_934_n N_A_1545_332#_M1005_g 0.00648937f $X=8.74 $Y=1.03
+ $X2=0 $Y2=0
cc_725 N_A_1091_21#_c_935_n N_A_1545_332#_M1005_g 0.00387931f $X=7.835 $Y=1.03
+ $X2=0 $Y2=0
cc_726 N_A_1091_21#_c_946_n N_A_1545_332#_M1027_g 2.92669e-19 $X=10.23 $Y=1.86
+ $X2=0 $Y2=0
cc_727 N_A_1091_21#_M1001_g N_A_1545_332#_c_1276_n 0.00158681f $X=9.45 $Y=2.57
+ $X2=0 $Y2=0
cc_728 N_A_1091_21#_M1001_g N_A_1545_332#_c_1263_n 0.0137656f $X=9.45 $Y=2.57
+ $X2=0 $Y2=0
cc_729 N_A_1091_21#_c_926_n N_A_1545_332#_c_1263_n 0.00708588f $X=9.375 $Y=1.51
+ $X2=0 $Y2=0
cc_730 N_A_1091_21#_c_938_n N_A_1545_332#_c_1263_n 0.0154334f $X=9.845 $Y=1.39
+ $X2=0 $Y2=0
cc_731 N_A_1091_21#_c_945_n N_A_1545_332#_c_1263_n 0.02413f $X=10.01 $Y=1.86
+ $X2=0 $Y2=0
cc_732 N_A_1091_21#_M1025_s N_A_1545_332#_c_1279_n 0.00328558f $X=10.085
+ $Y=1.715 $X2=0 $Y2=0
cc_733 N_A_1091_21#_M1001_g N_A_1545_332#_c_1279_n 0.00738985f $X=9.45 $Y=2.57
+ $X2=0 $Y2=0
cc_734 N_A_1091_21#_c_926_n N_A_1545_332#_c_1279_n 0.00343408f $X=9.375 $Y=1.51
+ $X2=0 $Y2=0
cc_735 N_A_1091_21#_c_939_n N_A_1545_332#_c_1279_n 0.00106768f $X=9.845 $Y=1.39
+ $X2=0 $Y2=0
cc_736 N_A_1091_21#_c_945_n N_A_1545_332#_c_1279_n 0.0265884f $X=10.01 $Y=1.86
+ $X2=0 $Y2=0
cc_737 N_A_1091_21#_c_946_n N_A_1545_332#_c_1279_n 0.0240404f $X=10.23 $Y=1.86
+ $X2=0 $Y2=0
cc_738 N_A_1091_21#_c_946_n N_A_1545_332#_c_1264_n 0.0151658f $X=10.23 $Y=1.86
+ $X2=0 $Y2=0
cc_739 N_A_1091_21#_M1001_g N_A_1545_332#_c_1281_n 6.08907e-19 $X=9.45 $Y=2.57
+ $X2=0 $Y2=0
cc_740 N_A_1091_21#_M1014_g N_A_1545_332#_c_1265_n 0.00427829f $X=9.465 $Y=0.59
+ $X2=0 $Y2=0
cc_741 N_A_1091_21#_c_926_n N_A_1545_332#_c_1265_n 0.00905234f $X=9.375 $Y=1.51
+ $X2=0 $Y2=0
cc_742 N_A_1091_21#_c_936_n N_A_1545_332#_c_1265_n 0.0286714f $X=9.68 $Y=0.86
+ $X2=0 $Y2=0
cc_743 N_A_1091_21#_c_938_n N_A_1545_332#_c_1265_n 0.0228394f $X=9.845 $Y=1.39
+ $X2=0 $Y2=0
cc_744 N_A_1091_21#_M1001_g N_A_1545_332#_c_1328_n 0.0131285f $X=9.45 $Y=2.57
+ $X2=0 $Y2=0
cc_745 N_A_1091_21#_c_931_n N_A_1307_428#_M1013_d 0.00241744f $X=7.665 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_746 N_A_1091_21#_M1014_g N_A_1307_428#_M1029_g 0.0357109f $X=9.465 $Y=0.59
+ $X2=0 $Y2=0
cc_747 N_A_1091_21#_c_926_n N_A_1307_428#_M1029_g 0.00301135f $X=9.375 $Y=1.51
+ $X2=0 $Y2=0
cc_748 N_A_1091_21#_c_934_n N_A_1307_428#_M1029_g 3.0806e-19 $X=8.74 $Y=1.03
+ $X2=0 $Y2=0
cc_749 N_A_1091_21#_c_936_n N_A_1307_428#_M1029_g 0.00655432f $X=9.68 $Y=0.86
+ $X2=0 $Y2=0
cc_750 N_A_1091_21#_c_940_n N_A_1307_428#_M1029_g 0.0112619f $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_751 N_A_1091_21#_M1001_g N_A_1307_428#_M1038_g 0.0539804f $X=9.45 $Y=2.57
+ $X2=0 $Y2=0
cc_752 N_A_1091_21#_c_929_n N_A_1307_428#_c_1438_n 0.0119004f $X=6.57 $Y=0.845
+ $X2=0 $Y2=0
cc_753 N_A_1091_21#_c_952_n N_A_1307_428#_c_1438_n 0.00904598f $X=6.655 $Y=0.76
+ $X2=0 $Y2=0
cc_754 N_A_1091_21#_c_931_n N_A_1307_428#_c_1438_n 0.0299123f $X=7.665 $Y=0.35
+ $X2=0 $Y2=0
cc_755 N_A_1091_21#_c_933_n N_A_1307_428#_c_1438_n 0.0232206f $X=7.75 $Y=0.945
+ $X2=0 $Y2=0
cc_756 N_A_1091_21#_c_933_n N_A_1307_428#_c_1439_n 9.5925e-19 $X=7.75 $Y=0.945
+ $X2=0 $Y2=0
cc_757 N_A_1091_21#_c_935_n N_A_1307_428#_c_1439_n 0.01314f $X=7.835 $Y=1.03
+ $X2=0 $Y2=0
cc_758 N_A_1091_21#_c_934_n N_A_1307_428#_c_1441_n 0.0602894f $X=8.74 $Y=1.03
+ $X2=0 $Y2=0
cc_759 N_A_1091_21#_c_935_n N_A_1307_428#_c_1441_n 0.0121865f $X=7.835 $Y=1.03
+ $X2=0 $Y2=0
cc_760 N_A_1091_21#_c_940_n N_A_1307_428#_c_1441_n 0.0119492f $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_761 N_A_1091_21#_c_926_n N_A_1307_428#_c_1444_n 3.74136e-19 $X=9.375 $Y=1.51
+ $X2=0 $Y2=0
cc_762 N_A_1091_21#_c_926_n N_A_1307_428#_c_1445_n 0.0180717f $X=9.375 $Y=1.51
+ $X2=0 $Y2=0
cc_763 N_A_1091_21#_c_936_n N_A_1307_428#_c_1445_n 0.00330102f $X=9.68 $Y=0.86
+ $X2=0 $Y2=0
cc_764 N_A_1091_21#_c_938_n N_RESET_B_M1025_g 0.00189804f $X=9.845 $Y=1.39 $X2=0
+ $Y2=0
cc_765 N_A_1091_21#_c_939_n N_RESET_B_M1025_g 0.00566261f $X=9.845 $Y=1.39 $X2=0
+ $Y2=0
cc_766 N_A_1091_21#_c_946_n N_RESET_B_M1025_g 0.00579214f $X=10.23 $Y=1.86 $X2=0
+ $Y2=0
cc_767 N_A_1091_21#_c_937_n RESET_B 0.0130519f $X=9.845 $Y=1 $X2=0 $Y2=0
cc_768 N_A_1091_21#_c_938_n RESET_B 0.0241509f $X=9.845 $Y=1.39 $X2=0 $Y2=0
cc_769 N_A_1091_21#_c_939_n RESET_B 0.00178487f $X=9.845 $Y=1.39 $X2=0 $Y2=0
cc_770 N_A_1091_21#_c_946_n RESET_B 0.0143797f $X=10.23 $Y=1.86 $X2=0 $Y2=0
cc_771 N_A_1091_21#_M1014_g N_RESET_B_c_1560_n 3.7931e-19 $X=9.465 $Y=0.59 $X2=0
+ $Y2=0
cc_772 N_A_1091_21#_c_937_n N_RESET_B_c_1560_n 9.81404e-19 $X=9.845 $Y=1 $X2=0
+ $Y2=0
cc_773 N_A_1091_21#_c_938_n N_RESET_B_c_1560_n 5.28667e-19 $X=9.845 $Y=1.39
+ $X2=0 $Y2=0
cc_774 N_A_1091_21#_c_939_n N_RESET_B_c_1560_n 0.0190891f $X=9.845 $Y=1.39 $X2=0
+ $Y2=0
cc_775 N_A_1091_21#_c_946_n N_RESET_B_c_1560_n 0.00339756f $X=10.23 $Y=1.86
+ $X2=0 $Y2=0
cc_776 N_A_1091_21#_c_937_n N_RESET_B_c_1561_n 0.00498607f $X=9.845 $Y=1 $X2=0
+ $Y2=0
cc_777 N_A_1091_21#_c_938_n N_RESET_B_c_1561_n 0.00530447f $X=9.845 $Y=1.39
+ $X2=0 $Y2=0
cc_778 N_A_1091_21#_M1016_g N_VPWR_c_1656_n 0.011889f $X=5.545 $Y=2.315 $X2=0
+ $Y2=0
cc_779 N_A_1091_21#_M1001_g N_VPWR_c_1658_n 0.0142303f $X=9.45 $Y=2.57 $X2=0
+ $Y2=0
cc_780 N_A_1091_21#_M1001_g N_VPWR_c_1665_n 0.0040395f $X=9.45 $Y=2.57 $X2=0
+ $Y2=0
cc_781 N_A_1091_21#_M1016_g N_VPWR_c_1651_n 7.88961e-19 $X=5.545 $Y=2.315 $X2=0
+ $Y2=0
cc_782 N_A_1091_21#_M1001_g N_VPWR_c_1651_n 0.00777113f $X=9.45 $Y=2.57 $X2=0
+ $Y2=0
cc_783 N_A_1091_21#_c_929_n N_VGND_M1012_s 0.00309765f $X=6.57 $Y=0.845 $X2=0
+ $Y2=0
cc_784 N_A_1091_21#_c_922_n N_VGND_c_1932_n 0.00224464f $X=5.53 $Y=0.985 $X2=0
+ $Y2=0
cc_785 N_A_1091_21#_c_929_n N_VGND_c_1932_n 0.0186154f $X=6.57 $Y=0.845 $X2=0
+ $Y2=0
cc_786 N_A_1091_21#_c_932_n N_VGND_c_1932_n 0.00699226f $X=6.74 $Y=0.35 $X2=0
+ $Y2=0
cc_787 N_A_1091_21#_c_931_n N_VGND_c_1933_n 0.0111412f $X=7.665 $Y=0.35 $X2=0
+ $Y2=0
cc_788 N_A_1091_21#_c_933_n N_VGND_c_1933_n 0.0186051f $X=7.75 $Y=0.945 $X2=0
+ $Y2=0
cc_789 N_A_1091_21#_c_934_n N_VGND_c_1933_n 0.0196257f $X=8.74 $Y=1.03 $X2=0
+ $Y2=0
cc_790 N_A_1091_21#_c_937_n N_VGND_c_1934_n 0.0148459f $X=9.845 $Y=1 $X2=0 $Y2=0
cc_791 N_A_1091_21#_c_922_n N_VGND_c_1938_n 0.00359964f $X=5.53 $Y=0.985 $X2=0
+ $Y2=0
cc_792 N_A_1091_21#_c_929_n N_VGND_c_1938_n 0.00176484f $X=6.57 $Y=0.845 $X2=0
+ $Y2=0
cc_793 N_A_1091_21#_c_930_n N_VGND_c_1938_n 0.00164511f $X=6.015 $Y=0.845 $X2=0
+ $Y2=0
cc_794 N_A_1091_21#_c_929_n N_VGND_c_1940_n 0.00192901f $X=6.57 $Y=0.845 $X2=0
+ $Y2=0
cc_795 N_A_1091_21#_c_931_n N_VGND_c_1940_n 0.0670649f $X=7.665 $Y=0.35 $X2=0
+ $Y2=0
cc_796 N_A_1091_21#_c_932_n N_VGND_c_1940_n 0.0113565f $X=6.74 $Y=0.35 $X2=0
+ $Y2=0
cc_797 N_A_1091_21#_M1014_g N_VGND_c_1943_n 0.00337062f $X=9.465 $Y=0.59 $X2=0
+ $Y2=0
cc_798 N_A_1091_21#_c_937_n N_VGND_c_1943_n 0.00632222f $X=9.845 $Y=1 $X2=0
+ $Y2=0
cc_799 N_A_1091_21#_c_922_n N_VGND_c_1946_n 0.007043f $X=5.53 $Y=0.985 $X2=0
+ $Y2=0
cc_800 N_A_1091_21#_M1014_g N_VGND_c_1946_n 0.0063727f $X=9.465 $Y=0.59 $X2=0
+ $Y2=0
cc_801 N_A_1091_21#_c_929_n N_VGND_c_1946_n 0.00827129f $X=6.57 $Y=0.845 $X2=0
+ $Y2=0
cc_802 N_A_1091_21#_c_930_n N_VGND_c_1946_n 0.00336579f $X=6.015 $Y=0.845 $X2=0
+ $Y2=0
cc_803 N_A_1091_21#_c_931_n N_VGND_c_1946_n 0.0404529f $X=7.665 $Y=0.35 $X2=0
+ $Y2=0
cc_804 N_A_1091_21#_c_932_n N_VGND_c_1946_n 0.00645868f $X=6.74 $Y=0.35 $X2=0
+ $Y2=0
cc_805 N_A_1091_21#_c_937_n N_VGND_c_1946_n 0.0192115f $X=9.845 $Y=1 $X2=0 $Y2=0
cc_806 N_A_1091_21#_c_930_n N_A_917_47#_M1019_d 0.00337953f $X=6.015 $Y=0.845
+ $X2=0 $Y2=0
cc_807 N_A_1091_21#_c_922_n N_A_917_47#_c_2075_n 9.44341e-19 $X=5.53 $Y=0.985
+ $X2=0 $Y2=0
cc_808 N_A_1091_21#_c_922_n N_A_917_47#_c_2076_n 0.00356091f $X=5.53 $Y=0.985
+ $X2=0 $Y2=0
cc_809 N_A_1091_21#_c_928_n N_A_917_47#_c_2076_n 0.00365957f $X=5.85 $Y=1.15
+ $X2=0 $Y2=0
cc_810 N_A_1091_21#_c_930_n N_A_917_47#_c_2076_n 0.0108688f $X=6.015 $Y=0.845
+ $X2=0 $Y2=0
cc_811 N_A_1091_21#_c_922_n N_A_917_47#_c_2077_n 0.00876745f $X=5.53 $Y=0.985
+ $X2=0 $Y2=0
cc_812 N_A_1091_21#_c_929_n A_1319_54# 0.00141319f $X=6.57 $Y=0.845 $X2=-0.19
+ $Y2=-0.245
cc_813 N_A_1091_21#_c_952_n A_1319_54# 0.00328555f $X=6.655 $Y=0.76 $X2=-0.19
+ $Y2=-0.245
cc_814 N_A_1091_21#_c_931_n A_1319_54# 0.00141176f $X=7.665 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_815 N_A_1091_21#_c_933_n A_1499_98# 0.00395864f $X=7.75 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_816 N_A_1091_21#_c_940_n N_A_1705_54#_M1020_d 0.00169355f $X=8.825 $Y=0.86
+ $X2=-0.19 $Y2=-0.245
cc_817 N_A_1091_21#_c_936_n N_A_1705_54#_M1014_d 8.77141e-19 $X=9.68 $Y=0.86
+ $X2=0 $Y2=0
cc_818 N_A_1091_21#_c_937_n N_A_1705_54#_M1014_d 0.00230654f $X=9.845 $Y=1 $X2=0
+ $Y2=0
cc_819 N_A_1091_21#_M1014_g N_A_1705_54#_c_2105_n 0.013256f $X=9.465 $Y=0.59
+ $X2=0 $Y2=0
cc_820 N_A_1091_21#_c_934_n N_A_1705_54#_c_2105_n 0.00961922f $X=8.74 $Y=1.03
+ $X2=0 $Y2=0
cc_821 N_A_1091_21#_c_936_n N_A_1705_54#_c_2105_n 0.0413196f $X=9.68 $Y=0.86
+ $X2=0 $Y2=0
cc_822 N_A_1091_21#_c_937_n N_A_1705_54#_c_2105_n 0.0130263f $X=9.845 $Y=1 $X2=0
+ $Y2=0
cc_823 N_A_1091_21#_c_939_n N_A_1705_54#_c_2105_n 6.04385e-19 $X=9.845 $Y=1.39
+ $X2=0 $Y2=0
cc_824 N_A_1091_21#_c_940_n N_A_1705_54#_c_2105_n 0.00771995f $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_825 N_A_114_57#_M1004_g N_A_1545_332#_M1005_g 0.0661932f $X=7.42 $Y=0.7 $X2=0
+ $Y2=0
cc_826 N_A_114_57#_M1004_g N_A_1545_332#_c_1273_n 0.00941943f $X=7.42 $Y=0.7
+ $X2=0 $Y2=0
cc_827 N_A_114_57#_M1004_g N_A_1307_428#_c_1438_n 0.0121832f $X=7.42 $Y=0.7
+ $X2=0 $Y2=0
cc_828 N_A_114_57#_M1004_g N_A_1307_428#_c_1439_n 0.00967373f $X=7.42 $Y=0.7
+ $X2=0 $Y2=0
cc_829 N_A_114_57#_c_1120_n N_A_1307_428#_c_1440_n 0.00647186f $X=7.345 $Y=1.755
+ $X2=0 $Y2=0
cc_830 N_A_114_57#_M1004_g N_A_1307_428#_c_1440_n 0.00437259f $X=7.42 $Y=0.7
+ $X2=0 $Y2=0
cc_831 N_A_114_57#_c_1118_n N_A_1307_428#_c_1448_n 0.00217592f $X=6.46 $Y=2.065
+ $X2=0 $Y2=0
cc_832 N_A_114_57#_M1017_g N_A_1307_428#_c_1448_n 0.0113227f $X=6.46 $Y=2.56
+ $X2=0 $Y2=0
cc_833 N_A_114_57#_c_1120_n N_A_1307_428#_c_1443_n 0.00117762f $X=7.345 $Y=1.755
+ $X2=0 $Y2=0
cc_834 N_A_114_57#_M1004_g N_A_1307_428#_c_1443_n 0.0071465f $X=7.42 $Y=0.7
+ $X2=0 $Y2=0
cc_835 N_A_114_57#_c_1124_n N_VPWR_c_1653_n 0.0258905f $X=0.86 $Y=2.55 $X2=0
+ $Y2=0
cc_836 N_A_114_57#_M1011_g N_VPWR_c_1654_n 0.00795579f $X=1.635 $Y=2.635 $X2=0
+ $Y2=0
cc_837 N_A_114_57#_c_1114_n N_VPWR_c_1654_n 0.0243149f $X=3.625 $Y=3.15 $X2=0
+ $Y2=0
cc_838 N_A_114_57#_M1034_g N_VPWR_c_1655_n 0.00585489f $X=3.7 $Y=2.525 $X2=0
+ $Y2=0
cc_839 N_A_114_57#_c_1117_n N_VPWR_c_1655_n 0.0252872f $X=6.385 $Y=3.15 $X2=0
+ $Y2=0
cc_840 N_A_114_57#_c_1117_n N_VPWR_c_1656_n 0.0254833f $X=6.385 $Y=3.15 $X2=0
+ $Y2=0
cc_841 N_A_114_57#_M1017_g N_VPWR_c_1656_n 0.00833493f $X=6.46 $Y=2.56 $X2=0
+ $Y2=0
cc_842 N_A_114_57#_c_1115_n N_VPWR_c_1661_n 0.00762896f $X=1.71 $Y=3.15 $X2=0
+ $Y2=0
cc_843 N_A_114_57#_c_1124_n N_VPWR_c_1661_n 0.0220321f $X=0.86 $Y=2.55 $X2=0
+ $Y2=0
cc_844 N_A_114_57#_c_1117_n N_VPWR_c_1663_n 0.0324598f $X=6.385 $Y=3.15 $X2=0
+ $Y2=0
cc_845 N_A_114_57#_c_1114_n N_VPWR_c_1667_n 0.0697509f $X=3.625 $Y=3.15 $X2=0
+ $Y2=0
cc_846 N_A_114_57#_c_1117_n N_VPWR_c_1668_n 0.0223877f $X=6.385 $Y=3.15 $X2=0
+ $Y2=0
cc_847 N_A_114_57#_c_1114_n N_VPWR_c_1651_n 0.0629818f $X=3.625 $Y=3.15 $X2=0
+ $Y2=0
cc_848 N_A_114_57#_c_1115_n N_VPWR_c_1651_n 0.0106041f $X=1.71 $Y=3.15 $X2=0
+ $Y2=0
cc_849 N_A_114_57#_c_1117_n N_VPWR_c_1651_n 0.086158f $X=6.385 $Y=3.15 $X2=0
+ $Y2=0
cc_850 N_A_114_57#_c_1122_n N_VPWR_c_1651_n 0.00671854f $X=3.7 $Y=3.15 $X2=0
+ $Y2=0
cc_851 N_A_114_57#_c_1124_n N_VPWR_c_1651_n 0.0125808f $X=0.86 $Y=2.55 $X2=0
+ $Y2=0
cc_852 N_A_114_57#_M1021_g N_A_531_47#_c_1799_n 0.00970231f $X=3.01 $Y=0.445
+ $X2=0 $Y2=0
cc_853 N_A_114_57#_c_1114_n N_A_531_47#_c_1796_n 0.00570991f $X=3.625 $Y=3.15
+ $X2=0 $Y2=0
cc_854 N_A_114_57#_M1034_g N_A_531_47#_c_1796_n 2.52091e-19 $X=3.7 $Y=2.525
+ $X2=0 $Y2=0
cc_855 N_A_114_57#_M1021_g N_A_531_47#_c_1793_n 0.00812597f $X=3.01 $Y=0.445
+ $X2=0 $Y2=0
cc_856 N_A_114_57#_c_1105_n N_A_531_47#_c_1794_n 0.00688772f $X=2.935 $Y=1.23
+ $X2=0 $Y2=0
cc_857 N_A_114_57#_M1021_g N_A_531_47#_c_1794_n 0.0035575f $X=3.01 $Y=0.445
+ $X2=0 $Y2=0
cc_858 N_A_114_57#_M1021_g N_A_531_47#_c_1795_n 0.00562216f $X=3.01 $Y=0.445
+ $X2=0 $Y2=0
cc_859 N_A_114_57#_c_1111_n N_VGND_c_1929_n 0.0179429f $X=0.71 $Y=0.495 $X2=0
+ $Y2=0
cc_860 N_A_114_57#_M1008_g N_VGND_c_1930_n 0.00666045f $X=1.485 $Y=0.445 $X2=0
+ $Y2=0
cc_861 N_A_114_57#_M1008_g N_VGND_c_1936_n 0.00359757f $X=1.485 $Y=0.445 $X2=0
+ $Y2=0
cc_862 N_A_114_57#_c_1111_n N_VGND_c_1936_n 0.0217479f $X=0.71 $Y=0.495 $X2=0
+ $Y2=0
cc_863 N_A_114_57#_M1004_g N_VGND_c_1940_n 7.36939e-19 $X=7.42 $Y=0.7 $X2=0
+ $Y2=0
cc_864 N_A_114_57#_M1021_g N_VGND_c_1942_n 0.00549284f $X=3.01 $Y=0.445 $X2=0
+ $Y2=0
cc_865 N_A_114_57#_M1008_g N_VGND_c_1946_n 0.00822274f $X=1.485 $Y=0.445 $X2=0
+ $Y2=0
cc_866 N_A_114_57#_M1021_g N_VGND_c_1946_n 0.00656797f $X=3.01 $Y=0.445 $X2=0
+ $Y2=0
cc_867 N_A_114_57#_c_1111_n N_VGND_c_1946_n 0.0125215f $X=0.71 $Y=0.495 $X2=0
+ $Y2=0
cc_868 N_A_1545_332#_c_1263_n N_A_1307_428#_M1029_g 0.00120994f $X=9.4 $Y=2.145
+ $X2=0 $Y2=0
cc_869 N_A_1545_332#_c_1265_n N_A_1307_428#_M1029_g 0.00618282f $X=9.4 $Y=1.29
+ $X2=0 $Y2=0
cc_870 N_A_1545_332#_c_1276_n N_A_1307_428#_M1038_g 0.0107209f $X=8.825 $Y=2.845
+ $X2=0 $Y2=0
cc_871 N_A_1545_332#_c_1277_n N_A_1307_428#_M1038_g 0.0125753f $X=9.315 $Y=2.26
+ $X2=0 $Y2=0
cc_872 N_A_1545_332#_c_1263_n N_A_1307_428#_M1038_g 0.00353264f $X=9.4 $Y=2.145
+ $X2=0 $Y2=0
cc_873 N_A_1545_332#_c_1281_n N_A_1307_428#_M1038_g 0.00332606f $X=8.825 $Y=2.31
+ $X2=0 $Y2=0
cc_874 N_A_1545_332#_M1005_g N_A_1307_428#_c_1438_n 3.47e-19 $X=7.81 $Y=0.7
+ $X2=0 $Y2=0
cc_875 N_A_1545_332#_M1036_g N_A_1307_428#_c_1453_n 0.00416807f $X=7.81 $Y=2.77
+ $X2=0 $Y2=0
cc_876 N_A_1545_332#_M1005_g N_A_1307_428#_c_1439_n 0.00144986f $X=7.81 $Y=0.7
+ $X2=0 $Y2=0
cc_877 N_A_1545_332#_M1005_g N_A_1307_428#_c_1440_n 0.00371296f $X=7.81 $Y=0.7
+ $X2=0 $Y2=0
cc_878 N_A_1545_332#_M1036_g N_A_1307_428#_c_1440_n 0.00664062f $X=7.81 $Y=2.77
+ $X2=0 $Y2=0
cc_879 N_A_1545_332#_c_1272_n N_A_1307_428#_c_1440_n 0.0466938f $X=7.89 $Y=1.825
+ $X2=0 $Y2=0
cc_880 N_A_1545_332#_c_1273_n N_A_1307_428#_c_1440_n 0.00461382f $X=7.89
+ $Y=1.825 $X2=0 $Y2=0
cc_881 N_A_1545_332#_c_1275_n N_A_1307_428#_c_1440_n 0.013007f $X=8.055 $Y=2.415
+ $X2=0 $Y2=0
cc_882 N_A_1545_332#_M1005_g N_A_1307_428#_c_1441_n 0.0115394f $X=7.81 $Y=0.7
+ $X2=0 $Y2=0
cc_883 N_A_1545_332#_c_1272_n N_A_1307_428#_c_1441_n 0.0207373f $X=7.89 $Y=1.825
+ $X2=0 $Y2=0
cc_884 N_A_1545_332#_c_1273_n N_A_1307_428#_c_1441_n 0.00154825f $X=7.89
+ $Y=1.825 $X2=0 $Y2=0
cc_885 N_A_1545_332#_c_1263_n N_A_1307_428#_c_1441_n 0.00103862f $X=9.4 $Y=2.145
+ $X2=0 $Y2=0
cc_886 N_A_1545_332#_c_1265_n N_A_1307_428#_c_1441_n 0.0115854f $X=9.4 $Y=1.29
+ $X2=0 $Y2=0
cc_887 N_A_1545_332#_c_1263_n N_A_1307_428#_c_1442_n 0.00577504f $X=9.4 $Y=2.145
+ $X2=0 $Y2=0
cc_888 N_A_1545_332#_c_1277_n N_A_1307_428#_c_1444_n 0.010159f $X=9.315 $Y=2.26
+ $X2=0 $Y2=0
cc_889 N_A_1545_332#_c_1263_n N_A_1307_428#_c_1444_n 0.0240502f $X=9.4 $Y=2.145
+ $X2=0 $Y2=0
cc_890 N_A_1545_332#_c_1281_n N_A_1307_428#_c_1444_n 0.0203521f $X=8.825 $Y=2.31
+ $X2=0 $Y2=0
cc_891 N_A_1545_332#_c_1265_n N_A_1307_428#_c_1444_n 0.00341162f $X=9.4 $Y=1.29
+ $X2=0 $Y2=0
cc_892 N_A_1545_332#_c_1277_n N_A_1307_428#_c_1445_n 4.48803e-19 $X=9.315
+ $Y=2.26 $X2=0 $Y2=0
cc_893 N_A_1545_332#_c_1263_n N_A_1307_428#_c_1445_n 0.00100302f $X=9.4 $Y=2.145
+ $X2=0 $Y2=0
cc_894 N_A_1545_332#_c_1281_n N_A_1307_428#_c_1445_n 0.00429421f $X=8.825
+ $Y=2.31 $X2=0 $Y2=0
cc_895 N_A_1545_332#_c_1265_n N_A_1307_428#_c_1445_n 0.00111671f $X=9.4 $Y=1.29
+ $X2=0 $Y2=0
cc_896 N_A_1545_332#_M1027_g N_RESET_B_M1025_g 0.0293818f $X=10.955 $Y=2.345
+ $X2=0 $Y2=0
cc_897 N_A_1545_332#_c_1279_n N_RESET_B_M1025_g 0.0203764f $X=10.735 $Y=2.29
+ $X2=0 $Y2=0
cc_898 N_A_1545_332#_c_1264_n N_RESET_B_M1025_g 0.00982587f $X=10.82 $Y=2.205
+ $X2=0 $Y2=0
cc_899 N_A_1545_332#_c_1266_n RESET_B 0.024833f $X=10.93 $Y=1.35 $X2=0 $Y2=0
cc_900 N_A_1545_332#_c_1267_n RESET_B 3.86988e-19 $X=10.93 $Y=1.26 $X2=0 $Y2=0
cc_901 N_A_1545_332#_c_1266_n N_RESET_B_c_1560_n 0.00112541f $X=10.93 $Y=1.35
+ $X2=0 $Y2=0
cc_902 N_A_1545_332#_c_1267_n N_RESET_B_c_1560_n 0.0208524f $X=10.93 $Y=1.26
+ $X2=0 $Y2=0
cc_903 N_A_1545_332#_c_1268_n N_RESET_B_c_1561_n 0.0133137f $X=10.93 $Y=1.185
+ $X2=0 $Y2=0
cc_904 N_A_1545_332#_c_1260_n N_A_2317_367#_M1039_g 0.0154614f $X=11.945
+ $Y=1.185 $X2=0 $Y2=0
cc_905 N_A_1545_332#_M1022_g N_A_2317_367#_M1024_g 0.0167559f $X=11.945 $Y=2.155
+ $X2=0 $Y2=0
cc_906 N_A_1545_332#_c_1260_n N_A_2317_367#_c_1592_n 0.00864467f $X=11.945
+ $Y=1.185 $X2=0 $Y2=0
cc_907 N_A_1545_332#_c_1268_n N_A_2317_367#_c_1592_n 8.38288e-19 $X=10.93
+ $Y=1.185 $X2=0 $Y2=0
cc_908 N_A_1545_332#_M1027_g N_A_2317_367#_c_1600_n 0.00160847f $X=10.955
+ $Y=2.345 $X2=0 $Y2=0
cc_909 N_A_1545_332#_M1022_g N_A_2317_367#_c_1600_n 0.0151894f $X=11.945
+ $Y=2.155 $X2=0 $Y2=0
cc_910 N_A_1545_332#_c_1260_n N_A_2317_367#_c_1593_n 0.00688256f $X=11.945
+ $Y=1.185 $X2=0 $Y2=0
cc_911 N_A_1545_332#_c_1262_n N_A_2317_367#_c_1593_n 0.00388801f $X=11.945
+ $Y=1.26 $X2=0 $Y2=0
cc_912 N_A_1545_332#_c_1259_n N_A_2317_367#_c_1594_n 0.00820827f $X=11.87
+ $Y=1.26 $X2=0 $Y2=0
cc_913 N_A_1545_332#_c_1260_n N_A_2317_367#_c_1594_n 0.00146351f $X=11.945
+ $Y=1.185 $X2=0 $Y2=0
cc_914 N_A_1545_332#_c_1262_n N_A_2317_367#_c_1594_n 5.27884e-19 $X=11.945
+ $Y=1.26 $X2=0 $Y2=0
cc_915 N_A_1545_332#_M1022_g N_A_2317_367#_c_1595_n 0.0104731f $X=11.945
+ $Y=2.155 $X2=0 $Y2=0
cc_916 N_A_1545_332#_c_1259_n N_A_2317_367#_c_1596_n 0.00541284f $X=11.87
+ $Y=1.26 $X2=0 $Y2=0
cc_917 N_A_1545_332#_M1022_g N_A_2317_367#_c_1596_n 0.0039104f $X=11.945
+ $Y=2.155 $X2=0 $Y2=0
cc_918 N_A_1545_332#_c_1262_n N_A_2317_367#_c_1597_n 0.00198978f $X=11.945
+ $Y=1.26 $X2=0 $Y2=0
cc_919 N_A_1545_332#_c_1262_n N_A_2317_367#_c_1598_n 0.0209917f $X=11.945
+ $Y=1.26 $X2=0 $Y2=0
cc_920 N_A_1545_332#_c_1274_n N_VPWR_M1036_d 0.00587974f $X=8.74 $Y=2.415 $X2=0
+ $Y2=0
cc_921 N_A_1545_332#_c_1279_n N_VPWR_M1001_d 0.00629221f $X=10.735 $Y=2.29 $X2=0
+ $Y2=0
cc_922 N_A_1545_332#_c_1279_n N_VPWR_M1025_d 0.00849026f $X=10.735 $Y=2.29 $X2=0
+ $Y2=0
cc_923 N_A_1545_332#_c_1264_n N_VPWR_M1025_d 0.0056513f $X=10.82 $Y=2.205 $X2=0
+ $Y2=0
cc_924 N_A_1545_332#_M1036_g N_VPWR_c_1657_n 0.00910848f $X=7.81 $Y=2.77 $X2=0
+ $Y2=0
cc_925 N_A_1545_332#_c_1274_n N_VPWR_c_1657_n 0.0196305f $X=8.74 $Y=2.415 $X2=0
+ $Y2=0
cc_926 N_A_1545_332#_c_1276_n N_VPWR_c_1657_n 0.0176165f $X=8.825 $Y=2.845 $X2=0
+ $Y2=0
cc_927 N_A_1545_332#_c_1276_n N_VPWR_c_1658_n 0.0136293f $X=8.825 $Y=2.845 $X2=0
+ $Y2=0
cc_928 N_A_1545_332#_c_1279_n N_VPWR_c_1658_n 0.0210602f $X=10.735 $Y=2.29 $X2=0
+ $Y2=0
cc_929 N_A_1545_332#_M1027_g N_VPWR_c_1659_n 0.0132198f $X=10.955 $Y=2.345 $X2=0
+ $Y2=0
cc_930 N_A_1545_332#_c_1279_n N_VPWR_c_1659_n 0.021916f $X=10.735 $Y=2.29 $X2=0
+ $Y2=0
cc_931 N_A_1545_332#_M1022_g N_VPWR_c_1660_n 0.00526768f $X=11.945 $Y=2.155
+ $X2=0 $Y2=0
cc_932 N_A_1545_332#_c_1276_n N_VPWR_c_1665_n 0.0124998f $X=8.825 $Y=2.845 $X2=0
+ $Y2=0
cc_933 N_A_1545_332#_M1036_g N_VPWR_c_1668_n 0.00478016f $X=7.81 $Y=2.77 $X2=0
+ $Y2=0
cc_934 N_A_1545_332#_M1027_g N_VPWR_c_1670_n 0.00393414f $X=10.955 $Y=2.345
+ $X2=0 $Y2=0
cc_935 N_A_1545_332#_M1022_g N_VPWR_c_1670_n 0.00312414f $X=11.945 $Y=2.155
+ $X2=0 $Y2=0
cc_936 N_A_1545_332#_M1036_g N_VPWR_c_1651_n 0.00611078f $X=7.81 $Y=2.77 $X2=0
+ $Y2=0
cc_937 N_A_1545_332#_M1027_g N_VPWR_c_1651_n 0.00787963f $X=10.955 $Y=2.345
+ $X2=0 $Y2=0
cc_938 N_A_1545_332#_M1022_g N_VPWR_c_1651_n 0.00410284f $X=11.945 $Y=2.155
+ $X2=0 $Y2=0
cc_939 N_A_1545_332#_c_1274_n N_VPWR_c_1651_n 0.0125941f $X=8.74 $Y=2.415 $X2=0
+ $Y2=0
cc_940 N_A_1545_332#_c_1275_n N_VPWR_c_1651_n 0.0105924f $X=8.055 $Y=2.415 $X2=0
+ $Y2=0
cc_941 N_A_1545_332#_c_1276_n N_VPWR_c_1651_n 0.00920722f $X=8.825 $Y=2.845
+ $X2=0 $Y2=0
cc_942 N_A_1545_332#_c_1277_n A_1823_430# 0.00561991f $X=9.315 $Y=2.26 $X2=-0.19
+ $Y2=-0.245
cc_943 N_A_1545_332#_c_1260_n N_Q_N_c_1865_n 0.00348491f $X=11.945 $Y=1.185
+ $X2=0 $Y2=0
cc_944 N_A_1545_332#_c_1268_n N_Q_N_c_1865_n 0.00622098f $X=10.93 $Y=1.185 $X2=0
+ $Y2=0
cc_945 N_A_1545_332#_c_1259_n N_Q_N_c_1866_n 0.00609999f $X=11.87 $Y=1.26 $X2=0
+ $Y2=0
cc_946 N_A_1545_332#_c_1266_n N_Q_N_c_1866_n 0.00407834f $X=10.93 $Y=1.35 $X2=0
+ $Y2=0
cc_947 N_A_1545_332#_c_1268_n N_Q_N_c_1866_n 0.00260315f $X=10.93 $Y=1.185 $X2=0
+ $Y2=0
cc_948 N_A_1545_332#_M1027_g N_Q_N_c_1868_n 0.00453786f $X=10.955 $Y=2.345 $X2=0
+ $Y2=0
cc_949 N_A_1545_332#_c_1259_n N_Q_N_c_1868_n 0.00620508f $X=11.87 $Y=1.26 $X2=0
+ $Y2=0
cc_950 N_A_1545_332#_c_1264_n N_Q_N_c_1868_n 0.0172466f $X=10.82 $Y=2.205 $X2=0
+ $Y2=0
cc_951 N_A_1545_332#_c_1266_n N_Q_N_c_1868_n 7.27024e-19 $X=10.93 $Y=1.35 $X2=0
+ $Y2=0
cc_952 N_A_1545_332#_c_1267_n N_Q_N_c_1868_n 2.43744e-19 $X=10.93 $Y=1.26 $X2=0
+ $Y2=0
cc_953 N_A_1545_332#_M1027_g N_Q_N_c_1867_n 0.00250731f $X=10.955 $Y=2.345 $X2=0
+ $Y2=0
cc_954 N_A_1545_332#_c_1259_n N_Q_N_c_1867_n 0.0161478f $X=11.87 $Y=1.26 $X2=0
+ $Y2=0
cc_955 N_A_1545_332#_M1022_g N_Q_N_c_1867_n 0.00632993f $X=11.945 $Y=2.155 $X2=0
+ $Y2=0
cc_956 N_A_1545_332#_c_1264_n N_Q_N_c_1867_n 0.00519375f $X=10.82 $Y=2.205 $X2=0
+ $Y2=0
cc_957 N_A_1545_332#_c_1266_n N_Q_N_c_1867_n 0.0233178f $X=10.93 $Y=1.35 $X2=0
+ $Y2=0
cc_958 N_A_1545_332#_c_1267_n N_Q_N_c_1867_n 0.00124625f $X=10.93 $Y=1.26 $X2=0
+ $Y2=0
cc_959 N_A_1545_332#_c_1268_n N_Q_N_c_1867_n 0.00411273f $X=10.93 $Y=1.185 $X2=0
+ $Y2=0
cc_960 N_A_1545_332#_M1022_g Q_N 0.00198823f $X=11.945 $Y=2.155 $X2=0 $Y2=0
cc_961 N_A_1545_332#_c_1260_n N_Q_c_1902_n 5.92037e-19 $X=11.945 $Y=1.185 $X2=0
+ $Y2=0
cc_962 N_A_1545_332#_M1005_g N_VGND_c_1933_n 0.00339422f $X=7.81 $Y=0.7 $X2=0
+ $Y2=0
cc_963 N_A_1545_332#_c_1266_n N_VGND_c_1934_n 0.00735348f $X=10.93 $Y=1.35 $X2=0
+ $Y2=0
cc_964 N_A_1545_332#_c_1267_n N_VGND_c_1934_n 0.00147662f $X=10.93 $Y=1.26 $X2=0
+ $Y2=0
cc_965 N_A_1545_332#_c_1268_n N_VGND_c_1934_n 0.00483983f $X=10.93 $Y=1.185
+ $X2=0 $Y2=0
cc_966 N_A_1545_332#_c_1260_n N_VGND_c_1935_n 0.00321894f $X=11.945 $Y=1.185
+ $X2=0 $Y2=0
cc_967 N_A_1545_332#_M1005_g N_VGND_c_1940_n 0.00213742f $X=7.81 $Y=0.7 $X2=0
+ $Y2=0
cc_968 N_A_1545_332#_c_1260_n N_VGND_c_1944_n 0.00385415f $X=11.945 $Y=1.185
+ $X2=0 $Y2=0
cc_969 N_A_1545_332#_c_1268_n N_VGND_c_1944_n 0.00549284f $X=10.93 $Y=1.185
+ $X2=0 $Y2=0
cc_970 N_A_1545_332#_M1005_g N_VGND_c_1946_n 0.0016946f $X=7.81 $Y=0.7 $X2=0
+ $Y2=0
cc_971 N_A_1545_332#_c_1260_n N_VGND_c_1946_n 0.0046122f $X=11.945 $Y=1.185
+ $X2=0 $Y2=0
cc_972 N_A_1545_332#_c_1268_n N_VGND_c_1946_n 0.0123926f $X=10.93 $Y=1.185 $X2=0
+ $Y2=0
cc_973 N_A_1545_332#_M1029_d N_A_1705_54#_c_2105_n 0.00492093f $X=8.955 $Y=0.27
+ $X2=0 $Y2=0
cc_974 N_A_1307_428#_M1038_g N_VPWR_c_1657_n 7.13137e-19 $X=9.04 $Y=2.57 $X2=0
+ $Y2=0
cc_975 N_A_1307_428#_c_1453_n N_VPWR_c_1657_n 0.00243483f $X=7.415 $Y=2.665
+ $X2=0 $Y2=0
cc_976 N_A_1307_428#_M1038_g N_VPWR_c_1658_n 0.00196142f $X=9.04 $Y=2.57 $X2=0
+ $Y2=0
cc_977 N_A_1307_428#_M1038_g N_VPWR_c_1665_n 0.00457319f $X=9.04 $Y=2.57 $X2=0
+ $Y2=0
cc_978 N_A_1307_428#_c_1453_n N_VPWR_c_1668_n 0.0118615f $X=7.415 $Y=2.665 $X2=0
+ $Y2=0
cc_979 N_A_1307_428#_c_1448_n N_VPWR_c_1668_n 0.0152961f $X=6.805 $Y=2.665 $X2=0
+ $Y2=0
cc_980 N_A_1307_428#_M1038_g N_VPWR_c_1651_n 0.00880519f $X=9.04 $Y=2.57 $X2=0
+ $Y2=0
cc_981 N_A_1307_428#_c_1453_n N_VPWR_c_1651_n 0.0179941f $X=7.415 $Y=2.665 $X2=0
+ $Y2=0
cc_982 N_A_1307_428#_c_1448_n N_VPWR_c_1651_n 0.0119585f $X=6.805 $Y=2.665 $X2=0
+ $Y2=0
cc_983 N_A_1307_428#_c_1453_n A_1419_512# 0.0157389f $X=7.415 $Y=2.665 $X2=-0.19
+ $Y2=-0.245
cc_984 N_A_1307_428#_c_1440_n A_1419_512# 6.42998e-19 $X=7.5 $Y=2.58 $X2=-0.19
+ $Y2=-0.245
cc_985 N_A_1307_428#_M1029_g N_VGND_c_1943_n 0.00337062f $X=8.88 $Y=0.59 $X2=0
+ $Y2=0
cc_986 N_A_1307_428#_M1029_g N_VGND_c_1946_n 0.00533431f $X=8.88 $Y=0.59 $X2=0
+ $Y2=0
cc_987 N_A_1307_428#_M1029_g N_A_1705_54#_c_2105_n 0.0132372f $X=8.88 $Y=0.59
+ $X2=0 $Y2=0
cc_988 N_RESET_B_M1025_g N_VPWR_c_1651_n 0.0038268f $X=10.445 $Y=2.035 $X2=0
+ $Y2=0
cc_989 N_RESET_B_c_1561_n N_VGND_c_1934_n 0.00490854f $X=10.385 $Y=1.185 $X2=0
+ $Y2=0
cc_990 N_RESET_B_c_1561_n N_VGND_c_1943_n 0.00384813f $X=10.385 $Y=1.185 $X2=0
+ $Y2=0
cc_991 N_RESET_B_c_1561_n N_VGND_c_1946_n 0.0046122f $X=10.385 $Y=1.185 $X2=0
+ $Y2=0
cc_992 N_RESET_B_c_1561_n N_A_1705_54#_c_2105_n 0.00194668f $X=10.385 $Y=1.185
+ $X2=0 $Y2=0
cc_993 N_A_2317_367#_M1024_g N_VPWR_c_1660_n 0.00698192f $X=12.455 $Y=2.465
+ $X2=0 $Y2=0
cc_994 N_A_2317_367#_c_1600_n N_VPWR_c_1660_n 0.0248129f $X=11.73 $Y=1.98 $X2=0
+ $Y2=0
cc_995 N_A_2317_367#_c_1595_n N_VPWR_c_1660_n 0.00637101f $X=12.155 $Y=1.55
+ $X2=0 $Y2=0
cc_996 N_A_2317_367#_c_1597_n N_VPWR_c_1660_n 0.0144853f $X=12.395 $Y=1.47 $X2=0
+ $Y2=0
cc_997 N_A_2317_367#_c_1598_n N_VPWR_c_1660_n 7.38452e-19 $X=12.395 $Y=1.47
+ $X2=0 $Y2=0
cc_998 N_A_2317_367#_M1024_g N_VPWR_c_1671_n 0.00549284f $X=12.455 $Y=2.465
+ $X2=0 $Y2=0
cc_999 N_A_2317_367#_M1024_g N_VPWR_c_1651_n 0.0120527f $X=12.455 $Y=2.465 $X2=0
+ $Y2=0
cc_1000 N_A_2317_367#_c_1600_n N_VPWR_c_1651_n 0.00972751f $X=11.73 $Y=1.98
+ $X2=0 $Y2=0
cc_1001 N_A_2317_367#_c_1592_n N_Q_N_c_1865_n 0.0347646f $X=11.73 $Y=0.865 $X2=0
+ $Y2=0
cc_1002 N_A_2317_367#_c_1600_n N_Q_N_c_1867_n 0.0620686f $X=11.73 $Y=1.98 $X2=0
+ $Y2=0
cc_1003 N_A_2317_367#_c_1594_n N_Q_N_c_1867_n 0.0119545f $X=11.895 $Y=1.2 $X2=0
+ $Y2=0
cc_1004 N_A_2317_367#_c_1596_n N_Q_N_c_1867_n 0.0128012f $X=11.895 $Y=1.55 $X2=0
+ $Y2=0
cc_1005 N_A_2317_367#_M1024_g N_Q_c_1904_n 0.0144925f $X=12.455 $Y=2.465 $X2=0
+ $Y2=0
cc_1006 N_A_2317_367#_M1024_g N_Q_c_1905_n 0.0030281f $X=12.455 $Y=2.465 $X2=0
+ $Y2=0
cc_1007 N_A_2317_367#_c_1597_n N_Q_c_1905_n 0.00107246f $X=12.395 $Y=1.47 $X2=0
+ $Y2=0
cc_1008 N_A_2317_367#_c_1598_n N_Q_c_1905_n 0.00131892f $X=12.395 $Y=1.47 $X2=0
+ $Y2=0
cc_1009 N_A_2317_367#_M1039_g N_Q_c_1901_n 0.00339687f $X=12.455 $Y=0.655 $X2=0
+ $Y2=0
cc_1010 N_A_2317_367#_M1024_g N_Q_c_1901_n 0.00443387f $X=12.455 $Y=2.465 $X2=0
+ $Y2=0
cc_1011 N_A_2317_367#_c_1597_n N_Q_c_1901_n 0.0327221f $X=12.395 $Y=1.47 $X2=0
+ $Y2=0
cc_1012 N_A_2317_367#_c_1598_n N_Q_c_1901_n 0.00770157f $X=12.395 $Y=1.47 $X2=0
+ $Y2=0
cc_1013 N_A_2317_367#_M1039_g N_Q_c_1902_n 0.00938329f $X=12.455 $Y=0.655 $X2=0
+ $Y2=0
cc_1014 N_A_2317_367#_M1039_g Q 0.00443358f $X=12.455 $Y=0.655 $X2=0 $Y2=0
cc_1015 N_A_2317_367#_c_1592_n Q 0.00411089f $X=11.73 $Y=0.865 $X2=0 $Y2=0
cc_1016 N_A_2317_367#_c_1597_n Q 9.46903e-19 $X=12.395 $Y=1.47 $X2=0 $Y2=0
cc_1017 N_A_2317_367#_c_1598_n Q 0.00127702f $X=12.395 $Y=1.47 $X2=0 $Y2=0
cc_1018 N_A_2317_367#_M1039_g N_VGND_c_1935_n 0.00449979f $X=12.455 $Y=0.655
+ $X2=0 $Y2=0
cc_1019 N_A_2317_367#_c_1592_n N_VGND_c_1935_n 0.0110325f $X=11.73 $Y=0.865
+ $X2=0 $Y2=0
cc_1020 N_A_2317_367#_c_1593_n N_VGND_c_1935_n 0.00618613f $X=12.155 $Y=1.2
+ $X2=0 $Y2=0
cc_1021 N_A_2317_367#_c_1597_n N_VGND_c_1935_n 0.0145552f $X=12.395 $Y=1.47
+ $X2=0 $Y2=0
cc_1022 N_A_2317_367#_c_1598_n N_VGND_c_1935_n 4.77677e-19 $X=12.395 $Y=1.47
+ $X2=0 $Y2=0
cc_1023 N_A_2317_367#_c_1592_n N_VGND_c_1944_n 0.00494947f $X=11.73 $Y=0.865
+ $X2=0 $Y2=0
cc_1024 N_A_2317_367#_M1039_g N_VGND_c_1945_n 0.00549284f $X=12.455 $Y=0.655
+ $X2=0 $Y2=0
cc_1025 N_A_2317_367#_M1039_g N_VGND_c_1946_n 0.0120527f $X=12.455 $Y=0.655
+ $X2=0 $Y2=0
cc_1026 N_A_2317_367#_c_1592_n N_VGND_c_1946_n 0.00748098f $X=11.73 $Y=0.865
+ $X2=0 $Y2=0
cc_1027 N_VPWR_c_1667_n N_A_531_47#_c_1796_n 0.00729809f $X=4.265 $Y=3.33 $X2=0
+ $Y2=0
cc_1028 N_VPWR_c_1651_n N_A_531_47#_c_1796_n 0.00892727f $X=12.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1029 N_VPWR_c_1659_n Q_N 0.0165395f $X=10.74 $Y=2.775 $X2=0 $Y2=0
cc_1030 N_VPWR_c_1660_n Q_N 0.0164451f $X=12.24 $Y=1.98 $X2=0 $Y2=0
cc_1031 N_VPWR_c_1670_n Q_N 0.0169956f $X=12.075 $Y=3.33 $X2=0 $Y2=0
cc_1032 N_VPWR_c_1651_n Q_N 0.0133402f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_1033 N_VPWR_c_1651_n N_Q_M1024_d 0.0023218f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_1034 N_VPWR_c_1671_n N_Q_c_1904_n 0.0221179f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_1035 N_VPWR_c_1651_n N_Q_c_1904_n 0.0138623f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_1036 N_VPWR_c_1660_n N_Q_c_1905_n 0.0461898f $X=12.24 $Y=1.98 $X2=0 $Y2=0
cc_1037 N_A_531_47#_c_1799_n N_VGND_c_1930_n 0.0101653f $X=2.795 $Y=0.47 $X2=0
+ $Y2=0
cc_1038 N_A_531_47#_c_1799_n N_VGND_c_1942_n 0.0178561f $X=2.795 $Y=0.47 $X2=0
+ $Y2=0
cc_1039 N_A_531_47#_M1002_d N_VGND_c_1946_n 0.0022543f $X=2.655 $Y=0.235 $X2=0
+ $Y2=0
cc_1040 N_A_531_47#_c_1799_n N_VGND_c_1946_n 0.0124703f $X=2.795 $Y=0.47 $X2=0
+ $Y2=0
cc_1041 N_A_531_47#_c_1793_n N_VGND_c_1946_n 0.00542338f $X=3.18 $Y=0.915 $X2=0
+ $Y2=0
cc_1042 N_Q_N_c_1865_n N_VGND_c_1935_n 0.0123407f $X=11.175 $Y=0.43 $X2=0 $Y2=0
cc_1043 N_Q_N_c_1865_n N_VGND_c_1944_n 0.0268376f $X=11.175 $Y=0.43 $X2=0 $Y2=0
cc_1044 N_Q_N_M1037_d N_VGND_c_1946_n 0.0023218f $X=11.035 $Y=0.235 $X2=0 $Y2=0
cc_1045 N_Q_N_c_1865_n N_VGND_c_1946_n 0.0165708f $X=11.175 $Y=0.43 $X2=0 $Y2=0
cc_1046 N_Q_c_1902_n N_VGND_c_1945_n 0.0221179f $X=12.67 $Y=0.43 $X2=0 $Y2=0
cc_1047 N_Q_M1039_d N_VGND_c_1946_n 0.0023218f $X=12.53 $Y=0.235 $X2=0 $Y2=0
cc_1048 N_Q_c_1902_n N_VGND_c_1946_n 0.0138623f $X=12.67 $Y=0.43 $X2=0 $Y2=0
cc_1049 N_VGND_c_1946_n A_719_47# 0.00678611f $X=12.72 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1050 N_VGND_c_1946_n N_A_917_47#_M1003_d 0.0022543f $X=12.72 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1051 N_VGND_c_1946_n N_A_917_47#_M1019_d 0.00232217f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_1052 N_VGND_c_1938_n N_A_917_47#_c_2080_n 0.0178736f $X=6.14 $Y=0 $X2=0 $Y2=0
cc_1053 N_VGND_c_1946_n N_A_917_47#_c_2080_n 0.0125011f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_1054 N_VGND_c_1932_n N_A_917_47#_c_2076_n 0.0177521f $X=6.305 $Y=0.415 $X2=0
+ $Y2=0
cc_1055 N_VGND_c_1938_n N_A_917_47#_c_2077_n 0.0562164f $X=6.14 $Y=0 $X2=0 $Y2=0
cc_1056 N_VGND_c_1946_n N_A_917_47#_c_2077_n 0.0369028f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_1057 N_VGND_c_1933_n N_A_1705_54#_c_2105_n 0.0133095f $X=8.155 $Y=0.505 $X2=0
+ $Y2=0
cc_1058 N_VGND_c_1943_n N_A_1705_54#_c_2105_n 0.0844231f $X=10.58 $Y=0 $X2=0
+ $Y2=0
cc_1059 N_VGND_c_1946_n N_A_1705_54#_c_2105_n 0.0495512f $X=12.72 $Y=0 $X2=0
+ $Y2=0
