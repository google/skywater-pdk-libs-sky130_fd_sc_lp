* File: sky130_fd_sc_lp__a32oi_lp.pxi.spice
* Created: Wed Sep  2 09:28:34 2020
* 
x_PM_SKY130_FD_SC_LP__A32OI_LP%B2 N_B2_M1008_g N_B2_c_68_n N_B2_M1005_g
+ N_B2_c_69_n B2 B2 N_B2_c_71_n PM_SKY130_FD_SC_LP__A32OI_LP%B2
x_PM_SKY130_FD_SC_LP__A32OI_LP%B1 N_B1_c_106_n N_B1_M1006_g N_B1_M1000_g
+ N_B1_c_107_n N_B1_c_108_n N_B1_c_109_n N_B1_c_110_n B1 B1 N_B1_c_112_n
+ PM_SKY130_FD_SC_LP__A32OI_LP%B1
x_PM_SKY130_FD_SC_LP__A32OI_LP%A1 N_A1_M1007_g N_A1_M1001_g N_A1_c_166_n
+ N_A1_c_167_n N_A1_c_168_n A1 A1 A1 A1 N_A1_c_170_n
+ PM_SKY130_FD_SC_LP__A32OI_LP%A1
x_PM_SKY130_FD_SC_LP__A32OI_LP%A2 N_A2_M1002_g N_A2_M1004_g A2 N_A2_c_221_n
+ PM_SKY130_FD_SC_LP__A32OI_LP%A2
x_PM_SKY130_FD_SC_LP__A32OI_LP%A3 N_A3_M1003_g N_A3_M1009_g A3 A3 N_A3_c_256_n
+ PM_SKY130_FD_SC_LP__A32OI_LP%A3
x_PM_SKY130_FD_SC_LP__A32OI_LP%A_56_409# N_A_56_409#_M1005_s N_A_56_409#_M1000_d
+ N_A_56_409#_M1002_d N_A_56_409#_c_279_n N_A_56_409#_c_280_n
+ N_A_56_409#_c_281_n N_A_56_409#_c_282_n N_A_56_409#_c_289_n
+ N_A_56_409#_c_283_n N_A_56_409#_c_284_n N_A_56_409#_c_285_n
+ PM_SKY130_FD_SC_LP__A32OI_LP%A_56_409#
x_PM_SKY130_FD_SC_LP__A32OI_LP%Y N_Y_M1006_d N_Y_M1005_d N_Y_c_336_n N_Y_c_340_n
+ N_Y_c_341_n N_Y_c_349_n N_Y_c_337_n Y Y Y N_Y_c_339_n
+ PM_SKY130_FD_SC_LP__A32OI_LP%Y
x_PM_SKY130_FD_SC_LP__A32OI_LP%VPWR N_VPWR_M1007_d N_VPWR_M1009_d N_VPWR_c_391_n
+ N_VPWR_c_392_n N_VPWR_c_393_n N_VPWR_c_394_n N_VPWR_c_395_n VPWR
+ N_VPWR_c_396_n N_VPWR_c_390_n PM_SKY130_FD_SC_LP__A32OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A32OI_LP%VGND N_VGND_M1008_s N_VGND_M1003_d N_VGND_c_428_n
+ N_VGND_c_429_n N_VGND_c_430_n N_VGND_c_431_n N_VGND_c_432_n VGND
+ N_VGND_c_433_n N_VGND_c_434_n PM_SKY130_FD_SC_LP__A32OI_LP%VGND
cc_1 VNB N_B2_M1008_g 0.0420309f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.445
cc_2 VNB N_B2_c_68_n 0.00227792f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.79
cc_3 VNB N_B2_c_69_n 0.0256646f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.625
cc_4 VNB B2 0.00173674f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_B2_c_71_n 0.0176088f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_6 VNB N_B1_c_106_n 0.0156507f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.12
cc_7 VNB N_B1_c_107_n 0.016022f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_B1_c_108_n 0.0133579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_109_n 0.0232004f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_10 VNB N_B1_c_110_n 0.00276104f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_11 VNB B1 0.00171029f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_12 VNB N_B1_c_112_n 0.0164244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1007_g 0.0110861f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.445
cc_14 VNB N_A1_c_166_n 0.0180554f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_15 VNB N_A1_c_167_n 0.0226054f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.12
cc_16 VNB N_A1_c_168_n 0.012682f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.625
cc_17 VNB A1 0.0102711f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_18 VNB N_A1_c_170_n 0.0167019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_M1004_g 0.0534506f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.545
cc_20 VNB A2 0.00470379f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_21 VNB N_A2_c_221_n 0.0215f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_22 VNB N_A3_M1003_g 0.024692f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.445
cc_23 VNB N_A3_M1009_g 0.0481384f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.545
cc_24 VNB A3 0.0351865f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.12
cc_25 VNB N_A3_c_256_n 0.0353788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_336_n 0.0221972f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.545
cc_27 VNB N_Y_c_337_n 6.658e-19 $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_28 VNB Y 0.0367309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_339_n 0.0110226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_390_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_428_n 0.0147066f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.545
cc_32 VNB N_VGND_c_429_n 0.0158836f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_33 VNB N_VGND_c_430_n 0.0177827f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_34 VNB N_VGND_c_431_n 0.0580711f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_35 VNB N_VGND_c_432_n 0.00511011f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.285
cc_36 VNB N_VGND_c_433_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_434_n 0.194577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_B2_c_68_n 0.0124909f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.79
cc_39 VPB N_B2_M1005_g 0.0360101f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.545
cc_40 VPB B2 7.45984e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_41 VPB N_B1_M1000_g 0.0319548f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_B1_c_110_n 0.0108545f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.285
cc_43 VPB B1 7.50599e-19 $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.285
cc_44 VPB N_A1_M1007_g 0.0379571f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.445
cc_45 VPB A1 0.00263147f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_46 VPB N_A2_M1002_g 0.0315788f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.445
cc_47 VPB A2 0.0028409f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.285
cc_48 VPB N_A2_c_221_n 0.00918451f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_49 VPB N_A3_M1009_g 0.0528141f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.545
cc_50 VPB N_A_56_409#_c_279_n 0.0219771f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_51 VPB N_A_56_409#_c_280_n 0.00202865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_56_409#_c_281_n 0.00938685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_56_409#_c_282_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.285
cc_54 VPB N_A_56_409#_c_283_n 0.010195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_56_409#_c_284_n 0.00814719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_56_409#_c_285_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_340_n 0.0155937f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.285
cc_58 VPB N_Y_c_341_n 0.0137584f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.12
cc_59 VPB Y 0.016339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_391_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.285
cc_61 VPB N_VPWR_c_392_n 0.0108116f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.625
cc_62 VPB N_VPWR_c_393_n 0.0555303f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_63 VPB N_VPWR_c_394_n 0.0474858f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.285
cc_64 VPB N_VPWR_c_395_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.285
cc_65 VPB N_VPWR_c_396_n 0.0219685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_390_n 0.0619474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 N_B2_M1008_g N_B1_c_106_n 0.040928f $X=0.625 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_68 N_B2_c_68_n N_B1_M1000_g 5.52405e-19 $X=0.69 $Y=1.79 $X2=0 $Y2=0
cc_69 N_B2_M1005_g N_B1_M1000_g 0.0334594f $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_70 N_B2_M1008_g N_B1_c_108_n 0.00909334f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_71 N_B2_c_69_n N_B1_c_109_n 0.0133663f $X=0.69 $Y=1.625 $X2=0 $Y2=0
cc_72 N_B2_c_68_n N_B1_c_110_n 0.0133663f $X=0.69 $Y=1.79 $X2=0 $Y2=0
cc_73 B2 B1 0.0416998f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_B2_c_71_n B1 0.00229175f $X=0.69 $Y=1.285 $X2=0 $Y2=0
cc_75 B2 N_B1_c_112_n 0.00229175f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B2_c_71_n N_B1_c_112_n 0.0133663f $X=0.69 $Y=1.285 $X2=0 $Y2=0
cc_77 N_B2_M1005_g N_A_56_409#_c_279_n 0.0110936f $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_78 N_B2_M1005_g N_A_56_409#_c_280_n 0.0164696f $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_79 N_B2_M1005_g N_A_56_409#_c_281_n 9.65935e-19 $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_80 N_B2_M1005_g N_A_56_409#_c_289_n 7.1089e-19 $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_81 N_B2_M1008_g N_Y_c_336_n 0.0137253f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_82 B2 N_Y_c_336_n 0.0234911f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 N_B2_c_71_n N_Y_c_336_n 0.00120985f $X=0.69 $Y=1.285 $X2=0 $Y2=0
cc_84 N_B2_c_68_n N_Y_c_340_n 5.7132e-19 $X=0.69 $Y=1.79 $X2=0 $Y2=0
cc_85 N_B2_M1005_g N_Y_c_340_n 0.0211953f $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_86 B2 N_Y_c_340_n 0.0246384f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 N_B2_M1005_g N_Y_c_349_n 0.0152285f $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_88 N_B2_M1008_g N_Y_c_337_n 0.00177798f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_89 N_B2_M1008_g Y 0.00642454f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_90 N_B2_M1005_g Y 0.00634172f $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_91 B2 Y 0.0491281f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_92 N_B2_c_71_n Y 0.0149783f $X=0.69 $Y=1.285 $X2=0 $Y2=0
cc_93 N_B2_M1005_g N_VPWR_c_394_n 0.00546179f $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_94 N_B2_M1005_g N_VPWR_c_390_n 0.00813499f $X=0.69 $Y=2.545 $X2=0 $Y2=0
cc_95 N_B2_M1008_g N_VGND_c_429_n 0.0119757f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_96 N_B2_M1008_g N_VGND_c_431_n 0.00367954f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_97 N_B2_M1008_g N_VGND_c_434_n 0.0043701f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_98 N_B1_M1000_g N_A1_M1007_g 0.0202091f $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_99 N_B1_c_109_n N_A1_M1007_g 0.0191489f $X=1.23 $Y=1.615 $X2=0 $Y2=0
cc_100 B1 N_A1_M1007_g 3.9656e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B1_c_106_n N_A1_c_166_n 0.00792792f $X=1.015 $Y=0.73 $X2=0 $Y2=0
cc_102 N_B1_c_107_n N_A1_c_166_n 8.87692e-19 $X=1.14 $Y=0.805 $X2=0 $Y2=0
cc_103 N_B1_c_108_n N_A1_c_167_n 0.00478705f $X=1.23 $Y=1.11 $X2=0 $Y2=0
cc_104 B1 N_A1_c_167_n 3.82958e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B1_c_112_n N_A1_c_167_n 0.0101427f $X=1.23 $Y=1.275 $X2=0 $Y2=0
cc_106 N_B1_c_109_n N_A1_c_168_n 0.0101427f $X=1.23 $Y=1.615 $X2=0 $Y2=0
cc_107 N_B1_c_106_n A1 4.94388e-19 $X=1.015 $Y=0.73 $X2=0 $Y2=0
cc_108 N_B1_c_107_n A1 5.22018e-19 $X=1.14 $Y=0.805 $X2=0 $Y2=0
cc_109 N_B1_c_108_n A1 0.00359436f $X=1.23 $Y=1.11 $X2=0 $Y2=0
cc_110 B1 A1 0.0510783f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B1_c_112_n A1 0.00391221f $X=1.23 $Y=1.275 $X2=0 $Y2=0
cc_112 N_B1_c_107_n N_A1_c_170_n 0.00478705f $X=1.14 $Y=0.805 $X2=0 $Y2=0
cc_113 N_B1_M1000_g N_A_56_409#_c_279_n 7.1089e-19 $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_114 N_B1_M1000_g N_A_56_409#_c_280_n 0.0164696f $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_115 N_B1_M1000_g N_A_56_409#_c_282_n 8.05528e-19 $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_116 N_B1_M1000_g N_A_56_409#_c_289_n 0.0134077f $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_117 N_B1_M1000_g N_A_56_409#_c_284_n 0.00434405f $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_118 N_B1_c_110_n N_A_56_409#_c_284_n 3.80871e-19 $X=1.23 $Y=1.78 $X2=0 $Y2=0
cc_119 B1 N_A_56_409#_c_284_n 0.00619639f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B1_c_107_n N_Y_c_336_n 0.0106693f $X=1.14 $Y=0.805 $X2=0 $Y2=0
cc_121 N_B1_c_108_n N_Y_c_336_n 0.00412273f $X=1.23 $Y=1.11 $X2=0 $Y2=0
cc_122 B1 N_Y_c_336_n 0.027244f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_123 N_B1_c_112_n N_Y_c_336_n 0.00138018f $X=1.23 $Y=1.275 $X2=0 $Y2=0
cc_124 N_B1_M1000_g N_Y_c_340_n 0.00418961f $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_125 N_B1_c_110_n N_Y_c_340_n 2.23711e-19 $X=1.23 $Y=1.78 $X2=0 $Y2=0
cc_126 B1 N_Y_c_340_n 0.00430536f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B1_M1000_g N_Y_c_349_n 0.00995048f $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_128 N_B1_c_106_n N_Y_c_337_n 0.00934714f $X=1.015 $Y=0.73 $X2=0 $Y2=0
cc_129 N_B1_c_107_n N_Y_c_337_n 0.00394925f $X=1.14 $Y=0.805 $X2=0 $Y2=0
cc_130 N_B1_M1000_g N_VPWR_c_391_n 8.65588e-19 $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_131 N_B1_M1000_g N_VPWR_c_394_n 0.00546179f $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_132 N_B1_M1000_g N_VPWR_c_390_n 0.00742485f $X=1.22 $Y=2.545 $X2=0 $Y2=0
cc_133 N_B1_c_106_n N_VGND_c_429_n 0.00212811f $X=1.015 $Y=0.73 $X2=0 $Y2=0
cc_134 N_B1_c_106_n N_VGND_c_431_n 0.00430243f $X=1.015 $Y=0.73 $X2=0 $Y2=0
cc_135 N_B1_c_107_n N_VGND_c_431_n 2.88546e-19 $X=1.14 $Y=0.805 $X2=0 $Y2=0
cc_136 N_B1_c_106_n N_VGND_c_434_n 0.00666884f $X=1.015 $Y=0.73 $X2=0 $Y2=0
cc_137 N_A1_M1007_g N_A2_M1002_g 0.0318804f $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_138 N_A1_M1007_g N_A2_M1004_g 5.27058e-19 $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_139 N_A1_c_166_n N_A2_M1004_g 0.0205783f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_140 A1 N_A2_M1004_g 0.0113086f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_141 N_A1_c_170_n N_A2_M1004_g 0.0362806f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_142 N_A1_M1007_g A2 3.78364e-19 $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_143 A1 A2 0.0234319f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_144 N_A1_M1007_g N_A2_c_221_n 0.0156685f $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_145 A1 N_A2_c_221_n 0.0012155f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_146 A1 A3 0.0108459f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_147 N_A1_M1007_g N_A_56_409#_c_282_n 0.00335672f $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_148 N_A1_M1007_g N_A_56_409#_c_289_n 0.013408f $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_149 N_A1_M1007_g N_A_56_409#_c_283_n 0.0178513f $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_150 A1 N_A_56_409#_c_283_n 0.0211197f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_151 N_A1_M1007_g N_A_56_409#_c_284_n 0.00175233f $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_152 A1 N_A_56_409#_c_284_n 0.00642801f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_153 N_A1_M1007_g N_A_56_409#_c_285_n 9.22443e-19 $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_154 A1 N_Y_M1006_d 0.00212073f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_155 A1 N_Y_c_336_n 0.014528f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_156 N_A1_c_170_n N_Y_c_336_n 6.71456e-19 $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_157 N_A1_c_166_n N_Y_c_337_n 0.00535186f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_158 A1 N_Y_c_337_n 0.0250478f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_159 N_A1_M1007_g N_VPWR_c_391_n 0.0178519f $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_160 N_A1_M1007_g N_VPWR_c_394_n 0.00767656f $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_161 N_A1_M1007_g N_VPWR_c_390_n 0.0134103f $X=1.75 $Y=2.545 $X2=0 $Y2=0
cc_162 N_A1_c_166_n N_VGND_c_431_n 0.00393362f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_163 A1 N_VGND_c_431_n 0.00938196f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_164 N_A1_c_170_n N_VGND_c_431_n 4.68429e-19 $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_165 N_A1_c_166_n N_VGND_c_434_n 0.00646985f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_166 A1 N_VGND_c_434_n 0.0117206f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_167 A1 A_357_47# 0.00415398f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_168 N_A2_M1004_g N_A3_M1003_g 0.0549862f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A2_M1002_g N_A3_M1009_g 0.0201312f $X=2.28 $Y=2.545 $X2=0 $Y2=0
cc_170 N_A2_M1004_g N_A3_M1009_g 0.0130093f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_171 A2 N_A3_M1009_g 0.0237525f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_172 N_A2_c_221_n N_A3_M1009_g 0.0213979f $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_173 N_A2_M1004_g A3 0.00368567f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_174 A2 A3 0.011522f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_175 A2 N_A3_c_256_n 0.00290268f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A2_M1002_g N_A_56_409#_c_289_n 8.71905e-19 $X=2.28 $Y=2.545 $X2=0 $Y2=0
cc_177 N_A2_M1002_g N_A_56_409#_c_283_n 0.0196138f $X=2.28 $Y=2.545 $X2=0 $Y2=0
cc_178 A2 N_A_56_409#_c_283_n 0.0433404f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A2_c_221_n N_A_56_409#_c_283_n 0.00184542f $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_180 N_A2_M1002_g N_A_56_409#_c_285_n 0.016685f $X=2.28 $Y=2.545 $X2=0 $Y2=0
cc_181 N_A2_M1002_g N_VPWR_c_391_n 0.0178582f $X=2.28 $Y=2.545 $X2=0 $Y2=0
cc_182 N_A2_M1002_g N_VPWR_c_396_n 0.00769046f $X=2.28 $Y=2.545 $X2=0 $Y2=0
cc_183 N_A2_M1002_g N_VPWR_c_390_n 0.0134474f $X=2.28 $Y=2.545 $X2=0 $Y2=0
cc_184 N_A2_M1004_g N_VGND_c_430_n 0.00304577f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A2_M1004_g N_VGND_c_431_n 0.00585385f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A2_M1004_g N_VGND_c_434_n 0.0111877f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A3_M1009_g N_A_56_409#_c_283_n 0.00617417f $X=2.81 $Y=2.545 $X2=0 $Y2=0
cc_188 N_A3_M1009_g N_A_56_409#_c_285_n 0.0151466f $X=2.81 $Y=2.545 $X2=0 $Y2=0
cc_189 N_A3_M1009_g N_VPWR_c_391_n 8.6579e-19 $X=2.81 $Y=2.545 $X2=0 $Y2=0
cc_190 N_A3_M1009_g N_VPWR_c_393_n 0.00505795f $X=2.81 $Y=2.545 $X2=0 $Y2=0
cc_191 N_A3_M1009_g N_VPWR_c_396_n 0.0086001f $X=2.81 $Y=2.545 $X2=0 $Y2=0
cc_192 N_A3_M1009_g N_VPWR_c_390_n 0.0163182f $X=2.81 $Y=2.545 $X2=0 $Y2=0
cc_193 N_A3_M1003_g N_VGND_c_430_n 0.0135345f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_194 A3 N_VGND_c_430_n 0.0230834f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_195 N_A3_c_256_n N_VGND_c_430_n 0.00577783f $X=2.73 $Y=0.975 $X2=0 $Y2=0
cc_196 N_A3_M1003_g N_VGND_c_431_n 0.00486043f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_197 N_A3_M1003_g N_VGND_c_434_n 0.00447521f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_198 A3 N_VGND_c_434_n 0.014566f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_199 N_A_56_409#_c_280_n N_Y_M1005_d 0.00180746f $X=1.32 $Y=2.98 $X2=0 $Y2=0
cc_200 N_A_56_409#_M1005_s N_Y_c_340_n 0.00196682f $X=0.28 $Y=2.045 $X2=0 $Y2=0
cc_201 N_A_56_409#_c_279_n N_Y_c_340_n 0.0143771f $X=0.425 $Y=2.485 $X2=0 $Y2=0
cc_202 N_A_56_409#_c_289_n N_Y_c_340_n 6.67284e-19 $X=1.485 $Y=2.19 $X2=0 $Y2=0
cc_203 N_A_56_409#_c_284_n N_Y_c_340_n 0.0118744f $X=1.65 $Y=2.045 $X2=0 $Y2=0
cc_204 N_A_56_409#_M1005_s N_Y_c_341_n 0.00107873f $X=0.28 $Y=2.045 $X2=0 $Y2=0
cc_205 N_A_56_409#_c_279_n N_Y_c_341_n 0.00732286f $X=0.425 $Y=2.485 $X2=0 $Y2=0
cc_206 N_A_56_409#_c_279_n N_Y_c_349_n 0.0260268f $X=0.425 $Y=2.485 $X2=0 $Y2=0
cc_207 N_A_56_409#_c_280_n N_Y_c_349_n 0.015238f $X=1.32 $Y=2.98 $X2=0 $Y2=0
cc_208 N_A_56_409#_c_289_n N_Y_c_349_n 0.0378542f $X=1.485 $Y=2.19 $X2=0 $Y2=0
cc_209 N_A_56_409#_c_283_n N_VPWR_M1007_d 0.00180746f $X=2.38 $Y=2.045 $X2=-0.19
+ $Y2=1.655
cc_210 N_A_56_409#_c_282_n N_VPWR_c_391_n 0.0119061f $X=1.485 $Y=2.895 $X2=0
+ $Y2=0
cc_211 N_A_56_409#_c_289_n N_VPWR_c_391_n 0.0385131f $X=1.485 $Y=2.19 $X2=0
+ $Y2=0
cc_212 N_A_56_409#_c_283_n N_VPWR_c_391_n 0.0163515f $X=2.38 $Y=2.045 $X2=0
+ $Y2=0
cc_213 N_A_56_409#_c_285_n N_VPWR_c_391_n 0.0497475f $X=2.545 $Y=2.19 $X2=0
+ $Y2=0
cc_214 N_A_56_409#_c_283_n N_VPWR_c_393_n 0.00349942f $X=2.38 $Y=2.045 $X2=0
+ $Y2=0
cc_215 N_A_56_409#_c_285_n N_VPWR_c_393_n 0.024056f $X=2.545 $Y=2.19 $X2=0 $Y2=0
cc_216 N_A_56_409#_c_280_n N_VPWR_c_394_n 0.0429254f $X=1.32 $Y=2.98 $X2=0 $Y2=0
cc_217 N_A_56_409#_c_281_n N_VPWR_c_394_n 0.0221635f $X=0.59 $Y=2.98 $X2=0 $Y2=0
cc_218 N_A_56_409#_c_282_n N_VPWR_c_394_n 0.0220769f $X=1.485 $Y=2.895 $X2=0
+ $Y2=0
cc_219 N_A_56_409#_c_285_n N_VPWR_c_396_n 0.021949f $X=2.545 $Y=2.19 $X2=0 $Y2=0
cc_220 N_A_56_409#_c_280_n N_VPWR_c_390_n 0.0252151f $X=1.32 $Y=2.98 $X2=0 $Y2=0
cc_221 N_A_56_409#_c_281_n N_VPWR_c_390_n 0.0126536f $X=0.59 $Y=2.98 $X2=0 $Y2=0
cc_222 N_A_56_409#_c_282_n N_VPWR_c_390_n 0.0125384f $X=1.485 $Y=2.895 $X2=0
+ $Y2=0
cc_223 N_A_56_409#_c_285_n N_VPWR_c_390_n 0.0124703f $X=2.545 $Y=2.19 $X2=0
+ $Y2=0
cc_224 N_Y_c_339_n N_VGND_c_428_n 0.00191638f $X=0.235 $Y=0.93 $X2=0 $Y2=0
cc_225 N_Y_c_336_n N_VGND_c_429_n 0.0148247f $X=1.065 $Y=0.845 $X2=0 $Y2=0
cc_226 N_Y_c_337_n N_VGND_c_429_n 0.00997941f $X=1.23 $Y=0.47 $X2=0 $Y2=0
cc_227 N_Y_c_339_n N_VGND_c_429_n 0.00840986f $X=0.235 $Y=0.93 $X2=0 $Y2=0
cc_228 N_Y_c_336_n N_VGND_c_431_n 0.00650557f $X=1.065 $Y=0.845 $X2=0 $Y2=0
cc_229 N_Y_c_337_n N_VGND_c_431_n 0.0197336f $X=1.23 $Y=0.47 $X2=0 $Y2=0
cc_230 N_Y_M1006_d N_VGND_c_434_n 0.0108431f $X=1.09 $Y=0.235 $X2=0 $Y2=0
cc_231 N_Y_c_336_n N_VGND_c_434_n 0.0123265f $X=1.065 $Y=0.845 $X2=0 $Y2=0
cc_232 N_Y_c_337_n N_VGND_c_434_n 0.0125731f $X=1.23 $Y=0.47 $X2=0 $Y2=0
cc_233 N_Y_c_339_n N_VGND_c_434_n 0.0037794f $X=0.235 $Y=0.93 $X2=0 $Y2=0
cc_234 N_VGND_c_434_n A_140_47# 0.00323414f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_235 N_VGND_c_434_n A_357_47# 0.0116489f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_236 N_VGND_c_434_n A_465_47# 0.00913486f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
