* File: sky130_fd_sc_lp__einvp_8.pxi.spice
* Created: Wed Sep  2 09:52:42 2020
* 
x_PM_SKY130_FD_SC_LP__EINVP_8%A_182_367# N_A_182_367#_M1027_d
+ N_A_182_367#_M1026_d N_A_182_367#_c_175_n N_A_182_367#_c_176_n
+ N_A_182_367#_c_194_n N_A_182_367#_M1000_g N_A_182_367#_c_177_n
+ N_A_182_367#_c_196_n N_A_182_367#_M1005_g N_A_182_367#_c_178_n
+ N_A_182_367#_c_198_n N_A_182_367#_M1007_g N_A_182_367#_c_179_n
+ N_A_182_367#_c_200_n N_A_182_367#_M1016_g N_A_182_367#_c_180_n
+ N_A_182_367#_c_202_n N_A_182_367#_M1019_g N_A_182_367#_c_181_n
+ N_A_182_367#_c_204_n N_A_182_367#_M1020_g N_A_182_367#_c_182_n
+ N_A_182_367#_c_206_n N_A_182_367#_M1021_g N_A_182_367#_c_183_n
+ N_A_182_367#_c_208_n N_A_182_367#_M1033_g N_A_182_367#_c_209_n
+ N_A_182_367#_c_210_n N_A_182_367#_c_184_n N_A_182_367#_c_185_n
+ N_A_182_367#_c_186_n N_A_182_367#_c_187_n N_A_182_367#_c_188_n
+ N_A_182_367#_c_189_n N_A_182_367#_c_190_n N_A_182_367#_c_218_n
+ N_A_182_367#_c_219_n N_A_182_367#_c_191_n N_A_182_367#_c_221_n
+ PM_SKY130_FD_SC_LP__EINVP_8%A_182_367#
x_PM_SKY130_FD_SC_LP__EINVP_8%TE N_TE_M1026_g N_TE_c_338_n N_TE_M1027_g
+ N_TE_c_339_n N_TE_c_340_n N_TE_c_341_n N_TE_M1001_g N_TE_c_342_n N_TE_c_343_n
+ N_TE_c_344_n N_TE_M1004_g N_TE_c_345_n N_TE_c_346_n N_TE_M1010_g N_TE_c_347_n
+ N_TE_c_348_n N_TE_M1014_g N_TE_c_349_n N_TE_c_350_n N_TE_M1017_g N_TE_c_351_n
+ N_TE_c_352_n N_TE_M1024_g N_TE_c_353_n N_TE_c_354_n N_TE_M1028_g N_TE_c_355_n
+ N_TE_c_356_n N_TE_M1030_g N_TE_c_357_n N_TE_c_358_n N_TE_c_359_n N_TE_c_360_n
+ N_TE_c_361_n N_TE_c_362_n N_TE_c_363_n TE TE PM_SKY130_FD_SC_LP__EINVP_8%TE
x_PM_SKY130_FD_SC_LP__EINVP_8%A N_A_M1003_g N_A_M1002_g N_A_M1006_g N_A_M1008_g
+ N_A_M1009_g N_A_M1011_g N_A_M1012_g N_A_M1015_g N_A_M1013_g N_A_M1022_g
+ N_A_M1018_g N_A_M1025_g N_A_M1023_g N_A_M1029_g N_A_M1032_g N_A_M1031_g
+ N_A_c_559_p N_A_c_493_n N_A_c_494_n A A N_A_c_495_n
+ PM_SKY130_FD_SC_LP__EINVP_8%A
x_PM_SKY130_FD_SC_LP__EINVP_8%VPWR N_VPWR_M1026_s N_VPWR_M1000_d N_VPWR_M1007_d
+ N_VPWR_M1019_d N_VPWR_M1021_d N_VPWR_c_644_n N_VPWR_c_645_n N_VPWR_c_646_n
+ N_VPWR_c_647_n N_VPWR_c_648_n N_VPWR_c_649_n N_VPWR_c_650_n N_VPWR_c_651_n
+ VPWR N_VPWR_c_652_n N_VPWR_c_653_n N_VPWR_c_654_n N_VPWR_c_655_n
+ N_VPWR_c_643_n N_VPWR_c_657_n N_VPWR_c_658_n N_VPWR_c_659_n N_VPWR_c_660_n
+ PM_SKY130_FD_SC_LP__EINVP_8%VPWR
x_PM_SKY130_FD_SC_LP__EINVP_8%A_365_367# N_A_365_367#_M1000_s
+ N_A_365_367#_M1005_s N_A_365_367#_M1016_s N_A_365_367#_M1020_s
+ N_A_365_367#_M1033_s N_A_365_367#_M1006_d N_A_365_367#_M1012_d
+ N_A_365_367#_M1018_d N_A_365_367#_M1032_d N_A_365_367#_c_766_n
+ N_A_365_367#_c_758_n N_A_365_367#_c_759_n N_A_365_367#_c_767_n
+ N_A_365_367#_c_760_n N_A_365_367#_c_768_n N_A_365_367#_c_761_n
+ N_A_365_367#_c_769_n N_A_365_367#_c_762_n N_A_365_367#_c_871_n
+ N_A_365_367#_c_771_n N_A_365_367#_c_822_n N_A_365_367#_c_824_n
+ N_A_365_367#_c_828_n N_A_365_367#_c_830_n N_A_365_367#_c_834_n
+ N_A_365_367#_c_836_n N_A_365_367#_c_840_n N_A_365_367#_c_772_n
+ N_A_365_367#_c_773_n N_A_365_367#_c_763_n N_A_365_367#_c_764_n
+ N_A_365_367#_c_765_n N_A_365_367#_c_844_n N_A_365_367#_c_846_n
+ N_A_365_367#_c_848_n PM_SKY130_FD_SC_LP__EINVP_8%A_365_367#
x_PM_SKY130_FD_SC_LP__EINVP_8%Z N_Z_M1002_s N_Z_M1011_s N_Z_M1022_s N_Z_M1029_s
+ N_Z_M1003_s N_Z_M1009_s N_Z_M1013_s N_Z_M1023_s N_Z_c_995_n N_Z_c_933_n
+ N_Z_c_925_n N_Z_c_998_n N_Z_c_926_n N_Z_c_1001_n N_Z_c_927_n N_Z_c_920_n
+ N_Z_c_921_n N_Z_c_1004_n N_Z_c_1026_p N_Z_c_929_n N_Z_c_930_n N_Z_c_922_n
+ N_Z_c_931_n N_Z_c_923_n N_Z_c_932_n Z Z N_Z_c_986_n
+ PM_SKY130_FD_SC_LP__EINVP_8%Z
x_PM_SKY130_FD_SC_LP__EINVP_8%VGND N_VGND_M1027_s N_VGND_M1001_d N_VGND_M1010_d
+ N_VGND_M1017_d N_VGND_M1028_d N_VGND_c_1031_n N_VGND_c_1032_n N_VGND_c_1033_n
+ N_VGND_c_1034_n N_VGND_c_1035_n N_VGND_c_1036_n N_VGND_c_1037_n
+ N_VGND_c_1038_n VGND N_VGND_c_1039_n N_VGND_c_1040_n N_VGND_c_1041_n
+ N_VGND_c_1042_n N_VGND_c_1043_n N_VGND_c_1044_n N_VGND_c_1045_n
+ N_VGND_c_1046_n N_VGND_c_1047_n PM_SKY130_FD_SC_LP__EINVP_8%VGND
x_PM_SKY130_FD_SC_LP__EINVP_8%A_371_47# N_A_371_47#_M1001_s N_A_371_47#_M1004_s
+ N_A_371_47#_M1014_s N_A_371_47#_M1024_s N_A_371_47#_M1030_s
+ N_A_371_47#_M1008_d N_A_371_47#_M1015_d N_A_371_47#_M1025_d
+ N_A_371_47#_M1031_d N_A_371_47#_c_1140_n N_A_371_47#_c_1141_n
+ N_A_371_47#_c_1142_n N_A_371_47#_c_1143_n N_A_371_47#_c_1144_n
+ N_A_371_47#_c_1145_n N_A_371_47#_c_1146_n N_A_371_47#_c_1147_n
+ N_A_371_47#_c_1148_n N_A_371_47#_c_1192_n N_A_371_47#_c_1193_n
+ N_A_371_47#_c_1204_n N_A_371_47#_c_1210_n N_A_371_47#_c_1149_n
+ N_A_371_47#_c_1150_n N_A_371_47#_c_1151_n N_A_371_47#_c_1212_n
+ N_A_371_47#_c_1152_n PM_SKY130_FD_SC_LP__EINVP_8%A_371_47#
cc_1 VNB N_A_182_367#_c_175_n 0.00583057f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=1.685
cc_2 VNB N_A_182_367#_c_176_n 0.00487805f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=1.685
cc_3 VNB N_A_182_367#_c_177_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=2.52 $Y2=1.65
cc_4 VNB N_A_182_367#_c_178_n 0.00513635f $X=-0.19 $Y=-0.245 $X2=2.95 $Y2=1.65
cc_5 VNB N_A_182_367#_c_179_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=1.65
cc_6 VNB N_A_182_367#_c_180_n 0.0051668f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.65
cc_7 VNB N_A_182_367#_c_181_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=4.24 $Y2=1.65
cc_8 VNB N_A_182_367#_c_182_n 0.00513635f $X=-0.19 $Y=-0.245 $X2=4.67 $Y2=1.65
cc_9 VNB N_A_182_367#_c_183_n 0.00904747f $X=-0.19 $Y=-0.245 $X2=5.1 $Y2=1.65
cc_10 VNB N_A_182_367#_c_184_n 0.00379509f $X=-0.19 $Y=-0.245 $X2=2.165
+ $Y2=1.667
cc_11 VNB N_A_182_367#_c_185_n 0.00279623f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=1.65
cc_12 VNB N_A_182_367#_c_186_n 0.00279623f $X=-0.19 $Y=-0.245 $X2=3.025 $Y2=1.65
cc_13 VNB N_A_182_367#_c_187_n 0.00279623f $X=-0.19 $Y=-0.245 $X2=3.455 $Y2=1.65
cc_14 VNB N_A_182_367#_c_188_n 0.00279623f $X=-0.19 $Y=-0.245 $X2=3.885 $Y2=1.65
cc_15 VNB N_A_182_367#_c_189_n 0.00279623f $X=-0.19 $Y=-0.245 $X2=4.315 $Y2=1.65
cc_16 VNB N_A_182_367#_c_190_n 0.00279623f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=1.65
cc_17 VNB N_A_182_367#_c_191_n 0.0281322f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.49
cc_18 VNB N_TE_M1026_g 0.00214287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_TE_c_338_n 0.0187544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_TE_c_339_n 0.025559f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.93
cc_21 VNB N_TE_c_340_n 0.0222535f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=1.685
cc_22 VNB N_TE_c_341_n 0.0190592f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=1.685
cc_23 VNB N_TE_c_342_n 0.0103769f $X=-0.19 $Y=-0.245 $X2=2.165 $Y2=2.465
cc_24 VNB N_TE_c_343_n 0.0689868f $X=-0.19 $Y=-0.245 $X2=2.52 $Y2=1.65
cc_25 VNB N_TE_c_344_n 0.0159665f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=1.65
cc_26 VNB N_TE_c_345_n 0.0109794f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=2.465
cc_27 VNB N_TE_c_346_n 0.0159665f $X=-0.19 $Y=-0.245 $X2=2.67 $Y2=1.65
cc_28 VNB N_TE_c_347_n 0.0103769f $X=-0.19 $Y=-0.245 $X2=3.025 $Y2=2.465
cc_29 VNB N_TE_c_348_n 0.0159665f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=1.65
cc_30 VNB N_TE_c_349_n 0.0109388f $X=-0.19 $Y=-0.245 $X2=3.455 $Y2=2.465
cc_31 VNB N_TE_c_350_n 0.0159665f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=1.65
cc_32 VNB N_TE_c_351_n 0.0103769f $X=-0.19 $Y=-0.245 $X2=3.885 $Y2=2.465
cc_33 VNB N_TE_c_352_n 0.0159665f $X=-0.19 $Y=-0.245 $X2=3.96 $Y2=1.65
cc_34 VNB N_TE_c_353_n 0.0109794f $X=-0.19 $Y=-0.245 $X2=4.315 $Y2=2.465
cc_35 VNB N_TE_c_354_n 0.0161619f $X=-0.19 $Y=-0.245 $X2=4.39 $Y2=1.65
cc_36 VNB N_TE_c_355_n 0.0175038f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=2.465
cc_37 VNB N_TE_c_356_n 0.0157884f $X=-0.19 $Y=-0.245 $X2=4.82 $Y2=1.65
cc_38 VNB N_TE_c_357_n 0.0766705f $X=-0.19 $Y=-0.245 $X2=5.175 $Y2=2.465
cc_39 VNB N_TE_c_358_n 0.00438817f $X=-0.19 $Y=-0.245 $X2=2.165 $Y2=1.667
cc_40 VNB N_TE_c_359_n 0.00438817f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=1.65
cc_41 VNB N_TE_c_360_n 0.00438817f $X=-0.19 $Y=-0.245 $X2=3.025 $Y2=1.65
cc_42 VNB N_TE_c_361_n 0.00438817f $X=-0.19 $Y=-0.245 $X2=3.455 $Y2=1.65
cc_43 VNB N_TE_c_362_n 0.00438817f $X=-0.19 $Y=-0.245 $X2=3.885 $Y2=1.65
cc_44 VNB N_TE_c_363_n 0.00438817f $X=-0.19 $Y=-0.245 $X2=4.315 $Y2=1.65
cc_45 VNB TE 0.0233322f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.91
cc_46 VNB N_A_M1002_g 0.0222464f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.76
cc_47 VNB N_A_M1008_g 0.0222278f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=1.65
cc_48 VNB N_A_M1011_g 0.0223615f $X=-0.19 $Y=-0.245 $X2=3.025 $Y2=2.465
cc_49 VNB N_A_M1015_g 0.0223561f $X=-0.19 $Y=-0.245 $X2=3.885 $Y2=1.725
cc_50 VNB N_A_M1022_g 0.0228425f $X=-0.19 $Y=-0.245 $X2=4.67 $Y2=1.65
cc_51 VNB N_A_M1025_g 0.0224111f $X=-0.19 $Y=-0.245 $X2=5.175 $Y2=2.465
cc_52 VNB N_A_M1029_g 0.0218146f $X=-0.19 $Y=-0.245 $X2=3.455 $Y2=1.65
cc_53 VNB N_A_M1031_g 0.0327484f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.855
cc_54 VNB N_A_c_493_n 0.00532422f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=2.095
cc_55 VNB N_A_c_494_n 0.00316678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_c_495_n 0.162399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_643_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_365_367#_c_758_n 0.0036176f $X=-0.19 $Y=-0.245 $X2=4.24 $Y2=1.65
cc_59 VNB N_A_365_367#_c_759_n 0.00281705f $X=-0.19 $Y=-0.245 $X2=3.96 $Y2=1.65
cc_60 VNB N_A_365_367#_c_760_n 0.00364785f $X=-0.19 $Y=-0.245 $X2=4.745
+ $Y2=2.465
cc_61 VNB N_A_365_367#_c_761_n 0.00358736f $X=-0.19 $Y=-0.245 $X2=1.542 $Y2=1.93
cc_62 VNB N_A_365_367#_c_762_n 0.00680459f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=1.65
cc_63 VNB N_A_365_367#_c_763_n 0.0016053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_365_367#_c_764_n 0.0016053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_365_367#_c_765_n 0.00163616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Z_c_920_n 0.00344658f $X=-0.19 $Y=-0.245 $X2=5.175 $Y2=2.465
cc_67 VNB N_Z_c_921_n 0.00148732f $X=-0.19 $Y=-0.245 $X2=1.542 $Y2=1.93
cc_68 VNB N_Z_c_922_n 0.00203693f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.49
cc_69 VNB N_Z_c_923_n 0.00215318f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=2.095
cc_70 VNB Z 0.00157368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1031_n 0.0374522f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=2.465
cc_72 VNB N_VGND_c_1032_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=3.025 $Y2=2.465
cc_73 VNB N_VGND_c_1033_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=1.65
cc_74 VNB N_VGND_c_1034_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=3.455 $Y2=2.465
cc_75 VNB N_VGND_c_1035_n 3.14366e-19 $X=-0.19 $Y=-0.245 $X2=3.885 $Y2=2.465
cc_76 VNB N_VGND_c_1036_n 0.0043524f $X=-0.19 $Y=-0.245 $X2=4.315 $Y2=1.725
cc_77 VNB N_VGND_c_1037_n 0.0379344f $X=-0.19 $Y=-0.245 $X2=4.315 $Y2=2.465
cc_78 VNB N_VGND_c_1038_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=4.67 $Y2=1.65
cc_79 VNB N_VGND_c_1039_n 0.0198045f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=2.465
cc_80 VNB N_VGND_c_1040_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=3.025 $Y2=1.65
cc_81 VNB N_VGND_c_1041_n 0.0146078f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.265
cc_82 VNB N_VGND_c_1042_n 0.0964758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1043_n 0.471068f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.02
cc_84 VNB N_VGND_c_1044_n 0.00577043f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=2.095
cc_85 VNB N_VGND_c_1045_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1046_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1047_n 0.00442399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_371_47#_c_1140_n 0.0159055f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=1.65
cc_89 VNB N_A_371_47#_c_1141_n 0.00406129f $X=-0.19 $Y=-0.245 $X2=3.885
+ $Y2=2.465
cc_90 VNB N_A_371_47#_c_1142_n 0.00178925f $X=-0.19 $Y=-0.245 $X2=3.885
+ $Y2=2.465
cc_91 VNB N_A_371_47#_c_1143_n 0.00187197f $X=-0.19 $Y=-0.245 $X2=4.315
+ $Y2=1.725
cc_92 VNB N_A_371_47#_c_1144_n 0.00405982f $X=-0.19 $Y=-0.245 $X2=4.315
+ $Y2=2.465
cc_93 VNB N_A_371_47#_c_1145_n 0.00187197f $X=-0.19 $Y=-0.245 $X2=4.745
+ $Y2=2.465
cc_94 VNB N_A_371_47#_c_1146_n 0.00403545f $X=-0.19 $Y=-0.245 $X2=5.1 $Y2=1.65
cc_95 VNB N_A_371_47#_c_1147_n 0.00179503f $X=-0.19 $Y=-0.245 $X2=5.175
+ $Y2=2.465
cc_96 VNB N_A_371_47#_c_1148_n 0.00647603f $X=-0.19 $Y=-0.245 $X2=1.542 $Y2=1.93
cc_97 VNB N_A_371_47#_c_1149_n 0.00117816f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.49
cc_98 VNB N_A_371_47#_c_1150_n 0.00117816f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.49
cc_99 VNB N_A_371_47#_c_1151_n 0.00136446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_371_47#_c_1152_n 0.0444999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VPB N_A_182_367#_c_175_n 0.0083488f $X=-0.19 $Y=1.655 $X2=2.09 $Y2=1.685
cc_102 VPB N_A_182_367#_c_176_n 0.00498378f $X=-0.19 $Y=1.655 $X2=1.75 $Y2=1.685
cc_103 VPB N_A_182_367#_c_194_n 0.0172093f $X=-0.19 $Y=1.655 $X2=2.165 $Y2=1.76
cc_104 VPB N_A_182_367#_c_177_n 0.00428737f $X=-0.19 $Y=1.655 $X2=2.52 $Y2=1.65
cc_105 VPB N_A_182_367#_c_196_n 0.0161637f $X=-0.19 $Y=1.655 $X2=2.595 $Y2=1.725
cc_106 VPB N_A_182_367#_c_178_n 0.0049292f $X=-0.19 $Y=1.655 $X2=2.95 $Y2=1.65
cc_107 VPB N_A_182_367#_c_198_n 0.0161636f $X=-0.19 $Y=1.655 $X2=3.025 $Y2=1.725
cc_108 VPB N_A_182_367#_c_179_n 0.00428737f $X=-0.19 $Y=1.655 $X2=3.38 $Y2=1.65
cc_109 VPB N_A_182_367#_c_200_n 0.0161637f $X=-0.19 $Y=1.655 $X2=3.455 $Y2=1.725
cc_110 VPB N_A_182_367#_c_180_n 0.0049292f $X=-0.19 $Y=1.655 $X2=3.81 $Y2=1.65
cc_111 VPB N_A_182_367#_c_202_n 0.0161633f $X=-0.19 $Y=1.655 $X2=3.885 $Y2=1.725
cc_112 VPB N_A_182_367#_c_181_n 0.00428737f $X=-0.19 $Y=1.655 $X2=4.24 $Y2=1.65
cc_113 VPB N_A_182_367#_c_204_n 0.0161635f $X=-0.19 $Y=1.655 $X2=4.315 $Y2=1.725
cc_114 VPB N_A_182_367#_c_182_n 0.0049292f $X=-0.19 $Y=1.655 $X2=4.67 $Y2=1.65
cc_115 VPB N_A_182_367#_c_206_n 0.0161635f $X=-0.19 $Y=1.655 $X2=4.745 $Y2=1.725
cc_116 VPB N_A_182_367#_c_183_n 0.00635142f $X=-0.19 $Y=1.655 $X2=5.1 $Y2=1.65
cc_117 VPB N_A_182_367#_c_208_n 0.0163984f $X=-0.19 $Y=1.655 $X2=5.175 $Y2=1.725
cc_118 VPB N_A_182_367#_c_209_n 0.0109757f $X=-0.19 $Y=1.655 $X2=1.542 $Y2=1.93
cc_119 VPB N_A_182_367#_c_210_n 0.0223043f $X=-0.19 $Y=1.655 $X2=1.542 $Y2=2.08
cc_120 VPB N_A_182_367#_c_184_n 0.00228082f $X=-0.19 $Y=1.655 $X2=2.165
+ $Y2=1.667
cc_121 VPB N_A_182_367#_c_185_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.595 $Y2=1.65
cc_122 VPB N_A_182_367#_c_186_n 0.00111435f $X=-0.19 $Y=1.655 $X2=3.025 $Y2=1.65
cc_123 VPB N_A_182_367#_c_187_n 0.00111435f $X=-0.19 $Y=1.655 $X2=3.455 $Y2=1.65
cc_124 VPB N_A_182_367#_c_188_n 0.00111435f $X=-0.19 $Y=1.655 $X2=3.885 $Y2=1.65
cc_125 VPB N_A_182_367#_c_189_n 0.00111435f $X=-0.19 $Y=1.655 $X2=4.315 $Y2=1.65
cc_126 VPB N_A_182_367#_c_190_n 0.00111435f $X=-0.19 $Y=1.655 $X2=4.745 $Y2=1.65
cc_127 VPB N_A_182_367#_c_218_n 0.00517179f $X=-0.19 $Y=1.655 $X2=1.28 $Y2=2.265
cc_128 VPB N_A_182_367#_c_219_n 0.0114277f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=2.91
cc_129 VPB N_A_182_367#_c_191_n 0.00472536f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=0.49
cc_130 VPB N_A_182_367#_c_221_n 0.049013f $X=-0.19 $Y=1.655 $X2=1.5 $Y2=2.095
cc_131 VPB N_TE_M1026_g 0.0308444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB TE 0.0196533f $X=-0.19 $Y=1.655 $X2=1.28 $Y2=2.91
cc_133 VPB N_A_M1003_g 0.0200003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_M1006_g 0.0182261f $X=-0.19 $Y=1.655 $X2=2.165 $Y2=1.76
cc_135 VPB N_A_M1009_g 0.0191281f $X=-0.19 $Y=1.655 $X2=2.95 $Y2=1.65
cc_136 VPB N_A_M1012_g 0.0191449f $X=-0.19 $Y=1.655 $X2=3.455 $Y2=2.465
cc_137 VPB N_A_M1013_g 0.0191459f $X=-0.19 $Y=1.655 $X2=3.96 $Y2=1.65
cc_138 VPB N_A_M1018_g 0.0191155f $X=-0.19 $Y=1.655 $X2=4.745 $Y2=2.465
cc_139 VPB N_A_M1023_g 0.0186727f $X=-0.19 $Y=1.655 $X2=1.542 $Y2=2.08
cc_140 VPB N_A_M1032_g 0.0271375f $X=-0.19 $Y=1.655 $X2=1.28 $Y2=2.265
cc_141 VPB N_A_c_495_n 0.0189846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_644_n 0.0497352f $X=-0.19 $Y=1.655 $X2=2.595 $Y2=2.465
cc_143 VPB N_VPWR_c_645_n 0.00461568f $X=-0.19 $Y=1.655 $X2=3.38 $Y2=1.65
cc_144 VPB N_VPWR_c_646_n 0.0165512f $X=-0.19 $Y=1.655 $X2=3.455 $Y2=2.465
cc_145 VPB N_VPWR_c_647_n 0.00403733f $X=-0.19 $Y=1.655 $X2=3.885 $Y2=2.465
cc_146 VPB N_VPWR_c_648_n 0.00398868f $X=-0.19 $Y=1.655 $X2=4.315 $Y2=2.465
cc_147 VPB N_VPWR_c_649_n 0.00462176f $X=-0.19 $Y=1.655 $X2=5.1 $Y2=1.65
cc_148 VPB N_VPWR_c_650_n 0.0392609f $X=-0.19 $Y=1.655 $X2=5.175 $Y2=2.465
cc_149 VPB N_VPWR_c_651_n 0.00497514f $X=-0.19 $Y=1.655 $X2=1.5 $Y2=2.08
cc_150 VPB N_VPWR_c_652_n 0.0166223f $X=-0.19 $Y=1.655 $X2=2.165 $Y2=1.667
cc_151 VPB N_VPWR_c_653_n 0.0166024f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=2.91
cc_152 VPB N_VPWR_c_654_n 0.0167145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_655_n 0.0941712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_643_n 0.0714363f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_657_n 0.00516749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_658_n 0.00507132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_659_n 0.00487897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_660_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_365_367#_c_766_n 0.0120391f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=1.65
cc_160 VPB N_A_365_367#_c_767_n 0.00176793f $X=-0.19 $Y=1.655 $X2=4.315
+ $Y2=2.465
cc_161 VPB N_A_365_367#_c_768_n 0.00176405f $X=-0.19 $Y=1.655 $X2=5.175
+ $Y2=1.725
cc_162 VPB N_A_365_367#_c_769_n 0.00176014f $X=-0.19 $Y=1.655 $X2=3.025 $Y2=1.65
cc_163 VPB N_A_365_367#_c_762_n 8.74815e-19 $X=-0.19 $Y=1.655 $X2=4.745 $Y2=1.65
cc_164 VPB N_A_365_367#_c_771_n 0.00185697f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.855
cc_165 VPB N_A_365_367#_c_772_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_365_367#_c_773_n 0.0531237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_Z_c_925_n 0.00484398f $X=-0.19 $Y=1.655 $X2=3.885 $Y2=2.465
cc_168 VPB N_Z_c_926_n 0.00304888f $X=-0.19 $Y=1.655 $X2=4.67 $Y2=1.65
cc_169 VPB N_Z_c_927_n 0.00315127f $X=-0.19 $Y=1.655 $X2=4.82 $Y2=1.65
cc_170 VPB N_Z_c_921_n 0.00108488f $X=-0.19 $Y=1.655 $X2=1.542 $Y2=1.93
cc_171 VPB N_Z_c_929_n 0.00246915f $X=-0.19 $Y=1.655 $X2=1.28 $Y2=2.91
cc_172 VPB N_Z_c_930_n 0.00144499f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.855
cc_173 VPB N_Z_c_931_n 0.00144499f $X=-0.19 $Y=1.655 $X2=1.5 $Y2=2.095
cc_174 VPB N_Z_c_932_n 6.46409e-19 $X=-0.19 $Y=1.655 $X2=1.5 $Y2=2.095
cc_175 N_A_182_367#_c_176_n N_TE_M1026_g 0.00248659f $X=1.75 $Y=1.685 $X2=0
+ $Y2=0
cc_176 N_A_182_367#_c_210_n N_TE_M1026_g 0.00892181f $X=1.542 $Y=2.08 $X2=0
+ $Y2=0
cc_177 N_A_182_367#_c_191_n N_TE_M1026_g 0.00425473f $X=1.15 $Y=0.49 $X2=0 $Y2=0
cc_178 N_A_182_367#_c_191_n N_TE_c_338_n 0.00659077f $X=1.15 $Y=0.49 $X2=0 $Y2=0
cc_179 N_A_182_367#_c_210_n N_TE_c_339_n 0.00303025f $X=1.542 $Y=2.08 $X2=0
+ $Y2=0
cc_180 N_A_182_367#_c_218_n N_TE_c_339_n 0.00190957f $X=1.28 $Y=2.265 $X2=0
+ $Y2=0
cc_181 N_A_182_367#_c_191_n N_TE_c_339_n 0.0243318f $X=1.15 $Y=0.49 $X2=0 $Y2=0
cc_182 N_A_182_367#_c_176_n N_TE_c_340_n 2.20331e-19 $X=1.75 $Y=1.685 $X2=0
+ $Y2=0
cc_183 N_A_182_367#_c_218_n N_TE_c_340_n 0.00244958f $X=1.28 $Y=2.265 $X2=0
+ $Y2=0
cc_184 N_A_182_367#_c_191_n N_TE_c_340_n 0.00683262f $X=1.15 $Y=0.49 $X2=0 $Y2=0
cc_185 N_A_182_367#_c_177_n N_TE_c_342_n 0.0146492f $X=2.52 $Y=1.65 $X2=0 $Y2=0
cc_186 N_A_182_367#_c_176_n N_TE_c_343_n 0.0280386f $X=1.75 $Y=1.685 $X2=0 $Y2=0
cc_187 N_A_182_367#_c_210_n N_TE_c_343_n 0.00159416f $X=1.542 $Y=2.08 $X2=0
+ $Y2=0
cc_188 N_A_182_367#_c_184_n N_TE_c_343_n 0.0146492f $X=2.165 $Y=1.667 $X2=0
+ $Y2=0
cc_189 N_A_182_367#_c_218_n N_TE_c_343_n 5.61566e-19 $X=1.28 $Y=2.265 $X2=0
+ $Y2=0
cc_190 N_A_182_367#_c_191_n N_TE_c_343_n 0.00108307f $X=1.15 $Y=0.49 $X2=0 $Y2=0
cc_191 N_A_182_367#_c_178_n N_TE_c_345_n 0.0146492f $X=2.95 $Y=1.65 $X2=0 $Y2=0
cc_192 N_A_182_367#_c_179_n N_TE_c_347_n 0.0146492f $X=3.38 $Y=1.65 $X2=0 $Y2=0
cc_193 N_A_182_367#_c_180_n N_TE_c_349_n 0.0146492f $X=3.81 $Y=1.65 $X2=0 $Y2=0
cc_194 N_A_182_367#_c_181_n N_TE_c_351_n 0.0146492f $X=4.24 $Y=1.65 $X2=0 $Y2=0
cc_195 N_A_182_367#_c_182_n N_TE_c_353_n 0.0146492f $X=4.67 $Y=1.65 $X2=0 $Y2=0
cc_196 N_A_182_367#_c_183_n N_TE_c_355_n 0.0146492f $X=5.1 $Y=1.65 $X2=0 $Y2=0
cc_197 N_A_182_367#_c_185_n N_TE_c_358_n 0.0146492f $X=2.595 $Y=1.65 $X2=0 $Y2=0
cc_198 N_A_182_367#_c_186_n N_TE_c_359_n 0.0146492f $X=3.025 $Y=1.65 $X2=0 $Y2=0
cc_199 N_A_182_367#_c_187_n N_TE_c_360_n 0.0146492f $X=3.455 $Y=1.65 $X2=0 $Y2=0
cc_200 N_A_182_367#_c_188_n N_TE_c_361_n 0.0146492f $X=3.885 $Y=1.65 $X2=0 $Y2=0
cc_201 N_A_182_367#_c_189_n N_TE_c_362_n 0.0146492f $X=4.315 $Y=1.65 $X2=0 $Y2=0
cc_202 N_A_182_367#_c_190_n N_TE_c_363_n 0.0146492f $X=4.745 $Y=1.65 $X2=0 $Y2=0
cc_203 N_A_182_367#_c_191_n TE 0.0364062f $X=1.15 $Y=0.49 $X2=0 $Y2=0
cc_204 N_A_182_367#_c_208_n N_A_M1003_g 0.0109851f $X=5.175 $Y=1.725 $X2=0 $Y2=0
cc_205 N_A_182_367#_c_183_n N_A_c_495_n 0.0109851f $X=5.1 $Y=1.65 $X2=0 $Y2=0
cc_206 N_A_182_367#_c_194_n N_VPWR_c_645_n 0.00366503f $X=2.165 $Y=1.76 $X2=0
+ $Y2=0
cc_207 N_A_182_367#_c_177_n N_VPWR_c_645_n 0.00200847f $X=2.52 $Y=1.65 $X2=0
+ $Y2=0
cc_208 N_A_182_367#_c_196_n N_VPWR_c_645_n 0.00213876f $X=2.595 $Y=1.725 $X2=0
+ $Y2=0
cc_209 N_A_182_367#_c_196_n N_VPWR_c_646_n 0.00585385f $X=2.595 $Y=1.725 $X2=0
+ $Y2=0
cc_210 N_A_182_367#_c_198_n N_VPWR_c_646_n 0.00585385f $X=3.025 $Y=1.725 $X2=0
+ $Y2=0
cc_211 N_A_182_367#_c_198_n N_VPWR_c_647_n 0.00219639f $X=3.025 $Y=1.725 $X2=0
+ $Y2=0
cc_212 N_A_182_367#_c_179_n N_VPWR_c_647_n 0.00200847f $X=3.38 $Y=1.65 $X2=0
+ $Y2=0
cc_213 N_A_182_367#_c_200_n N_VPWR_c_647_n 0.00216866f $X=3.455 $Y=1.725 $X2=0
+ $Y2=0
cc_214 N_A_182_367#_c_202_n N_VPWR_c_648_n 0.00216341f $X=3.885 $Y=1.725 $X2=0
+ $Y2=0
cc_215 N_A_182_367#_c_181_n N_VPWR_c_648_n 0.00200847f $X=4.24 $Y=1.65 $X2=0
+ $Y2=0
cc_216 N_A_182_367#_c_204_n N_VPWR_c_648_n 0.00214286f $X=4.315 $Y=1.725 $X2=0
+ $Y2=0
cc_217 N_A_182_367#_c_206_n N_VPWR_c_649_n 0.00217286f $X=4.745 $Y=1.725 $X2=0
+ $Y2=0
cc_218 N_A_182_367#_c_183_n N_VPWR_c_649_n 0.00200847f $X=5.1 $Y=1.65 $X2=0
+ $Y2=0
cc_219 N_A_182_367#_c_208_n N_VPWR_c_649_n 0.0036292f $X=5.175 $Y=1.725 $X2=0
+ $Y2=0
cc_220 N_A_182_367#_c_194_n N_VPWR_c_650_n 0.00585385f $X=2.165 $Y=1.76 $X2=0
+ $Y2=0
cc_221 N_A_182_367#_c_219_n N_VPWR_c_650_n 0.0468406f $X=1.05 $Y=2.91 $X2=0
+ $Y2=0
cc_222 N_A_182_367#_c_221_n N_VPWR_c_650_n 0.00169265f $X=1.5 $Y=2.095 $X2=0
+ $Y2=0
cc_223 N_A_182_367#_c_200_n N_VPWR_c_653_n 0.00585385f $X=3.455 $Y=1.725 $X2=0
+ $Y2=0
cc_224 N_A_182_367#_c_202_n N_VPWR_c_653_n 0.00585385f $X=3.885 $Y=1.725 $X2=0
+ $Y2=0
cc_225 N_A_182_367#_c_204_n N_VPWR_c_654_n 0.00585385f $X=4.315 $Y=1.725 $X2=0
+ $Y2=0
cc_226 N_A_182_367#_c_206_n N_VPWR_c_654_n 0.00585385f $X=4.745 $Y=1.725 $X2=0
+ $Y2=0
cc_227 N_A_182_367#_c_208_n N_VPWR_c_655_n 0.00585385f $X=5.175 $Y=1.725 $X2=0
+ $Y2=0
cc_228 N_A_182_367#_M1026_d N_VPWR_c_643_n 0.00336915f $X=0.91 $Y=1.835 $X2=0
+ $Y2=0
cc_229 N_A_182_367#_c_194_n N_VPWR_c_643_n 0.0118084f $X=2.165 $Y=1.76 $X2=0
+ $Y2=0
cc_230 N_A_182_367#_c_196_n N_VPWR_c_643_n 0.0105361f $X=2.595 $Y=1.725 $X2=0
+ $Y2=0
cc_231 N_A_182_367#_c_198_n N_VPWR_c_643_n 0.0105087f $X=3.025 $Y=1.725 $X2=0
+ $Y2=0
cc_232 N_A_182_367#_c_200_n N_VPWR_c_643_n 0.0105224f $X=3.455 $Y=1.725 $X2=0
+ $Y2=0
cc_233 N_A_182_367#_c_202_n N_VPWR_c_643_n 0.0105224f $X=3.885 $Y=1.725 $X2=0
+ $Y2=0
cc_234 N_A_182_367#_c_204_n N_VPWR_c_643_n 0.0105361f $X=4.315 $Y=1.725 $X2=0
+ $Y2=0
cc_235 N_A_182_367#_c_206_n N_VPWR_c_643_n 0.0105224f $X=4.745 $Y=1.725 $X2=0
+ $Y2=0
cc_236 N_A_182_367#_c_208_n N_VPWR_c_643_n 0.0105477f $X=5.175 $Y=1.725 $X2=0
+ $Y2=0
cc_237 N_A_182_367#_c_219_n N_VPWR_c_643_n 0.0259703f $X=1.05 $Y=2.91 $X2=0
+ $Y2=0
cc_238 N_A_182_367#_c_221_n N_VPWR_c_643_n 0.00139091f $X=1.5 $Y=2.095 $X2=0
+ $Y2=0
cc_239 N_A_182_367#_c_175_n N_A_365_367#_c_766_n 0.0061983f $X=2.09 $Y=1.685
+ $X2=0 $Y2=0
cc_240 N_A_182_367#_c_194_n N_A_365_367#_c_766_n 0.00285595f $X=2.165 $Y=1.76
+ $X2=0 $Y2=0
cc_241 N_A_182_367#_c_209_n N_A_365_367#_c_766_n 0.00368672f $X=1.542 $Y=1.93
+ $X2=0 $Y2=0
cc_242 N_A_182_367#_c_218_n N_A_365_367#_c_766_n 0.0308398f $X=1.28 $Y=2.265
+ $X2=0 $Y2=0
cc_243 N_A_182_367#_c_219_n N_A_365_367#_c_766_n 0.069037f $X=1.05 $Y=2.91 $X2=0
+ $Y2=0
cc_244 N_A_182_367#_c_191_n N_A_365_367#_c_766_n 0.00523045f $X=1.15 $Y=0.49
+ $X2=0 $Y2=0
cc_245 N_A_182_367#_c_221_n N_A_365_367#_c_766_n 0.00470837f $X=1.5 $Y=2.095
+ $X2=0 $Y2=0
cc_246 N_A_182_367#_c_175_n N_A_365_367#_c_758_n 7.60673e-19 $X=2.09 $Y=1.685
+ $X2=0 $Y2=0
cc_247 N_A_182_367#_c_177_n N_A_365_367#_c_758_n 0.00784018f $X=2.52 $Y=1.65
+ $X2=0 $Y2=0
cc_248 N_A_182_367#_c_184_n N_A_365_367#_c_758_n 0.00966608f $X=2.165 $Y=1.667
+ $X2=0 $Y2=0
cc_249 N_A_182_367#_c_185_n N_A_365_367#_c_758_n 0.00895896f $X=2.595 $Y=1.65
+ $X2=0 $Y2=0
cc_250 N_A_182_367#_c_175_n N_A_365_367#_c_759_n 0.00608319f $X=2.09 $Y=1.685
+ $X2=0 $Y2=0
cc_251 N_A_182_367#_c_191_n N_A_365_367#_c_759_n 0.00683888f $X=1.15 $Y=0.49
+ $X2=0 $Y2=0
cc_252 N_A_182_367#_c_196_n N_A_365_367#_c_767_n 0.00228772f $X=2.595 $Y=1.725
+ $X2=0 $Y2=0
cc_253 N_A_182_367#_c_178_n N_A_365_367#_c_767_n 0.00250619f $X=2.95 $Y=1.65
+ $X2=0 $Y2=0
cc_254 N_A_182_367#_c_198_n N_A_365_367#_c_767_n 0.00224781f $X=3.025 $Y=1.725
+ $X2=0 $Y2=0
cc_255 N_A_182_367#_c_178_n N_A_365_367#_c_760_n 7.76443e-19 $X=2.95 $Y=1.65
+ $X2=0 $Y2=0
cc_256 N_A_182_367#_c_179_n N_A_365_367#_c_760_n 0.00768727f $X=3.38 $Y=1.65
+ $X2=0 $Y2=0
cc_257 N_A_182_367#_c_180_n N_A_365_367#_c_760_n 4.77811e-19 $X=3.81 $Y=1.65
+ $X2=0 $Y2=0
cc_258 N_A_182_367#_c_186_n N_A_365_367#_c_760_n 0.00895896f $X=3.025 $Y=1.65
+ $X2=0 $Y2=0
cc_259 N_A_182_367#_c_187_n N_A_365_367#_c_760_n 0.00895896f $X=3.455 $Y=1.65
+ $X2=0 $Y2=0
cc_260 N_A_182_367#_c_200_n N_A_365_367#_c_768_n 0.00227094f $X=3.455 $Y=1.725
+ $X2=0 $Y2=0
cc_261 N_A_182_367#_c_180_n N_A_365_367#_c_768_n 0.00250619f $X=3.81 $Y=1.65
+ $X2=0 $Y2=0
cc_262 N_A_182_367#_c_202_n N_A_365_367#_c_768_n 0.00225773f $X=3.885 $Y=1.725
+ $X2=0 $Y2=0
cc_263 N_A_182_367#_c_180_n N_A_365_367#_c_761_n 4.77811e-19 $X=3.81 $Y=1.65
+ $X2=0 $Y2=0
cc_264 N_A_182_367#_c_181_n N_A_365_367#_c_761_n 0.0079931f $X=4.24 $Y=1.65
+ $X2=0 $Y2=0
cc_265 N_A_182_367#_c_188_n N_A_365_367#_c_761_n 0.00895896f $X=3.885 $Y=1.65
+ $X2=0 $Y2=0
cc_266 N_A_182_367#_c_189_n N_A_365_367#_c_761_n 0.00895896f $X=4.315 $Y=1.65
+ $X2=0 $Y2=0
cc_267 N_A_182_367#_c_204_n N_A_365_367#_c_769_n 0.00228574f $X=4.315 $Y=1.725
+ $X2=0 $Y2=0
cc_268 N_A_182_367#_c_182_n N_A_365_367#_c_769_n 0.00250807f $X=4.67 $Y=1.65
+ $X2=0 $Y2=0
cc_269 N_A_182_367#_c_206_n N_A_365_367#_c_769_n 0.00226903f $X=4.745 $Y=1.725
+ $X2=0 $Y2=0
cc_270 N_A_182_367#_c_182_n N_A_365_367#_c_762_n 4.77811e-19 $X=4.67 $Y=1.65
+ $X2=0 $Y2=0
cc_271 N_A_182_367#_c_183_n N_A_365_367#_c_762_n 0.0182127f $X=5.1 $Y=1.65 $X2=0
+ $Y2=0
cc_272 N_A_182_367#_c_190_n N_A_365_367#_c_762_n 0.00895896f $X=4.745 $Y=1.65
+ $X2=0 $Y2=0
cc_273 N_A_182_367#_c_183_n N_A_365_367#_c_771_n 0.00233164f $X=5.1 $Y=1.65
+ $X2=0 $Y2=0
cc_274 N_A_182_367#_c_178_n N_A_365_367#_c_763_n 0.00406286f $X=2.95 $Y=1.65
+ $X2=0 $Y2=0
cc_275 N_A_182_367#_c_180_n N_A_365_367#_c_764_n 0.00406286f $X=3.81 $Y=1.65
+ $X2=0 $Y2=0
cc_276 N_A_182_367#_c_182_n N_A_365_367#_c_765_n 0.00414099f $X=4.67 $Y=1.65
+ $X2=0 $Y2=0
cc_277 N_A_182_367#_c_191_n N_VGND_c_1031_n 0.0072808f $X=1.15 $Y=0.49 $X2=0
+ $Y2=0
cc_278 N_A_182_367#_c_191_n N_VGND_c_1037_n 0.0206458f $X=1.15 $Y=0.49 $X2=0
+ $Y2=0
cc_279 N_A_182_367#_c_191_n N_VGND_c_1043_n 0.0111968f $X=1.15 $Y=0.49 $X2=0
+ $Y2=0
cc_280 N_A_182_367#_c_191_n N_A_371_47#_c_1140_n 0.0365494f $X=1.15 $Y=0.49
+ $X2=0 $Y2=0
cc_281 N_A_182_367#_c_184_n N_A_371_47#_c_1141_n 0.0017973f $X=2.165 $Y=1.667
+ $X2=0 $Y2=0
cc_282 N_A_182_367#_c_175_n N_A_371_47#_c_1142_n 8.76984e-19 $X=2.09 $Y=1.685
+ $X2=0 $Y2=0
cc_283 N_A_182_367#_c_191_n N_A_371_47#_c_1142_n 0.00582532f $X=1.15 $Y=0.49
+ $X2=0 $Y2=0
cc_284 N_A_182_367#_c_178_n N_A_371_47#_c_1144_n 0.00183861f $X=2.95 $Y=1.65
+ $X2=0 $Y2=0
cc_285 N_A_182_367#_c_180_n N_A_371_47#_c_1146_n 0.0018385f $X=3.81 $Y=1.65
+ $X2=0 $Y2=0
cc_286 N_A_182_367#_c_190_n N_A_371_47#_c_1148_n 0.00154902f $X=4.745 $Y=1.65
+ $X2=0 $Y2=0
cc_287 N_A_182_367#_c_178_n N_A_371_47#_c_1149_n 6.75551e-19 $X=2.95 $Y=1.65
+ $X2=0 $Y2=0
cc_288 N_A_182_367#_c_180_n N_A_371_47#_c_1150_n 6.75551e-19 $X=3.81 $Y=1.65
+ $X2=0 $Y2=0
cc_289 N_A_182_367#_c_182_n N_A_371_47#_c_1151_n 7.84392e-19 $X=4.67 $Y=1.65
+ $X2=0 $Y2=0
cc_290 N_TE_c_356_n N_A_M1002_g 0.0250117f $X=5.205 $Y=1.185 $X2=0 $Y2=0
cc_291 N_TE_c_355_n N_A_c_495_n 0.00210865f $X=5.13 $Y=1.275 $X2=0 $Y2=0
cc_292 N_TE_M1026_g N_VPWR_c_644_n 0.00634905f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_293 N_TE_c_357_n N_VPWR_c_644_n 0.00151315f $X=0.76 $Y=1.46 $X2=0 $Y2=0
cc_294 TE N_VPWR_c_644_n 0.0232247f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_295 N_TE_M1026_g N_VPWR_c_650_n 0.00585385f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_296 N_TE_M1026_g N_VPWR_c_643_n 0.0131901f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_297 N_TE_c_343_n N_A_365_367#_c_758_n 0.00168865f $X=2.27 $Y=1.275 $X2=0
+ $Y2=0
cc_298 N_TE_c_343_n N_A_365_367#_c_759_n 0.00178131f $X=2.27 $Y=1.275 $X2=0
+ $Y2=0
cc_299 N_TE_c_345_n N_A_365_367#_c_760_n 0.00170005f $X=2.98 $Y=1.275 $X2=0
+ $Y2=0
cc_300 N_TE_c_349_n N_A_365_367#_c_761_n 0.00166904f $X=3.84 $Y=1.275 $X2=0
+ $Y2=0
cc_301 N_TE_c_353_n N_A_365_367#_c_762_n 0.00174349f $X=4.7 $Y=1.275 $X2=0 $Y2=0
cc_302 N_TE_c_358_n N_A_365_367#_c_763_n 9.48633e-19 $X=2.625 $Y=1.275 $X2=0
+ $Y2=0
cc_303 N_TE_c_360_n N_A_365_367#_c_764_n 9.51527e-19 $X=3.485 $Y=1.275 $X2=0
+ $Y2=0
cc_304 N_TE_c_362_n N_A_365_367#_c_765_n 9.66765e-19 $X=4.345 $Y=1.275 $X2=0
+ $Y2=0
cc_305 N_TE_c_338_n N_VGND_c_1031_n 0.00370214f $X=0.935 $Y=1.26 $X2=0 $Y2=0
cc_306 N_TE_c_357_n N_VGND_c_1031_n 0.0015761f $X=0.76 $Y=1.46 $X2=0 $Y2=0
cc_307 TE N_VGND_c_1031_n 0.0223336f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_308 N_TE_c_341_n N_VGND_c_1032_n 0.0162749f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_309 N_TE_c_342_n N_VGND_c_1032_n 0.00213216f $X=2.55 $Y=1.275 $X2=0 $Y2=0
cc_310 N_TE_c_344_n N_VGND_c_1032_n 0.0144015f $X=2.625 $Y=1.185 $X2=0 $Y2=0
cc_311 N_TE_c_346_n N_VGND_c_1032_n 6.72004e-19 $X=3.055 $Y=1.185 $X2=0 $Y2=0
cc_312 N_TE_c_344_n N_VGND_c_1033_n 0.00486043f $X=2.625 $Y=1.185 $X2=0 $Y2=0
cc_313 N_TE_c_346_n N_VGND_c_1033_n 0.00486043f $X=3.055 $Y=1.185 $X2=0 $Y2=0
cc_314 N_TE_c_344_n N_VGND_c_1034_n 6.72004e-19 $X=2.625 $Y=1.185 $X2=0 $Y2=0
cc_315 N_TE_c_346_n N_VGND_c_1034_n 0.0144015f $X=3.055 $Y=1.185 $X2=0 $Y2=0
cc_316 N_TE_c_347_n N_VGND_c_1034_n 0.00213216f $X=3.41 $Y=1.275 $X2=0 $Y2=0
cc_317 N_TE_c_348_n N_VGND_c_1034_n 0.0144015f $X=3.485 $Y=1.185 $X2=0 $Y2=0
cc_318 N_TE_c_350_n N_VGND_c_1034_n 6.72004e-19 $X=3.915 $Y=1.185 $X2=0 $Y2=0
cc_319 N_TE_c_348_n N_VGND_c_1035_n 6.72004e-19 $X=3.485 $Y=1.185 $X2=0 $Y2=0
cc_320 N_TE_c_350_n N_VGND_c_1035_n 0.0144015f $X=3.915 $Y=1.185 $X2=0 $Y2=0
cc_321 N_TE_c_351_n N_VGND_c_1035_n 0.00213216f $X=4.27 $Y=1.275 $X2=0 $Y2=0
cc_322 N_TE_c_352_n N_VGND_c_1035_n 0.0144708f $X=4.345 $Y=1.185 $X2=0 $Y2=0
cc_323 N_TE_c_354_n N_VGND_c_1035_n 6.84211e-19 $X=4.775 $Y=1.185 $X2=0 $Y2=0
cc_324 N_TE_c_354_n N_VGND_c_1036_n 0.00216829f $X=4.775 $Y=1.185 $X2=0 $Y2=0
cc_325 N_TE_c_355_n N_VGND_c_1036_n 0.00213216f $X=5.13 $Y=1.275 $X2=0 $Y2=0
cc_326 N_TE_c_356_n N_VGND_c_1036_n 0.00339569f $X=5.205 $Y=1.185 $X2=0 $Y2=0
cc_327 N_TE_c_338_n N_VGND_c_1037_n 0.00482246f $X=0.935 $Y=1.26 $X2=0 $Y2=0
cc_328 N_TE_c_341_n N_VGND_c_1037_n 0.00486043f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_329 N_TE_c_348_n N_VGND_c_1040_n 0.00486043f $X=3.485 $Y=1.185 $X2=0 $Y2=0
cc_330 N_TE_c_350_n N_VGND_c_1040_n 0.00486043f $X=3.915 $Y=1.185 $X2=0 $Y2=0
cc_331 N_TE_c_352_n N_VGND_c_1041_n 0.00486043f $X=4.345 $Y=1.185 $X2=0 $Y2=0
cc_332 N_TE_c_354_n N_VGND_c_1041_n 0.00585385f $X=4.775 $Y=1.185 $X2=0 $Y2=0
cc_333 N_TE_c_356_n N_VGND_c_1042_n 0.00548125f $X=5.205 $Y=1.185 $X2=0 $Y2=0
cc_334 N_TE_c_338_n N_VGND_c_1043_n 0.0100187f $X=0.935 $Y=1.26 $X2=0 $Y2=0
cc_335 N_TE_c_341_n N_VGND_c_1043_n 0.00954696f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_336 N_TE_c_344_n N_VGND_c_1043_n 0.00824727f $X=2.625 $Y=1.185 $X2=0 $Y2=0
cc_337 N_TE_c_346_n N_VGND_c_1043_n 0.00824727f $X=3.055 $Y=1.185 $X2=0 $Y2=0
cc_338 N_TE_c_348_n N_VGND_c_1043_n 0.00824727f $X=3.485 $Y=1.185 $X2=0 $Y2=0
cc_339 N_TE_c_350_n N_VGND_c_1043_n 0.00824727f $X=3.915 $Y=1.185 $X2=0 $Y2=0
cc_340 N_TE_c_352_n N_VGND_c_1043_n 0.00824727f $X=4.345 $Y=1.185 $X2=0 $Y2=0
cc_341 N_TE_c_354_n N_VGND_c_1043_n 0.0105087f $X=4.775 $Y=1.185 $X2=0 $Y2=0
cc_342 N_TE_c_356_n N_VGND_c_1043_n 0.00975463f $X=5.205 $Y=1.185 $X2=0 $Y2=0
cc_343 N_TE_c_341_n N_A_371_47#_c_1140_n 0.00551568f $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_344 N_TE_c_343_n N_A_371_47#_c_1140_n 0.00796101f $X=2.27 $Y=1.275 $X2=0
+ $Y2=0
cc_345 N_TE_c_342_n N_A_371_47#_c_1141_n 0.00745675f $X=2.55 $Y=1.275 $X2=0
+ $Y2=0
cc_346 N_TE_c_343_n N_A_371_47#_c_1141_n 0.0106511f $X=2.27 $Y=1.275 $X2=0 $Y2=0
cc_347 N_TE_c_345_n N_A_371_47#_c_1141_n 0.00259328f $X=2.98 $Y=1.275 $X2=0
+ $Y2=0
cc_348 N_TE_c_358_n N_A_371_47#_c_1141_n 0.00831233f $X=2.625 $Y=1.275 $X2=0
+ $Y2=0
cc_349 N_TE_c_343_n N_A_371_47#_c_1142_n 0.00871339f $X=2.27 $Y=1.275 $X2=0
+ $Y2=0
cc_350 N_TE_c_344_n N_A_371_47#_c_1143_n 0.00198932f $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_351 N_TE_c_345_n N_A_371_47#_c_1143_n 0.00421045f $X=2.98 $Y=1.275 $X2=0
+ $Y2=0
cc_352 N_TE_c_346_n N_A_371_47#_c_1143_n 0.00198932f $X=3.055 $Y=1.185 $X2=0
+ $Y2=0
cc_353 N_TE_c_345_n N_A_371_47#_c_1144_n 0.00259328f $X=2.98 $Y=1.275 $X2=0
+ $Y2=0
cc_354 N_TE_c_347_n N_A_371_47#_c_1144_n 0.00745675f $X=3.41 $Y=1.275 $X2=0
+ $Y2=0
cc_355 N_TE_c_349_n N_A_371_47#_c_1144_n 0.00259328f $X=3.84 $Y=1.275 $X2=0
+ $Y2=0
cc_356 N_TE_c_359_n N_A_371_47#_c_1144_n 0.00831233f $X=3.055 $Y=1.275 $X2=0
+ $Y2=0
cc_357 N_TE_c_360_n N_A_371_47#_c_1144_n 0.00831233f $X=3.485 $Y=1.275 $X2=0
+ $Y2=0
cc_358 N_TE_c_348_n N_A_371_47#_c_1145_n 0.00198932f $X=3.485 $Y=1.185 $X2=0
+ $Y2=0
cc_359 N_TE_c_349_n N_A_371_47#_c_1145_n 0.00421045f $X=3.84 $Y=1.275 $X2=0
+ $Y2=0
cc_360 N_TE_c_350_n N_A_371_47#_c_1145_n 0.00198932f $X=3.915 $Y=1.185 $X2=0
+ $Y2=0
cc_361 N_TE_c_349_n N_A_371_47#_c_1146_n 0.00258696f $X=3.84 $Y=1.275 $X2=0
+ $Y2=0
cc_362 N_TE_c_351_n N_A_371_47#_c_1146_n 0.00745675f $X=4.27 $Y=1.275 $X2=0
+ $Y2=0
cc_363 N_TE_c_353_n N_A_371_47#_c_1146_n 0.00259328f $X=4.7 $Y=1.275 $X2=0 $Y2=0
cc_364 N_TE_c_361_n N_A_371_47#_c_1146_n 0.00831233f $X=3.915 $Y=1.275 $X2=0
+ $Y2=0
cc_365 N_TE_c_362_n N_A_371_47#_c_1146_n 0.00831233f $X=4.345 $Y=1.275 $X2=0
+ $Y2=0
cc_366 N_TE_c_352_n N_A_371_47#_c_1147_n 0.00202385f $X=4.345 $Y=1.185 $X2=0
+ $Y2=0
cc_367 N_TE_c_353_n N_A_371_47#_c_1147_n 0.00421795f $X=4.7 $Y=1.275 $X2=0 $Y2=0
cc_368 N_TE_c_354_n N_A_371_47#_c_1147_n 0.00202583f $X=4.775 $Y=1.185 $X2=0
+ $Y2=0
cc_369 N_TE_c_353_n N_A_371_47#_c_1148_n 7.84014e-19 $X=4.7 $Y=1.275 $X2=0 $Y2=0
cc_370 N_TE_c_355_n N_A_371_47#_c_1148_n 0.0189841f $X=5.13 $Y=1.275 $X2=0 $Y2=0
cc_371 N_TE_c_363_n N_A_371_47#_c_1148_n 0.00904631f $X=4.775 $Y=1.275 $X2=0
+ $Y2=0
cc_372 N_TE_c_356_n N_A_371_47#_c_1192_n 0.00306942f $X=5.205 $Y=1.185 $X2=0
+ $Y2=0
cc_373 N_TE_c_354_n N_A_371_47#_c_1193_n 5.0305e-19 $X=4.775 $Y=1.185 $X2=0
+ $Y2=0
cc_374 N_TE_c_355_n N_A_371_47#_c_1193_n 9.63251e-19 $X=5.13 $Y=1.275 $X2=0
+ $Y2=0
cc_375 N_TE_c_356_n N_A_371_47#_c_1193_n 0.0106477f $X=5.205 $Y=1.185 $X2=0
+ $Y2=0
cc_376 N_TE_c_345_n N_A_371_47#_c_1149_n 0.00307987f $X=2.98 $Y=1.275 $X2=0
+ $Y2=0
cc_377 N_TE_c_349_n N_A_371_47#_c_1150_n 0.00307987f $X=3.84 $Y=1.275 $X2=0
+ $Y2=0
cc_378 N_TE_c_353_n N_A_371_47#_c_1151_n 0.00356616f $X=4.7 $Y=1.275 $X2=0 $Y2=0
cc_379 N_A_M1003_g N_VPWR_c_655_n 0.00357877f $X=5.605 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A_M1006_g N_VPWR_c_655_n 0.00357842f $X=6.035 $Y=2.465 $X2=0 $Y2=0
cc_381 N_A_M1009_g N_VPWR_c_655_n 0.00357842f $X=6.465 $Y=2.465 $X2=0 $Y2=0
cc_382 N_A_M1012_g N_VPWR_c_655_n 0.00357842f $X=6.895 $Y=2.465 $X2=0 $Y2=0
cc_383 N_A_M1013_g N_VPWR_c_655_n 0.00357842f $X=7.325 $Y=2.465 $X2=0 $Y2=0
cc_384 N_A_M1018_g N_VPWR_c_655_n 0.00357842f $X=7.755 $Y=2.465 $X2=0 $Y2=0
cc_385 N_A_M1023_g N_VPWR_c_655_n 0.00357842f $X=8.185 $Y=2.465 $X2=0 $Y2=0
cc_386 N_A_M1032_g N_VPWR_c_655_n 0.00357877f $X=8.615 $Y=2.465 $X2=0 $Y2=0
cc_387 N_A_M1003_g N_VPWR_c_643_n 0.00537654f $X=5.605 $Y=2.465 $X2=0 $Y2=0
cc_388 N_A_M1006_g N_VPWR_c_643_n 0.00535118f $X=6.035 $Y=2.465 $X2=0 $Y2=0
cc_389 N_A_M1009_g N_VPWR_c_643_n 0.00535118f $X=6.465 $Y=2.465 $X2=0 $Y2=0
cc_390 N_A_M1012_g N_VPWR_c_643_n 0.00535118f $X=6.895 $Y=2.465 $X2=0 $Y2=0
cc_391 N_A_M1013_g N_VPWR_c_643_n 0.00535118f $X=7.325 $Y=2.465 $X2=0 $Y2=0
cc_392 N_A_M1018_g N_VPWR_c_643_n 0.00535118f $X=7.755 $Y=2.465 $X2=0 $Y2=0
cc_393 N_A_M1023_g N_VPWR_c_643_n 0.00535118f $X=8.185 $Y=2.465 $X2=0 $Y2=0
cc_394 N_A_M1032_g N_VPWR_c_643_n 0.00631099f $X=8.615 $Y=2.465 $X2=0 $Y2=0
cc_395 N_A_c_495_n N_A_365_367#_c_762_n 0.00224981f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_396 N_A_M1003_g N_A_365_367#_c_771_n 0.00158827f $X=5.605 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_A_M1003_g N_A_365_367#_c_822_n 0.012237f $X=5.605 $Y=2.465 $X2=0 $Y2=0
cc_398 N_A_M1006_g N_A_365_367#_c_822_n 0.010474f $X=6.035 $Y=2.465 $X2=0 $Y2=0
cc_399 N_A_M1003_g N_A_365_367#_c_824_n 6.21331e-19 $X=5.605 $Y=2.465 $X2=0
+ $Y2=0
cc_400 N_A_M1006_g N_A_365_367#_c_824_n 0.00975565f $X=6.035 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_A_M1009_g N_A_365_367#_c_824_n 0.00964814f $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_402 N_A_M1012_g N_A_365_367#_c_824_n 6.13082e-19 $X=6.895 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A_M1009_g N_A_365_367#_c_828_n 0.0105205f $X=6.465 $Y=2.465 $X2=0 $Y2=0
cc_404 N_A_M1012_g N_A_365_367#_c_828_n 0.0105205f $X=6.895 $Y=2.465 $X2=0 $Y2=0
cc_405 N_A_M1009_g N_A_365_367#_c_830_n 6.13082e-19 $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_406 N_A_M1012_g N_A_365_367#_c_830_n 0.00964814f $X=6.895 $Y=2.465 $X2=0
+ $Y2=0
cc_407 N_A_M1013_g N_A_365_367#_c_830_n 0.00964814f $X=7.325 $Y=2.465 $X2=0
+ $Y2=0
cc_408 N_A_M1018_g N_A_365_367#_c_830_n 6.13082e-19 $X=7.755 $Y=2.465 $X2=0
+ $Y2=0
cc_409 N_A_M1013_g N_A_365_367#_c_834_n 0.0105205f $X=7.325 $Y=2.465 $X2=0 $Y2=0
cc_410 N_A_M1018_g N_A_365_367#_c_834_n 0.0105205f $X=7.755 $Y=2.465 $X2=0 $Y2=0
cc_411 N_A_M1013_g N_A_365_367#_c_836_n 6.13082e-19 $X=7.325 $Y=2.465 $X2=0
+ $Y2=0
cc_412 N_A_M1018_g N_A_365_367#_c_836_n 0.00964814f $X=7.755 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_A_M1023_g N_A_365_367#_c_836_n 0.00975666f $X=8.185 $Y=2.465 $X2=0
+ $Y2=0
cc_414 N_A_M1032_g N_A_365_367#_c_836_n 6.21331e-19 $X=8.615 $Y=2.465 $X2=0
+ $Y2=0
cc_415 N_A_M1023_g N_A_365_367#_c_840_n 0.0105205f $X=8.185 $Y=2.465 $X2=0 $Y2=0
cc_416 N_A_M1032_g N_A_365_367#_c_840_n 0.012237f $X=8.615 $Y=2.465 $X2=0 $Y2=0
cc_417 N_A_M1032_g N_A_365_367#_c_773_n 0.00346806f $X=8.615 $Y=2.465 $X2=0
+ $Y2=0
cc_418 N_A_c_495_n N_A_365_367#_c_773_n 6.84763e-19 $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_419 N_A_M1006_g N_A_365_367#_c_844_n 5.89773e-19 $X=6.035 $Y=2.465 $X2=0
+ $Y2=0
cc_420 N_A_M1009_g N_A_365_367#_c_844_n 5.89773e-19 $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_421 N_A_M1012_g N_A_365_367#_c_846_n 5.89773e-19 $X=6.895 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_M1013_g N_A_365_367#_c_846_n 5.89773e-19 $X=7.325 $Y=2.465 $X2=0
+ $Y2=0
cc_423 N_A_M1018_g N_A_365_367#_c_848_n 5.89773e-19 $X=7.755 $Y=2.465 $X2=0
+ $Y2=0
cc_424 N_A_M1023_g N_A_365_367#_c_848_n 5.89773e-19 $X=8.185 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_M1008_g N_Z_c_933_n 0.00440183f $X=6.065 $Y=0.655 $X2=0 $Y2=0
cc_426 N_A_M1011_g N_Z_c_933_n 0.0113095f $X=6.495 $Y=0.655 $X2=0 $Y2=0
cc_427 N_A_M1015_g N_Z_c_933_n 0.0113838f $X=6.925 $Y=0.655 $X2=0 $Y2=0
cc_428 N_A_M1022_g N_Z_c_933_n 0.0125519f $X=7.355 $Y=0.655 $X2=0 $Y2=0
cc_429 N_A_c_559_p N_Z_c_933_n 0.0061577f $X=7.82 $Y=1.49 $X2=0 $Y2=0
cc_430 N_A_c_493_n N_Z_c_933_n 0.05509f $X=7.053 $Y=1.402 $X2=0 $Y2=0
cc_431 N_A_c_495_n N_Z_c_933_n 0.00342994f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_432 N_A_M1006_g N_Z_c_925_n 6.34533e-19 $X=6.035 $Y=2.465 $X2=0 $Y2=0
cc_433 N_A_M1009_g N_Z_c_925_n 0.0127344f $X=6.465 $Y=2.465 $X2=0 $Y2=0
cc_434 N_A_c_493_n N_Z_c_925_n 0.0214581f $X=7.053 $Y=1.402 $X2=0 $Y2=0
cc_435 N_A_c_495_n N_Z_c_925_n 0.00405554f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_436 N_A_M1012_g N_Z_c_926_n 0.013073f $X=6.895 $Y=2.465 $X2=0 $Y2=0
cc_437 N_A_M1013_g N_Z_c_926_n 0.0130918f $X=7.325 $Y=2.465 $X2=0 $Y2=0
cc_438 N_A_c_493_n N_Z_c_926_n 0.0491942f $X=7.053 $Y=1.402 $X2=0 $Y2=0
cc_439 N_A_c_495_n N_Z_c_926_n 0.00253271f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_440 N_A_M1018_g N_Z_c_927_n 0.0130453f $X=7.755 $Y=2.465 $X2=0 $Y2=0
cc_441 N_A_M1023_g N_Z_c_927_n 0.00507842f $X=8.185 $Y=2.465 $X2=0 $Y2=0
cc_442 N_A_c_559_p N_Z_c_927_n 0.0251603f $X=7.82 $Y=1.49 $X2=0 $Y2=0
cc_443 N_A_c_495_n N_Z_c_927_n 0.00269875f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_444 N_A_M1025_g N_Z_c_920_n 0.010047f $X=7.785 $Y=0.655 $X2=0 $Y2=0
cc_445 N_A_M1029_g N_Z_c_920_n 0.00274854f $X=8.215 $Y=0.655 $X2=0 $Y2=0
cc_446 N_A_c_559_p N_Z_c_920_n 0.0229905f $X=7.82 $Y=1.49 $X2=0 $Y2=0
cc_447 N_A_c_495_n N_Z_c_920_n 0.00270304f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_448 N_A_M1018_g N_Z_c_921_n 6.16809e-19 $X=7.755 $Y=2.465 $X2=0 $Y2=0
cc_449 N_A_M1025_g N_Z_c_921_n 8.98846e-19 $X=7.785 $Y=0.655 $X2=0 $Y2=0
cc_450 N_A_M1023_g N_Z_c_921_n 0.00373693f $X=8.185 $Y=2.465 $X2=0 $Y2=0
cc_451 N_A_M1029_g N_Z_c_921_n 0.00537963f $X=8.215 $Y=0.655 $X2=0 $Y2=0
cc_452 N_A_M1032_g N_Z_c_921_n 0.00323386f $X=8.615 $Y=2.465 $X2=0 $Y2=0
cc_453 N_A_M1031_g N_Z_c_921_n 0.0042563f $X=8.645 $Y=0.655 $X2=0 $Y2=0
cc_454 N_A_c_559_p N_Z_c_921_n 0.0200006f $X=7.82 $Y=1.49 $X2=0 $Y2=0
cc_455 N_A_c_495_n N_Z_c_921_n 0.0381556f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_456 N_A_M1003_g N_Z_c_929_n 0.00245936f $X=5.605 $Y=2.465 $X2=0 $Y2=0
cc_457 N_A_M1006_g N_Z_c_929_n 0.0134669f $X=6.035 $Y=2.465 $X2=0 $Y2=0
cc_458 N_A_M1009_g N_Z_c_929_n 0.00258592f $X=6.465 $Y=2.465 $X2=0 $Y2=0
cc_459 N_A_c_495_n N_Z_c_929_n 0.0174107f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_460 N_A_c_493_n N_Z_c_930_n 0.0161954f $X=7.053 $Y=1.402 $X2=0 $Y2=0
cc_461 N_A_c_495_n N_Z_c_930_n 0.00263158f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_462 N_A_M1015_g N_Z_c_922_n 9.88689e-19 $X=6.925 $Y=0.655 $X2=0 $Y2=0
cc_463 N_A_M1022_g N_Z_c_922_n 0.00551635f $X=7.355 $Y=0.655 $X2=0 $Y2=0
cc_464 N_A_M1025_g N_Z_c_922_n 2.17703e-19 $X=7.785 $Y=0.655 $X2=0 $Y2=0
cc_465 N_A_c_559_p N_Z_c_922_n 0.0197717f $X=7.82 $Y=1.49 $X2=0 $Y2=0
cc_466 N_A_c_495_n N_Z_c_922_n 0.00247501f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_467 N_A_c_559_p N_Z_c_931_n 0.015726f $X=7.82 $Y=1.49 $X2=0 $Y2=0
cc_468 N_A_c_495_n N_Z_c_931_n 0.00263158f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_469 N_A_M1029_g N_Z_c_923_n 0.00748259f $X=8.215 $Y=0.655 $X2=0 $Y2=0
cc_470 N_A_M1031_g N_Z_c_923_n 0.00317458f $X=8.645 $Y=0.655 $X2=0 $Y2=0
cc_471 N_A_M1023_g N_Z_c_932_n 0.00770792f $X=8.185 $Y=2.465 $X2=0 $Y2=0
cc_472 N_A_M1032_g N_Z_c_932_n 0.00185876f $X=8.615 $Y=2.465 $X2=0 $Y2=0
cc_473 N_A_M1002_g Z 0.001913f $X=5.635 $Y=0.655 $X2=0 $Y2=0
cc_474 N_A_M1008_g Z 0.0100286f $X=6.065 $Y=0.655 $X2=0 $Y2=0
cc_475 N_A_M1011_g Z 0.00141925f $X=6.495 $Y=0.655 $X2=0 $Y2=0
cc_476 N_A_c_493_n Z 0.0313361f $X=7.053 $Y=1.402 $X2=0 $Y2=0
cc_477 N_A_c_495_n Z 0.0189655f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_478 N_A_M1008_g N_Z_c_986_n 0.00533678f $X=6.065 $Y=0.655 $X2=0 $Y2=0
cc_479 N_A_M1002_g N_VGND_c_1042_n 0.00361998f $X=5.635 $Y=0.655 $X2=0 $Y2=0
cc_480 N_A_M1008_g N_VGND_c_1042_n 0.00362032f $X=6.065 $Y=0.655 $X2=0 $Y2=0
cc_481 N_A_M1011_g N_VGND_c_1042_n 0.00362032f $X=6.495 $Y=0.655 $X2=0 $Y2=0
cc_482 N_A_M1015_g N_VGND_c_1042_n 0.00362032f $X=6.925 $Y=0.655 $X2=0 $Y2=0
cc_483 N_A_M1022_g N_VGND_c_1042_n 0.00362032f $X=7.355 $Y=0.655 $X2=0 $Y2=0
cc_484 N_A_M1025_g N_VGND_c_1042_n 0.00363488f $X=7.785 $Y=0.655 $X2=0 $Y2=0
cc_485 N_A_M1029_g N_VGND_c_1042_n 0.00363488f $X=8.215 $Y=0.655 $X2=0 $Y2=0
cc_486 N_A_M1031_g N_VGND_c_1042_n 0.00362032f $X=8.645 $Y=0.655 $X2=0 $Y2=0
cc_487 N_A_M1002_g N_VGND_c_1043_n 0.00538087f $X=5.635 $Y=0.655 $X2=0 $Y2=0
cc_488 N_A_M1008_g N_VGND_c_1043_n 0.00541723f $X=6.065 $Y=0.655 $X2=0 $Y2=0
cc_489 N_A_M1011_g N_VGND_c_1043_n 0.00541723f $X=6.495 $Y=0.655 $X2=0 $Y2=0
cc_490 N_A_M1015_g N_VGND_c_1043_n 0.00541723f $X=6.925 $Y=0.655 $X2=0 $Y2=0
cc_491 N_A_M1022_g N_VGND_c_1043_n 0.00540811f $X=7.355 $Y=0.655 $X2=0 $Y2=0
cc_492 N_A_M1025_g N_VGND_c_1043_n 0.00534642f $X=7.785 $Y=0.655 $X2=0 $Y2=0
cc_493 N_A_M1029_g N_VGND_c_1043_n 0.00534642f $X=8.215 $Y=0.655 $X2=0 $Y2=0
cc_494 N_A_M1031_g N_VGND_c_1043_n 0.00642157f $X=8.645 $Y=0.655 $X2=0 $Y2=0
cc_495 N_A_M1002_g N_A_371_47#_c_1148_n 0.0024979f $X=5.635 $Y=0.655 $X2=0 $Y2=0
cc_496 N_A_c_495_n N_A_371_47#_c_1148_n 0.0055018f $X=8.645 $Y=1.49 $X2=0 $Y2=0
cc_497 N_A_M1002_g N_A_371_47#_c_1192_n 8.601e-19 $X=5.635 $Y=0.655 $X2=0 $Y2=0
cc_498 N_A_M1002_g N_A_371_47#_c_1193_n 0.0114023f $X=5.635 $Y=0.655 $X2=0 $Y2=0
cc_499 N_A_M1008_g N_A_371_47#_c_1193_n 9.59241e-19 $X=6.065 $Y=0.655 $X2=0
+ $Y2=0
cc_500 N_A_M1002_g N_A_371_47#_c_1204_n 0.0135568f $X=5.635 $Y=0.655 $X2=0 $Y2=0
cc_501 N_A_M1008_g N_A_371_47#_c_1204_n 0.0107175f $X=6.065 $Y=0.655 $X2=0 $Y2=0
cc_502 N_A_M1011_g N_A_371_47#_c_1204_n 0.0107232f $X=6.495 $Y=0.655 $X2=0 $Y2=0
cc_503 N_A_M1015_g N_A_371_47#_c_1204_n 0.0107232f $X=6.925 $Y=0.655 $X2=0 $Y2=0
cc_504 N_A_M1022_g N_A_371_47#_c_1204_n 0.0107086f $X=7.355 $Y=0.655 $X2=0 $Y2=0
cc_505 N_A_M1025_g N_A_371_47#_c_1204_n 0.0119073f $X=7.785 $Y=0.655 $X2=0 $Y2=0
cc_506 N_A_M1029_g N_A_371_47#_c_1210_n 0.00895842f $X=8.215 $Y=0.655 $X2=0
+ $Y2=0
cc_507 N_A_M1031_g N_A_371_47#_c_1210_n 0.0123718f $X=8.645 $Y=0.655 $X2=0 $Y2=0
cc_508 N_A_M1022_g N_A_371_47#_c_1212_n 8.95744e-19 $X=7.355 $Y=0.655 $X2=0
+ $Y2=0
cc_509 N_A_M1025_g N_A_371_47#_c_1212_n 0.0061282f $X=7.785 $Y=0.655 $X2=0 $Y2=0
cc_510 N_A_M1029_g N_A_371_47#_c_1212_n 0.00661712f $X=8.215 $Y=0.655 $X2=0
+ $Y2=0
cc_511 N_A_M1031_g N_A_371_47#_c_1212_n 5.83772e-19 $X=8.645 $Y=0.655 $X2=0
+ $Y2=0
cc_512 N_A_M1031_g N_A_371_47#_c_1152_n 0.00248138f $X=8.645 $Y=0.655 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_643_n N_A_365_367#_M1000_s 0.0026734f $X=8.88 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_514 N_VPWR_c_643_n N_A_365_367#_M1005_s 0.00293134f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_643_n N_A_365_367#_M1016_s 0.00293134f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_643_n N_A_365_367#_M1020_s 0.0027574f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_643_n N_A_365_367#_M1033_s 0.00254869f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_643_n N_A_365_367#_M1006_d 0.00223559f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_643_n N_A_365_367#_M1012_d 0.00223559f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_643_n N_A_365_367#_M1018_d 0.00223559f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_643_n N_A_365_367#_M1032_d 0.00215159f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_650_n N_A_365_367#_c_766_n 0.0188755f $X=2.245 $Y=3.33 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_643_n N_A_365_367#_c_766_n 0.0111968f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_645_n N_A_365_367#_c_758_n 0.0162354f $X=2.38 $Y=2.055 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_646_n N_A_365_367#_c_767_n 0.0149362f $X=3.105 $Y=3.33 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_643_n N_A_365_367#_c_767_n 0.0100304f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_647_n N_A_365_367#_c_760_n 0.0164056f $X=3.24 $Y=2.055 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_653_n N_A_365_367#_c_768_n 0.0149362f $X=3.97 $Y=3.33 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_643_n N_A_365_367#_c_768_n 0.0100304f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_648_n N_A_365_367#_c_761_n 0.0160651f $X=4.1 $Y=2.055 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_654_n N_A_365_367#_c_769_n 0.0151136f $X=4.83 $Y=3.33 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_643_n N_A_365_367#_c_769_n 0.0102248f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_649_n N_A_365_367#_c_762_n 0.0162354f $X=4.96 $Y=2.055 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_655_n N_A_365_367#_c_871_n 0.0148297f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_643_n N_A_365_367#_c_871_n 0.00990325f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_655_n N_A_365_367#_c_822_n 0.0319341f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_643_n N_A_365_367#_c_822_n 0.0201012f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_655_n N_A_365_367#_c_828_n 0.0298674f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_643_n N_A_365_367#_c_828_n 0.0187823f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_655_n N_A_365_367#_c_834_n 0.0298674f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_643_n N_A_365_367#_c_834_n 0.0187823f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_655_n N_A_365_367#_c_840_n 0.0319341f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_643_n N_A_365_367#_c_840_n 0.0201012f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_655_n N_A_365_367#_c_772_n 0.0189827f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_643_n N_A_365_367#_c_772_n 0.0112692f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_655_n N_A_365_367#_c_844_n 0.01906f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_547 N_VPWR_c_643_n N_A_365_367#_c_844_n 0.0124545f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_655_n N_A_365_367#_c_846_n 0.01906f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_549 N_VPWR_c_643_n N_A_365_367#_c_846_n 0.0124545f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_655_n N_A_365_367#_c_848_n 0.01906f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_551 N_VPWR_c_643_n N_A_365_367#_c_848_n 0.0124545f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_643_n N_Z_M1003_s 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_553 N_VPWR_c_643_n N_Z_M1009_s 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_554 N_VPWR_c_643_n N_Z_M1013_s 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_555 N_VPWR_c_643_n N_Z_M1023_s 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_556 N_A_365_367#_c_822_n N_Z_M1003_s 0.00332344f $X=6.085 $Y=2.99 $X2=0 $Y2=0
cc_557 N_A_365_367#_c_828_n N_Z_M1009_s 0.00332344f $X=6.945 $Y=2.99 $X2=0 $Y2=0
cc_558 N_A_365_367#_c_834_n N_Z_M1013_s 0.00332344f $X=7.805 $Y=2.99 $X2=0 $Y2=0
cc_559 N_A_365_367#_c_840_n N_Z_M1023_s 0.00332344f $X=8.705 $Y=2.99 $X2=0 $Y2=0
cc_560 N_A_365_367#_c_822_n N_Z_c_995_n 0.0126348f $X=6.085 $Y=2.99 $X2=0 $Y2=0
cc_561 N_A_365_367#_M1006_d N_Z_c_925_n 0.00176461f $X=6.11 $Y=1.835 $X2=0 $Y2=0
cc_562 N_A_365_367#_c_824_n N_Z_c_925_n 0.0152916f $X=6.25 $Y=2.19 $X2=0 $Y2=0
cc_563 N_A_365_367#_c_828_n N_Z_c_998_n 0.0126348f $X=6.945 $Y=2.99 $X2=0 $Y2=0
cc_564 N_A_365_367#_M1012_d N_Z_c_926_n 0.00176461f $X=6.97 $Y=1.835 $X2=0 $Y2=0
cc_565 N_A_365_367#_c_830_n N_Z_c_926_n 0.0170777f $X=7.11 $Y=2.19 $X2=0 $Y2=0
cc_566 N_A_365_367#_c_834_n N_Z_c_1001_n 0.0126348f $X=7.805 $Y=2.99 $X2=0 $Y2=0
cc_567 N_A_365_367#_M1018_d N_Z_c_927_n 0.00176461f $X=7.83 $Y=1.835 $X2=0 $Y2=0
cc_568 N_A_365_367#_c_836_n N_Z_c_927_n 0.0170777f $X=7.97 $Y=2.19 $X2=0 $Y2=0
cc_569 N_A_365_367#_c_840_n N_Z_c_1004_n 0.0126348f $X=8.705 $Y=2.99 $X2=0 $Y2=0
cc_570 N_A_365_367#_c_762_n N_Z_c_929_n 0.0148981f $X=5.26 $Y=1.635 $X2=0 $Y2=0
cc_571 N_A_365_367#_c_771_n N_Z_c_929_n 0.00947493f $X=5.39 $Y=1.98 $X2=0 $Y2=0
cc_572 N_A_365_367#_c_824_n N_Z_c_929_n 0.0019893f $X=6.25 $Y=2.19 $X2=0 $Y2=0
cc_573 N_A_365_367#_c_773_n N_Z_c_932_n 0.00166417f $X=8.83 $Y=1.98 $X2=0 $Y2=0
cc_574 N_A_365_367#_c_758_n N_A_371_47#_c_1141_n 0.0450506f $X=2.675 $Y=1.635
+ $X2=0 $Y2=0
cc_575 N_A_365_367#_c_763_n N_A_371_47#_c_1141_n 0.00587222f $X=2.805 $Y=1.635
+ $X2=0 $Y2=0
cc_576 N_A_365_367#_c_759_n N_A_371_47#_c_1142_n 0.0243534f $X=2.075 $Y=1.635
+ $X2=0 $Y2=0
cc_577 N_A_365_367#_c_760_n N_A_371_47#_c_1144_n 0.045427f $X=3.54 $Y=1.635
+ $X2=0 $Y2=0
cc_578 N_A_365_367#_c_764_n N_A_371_47#_c_1144_n 0.00545007f $X=3.67 $Y=1.635
+ $X2=0 $Y2=0
cc_579 N_A_365_367#_c_761_n N_A_371_47#_c_1146_n 0.0447119f $X=4.395 $Y=1.635
+ $X2=0 $Y2=0
cc_580 N_A_365_367#_c_764_n N_A_371_47#_c_1146_n 3.8435e-19 $X=3.67 $Y=1.635
+ $X2=0 $Y2=0
cc_581 N_A_365_367#_c_765_n N_A_371_47#_c_1146_n 0.00587222f $X=4.527 $Y=1.635
+ $X2=0 $Y2=0
cc_582 N_A_365_367#_c_762_n N_A_371_47#_c_1148_n 0.0671071f $X=5.26 $Y=1.635
+ $X2=0 $Y2=0
cc_583 N_A_365_367#_c_763_n N_A_371_47#_c_1149_n 0.017796f $X=2.805 $Y=1.635
+ $X2=0 $Y2=0
cc_584 N_A_365_367#_c_764_n N_A_371_47#_c_1150_n 0.017796f $X=3.67 $Y=1.635
+ $X2=0 $Y2=0
cc_585 N_A_365_367#_c_762_n N_A_371_47#_c_1151_n 0.00207293f $X=5.26 $Y=1.635
+ $X2=0 $Y2=0
cc_586 N_A_365_367#_c_765_n N_A_371_47#_c_1151_n 0.0182643f $X=4.527 $Y=1.635
+ $X2=0 $Y2=0
cc_587 N_Z_M1002_s N_VGND_c_1043_n 0.00225919f $X=5.71 $Y=0.235 $X2=0 $Y2=0
cc_588 N_Z_M1011_s N_VGND_c_1043_n 0.00225919f $X=6.57 $Y=0.235 $X2=0 $Y2=0
cc_589 N_Z_M1022_s N_VGND_c_1043_n 0.00225919f $X=7.43 $Y=0.235 $X2=0 $Y2=0
cc_590 N_Z_M1029_s N_VGND_c_1043_n 0.00225919f $X=8.29 $Y=0.235 $X2=0 $Y2=0
cc_591 N_Z_c_933_n N_A_371_47#_M1008_d 0.004731f $X=7.415 $Y=0.86 $X2=0 $Y2=0
cc_592 N_Z_c_933_n N_A_371_47#_M1015_d 0.00353077f $X=7.415 $Y=0.86 $X2=0 $Y2=0
cc_593 N_Z_c_920_n N_A_371_47#_M1025_d 0.00180746f $X=8.155 $Y=1.09 $X2=0 $Y2=0
cc_594 Z N_A_371_47#_c_1148_n 0.0141176f $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_595 Z N_A_371_47#_c_1193_n 0.0137022f $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_596 N_Z_M1002_s N_A_371_47#_c_1204_n 0.00344536f $X=5.71 $Y=0.235 $X2=0 $Y2=0
cc_597 N_Z_M1011_s N_A_371_47#_c_1204_n 0.00344973f $X=6.57 $Y=0.235 $X2=0 $Y2=0
cc_598 N_Z_M1022_s N_A_371_47#_c_1204_n 0.00344536f $X=7.43 $Y=0.235 $X2=0 $Y2=0
cc_599 N_Z_c_933_n N_A_371_47#_c_1204_n 0.0687437f $X=7.415 $Y=0.86 $X2=0 $Y2=0
cc_600 N_Z_c_920_n N_A_371_47#_c_1204_n 0.00398821f $X=8.155 $Y=1.09 $X2=0 $Y2=0
cc_601 N_Z_c_922_n N_A_371_47#_c_1204_n 0.013996f $X=7.54 $Y=0.86 $X2=0 $Y2=0
cc_602 N_Z_c_986_n N_A_371_47#_c_1204_n 0.0235983f $X=5.94 $Y=0.995 $X2=0 $Y2=0
cc_603 N_Z_M1029_s N_A_371_47#_c_1210_n 0.00339264f $X=8.29 $Y=0.235 $X2=0 $Y2=0
cc_604 N_Z_c_1026_p N_A_371_47#_c_1210_n 0.0126887f $X=8.43 $Y=0.78 $X2=0 $Y2=0
cc_605 N_Z_c_923_n N_A_371_47#_c_1210_n 0.00356188f $X=8.357 $Y=1.09 $X2=0 $Y2=0
cc_606 N_Z_c_920_n N_A_371_47#_c_1212_n 0.0153958f $X=8.155 $Y=1.09 $X2=0 $Y2=0
cc_607 N_Z_c_923_n N_A_371_47#_c_1212_n 7.1577e-19 $X=8.357 $Y=1.09 $X2=0 $Y2=0
cc_608 N_Z_c_923_n N_A_371_47#_c_1152_n 0.00166618f $X=8.357 $Y=1.09 $X2=0 $Y2=0
cc_609 N_VGND_c_1043_n N_A_371_47#_M1001_s 0.00371702f $X=8.88 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_610 N_VGND_c_1043_n N_A_371_47#_M1004_s 0.00536646f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_c_1043_n N_A_371_47#_M1014_s 0.00536646f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_612 N_VGND_c_1043_n N_A_371_47#_M1024_s 0.00432284f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_613 N_VGND_c_1043_n N_A_371_47#_M1030_s 0.00224253f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_c_1043_n N_A_371_47#_M1008_d 0.00224306f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_615 N_VGND_c_1043_n N_A_371_47#_M1015_d 0.00224306f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_616 N_VGND_c_1043_n N_A_371_47#_M1025_d 0.00224253f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_617 N_VGND_c_1043_n N_A_371_47#_M1031_d 0.00215819f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_618 N_VGND_c_1037_n N_A_371_47#_c_1140_n 0.0178111f $X=2.245 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_c_1043_n N_A_371_47#_c_1140_n 0.0100304f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_620 N_VGND_c_1032_n N_A_371_47#_c_1141_n 0.0204885f $X=2.41 $Y=0.38 $X2=0
+ $Y2=0
cc_621 N_VGND_c_1033_n N_A_371_47#_c_1143_n 0.0124525f $X=3.105 $Y=0 $X2=0 $Y2=0
cc_622 N_VGND_c_1043_n N_A_371_47#_c_1143_n 0.00730901f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_623 N_VGND_c_1034_n N_A_371_47#_c_1144_n 0.0204885f $X=3.27 $Y=0.38 $X2=0
+ $Y2=0
cc_624 N_VGND_c_1040_n N_A_371_47#_c_1145_n 0.0124525f $X=3.965 $Y=0 $X2=0 $Y2=0
cc_625 N_VGND_c_1043_n N_A_371_47#_c_1145_n 0.00730901f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_626 N_VGND_c_1035_n N_A_371_47#_c_1146_n 0.0204885f $X=4.13 $Y=0.38 $X2=0
+ $Y2=0
cc_627 N_VGND_c_1041_n N_A_371_47#_c_1147_n 0.0135169f $X=4.855 $Y=0 $X2=0 $Y2=0
cc_628 N_VGND_c_1043_n N_A_371_47#_c_1147_n 0.00847534f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_629 N_VGND_c_1036_n N_A_371_47#_c_1148_n 0.0152138f $X=4.99 $Y=0.36 $X2=0
+ $Y2=0
cc_630 N_VGND_c_1042_n N_A_371_47#_c_1192_n 0.0169136f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_631 N_VGND_c_1043_n N_A_371_47#_c_1192_n 0.0123294f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_632 N_VGND_c_1042_n N_A_371_47#_c_1204_n 0.113988f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_633 N_VGND_c_1043_n N_A_371_47#_c_1204_n 0.0803546f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_634 N_VGND_c_1042_n N_A_371_47#_c_1210_n 0.0282056f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_635 N_VGND_c_1043_n N_A_371_47#_c_1210_n 0.0196468f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_636 N_VGND_c_1042_n N_A_371_47#_c_1212_n 0.0165945f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_637 N_VGND_c_1043_n N_A_371_47#_c_1212_n 0.0121884f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_638 N_VGND_c_1042_n N_A_371_47#_c_1152_n 0.0169934f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_639 N_VGND_c_1043_n N_A_371_47#_c_1152_n 0.0113583f $X=8.88 $Y=0 $X2=0 $Y2=0
