* NGSPICE file created from sky130_fd_sc_lp__and4_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and4_2 A B C D VGND VNB VPB VPWR X
M1000 VPWR D a_72_49# VPB phighvt w=420000u l=150000u
+  ad=1.1067e+12p pd=9.87e+06u as=2.352e+11p ps=2.8e+06u
M1001 a_335_49# C a_227_49# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.638e+11p ps=1.62e+06u
M1002 X a_72_49# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=5.922e+11p ps=5.12e+06u
M1003 VPWR B a_72_49# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_72_49# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1005 a_72_49# C VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND D a_335_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_227_49# B a_155_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1008 VGND a_72_49# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_72_49# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_155_49# A a_72_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 VPWR a_72_49# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

