* File: sky130_fd_sc_lp__clkbuflp_2.spice
* Created: Fri Aug 28 10:15:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkbuflp_2.pex.spice"
.subckt sky130_fd_sc_lp__clkbuflp_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 A_110_47# N_A_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g A_110_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1000_d N_A_27_47#_M1005_g A_268_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 A_268_47# N_A_27_47#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1006 A_426_47# N_A_27_47#_M1006_g N_X_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_27_47#_M1007_g A_426_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1002 N_VPWR_M1001_d N_A_27_47#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_A_27_47#_M1008_g N_X_M1002_s VPB PHIGHVT L=0.25 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX9_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__clkbuflp_2.pxi.spice"
*
.ends
*
*
