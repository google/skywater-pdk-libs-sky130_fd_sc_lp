* File: sky130_fd_sc_lp__xnor2_lp.pex.spice
* Created: Fri Aug 28 11:35:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XNOR2_LP%A_82_66# 1 2 9 13 15 21 22 23 26 28 31 32
+ 34 40
c79 40 0 1.28604e-19 $X=0.745 $Y=1.63
r80 34 36 10.6092 $w=3.53e-07 $l=2.3e-07 $layer=LI1_cond $X=3.092 $Y=0.835
+ $X2=3.092 $Y2=1.065
r81 31 36 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.185 $Y=2.02
+ $X2=3.185 $Y2=1.065
r82 29 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=2.105
+ $X2=2.56 $Y2=2.105
r83 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.105
+ $X2=3.185 $Y2=2.02
r84 28 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.1 $Y=2.105
+ $X2=2.725 $Y2=2.105
r85 24 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=2.19 $X2=2.56
+ $Y2=2.105
r86 24 26 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.56 $Y=2.19 $X2=2.56
+ $Y2=2.24
r87 22 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=2.105
+ $X2=2.56 $Y2=2.105
r88 22 23 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.395 $Y=2.105
+ $X2=1.525 $Y2=2.105
r89 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.44 $Y=2.02
+ $X2=1.525 $Y2=2.105
r90 20 21 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.44 $Y=1.795
+ $X2=1.44 $Y2=2.02
r91 18 40 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.705 $Y=1.63
+ $X2=0.745 $Y2=1.63
r92 18 37 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.705 $Y=1.63
+ $X2=0.485 $Y2=1.63
r93 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.705
+ $Y=1.63 $X2=0.705 $Y2=1.63
r94 15 20 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.355 $Y=1.63
+ $X2=1.44 $Y2=1.795
r95 15 17 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=1.355 $Y=1.63
+ $X2=0.705 $Y2=1.63
r96 11 40 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.745 $Y=1.795
+ $X2=0.745 $Y2=1.63
r97 11 13 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=0.745 $Y=1.795
+ $X2=0.745 $Y2=2.595
r98 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.465
+ $X2=0.485 $Y2=1.63
r99 7 9 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.485 $Y=1.465
+ $X2=0.485 $Y2=0.67
r100 2 26 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.42
+ $Y=2.095 $X2=2.56 $Y2=2.24
r101 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.625 $X2=3.08 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_LP%A 3 5 7 10 12 14 15 21 22
c51 21 0 1.29497e-20 $X=2.18 $Y=1.41
c52 5 0 1.46822e-19 $X=2.045 $Y=1.12
c53 3 0 8.55262e-20 $X=1.765 $Y=2.595
r54 20 22 13.7203 $w=4.04e-07 $l=1.15e-07 $layer=POLY_cond $X=2.18 $Y=1.41
+ $X2=2.295 $Y2=1.41
r55 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.18
+ $Y=1.41 $X2=2.18 $Y2=1.41
r56 18 20 16.1064 $w=4.04e-07 $l=1.35e-07 $layer=POLY_cond $X=2.045 $Y=1.41
+ $X2=2.18 $Y2=1.41
r57 17 18 33.4059 $w=4.04e-07 $l=2.8e-07 $layer=POLY_cond $X=1.765 $Y=1.41
+ $X2=2.045 $Y2=1.41
r58 15 21 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.18 $Y=1.665
+ $X2=2.18 $Y2=1.41
r59 12 22 21.4752 $w=4.04e-07 $l=3.69188e-07 $layer=POLY_cond $X=2.475 $Y=1.12
+ $X2=2.295 $Y2=1.41
r60 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.475 $Y=1.12
+ $X2=2.475 $Y2=0.835
r61 8 22 14.0064 $w=2.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.295 $Y=1.7
+ $X2=2.295 $Y2=1.41
r62 8 10 222.366 $w=2.5e-07 $l=8.95e-07 $layer=POLY_cond $X=2.295 $Y=1.7
+ $X2=2.295 $Y2=2.595
r63 5 18 26.1054 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.045 $Y=1.12
+ $X2=2.045 $Y2=1.41
r64 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.045 $Y=1.12 $X2=2.045
+ $Y2=0.835
r65 1 17 14.0064 $w=2.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.765 $Y=1.7
+ $X2=1.765 $Y2=1.41
r66 1 3 222.366 $w=2.5e-07 $l=8.95e-07 $layer=POLY_cond $X=1.765 $Y=1.7
+ $X2=1.765 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_LP%B 3 8 9 10 13 18 21 23 26 27
c71 21 0 1.29497e-20 $X=1.455 $Y=1.195
r72 26 29 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.675
+ $X2=2.795 $Y2=1.84
r73 26 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.675
+ $X2=2.795 $Y2=1.51
r74 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.795
+ $Y=1.675 $X2=2.795 $Y2=1.675
r75 23 27 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.64 $Y=1.675
+ $X2=2.795 $Y2=1.675
r76 18 28 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.865 $Y=0.835
+ $X2=2.865 $Y2=1.51
r77 15 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.865 $Y=0.255
+ $X2=2.865 $Y2=0.835
r78 13 29 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.825 $Y=2.595
+ $X2=2.825 $Y2=1.84
r79 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.79 $Y=0.18
+ $X2=2.865 $Y2=0.255
r80 9 10 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=2.79 $Y=0.18
+ $X2=1.53 $Y2=0.18
r81 6 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.455 $Y=1.12
+ $X2=1.455 $Y2=1.195
r82 6 8 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.455 $Y=1.12
+ $X2=1.455 $Y2=0.835
r83 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.455 $Y=0.255
+ $X2=1.53 $Y2=0.18
r84 5 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.455 $Y=0.255
+ $X2=1.455 $Y2=0.835
r85 1 21 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.275 $Y=1.195
+ $X2=1.455 $Y2=1.195
r86 1 3 329.201 $w=2.5e-07 $l=1.325e-06 $layer=POLY_cond $X=1.275 $Y=1.27
+ $X2=1.275 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_LP%VPWR 1 2 3 12 16 18 20 23 24 26 27 28 40 46
r47 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 40 45 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=3.142 $Y2=3.33
r51 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r53 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 32 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 28 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 28 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 28 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 26 38 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=2.03 $Y2=3.33
r61 25 42 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.03 $Y2=3.33
r63 23 31 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.315 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.315 $Y=3.33
+ $X2=0.48 $Y2=3.33
r65 22 35 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=0.48 $Y2=3.33
r67 18 45 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.09 $Y=3.245
+ $X2=3.142 $Y2=3.33
r68 18 20 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.09 $Y=3.245
+ $X2=3.09 $Y2=2.535
r69 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=3.33
r70 14 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=2.535
r71 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.48 $Y=3.245
+ $X2=0.48 $Y2=3.33
r72 10 12 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.48 $Y=3.245
+ $X2=0.48 $Y2=2.49
r73 3 20 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=2.95
+ $Y=2.095 $X2=3.09 $Y2=2.535
r74 2 16 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=1.89
+ $Y=2.095 $X2=2.03 $Y2=2.535
r75 1 12 300 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=2 $X=0.335
+ $Y=2.095 $X2=0.48 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_LP%Y 1 2 7 8 11 14 15 16 17 25
c32 7 0 8.55262e-20 $X=0.845 $Y=2.06
r33 25 37 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=0.23 $Y=0.925
+ $X2=0.23 $Y2=0.9
r34 16 17 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.665
r35 15 37 1.75234 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.27 $Y=0.87 $X2=0.27
+ $Y2=0.9
r36 15 35 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=0.87 $X2=0.27
+ $Y2=0.67
r37 15 16 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.23 $Y=0.955
+ $X2=0.23 $Y2=1.295
r38 15 25 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.955 $X2=0.23
+ $Y2=0.925
r39 14 35 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.27 $Y=0.555
+ $X2=0.27 $Y2=0.67
r40 13 17 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.23 $Y=1.975
+ $X2=0.23 $Y2=1.665
r41 9 11 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.01 $Y=2.145
+ $X2=1.01 $Y2=2.24
r42 8 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.355 $Y=2.06
+ $X2=0.23 $Y2=1.975
r43 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.845 $Y=2.06
+ $X2=1.01 $Y2=2.145
r44 7 8 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=0.845 $Y=2.06
+ $X2=0.355 $Y2=2.06
r45 2 11 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.87
+ $Y=2.095 $X2=1.01 $Y2=2.24
r46 1 35 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.46 $X2=0.27 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_LP%A_112_92# 1 2 9 11 12 15
c29 11 0 2.75425e-19 $X=1.585 $Y=1.2
r30 13 15 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.71 $Y=1.115
+ $X2=1.71 $Y2=0.835
r31 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.585 $Y=1.2
+ $X2=1.71 $Y2=1.115
r32 11 12 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.585 $Y=1.2
+ $X2=0.865 $Y2=1.2
r33 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.74 $Y=1.115
+ $X2=0.865 $Y2=1.2
r34 7 9 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.74 $Y=1.115
+ $X2=0.74 $Y2=0.67
r35 2 15 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.625 $X2=1.75 $Y2=0.835
r36 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.46 $X2=0.7 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_LP%VGND 1 2 9 11 15 17 19 26 27 30 33
r41 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 27 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r44 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 24 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.22
+ $Y2=0
r46 24 26 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=3.12
+ $Y2=0
r47 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r48 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=1.24
+ $Y2=0
r50 19 21 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=0.72
+ $Y2=0
r51 17 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r52 17 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r53 13 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=0.085
+ $X2=2.22 $Y2=0
r54 13 15 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=2.22 $Y=0.085
+ $X2=2.22 $Y2=0.835
r55 12 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.24
+ $Y2=0
r56 11 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.22
+ $Y2=0
r57 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=1.405
+ $Y2=0
r58 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=0.085 $X2=1.24
+ $Y2=0
r59 7 9 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=1.24 $Y=0.085
+ $X2=1.24 $Y2=0.77
r60 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.625 $X2=2.26 $Y2=0.835
r61 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.105
+ $Y=0.625 $X2=1.24 $Y2=0.77
.ends

