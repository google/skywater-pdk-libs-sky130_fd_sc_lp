* File: sky130_fd_sc_lp__iso1n_lp.pex.spice
* Created: Wed Sep  2 09:58:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__ISO1N_LP%SLEEP_B 3 7 11 15 17 18 25
c42 17 0 4.31101e-21 $X=0.75 $Y=1.295
c43 11 0 3.94423e-21 $X=0.835 $Y=0.675
r44 25 27 7.13487 $w=6.08e-07 $l=9e-08 $layer=POLY_cond $X=0.995 $Y=1.655
+ $X2=1.085 $Y2=1.655
r45 25 26 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=0.995
+ $Y=1.485 $X2=0.995 $Y2=1.485
r46 23 25 12.6842 $w=6.08e-07 $l=1.6e-07 $layer=POLY_cond $X=0.835 $Y=1.655
+ $X2=0.995 $Y2=1.655
r47 22 23 11.0987 $w=6.08e-07 $l=1.4e-07 $layer=POLY_cond $X=0.695 $Y=1.655
+ $X2=0.835 $Y2=1.655
r48 18 26 3.47249 $w=6.18e-07 $l=1.8e-07 $layer=LI1_cond $X=0.85 $Y=1.665
+ $X2=0.85 $Y2=1.485
r49 17 26 3.6654 $w=6.18e-07 $l=1.9e-07 $layer=LI1_cond $X=0.85 $Y=1.295
+ $X2=0.85 $Y2=1.485
r50 13 27 36.4184 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.085 $Y=1.99
+ $X2=1.085 $Y2=1.655
r51 13 15 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=1.085 $Y=1.99
+ $X2=1.085 $Y2=2.655
r52 9 23 36.4184 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.835 $Y=1.32
+ $X2=0.835 $Y2=1.655
r53 9 11 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.835 $Y=1.32
+ $X2=0.835 $Y2=0.675
r54 5 22 36.4184 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.695 $Y=1.99
+ $X2=0.695 $Y2=1.655
r55 5 7 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=0.695 $Y=1.99
+ $X2=0.695 $Y2=2.655
r56 1 22 17.4408 $w=6.08e-07 $l=4.3119e-07 $layer=POLY_cond $X=0.475 $Y=1.32
+ $X2=0.695 $Y2=1.655
r57 1 3 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.475 $Y=1.32
+ $X2=0.475 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP%A_27_93# 1 2 7 9 10 12 15 21 24 25 29 32 34
+ 35 38 39
c66 38 0 3.94423e-21 $X=1.535 $Y=1.48
c67 15 0 4.31101e-21 $X=1.625 $Y=2.655
r68 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.535
+ $Y=1.48 $X2=1.535 $Y2=1.48
r69 36 38 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.535 $Y=2.16
+ $X2=1.535 $Y2=1.48
r70 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.37 $Y=2.245
+ $X2=1.535 $Y2=2.16
r71 34 35 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.37 $Y=2.245
+ $X2=0.59 $Y2=2.245
r72 30 35 8.0246 $w=1.68e-07 $l=1.23e-07 $layer=LI1_cond $X=0.467 $Y=2.245
+ $X2=0.59 $Y2=2.245
r73 30 32 15.2875 $w=2.43e-07 $l=3.25e-07 $layer=LI1_cond $X=0.467 $Y=2.33
+ $X2=0.467 $Y2=2.655
r74 29 30 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.247 $Y=2.245
+ $X2=0.467 $Y2=2.245
r75 28 29 54.2354 $w=2.43e-07 $l=1.153e-06 $layer=LI1_cond $X=0.247 $Y=1.007
+ $X2=0.247 $Y2=2.16
r76 25 28 12.1502 $w=2.45e-07 $l=2.46487e-07 $layer=LI1_cond $X=0.242 $Y=0.763
+ $X2=0.247 $Y2=1.007
r77 25 27 2.14122 $w=2.45e-07 $l=4.3e-08 $layer=LI1_cond $X=0.242 $Y=0.763
+ $X2=0.242 $Y2=0.72
r78 23 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.535 $Y=1.82
+ $X2=1.535 $Y2=1.48
r79 23 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.535 $Y=1.82
+ $X2=1.535 $Y2=1.985
r80 20 39 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=1.535 $Y=1.11
+ $X2=1.535 $Y2=1.48
r81 20 21 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.535 $Y=1.035
+ $X2=1.625 $Y2=1.035
r82 17 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.265 $Y=1.035
+ $X2=1.535 $Y2=1.035
r83 15 24 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.625 $Y=2.655
+ $X2=1.625 $Y2=1.985
r84 10 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.625 $Y=0.96
+ $X2=1.625 $Y2=1.035
r85 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.625 $Y=0.96
+ $X2=1.625 $Y2=0.675
r86 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.265 $Y=0.96
+ $X2=1.265 $Y2=1.035
r87 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.265 $Y=0.96 $X2=1.265
+ $Y2=0.675
r88 2 32 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=2.445 $X2=0.48 $Y2=2.655
r89 1 27 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP%A 3 7 11 13 20 21
c46 20 0 8.05229e-20 $X=2.415 $Y=1.48
r47 19 21 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.415 $Y=1.48
+ $X2=2.475 $Y2=1.48
r48 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.415
+ $Y=1.48 $X2=2.415 $Y2=1.48
r49 17 19 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.115 $Y=1.48
+ $X2=2.415 $Y2=1.48
r50 15 17 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.985 $Y=1.48
+ $X2=2.115 $Y2=1.48
r51 13 20 3.3026 $w=6.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.245 $Y=1.665
+ $X2=2.245 $Y2=1.48
r52 9 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.475 $Y=1.315
+ $X2=2.475 $Y2=1.48
r53 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.475 $Y=1.315
+ $X2=2.475 $Y2=0.675
r54 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.115 $Y=1.315
+ $X2=2.115 $Y2=1.48
r55 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.115 $Y=1.315
+ $X2=2.115 $Y2=0.675
r56 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=1.645
+ $X2=1.985 $Y2=1.48
r57 1 3 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.985 $Y=1.645
+ $X2=1.985 $Y2=2.655
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP%A_340_93# 1 2 7 9 12 14 16 19 22 23 24 27
+ 29 30 31 32 34 39
r75 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.06
+ $Y=1.17 $X2=3.06 $Y2=1.17
r76 34 36 7.84973 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.9 $Y=0.715 $X2=1.9
+ $Y2=0.885
r77 31 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=1.225 $X2=3.06
+ $Y2=1.14
r78 31 32 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=3.06 $Y=1.225
+ $X2=3.06 $Y2=1.955
r79 29 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.895 $Y=2.04
+ $X2=3.06 $Y2=1.955
r80 29 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.895 $Y=2.04
+ $X2=2.305 $Y2=2.04
r81 25 30 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.2 $Y=2.125
+ $X2=2.305 $Y2=2.04
r82 25 27 30.1039 $w=2.08e-07 $l=5.7e-07 $layer=LI1_cond $X=2.2 $Y=2.125 $X2=2.2
+ $Y2=2.695
r83 23 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=1.14
+ $X2=3.06 $Y2=1.14
r84 23 24 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.895 $Y=1.14
+ $X2=2.065 $Y2=1.14
r85 22 24 6.85817 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=1.967 $Y=1.055
+ $X2=2.065 $Y2=1.14
r86 22 36 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=1.967 $Y=1.055
+ $X2=1.967 $Y2=0.885
r87 17 39 100.035 $w=2.55e-07 $l=6.03324e-07 $layer=POLY_cond $X=3.295 $Y=1.69
+ $X2=3.115 $Y2=1.17
r88 17 19 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=3.295 $Y=1.69
+ $X2=3.295 $Y2=2.465
r89 14 39 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=3.295 $Y=1.005
+ $X2=3.115 $Y2=1.17
r90 14 16 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.295 $Y=1.005
+ $X2=3.295 $Y2=0.675
r91 10 39 100.035 $w=2.55e-07 $l=6.03324e-07 $layer=POLY_cond $X=2.935 $Y=1.69
+ $X2=3.115 $Y2=1.17
r92 10 12 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=2.935 $Y=1.69
+ $X2=2.935 $Y2=2.465
r93 7 39 32.933 $w=2.55e-07 $l=1.8e-07 $layer=POLY_cond $X=2.935 $Y=1.17
+ $X2=3.115 $Y2=1.17
r94 7 9 106.04 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.935 $Y=1.17
+ $X2=2.935 $Y2=0.675
r95 2 27 600 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=2.06
+ $Y=2.445 $X2=2.2 $Y2=2.695
r96 1 34 182 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.465 $X2=1.9 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP%VPWR 1 2 9 13 15 17 22 29 30 33 36
r40 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 27 36 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.91 $Y=3.33
+ $X2=2.717 $Y2=3.33
r45 27 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.91 $Y=3.33 $X2=3.6
+ $Y2=3.33
r46 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=3.33
+ $X2=1.355 $Y2=3.33
r49 23 25 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.52 $Y=3.33 $X2=2.16
+ $Y2=3.33
r50 22 36 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.717 $Y2=3.33
r51 22 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 20 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=3.33
+ $X2=1.355 $Y2=3.33
r55 17 19 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=1.19 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 11 36 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.717 $Y=3.245
+ $X2=2.717 $Y2=3.33
r59 11 13 25.8926 $w=3.83e-07 $l=8.65e-07 $layer=LI1_cond $X=2.717 $Y=3.245
+ $X2=2.717 $Y2=2.38
r60 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=3.33
r61 7 9 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=2.655
r62 2 13 300 $w=1.7e-07 $l=6.04276e-07 $layer=licon1_PDIFF $count=2 $X=2.595
+ $Y=1.835 $X2=2.72 $Y2=2.38
r63 1 9 600 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=2.445 $X2=1.355 $Y2=2.655
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP%X 1 2 7 8 9 10 11 18
r13 11 33 16.1662 $w=3.58e-07 $l=5.05e-07 $layer=LI1_cond $X=3.575 $Y=2.405
+ $X2=3.575 $Y2=2.91
r14 10 11 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.575 $Y=2.035
+ $X2=3.575 $Y2=2.405
r15 10 27 1.76068 $w=3.58e-07 $l=5.5e-08 $layer=LI1_cond $X=3.575 $Y=2.035
+ $X2=3.575 $Y2=1.98
r16 9 27 10.0839 $w=3.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.575 $Y=1.665
+ $X2=3.575 $Y2=1.98
r17 8 9 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.575 $Y=1.295
+ $X2=3.575 $Y2=1.665
r18 7 8 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.575 $Y=0.925
+ $X2=3.575 $Y2=1.295
r19 7 18 6.56252 $w=3.58e-07 $l=2.05e-07 $layer=LI1_cond $X=3.575 $Y=0.925
+ $X2=3.575 $Y2=0.72
r20 2 33 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=1.835 $X2=3.51 $Y2=2.91
r21 2 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=1.835 $X2=3.51 $Y2=1.98
r22 1 18 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.465 $X2=3.51 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP%KAGND 1 2 7 10 17 18
r49 17 21 3.13259 $w=6.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=0.555
+ $X2=2.84 $Y2=0.72
r50 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.02 $Y=0.555
+ $X2=3.02 $Y2=0.555
r51 10 14 2.94273 $w=6.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=0.555
+ $X2=1.2 $Y2=0.71
r52 10 11 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.38 $Y=0.555
+ $X2=1.38 $Y2=0.555
r53 7 18 0.705765 $w=2.3e-07 $l=1.1e-06 $layer=MET1_cond $X=1.92 $Y=0.555
+ $X2=3.02 $Y2=0.555
r54 7 11 0.346466 $w=2.3e-07 $l=5.4e-07 $layer=MET1_cond $X=1.92 $Y=0.555
+ $X2=1.38 $Y2=0.555
r55 2 21 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.465 $X2=2.69 $Y2=0.72
r56 1 14 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.465 $X2=1.05 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP%VGND 1 5 8 15
r30 5 8 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r31 4 8 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r32 4 5 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 1 15 9.76563e-05 $w=3.84e-06 $l=3e-09 $layer=MET1_cond $X=1.92 $Y=0.122
+ $X2=1.92 $Y2=0.125
r34 1 5 0.00397135 $w=3.84e-06 $l=1.22e-07 $layer=MET1_cond $X=1.92 $Y=0.122
+ $X2=1.92 $Y2=0
.ends

