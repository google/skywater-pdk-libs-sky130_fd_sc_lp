# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a2111oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a2111oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465000 1.345000 4.185000 1.615000 ;
        RECT 3.465000 1.615000 5.155000 1.785000 ;
        RECT 4.895000 1.345000 5.155000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 1.210000 4.725000 1.435000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065000 1.425000 2.855000 1.775000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.295000 0.455000 1.605000 ;
        RECT 0.125000 1.605000 1.895000 1.775000 ;
        RECT 1.525000 1.295000 1.895000 1.605000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.210000 1.355000 1.435000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.541400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.255000 0.380000 0.870000 ;
        RECT 0.120000 0.870000 2.295000 1.040000 ;
        RECT 1.000000 1.945000 3.295000 1.955000 ;
        RECT 1.000000 1.955000 5.660000 2.125000 ;
        RECT 1.000000 2.125000 1.265000 2.355000 ;
        RECT 1.050000 0.265000 1.295000 0.870000 ;
        RECT 1.965000 0.255000 2.295000 0.870000 ;
        RECT 2.065000 1.040000 2.295000 1.085000 ;
        RECT 2.065000 1.085000 3.295000 1.255000 ;
        RECT 2.965000 0.255000 3.295000 1.085000 ;
        RECT 3.025000 1.255000 3.295000 1.945000 ;
        RECT 5.020000 0.255000 5.660000 1.095000 ;
        RECT 5.325000 1.095000 5.660000 1.955000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.120000  1.955000 0.400000 2.865000 ;
      RECT 0.120000  2.865000 3.070000 3.075000 ;
      RECT 0.550000  0.085000 0.880000 0.700000 ;
      RECT 0.570000  1.955000 0.830000 2.525000 ;
      RECT 0.570000  2.525000 1.700000 2.695000 ;
      RECT 1.450000  2.295000 1.700000 2.525000 ;
      RECT 1.465000  0.085000 1.795000 0.700000 ;
      RECT 1.870000  2.295000 2.165000 2.815000 ;
      RECT 1.870000  2.815000 3.070000 2.865000 ;
      RECT 2.335000  2.295000 5.350000 2.465000 ;
      RECT 2.335000  2.465000 3.520000 2.645000 ;
      RECT 2.465000  0.085000 2.795000 0.915000 ;
      RECT 3.260000  2.645000 3.520000 3.075000 ;
      RECT 3.530000  0.255000 3.860000 0.870000 ;
      RECT 3.530000  0.870000 4.850000 1.040000 ;
      RECT 3.690000  2.635000 4.020000 3.245000 ;
      RECT 4.125000  0.085000 4.455000 0.700000 ;
      RECT 4.190000  2.465000 4.400000 3.075000 ;
      RECT 4.570000  2.635000 4.900000 3.245000 ;
      RECT 4.625000  0.255000 4.850000 0.870000 ;
      RECT 5.070000  2.465000 5.350000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__a2111oi_2
