* File: sky130_fd_sc_lp__a2111oi_0.pex.spice
* Created: Wed Sep  2 09:16:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111OI_0%D1 2 3 4 5 6 9 11 13 16 17 18 19 20 26
r39 19 20 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=2.035
r40 18 19 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r41 17 18 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r42 17 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r43 15 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.005
r44 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.51
r45 14 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.99
+ $X2=0.27 $Y2=1.005
r46 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.795 $Y=2.29
+ $X2=0.795 $Y2=2.735
r47 7 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.725 $Y=0.84
+ $X2=0.725 $Y2=0.445
r48 5 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.72 $Y=2.215
+ $X2=0.795 $Y2=2.29
r49 5 6 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.72 $Y=2.215
+ $X2=0.435 $Y2=2.215
r50 4 14 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=0.915
+ $X2=0.27 $Y2=0.99
r51 3 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.65 $Y=0.915
+ $X2=0.725 $Y2=0.84
r52 3 4 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.65 $Y=0.915
+ $X2=0.435 $Y2=0.915
r53 2 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.36 $Y=2.14
+ $X2=0.435 $Y2=2.215
r54 2 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.36 $Y=2.14 $X2=0.36
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_0%C1 3 7 11 12 13 14 15 16 17 24
c44 7 0 1.52116e-19 $X=1.155 $Y=2.735
r45 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.065
+ $Y=1.395 $X2=1.065 $Y2=1.395
r46 16 17 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.165 $Y=2.405
+ $X2=1.165 $Y2=2.775
r47 15 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.165 $Y=2.035
+ $X2=1.165 $Y2=2.405
r48 14 15 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.165 $Y=1.665
+ $X2=1.165 $Y2=2.035
r49 14 25 8.40972 $w=3.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.165 $Y=1.665
+ $X2=1.165 $Y2=1.395
r50 13 25 3.11471 $w=3.68e-07 $l=1e-07 $layer=LI1_cond $X=1.165 $Y=1.295
+ $X2=1.165 $Y2=1.395
r51 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.065 $Y=1.735
+ $X2=1.065 $Y2=1.395
r52 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.735
+ $X2=1.065 $Y2=1.9
r53 10 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.23
+ $X2=1.065 $Y2=1.395
r54 7 12 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=1.155 $Y=2.735
+ $X2=1.155 $Y2=1.9
r55 3 10 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.155 $Y=0.445
+ $X2=1.155 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_0%B1 2 5 9 11 12 14 21
r42 21 23 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.355
+ $X2=1.62 $Y2=1.19
r43 12 14 9.37226 $w=6.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.635 $Y=1.525
+ $X2=2.16 $Y2=1.525
r44 12 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.635
+ $Y=1.355 $X2=1.635 $Y2=1.355
r45 9 23 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=1.655 $Y=0.445
+ $X2=1.655 $Y2=1.19
r46 5 11 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.515 $Y=2.735
+ $X2=1.515 $Y2=1.86
r47 2 11 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.62 $Y=1.68 $X2=1.62
+ $Y2=1.86
r48 1 21 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.62 $Y=1.37 $X2=1.62
+ $Y2=1.355
r49 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.62 $Y=1.37 $X2=1.62
+ $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_0%A1 3 7 10 15 16 17 22
c48 22 0 9.69801e-21 $X=2.52 $Y=1.37
c49 10 0 1.27929e-19 $X=2.1 $Y=2.1
c50 7 0 1.62485e-19 $X=2.085 $Y=0.445
r51 22 25 72.7041 $w=6.75e-07 $l=5.05e-07 $layer=POLY_cond $X=2.347 $Y=1.37
+ $X2=2.347 $Y2=1.875
r52 22 24 51.7148 $w=6.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.347 $Y=1.37
+ $X2=2.347 $Y2=1.205
r53 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.37 $X2=2.52 $Y2=1.37
r54 17 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.6 $Y=1.665
+ $X2=2.6 $Y2=1.37
r55 16 23 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=2.6 $Y=1.295 $X2=2.6
+ $Y2=1.37
r56 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.6 $Y=0.925 $X2=2.6
+ $Y2=1.295
r57 10 11 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.1 $Y=2.175
+ $X2=1.945 $Y2=2.175
r58 10 25 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=2.1 $Y=2.1 $X2=2.1
+ $Y2=1.875
r59 7 24 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.085 $Y=0.445
+ $X2=2.085 $Y2=1.205
r60 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.945 $Y=2.25
+ $X2=1.945 $Y2=2.175
r61 1 3 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.945 $Y=2.25
+ $X2=1.945 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_0%A2 3 7 9 10 11 12 14 17 18 19 20 21 27
r45 20 21 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=1.665
+ $X2=3.105 $Y2=2.035
r46 19 20 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=1.295
+ $X2=3.105 $Y2=1.665
r47 18 19 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=0.925
+ $X2=3.105 $Y2=1.295
r48 18 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.005 $X2=3.09 $Y2=1.005
r49 16 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.09 $Y=1.345
+ $X2=3.09 $Y2=1.005
r50 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.345
+ $X2=3.09 $Y2=1.51
r51 15 27 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.09 $Y=0.965 $X2=3.09
+ $Y2=1.005
r52 14 17 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=3 $Y=2.115 $X2=3
+ $Y2=1.51
r53 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.925 $Y=2.19
+ $X2=3 $Y2=2.115
r54 11 12 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.925 $Y=2.19
+ $X2=2.55 $Y2=2.19
r55 9 15 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.925 $Y=0.89
+ $X2=3.09 $Y2=0.965
r56 9 10 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.925 $Y=0.89
+ $X2=2.52 $Y2=0.89
r57 5 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.475 $Y=2.265
+ $X2=2.55 $Y2=2.19
r58 5 7 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.475 $Y=2.265 $X2=2.475
+ $Y2=2.735
r59 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.445 $Y=0.815
+ $X2=2.52 $Y2=0.89
r60 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.445 $Y=0.815
+ $X2=2.445 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_0%Y 1 2 3 10 12 18 20 21 22 23 30 31 36 43
c50 30 0 1.62485e-19 $X=1.735 $Y=0.9
r51 43 45 10.2682 $w=5.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2 $Y=0.445 $X2=2
+ $Y2=0.9
r52 31 41 6.14636 $w=2.38e-07 $l=1.28e-07 $layer=LI1_cond $X=1.065 $Y=0.9
+ $X2=0.937 $Y2=0.9
r53 30 45 5.39456 $w=2.4e-07 $l=2.65e-07 $layer=LI1_cond $X=1.735 $Y=0.9 $X2=2
+ $Y2=0.9
r54 30 36 2.64102 $w=2.38e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=0.9
+ $X2=1.68 $Y2=0.9
r55 23 45 0.564188 $w=5.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2 $Y=0.925 $X2=2
+ $Y2=0.9
r56 23 36 0.720277 $w=2.38e-07 $l=1.5e-08 $layer=LI1_cond $X=1.665 $Y=0.9
+ $X2=1.68 $Y2=0.9
r57 22 23 22.3286 $w=2.38e-07 $l=4.65e-07 $layer=LI1_cond $X=1.2 $Y=0.9
+ $X2=1.665 $Y2=0.9
r58 22 31 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=0.9
+ $X2=1.065 $Y2=0.9
r59 21 41 10.42 $w=2.38e-07 $l=2.17e-07 $layer=LI1_cond $X=0.72 $Y=0.9 $X2=0.937
+ $Y2=0.9
r60 21 37 4.80185 $w=2.38e-07 $l=1e-07 $layer=LI1_cond $X=0.72 $Y=0.9 $X2=0.62
+ $Y2=0.9
r61 16 41 0.368803 $w=2.55e-07 $l=1.2e-07 $layer=LI1_cond $X=0.937 $Y=0.78
+ $X2=0.937 $Y2=0.9
r62 16 18 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=0.937 $Y=0.78
+ $X2=0.937 $Y2=0.445
r63 14 37 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.62 $Y=1.02 $X2=0.62
+ $Y2=0.9
r64 14 20 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=0.62 $Y=1.02
+ $X2=0.62 $Y2=2.395
r65 10 20 8.28018 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.545 $Y=2.555
+ $X2=0.545 $Y2=2.395
r66 10 12 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=0.545 $Y=2.555
+ $X2=0.545 $Y2=2.56
r67 3 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.425
+ $Y=2.415 $X2=0.55 $Y2=2.56
r68 2 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.73
+ $Y=0.235 $X2=1.87 $Y2=0.445
r69 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.8
+ $Y=0.235 $X2=0.94 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_0%A_318_483# 1 2 9 11 12 15 17 19
c35 19 0 1.27929e-19 $X=2.697 $Y=2.395
c36 12 0 1.52116e-19 $X=1.86 $Y=2.135
r37 15 19 6.70178 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=2.697 $Y=2.552
+ $X2=2.697 $Y2=2.395
r38 15 17 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=2.697 $Y=2.552
+ $X2=2.697 $Y2=2.56
r39 13 19 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=2.652 $Y=2.225
+ $X2=2.652 $Y2=2.395
r40 11 13 6.92652 $w=1.8e-07 $l=1.50413e-07 $layer=LI1_cond $X=2.54 $Y=2.135
+ $X2=2.652 $Y2=2.225
r41 11 12 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.54 $Y=2.135
+ $X2=1.86 $Y2=2.135
r42 7 12 7.34943 $w=1.8e-07 $l=1.87681e-07 $layer=LI1_cond $X=1.712 $Y=2.225
+ $X2=1.86 $Y2=2.135
r43 7 9 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=1.712 $Y=2.225
+ $X2=1.712 $Y2=2.56
r44 2 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.55
+ $Y=2.415 $X2=2.69 $Y2=2.56
r45 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=2.415 $X2=1.73 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_0%VPWR 1 6 8 10 20 21 24
r30 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r33 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.205 $Y2=3.33
r34 18 20 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=2.205 $Y2=3.33
r38 10 16 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 8 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=3.245
+ $X2=2.205 $Y2=3.33
r43 4 6 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.205 $Y=3.245
+ $X2=2.205 $Y2=2.57
r44 1 6 300 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=2 $X=2.02
+ $Y=2.415 $X2=2.205 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_0%VGND 1 2 3 12 16 20 23 24 26 27 28 37 43
+ 44 47
c47 20 0 9.69801e-21 $X=2.66 $Y=0.445
r48 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r49 44 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r50 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r51 41 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.66
+ $Y2=0
r52 41 43 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=3.12
+ $Y2=0
r53 40 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r54 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r55 37 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.66
+ $Y2=0
r56 37 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.16
+ $Y2=0
r57 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r58 32 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r59 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r60 28 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r61 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r62 26 35 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.2
+ $Y2=0
r63 26 27 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.397
+ $Y2=0
r64 25 39 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=2.16
+ $Y2=0
r65 25 27 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.397
+ $Y2=0
r66 23 31 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.24
+ $Y2=0
r67 23 24 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.492
+ $Y2=0
r68 22 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.64 $Y=0 $X2=1.2
+ $Y2=0
r69 22 24 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.64 $Y=0 $X2=0.492
+ $Y2=0
r70 18 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0
r71 18 20 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0.445
r72 14 27 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.397 $Y=0.085
+ $X2=1.397 $Y2=0
r73 14 16 12.7655 $w=3.23e-07 $l=3.6e-07 $layer=LI1_cond $X=1.397 $Y=0.085
+ $X2=1.397 $Y2=0.445
r74 10 24 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.492 $Y=0.085
+ $X2=0.492 $Y2=0
r75 10 12 14.0637 $w=2.93e-07 $l=3.6e-07 $layer=LI1_cond $X=0.492 $Y=0.085
+ $X2=0.492 $Y2=0.445
r76 3 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.52
+ $Y=0.235 $X2=2.66 $Y2=0.445
r77 2 16 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=1.23
+ $Y=0.235 $X2=1.39 $Y2=0.445
r78 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.385
+ $Y=0.235 $X2=0.51 $Y2=0.445
.ends

