* File: sky130_fd_sc_lp__dfrbp_1.spice
* Created: Wed Sep  2 09:43:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfrbp_1.pex.spice"
.subckt sky130_fd_sc_lp__dfrbp_1  VNB VPB CLK D RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1027 N_VGND_M1027_d N_CLK_M1027_g N_A_28_108#_M1027_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1014 N_A_197_108#_M1014_d N_A_28_108#_M1014_g N_VGND_M1027_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_423_191# N_RESET_B_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.32025 PD=0.63 PS=2.69 NRD=14.28 NRS=202.14 M=1 R=2.8 SA=75000.3
+ SB=75004.7 A=0.063 P=1.14 MULT=1
MM1022 N_A_304_463#_M1022_d N_D_M1022_g A_423_191# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=17.136 NRS=14.28 M=1 R=2.8 SA=75000.7
+ SB=75004.3 A=0.063 P=1.14 MULT=1
MM1003 N_A_603_191#_M1003_d N_A_28_108#_M1003_g N_A_304_463#_M1022_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.13545 AS=0.0819 PD=1.065 PS=0.81 NRD=104.28 NRS=14.28 M=1
+ R=2.8 SA=75001.2 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1019 A_762_191# N_A_197_108#_M1019_g N_A_603_191#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.13545 PD=0.7 PS=1.065 NRD=24.276 NRS=0 M=1 R=2.8
+ SA=75002 SB=75003 A=0.063 P=1.14 MULT=1
MM1010 A_848_191# N_A_804_328#_M1010_g A_762_191# VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=24.276 M=1 R=2.8 SA=75002.5
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_RESET_B_M1026_g A_848_191# VNB NSHORT L=0.15 W=0.42
+ AD=0.23625 AS=0.0672 PD=1.56906 PS=0.74 NRD=144.996 NRS=30 M=1 R=2.8
+ SA=75002.9 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1020 N_A_804_328#_M1020_d N_A_603_191#_M1020_g N_VGND_M1026_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.36 PD=0.92 PS=2.39094 NRD=0 NRS=95.148 M=1
+ R=4.26667 SA=75002.3 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1021 N_A_1245_128#_M1021_d N_A_197_108#_M1021_g N_A_804_328#_M1020_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.26554 AS=0.0896 PD=1.6483 PS=0.92 NRD=63.744 NRS=0
+ M=1 R=4.26667 SA=75002.7 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1005 A_1420_128# N_A_28_108#_M1005_g N_A_1245_128#_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.17426 PD=0.63 PS=1.0817 NRD=14.28 NRS=30.708 M=1 R=2.8
+ SA=75002.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_A_1440_304#_M1033_g A_1420_128# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1017 A_1578_128# N_RESET_B_M1017_g N_VGND_M1033_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_A_1440_304#_M1024_d N_A_1245_128#_M1024_g A_1578_128# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75003.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_A_1245_128#_M1031_g N_A_1796_139#_M1031_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.117233 AS=0.1883 PD=0.936667 PS=1.78 NRD=64.032 NRS=34.284
+ M=1 R=2.8 SA=75000.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_Q_M1007_d N_A_1796_139#_M1007_g N_VGND_M1031_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.234467 PD=2.25 PS=1.87333 NRD=0 NRS=9.276 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_Q_N_M1008_d N_A_1245_128#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.2394 PD=2.21 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_28_108#_M1012_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1028 N_A_197_108#_M1028_d N_A_28_108#_M1028_g N_VPWR_M1012_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1025 N_VPWR_M1025_d N_RESET_B_M1025_g N_A_304_463#_M1025_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1125 AS=0.1113 PD=1.02 PS=1.37 NRD=35.1645 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1013 N_A_304_463#_M1013_d N_D_M1013_g N_VPWR_M1025_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1125 PD=1.41 PS=1.02 NRD=0 NRS=35.1645 M=1 R=2.8 SA=75000.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_603_191#_M1018_d N_A_197_108#_M1018_g N_A_304_463#_M1018_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1155 PD=0.7 PS=1.39 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1011 A_789_463# N_A_28_108#_M1011_g N_A_603_191#_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_804_328#_M1009_g A_789_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1065 AS=0.0441 PD=1 PS=0.63 NRD=30.4759 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 N_A_603_191#_M1015_d N_RESET_B_M1015_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1065 PD=1.37 PS=1 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 N_A_804_328#_M1032_d N_A_603_191#_M1032_g N_VPWR_M1032_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.234825 AS=0.2226 PD=1.515 PS=2.21 NRD=22.655 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1029 N_A_1245_128#_M1029_d N_A_28_108#_M1029_g N_A_804_328#_M1032_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1792 AS=0.234825 PD=1.62 PS=1.515 NRD=0 NRS=32.0322
+ M=1 R=5.6 SA=75000.7 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1002 A_1398_472# N_A_197_108#_M1002_g N_A_1245_128#_M1029_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0896 PD=0.63 PS=0.81 NRD=23.443 NRS=46.886 M=1 R=2.8
+ SA=75001.3 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_1440_304#_M1001_g A_1398_472# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1323 AS=0.0441 PD=1.05 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75001.7 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1016 N_A_1440_304#_M1016_d N_RESET_B_M1016_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1323 PD=0.7 PS=1.05 NRD=0 NRS=0 M=1 R=2.8 SA=75002.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_1245_128#_M1006_g N_A_1440_304#_M1016_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1030 N_VPWR_M1030_d N_A_1245_128#_M1030_g N_A_1796_139#_M1030_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1004_d N_A_1796_139#_M1004_g N_Q_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.21105 AS=0.3339 PD=1.595 PS=3.05 NRD=5.4569 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1023 N_Q_N_M1023_d N_A_1245_128#_M1023_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.21105 PD=3.09 PS=1.595 NRD=3.1126 NRS=3.1126 M=1 R=8.4
+ SA=75000.7 SB=75000.2 A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=21.9574 P=27.65
c_245 VPB 0 6.47584e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dfrbp_1.pxi.spice"
*
.ends
*
*
