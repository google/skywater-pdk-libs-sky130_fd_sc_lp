* File: sky130_fd_sc_lp__clkbuf_lp.spice
* Created: Fri Aug 28 10:15:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkbuf_lp.pex.spice"
.subckt sky130_fd_sc_lp__clkbuf_lp  VNB VPB A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1000 A_124_57# N_A_94_31#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_94_31#_M1005_g A_124_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0903 AS=0.0441 PD=0.85 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 A_312_57# N_A_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0903 PD=0.63 PS=0.85 NRD=14.28 NRS=42.852 M=1 R=2.8 SA=75001.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_94_31#_M1003_d N_A_M1003_g A_312_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_94_31#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.2625 AS=0.285 PD=1.525 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_A_94_31#_M1001_d N_A_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.2625 PD=2.57 PS=1.525 NRD=0 NRS=48.265 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__clkbuf_lp.pxi.spice"
*
.ends
*
*
