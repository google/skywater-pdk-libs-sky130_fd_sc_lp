* File: sky130_fd_sc_lp__a32o_2.pxi.spice
* Created: Wed Sep  2 09:27:41 2020
* 
x_PM_SKY130_FD_SC_LP__A32O_2%A_108_267# N_A_108_267#_M1010_d
+ N_A_108_267#_M1008_d N_A_108_267#_M1005_g N_A_108_267#_M1001_g
+ N_A_108_267#_M1006_g N_A_108_267#_M1011_g N_A_108_267#_c_74_n
+ N_A_108_267#_c_75_n N_A_108_267#_c_112_p N_A_108_267#_c_98_p
+ N_A_108_267#_c_76_n N_A_108_267#_c_77_n N_A_108_267#_c_78_n
+ PM_SKY130_FD_SC_LP__A32O_2%A_108_267#
x_PM_SKY130_FD_SC_LP__A32O_2%B2 N_B2_c_152_n N_B2_M1008_g N_B2_M1000_g B2
+ N_B2_c_150_n N_B2_c_151_n PM_SKY130_FD_SC_LP__A32O_2%B2
x_PM_SKY130_FD_SC_LP__A32O_2%B1 N_B1_c_187_n N_B1_M1010_g N_B1_M1003_g B1 B1 B1
+ B1 N_B1_c_190_n PM_SKY130_FD_SC_LP__A32O_2%B1
x_PM_SKY130_FD_SC_LP__A32O_2%A1 N_A1_M1002_g N_A1_M1007_g A1 A1 A1 N_A1_c_228_n
+ N_A1_c_229_n PM_SKY130_FD_SC_LP__A32O_2%A1
x_PM_SKY130_FD_SC_LP__A32O_2%A2 N_A2_M1009_g N_A2_M1004_g A2 A2 A2 N_A2_c_267_n
+ N_A2_c_268_n PM_SKY130_FD_SC_LP__A32O_2%A2
x_PM_SKY130_FD_SC_LP__A32O_2%A3 N_A3_M1013_g N_A3_M1012_g A3 A3 N_A3_c_302_n
+ PM_SKY130_FD_SC_LP__A32O_2%A3
x_PM_SKY130_FD_SC_LP__A32O_2%X N_X_M1001_s N_X_M1005_s N_X_M1006_s N_X_c_324_n
+ N_X_c_325_n N_X_c_361_p N_X_c_326_n N_X_c_322_n N_X_c_327_n X
+ PM_SKY130_FD_SC_LP__A32O_2%X
x_PM_SKY130_FD_SC_LP__A32O_2%VPWR N_VPWR_M1005_d N_VPWR_M1007_d N_VPWR_M1012_d
+ N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n
+ N_VPWR_c_370_n VPWR N_VPWR_c_371_n N_VPWR_c_372_n N_VPWR_c_364_n
+ PM_SKY130_FD_SC_LP__A32O_2%VPWR
x_PM_SKY130_FD_SC_LP__A32O_2%A_345_367# N_A_345_367#_M1008_s
+ N_A_345_367#_M1003_d N_A_345_367#_M1004_d N_A_345_367#_c_419_n
+ N_A_345_367#_c_420_n N_A_345_367#_c_433_n N_A_345_367#_c_421_n
+ N_A_345_367#_c_422_n N_A_345_367#_c_447_n N_A_345_367#_c_423_n
+ N_A_345_367#_c_430_n PM_SKY130_FD_SC_LP__A32O_2%A_345_367#
x_PM_SKY130_FD_SC_LP__A32O_2%VGND N_VGND_M1001_d N_VGND_M1011_d N_VGND_M1013_d
+ N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n
+ VGND N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n
+ PM_SKY130_FD_SC_LP__A32O_2%VGND
cc_1 VNB N_A_108_267#_M1005_g 0.009776f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_2 VNB N_A_108_267#_M1001_g 0.0273258f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.655
cc_3 VNB N_A_108_267#_M1011_g 0.0283796f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=0.655
cc_4 VNB N_A_108_267#_c_74_n 0.00221617f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.405
cc_5 VNB N_A_108_267#_c_75_n 0.010638f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.09
cc_6 VNB N_A_108_267#_c_76_n 0.00608371f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.98
cc_7 VNB N_A_108_267#_c_77_n 0.00124312f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.505
cc_8 VNB N_A_108_267#_c_78_n 0.047534f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.5
cc_9 VNB N_B2_M1000_g 0.0280013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B2_c_150_n 0.0060695f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.655
cc_11 VNB N_B2_c_151_n 0.0370275f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.655
cc_12 VNB N_B1_c_187_n 0.0169015f $X=-0.19 $Y=-0.245 $X2=2.52 $Y2=0.235
cc_13 VNB N_B1_M1003_g 0.00781712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB B1 0.00344939f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_15 VNB N_B1_c_190_n 0.0422081f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=2.465
cc_16 VNB N_A1_M1007_g 0.00919584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A1 0.00170702f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_18 VNB N_A1_c_228_n 0.0344932f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=1.665
cc_19 VNB N_A1_c_229_n 0.0185773f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=2.465
cc_20 VNB N_A2_M1004_g 0.00801241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A2 0.00945979f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_22 VNB N_A2_c_267_n 0.0285538f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=0.655
cc_23 VNB N_A2_c_268_n 0.0172487f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.175
cc_24 VNB N_A3_M1013_g 0.0244396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A3_M1012_g 0.00646773f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.485
cc_26 VNB A3 0.0252096f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_27 VNB N_A3_c_302_n 0.0536241f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=2.465
cc_28 VNB N_X_c_322_n 0.021596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB X 0.0224932f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.5
cc_30 VNB N_VPWR_c_364_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_468_n 0.0284267f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.655
cc_32 VNB N_VGND_c_469_n 0.0138045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_470_n 0.0354271f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=2.465
cc_34 VNB N_VGND_c_471_n 0.0143948f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.335
cc_35 VNB N_VGND_c_472_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=0.655
cc_36 VNB N_VGND_c_473_n 0.0129657f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.175
cc_37 VNB N_VGND_c_474_n 0.0584121f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.505
cc_38 VNB N_VGND_c_475_n 0.0152853f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.335
cc_39 VNB N_VGND_c_476_n 0.26424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_A_108_267#_M1005_g 0.0234232f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.465
cc_41 VPB N_A_108_267#_M1006_g 0.0234083f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=2.465
cc_42 VPB N_A_108_267#_c_76_n 0.00346902f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=1.98
cc_43 VPB N_A_108_267#_c_78_n 0.00803445f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=1.5
cc_44 VPB N_B2_c_152_n 0.0206104f $X=-0.19 $Y=1.655 $X2=2.52 $Y2=0.235
cc_45 VPB N_B2_c_150_n 0.00809068f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=0.655
cc_46 VPB N_B2_c_151_n 0.015912f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=0.655
cc_47 VPB N_B1_M1003_g 0.0219858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB B1 0.00171639f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.465
cc_49 VPB N_A1_M1007_g 0.0232217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A2_M1004_g 0.0206299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A3_M1012_g 0.024843f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.485
cc_52 VPB A3 0.0136741f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.465
cc_53 VPB N_X_c_324_n 0.0480658f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=0.655
cc_54 VPB N_X_c_325_n 0.00593056f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=2.465
cc_55 VPB N_X_c_326_n 0.0113011f $X=-0.19 $Y=1.655 $X2=1.33 $Y2=1.405
cc_56 VPB N_X_c_327_n 0.00786683f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=1.5
cc_57 VPB X 0.00708404f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=1.5
cc_58 VPB N_VPWR_c_365_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_366_n 0.00493725f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=0.655
cc_60 VPB N_VPWR_c_367_n 0.015603f $X=-0.19 $Y=1.655 $X2=1.33 $Y2=1.405
cc_61 VPB N_VPWR_c_368_n 0.0482736f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.09
cc_62 VPB N_VPWR_c_369_n 0.0560374f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=1.505
cc_63 VPB N_VPWR_c_370_n 0.00631825f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=1.5
cc_64 VPB N_VPWR_c_371_n 0.0149762f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=1.5
cc_65 VPB N_VPWR_c_372_n 0.023447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_364_n 0.0666718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_345_367#_c_419_n 0.00204872f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_345_367#_c_420_n 0.0101684f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=0.655
cc_69 VPB N_A_345_367#_c_421_n 0.00896518f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=0.655
cc_70 VPB N_A_345_367#_c_422_n 0.00578436f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=0.655
cc_71 N_A_108_267#_c_74_n N_B2_M1000_g 0.00355919f $X=1.33 $Y=1.405 $X2=0 $Y2=0
cc_72 N_A_108_267#_c_75_n N_B2_M1000_g 0.0202031f $X=2.185 $Y=1.09 $X2=0 $Y2=0
cc_73 N_A_108_267#_c_76_n N_B2_M1000_g 0.00540172f $X=2.28 $Y=1.98 $X2=0 $Y2=0
cc_74 N_A_108_267#_c_78_n N_B2_M1000_g 2.30293e-19 $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_75 N_A_108_267#_M1006_g N_B2_c_150_n 0.00213216f $X=1.045 $Y=2.465 $X2=0
+ $Y2=0
cc_76 N_A_108_267#_c_74_n N_B2_c_150_n 0.00463237f $X=1.33 $Y=1.405 $X2=0 $Y2=0
cc_77 N_A_108_267#_c_75_n N_B2_c_150_n 0.0331775f $X=2.185 $Y=1.09 $X2=0 $Y2=0
cc_78 N_A_108_267#_c_76_n N_B2_c_150_n 0.0320562f $X=2.28 $Y=1.98 $X2=0 $Y2=0
cc_79 N_A_108_267#_c_77_n N_B2_c_150_n 0.016084f $X=1.33 $Y=1.505 $X2=0 $Y2=0
cc_80 N_A_108_267#_c_78_n N_B2_c_150_n 0.00267292f $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_81 N_A_108_267#_M1006_g N_B2_c_151_n 0.00100504f $X=1.045 $Y=2.465 $X2=0
+ $Y2=0
cc_82 N_A_108_267#_c_75_n N_B2_c_151_n 0.00249493f $X=2.185 $Y=1.09 $X2=0 $Y2=0
cc_83 N_A_108_267#_c_76_n N_B2_c_151_n 0.00490003f $X=2.28 $Y=1.98 $X2=0 $Y2=0
cc_84 N_A_108_267#_c_77_n N_B2_c_151_n 2.18154e-19 $X=1.33 $Y=1.505 $X2=0 $Y2=0
cc_85 N_A_108_267#_c_78_n N_B2_c_151_n 0.0176464f $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_86 N_A_108_267#_c_98_p N_B1_c_187_n 0.039748f $X=2.28 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A_108_267#_c_76_n N_B1_c_187_n 2.025e-19 $X=2.28 $Y=1.98 $X2=-0.19
+ $Y2=-0.245
cc_88 N_A_108_267#_c_98_p B1 0.0143759f $X=2.28 $Y=1.175 $X2=0 $Y2=0
cc_89 N_A_108_267#_c_76_n B1 0.0721518f $X=2.28 $Y=1.98 $X2=0 $Y2=0
cc_90 N_A_108_267#_c_98_p N_B1_c_190_n 0.00405937f $X=2.28 $Y=1.175 $X2=0 $Y2=0
cc_91 N_A_108_267#_c_76_n N_B1_c_190_n 0.0076089f $X=2.28 $Y=1.98 $X2=0 $Y2=0
cc_92 N_A_108_267#_c_98_p A1 0.0559049f $X=2.28 $Y=1.175 $X2=0 $Y2=0
cc_93 N_A_108_267#_c_98_p N_A1_c_229_n 0.00938731f $X=2.28 $Y=1.175 $X2=0 $Y2=0
cc_94 N_A_108_267#_M1006_g N_X_c_325_n 0.0148266f $X=1.045 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A_108_267#_c_77_n N_X_c_325_n 0.0259714f $X=1.33 $Y=1.505 $X2=0 $Y2=0
cc_96 N_A_108_267#_c_78_n N_X_c_325_n 0.00810055f $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_97 N_A_108_267#_M1001_g N_X_c_322_n 0.0145838f $X=0.765 $Y=0.655 $X2=0 $Y2=0
cc_98 N_A_108_267#_M1011_g N_X_c_322_n 0.00183f $X=1.195 $Y=0.655 $X2=0 $Y2=0
cc_99 N_A_108_267#_c_74_n N_X_c_322_n 0.00478504f $X=1.33 $Y=1.405 $X2=0 $Y2=0
cc_100 N_A_108_267#_c_112_p N_X_c_322_n 0.0117765f $X=1.415 $Y=1.09 $X2=0 $Y2=0
cc_101 N_A_108_267#_c_78_n N_X_c_322_n 0.00356846f $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_102 N_A_108_267#_M1005_g N_X_c_327_n 0.0125148f $X=0.615 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_108_267#_M1005_g X 0.0125676f $X=0.615 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A_108_267#_M1001_g X 0.00401439f $X=0.765 $Y=0.655 $X2=0 $Y2=0
cc_105 N_A_108_267#_M1011_g X 8.12635e-19 $X=1.195 $Y=0.655 $X2=0 $Y2=0
cc_106 N_A_108_267#_c_74_n X 0.00735357f $X=1.33 $Y=1.405 $X2=0 $Y2=0
cc_107 N_A_108_267#_c_77_n X 0.0139528f $X=1.33 $Y=1.505 $X2=0 $Y2=0
cc_108 N_A_108_267#_c_78_n X 0.0220714f $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_109 N_A_108_267#_M1005_g N_VPWR_c_365_n 0.0159851f $X=0.615 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_108_267#_M1006_g N_VPWR_c_365_n 0.0159861f $X=1.045 $Y=2.465 $X2=0
+ $Y2=0
cc_111 N_A_108_267#_c_78_n N_VPWR_c_365_n 3.17289e-19 $X=1.195 $Y=1.5 $X2=0
+ $Y2=0
cc_112 N_A_108_267#_M1006_g N_VPWR_c_369_n 0.00486043f $X=1.045 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_108_267#_M1005_g N_VPWR_c_372_n 0.00486043f $X=0.615 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_108_267#_M1008_d N_VPWR_c_364_n 0.00225186f $X=2.14 $Y=1.835 $X2=0
+ $Y2=0
cc_115 N_A_108_267#_M1005_g N_VPWR_c_364_n 0.00928803f $X=0.615 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_108_267#_M1006_g N_VPWR_c_364_n 0.00954696f $X=1.045 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_108_267#_M1008_d N_A_345_367#_c_423_n 0.00332344f $X=2.14 $Y=1.835
+ $X2=0 $Y2=0
cc_118 N_A_108_267#_c_76_n N_A_345_367#_c_423_n 0.0126348f $X=2.28 $Y=1.98 $X2=0
+ $Y2=0
cc_119 N_A_108_267#_c_75_n N_VGND_M1011_d 0.0071597f $X=2.185 $Y=1.09 $X2=0
+ $Y2=0
cc_120 N_A_108_267#_c_112_p N_VGND_M1011_d 9.47307e-19 $X=1.415 $Y=1.09 $X2=0
+ $Y2=0
cc_121 N_A_108_267#_M1001_g N_VGND_c_468_n 0.0126571f $X=0.765 $Y=0.655 $X2=0
+ $Y2=0
cc_122 N_A_108_267#_M1011_g N_VGND_c_468_n 6.30983e-19 $X=1.195 $Y=0.655 $X2=0
+ $Y2=0
cc_123 N_A_108_267#_c_78_n N_VGND_c_468_n 5.44298e-19 $X=1.195 $Y=1.5 $X2=0
+ $Y2=0
cc_124 N_A_108_267#_M1001_g N_VGND_c_473_n 0.00486043f $X=0.765 $Y=0.655 $X2=0
+ $Y2=0
cc_125 N_A_108_267#_M1011_g N_VGND_c_473_n 0.00487821f $X=1.195 $Y=0.655 $X2=0
+ $Y2=0
cc_126 N_A_108_267#_c_98_p N_VGND_c_474_n 0.0416965f $X=2.28 $Y=1.175 $X2=0
+ $Y2=0
cc_127 N_A_108_267#_M1001_g N_VGND_c_475_n 6.29646e-19 $X=0.765 $Y=0.655 $X2=0
+ $Y2=0
cc_128 N_A_108_267#_M1011_g N_VGND_c_475_n 0.0117428f $X=1.195 $Y=0.655 $X2=0
+ $Y2=0
cc_129 N_A_108_267#_c_75_n N_VGND_c_475_n 0.0455205f $X=2.185 $Y=1.09 $X2=0
+ $Y2=0
cc_130 N_A_108_267#_c_112_p N_VGND_c_475_n 0.0095479f $X=1.415 $Y=1.09 $X2=0
+ $Y2=0
cc_131 N_A_108_267#_c_78_n N_VGND_c_475_n 4.72016e-19 $X=1.195 $Y=1.5 $X2=0
+ $Y2=0
cc_132 N_A_108_267#_M1010_d N_VGND_c_476_n 0.00881249f $X=2.52 $Y=0.235 $X2=0
+ $Y2=0
cc_133 N_A_108_267#_M1001_g N_VGND_c_476_n 0.00824727f $X=0.765 $Y=0.655 $X2=0
+ $Y2=0
cc_134 N_A_108_267#_M1011_g N_VGND_c_476_n 0.00824731f $X=1.195 $Y=0.655 $X2=0
+ $Y2=0
cc_135 N_A_108_267#_c_98_p N_VGND_c_476_n 0.0249729f $X=2.28 $Y=1.175 $X2=0
+ $Y2=0
cc_136 N_A_108_267#_c_98_p A_432_47# 9.38685e-19 $X=2.28 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_137 N_B2_M1000_g N_B1_c_187_n 0.0741757f $X=2.085 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_138 N_B2_c_152_n N_B1_M1003_g 0.0202732f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_139 N_B2_M1000_g N_B1_c_190_n 0.00722442f $X=2.085 $Y=0.655 $X2=0 $Y2=0
cc_140 N_B2_c_151_n N_B1_c_190_n 0.0202732f $X=2.065 $Y=1.535 $X2=0 $Y2=0
cc_141 N_B2_c_152_n N_X_c_325_n 0.0031258f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_142 N_B2_c_152_n N_X_c_326_n 0.00230071f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_143 N_B2_c_152_n N_VPWR_c_369_n 0.00357842f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_144 N_B2_c_152_n N_VPWR_c_364_n 0.00667816f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_145 N_B2_c_152_n N_A_345_367#_c_419_n 5.81207e-19 $X=2.065 $Y=1.725 $X2=0
+ $Y2=0
cc_146 N_B2_c_152_n N_A_345_367#_c_420_n 0.0145157f $X=2.065 $Y=1.725 $X2=0
+ $Y2=0
cc_147 N_B2_c_150_n N_A_345_367#_c_420_n 0.0263417f $X=1.82 $Y=1.51 $X2=0 $Y2=0
cc_148 N_B2_c_151_n N_A_345_367#_c_420_n 0.00202073f $X=2.065 $Y=1.535 $X2=0
+ $Y2=0
cc_149 N_B2_c_152_n N_A_345_367#_c_423_n 0.010474f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_150 N_B2_c_152_n N_A_345_367#_c_430_n 4.13013e-19 $X=2.065 $Y=1.725 $X2=0
+ $Y2=0
cc_151 N_B2_M1000_g N_VGND_c_474_n 0.00487821f $X=2.085 $Y=0.655 $X2=0 $Y2=0
cc_152 N_B2_M1000_g N_VGND_c_475_n 0.0128112f $X=2.085 $Y=0.655 $X2=0 $Y2=0
cc_153 N_B2_M1000_g N_VGND_c_476_n 0.00818716f $X=2.085 $Y=0.655 $X2=0 $Y2=0
cc_154 N_B1_M1003_g N_A1_M1007_g 0.0182584f $X=2.495 $Y=2.465 $X2=0 $Y2=0
cc_155 B1 N_A1_M1007_g 0.00464209f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B1_c_187_n A1 0.00115342f $X=2.445 $Y=1.185 $X2=0 $Y2=0
cc_157 B1 A1 0.0146112f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_158 N_B1_c_190_n A1 0.00118698f $X=2.495 $Y=1.35 $X2=0 $Y2=0
cc_159 B1 N_A1_c_228_n 0.00107513f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_160 N_B1_c_190_n N_A1_c_228_n 0.020726f $X=2.495 $Y=1.35 $X2=0 $Y2=0
cc_161 N_B1_c_187_n N_A1_c_229_n 0.0210987f $X=2.445 $Y=1.185 $X2=0 $Y2=0
cc_162 N_B1_M1003_g N_VPWR_c_369_n 0.00357877f $X=2.495 $Y=2.465 $X2=0 $Y2=0
cc_163 N_B1_M1003_g N_VPWR_c_364_n 0.00593675f $X=2.495 $Y=2.465 $X2=0 $Y2=0
cc_164 B1 N_A_345_367#_M1003_d 0.00793079f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_165 N_B1_M1003_g N_A_345_367#_c_420_n 6.87535e-19 $X=2.495 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_B1_M1003_g N_A_345_367#_c_433_n 0.00329609f $X=2.495 $Y=2.465 $X2=0
+ $Y2=0
cc_167 B1 N_A_345_367#_c_433_n 0.0485833f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_168 N_B1_M1003_g N_A_345_367#_c_422_n 5.49694e-19 $X=2.495 $Y=2.465 $X2=0
+ $Y2=0
cc_169 B1 N_A_345_367#_c_422_n 0.0141853f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_170 N_B1_M1003_g N_A_345_367#_c_423_n 0.011404f $X=2.495 $Y=2.465 $X2=0 $Y2=0
cc_171 B1 N_A_345_367#_c_423_n 7.12352e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_172 N_B1_M1003_g N_A_345_367#_c_430_n 0.00268135f $X=2.495 $Y=2.465 $X2=0
+ $Y2=0
cc_173 B1 N_A_345_367#_c_430_n 0.00913587f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_174 N_B1_c_187_n N_VGND_c_474_n 0.00357668f $X=2.445 $Y=1.185 $X2=0 $Y2=0
cc_175 N_B1_c_187_n N_VGND_c_475_n 0.00174663f $X=2.445 $Y=1.185 $X2=0 $Y2=0
cc_176 N_B1_c_187_n N_VGND_c_476_n 0.0057288f $X=2.445 $Y=1.185 $X2=0 $Y2=0
cc_177 N_A1_M1007_g N_A2_M1004_g 0.0212413f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_178 A1 A2 0.0953118f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_179 N_A1_c_228_n A2 0.00238186f $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_180 N_A1_c_229_n A2 0.00282389f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_181 A1 N_A2_c_267_n 2.89609e-19 $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_182 N_A1_c_228_n N_A2_c_267_n 0.0204266f $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_183 A1 N_A2_c_268_n 0.00222353f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_184 N_A1_c_229_n N_A2_c_268_n 0.0324108f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_185 N_A1_M1007_g N_VPWR_c_366_n 0.003261f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A1_M1007_g N_VPWR_c_369_n 0.00585385f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A1_M1007_g N_VPWR_c_364_n 0.011496f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A1_M1007_g N_A_345_367#_c_421_n 0.0145228f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_189 A1 N_A_345_367#_c_421_n 0.00713501f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_190 N_A1_c_228_n N_A_345_367#_c_421_n 0.0019165f $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_191 N_A1_M1007_g N_A_345_367#_c_422_n 0.00109436f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_192 A1 N_A_345_367#_c_422_n 0.00646303f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_193 N_A1_c_228_n N_A_345_367#_c_422_n 0.00209743f $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_194 N_A1_M1007_g N_A_345_367#_c_447_n 4.97528e-19 $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A1_M1007_g N_A_345_367#_c_430_n 0.00413324f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_196 A1 N_VGND_c_474_n 0.007766f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_197 N_A1_c_229_n N_VGND_c_474_n 0.00421391f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_198 A1 N_VGND_c_476_n 0.00742637f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_199 N_A1_c_229_n N_VGND_c_476_n 0.00738676f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_200 A1 A_631_47# 0.00682159f $X=3.035 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_201 A2 N_A3_M1013_g 0.0321678f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_202 N_A2_c_267_n N_A3_M1013_g 0.0214182f $X=3.71 $Y=1.35 $X2=0 $Y2=0
cc_203 N_A2_c_268_n N_A3_M1013_g 0.0323555f $X=3.71 $Y=1.185 $X2=0 $Y2=0
cc_204 A2 A3 0.023339f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_205 N_A2_M1004_g N_A3_c_302_n 0.0270747f $X=3.73 $Y=2.465 $X2=0 $Y2=0
cc_206 A2 N_A3_c_302_n 0.0137223f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_207 N_A2_M1004_g N_VPWR_c_366_n 0.00172006f $X=3.73 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A2_M1004_g N_VPWR_c_368_n 8.65002e-19 $X=3.73 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A2_M1004_g N_VPWR_c_371_n 0.00579312f $X=3.73 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A2_M1004_g N_VPWR_c_364_n 0.0106875f $X=3.73 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A2_M1004_g N_A_345_367#_c_421_n 0.0143589f $X=3.73 $Y=2.465 $X2=0 $Y2=0
cc_212 A2 N_A_345_367#_c_421_n 0.0402725f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_213 N_A2_c_267_n N_A_345_367#_c_421_n 0.00124391f $X=3.71 $Y=1.35 $X2=0 $Y2=0
cc_214 N_A2_M1004_g N_A_345_367#_c_447_n 0.0133505f $X=3.73 $Y=2.465 $X2=0 $Y2=0
cc_215 A2 N_VGND_c_470_n 0.0547487f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_216 A2 N_VGND_c_474_n 0.0270272f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_217 N_A2_c_268_n N_VGND_c_474_n 0.0037867f $X=3.71 $Y=1.185 $X2=0 $Y2=0
cc_218 A2 N_VGND_c_476_n 0.0259829f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_219 N_A2_c_268_n N_VGND_c_476_n 0.00606487f $X=3.71 $Y=1.185 $X2=0 $Y2=0
cc_220 A2 A_631_47# 0.00723399f $X=3.515 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_221 A2 A_739_47# 0.00440697f $X=3.515 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_222 N_A3_M1012_g N_VPWR_c_368_n 0.0213721f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_223 A3 N_VPWR_c_368_n 0.0175032f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_224 N_A3_c_302_n N_VPWR_c_368_n 0.00378877f $X=4.43 $Y=1.375 $X2=0 $Y2=0
cc_225 N_A3_M1012_g N_VPWR_c_371_n 0.00486043f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A3_M1012_g N_VPWR_c_364_n 0.0082726f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_227 N_A3_M1012_g N_A_345_367#_c_421_n 0.00253514f $X=4.16 $Y=2.465 $X2=0
+ $Y2=0
cc_228 N_A3_M1013_g N_VGND_c_470_n 0.0104161f $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_229 A3 N_VGND_c_470_n 0.020953f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_230 N_A3_c_302_n N_VGND_c_470_n 0.00236769f $X=4.43 $Y=1.375 $X2=0 $Y2=0
cc_231 N_A3_M1013_g N_VGND_c_474_n 0.00476515f $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_232 N_A3_M1013_g N_VGND_c_476_n 0.00932429f $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_233 N_X_c_325_n N_VPWR_M1005_d 3.93317e-19 $X=1.165 $Y=1.86 $X2=-0.19
+ $Y2=-0.245
cc_234 N_X_c_327_n N_VPWR_M1005_d 0.00141648f $X=0.515 $Y=1.86 $X2=-0.19
+ $Y2=-0.245
cc_235 N_X_c_325_n N_VPWR_c_365_n 0.00484123f $X=1.165 $Y=1.86 $X2=0 $Y2=0
cc_236 N_X_c_327_n N_VPWR_c_365_n 0.01353f $X=0.515 $Y=1.86 $X2=0 $Y2=0
cc_237 N_X_c_326_n N_VPWR_c_369_n 0.0170942f $X=1.26 $Y=1.98 $X2=0 $Y2=0
cc_238 N_X_c_324_n N_VPWR_c_372_n 0.023546f $X=0.4 $Y=1.98 $X2=0 $Y2=0
cc_239 N_X_M1005_s N_VPWR_c_364_n 0.00371702f $X=0.275 $Y=1.835 $X2=0 $Y2=0
cc_240 N_X_M1006_s N_VPWR_c_364_n 0.00371702f $X=1.12 $Y=1.835 $X2=0 $Y2=0
cc_241 N_X_c_324_n N_VPWR_c_364_n 0.0131407f $X=0.4 $Y=1.98 $X2=0 $Y2=0
cc_242 N_X_c_326_n N_VPWR_c_364_n 0.00964167f $X=1.26 $Y=1.98 $X2=0 $Y2=0
cc_243 N_X_c_326_n N_A_345_367#_c_419_n 0.0106732f $X=1.26 $Y=1.98 $X2=0 $Y2=0
cc_244 N_X_c_325_n N_A_345_367#_c_420_n 9.60437e-19 $X=1.165 $Y=1.86 $X2=0 $Y2=0
cc_245 N_X_c_326_n N_A_345_367#_c_420_n 0.0567024f $X=1.26 $Y=1.98 $X2=0 $Y2=0
cc_246 N_X_c_322_n N_VGND_M1001_d 0.00234883f $X=0.615 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_247 N_X_c_322_n N_VGND_c_468_n 0.0243971f $X=0.615 $Y=1.235 $X2=0 $Y2=0
cc_248 N_X_c_361_p N_VGND_c_473_n 0.0124525f $X=0.98 $Y=0.42 $X2=0 $Y2=0
cc_249 N_X_M1001_s N_VGND_c_476_n 0.00536646f $X=0.84 $Y=0.235 $X2=0 $Y2=0
cc_250 N_X_c_361_p N_VGND_c_476_n 0.00730901f $X=0.98 $Y=0.42 $X2=0 $Y2=0
cc_251 N_VPWR_c_364_n N_A_345_367#_M1008_s 0.00215158f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_252 N_VPWR_c_364_n N_A_345_367#_M1003_d 0.00455487f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_364_n N_A_345_367#_M1004_d 0.00380103f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_369_n N_A_345_367#_c_419_n 0.0211538f $X=3.3 $Y=3.33 $X2=0 $Y2=0
cc_255 N_VPWR_c_364_n N_A_345_367#_c_419_n 0.0126374f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_256 N_VPWR_M1007_d N_A_345_367#_c_421_n 0.00291574f $X=3.28 $Y=1.835 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_366_n N_A_345_367#_c_421_n 0.0203459f $X=3.465 $Y=2.19 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_371_n N_A_345_367#_c_447_n 0.0143246f $X=4.21 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_364_n N_A_345_367#_c_447_n 0.00916141f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_369_n N_A_345_367#_c_423_n 0.0649891f $X=3.3 $Y=3.33 $X2=0 $Y2=0
cc_261 N_VPWR_c_364_n N_A_345_367#_c_423_n 0.0409084f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_VGND_c_476_n A_432_47# 0.00325419f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
cc_263 N_VGND_c_476_n A_631_47# 0.00921635f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
cc_264 N_VGND_c_476_n A_739_47# 0.00330119f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
