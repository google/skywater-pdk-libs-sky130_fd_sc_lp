* NGSPICE file created from sky130_fd_sc_lp__a32o_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 VPWR A2 a_249_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3041e+12p pd=7.11e+06u as=1.0395e+12p ps=9.21e+06u
M1001 a_609_47# B1 a_80_21# VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=5.292e+11p ps=2.94e+06u
M1002 a_263_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=2.646e+11p pd=2.31e+06u as=7.392e+11p ps=5.12e+06u
M1003 a_80_21# B1 a_249_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.032e+11p pd=3.16e+06u as=0p ps=0u
M1004 a_80_21# A1 a_356_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.814e+11p ps=2.35e+06u
M1005 VPWR a_80_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1006 VGND a_80_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1007 a_356_47# A2 a_263_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_249_367# A3 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_249_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B2 a_609_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_249_367# B2 a_80_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

