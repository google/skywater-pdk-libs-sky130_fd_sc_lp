* File: sky130_fd_sc_lp__decap_8.pxi.spice
* Created: Fri Aug 28 10:20:12 2020
* 
x_PM_SKY130_FD_SC_LP__DECAP_8%VGND N_VGND_M1000_s N_VGND_c_27_n N_VGND_c_28_n
+ N_VGND_c_29_n N_VGND_c_30_n N_VGND_c_31_n VGND N_VGND_M1001_g N_VGND_c_32_n
+ N_VGND_c_33_n N_VGND_c_34_n N_VGND_c_35_n N_VGND_c_36_n
+ PM_SKY130_FD_SC_LP__DECAP_8%VGND
x_PM_SKY130_FD_SC_LP__DECAP_8%VPWR N_VPWR_M1001_s N_VPWR_c_57_n N_VPWR_c_54_n
+ N_VPWR_c_55_n N_VPWR_c_60_n N_VPWR_c_61_n N_VPWR_c_62_n VPWR N_VPWR_M1000_g
+ N_VPWR_c_63_n N_VPWR_c_64_n N_VPWR_c_56_n N_VPWR_c_66_n
+ PM_SKY130_FD_SC_LP__DECAP_8%VPWR
cc_1 VNB N_VGND_c_27_n 0.0651019f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=0.38
cc_2 VNB N_VGND_c_28_n 0.00211035f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.77
cc_3 VNB N_VGND_c_29_n 4.60769e-19 $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.77
cc_4 VNB N_VGND_c_30_n 0.0193278f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.77
cc_5 VNB N_VGND_c_31_n 0.0371702f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=0.36
cc_6 VNB N_VGND_c_32_n 0.0598957f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=0
cc_7 VNB N_VGND_c_33_n 0.0206f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=0
cc_8 VNB N_VGND_c_34_n 0.2505f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=0
cc_9 VNB N_VGND_c_35_n 0.0279619f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_10 VNB N_VGND_c_36_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=0
cc_11 VNB N_VPWR_c_54_n 0.0260329f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.06
cc_12 VNB N_VPWR_c_55_n 0.209886f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.77
cc_13 VNB N_VPWR_c_56_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=0
cc_14 VPB N_VGND_c_28_n 0.0140672f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.77
cc_15 VPB N_VGND_c_29_n 0.00877216f $X=-0.19 $Y=1.655 $X2=1.395 $Y2=1.77
cc_16 VPB N_VGND_c_30_n 0.220826f $X=-0.19 $Y=1.655 $X2=1.395 $Y2=1.77
cc_17 VPB N_VPWR_c_57_n 0.0425694f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=0.085
cc_18 VPB N_VPWR_c_54_n 0.0010302f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=1.06
cc_19 VPB N_VPWR_c_55_n 0.0210044f $X=-0.19 $Y=1.655 $X2=1.395 $Y2=1.77
cc_20 VPB N_VPWR_c_60_n 0.0654031f $X=-0.19 $Y=1.655 $X2=3.095 $Y2=1.04
cc_21 VPB N_VPWR_c_61_n 0.0602139f $X=-0.19 $Y=1.655 $X2=1.395 $Y2=1.77
cc_22 VPB N_VPWR_c_62_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=2.595
cc_23 VPB N_VPWR_c_63_n 0.0204409f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=0
cc_24 VPB N_VPWR_c_64_n 0.0226685f $X=-0.19 $Y=1.655 $X2=3.12 $Y2=0
cc_25 VPB N_VPWR_c_56_n 0.0864025f $X=-0.19 $Y=1.655 $X2=3.12 $Y2=0
cc_26 VPB N_VPWR_c_66_n 0.00516759f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=0
cc_27 N_VGND_c_28_n N_VPWR_c_57_n 0.0205458f $X=0.98 $Y=1.77 $X2=0 $Y2=0
cc_28 N_VGND_c_30_n N_VPWR_c_57_n 0.0546006f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_29 N_VGND_c_29_n N_VPWR_c_54_n 0.00290374f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_30 N_VGND_c_30_n N_VPWR_c_54_n 0.00707553f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_31 N_VGND_c_31_n N_VPWR_c_54_n 0.0180409f $X=3.095 $Y=0.36 $X2=0 $Y2=0
cc_32 N_VGND_c_27_n N_VPWR_c_55_n 0.0654854f $X=0.815 $Y=0.38 $X2=0 $Y2=0
cc_33 N_VGND_c_29_n N_VPWR_c_55_n 0.00447085f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_34 N_VGND_c_30_n N_VPWR_c_55_n 0.127128f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_35 N_VGND_c_31_n N_VPWR_c_55_n 0.0510144f $X=3.095 $Y=0.36 $X2=0 $Y2=0
cc_36 N_VGND_c_32_n N_VPWR_c_55_n 0.0760645f $X=2.93 $Y=0 $X2=0 $Y2=0
cc_37 N_VGND_c_34_n N_VPWR_c_55_n 0.120027f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_38 N_VGND_c_30_n N_VPWR_c_60_n 0.0710714f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_39 N_VGND_c_30_n N_VPWR_c_61_n 0.0764547f $X=1.395 $Y=1.77 $X2=0 $Y2=0
cc_40 N_VGND_c_30_n N_VPWR_c_56_n 0.120644f $X=1.395 $Y=1.77 $X2=0 $Y2=0
