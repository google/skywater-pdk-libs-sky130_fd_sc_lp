* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__clkbuf_lp A VGND VNB VPB VPWR X
X0 VGND A a_312_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR A a_94_31# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_124_57# a_94_31# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 X a_94_31# a_124_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_312_57# A a_94_31# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_94_31# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
