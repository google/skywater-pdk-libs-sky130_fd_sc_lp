* File: sky130_fd_sc_lp__a211o_0.spice
* Created: Fri Aug 28 09:47:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a211o_0.pex.spice"
.subckt sky130_fd_sc_lp__a211o_0  VNB VPB A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_80_172#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.1113 PD=1.04 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1001 A_265_60# N_A2_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1302 PD=0.63 PS=1.04 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_80_172#_M1002_d N_A1_M1002_g A_265_60# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_A_80_172#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0588 PD=1.04 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_80_172#_M1000_d N_C1_M1000_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1302 PD=1.37 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_80_172#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_224_482#_M1008_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.1696 PD=0.96 PS=1.81 NRD=3.0732 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1006 N_A_224_482#_M1006_d N_A1_M1006_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=9.2196 M=1 R=4.26667
+ SA=75000.7 SB=75001 A=0.096 P=1.58 MULT=1
MM1004 A_487_482# N_B1_M1004_g N_A_224_482#_M1006_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1005 N_A_80_172#_M1005_d N_C1_M1005_g A_487_482# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a211o_0.pxi.spice"
*
.ends
*
*
