* NGSPICE file created from sky130_fd_sc_lp__o21bai_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o21bai_m A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 a_320_78# A1 VGND VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.289e+11p ps=2.77e+06u
M1001 a_320_78# a_32_62# Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1002 VGND B1_N a_32_62# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 a_315_535# A2 Y VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1004 VPWR A1 a_315_535# VPB phighvt w=420000u l=150000u
+  ad=2.835e+11p pd=3.03e+06u as=0p ps=0u
M1005 VPWR B1_N a_32_62# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 VGND A2 a_320_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_32_62# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

