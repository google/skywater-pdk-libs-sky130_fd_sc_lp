* NGSPICE file created from sky130_fd_sc_lp__a2111oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_684_47# A1 Y VNB nshort w=840000u l=150000u
+  ad=6.972e+11p pd=5.02e+06u as=1.1886e+12p ps=1.123e+07u
M1001 a_467_367# B1 a_32_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3734e+12p pd=1.226e+07u as=1.071e+12p ps=9.26e+06u
M1002 VPWR A1 a_467_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.56e+11p pd=6.24e+06u as=0p ps=0u
M1003 VGND B1 Y VNB nshort w=840000u l=150000u
+  ad=1.1802e+12p pd=9.53e+06u as=0p ps=0u
M1004 a_684_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_32_367# C1 a_115_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.16e+06u
M1006 a_467_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND D1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_115_367# C1 a_32_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_115_367# D1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1010 a_32_367# B1 a_467_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A1 a_684_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_467_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y D1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y D1 a_115_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A2 a_467_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A2 a_684_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

