* File: sky130_fd_sc_lp__mux2_8.spice
* Created: Wed Sep  2 10:00:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2_8.pex.spice"
.subckt sky130_fd_sc_lp__mux2_8  VNB VPB S A1 A0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_84_21#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75006.7 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A_84_21#_M1005_g N_X_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75006.3 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1005_d N_A_84_21#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75005.9 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A_84_21#_M1011_g N_X_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75005.5 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1011_d N_A_84_21#_M1014_g N_X_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9 SB=75005
+ A=0.126 P=1.98 MULT=1
MM1025 N_VGND_M1025_d N_A_84_21#_M1025_g N_X_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4 SB=75004.6
+ A=0.126 P=1.98 MULT=1
MM1027 N_VGND_M1025_d N_A_84_21#_M1027_g N_X_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1033 N_VGND_M1033_d N_A_84_21#_M1033_g N_X_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.175832 AS=0.1176 PD=1.40189 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75003.7 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1033_d N_S_M1010_g N_A_839_47#_M1010_s VNB NSHORT L=0.15 W=0.64
+ AD=0.133968 AS=0.0896 PD=1.06811 PS=0.92 NRD=22.02 NRS=0 M=1 R=4.26667
+ SA=75003.8 SB=75004.2 A=0.096 P=1.58 MULT=1
MM1016 N_A_839_47#_M1010_s N_A1_M1016_g N_A_84_21#_M1016_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75004.3 SB=75003.8 A=0.096 P=1.58 MULT=1
MM1019 N_A_839_47#_M1019_d N_A1_M1019_g N_A_84_21#_M1016_s VNB NSHORT L=0.15
+ W=0.64 AD=0.112 AS=0.112 PD=0.99 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75004.8 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_S_M1018_g N_A_839_47#_M1019_d VNB NSHORT L=0.15 W=0.64
+ AD=0.14515 AS=0.112 PD=1.11 PS=0.99 NRD=14.988 NRS=0 M=1 R=4.26667 SA=75005.3
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1018_d N_A_1179_311#_M1001_g N_A_1243_47#_M1001_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.14515 AS=0.0896 PD=1.11 PS=0.92 NRD=14.988 NRS=0 M=1
+ R=4.26667 SA=75005.9 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_1243_47#_M1001_s N_A0_M1008_g N_A_84_21#_M1008_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75006.3 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1029 N_A_1243_47#_M1029_d N_A0_M1029_g N_A_84_21#_M1008_s VNB NSHORT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75006.7 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_A_1179_311#_M1020_g N_A_1243_47#_M1029_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.159395 AS=0.112 PD=1.12865 PS=0.99 NRD=21.552 NRS=0 M=1
+ R=4.26667 SA=75007.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1030 N_A_1179_311#_M1030_d N_S_M1030_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.209205 PD=2.25 PS=1.48135 NRD=0 NRS=9.996 M=1 R=5.6 SA=75006
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_X_M1006_d N_A_84_21#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75006.9 A=0.189 P=2.82 MULT=1
MM1012 N_X_M1006_d N_A_84_21#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75006.5 A=0.189 P=2.82 MULT=1
MM1015 N_X_M1015_d N_A_84_21#_M1015_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1 SB=75006
+ A=0.189 P=2.82 MULT=1
MM1021 N_X_M1015_d N_A_84_21#_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75005.6 A=0.189 P=2.82 MULT=1
MM1022 N_X_M1022_d N_A_84_21#_M1022_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75005.2 A=0.189 P=2.82 MULT=1
MM1024 N_X_M1022_d N_A_84_21#_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1031 N_X_M1031_d N_A_84_21#_M1031_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1032 N_X_M1031_d N_A_84_21#_M1032_g N_VPWR_M1032_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.311711 PD=1.54 PS=1.94575 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75003.9 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1032_s N_S_M1007_g N_A_843_419#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.247389 AS=0.175 PD=1.54425 PS=1.35 NRD=40.3653 NRS=0 M=1 R=6.66667
+ SA=75003.9 SB=75004.2 A=0.15 P=2.3 MULT=1
MM1002 N_A_843_419#_M1007_s N_A0_M1002_g N_A_84_21#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.14 PD=1.35 PS=1.28 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75004.4 SB=75003.7 A=0.15 P=2.3 MULT=1
MM1028 N_A_843_419#_M1028_d N_A0_M1028_g N_A_84_21#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.14 PD=1.35 PS=1.28 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75004.8 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1023 N_VPWR_M1023_d N_S_M1023_g N_A_843_419#_M1028_d VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.175 PD=1.42 PS=1.35 NRD=13.7703 NRS=0 M=1 R=6.66667 SA=75005.3
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1023_d N_A_1179_311#_M1003_g N_A_1243_419#_M1003_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.21 AS=0.14 PD=1.42 PS=1.28 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75005.9 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1017 N_A_84_21#_M1017_d N_A1_M1017_g N_A_1243_419#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.14 PD=1.35 PS=1.28 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75006.3 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1026 N_A_84_21#_M1017_d N_A1_M1026_g N_A_1243_419#_M1026_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.18 PD=1.35 PS=1.36 NRD=0 NRS=13.7703 M=1 R=6.66667
+ SA=75006.8 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A_1179_311#_M1013_g N_A_1243_419#_M1026_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.207566 AS=0.18 PD=1.4646 PS=1.36 NRD=22.6353 NRS=1.9503 M=1
+ R=6.66667 SA=75007.3 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1000 N_A_1179_311#_M1000_d N_S_M1000_g N_VPWR_M1013_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.261534 PD=3.09 PS=1.8454 NRD=0 NRS=0 M=1 R=8.4
+ SA=75006.3 SB=75000.2 A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=16.8223 P=21.77
c_91 VNB 0 1.75633e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__mux2_8.pxi.spice"
*
.ends
*
*
