* File: sky130_fd_sc_lp__a32oi_0.pxi.spice
* Created: Wed Sep  2 09:28:08 2020
* 
x_PM_SKY130_FD_SC_LP__A32OI_0%B2 N_B2_M1001_g N_B2_M1005_g N_B2_c_71_n
+ N_B2_c_72_n B2 B2 B2 N_B2_c_74_n PM_SKY130_FD_SC_LP__A32OI_0%B2
x_PM_SKY130_FD_SC_LP__A32OI_0%B1 N_B1_M1008_g N_B1_M1002_g N_B1_c_100_n
+ N_B1_c_101_n N_B1_c_102_n B1 B1 N_B1_c_104_n PM_SKY130_FD_SC_LP__A32OI_0%B1
x_PM_SKY130_FD_SC_LP__A32OI_0%A1 N_A1_M1003_g N_A1_M1009_g N_A1_c_137_n
+ N_A1_c_145_n N_A1_c_138_n N_A1_c_139_n N_A1_c_140_n A1 A1 A1 N_A1_c_142_n
+ PM_SKY130_FD_SC_LP__A32OI_0%A1
x_PM_SKY130_FD_SC_LP__A32OI_0%A2 N_A2_M1006_g N_A2_M1004_g N_A2_c_187_n
+ N_A2_c_195_n N_A2_c_188_n N_A2_c_189_n N_A2_c_190_n A2 A2 A2 N_A2_c_192_n
+ PM_SKY130_FD_SC_LP__A32OI_0%A2
x_PM_SKY130_FD_SC_LP__A32OI_0%A3 N_A3_M1000_g N_A3_M1007_g N_A3_c_238_n
+ N_A3_c_239_n N_A3_c_240_n A3 A3 A3 N_A3_c_242_n PM_SKY130_FD_SC_LP__A32OI_0%A3
x_PM_SKY130_FD_SC_LP__A32OI_0%A_37_397# N_A_37_397#_M1001_s N_A_37_397#_M1008_d
+ N_A_37_397#_M1006_d N_A_37_397#_c_274_n N_A_37_397#_c_275_n
+ N_A_37_397#_c_276_n N_A_37_397#_c_277_n N_A_37_397#_c_272_n
+ N_A_37_397#_c_273_n N_A_37_397#_c_279_n PM_SKY130_FD_SC_LP__A32OI_0%A_37_397#
x_PM_SKY130_FD_SC_LP__A32OI_0%Y N_Y_M1002_d N_Y_M1001_d N_Y_c_328_n Y Y Y Y Y Y
+ N_Y_c_327_n PM_SKY130_FD_SC_LP__A32OI_0%Y
x_PM_SKY130_FD_SC_LP__A32OI_0%VPWR N_VPWR_M1003_d N_VPWR_M1000_d N_VPWR_c_352_n
+ N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_355_n VPWR N_VPWR_c_356_n
+ N_VPWR_c_357_n N_VPWR_c_351_n N_VPWR_c_359_n PM_SKY130_FD_SC_LP__A32OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A32OI_0%VGND N_VGND_M1005_s N_VGND_M1007_d N_VGND_c_384_n
+ N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n
+ VGND N_VGND_c_390_n PM_SKY130_FD_SC_LP__A32OI_0%VGND
cc_1 VNB N_B2_M1001_g 0.0091255f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.305
cc_2 VNB N_B2_M1005_g 0.0268588f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.445
cc_3 VNB N_B2_c_71_n 0.0307317f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.99
cc_4 VNB N_B2_c_72_n 0.0285232f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.51
cc_5 VNB B2 0.036127f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_B2_c_74_n 0.0290225f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.005
cc_7 VNB N_B1_M1008_g 0.0124565f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.305
cc_8 VNB N_B1_c_100_n 0.0238775f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=0.99
cc_9 VNB N_B1_c_101_n 0.021514f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.84
cc_10 VNB N_B1_c_102_n 0.0179886f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.293
cc_11 VNB B1 0.00934654f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.51
cc_12 VNB N_B1_c_104_n 0.0157584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_137_n 0.0138471f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=0.99
cc_14 VNB N_A1_c_138_n 0.0183409f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_A1_c_139_n 0.0217696f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_A1_c_140_n 0.015765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A1 0.00668277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_142_n 0.015833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_187_n 0.0132237f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.84
cc_20 VNB N_A2_c_188_n 0.0174664f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.51
cc_21 VNB N_A2_c_189_n 0.0213758f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_22 VNB N_A2_c_190_n 0.0155442f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB A2 0.00843985f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A2_c_192_n 0.0155459f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.925
cc_25 VNB N_A3_M1007_g 0.0272053f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.445
cc_26 VNB N_A3_c_238_n 0.0256967f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.84
cc_27 VNB N_A3_c_239_n 0.0101927f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.293
cc_28 VNB N_A3_c_240_n 0.0206797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB A3 0.0451587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A3_c_242_n 0.0210116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_37_397#_c_272_n 0.0181619f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.005
cc_32 VNB N_A_37_397#_c_273_n 0.0017359f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.005
cc_33 VNB Y 0.014549f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.99
cc_34 VNB N_VPWR_c_351_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_384_n 0.01403f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.445
cc_36 VNB N_VGND_c_385_n 0.0049188f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=0.99
cc_37 VNB N_VGND_c_386_n 0.0174842f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.51
cc_38 VNB N_VGND_c_387_n 0.0110534f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_39 VNB N_VGND_c_388_n 0.0599415f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_40 VNB N_VGND_c_389_n 0.00510915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_390_n 0.191295f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_42 VPB N_B2_M1001_g 0.0358849f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.305
cc_43 VPB B2 0.0112985f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_44 VPB N_B1_M1008_g 0.025933f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.305
cc_45 VPB N_A1_M1003_g 0.0226413f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.305
cc_46 VPB N_A1_c_137_n 0.00156371f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=0.99
cc_47 VPB N_A1_c_145_n 0.021992f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=1.293
cc_48 VPB N_A2_M1006_g 0.0232652f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.305
cc_49 VPB N_A2_c_187_n 9.76223e-19 $X=-0.19 $Y=1.655 $X2=0.435 $Y2=0.84
cc_50 VPB N_A2_c_195_n 0.00789836f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=0.99
cc_51 VPB N_A3_M1000_g 0.02468f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.305
cc_52 VPB N_A3_c_239_n 0.0238911f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=1.293
cc_53 VPB A3 0.0210094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_37_397#_c_274_n 0.0363045f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=1.293
cc_55 VPB N_A_37_397#_c_275_n 0.018019f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_56 VPB N_A_37_397#_c_276_n 0.0106885f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_57 VPB N_A_37_397#_c_277_n 0.00448712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_37_397#_c_272_n 0.00603665f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=1.005
cc_59 VPB N_A_37_397#_c_279_n 0.00775761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB Y 0.00931857f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=0.99
cc_61 VPB N_VPWR_c_352_n 0.0348565f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=0.99
cc_62 VPB N_VPWR_c_353_n 0.0604329f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=1.51
cc_63 VPB N_VPWR_c_354_n 0.0175089f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_64 VPB N_VPWR_c_355_n 0.00584071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_356_n 0.039809f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=1.005
cc_66 VPB N_VPWR_c_357_n 0.014713f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_351_n 0.0816147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_359_n 0.0116111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 N_B2_M1001_g N_B1_M1008_g 0.015125f $X=0.525 $Y=2.305 $X2=0 $Y2=0
cc_70 N_B2_c_74_n N_B1_c_100_n 0.00899992f $X=0.33 $Y=1.005 $X2=0 $Y2=0
cc_71 N_B2_c_72_n N_B1_c_101_n 0.015125f $X=0.382 $Y=1.51 $X2=0 $Y2=0
cc_72 N_B2_M1005_g N_B1_c_102_n 0.02371f $X=0.63 $Y=0.445 $X2=0 $Y2=0
cc_73 N_B2_c_71_n N_B1_c_104_n 0.02371f $X=0.435 $Y=0.99 $X2=0 $Y2=0
cc_74 N_B2_M1001_g N_A_37_397#_c_274_n 0.0107745f $X=0.525 $Y=2.305 $X2=0 $Y2=0
cc_75 N_B2_c_72_n N_A_37_397#_c_274_n 0.00120035f $X=0.382 $Y=1.51 $X2=0 $Y2=0
cc_76 B2 N_A_37_397#_c_274_n 0.0288223f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_77 N_B2_M1001_g N_A_37_397#_c_275_n 0.00676567f $X=0.525 $Y=2.305 $X2=0 $Y2=0
cc_78 N_B2_M1001_g N_A_37_397#_c_277_n 5.45526e-19 $X=0.525 $Y=2.305 $X2=0 $Y2=0
cc_79 N_B2_M1005_g Y 0.0123401f $X=0.63 $Y=0.445 $X2=0 $Y2=0
cc_80 N_B2_c_71_n Y 0.00614536f $X=0.435 $Y=0.99 $X2=0 $Y2=0
cc_81 B2 Y 0.073387f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_82 N_B2_c_74_n Y 0.0118956f $X=0.33 $Y=1.005 $X2=0 $Y2=0
cc_83 N_B2_M1005_g N_Y_c_327_n 0.00883332f $X=0.63 $Y=0.445 $X2=0 $Y2=0
cc_84 N_B2_M1005_g N_VGND_c_385_n 0.0123086f $X=0.63 $Y=0.445 $X2=0 $Y2=0
cc_85 N_B2_c_71_n N_VGND_c_385_n 0.00156551f $X=0.435 $Y=0.99 $X2=0 $Y2=0
cc_86 B2 N_VGND_c_385_n 0.0136703f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_87 N_B2_M1005_g N_VGND_c_388_n 0.0046505f $X=0.63 $Y=0.445 $X2=0 $Y2=0
cc_88 N_B2_M1005_g N_VGND_c_390_n 0.00906625f $X=0.63 $Y=0.445 $X2=0 $Y2=0
cc_89 N_B2_c_71_n N_VGND_c_390_n 0.00258418f $X=0.435 $Y=0.99 $X2=0 $Y2=0
cc_90 B2 N_VGND_c_390_n 0.00677726f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_91 N_B1_M1008_g N_A1_c_137_n 0.0058613f $X=0.955 $Y=2.305 $X2=0 $Y2=0
cc_92 N_B1_M1008_g N_A1_c_145_n 0.0178285f $X=0.955 $Y=2.305 $X2=0 $Y2=0
cc_93 B1 N_A1_c_145_n 3.17923e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_94 N_B1_c_102_n N_A1_c_138_n 0.0120136f $X=1.11 $Y=0.775 $X2=0 $Y2=0
cc_95 N_B1_c_100_n N_A1_c_139_n 0.0116888f $X=1.077 $Y=1.295 $X2=0 $Y2=0
cc_96 N_B1_c_101_n N_A1_c_140_n 0.0116888f $X=1.077 $Y=1.445 $X2=0 $Y2=0
cc_97 N_B1_c_102_n A1 6.00263e-19 $X=1.11 $Y=0.775 $X2=0 $Y2=0
cc_98 B1 A1 0.0528556f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_99 N_B1_c_104_n A1 7.01255e-19 $X=1.11 $Y=0.94 $X2=0 $Y2=0
cc_100 B1 N_A1_c_142_n 0.00415564f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_101 N_B1_c_104_n N_A1_c_142_n 0.0116888f $X=1.11 $Y=0.94 $X2=0 $Y2=0
cc_102 N_B1_M1008_g N_A_37_397#_c_274_n 4.9918e-19 $X=0.955 $Y=2.305 $X2=0 $Y2=0
cc_103 N_B1_M1008_g N_A_37_397#_c_275_n 0.00676567f $X=0.955 $Y=2.305 $X2=0
+ $Y2=0
cc_104 N_B1_M1008_g N_A_37_397#_c_277_n 0.0124109f $X=0.955 $Y=2.305 $X2=0 $Y2=0
cc_105 B1 N_A_37_397#_c_272_n 0.00495779f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_106 N_B1_M1008_g N_A_37_397#_c_273_n 0.00408763f $X=0.955 $Y=2.305 $X2=0
+ $Y2=0
cc_107 N_B1_c_101_n N_A_37_397#_c_273_n 0.00191752f $X=1.077 $Y=1.445 $X2=0
+ $Y2=0
cc_108 B1 N_A_37_397#_c_273_n 0.0244976f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_109 N_B1_c_102_n N_Y_c_328_n 0.0141437f $X=1.11 $Y=0.775 $X2=0 $Y2=0
cc_110 B1 N_Y_c_328_n 0.0231819f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_111 N_B1_c_104_n N_Y_c_328_n 0.0011555f $X=1.11 $Y=0.94 $X2=0 $Y2=0
cc_112 N_B1_c_101_n Y 0.00875198f $X=1.077 $Y=1.445 $X2=0 $Y2=0
cc_113 N_B1_c_102_n Y 0.00622783f $X=1.11 $Y=0.775 $X2=0 $Y2=0
cc_114 B1 Y 0.0515164f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_115 N_B1_c_102_n N_VGND_c_388_n 0.00359964f $X=1.11 $Y=0.775 $X2=0 $Y2=0
cc_116 N_B1_c_102_n N_VGND_c_390_n 0.00559721f $X=1.11 $Y=0.775 $X2=0 $Y2=0
cc_117 N_A1_M1003_g N_A2_M1006_g 0.00465302f $X=1.385 $Y=2.305 $X2=0 $Y2=0
cc_118 N_A1_c_145_n N_A2_M1006_g 0.00221895f $X=1.59 $Y=1.76 $X2=0 $Y2=0
cc_119 N_A1_c_137_n N_A2_c_187_n 0.00774804f $X=1.59 $Y=1.685 $X2=0 $Y2=0
cc_120 N_A1_c_137_n N_A2_c_195_n 0.00221895f $X=1.59 $Y=1.685 $X2=0 $Y2=0
cc_121 N_A1_c_138_n N_A2_c_188_n 0.0190693f $X=1.68 $Y=0.765 $X2=0 $Y2=0
cc_122 A1 N_A2_c_188_n 0.00322392f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_123 N_A1_c_139_n N_A2_c_189_n 0.0122475f $X=1.68 $Y=1.27 $X2=0 $Y2=0
cc_124 N_A1_c_140_n N_A2_c_190_n 0.0122475f $X=1.68 $Y=1.435 $X2=0 $Y2=0
cc_125 N_A1_c_138_n A2 9.94648e-19 $X=1.68 $Y=0.765 $X2=0 $Y2=0
cc_126 A1 A2 0.0884168f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_127 N_A1_c_142_n A2 0.00231413f $X=1.68 $Y=0.93 $X2=0 $Y2=0
cc_128 N_A1_c_142_n N_A2_c_192_n 0.0122475f $X=1.68 $Y=0.93 $X2=0 $Y2=0
cc_129 N_A1_c_145_n N_A_37_397#_c_277_n 0.00592164f $X=1.59 $Y=1.76 $X2=0 $Y2=0
cc_130 N_A1_c_137_n N_A_37_397#_c_272_n 0.0057537f $X=1.59 $Y=1.685 $X2=0 $Y2=0
cc_131 N_A1_c_145_n N_A_37_397#_c_272_n 0.0181057f $X=1.59 $Y=1.76 $X2=0 $Y2=0
cc_132 N_A1_c_140_n N_A_37_397#_c_272_n 0.00122246f $X=1.68 $Y=1.435 $X2=0 $Y2=0
cc_133 A1 N_A_37_397#_c_272_n 0.0258465f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_134 N_A1_c_138_n N_Y_c_328_n 0.00518981f $X=1.68 $Y=0.765 $X2=0 $Y2=0
cc_135 A1 N_Y_c_328_n 0.0172223f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 A1 Y 0.00465721f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_137 N_A1_M1003_g N_VPWR_c_352_n 0.00193181f $X=1.385 $Y=2.305 $X2=0 $Y2=0
cc_138 N_A1_c_145_n N_VPWR_c_352_n 0.00520779f $X=1.59 $Y=1.76 $X2=0 $Y2=0
cc_139 N_A1_M1003_g N_VPWR_c_356_n 0.00375548f $X=1.385 $Y=2.305 $X2=0 $Y2=0
cc_140 N_A1_M1003_g N_VPWR_c_351_n 0.00447875f $X=1.385 $Y=2.305 $X2=0 $Y2=0
cc_141 N_A1_c_138_n N_VGND_c_388_n 0.00404925f $X=1.68 $Y=0.765 $X2=0 $Y2=0
cc_142 A1 N_VGND_c_388_n 0.0108361f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A1_c_142_n N_VGND_c_388_n 4.47052e-19 $X=1.68 $Y=0.93 $X2=0 $Y2=0
cc_144 N_A1_c_138_n N_VGND_c_390_n 0.00680344f $X=1.68 $Y=0.765 $X2=0 $Y2=0
cc_145 A1 N_VGND_c_390_n 0.010838f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_146 A1 A_333_47# 0.00400992f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_147 N_A2_M1006_g N_A3_M1000_g 0.0107363f $X=2.155 $Y=2.305 $X2=0 $Y2=0
cc_148 N_A2_c_188_n N_A3_M1007_g 0.0191364f $X=2.25 $Y=0.765 $X2=0 $Y2=0
cc_149 A2 N_A3_M1007_g 0.00815601f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_150 N_A2_c_192_n N_A3_M1007_g 0.0136711f $X=2.25 $Y=0.93 $X2=0 $Y2=0
cc_151 N_A2_c_190_n N_A3_c_238_n 0.0136711f $X=2.25 $Y=1.435 $X2=0 $Y2=0
cc_152 N_A2_c_195_n N_A3_c_239_n 0.00627351f $X=2.157 $Y=1.825 $X2=0 $Y2=0
cc_153 N_A2_c_187_n N_A3_c_240_n 0.00737955f $X=2.157 $Y=1.675 $X2=0 $Y2=0
cc_154 N_A2_c_187_n A3 0.00105496f $X=2.157 $Y=1.675 $X2=0 $Y2=0
cc_155 A2 A3 0.0395404f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_156 N_A2_c_192_n A3 0.00215137f $X=2.25 $Y=0.93 $X2=0 $Y2=0
cc_157 N_A2_c_189_n N_A3_c_242_n 0.0136711f $X=2.25 $Y=1.27 $X2=0 $Y2=0
cc_158 N_A2_c_187_n N_A_37_397#_c_272_n 0.00448095f $X=2.157 $Y=1.675 $X2=0
+ $Y2=0
cc_159 N_A2_c_195_n N_A_37_397#_c_272_n 0.011677f $X=2.157 $Y=1.825 $X2=0 $Y2=0
cc_160 N_A2_c_190_n N_A_37_397#_c_272_n 0.00135185f $X=2.25 $Y=1.435 $X2=0 $Y2=0
cc_161 A2 N_A_37_397#_c_272_n 0.0335394f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_162 N_A2_M1006_g N_A_37_397#_c_279_n 0.00407311f $X=2.155 $Y=2.305 $X2=0
+ $Y2=0
cc_163 N_A2_c_195_n N_A_37_397#_c_279_n 7.89312e-19 $X=2.157 $Y=1.825 $X2=0
+ $Y2=0
cc_164 N_A2_M1006_g N_VPWR_c_352_n 0.00279061f $X=2.155 $Y=2.305 $X2=0 $Y2=0
cc_165 N_A2_M1006_g N_VPWR_c_354_n 0.00375548f $X=2.155 $Y=2.305 $X2=0 $Y2=0
cc_166 N_A2_M1006_g N_VPWR_c_351_n 0.00447875f $X=2.155 $Y=2.305 $X2=0 $Y2=0
cc_167 N_A2_c_188_n N_VGND_c_386_n 0.00177342f $X=2.25 $Y=0.765 $X2=0 $Y2=0
cc_168 A2 N_VGND_c_386_n 0.0105298f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_169 N_A2_c_188_n N_VGND_c_388_n 0.00383378f $X=2.25 $Y=0.765 $X2=0 $Y2=0
cc_170 A2 N_VGND_c_388_n 0.0126457f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_171 N_A2_c_192_n N_VGND_c_388_n 4.44569e-19 $X=2.25 $Y=0.93 $X2=0 $Y2=0
cc_172 N_A2_c_188_n N_VGND_c_390_n 0.00615839f $X=2.25 $Y=0.765 $X2=0 $Y2=0
cc_173 A2 N_VGND_c_390_n 0.0134705f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_174 A2 A_333_47# 0.00258003f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_175 A2 A_447_47# 0.0047341f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_176 N_A3_c_239_n N_A_37_397#_c_272_n 0.00161511f $X=2.715 $Y=1.675 $X2=0
+ $Y2=0
cc_177 A3 N_A_37_397#_c_272_n 0.0158141f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_178 N_A3_c_239_n N_A_37_397#_c_279_n 0.00484644f $X=2.715 $Y=1.675 $X2=0
+ $Y2=0
cc_179 N_A3_M1000_g N_VPWR_c_353_n 0.00426613f $X=2.585 $Y=2.305 $X2=0 $Y2=0
cc_180 N_A3_c_239_n N_VPWR_c_353_n 0.00406235f $X=2.715 $Y=1.675 $X2=0 $Y2=0
cc_181 N_A3_c_240_n N_VPWR_c_353_n 6.69666e-19 $X=2.805 $Y=1.51 $X2=0 $Y2=0
cc_182 A3 N_VPWR_c_353_n 0.0277354f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_183 N_A3_M1000_g N_VPWR_c_354_n 0.00374771f $X=2.585 $Y=2.305 $X2=0 $Y2=0
cc_184 N_A3_M1000_g N_VPWR_c_351_n 0.00447875f $X=2.585 $Y=2.305 $X2=0 $Y2=0
cc_185 N_A3_M1007_g N_VGND_c_386_n 0.0126738f $X=2.7 $Y=0.445 $X2=0 $Y2=0
cc_186 A3 N_VGND_c_386_n 0.0265516f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_187 N_A3_c_242_n N_VGND_c_386_n 0.0012464f $X=2.82 $Y=1.005 $X2=0 $Y2=0
cc_188 N_A3_M1007_g N_VGND_c_388_n 0.00486043f $X=2.7 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A3_M1007_g N_VGND_c_390_n 0.0058833f $X=2.7 $Y=0.445 $X2=0 $Y2=0
cc_190 A3 N_VGND_c_390_n 0.0124473f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_191 N_A_37_397#_c_274_n Y 0.0267689f $X=0.31 $Y=2.13 $X2=0 $Y2=0
cc_192 N_A_37_397#_c_275_n Y 0.0183356f $X=1.025 $Y=2.9 $X2=0 $Y2=0
cc_193 N_A_37_397#_c_277_n Y 0.0391723f $X=1.17 $Y=2.13 $X2=0 $Y2=0
cc_194 N_A_37_397#_c_273_n Y 0.0147023f $X=1.3 $Y=1.705 $X2=0 $Y2=0
cc_195 N_A_37_397#_c_275_n N_VPWR_c_352_n 0.0157199f $X=1.025 $Y=2.9 $X2=0 $Y2=0
cc_196 N_A_37_397#_c_277_n N_VPWR_c_352_n 0.0178647f $X=1.17 $Y=2.13 $X2=0 $Y2=0
cc_197 N_A_37_397#_c_272_n N_VPWR_c_352_n 0.0503893f $X=2.245 $Y=1.705 $X2=0
+ $Y2=0
cc_198 N_A_37_397#_c_279_n N_VPWR_c_352_n 0.00324376f $X=2.37 $Y=2.13 $X2=0
+ $Y2=0
cc_199 N_A_37_397#_c_279_n N_VPWR_c_353_n 0.0293845f $X=2.37 $Y=2.13 $X2=0 $Y2=0
cc_200 N_A_37_397#_c_279_n N_VPWR_c_354_n 0.00445166f $X=2.37 $Y=2.13 $X2=0
+ $Y2=0
cc_201 N_A_37_397#_c_275_n N_VPWR_c_356_n 0.0359482f $X=1.025 $Y=2.9 $X2=0 $Y2=0
cc_202 N_A_37_397#_c_276_n N_VPWR_c_356_n 0.0141155f $X=0.455 $Y=2.9 $X2=0 $Y2=0
cc_203 N_A_37_397#_c_275_n N_VPWR_c_351_n 0.0304026f $X=1.025 $Y=2.9 $X2=0 $Y2=0
cc_204 N_A_37_397#_c_276_n N_VPWR_c_351_n 0.0114836f $X=0.455 $Y=2.9 $X2=0 $Y2=0
cc_205 N_A_37_397#_c_279_n N_VPWR_c_351_n 0.00710663f $X=2.37 $Y=2.13 $X2=0
+ $Y2=0
cc_206 Y N_VGND_c_385_n 0.00105928f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_207 N_Y_c_327_n N_VGND_c_385_n 0.0263248f $X=0.74 $Y=0.595 $X2=0 $Y2=0
cc_208 N_Y_c_328_n N_VGND_c_388_n 0.0278274f $X=1.26 $Y=0.43 $X2=0 $Y2=0
cc_209 N_Y_c_327_n N_VGND_c_388_n 0.0131705f $X=0.74 $Y=0.595 $X2=0 $Y2=0
cc_210 N_Y_M1002_d N_VGND_c_390_n 0.00877646f $X=1.095 $Y=0.235 $X2=0 $Y2=0
cc_211 N_Y_c_328_n N_VGND_c_390_n 0.0184001f $X=1.26 $Y=0.43 $X2=0 $Y2=0
cc_212 N_Y_c_327_n N_VGND_c_390_n 0.00853094f $X=0.74 $Y=0.595 $X2=0 $Y2=0
cc_213 N_Y_c_328_n A_141_47# 0.00163637f $X=1.26 $Y=0.43 $X2=-0.19 $Y2=-0.245
cc_214 Y A_141_47# 8.59879e-19 $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_215 N_Y_c_327_n A_141_47# 9.29739e-19 $X=0.74 $Y=0.595 $X2=-0.19 $Y2=-0.245
cc_216 N_VGND_c_390_n A_141_47# 0.00193237f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_217 N_VGND_c_390_n A_333_47# 0.00949073f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_218 N_VGND_c_390_n A_447_47# 0.0105477f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
