* File: sky130_fd_sc_lp__o211a_0.pxi.spice
* Created: Fri Aug 28 11:01:37 2020
* 
x_PM_SKY130_FD_SC_LP__O211A_0%A_80_21# N_A_80_21#_M1008_d N_A_80_21#_M1000_d
+ N_A_80_21#_M1006_d N_A_80_21#_M1003_g N_A_80_21#_c_81_n N_A_80_21#_c_82_n
+ N_A_80_21#_c_83_n N_A_80_21#_M1005_g N_A_80_21#_c_85_n N_A_80_21#_c_86_n
+ N_A_80_21#_c_87_n N_A_80_21#_c_88_n N_A_80_21#_c_75_n N_A_80_21#_c_118_p
+ N_A_80_21#_c_76_n N_A_80_21#_c_77_n N_A_80_21#_c_78_n N_A_80_21#_c_79_n
+ N_A_80_21#_c_90_n N_A_80_21#_c_91_n N_A_80_21#_c_92_n N_A_80_21#_c_93_n
+ PM_SKY130_FD_SC_LP__O211A_0%A_80_21#
x_PM_SKY130_FD_SC_LP__O211A_0%A1 N_A1_M1007_g N_A1_M1002_g N_A1_c_179_n
+ N_A1_c_180_n A1 N_A1_c_181_n PM_SKY130_FD_SC_LP__O211A_0%A1
x_PM_SKY130_FD_SC_LP__O211A_0%A2 N_A2_M1000_g N_A2_M1001_g N_A2_c_217_n
+ N_A2_c_222_n A2 A2 N_A2_c_219_n PM_SKY130_FD_SC_LP__O211A_0%A2
x_PM_SKY130_FD_SC_LP__O211A_0%B1 N_B1_M1009_g N_B1_M1004_g N_B1_c_266_n
+ N_B1_c_267_n B1 N_B1_c_264_n PM_SKY130_FD_SC_LP__O211A_0%B1
x_PM_SKY130_FD_SC_LP__O211A_0%C1 N_C1_c_315_n N_C1_M1008_g N_C1_M1006_g
+ N_C1_c_316_n N_C1_c_321_n C1 N_C1_c_318_n PM_SKY130_FD_SC_LP__O211A_0%C1
x_PM_SKY130_FD_SC_LP__O211A_0%X N_X_M1003_s N_X_M1005_s N_X_c_353_n X X X X X X
+ N_X_c_352_n PM_SKY130_FD_SC_LP__O211A_0%X
x_PM_SKY130_FD_SC_LP__O211A_0%VPWR N_VPWR_M1005_d N_VPWR_M1009_d N_VPWR_c_372_n
+ N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_375_n VPWR N_VPWR_c_376_n
+ N_VPWR_c_377_n N_VPWR_c_371_n N_VPWR_c_379_n PM_SKY130_FD_SC_LP__O211A_0%VPWR
x_PM_SKY130_FD_SC_LP__O211A_0%VGND N_VGND_M1003_d N_VGND_M1007_d N_VGND_c_411_n
+ N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n VGND N_VGND_c_415_n
+ N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n PM_SKY130_FD_SC_LP__O211A_0%VGND
x_PM_SKY130_FD_SC_LP__O211A_0%A_257_47# N_A_257_47#_M1007_s N_A_257_47#_M1001_d
+ N_A_257_47#_c_452_n N_A_257_47#_c_453_n N_A_257_47#_c_454_n
+ N_A_257_47#_c_455_n PM_SKY130_FD_SC_LP__O211A_0%A_257_47#
cc_1 VNB N_A_80_21#_M1003_g 0.0900101f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_80_21#_c_75_n 0.00629264f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=1.19
cc_3 VNB N_A_80_21#_c_76_n 0.0143447f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=0.445
cc_4 VNB N_A_80_21#_c_77_n 0.0137079f $X=-0.19 $Y=-0.245 $X2=2.935 $Y2=1.275
cc_5 VNB N_A_80_21#_c_78_n 8.77593e-19 $X=-0.19 $Y=-0.245 $X2=2.745 $Y2=1.275
cc_6 VNB N_A_80_21#_c_79_n 0.0135033f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=2.05
cc_7 VNB N_A1_M1007_g 0.0517292f $X=-0.19 $Y=-0.245 $X2=2.96 $Y2=2.425
cc_8 VNB N_A1_M1002_g 0.00705502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_c_179_n 0.0529879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_180_n 0.00859385f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.935
cc_11 VNB N_A1_c_181_n 0.0203069f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.1
cc_12 VNB N_A2_M1001_g 0.0371011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_217_n 0.0200345f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_14 VNB A2 0.00559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_219_n 0.0152508f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.745
cc_16 VNB N_B1_M1004_g 0.0536712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_264_n 0.0191311f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.265
cc_18 VNB N_C1_c_315_n 0.0216031f $X=-0.19 $Y=-0.245 $X2=2.96 $Y2=0.235
cc_19 VNB N_C1_c_316_n 0.0352659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB C1 0.00906297f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=2.1
cc_21 VNB N_C1_c_318_n 0.0462317f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=2.085
cc_22 VNB N_X_c_352_n 0.0717009f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=2.55
cc_23 VNB N_VPWR_c_371_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=1.19
cc_24 VNB N_VGND_c_411_n 0.0104144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_412_n 0.00245823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_413_n 0.0247725f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.265
cc_27 VNB N_VGND_c_414_n 0.00382174f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.745
cc_28 VNB N_VGND_c_415_n 0.0158747f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=2.085
cc_29 VNB N_VGND_c_416_n 0.0359999f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.605
cc_30 VNB N_VGND_c_417_n 0.204189f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=1.19
cc_31 VNB N_VGND_c_418_n 0.00522775f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=0.445
cc_32 VNB N_A_257_47#_c_452_n 0.0115434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_257_47#_c_453_n 0.0189335f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_34 VNB N_A_257_47#_c_454_n 0.00956178f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_35 VNB N_A_257_47#_c_455_n 0.00205578f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.1
cc_36 VPB N_A_80_21#_M1003_g 0.0234929f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_37 VPB N_A_80_21#_c_81_n 0.0533484f $X=-0.19 $Y=1.655 $X2=1.04 $Y2=2.1
cc_38 VPB N_A_80_21#_c_82_n 0.0173283f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.1
cc_39 VPB N_A_80_21#_c_83_n 0.0167418f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.265
cc_40 VPB N_A_80_21#_M1005_g 0.0248424f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.745
cc_41 VPB N_A_80_21#_c_85_n 0.00693875f $X=-0.19 $Y=1.655 $X2=1.64 $Y2=2.085
cc_42 VPB N_A_80_21#_c_86_n 0.00826171f $X=-0.19 $Y=1.655 $X2=2.065 $Y2=2.142
cc_43 VPB N_A_80_21#_c_87_n 0.00553454f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=2.55
cc_44 VPB N_A_80_21#_c_88_n 0.0131496f $X=-0.19 $Y=1.655 $X2=2.935 $Y2=2.142
cc_45 VPB N_A_80_21#_c_79_n 0.0181406f $X=-0.19 $Y=1.655 $X2=3.1 $Y2=2.05
cc_46 VPB N_A_80_21#_c_90_n 0.0345651f $X=-0.19 $Y=1.655 $X2=3.1 $Y2=2.57
cc_47 VPB N_A_80_21#_c_91_n 0.00788871f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=2.085
cc_48 VPB N_A_80_21#_c_92_n 0.00385957f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=2.142
cc_49 VPB N_A_80_21#_c_93_n 0.00753458f $X=-0.19 $Y=1.655 $X2=3.1 $Y2=2.142
cc_50 VPB N_A1_M1002_g 0.0554373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A2_M1000_g 0.040205f $X=-0.19 $Y=1.655 $X2=2.96 $Y2=2.425
cc_52 VPB N_A2_c_217_n 8.67025e-19 $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_53 VPB N_A2_c_222_n 0.015356f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_54 VPB A2 0.00332574f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B1_M1009_g 0.0215558f $X=-0.19 $Y=1.655 $X2=2.96 $Y2=2.425
cc_56 VPB N_B1_c_266_n 0.0135195f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_57 VPB N_B1_c_267_n 0.0112617f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_58 VPB B1 0.00158058f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_B1_c_264_n 0.0235502f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.265
cc_60 VPB N_C1_M1006_g 0.0262892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_C1_c_316_n 0.0229135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_C1_c_321_n 0.0276222f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_63 VPB N_X_c_353_n 0.0129164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB X 0.0362498f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.265
cc_65 VPB N_X_c_352_n 0.0420192f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=2.55
cc_66 VPB N_VPWR_c_372_n 0.00666645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_373_n 0.00491245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_374_n 0.0324346f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.265
cc_69 VPB N_VPWR_c_375_n 0.00533588f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.745
cc_70 VPB N_VPWR_c_376_n 0.025311f $X=-0.19 $Y=1.655 $X2=2.2 $Y2=2.235
cc_71 VPB N_VPWR_c_377_n 0.0178672f $X=-0.19 $Y=1.655 $X2=2.66 $Y2=0.605
cc_72 VPB N_VPWR_c_371_n 0.0699969f $X=-0.19 $Y=1.655 $X2=2.66 $Y2=1.19
cc_73 VPB N_VPWR_c_379_n 0.00398612f $X=-0.19 $Y=1.655 $X2=3.1 $Y2=0.445
cc_74 N_A_80_21#_c_83_n N_A1_M1002_g 0.0122671f $X=1.115 $Y=2.265 $X2=0 $Y2=0
cc_75 N_A_80_21#_M1005_g N_A1_M1002_g 0.0183511f $X=1.115 $Y=2.745 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_85_n N_A1_M1002_g 0.0118312f $X=1.64 $Y=2.085 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_91_n N_A1_M1002_g 0.00791788f $X=1.79 $Y=2.085 $X2=0 $Y2=0
cc_78 N_A_80_21#_M1003_g N_A1_c_179_n 0.00673588f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_81_n N_A1_c_179_n 0.00590616f $X=1.04 $Y=2.1 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_85_n N_A1_c_179_n 0.00739601f $X=1.64 $Y=2.085 $X2=0 $Y2=0
cc_81 N_A_80_21#_M1003_g N_A1_c_181_n 0.00330558f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_81_n N_A1_c_181_n 8.69649e-19 $X=1.04 $Y=2.1 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_85_n N_A1_c_181_n 0.0286844f $X=1.64 $Y=2.085 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_86_n N_A2_M1000_g 0.0171659f $X=2.065 $Y=2.142 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_87_n N_A2_M1000_g 0.00519389f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_91_n N_A2_M1000_g 0.00323658f $X=1.79 $Y=2.085 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_75_n N_A2_M1001_g 0.00121488f $X=2.66 $Y=1.19 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_92_n N_A2_c_222_n 0.00133168f $X=2.2 $Y=2.142 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_86_n A2 0.00657631f $X=2.065 $Y=2.142 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_75_n A2 0.00122911f $X=2.66 $Y=1.19 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_78_n A2 0.0094194f $X=2.745 $Y=1.275 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_79_n A2 0.00542422f $X=3.1 $Y=2.05 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_92_n A2 0.016142f $X=2.2 $Y=2.142 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_87_n N_B1_M1009_g 0.00261146f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_88_n N_B1_M1009_g 0.00626693f $X=2.935 $Y=2.142 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_90_n N_B1_M1009_g 7.17137e-19 $X=3.1 $Y=2.57 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_75_n N_B1_M1004_g 0.011804f $X=2.66 $Y=1.19 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_118_p N_B1_M1004_g 0.00646562f $X=2.745 $Y=0.442 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_78_n N_B1_M1004_g 0.00551928f $X=2.745 $Y=1.275 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_79_n N_B1_M1004_g 0.00140705f $X=3.1 $Y=2.05 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_88_n N_B1_c_266_n 0.00328243f $X=2.935 $Y=2.142 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_79_n N_B1_c_266_n 0.00467493f $X=3.1 $Y=2.05 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_88_n N_B1_c_267_n 0.00840444f $X=2.935 $Y=2.142 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_88_n B1 0.0213007f $X=2.935 $Y=2.142 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_77_n B1 0.00139717f $X=2.935 $Y=1.275 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_78_n B1 0.0142935f $X=2.745 $Y=1.275 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_79_n B1 0.0260243f $X=3.1 $Y=2.05 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_88_n N_B1_c_264_n 0.00438364f $X=2.935 $Y=2.142 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_77_n N_B1_c_264_n 0.00404167f $X=2.935 $Y=1.275 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_78_n N_B1_c_264_n 0.00356057f $X=2.745 $Y=1.275 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_79_n N_B1_c_264_n 0.00289406f $X=3.1 $Y=2.05 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_75_n N_C1_c_315_n 0.00728647f $X=2.66 $Y=1.19 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_80_21#_c_76_n N_C1_c_315_n 0.0120417f $X=3.1 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_80_21#_c_88_n N_C1_M1006_g 0.00579527f $X=2.935 $Y=2.142 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_90_n N_C1_M1006_g 0.0140893f $X=3.1 $Y=2.57 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_93_n N_C1_M1006_g 3.15806e-19 $X=3.1 $Y=2.142 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_77_n N_C1_c_316_n 0.00996861f $X=2.935 $Y=1.275 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_79_n N_C1_c_316_n 0.0246505f $X=3.1 $Y=2.05 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_93_n N_C1_c_316_n 5.39195e-19 $X=3.1 $Y=2.142 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_88_n N_C1_c_321_n 0.00394658f $X=2.935 $Y=2.142 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_93_n N_C1_c_321_n 0.0174202f $X=3.1 $Y=2.142 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_75_n C1 0.0183508f $X=2.66 $Y=1.19 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_76_n C1 0.0218795f $X=3.1 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_77_n C1 0.026376f $X=2.935 $Y=1.275 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_76_n N_C1_c_318_n 0.00701705f $X=3.1 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_77_n N_C1_c_318_n 0.00689647f $X=2.935 $Y=1.275 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_82_n N_X_c_353_n 0.0190802f $X=0.55 $Y=2.1 $X2=0 $Y2=0
cc_128 N_A_80_21#_M1005_g N_X_c_353_n 0.00821273f $X=1.115 $Y=2.745 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_85_n N_X_c_353_n 0.043124f $X=1.64 $Y=2.085 $X2=0 $Y2=0
cc_130 N_A_80_21#_M1003_g N_X_c_352_n 0.0596873f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_80_21#_M1005_g N_X_c_352_n 0.00300342f $X=1.115 $Y=2.745 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_85_n N_X_c_352_n 0.0236481f $X=1.64 $Y=2.085 $X2=0 $Y2=0
cc_133 N_A_80_21#_M1005_g N_VPWR_c_372_n 0.00641097f $X=1.115 $Y=2.745 $X2=0
+ $Y2=0
cc_134 N_A_80_21#_c_85_n N_VPWR_c_372_n 0.028613f $X=1.64 $Y=2.085 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_87_n N_VPWR_c_372_n 0.0111501f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_87_n N_VPWR_c_373_n 0.0253683f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_88_n N_VPWR_c_373_n 0.0217158f $X=2.935 $Y=2.142 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_90_n N_VPWR_c_373_n 0.0262636f $X=3.1 $Y=2.57 $X2=0 $Y2=0
cc_139 N_A_80_21#_M1005_g N_VPWR_c_374_n 0.0051909f $X=1.115 $Y=2.745 $X2=0
+ $Y2=0
cc_140 N_A_80_21#_c_87_n N_VPWR_c_376_n 0.019212f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_141 N_A_80_21#_c_90_n N_VPWR_c_377_n 0.0234289f $X=3.1 $Y=2.57 $X2=0 $Y2=0
cc_142 N_A_80_21#_M1005_g N_VPWR_c_371_n 0.0108775f $X=1.115 $Y=2.745 $X2=0
+ $Y2=0
cc_143 N_A_80_21#_c_87_n N_VPWR_c_371_n 0.0104192f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_144 N_A_80_21#_c_90_n N_VPWR_c_371_n 0.0126421f $X=3.1 $Y=2.57 $X2=0 $Y2=0
cc_145 N_A_80_21#_M1003_g N_VGND_c_411_n 0.00993967f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_146 N_A_80_21#_M1003_g N_VGND_c_415_n 0.00564095f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_147 N_A_80_21#_c_118_p N_VGND_c_416_n 0.00855533f $X=2.745 $Y=0.442 $X2=0
+ $Y2=0
cc_148 N_A_80_21#_c_76_n N_VGND_c_416_n 0.02642f $X=3.1 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_80_21#_M1008_d N_VGND_c_417_n 0.0021695f $X=2.96 $Y=0.235 $X2=0 $Y2=0
cc_150 N_A_80_21#_M1003_g N_VGND_c_417_n 0.010595f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_151 N_A_80_21#_c_118_p N_VGND_c_417_n 0.00641269f $X=2.745 $Y=0.442 $X2=0
+ $Y2=0
cc_152 N_A_80_21#_c_76_n N_VGND_c_417_n 0.0188517f $X=3.1 $Y=0.445 $X2=0 $Y2=0
cc_153 N_A_80_21#_c_75_n N_A_257_47#_c_453_n 0.013714f $X=2.66 $Y=1.19 $X2=0
+ $Y2=0
cc_154 N_A_80_21#_c_75_n N_A_257_47#_c_455_n 0.010742f $X=2.66 $Y=1.19 $X2=0
+ $Y2=0
cc_155 N_A_80_21#_c_75_n A_520_47# 5.39753e-19 $X=2.66 $Y=1.19 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_80_21#_c_118_p A_520_47# 9.08637e-19 $X=2.745 $Y=0.442 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A1_M1007_g N_A2_M1001_g 0.0295778f $X=1.625 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A1_c_181_n N_A2_M1001_g 2.68738e-19 $X=1.535 $Y=1.4 $X2=0 $Y2=0
cc_159 N_A1_c_180_n N_A2_c_217_n 0.0415362f $X=1.625 $Y=1.4 $X2=0 $Y2=0
cc_160 N_A1_M1002_g N_A2_c_222_n 0.0415362f $X=1.625 $Y=2.745 $X2=0 $Y2=0
cc_161 N_A1_M1007_g A2 4.63497e-19 $X=1.625 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A1_c_180_n A2 0.00159504f $X=1.625 $Y=1.4 $X2=0 $Y2=0
cc_163 N_A1_c_181_n A2 0.0225106f $X=1.535 $Y=1.4 $X2=0 $Y2=0
cc_164 N_A1_M1007_g N_A2_c_219_n 0.0415362f $X=1.625 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A1_c_181_n N_A2_c_219_n 0.00143705f $X=1.535 $Y=1.4 $X2=0 $Y2=0
cc_166 N_A1_c_181_n N_X_c_352_n 0.0132415f $X=1.535 $Y=1.4 $X2=0 $Y2=0
cc_167 N_A1_M1002_g N_VPWR_c_372_n 0.0161481f $X=1.625 $Y=2.745 $X2=0 $Y2=0
cc_168 N_A1_M1002_g N_VPWR_c_376_n 0.00461019f $X=1.625 $Y=2.745 $X2=0 $Y2=0
cc_169 N_A1_M1002_g N_VPWR_c_371_n 0.00806991f $X=1.625 $Y=2.745 $X2=0 $Y2=0
cc_170 N_A1_M1007_g N_VGND_c_411_n 0.00209611f $X=1.625 $Y=0.445 $X2=0 $Y2=0
cc_171 N_A1_M1007_g N_VGND_c_412_n 0.0029706f $X=1.625 $Y=0.445 $X2=0 $Y2=0
cc_172 N_A1_M1007_g N_VGND_c_413_n 0.0054978f $X=1.625 $Y=0.445 $X2=0 $Y2=0
cc_173 N_A1_M1007_g N_VGND_c_417_n 0.0075204f $X=1.625 $Y=0.445 $X2=0 $Y2=0
cc_174 N_A1_M1007_g N_A_257_47#_c_452_n 0.00950528f $X=1.625 $Y=0.445 $X2=0
+ $Y2=0
cc_175 N_A1_M1007_g N_A_257_47#_c_453_n 0.00842533f $X=1.625 $Y=0.445 $X2=0
+ $Y2=0
cc_176 N_A1_c_181_n N_A_257_47#_c_453_n 0.00911218f $X=1.535 $Y=1.4 $X2=0 $Y2=0
cc_177 N_A1_M1007_g N_A_257_47#_c_454_n 0.00415614f $X=1.625 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_A1_c_179_n N_A_257_47#_c_454_n 0.00174359f $X=1.55 $Y=1.4 $X2=0 $Y2=0
cc_179 N_A1_c_181_n N_A_257_47#_c_454_n 0.0286708f $X=1.535 $Y=1.4 $X2=0 $Y2=0
cc_180 N_A2_M1001_g N_B1_M1004_g 0.0254429f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_181 A2 N_B1_M1004_g 0.00492029f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A2_c_219_n N_B1_M1004_g 0.020545f $X=2.075 $Y=1.33 $X2=0 $Y2=0
cc_183 N_A2_M1000_g N_B1_c_267_n 0.0169673f $X=1.985 $Y=2.745 $X2=0 $Y2=0
cc_184 N_A2_c_217_n B1 3.51399e-19 $X=2.075 $Y=1.67 $X2=0 $Y2=0
cc_185 A2 B1 0.0239973f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A2_M1000_g N_B1_c_264_n 0.00823265f $X=1.985 $Y=2.745 $X2=0 $Y2=0
cc_187 N_A2_c_217_n N_B1_c_264_n 0.020545f $X=2.075 $Y=1.67 $X2=0 $Y2=0
cc_188 N_A2_M1000_g N_VPWR_c_372_n 0.00283315f $X=1.985 $Y=2.745 $X2=0 $Y2=0
cc_189 N_A2_M1000_g N_VPWR_c_373_n 0.00101021f $X=1.985 $Y=2.745 $X2=0 $Y2=0
cc_190 N_A2_M1000_g N_VPWR_c_376_n 0.00555245f $X=1.985 $Y=2.745 $X2=0 $Y2=0
cc_191 N_A2_M1000_g N_VPWR_c_371_n 0.0106189f $X=1.985 $Y=2.745 $X2=0 $Y2=0
cc_192 N_A2_M1001_g N_VGND_c_412_n 0.00849104f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_193 N_A2_M1001_g N_VGND_c_416_n 0.00525069f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A2_M1001_g N_VGND_c_417_n 0.00490838f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_195 N_A2_M1001_g N_A_257_47#_c_452_n 4.49912e-19 $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_196 N_A2_M1001_g N_A_257_47#_c_453_n 0.0116775f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_197 A2 N_A_257_47#_c_453_n 0.0216226f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_198 N_A2_c_219_n N_A_257_47#_c_453_n 0.00292972f $X=2.075 $Y=1.33 $X2=0 $Y2=0
cc_199 N_A2_M1001_g N_A_257_47#_c_455_n 0.00178535f $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_200 N_B1_M1004_g N_C1_c_315_n 0.0629153f $X=2.525 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_201 N_B1_M1009_g N_C1_M1006_g 0.0142594f $X=2.455 $Y=2.745 $X2=0 $Y2=0
cc_202 N_B1_c_267_n N_C1_M1006_g 0.004992f $X=2.49 $Y=2.225 $X2=0 $Y2=0
cc_203 N_B1_M1004_g N_C1_c_316_n 0.00598168f $X=2.525 $Y=0.445 $X2=0 $Y2=0
cc_204 N_B1_c_266_n N_C1_c_316_n 0.00218755f $X=2.49 $Y=2.075 $X2=0 $Y2=0
cc_205 B1 N_C1_c_316_n 2.57692e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_206 N_B1_c_264_n N_C1_c_316_n 0.0225734f $X=2.615 $Y=1.695 $X2=0 $Y2=0
cc_207 N_B1_c_266_n N_C1_c_321_n 0.004992f $X=2.49 $Y=2.075 $X2=0 $Y2=0
cc_208 N_B1_c_264_n N_C1_c_321_n 0.00475274f $X=2.615 $Y=1.695 $X2=0 $Y2=0
cc_209 N_B1_c_264_n N_C1_c_318_n 0.00185094f $X=2.615 $Y=1.695 $X2=0 $Y2=0
cc_210 N_B1_M1009_g N_VPWR_c_373_n 0.0115393f $X=2.455 $Y=2.745 $X2=0 $Y2=0
cc_211 N_B1_c_267_n N_VPWR_c_373_n 5.33265e-19 $X=2.49 $Y=2.225 $X2=0 $Y2=0
cc_212 N_B1_M1009_g N_VPWR_c_376_n 0.00461019f $X=2.455 $Y=2.745 $X2=0 $Y2=0
cc_213 N_B1_M1009_g N_VPWR_c_371_n 0.00830259f $X=2.455 $Y=2.745 $X2=0 $Y2=0
cc_214 N_B1_M1004_g N_VGND_c_412_n 0.00118445f $X=2.525 $Y=0.445 $X2=0 $Y2=0
cc_215 N_B1_M1004_g N_VGND_c_416_n 0.00548296f $X=2.525 $Y=0.445 $X2=0 $Y2=0
cc_216 N_B1_M1004_g N_VGND_c_417_n 0.00999102f $X=2.525 $Y=0.445 $X2=0 $Y2=0
cc_217 N_B1_M1004_g N_A_257_47#_c_453_n 0.00147037f $X=2.525 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_B1_M1004_g N_A_257_47#_c_455_n 0.00103182f $X=2.525 $Y=0.445 $X2=0
+ $Y2=0
cc_219 N_C1_M1006_g N_VPWR_c_373_n 0.00286f $X=2.885 $Y=2.745 $X2=0 $Y2=0
cc_220 N_C1_M1006_g N_VPWR_c_377_n 0.00520505f $X=2.885 $Y=2.745 $X2=0 $Y2=0
cc_221 N_C1_M1006_g N_VPWR_c_371_n 0.0104236f $X=2.885 $Y=2.745 $X2=0 $Y2=0
cc_222 N_C1_c_315_n N_VGND_c_416_n 0.00363059f $X=2.885 $Y=0.765 $X2=0 $Y2=0
cc_223 N_C1_c_315_n N_VGND_c_417_n 0.0062645f $X=2.885 $Y=0.765 $X2=0 $Y2=0
cc_224 N_X_c_353_n N_VPWR_c_372_n 0.0279139f $X=0.9 $Y=2.57 $X2=0 $Y2=0
cc_225 N_X_c_353_n N_VPWR_c_374_n 0.0496752f $X=0.9 $Y=2.57 $X2=0 $Y2=0
cc_226 X N_VPWR_c_374_n 0.0199999f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_227 N_X_c_353_n N_VPWR_c_371_n 0.0270691f $X=0.9 $Y=2.57 $X2=0 $Y2=0
cc_228 X N_VPWR_c_371_n 0.0108752f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_229 N_X_c_352_n N_VGND_c_415_n 0.0177488f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_230 N_X_M1003_s N_VGND_c_417_n 0.00341412f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_231 N_X_c_352_n N_VGND_c_417_n 0.0107567f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_232 N_VGND_c_417_n N_A_257_47#_M1007_s 0.00216892f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_233 N_VGND_c_417_n N_A_257_47#_M1001_d 0.00429378f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_411_n N_A_257_47#_c_452_n 0.015964f $X=0.69 $Y=0.445 $X2=0 $Y2=0
cc_235 N_VGND_c_413_n N_A_257_47#_c_452_n 0.0175133f $X=1.745 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_c_417_n N_A_257_47#_c_452_n 0.0120855f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_412_n N_A_257_47#_c_453_n 0.0175816f $X=1.85 $Y=0.445 $X2=0
+ $Y2=0
cc_238 N_VGND_c_417_n N_A_257_47#_c_453_n 0.011396f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_416_n N_A_257_47#_c_455_n 0.0128458f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_c_417_n N_A_257_47#_c_455_n 0.00875273f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_417_n A_520_47# 0.00169626f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
