* File: sky130_fd_sc_lp__a2bb2oi_0.pex.spice
* Created: Wed Sep  2 09:24:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2OI_0%A1_N 2 5 9 11 12 13 14 19
c28 12 0 1.62788e-19 $X=0.24 $Y=0.925
r29 19 21 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.327 $Y=1.005
+ $X2=0.327 $Y2=0.84
r30 13 14 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.665
r31 12 13 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=0.925
+ $X2=0.27 $Y2=1.295
r32 12 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r33 9 11 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=0.475 $Y=2.455
+ $X2=0.475 $Y2=1.51
r34 5 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.84
r35 2 11 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=0.327 $Y=1.288
+ $X2=0.327 $Y2=1.51
r36 1 19 7.12377 $w=4.45e-07 $l=5.7e-08 $layer=POLY_cond $X=0.327 $Y=1.062
+ $X2=0.327 $Y2=1.005
r37 1 2 28.2451 $w=4.45e-07 $l=2.26e-07 $layer=POLY_cond $X=0.327 $Y=1.062
+ $X2=0.327 $Y2=1.288
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_0%A2_N 3 7 8 9 13 15
c36 3 0 1.62788e-19 $X=0.835 $Y=2.455
r37 13 16 79.7055 $w=6.05e-07 $l=5.05e-07 $layer=POLY_cond $X=1.062 $Y=0.93
+ $X2=1.062 $Y2=1.435
r38 13 15 49.6377 $w=6.05e-07 $l=1.65e-07 $layer=POLY_cond $X=1.062 $Y=0.93
+ $X2=1.062 $Y2=0.765
r39 8 9 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.182 $Y=0.925
+ $X2=1.182 $Y2=1.295
r40 8 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2 $Y=0.93
+ $X2=1.2 $Y2=0.93
r41 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.905 $Y=0.445
+ $X2=0.905 $Y2=0.765
r42 3 16 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=0.835 $Y=2.455
+ $X2=0.835 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_0%A_110_47# 1 2 7 11 13 15 17 20 23 26 33 38
c62 11 0 1.78466e-19 $X=1.9 $Y=0.445
r63 34 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.315 $Y=1.81
+ $X2=1.48 $Y2=1.81
r64 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.315
+ $Y=1.81 $X2=1.315 $Y2=1.81
r65 31 33 6.21492 $w=5.08e-07 $l=2.65e-07 $layer=LI1_cond $X=1.05 $Y=1.9
+ $X2=1.315 $Y2=1.9
r66 29 31 7.57516 $w=5.08e-07 $l=3.23e-07 $layer=LI1_cond $X=0.727 $Y=1.9
+ $X2=1.05 $Y2=1.9
r67 26 28 7.68624 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.692 $Y=0.445
+ $X2=0.692 $Y2=0.61
r68 21 31 3.28461 $w=3.3e-07 $l=2.55e-07 $layer=LI1_cond $X=1.05 $Y=2.155
+ $X2=1.05 $Y2=1.9
r69 21 23 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.05 $Y=2.155
+ $X2=1.05 $Y2=2.29
r70 20 29 6.13047 $w=2.05e-07 $l=2.55e-07 $layer=LI1_cond $X=0.727 $Y=1.645
+ $X2=0.727 $Y2=1.9
r71 20 28 55.9956 $w=2.03e-07 $l=1.035e-06 $layer=LI1_cond $X=0.727 $Y=1.645
+ $X2=0.727 $Y2=0.61
r72 16 17 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.9 $Y=1.74
+ $X2=2.025 $Y2=1.74
r73 13 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.025 $Y=1.815
+ $X2=2.025 $Y2=1.74
r74 13 15 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.025 $Y=1.815
+ $X2=2.025 $Y2=2.255
r75 9 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.9 $Y=1.665 $X2=1.9
+ $Y2=1.74
r76 9 11 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=1.9 $Y=1.665 $X2=1.9
+ $Y2=0.445
r77 7 16 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.825 $Y=1.74 $X2=1.9
+ $Y2=1.74
r78 7 38 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.825 $Y=1.74
+ $X2=1.48 $Y2=1.74
r79 2 23 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=2.135 $X2=1.05 $Y2=2.29
r80 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_0%B2 3 7 11 12 13 14 18
c41 3 0 4.25579e-20 $X=2.33 $Y=0.445
r42 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.38
+ $Y=0.97 $X2=2.38 $Y2=0.97
r43 14 19 7.85304 $w=4.93e-07 $l=3.25e-07 $layer=LI1_cond $X=2.302 $Y=1.295
+ $X2=2.302 $Y2=0.97
r44 13 19 1.08734 $w=4.93e-07 $l=4.5e-08 $layer=LI1_cond $X=2.302 $Y=0.925
+ $X2=2.302 $Y2=0.97
r45 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.38 $Y=1.31
+ $X2=2.38 $Y2=0.97
r46 11 12 43.7316 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.31
+ $X2=2.38 $Y2=1.475
r47 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=0.805
+ $X2=2.38 $Y2=0.97
r48 7 12 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.455 $Y=2.255
+ $X2=2.455 $Y2=1.475
r49 3 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.33 $Y=0.445
+ $X2=2.33 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_0%B1 3 7 11 12 13 14 18
c29 13 0 2.27637e-20 $X=3.12 $Y=0.925
r30 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=0.97 $X2=2.95 $Y2=0.97
r31 14 19 9.13522 $w=4.08e-07 $l=3.25e-07 $layer=LI1_cond $X=3.07 $Y=1.295
+ $X2=3.07 $Y2=0.97
r32 13 19 1.26488 $w=4.08e-07 $l=4.5e-08 $layer=LI1_cond $X=3.07 $Y=0.925
+ $X2=3.07 $Y2=0.97
r33 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.95 $Y=1.31
+ $X2=2.95 $Y2=0.97
r34 11 12 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.31
+ $X2=2.95 $Y2=1.475
r35 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=0.805
+ $X2=2.95 $Y2=0.97
r36 7 12 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.885 $Y=2.255
+ $X2=2.885 $Y2=1.475
r37 3 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.86 $Y=0.445
+ $X2=2.86 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_0%VPWR 1 2 7 9 13 15 17 27 28 34
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.67 $Y2=3.33
r44 25 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 18 31 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r51 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.67 $Y2=3.33
r53 17 23 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=3.33
r57 11 13 41.034 $w=3.28e-07 $l=1.175e-06 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=2.07
r58 7 31 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r59 7 9 33.7002 $w=3.28e-07 $l=9.65e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.28
r60 2 13 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=2.53
+ $Y=1.935 $X2=2.67 $Y2=2.07
r61 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.135 $X2=0.26 $Y2=2.28
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_0%Y 1 2 12 14 15 16 17 18 19 43 45 49
c42 14 0 1.97942e-20 $X=1.595 $Y=0.84
r43 49 51 1.42082 $w=3.63e-07 $l=4.5e-08 $layer=LI1_cond $X=1.752 $Y=2.035
+ $X2=1.752 $Y2=2.08
r44 35 51 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=1.752 $Y=2.097
+ $X2=1.752 $Y2=2.08
r45 28 45 0.439026 $w=3.13e-07 $l=1.2e-08 $layer=LI1_cond $X=1.727 $Y=0.937
+ $X2=1.727 $Y2=0.925
r46 18 19 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.752 $Y=2.405
+ $X2=1.752 $Y2=2.775
r47 17 49 0.378885 $w=3.63e-07 $l=1.2e-08 $layer=LI1_cond $X=1.752 $Y=2.023
+ $X2=1.752 $Y2=2.035
r48 17 47 3.65793 $w=3.63e-07 $l=1.08e-07 $layer=LI1_cond $X=1.752 $Y=2.023
+ $X2=1.752 $Y2=1.915
r49 17 18 9.37741 $w=3.63e-07 $l=2.97e-07 $layer=LI1_cond $X=1.752 $Y=2.108
+ $X2=1.752 $Y2=2.405
r50 17 35 0.347312 $w=3.63e-07 $l=1.1e-08 $layer=LI1_cond $X=1.752 $Y=2.108
+ $X2=1.752 $Y2=2.097
r51 16 47 9.14637 $w=3.13e-07 $l=2.5e-07 $layer=LI1_cond $X=1.727 $Y=1.665
+ $X2=1.727 $Y2=1.915
r52 15 16 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.727 $Y=1.295
+ $X2=1.727 $Y2=1.665
r53 14 45 1.35366 $w=3.13e-07 $l=3.7e-08 $layer=LI1_cond $X=1.727 $Y=0.888
+ $X2=1.727 $Y2=0.925
r54 14 43 6.3772 $w=3.13e-07 $l=1.08e-07 $layer=LI1_cond $X=1.727 $Y=0.888
+ $X2=1.727 $Y2=0.78
r55 14 15 11.7805 $w=3.13e-07 $l=3.22e-07 $layer=LI1_cond $X=1.727 $Y=0.973
+ $X2=1.727 $Y2=1.295
r56 14 28 1.31708 $w=3.13e-07 $l=3.6e-08 $layer=LI1_cond $X=1.727 $Y=0.973
+ $X2=1.727 $Y2=0.937
r57 9 12 10.8364 $w=3.33e-07 $l=3.15e-07 $layer=LI1_cond $X=1.8 $Y=0.442
+ $X2=2.115 $Y2=0.442
r58 7 9 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.8 $Y=0.61 $X2=1.8
+ $Y2=0.442
r59 7 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.8 $Y=0.61 $X2=1.8
+ $Y2=0.78
r60 2 51 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.685
+ $Y=1.935 $X2=1.81 $Y2=2.08
r61 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.115 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_0%A_420_387# 1 2 9 11 12 15
c28 12 0 1.78466e-19 $X=2.335 $Y=1.73
r29 13 15 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=3.14 $Y=1.815
+ $X2=3.14 $Y2=2.08
r30 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.015 $Y=1.73
+ $X2=3.14 $Y2=1.815
r31 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.015 $Y=1.73
+ $X2=2.335 $Y2=1.73
r32 7 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.22 $Y=1.815
+ $X2=2.335 $Y2=1.73
r33 7 9 13.2781 $w=2.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.22 $Y=1.815
+ $X2=2.22 $Y2=2.08
r34 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.96
+ $Y=1.935 $X2=3.1 $Y2=2.08
r35 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.1
+ $Y=1.935 $X2=2.24 $Y2=2.08
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_0%VGND 1 2 3 10 12 14 16 18 20 25 45
r44 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 32 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r47 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 28 31 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r49 26 28 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.68
+ $Y2=0
r50 25 44 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=3.135
+ $Y2=0
r51 25 31 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=2.64
+ $Y2=0
r52 24 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r53 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r54 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 21 34 4.40339 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.192
+ $Y2=0
r56 21 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.72
+ $Y2=0
r57 20 41 9.76614 $w=5.43e-07 $l=4.45e-07 $layer=LI1_cond $X=1.272 $Y=0
+ $X2=1.272 $Y2=0.445
r58 20 26 7.70116 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=1.272 $Y=0 $X2=1.545
+ $Y2=0
r59 20 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r60 20 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.72
+ $Y2=0
r61 18 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r62 18 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r63 18 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 14 44 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.075 $Y=0.085
+ $X2=3.135 $Y2=0
r65 14 16 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.075 $Y=0.085
+ $X2=3.075 $Y2=0.445
r66 10 34 3.03446 $w=2.9e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.192 $Y2=0
r67 10 12 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.445
r68 3 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.935
+ $Y=0.235 $X2=3.075 $Y2=0.445
r69 2 41 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.235 $X2=1.46 $Y2=0.445
r70 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

