* File: sky130_fd_sc_lp__a41o_1.pex.spice
* Created: Wed Sep  2 09:28:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41O_1%A_113_237# 1 2 9 11 13 17 18 19 20 21 22 25
+ 31
r57 33 35 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.64 $Y=1.35 $X2=0.68
+ $Y2=1.35
r58 29 31 27.7273 $w=1.78e-07 $l=4.5e-07 $layer=LI1_cond $X=1.815 $Y=0.87
+ $X2=1.815 $Y2=0.42
r59 25 27 36.3313 $w=2.93e-07 $l=9.3e-07 $layer=LI1_cond $X=1.422 $Y=1.98
+ $X2=1.422 $Y2=2.91
r60 23 25 8.0085 $w=2.93e-07 $l=2.05e-07 $layer=LI1_cond $X=1.422 $Y=1.775
+ $X2=1.422 $Y2=1.98
r61 21 23 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=1.275 $Y=1.69
+ $X2=1.422 $Y2=1.775
r62 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.275 $Y=1.69
+ $X2=0.945 $Y2=1.69
r63 19 29 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.725 $Y=0.955
+ $X2=1.815 $Y2=0.87
r64 19 20 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.725 $Y=0.955
+ $X2=0.945 $Y2=0.955
r65 18 35 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.835 $Y=1.35
+ $X2=0.68 $Y2=1.35
r66 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.835
+ $Y=1.35 $X2=0.835 $Y2=1.35
r67 15 22 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.842 $Y=1.605
+ $X2=0.945 $Y2=1.69
r68 15 17 13.796 $w=2.03e-07 $l=2.55e-07 $layer=LI1_cond $X=0.842 $Y=1.605
+ $X2=0.842 $Y2=1.35
r69 14 20 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.842 $Y=1.04
+ $X2=0.945 $Y2=0.955
r70 14 17 16.7716 $w=2.03e-07 $l=3.1e-07 $layer=LI1_cond $X=0.842 $Y=1.04
+ $X2=0.842 $Y2=1.35
r71 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.68 $Y=1.185
+ $X2=0.68 $Y2=1.35
r72 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.68 $Y=1.185
+ $X2=0.68 $Y2=0.655
r73 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=1.515
+ $X2=0.64 $Y2=1.35
r74 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.64 $Y=1.515 $X2=0.64
+ $Y2=2.465
r75 2 27 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.835 $X2=1.44 $Y2=2.91
r76 2 25 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.835 $X2=1.44 $Y2=1.98
r77 1 31 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.68
+ $Y=0.235 $X2=1.82 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_1%B1 3 6 8 9 13 15
r35 13 16 47.4091 $w=5.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.535 $Y=1.35
+ $X2=1.535 $Y2=1.515
r36 13 15 47.4091 $w=5.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.535 $Y=1.35
+ $X2=1.535 $Y2=1.185
r37 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=1.35 $X2=1.635 $Y2=1.35
r38 8 9 22.2806 $w=2.23e-07 $l=4.35e-07 $layer=LI1_cond $X=1.2 $Y=1.322
+ $X2=1.635 $Y2=1.322
r39 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.655 $Y=2.465
+ $X2=1.655 $Y2=1.515
r40 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.605 $Y=0.655
+ $X2=1.605 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_1%A1 3 5 7 8 9 10 19
r35 17 19 14.4261 $w=3.6e-07 $l=9e-08 $layer=POLY_cond $X=2.225 $Y=1.365
+ $X2=2.315 $Y2=1.365
r36 14 17 22.4405 $w=3.6e-07 $l=1.4e-07 $layer=POLY_cond $X=2.085 $Y=1.365
+ $X2=2.225 $Y2=1.365
r37 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.225
+ $Y=1.35 $X2=2.225 $Y2=1.35
r38 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.21 $Y=0.925
+ $X2=2.21 $Y2=1.295
r39 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.21 $Y=0.555 $X2=2.21
+ $Y2=0.925
r40 5 19 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.315 $Y=1.185
+ $X2=2.315 $Y2=1.365
r41 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.315 $Y=1.185
+ $X2=2.315 $Y2=0.655
r42 1 14 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.085 $Y=1.545
+ $X2=2.085 $Y2=1.365
r43 1 3 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=2.085 $Y=1.545
+ $X2=2.085 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_1%A2 3 6 8 9 10 15 17
r33 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.35
+ $X2=2.765 $Y2=1.515
r34 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.35
+ $X2=2.765 $Y2=1.185
r35 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.35 $X2=2.765 $Y2=1.35
r36 10 16 1.89207 $w=3.33e-07 $l=5.5e-08 $layer=LI1_cond $X=2.682 $Y=1.295
+ $X2=2.682 $Y2=1.35
r37 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.682 $Y=0.925
+ $X2=2.682 $Y2=1.295
r38 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.682 $Y=0.555
+ $X2=2.682 $Y2=0.925
r39 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.855 $Y=2.465
+ $X2=2.855 $Y2=1.515
r40 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.675 $Y=0.655
+ $X2=2.675 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_1%A3 3 6 8 9 10 21 23
r35 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.35
+ $X2=3.305 $Y2=1.515
r36 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.35
+ $X2=3.305 $Y2=1.185
r37 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.305
+ $Y=1.35 $X2=3.305 $Y2=1.35
r38 10 22 0.989238 $w=6.63e-07 $l=5.5e-08 $layer=LI1_cond $X=3.352 $Y=1.295
+ $X2=3.352 $Y2=1.35
r39 9 10 6.65487 $w=6.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.352 $Y=0.925
+ $X2=3.352 $Y2=1.295
r40 8 9 6.65487 $w=6.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.352 $Y=0.555
+ $X2=3.352 $Y2=0.925
r41 6 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.285 $Y=2.465
+ $X2=3.285 $Y2=1.515
r42 3 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.215 $Y=0.655
+ $X2=3.215 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_1%A4 1 3 6 8 13
r23 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.35 $X2=3.95 $Y2=1.35
r24 10 13 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=3.755 $Y=1.35
+ $X2=3.95 $Y2=1.35
r25 8 14 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.08 $Y=1.35 $X2=3.95
+ $Y2=1.35
r26 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=1.515
+ $X2=3.755 $Y2=1.35
r27 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.755 $Y=1.515
+ $X2=3.755 $Y2=2.465
r28 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=1.185
+ $X2=3.755 $Y2=1.35
r29 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.755 $Y=1.185
+ $X2=3.755 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_1%X 1 2 7 8 9 10 11 12 13 22
r13 13 41 3.32929 $w=4.83e-07 $l=1.35e-07 $layer=LI1_cond $X=0.327 $Y=2.775
+ $X2=0.327 $Y2=2.91
r14 12 13 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.327 $Y=2.405
+ $X2=0.327 $Y2=2.775
r15 11 12 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.327 $Y=2.035
+ $X2=0.327 $Y2=2.405
r16 11 33 1.35638 $w=4.83e-07 $l=5.5e-08 $layer=LI1_cond $X=0.327 $Y=2.035
+ $X2=0.327 $Y2=1.98
r17 10 33 7.76834 $w=4.83e-07 $l=3.15e-07 $layer=LI1_cond $X=0.327 $Y=1.665
+ $X2=0.327 $Y2=1.98
r18 9 10 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.327 $Y=1.295
+ $X2=0.327 $Y2=1.665
r19 8 9 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.327 $Y=0.925
+ $X2=0.327 $Y2=1.295
r20 7 8 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.327 $Y=0.555
+ $X2=0.327 $Y2=0.925
r21 7 22 3.32929 $w=4.83e-07 $l=1.35e-07 $layer=LI1_cond $X=0.327 $Y=0.555
+ $X2=0.327 $Y2=0.42
r22 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.835 $X2=0.425 $Y2=2.91
r23 2 33 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.835 $X2=0.425 $Y2=1.98
r24 1 22 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.34
+ $Y=0.235 $X2=0.465 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_1%VPWR 1 2 3 12 18 24 29 30 31 37 41 48 49 52
+ 57
r56 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 49 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 46 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.52 $Y2=3.33
r61 46 48 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r63 45 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r65 42 52 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.47 $Y2=3.33
r66 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 41 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.52 $Y2=3.33
r68 41 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.12 $Y2=3.33
r69 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r70 37 52 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=2.47 $Y2=3.33
r71 37 39 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.135 $Y=3.33 $X2=1.2
+ $Y2=3.33
r72 35 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 31 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r75 31 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r76 31 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 29 34 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.75 $Y=3.33 $X2=0.72
+ $Y2=3.33
r78 29 30 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.75 $Y=3.33
+ $X2=0.885 $Y2=3.33
r79 28 39 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.02 $Y=3.33 $X2=1.2
+ $Y2=3.33
r80 28 30 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.02 $Y=3.33
+ $X2=0.885 $Y2=3.33
r81 24 27 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=3.52 $Y=2.11
+ $X2=3.52 $Y2=2.95
r82 22 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=3.33
r83 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=2.95
r84 18 21 14.9956 $w=6.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.47 $Y=2.11
+ $X2=2.47 $Y2=2.95
r85 16 52 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=3.245
+ $X2=2.47 $Y2=3.33
r86 16 21 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.47 $Y=3.245
+ $X2=2.47 $Y2=2.95
r87 12 15 35.8538 $w=2.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.885 $Y=2.11
+ $X2=0.885 $Y2=2.95
r88 10 30 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=3.245
+ $X2=0.885 $Y2=3.33
r89 10 15 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.885 $Y=3.245
+ $X2=0.885 $Y2=2.95
r90 3 27 400 $w=1.7e-07 $l=1.19232e-06 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.835 $X2=3.52 $Y2=2.95
r91 3 24 400 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.835 $X2=3.52 $Y2=2.11
r92 2 21 200 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=3 $X=2.16
+ $Y=1.835 $X2=2.3 $Y2=2.95
r93 2 18 200 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=3 $X=2.16
+ $Y=1.835 $X2=2.3 $Y2=2.11
r94 1 15 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=1.835 $X2=0.855 $Y2=2.95
r95 1 12 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=1.835 $X2=0.855 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_1%A_346_367# 1 2 3 12 16 17 20 24 28 32
r37 28 30 38.2776 $w=2.78e-07 $l=9.3e-07 $layer=LI1_cond $X=3.995 $Y=1.98
+ $X2=3.995 $Y2=2.91
r38 26 28 5.14483 $w=2.78e-07 $l=1.25e-07 $layer=LI1_cond $X=3.995 $Y=1.855
+ $X2=3.995 $Y2=1.98
r39 25 32 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.185 $Y=1.77
+ $X2=3.08 $Y2=1.77
r40 24 26 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.855 $Y=1.77
+ $X2=3.995 $Y2=1.855
r41 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.855 $Y=1.77
+ $X2=3.185 $Y2=1.77
r42 20 22 49.1169 $w=2.08e-07 $l=9.3e-07 $layer=LI1_cond $X=3.08 $Y=1.98
+ $X2=3.08 $Y2=2.91
r43 18 32 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=1.855
+ $X2=3.08 $Y2=1.77
r44 18 20 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=3.08 $Y=1.855
+ $X2=3.08 $Y2=1.98
r45 16 32 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.975 $Y=1.77
+ $X2=3.08 $Y2=1.77
r46 16 17 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.975 $Y=1.77
+ $X2=1.965 $Y2=1.77
r47 12 14 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=1.852 $Y=1.98
+ $X2=1.852 $Y2=2.91
r48 10 17 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.852 $Y=1.855
+ $X2=1.965 $Y2=1.77
r49 10 12 6.40246 $w=2.23e-07 $l=1.25e-07 $layer=LI1_cond $X=1.852 $Y=1.855
+ $X2=1.852 $Y2=1.98
r50 3 30 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.835 $X2=3.97 $Y2=2.91
r51 3 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.835 $X2=3.97 $Y2=1.98
r52 2 22 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.835 $X2=3.07 $Y2=2.91
r53 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.835 $X2=3.07 $Y2=1.98
r54 1 14 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.73
+ $Y=1.835 $X2=1.87 $Y2=2.91
r55 1 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.73
+ $Y=1.835 $X2=1.87 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_1%VGND 1 2 7 9 11 18 29 32 35
r45 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r46 31 32 11.3415 $w=7.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0.307
+ $X2=1.555 $Y2=0.307
r47 27 31 2.89497 $w=7.83e-07 $l=1.9e-07 $layer=LI1_cond $X=1.2 $Y=0.307
+ $X2=1.39 $Y2=0.307
r48 27 29 15.6839 $w=7.83e-07 $l=4.5e-07 $layer=LI1_cond $X=1.2 $Y=0.307
+ $X2=0.75 $Y2=0.307
r49 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r51 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r52 22 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r53 21 24 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r54 21 32 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.555
+ $Y2=0
r55 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 18 34 4.1749 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=4.087
+ $Y2=0
r57 18 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=3.6
+ $Y2=0
r58 16 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r59 15 29 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.75
+ $Y2=0
r60 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 11 25 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r62 11 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r63 7 34 3.18516 $w=2.8e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.995 $Y=0.085
+ $X2=4.087 $Y2=0
r64 7 9 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.995 $Y=0.085
+ $X2=3.995 $Y2=0.38
r65 2 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.83
+ $Y=0.235 $X2=3.97 $Y2=0.38
r66 1 31 91 $w=1.7e-07 $l=7.86845e-07 $layer=licon1_NDIFF $count=2 $X=0.755
+ $Y=0.235 $X2=1.39 $Y2=0.575
.ends

