* File: sky130_fd_sc_lp__a41o_0.spice
* Created: Fri Aug 28 10:02:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41o_0.pex.spice"
.subckt sky130_fd_sc_lp__a41o_0  VNB VPB B1 A1 A2 A3 A4 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_80_309#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_80_309#_M1006_d N_B1_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0588 PD=1.04 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1011 A_385_47# N_A1_M1011_g N_A_80_309#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.1302 PD=0.73 PS=1.04 NRD=28.56 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1007 A_477_47# N_A2_M1007_g A_385_47# VNB NSHORT L=0.15 W=0.42 AD=0.0609
+ AS=0.0651 PD=0.71 PS=0.73 NRD=25.704 NRS=28.56 M=1 R=2.8 SA=75001.8 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1003 A_565_47# N_A3_M1003_g A_477_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0609 PD=0.63 PS=0.71 NRD=14.28 NRS=25.704 M=1 R=2.8 SA=75002.3 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A4_M1004_g A_565_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_80_309#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_321_473#_M1008_d N_B1_M1008_g N_A_80_309#_M1008_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_321_473#_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1000 N_A_321_473#_M1000_d N_A2_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_A3_M1009_g N_A_321_473#_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0976 AS=0.0896 PD=0.945 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1010 N_A_321_473#_M1010_d N_A4_M1010_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0976 PD=1.81 PS=0.945 NRD=0 NRS=7.683 M=1 R=4.26667
+ SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a41o_0.pxi.spice"
*
.ends
*
*
