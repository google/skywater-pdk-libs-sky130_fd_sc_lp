* File: sky130_fd_sc_lp__or4bb_m.pex.spice
* Created: Fri Aug 28 11:27:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4BB_M%C_N 3 7 9 10 11 12 13 17
r33 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.54
+ $Y=0.94 $X2=0.54 $Y2=0.94
r34 13 18 11.6891 $w=3.48e-07 $l=3.55e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=0.94
r35 12 18 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=0.63 $Y=0.925
+ $X2=0.63 $Y2=0.94
r36 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.54 $Y=1.28
+ $X2=0.54 $Y2=0.94
r37 10 11 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.28
+ $X2=0.54 $Y2=1.445
r38 9 17 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=0.775
+ $X2=0.54 $Y2=0.94
r39 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.59 $Y=0.455 $X2=0.59
+ $Y2=0.775
r40 3 11 725.564 $w=1.5e-07 $l=1.415e-06 $layer=POLY_cond $X=0.475 $Y=2.86
+ $X2=0.475 $Y2=1.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_M%D_N 3 7 9 12 13
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=2.17
+ $X2=0.995 $Y2=2.335
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=2.17
+ $X2=0.995 $Y2=2.005
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=2.17 $X2=0.995 $Y2=2.17
r39 9 13 6.32541 $w=5.18e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=2.265
+ $X2=0.995 $Y2=2.265
r40 7 14 794.787 $w=1.5e-07 $l=1.55e-06 $layer=POLY_cond $X=1.02 $Y=0.455
+ $X2=1.02 $Y2=2.005
r41 3 15 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=0.905 $Y=2.86
+ $X2=0.905 $Y2=2.335
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_M%A_196_530# 1 2 8 11 13 15 16 18 22 25 26 31
+ 32 36 38 39 42 43 47
c71 32 0 1.31411e-19 $X=1.57 $Y=2.94
r72 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.62
+ $Y=0.94 $X2=1.62 $Y2=0.94
r73 40 42 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.62 $Y=0.905
+ $X2=1.62 $Y2=0.94
r74 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.535 $Y=0.82
+ $X2=1.62 $Y2=0.905
r75 38 39 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.535 $Y=0.82
+ $X2=1.34 $Y2=0.82
r76 34 39 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.235 $Y=0.735
+ $X2=1.34 $Y2=0.82
r77 34 36 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.235 $Y=0.735
+ $X2=1.235 $Y2=0.52
r78 32 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=2.94
+ $X2=1.57 $Y2=2.775
r79 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=2.94 $X2=1.57 $Y2=2.94
r80 28 31 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=2.86
+ $X2=1.57 $Y2=2.86
r81 24 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.62 $Y=1.28
+ $X2=1.62 $Y2=0.94
r82 24 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.28
+ $X2=1.62 $Y2=1.445
r83 20 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.62 $Y=0.925
+ $X2=1.62 $Y2=0.94
r84 20 22 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.62 $Y=0.85
+ $X2=1.97 $Y2=0.85
r85 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.02 $Y=2.085
+ $X2=2.02 $Y2=2.405
r86 13 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.97 $Y=0.775
+ $X2=1.97 $Y2=0.85
r87 13 15 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.97 $Y=0.775
+ $X2=1.97 $Y2=0.445
r88 12 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.605 $Y=2.01
+ $X2=1.53 $Y2=2.01
r89 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.945 $Y=2.01
+ $X2=2.02 $Y2=2.085
r90 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.945 $Y=2.01
+ $X2=1.605 $Y2=2.01
r91 9 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.53 $Y=2.085
+ $X2=1.53 $Y2=2.01
r92 9 47 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.53 $Y=2.085
+ $X2=1.53 $Y2=2.775
r93 8 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.53 $Y=1.935
+ $X2=1.53 $Y2=2.01
r94 8 25 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.53 $Y=1.935
+ $X2=1.53 $Y2=1.445
r95 2 28 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.65 $X2=1.12 $Y2=2.86
r96 1 36 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.245 $X2=1.235 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_M%A_27_530# 1 2 7 9 13 16 19 21 26 28 30
c74 30 0 1.00136e-19 $X=2.29 $Y=1.53
c75 7 0 1.80476e-19 $X=2.38 $Y=1.695
r76 30 33 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.29 $Y=1.53
+ $X2=2.29 $Y2=1.71
r77 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.53 $X2=2.29 $Y2=1.53
r78 23 26 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.19 $Y=0.43
+ $X2=0.375 $Y2=0.43
r79 22 28 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.365 $Y=1.71
+ $X2=0.235 $Y2=1.71
r80 21 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=1.71
+ $X2=2.29 $Y2=1.71
r81 21 22 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.205 $Y=1.71
+ $X2=0.365 $Y2=1.71
r82 17 28 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=1.795
+ $X2=0.235 $Y2=1.71
r83 17 19 44.3247 $w=2.58e-07 $l=1e-06 $layer=LI1_cond $X=0.235 $Y=1.795
+ $X2=0.235 $Y2=2.795
r84 16 28 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.19 $Y=1.625
+ $X2=0.235 $Y2=1.71
r85 15 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.19 $Y=0.595
+ $X2=0.19 $Y2=0.43
r86 15 16 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.19 $Y=0.595
+ $X2=0.19 $Y2=1.625
r87 11 31 38.6704 $w=3.39e-07 $l=2.09105e-07 $layer=POLY_cond $X=2.4 $Y=1.365
+ $X2=2.3 $Y2=1.53
r88 11 13 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=2.4 $Y=1.365 $X2=2.4
+ $Y2=0.445
r89 7 31 38.6704 $w=3.39e-07 $l=2.0106e-07 $layer=POLY_cond $X=2.38 $Y=1.695
+ $X2=2.3 $Y2=1.53
r90 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.38 $Y=1.695 $X2=2.38
+ $Y2=2.405
r91 2 19 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.65 $X2=0.26 $Y2=2.795
r92 1 26 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.25
+ $Y=0.245 $X2=0.375 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_M%B 3 7 11 12 13 16 17
c45 11 0 1.00136e-19 $X=2.85 $Y=1.4
r46 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.85
+ $Y=1.06 $X2=2.85 $Y2=1.06
r47 13 17 4.92503 $w=5.08e-07 $l=2.1e-07 $layer=LI1_cond $X=2.64 $Y=1.23
+ $X2=2.85 $Y2=1.23
r48 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.85 $Y=1.4 $X2=2.85
+ $Y2=1.06
r49 11 12 40.0117 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.4
+ $X2=2.85 $Y2=1.565
r50 10 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=0.895
+ $X2=2.85 $Y2=1.06
r51 7 10 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.91 $Y=0.445
+ $X2=2.91 $Y2=0.895
r52 3 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.89 $Y=2.635
+ $X2=2.89 $Y2=1.565
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_M%A 3 7 9 10 15 16
c49 15 0 1.16165e-19 $X=3.34 $Y=2.1
c50 7 0 1.04876e-19 $X=3.34 $Y=0.445
c51 3 0 1.51175e-19 $X=3.25 $Y=2.635
r52 18 24 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.12 $Y=2.32
+ $X2=3.12 $Y2=2.167
r53 16 24 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=3.34 $Y=2.167
+ $X2=3.12 $Y2=2.167
r54 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.34 $Y=2.1
+ $X2=3.34 $Y2=2.265
r55 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.34
+ $Y=2.1 $X2=3.34 $Y2=2.1
r56 9 24 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.12 $Y=2.32 $X2=3.12
+ $Y2=2.167
r57 9 10 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=2.405 $X2=3.12
+ $Y2=2.775
r58 9 18 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=2.405
+ $X2=3.12 $Y2=2.32
r59 5 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.34 $Y=1.935
+ $X2=3.34 $Y2=2.1
r60 5 7 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=3.34 $Y=1.935
+ $X2=3.34 $Y2=0.445
r61 3 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.25 $Y=2.635
+ $X2=3.25 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_M%A_336_439# 1 2 3 12 16 20 21 22 26 29 30 31
+ 33 34 38 39 42 47 51
c107 33 0 9.03474e-20 $X=3.28 $Y=1.665
c108 26 0 2.85353e-19 $X=3.02 $Y=0.71
c109 22 0 3.98751e-19 $X=2.685 $Y=2.34
r110 42 44 9.50649 $w=2.08e-07 $l=1.8e-07 $layer=LI1_cond $X=2.185 $Y=0.53
+ $X2=2.185 $Y2=0.71
r111 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.79
+ $Y=1.19 $X2=3.79 $Y2=1.19
r112 36 38 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.79 $Y=1.665
+ $X2=3.79 $Y2=1.19
r113 35 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=1.75
+ $X2=3.28 $Y2=1.75
r114 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.705 $Y=1.75
+ $X2=3.79 $Y2=1.665
r115 34 35 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.705 $Y=1.75
+ $X2=3.365 $Y2=1.75
r116 33 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=1.665
+ $X2=3.28 $Y2=1.75
r117 33 50 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.28 $Y=1.665
+ $X2=3.28 $Y2=0.795
r118 30 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=1.75
+ $X2=3.28 $Y2=1.75
r119 30 31 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.195 $Y=1.75
+ $X2=2.855 $Y2=1.75
r120 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=1.835
+ $X2=2.855 $Y2=1.75
r121 28 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.77 $Y=1.835
+ $X2=2.77 $Y2=2.175
r122 27 44 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.29 $Y=0.71
+ $X2=2.185 $Y2=0.71
r123 26 50 5.80707 $w=3.43e-07 $l=8.5e-08 $layer=LI1_cond $X=3.192 $Y=0.71
+ $X2=3.192 $Y2=0.795
r124 26 47 6.68083 $w=3.43e-07 $l=2e-07 $layer=LI1_cond $X=3.192 $Y=0.71
+ $X2=3.192 $Y2=0.51
r125 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.02 $Y=0.71
+ $X2=2.29 $Y2=0.71
r126 22 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.685 $Y=2.34
+ $X2=2.77 $Y2=2.175
r127 22 24 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=2.685 $Y=2.34
+ $X2=1.805 $Y2=2.34
r128 20 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.79 $Y=1.53
+ $X2=3.79 $Y2=1.19
r129 20 21 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=1.53
+ $X2=3.79 $Y2=1.695
r130 19 39 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=1.025
+ $X2=3.79 $Y2=1.19
r131 16 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.845 $Y=0.445
+ $X2=3.845 $Y2=1.025
r132 12 21 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.825 $Y=2.635
+ $X2=3.825 $Y2=1.695
r133 3 24 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=2.195 $X2=1.805 $Y2=2.34
r134 2 47 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.985
+ $Y=0.235 $X2=3.125 $Y2=0.51
r135 1 42 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.235 $X2=2.185 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_M%VPWR 1 2 9 13 15 17 22 29 30 33 36
r44 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 33 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=3.55 $Y2=3.33
r49 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r51 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 23 33 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.775 $Y=3.33
+ $X2=0.68 $Y2=3.33
r53 23 25 152.989 $w=1.68e-07 $l=2.345e-06 $layer=LI1_cond $X=0.775 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.55 $Y2=3.33
r55 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 17 33 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.68 $Y2=3.33
r59 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 15 34 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.55 $Y2=3.33
r63 11 13 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.55 $Y2=2.7
r64 7 33 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=3.33
r65 7 9 18.6794 $w=1.88e-07 $l=3.2e-07 $layer=LI1_cond $X=0.68 $Y=3.245 $X2=0.68
+ $Y2=2.925
r66 2 13 600 $w=1.7e-07 $l=3.7081e-07 $layer=licon1_PDIFF $count=1 $X=3.325
+ $Y=2.425 $X2=3.55 $Y2=2.7
r67 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.65 $X2=0.69 $Y2=2.925
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_M%X 1 2 9 12 13 30
r18 18 30 2.38436 $w=2.88e-07 $l=6e-08 $layer=LI1_cond $X=4.08 $Y=2.465 $X2=4.08
+ $Y2=2.405
r19 13 21 8.14658 $w=2.88e-07 $l=2.05e-07 $layer=LI1_cond $X=4.08 $Y=2.775
+ $X2=4.08 $Y2=2.57
r20 12 30 0.516612 $w=2.88e-07 $l=1.3e-08 $layer=LI1_cond $X=4.08 $Y=2.392
+ $X2=4.08 $Y2=2.405
r21 12 21 3.69577 $w=2.88e-07 $l=9.3e-08 $layer=LI1_cond $X=4.08 $Y=2.477
+ $X2=4.08 $Y2=2.57
r22 12 18 0.476873 $w=2.88e-07 $l=1.2e-08 $layer=LI1_cond $X=4.08 $Y=2.477
+ $X2=4.08 $Y2=2.465
r23 11 12 68.92 $w=2.78e-07 $l=1.645e-06 $layer=LI1_cond $X=4.14 $Y=0.675
+ $X2=4.14 $Y2=2.32
r24 9 11 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0.51
+ $X2=4.09 $Y2=0.675
r25 2 21 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=2.425 $X2=4.04 $Y2=2.57
r26 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.235 $X2=4.06 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_M%VGND 1 2 3 4 17 19 23 27 29 33 35 37 44 45
+ 48 51 54 57
r70 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r71 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r72 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r73 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 49 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r75 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r76 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r77 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r78 42 57 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.64
+ $Y2=0
r79 42 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=4.08
+ $Y2=0
r80 38 51 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.755
+ $Y2=0
r81 38 40 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=2.16
+ $Y2=0
r82 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.635
+ $Y2=0
r83 37 40 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.16
+ $Y2=0
r84 35 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r85 35 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r86 35 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r87 31 57 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0
r88 31 33 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0.38
r89 30 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.635
+ $Y2=0
r90 29 57 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.545 $Y=0 $X2=3.64
+ $Y2=0
r91 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.545 $Y=0 $X2=2.8
+ $Y2=0
r92 25 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0
r93 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0.36
r94 21 51 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0.085
+ $X2=1.755 $Y2=0
r95 21 23 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.755 $Y=0.085
+ $X2=1.755 $Y2=0.38
r96 20 48 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.805
+ $Y2=0
r97 19 51 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.755
+ $Y2=0
r98 19 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.65 $Y=0 $X2=0.91
+ $Y2=0
r99 15 48 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0
r100 15 17 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0.39
r101 4 33 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.63 $Y2=0.38
r102 3 27 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.635 $Y2=0.36
r103 2 23 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.63
+ $Y=0.235 $X2=1.755 $Y2=0.38
r104 1 17 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.665
+ $Y=0.245 $X2=0.805 $Y2=0.39
.ends

