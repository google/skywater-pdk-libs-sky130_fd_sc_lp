* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or3_0 A B C VGND VNB VPB VPWR X
X0 a_29_55# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND B a_29_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_29_55# C a_191_481# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_191_481# B a_263_481# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_263_481# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_29_55# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_29_55# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_29_55# X VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
