* File: sky130_fd_sc_lp__dfbbp_1.pex.spice
* Created: Fri Aug 28 10:21:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFBBP_1%CLK 2 5 7 9 12 14 17 19 20 21 26 27
c37 5 0 1.65835e-19 $X=0.495 $Y=0.495
r38 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=1.07 $X2=0.29 $Y2=1.07
r39 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=2.035
r40 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r41 19 27 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.07
r42 15 17 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.38 $Y=2.255
+ $X2=0.645 $Y2=2.255
r43 13 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.29 $Y=1.41
+ $X2=0.29 $Y2=1.07
r44 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.29 $Y=1.41
+ $X2=0.29 $Y2=1.575
r45 12 26 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.29 $Y=1.03 $X2=0.29
+ $Y2=1.07
r46 11 12 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.347 $Y=0.88
+ $X2=0.347 $Y2=1.03
r47 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.645 $Y=2.33
+ $X2=0.645 $Y2=2.255
r48 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.645 $Y=2.33
+ $X2=0.645 $Y2=2.725
r49 5 11 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.495 $Y=0.495
+ $X2=0.495 $Y2=0.88
r50 2 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.38 $Y=2.18 $X2=0.38
+ $Y2=2.255
r51 2 14 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=0.38 $Y=2.18
+ $X2=0.38 $Y2=1.575
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%D 1 3 5 7 8 10 11 12 13 17 24
c62 1 0 1.35289e-20 $X=2.505 $Y=0.84
r63 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=1.89 $X2=2.115 $Y2=1.89
r64 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=0.93 $X2=1.935 $Y2=0.93
r65 17 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.935 $Y=0.84
+ $X2=1.935 $Y2=0.93
r66 13 25 5.27682 $w=5.08e-07 $l=2.25e-07 $layer=LI1_cond $X=2.025 $Y=1.665
+ $X2=2.025 $Y2=1.89
r67 12 13 8.67743 $w=5.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.025 $Y=1.295
+ $X2=2.025 $Y2=1.665
r68 12 21 8.56017 $w=5.08e-07 $l=3.65e-07 $layer=LI1_cond $X=2.025 $Y=1.295
+ $X2=2.025 $Y2=0.93
r69 11 21 0.117263 $w=5.08e-07 $l=5e-09 $layer=LI1_cond $X=2.025 $Y=0.925
+ $X2=2.025 $Y2=0.93
r70 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.76 $Y=2.24 $X2=2.76
+ $Y2=2.525
r71 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.58 $Y=0.765 $X2=2.58
+ $Y2=0.445
r72 4 24 50.0189 $w=2.65e-07 $l=3.47851e-07 $layer=POLY_cond $X=2.28 $Y=2.165
+ $X2=2.115 $Y2=1.89
r73 3 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.685 $Y=2.165
+ $X2=2.76 $Y2=2.24
r74 3 4 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.685 $Y=2.165
+ $X2=2.28 $Y2=2.165
r75 2 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.1 $Y=0.84
+ $X2=1.935 $Y2=0.84
r76 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.505 $Y=0.84
+ $X2=2.58 $Y2=0.765
r77 1 2 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.505 $Y=0.84 $X2=2.1
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_225_47# 1 2 9 13 17 21 23 25 28 31 33 36
+ 38 41 47 52 53 56 57 60 63 69 70
c197 56 0 3.00867e-20 $X=6.815 $Y=1.295
c198 53 0 1.69381e-19 $X=7.11 $Y=2.235
c199 47 0 1.35289e-20 $X=2.835 $Y=1.715
c200 28 0 1.65835e-19 $X=1.42 $Y=2.235
c201 23 0 5.88079e-20 $X=3.115 $Y=1.715
r202 69 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=1.275
+ $X2=6.97 $Y2=1.11
r203 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.97
+ $Y=1.275 $X2=6.97 $Y2=1.275
r204 63 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.295
+ $X2=6.96 $Y2=1.295
r205 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.295
r206 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.295
+ $X2=2.64 $Y2=1.295
r207 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=1.295
+ $X2=6.96 $Y2=1.295
r208 56 57 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=6.815 $Y=1.295
+ $X2=2.785 $Y2=1.295
r209 54 70 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=6.97 $Y=2.07
+ $X2=6.97 $Y2=1.275
r210 53 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.11 $Y=2.235
+ $X2=7.11 $Y2=2.4
r211 52 54 5.07461 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.02 $Y=2.235
+ $X2=7.02 $Y2=2.07
r212 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.11
+ $Y=2.235 $X2=7.11 $Y2=2.235
r213 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.835
+ $Y=1.715 $X2=2.835 $Y2=1.715
r214 45 60 10.3525 $w=2.93e-07 $l=2.65e-07 $layer=LI1_cond $X=2.607 $Y=1.56
+ $X2=2.607 $Y2=1.295
r215 44 47 8.21116 $w=3.18e-07 $l=2.28e-07 $layer=LI1_cond $X=2.607 $Y=1.72
+ $X2=2.835 $Y2=1.72
r216 44 45 1.22678 $w=2.95e-07 $l=1.6e-07 $layer=LI1_cond $X=2.607 $Y=1.72
+ $X2=2.607 $Y2=1.56
r217 42 44 2.23286 $w=3.18e-07 $l=6.2e-08 $layer=LI1_cond $X=2.545 $Y=1.72
+ $X2=2.607 $Y2=1.72
r218 38 40 6.28597 $w=4.78e-07 $l=2.05e-07 $layer=LI1_cond $X=1.345 $Y=0.47
+ $X2=1.345 $Y2=0.675
r219 35 42 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.545 $Y=1.88
+ $X2=2.545 $Y2=1.72
r220 35 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.545 $Y=1.88
+ $X2=2.545 $Y2=2.235
r221 34 41 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=2.32
+ $X2=1.42 $Y2=2.32
r222 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=2.32
+ $X2=2.545 $Y2=2.235
r223 33 34 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.46 $Y=2.32
+ $X2=1.585 $Y2=2.32
r224 29 41 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=2.405
+ $X2=1.42 $Y2=2.32
r225 29 31 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.42 $Y=2.405
+ $X2=1.42 $Y2=2.46
r226 28 41 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=2.235
+ $X2=1.42 $Y2=2.32
r227 28 40 54.4791 $w=3.28e-07 $l=1.56e-06 $layer=LI1_cond $X=1.42 $Y=2.235
+ $X2=1.42 $Y2=0.675
r228 24 25 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.19 $Y=1.715
+ $X2=3.52 $Y2=1.715
r229 23 48 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=3.115 $Y=1.715
+ $X2=2.835 $Y2=1.715
r230 23 24 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.115 $Y=1.715
+ $X2=3.19 $Y2=1.715
r231 21 75 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.02 $Y=2.77
+ $X2=7.02 $Y2=2.4
r232 17 71 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.91 $Y=0.59
+ $X2=6.91 $Y2=1.11
r233 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.55
+ $X2=3.52 $Y2=1.715
r234 11 13 566.606 $w=1.5e-07 $l=1.105e-06 $layer=POLY_cond $X=3.52 $Y=1.55
+ $X2=3.52 $Y2=0.445
r235 7 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.88
+ $X2=3.19 $Y2=1.715
r236 7 9 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.19 $Y=1.88
+ $X2=3.19 $Y2=2.525
r237 2 31 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.275
+ $Y=2.315 $X2=1.42 $Y2=2.46
r238 1 38 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.27 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_767_21# 1 2 9 13 17 19 20 23 27 28 30 31
+ 32 33 34 38 41 42 46 47 51 55
c159 51 0 1.68735e-19 $X=4.98 $Y=2.415
c160 42 0 1.69381e-19 $X=6.225 $Y=2.045
c161 28 0 3.00867e-20 $X=4 $Y=1.57
c162 27 0 1.19365e-19 $X=4 $Y=1.57
r163 51 53 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=4.98 $Y=2.415
+ $X2=4.98 $Y2=2.59
r164 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.39
+ $Y=1.275 $X2=6.39 $Y2=1.275
r165 44 46 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=6.39 $Y=1.96
+ $X2=6.39 $Y2=1.275
r166 43 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=2.045
+ $X2=5.465 $Y2=2.045
r167 42 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.225 $Y=2.045
+ $X2=6.39 $Y2=1.96
r168 42 43 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.225 $Y=2.045
+ $X2=5.55 $Y2=2.045
r169 41 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=1.96
+ $X2=5.465 $Y2=2.045
r170 40 41 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=5.465 $Y=0.875
+ $X2=5.465 $Y2=1.96
r171 39 50 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.105 $Y=2.045
+ $X2=4.98 $Y2=2.045
r172 38 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.38 $Y=2.045
+ $X2=5.465 $Y2=2.045
r173 38 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.38 $Y=2.045
+ $X2=5.105 $Y2=2.045
r174 34 40 6.78935 $w=2.28e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.38 $Y=0.745
+ $X2=5.465 $Y2=0.875
r175 34 36 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=5.38 $Y=0.745
+ $X2=5.235 $Y2=0.745
r176 33 51 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.33
+ $X2=4.98 $Y2=2.415
r177 32 50 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.13
+ $X2=4.98 $Y2=2.045
r178 32 33 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=4.98 $Y=2.13 $X2=4.98
+ $Y2=2.33
r179 30 51 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=2.415
+ $X2=4.98 $Y2=2.415
r180 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.855 $Y=2.415
+ $X2=4.165 $Y2=2.415
r181 28 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4 $Y=1.57 $X2=4
+ $Y2=1.735
r182 28 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4 $Y=1.57 $X2=4
+ $Y2=1.405
r183 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4 $Y=1.57
+ $X2=4 $Y2=1.57
r184 25 31 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=4.022 $Y=2.33
+ $X2=4.165 $Y2=2.415
r185 25 27 30.7318 $w=2.83e-07 $l=7.6e-07 $layer=LI1_cond $X=4.022 $Y=2.33
+ $X2=4.022 $Y2=1.57
r186 21 47 38.7595 $w=2.78e-07 $l=2.13014e-07 $layer=POLY_cond $X=6.52 $Y=1.11
+ $X2=6.41 $Y2=1.275
r187 21 23 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.52 $Y=1.11
+ $X2=6.52 $Y2=0.59
r188 19 47 56.3489 $w=2.78e-07 $l=4.07124e-07 $layer=POLY_cond $X=6.225 $Y=1.6
+ $X2=6.41 $Y2=1.275
r189 19 20 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.225 $Y=1.6
+ $X2=6.06 $Y2=1.6
r190 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.985 $Y=1.675
+ $X2=6.06 $Y2=1.6
r191 15 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.985 $Y=1.675
+ $X2=5.985 $Y2=2.315
r192 13 58 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.09 $Y=2.525
+ $X2=4.09 $Y2=1.735
r193 9 57 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=3.91 $Y=0.445
+ $X2=3.91 $Y2=1.405
r194 2 53 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=4.8
+ $Y=1.895 $X2=4.94 $Y2=2.59
r195 2 50 600 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_PDIFF $count=1 $X=4.8
+ $Y=1.895 $X2=4.94 $Y2=2.125
r196 1 36 182 $w=1.7e-07 $l=5.79655e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.235 $X2=5.235 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%SET_B 3 5 7 10 14 16 18 19 22 25 30 32 33
c119 30 0 3.30925e-20 $X=4.54 $Y=1.57
c120 25 0 4.06414e-20 $X=8.4 $Y=2.035
c121 19 0 1.40216e-19 $X=4.705 $Y=2.035
c122 5 0 1.68735e-19 $X=4.725 $Y=1.775
r123 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.43 $Y=1.825
+ $X2=8.43 $Y2=1.99
r124 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.43 $Y=1.825
+ $X2=8.43 $Y2=1.66
r125 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.43
+ $Y=1.825 $X2=8.43 $Y2=1.825
r126 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.54
+ $Y=1.57 $X2=4.54 $Y2=1.57
r127 26 33 8.20383 $w=2.93e-07 $l=2.1e-07 $layer=LI1_cond $X=8.412 $Y=2.035
+ $X2=8.412 $Y2=1.825
r128 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r129 22 47 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=4.525 $Y=2.035
+ $X2=4.525 $Y2=1.78
r130 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=2.035
+ $X2=4.56 $Y2=2.035
r131 19 21 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=2.035
+ $X2=4.56 $Y2=2.035
r132 18 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=8.4 $Y2=2.035
r133 18 19 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=4.705 $Y2=2.035
r134 16 47 4.13427 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.54 $Y=1.665
+ $X2=4.54 $Y2=1.78
r135 16 30 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.54 $Y=1.665
+ $X2=4.54 $Y2=1.57
r136 14 35 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.52 $Y=2.57
+ $X2=8.52 $Y2=1.99
r137 10 34 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=8.45 $Y=0.59
+ $X2=8.45 $Y2=1.66
r138 5 29 44.2644 $w=3.68e-07 $l=2.6517e-07 $layer=POLY_cond $X=4.725 $Y=1.775
+ $X2=4.587 $Y2=1.57
r139 5 7 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=4.725 $Y=1.775
+ $X2=4.725 $Y2=2.315
r140 1 29 39.0253 $w=3.68e-07 $l=1.99825e-07 $layer=POLY_cond $X=4.51 $Y=1.405
+ $X2=4.587 $Y2=1.57
r141 1 3 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=4.51 $Y=1.405
+ $X2=4.51 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_617_47# 1 2 9 11 13 16 18 19 22 29
c89 19 0 9.56299e-20 $X=4.915 $Y=1.14
c90 13 0 1.40216e-19 $X=5.155 $Y=2.315
r91 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.08
+ $Y=1.22 $X2=5.08 $Y2=1.22
r92 20 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=1.14 $X2=3.615
+ $Y2=1.14
r93 19 33 3.23493 $w=2.83e-07 $l=8e-08 $layer=LI1_cond $X=5.057 $Y=1.14
+ $X2=5.057 $Y2=1.22
r94 19 20 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=4.915 $Y=1.14
+ $X2=3.7 $Y2=1.14
r95 18 25 4.34254 $w=3.43e-07 $l=1.3e-07 $layer=LI1_cond $X=3.615 $Y=2.582
+ $X2=3.485 $Y2=2.582
r96 17 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=1.225
+ $X2=3.615 $Y2=1.14
r97 17 18 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=3.615 $Y=1.225
+ $X2=3.615 $Y2=2.41
r98 16 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=1.055
+ $X2=3.615 $Y2=1.14
r99 15 22 12.777 $w=2.96e-07 $l=3.9488e-07 $layer=LI1_cond $X=3.615 $Y=0.65
+ $X2=3.305 $Y2=0.457
r100 15 16 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.615 $Y=0.65
+ $X2=3.615 $Y2=1.055
r101 11 34 38.7839 $w=3.5e-07 $l=2.09105e-07 $layer=POLY_cond $X=5.155 $Y=1.385
+ $X2=5.055 $Y2=1.22
r102 11 13 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=5.155 $Y=1.385
+ $X2=5.155 $Y2=2.315
r103 7 34 44.2925 $w=3.5e-07 $l=2.56125e-07 $layer=POLY_cond $X=4.94 $Y=1.015
+ $X2=5.055 $Y2=1.22
r104 7 9 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.94 $Y=1.015
+ $X2=4.94 $Y2=0.555
r105 2 25 600 $w=1.7e-07 $l=3.58504e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=2.315 $X2=3.485 $Y2=2.58
r106 1 22 182 $w=1.7e-07 $l=3.11127e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.305 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_1091_21# 1 2 7 9 12 16 20 23 26 27 29 30
+ 32 33 34 36 37 38 39 41 44 45 46 48 50
c178 23 0 3.03962e-19 $X=9.375 $Y=1.51
c179 12 0 9.56299e-20 $X=5.545 $Y=2.315
r180 59 61 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.53 $Y=1.15
+ $X2=5.545 $Y2=1.15
r181 50 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.825 $Y=0.86
+ $X2=8.825 $Y2=1.03
r182 46 48 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=10.01 $Y=1.86
+ $X2=10.23 $Y2=1.86
r183 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.845
+ $Y=1.39 $X2=9.845 $Y2=1.39
r184 42 46 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=9.845 $Y=1.695
+ $X2=10.01 $Y2=1.86
r185 42 44 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=9.845 $Y=1.695
+ $X2=9.845 $Y2=1.39
r186 41 56 16.4637 $w=2.89e-07 $l=3.9e-07 $layer=LI1_cond $X=9.845 $Y=0.817
+ $X2=10.235 $Y2=0.817
r187 41 44 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=9.845 $Y=1
+ $X2=9.845 $Y2=1.39
r188 40 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=0.86
+ $X2=8.825 $Y2=0.86
r189 39 41 9.01683 $w=2.89e-07 $l=1.85257e-07 $layer=LI1_cond $X=9.68 $Y=0.86
+ $X2=9.845 $Y2=0.817
r190 39 40 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=9.68 $Y=0.86
+ $X2=8.91 $Y2=0.86
r191 37 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.74 $Y=1.03
+ $X2=8.825 $Y2=1.03
r192 37 38 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=8.74 $Y=1.03
+ $X2=7.835 $Y2=1.03
r193 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.75 $Y=0.945
+ $X2=7.835 $Y2=1.03
r194 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.75 $Y=0.435
+ $X2=7.75 $Y2=0.945
r195 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.665 $Y=0.35
+ $X2=7.75 $Y2=0.435
r196 33 34 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=7.665 $Y=0.35
+ $X2=6.74 $Y2=0.35
r197 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.655 $Y=0.435
+ $X2=6.74 $Y2=0.35
r198 31 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.655 $Y=0.435
+ $X2=6.655 $Y2=0.76
r199 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.57 $Y=0.845
+ $X2=6.655 $Y2=0.76
r200 29 30 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=6.57 $Y=0.845
+ $X2=6.015 $Y2=0.845
r201 27 61 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=5.85 $Y=1.15
+ $X2=5.545 $Y2=1.15
r202 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.85
+ $Y=1.15 $X2=5.85 $Y2=1.15
r203 24 30 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=5.872 $Y=0.93
+ $X2=6.015 $Y2=0.845
r204 24 26 8.89605 $w=2.83e-07 $l=2.2e-07 $layer=LI1_cond $X=5.872 $Y=0.93
+ $X2=5.872 $Y2=1.15
r205 22 45 38.9947 $w=4.35e-07 $l=3.05e-07 $layer=POLY_cond $X=9.54 $Y=1.442
+ $X2=9.845 $Y2=1.442
r206 22 23 8.05214 $w=4.35e-07 $l=1.96074e-07 $layer=POLY_cond $X=9.54 $Y=1.442
+ $X2=9.375 $Y2=1.51
r207 18 23 44.2338 $w=1.5e-07 $l=3.26917e-07 $layer=POLY_cond $X=9.465 $Y=1.225
+ $X2=9.375 $Y2=1.51
r208 18 20 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.465 $Y=1.225
+ $X2=9.465 $Y2=0.59
r209 14 23 44.2338 $w=1.5e-07 $l=1.83712e-07 $layer=POLY_cond $X=9.45 $Y=1.66
+ $X2=9.375 $Y2=1.51
r210 14 16 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=9.45 $Y=1.66
+ $X2=9.45 $Y2=2.57
r211 10 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.545 $Y=1.315
+ $X2=5.545 $Y2=1.15
r212 10 12 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=5.545 $Y=1.315
+ $X2=5.545 $Y2=2.315
r213 7 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.53 $Y=0.985
+ $X2=5.53 $Y2=1.15
r214 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.53 $Y=0.985
+ $X2=5.53 $Y2=0.555
r215 2 48 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.085
+ $Y=1.715 $X2=10.23 $Y2=1.86
r216 1 56 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=10.09
+ $Y=0.655 $X2=10.235 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_114_57# 1 2 9 13 18 19 20 21 22 23 27 31
+ 33 35 38 39 43 47 51 57 58 60 63 66
c157 43 0 1.68286e-19 $X=7.42 $Y=0.7
c158 31 0 1.44713e-19 $X=3.7 $Y=2.525
r159 65 66 33.5808 $w=1.78e-07 $l=5.45e-07 $layer=LI1_cond $X=0.785 $Y=0.725
+ $X2=0.785 $Y2=1.27
r160 63 65 10.3964 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.71 $Y=0.495
+ $X2=0.71 $Y2=0.725
r161 57 66 8.12648 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=1.435
+ $X2=0.86 $Y2=1.27
r162 57 60 38.9386 $w=3.28e-07 $l=1.115e-06 $layer=LI1_cond $X=0.86 $Y=1.435
+ $X2=0.86 $Y2=2.55
r163 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.86
+ $Y=1.435 $X2=0.86 $Y2=1.435
r164 47 49 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.385 $Y=1.23
+ $X2=2.385 $Y2=1.41
r165 45 46 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.635 $Y2=1.41
r166 41 43 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=7.42 $Y=1.68
+ $X2=7.42 $Y2=0.7
r167 40 52 12.4931 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.735 $Y=1.755
+ $X2=6.585 $Y2=1.755
r168 39 41 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.345 $Y=1.755
+ $X2=7.42 $Y2=1.68
r169 39 40 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.345 $Y=1.755
+ $X2=6.735 $Y2=1.755
r170 36 38 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=6.46 $Y=3.075
+ $X2=6.46 $Y2=2.56
r171 35 52 71.3749 $w=2.27e-07 $l=3.67219e-07 $layer=POLY_cond $X=6.46 $Y=2.065
+ $X2=6.585 $Y2=1.755
r172 35 38 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.46 $Y=2.065
+ $X2=6.46 $Y2=2.56
r173 34 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.775 $Y=3.15
+ $X2=3.7 $Y2=3.15
r174 33 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.385 $Y=3.15
+ $X2=6.46 $Y2=3.075
r175 33 34 1338.32 $w=1.5e-07 $l=2.61e-06 $layer=POLY_cond $X=6.385 $Y=3.15
+ $X2=3.775 $Y2=3.15
r176 29 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.7 $Y=3.075
+ $X2=3.7 $Y2=3.15
r177 29 31 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.7 $Y=3.075
+ $X2=3.7 $Y2=2.525
r178 25 27 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.01 $Y=1.155
+ $X2=3.01 $Y2=0.445
r179 24 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.46 $Y=1.23
+ $X2=2.385 $Y2=1.23
r180 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.935 $Y=1.23
+ $X2=3.01 $Y2=1.155
r181 23 24 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=2.935 $Y=1.23
+ $X2=2.46 $Y2=1.23
r182 21 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.625 $Y=3.15
+ $X2=3.7 $Y2=3.15
r183 21 22 981.947 $w=1.5e-07 $l=1.915e-06 $layer=POLY_cond $X=3.625 $Y=3.15
+ $X2=1.71 $Y2=3.15
r184 20 46 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.71 $Y=1.41
+ $X2=1.635 $Y2=1.41
r185 19 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.31 $Y=1.41
+ $X2=2.385 $Y2=1.41
r186 19 20 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.31 $Y=1.41 $X2=1.71
+ $Y2=1.41
r187 16 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.635 $Y=3.075
+ $X2=1.71 $Y2=3.15
r188 16 18 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.635 $Y=3.075
+ $X2=1.635 $Y2=2.635
r189 15 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.635 $Y=1.485
+ $X2=1.635 $Y2=1.41
r190 15 18 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=1.635 $Y=1.485
+ $X2=1.635 $Y2=2.635
r191 11 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.485 $Y=1.335
+ $X2=1.485 $Y2=1.41
r192 11 13 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.485 $Y=1.335
+ $X2=1.485 $Y2=0.445
r193 10 58 20.8207 $w=1.5e-07 $l=1.80748e-07 $layer=POLY_cond $X=1.025 $Y=1.41
+ $X2=0.86 $Y2=1.377
r194 9 45 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.41
+ $X2=1.485 $Y2=1.41
r195 9 10 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.41 $Y=1.41
+ $X2=1.025 $Y2=1.41
r196 2 60 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.72
+ $Y=2.405 $X2=0.86 $Y2=2.55
r197 1 63 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.285 $X2=0.71 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_1545_332# 1 2 9 13 17 21 22 24 26 29 31 34
+ 35 37 38 41 43 46 47 50 52 56 58 62 68 69
c180 52 0 4.06414e-20 $X=8.825 $Y=2.31
c181 34 0 1.68286e-19 $X=7.89 $Y=1.825
c182 9 0 6.36774e-20 $X=7.81 $Y=0.7
r183 68 69 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.93 $Y=1.26
+ $X2=10.93 $Y2=1.185
r184 63 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.93 $Y=1.35
+ $X2=10.93 $Y2=1.515
r185 63 68 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.93 $Y=1.35
+ $X2=10.93 $Y2=1.26
r186 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.93
+ $Y=1.35 $X2=10.93 $Y2=1.35
r187 59 62 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=10.82 $Y=1.35
+ $X2=10.93 $Y2=1.35
r188 54 56 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=9.175 $Y=1.29
+ $X2=9.4 $Y2=1.29
r189 49 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.82 $Y=1.515
+ $X2=10.82 $Y2=1.35
r190 49 50 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.82 $Y=1.515
+ $X2=10.82 $Y2=2.205
r191 48 58 4.50329 $w=2e-07 $l=9.88686e-08 $layer=LI1_cond $X=9.485 $Y=2.29
+ $X2=9.4 $Y2=2.26
r192 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.735 $Y=2.29
+ $X2=10.82 $Y2=2.205
r193 47 48 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=10.735 $Y=2.29
+ $X2=9.485 $Y2=2.29
r194 46 58 1.93381 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.4 $Y=2.145
+ $X2=9.4 $Y2=2.26
r195 45 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.4 $Y=1.455
+ $X2=9.4 $Y2=1.29
r196 45 46 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.4 $Y=1.455 $X2=9.4
+ $Y2=2.145
r197 44 52 6.19399 $w=2e-07 $l=1.52889e-07 $layer=LI1_cond $X=8.99 $Y=2.26
+ $X2=8.865 $Y2=2.322
r198 43 58 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=9.315 $Y=2.26 $X2=9.4
+ $Y2=2.26
r199 43 44 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=9.315 $Y=2.26
+ $X2=8.99 $Y2=2.26
r200 39 52 0.552779 $w=2.5e-07 $l=1.78e-07 $layer=LI1_cond $X=8.865 $Y=2.5
+ $X2=8.865 $Y2=2.322
r201 39 41 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=8.865 $Y=2.5
+ $X2=8.865 $Y2=2.845
r202 37 52 6.19399 $w=2e-07 $l=1.65076e-07 $layer=LI1_cond $X=8.74 $Y=2.415
+ $X2=8.865 $Y2=2.322
r203 37 38 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=8.74 $Y=2.415
+ $X2=8.055 $Y2=2.415
r204 35 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.89 $Y=1.825
+ $X2=7.89 $Y2=1.99
r205 35 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.89 $Y=1.825
+ $X2=7.89 $Y2=1.66
r206 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.89
+ $Y=1.825 $X2=7.89 $Y2=1.825
r207 32 38 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=7.91 $Y=2.33
+ $X2=8.055 $Y2=2.415
r208 32 34 20.0684 $w=2.88e-07 $l=5.05e-07 $layer=LI1_cond $X=7.91 $Y=2.33
+ $X2=7.91 $Y2=1.825
r209 27 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.945 $Y=1.335
+ $X2=11.945 $Y2=1.26
r210 27 29 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=11.945 $Y=1.335
+ $X2=11.945 $Y2=2.155
r211 24 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.945 $Y=1.185
+ $X2=11.945 $Y2=1.26
r212 24 26 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.945 $Y=1.185
+ $X2=11.945 $Y2=0.865
r213 23 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.095 $Y=1.26
+ $X2=10.93 $Y2=1.26
r214 22 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.87 $Y=1.26
+ $X2=11.945 $Y2=1.26
r215 22 23 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=11.87 $Y=1.26
+ $X2=11.095 $Y2=1.26
r216 21 69 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.96 $Y=0.655
+ $X2=10.96 $Y2=1.185
r217 17 71 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=10.955 $Y=2.345
+ $X2=10.955 $Y2=1.515
r218 13 67 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.81 $Y=2.77
+ $X2=7.81 $Y2=1.99
r219 9 66 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=7.81 $Y=0.7 $X2=7.81
+ $Y2=1.66
r220 2 52 600 $w=1.7e-07 $l=2.995e-07 $layer=licon1_PDIFF $count=1 $X=8.595
+ $Y=2.15 $X2=8.825 $Y2=2.31
r221 2 41 600 $w=1.7e-07 $l=8.01795e-07 $layer=licon1_PDIFF $count=1 $X=8.595
+ $Y=2.15 $X2=8.825 $Y2=2.845
r222 1 54 182 $w=1.7e-07 $l=1.12463e-06 $layer=licon1_NDIFF $count=1 $X=8.955
+ $Y=0.27 $X2=9.175 $Y2=1.29
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_1307_428# 1 2 9 13 15 19 22 24 25 28 29 34
+ 38 39
c121 28 0 1.66022e-19 $X=8.825 $Y=1.635
c122 25 0 1.3794e-19 $X=8.74 $Y=1.395
c123 13 0 6.36774e-20 $X=9.04 $Y=2.57
r124 39 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.97 $Y=1.8
+ $X2=8.97 $Y2=1.965
r125 39 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.97 $Y=1.8
+ $X2=8.97 $Y2=1.635
r126 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.97
+ $Y=1.8 $X2=8.97 $Y2=1.8
r127 35 38 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.825 $Y=1.8
+ $X2=8.97 $Y2=1.8
r128 29 32 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=6.805 $Y=2.665
+ $X2=6.805 $Y2=2.79
r129 28 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.825 $Y=1.635
+ $X2=8.825 $Y2=1.8
r130 27 28 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.825 $Y=1.48
+ $X2=8.825 $Y2=1.635
r131 26 34 1.34256 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.585 $Y=1.395
+ $X2=7.45 $Y2=1.395
r132 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.74 $Y=1.395
+ $X2=8.825 $Y2=1.48
r133 25 26 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=8.74 $Y=1.395
+ $X2=7.585 $Y2=1.395
r134 23 34 5.16603 $w=1.7e-07 $l=1.07121e-07 $layer=LI1_cond $X=7.5 $Y=1.48
+ $X2=7.45 $Y2=1.395
r135 23 24 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=7.5 $Y=1.48 $X2=7.5
+ $Y2=2.58
r136 22 34 5.16603 $w=1.7e-07 $l=1.07121e-07 $layer=LI1_cond $X=7.4 $Y=1.31
+ $X2=7.45 $Y2=1.395
r137 21 22 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.4 $Y=0.93 $X2=7.4
+ $Y2=1.31
r138 20 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.97 $Y=2.665
+ $X2=6.805 $Y2=2.665
r139 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.415 $Y=2.665
+ $X2=7.5 $Y2=2.58
r140 19 20 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7.415 $Y=2.665
+ $X2=6.97 $Y2=2.665
r141 15 21 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.315 $Y=0.772
+ $X2=7.4 $Y2=0.93
r142 15 17 6.95124 $w=3.13e-07 $l=1.9e-07 $layer=LI1_cond $X=7.315 $Y=0.772
+ $X2=7.125 $Y2=0.772
r143 13 43 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=9.04 $Y=2.57
+ $X2=9.04 $Y2=1.965
r144 9 42 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=8.88 $Y=0.59
+ $X2=8.88 $Y2=1.635
r145 2 32 600 $w=1.7e-07 $l=7.73305e-07 $layer=licon1_PDIFF $count=1 $X=6.535
+ $Y=2.14 $X2=6.805 $Y2=2.79
r146 1 17 182 $w=1.7e-07 $l=5.25357e-07 $layer=licon1_NDIFF $count=1 $X=6.985
+ $Y=0.27 $X2=7.125 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%RESET_B 3 7 8 11 13
c32 13 0 1.37641e-19 $X=10.385 $Y=1.185
r33 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.385 $Y=1.35
+ $X2=10.385 $Y2=1.515
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.385 $Y=1.35
+ $X2=10.385 $Y2=1.185
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.385
+ $Y=1.35 $X2=10.385 $Y2=1.35
r36 7 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.45 $Y=0.865
+ $X2=10.45 $Y2=1.185
r37 3 14 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=10.445 $Y=2.035
+ $X2=10.445 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_2317_367# 1 2 9 13 17 21 23 24 25 26 29 30
c61 21 0 1.83005e-19 $X=11.73 $Y=1.98
r62 30 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.395 $Y=1.47
+ $X2=12.395 $Y2=1.635
r63 30 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.395 $Y=1.47
+ $X2=12.395 $Y2=1.305
r64 29 31 3.33106 $w=2.93e-07 $l=8e-08 $layer=LI1_cond $X=12.337 $Y=1.47
+ $X2=12.337 $Y2=1.55
r65 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.395
+ $Y=1.47 $X2=12.395 $Y2=1.47
r66 25 31 3.92235 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=12.155 $Y=1.55
+ $X2=12.337 $Y2=1.55
r67 25 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.155 $Y=1.55
+ $X2=11.895 $Y2=1.55
r68 23 29 11.2423 $w=2.93e-07 $l=3.49342e-07 $layer=LI1_cond $X=12.155 $Y=1.2
+ $X2=12.337 $Y2=1.47
r69 23 24 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.155 $Y=1.2
+ $X2=11.895 $Y2=1.2
r70 19 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.77 $Y=1.635
+ $X2=11.895 $Y2=1.55
r71 19 21 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=11.77 $Y=1.635
+ $X2=11.77 $Y2=1.98
r72 15 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.77 $Y=1.115
+ $X2=11.895 $Y2=1.2
r73 15 17 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=11.77 $Y=1.115
+ $X2=11.77 $Y2=0.865
r74 13 34 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=12.455 $Y=2.465
+ $X2=12.455 $Y2=1.635
r75 9 33 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=12.455 $Y=0.655
+ $X2=12.455 $Y2=1.305
r76 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=11.585
+ $Y=1.835 $X2=11.73 $Y2=1.98
r77 1 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.59
+ $Y=0.655 $X2=11.73 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 43 47 51
+ 55 60 61 63 64 66 67 68 77 88 99 103 110 111 117 120 123 126
r142 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r143 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r144 120 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r145 117 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r146 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r147 111 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r148 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r149 108 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.2 $Y2=3.33
r150 108 110 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.72 $Y2=3.33
r151 107 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r152 107 124 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=10.8 $Y2=3.33
r153 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r154 104 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=10.74 $Y2=3.33
r155 104 106 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=11.76 $Y2=3.33
r156 103 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.075 $Y=3.33
+ $X2=12.2 $Y2=3.33
r157 103 106 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.075 $Y=3.33
+ $X2=11.76 $Y2=3.33
r158 102 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r159 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r160 99 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.575 $Y=3.33
+ $X2=10.74 $Y2=3.33
r161 99 101 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.575 $Y=3.33
+ $X2=10.32 $Y2=3.33
r162 98 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r163 98 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.4 $Y2=3.33
r164 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r165 95 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=8.305 $Y2=3.33
r166 95 97 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=9.36 $Y2=3.33
r167 94 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r168 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r169 90 93 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.92
+ $Y2=3.33
r170 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r171 88 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=8.305 $Y2=3.33
r172 88 93 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=7.92 $Y2=3.33
r173 87 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r174 87 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r175 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r176 84 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.595 $Y=3.33
+ $X2=4.43 $Y2=3.33
r177 84 86 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.595 $Y=3.33
+ $X2=5.52 $Y2=3.33
r178 83 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r179 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r180 80 83 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r181 79 82 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r182 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r183 77 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.265 $Y=3.33
+ $X2=4.43 $Y2=3.33
r184 77 82 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.265 $Y=3.33
+ $X2=4.08 $Y2=3.33
r185 76 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r186 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r187 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r188 73 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r189 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r190 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r191 70 114 4.59558 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=0.515 $Y=3.33
+ $X2=0.257 $Y2=3.33
r192 70 72 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.515 $Y=3.33
+ $X2=0.72 $Y2=3.33
r193 68 94 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r194 68 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r195 66 97 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=9.5 $Y=3.33
+ $X2=9.36 $Y2=3.33
r196 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.5 $Y=3.33
+ $X2=9.665 $Y2=3.33
r197 65 101 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=9.83 $Y=3.33
+ $X2=10.32 $Y2=3.33
r198 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.83 $Y=3.33
+ $X2=9.665 $Y2=3.33
r199 63 86 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.595 $Y=3.33
+ $X2=5.52 $Y2=3.33
r200 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.595 $Y=3.33
+ $X2=5.76 $Y2=3.33
r201 62 90 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.925 $Y=3.33 $X2=6
+ $Y2=3.33
r202 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.925 $Y=3.33
+ $X2=5.76 $Y2=3.33
r203 60 75 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.68 $Y2=3.33
r204 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.93 $Y2=3.33
r205 59 79 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=2.16 $Y2=3.33
r206 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=1.93 $Y2=3.33
r207 55 58 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=12.2 $Y=1.98
+ $X2=12.2 $Y2=2.465
r208 53 126 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.2 $Y=3.245
+ $X2=12.2 $Y2=3.33
r209 53 58 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=12.2 $Y=3.245
+ $X2=12.2 $Y2=2.465
r210 49 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=3.245
+ $X2=10.74 $Y2=3.33
r211 49 51 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=10.74 $Y=3.245
+ $X2=10.74 $Y2=2.775
r212 45 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.665 $Y=3.245
+ $X2=9.665 $Y2=3.33
r213 45 47 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.665 $Y=3.245
+ $X2=9.665 $Y2=2.78
r214 41 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.305 $Y=3.245
+ $X2=8.305 $Y2=3.33
r215 41 43 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=8.305 $Y=3.245
+ $X2=8.305 $Y2=2.845
r216 37 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=3.245
+ $X2=5.76 $Y2=3.33
r217 37 39 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=5.76 $Y=3.245
+ $X2=5.76 $Y2=2.53
r218 33 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.43 $Y=3.245
+ $X2=4.43 $Y2=3.33
r219 33 35 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.43 $Y=3.245 $X2=4.43
+ $Y2=2.845
r220 29 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r221 29 31 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.78
r222 25 114 3.17059 $w=3.3e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.35 $Y=3.245
+ $X2=0.257 $Y2=3.33
r223 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.35 $Y=3.245
+ $X2=0.35 $Y2=2.55
r224 8 58 300 $w=1.7e-07 $l=7.31779e-07 $layer=licon1_PDIFF $count=2 $X=12.02
+ $Y=1.835 $X2=12.24 $Y2=2.465
r225 8 55 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=12.02
+ $Y=1.835 $X2=12.24 $Y2=1.98
r226 7 51 600 $w=1.7e-07 $l=1.16482e-06 $layer=licon1_PDIFF $count=1 $X=10.52
+ $Y=1.715 $X2=10.74 $Y2=2.775
r227 6 47 600 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=1 $X=9.525
+ $Y=2.15 $X2=9.665 $Y2=2.78
r228 5 43 600 $w=1.7e-07 $l=5.44151e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=2.56 $X2=8.305 $Y2=2.845
r229 4 39 600 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=1 $X=5.62
+ $Y=1.895 $X2=5.76 $Y2=2.53
r230 3 35 600 $w=1.7e-07 $l=6.49115e-07 $layer=licon1_PDIFF $count=1 $X=4.165
+ $Y=2.315 $X2=4.43 $Y2=2.845
r231 2 31 600 $w=1.7e-07 $l=5.6438e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.315 $X2=1.93 $Y2=2.78
r232 1 27 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.205
+ $Y=2.405 $X2=0.35 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_531_47# 1 2 9 13 15 16 18 21
c62 21 0 1.44713e-19 $X=3.265 $Y=2.145
c63 16 0 5.88079e-20 $X=2.96 $Y=0.915
r64 18 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=2.06
+ $X2=3.265 $Y2=2.145
r65 17 18 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.265 $Y=1
+ $X2=3.265 $Y2=2.06
r66 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.18 $Y=0.915
+ $X2=3.265 $Y2=1
r67 15 16 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.18 $Y=0.915
+ $X2=2.96 $Y2=0.915
r68 11 21 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.975 $Y=2.145
+ $X2=3.265 $Y2=2.145
r69 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.975 $Y=2.23
+ $X2=2.975 $Y2=2.525
r70 7 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.795 $Y=0.83
+ $X2=2.96 $Y2=0.915
r71 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.795 $Y=0.83
+ $X2=2.795 $Y2=0.47
r72 2 13 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.835
+ $Y=2.315 $X2=2.975 $Y2=2.525
r73 1 9 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.655
+ $Y=0.235 $X2=2.795 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%Q_N 1 2 9 13 16 17 18 19 20
c36 9 0 1.37641e-19 $X=11.175 $Y=0.43
r37 20 31 1.76068 $w=3.58e-07 $l=5.5e-08 $layer=LI1_cond $X=11.265 $Y=2.775
+ $X2=11.265 $Y2=2.83
r38 19 20 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=11.265 $Y=2.405
+ $X2=11.265 $Y2=2.775
r39 18 19 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=11.265 $Y=2.035
+ $X2=11.265 $Y2=2.405
r40 16 17 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=11.265 $Y=1.86
+ $X2=11.265 $Y2=1.695
r41 14 18 5.12197 $w=3.58e-07 $l=1.6e-07 $layer=LI1_cond $X=11.265 $Y=1.875
+ $X2=11.265 $Y2=2.035
r42 14 16 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=11.265 $Y=1.875
+ $X2=11.265 $Y2=1.86
r43 13 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.36 $Y=1.005
+ $X2=11.36 $Y2=1.695
r44 7 13 10.1875 $w=4.33e-07 $l=2.17e-07 $layer=LI1_cond $X=11.227 $Y=0.788
+ $X2=11.227 $Y2=1.005
r45 7 9 9.48447 $w=4.33e-07 $l=3.58e-07 $layer=LI1_cond $X=11.227 $Y=0.788
+ $X2=11.227 $Y2=0.43
r46 2 31 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=11.03
+ $Y=1.715 $X2=11.17 $Y2=2.83
r47 2 16 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.03
+ $Y=1.715 $X2=11.17 $Y2=1.86
r48 1 9 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=11.035
+ $Y=0.235 $X2=11.175 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%Q 1 2 9 14 15 16 17 23 29
r27 21 29 0.378885 $w=3.63e-07 $l=1.2e-08 $layer=LI1_cond $X=12.687 $Y=0.913
+ $X2=12.687 $Y2=0.925
r28 17 31 7.54552 $w=3.63e-07 $l=1.34e-07 $layer=LI1_cond $X=12.687 $Y=0.961
+ $X2=12.687 $Y2=1.095
r29 17 29 1.13666 $w=3.63e-07 $l=3.6e-08 $layer=LI1_cond $X=12.687 $Y=0.961
+ $X2=12.687 $Y2=0.925
r30 17 21 1.16823 $w=3.63e-07 $l=3.7e-08 $layer=LI1_cond $X=12.687 $Y=0.876
+ $X2=12.687 $Y2=0.913
r31 16 17 10.1352 $w=3.63e-07 $l=3.21e-07 $layer=LI1_cond $X=12.687 $Y=0.555
+ $X2=12.687 $Y2=0.876
r32 16 23 3.94672 $w=3.63e-07 $l=1.25e-07 $layer=LI1_cond $X=12.687 $Y=0.555
+ $X2=12.687 $Y2=0.43
r33 15 31 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=12.785 $Y=1.815
+ $X2=12.785 $Y2=1.095
r34 14 15 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=12.687 $Y=1.98
+ $X2=12.687 $Y2=1.815
r35 7 14 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=12.687 $Y=1.997
+ $X2=12.687 $Y2=1.98
r36 7 9 28.5111 $w=3.63e-07 $l=9.03e-07 $layer=LI1_cond $X=12.687 $Y=1.997
+ $X2=12.687 $Y2=2.9
r37 2 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.835 $X2=12.67 $Y2=1.98
r38 2 9 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.835 $X2=12.67 $Y2=2.9
r39 1 23 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=12.53
+ $Y=0.235 $X2=12.67 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 50
+ 55 56 58 59 61 62 63 72 89 96 103 104 110 113 116
r145 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r146 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r147 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r148 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r149 104 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r150 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r151 101 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.325 $Y=0
+ $X2=12.2 $Y2=0
r152 101 103 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.325 $Y=0
+ $X2=12.72 $Y2=0
r153 100 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r154 100 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=10.8 $Y2=0
r155 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r156 97 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.83 $Y=0
+ $X2=10.705 $Y2=0
r157 97 99 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=10.83 $Y=0
+ $X2=11.76 $Y2=0
r158 96 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=12.2 $Y2=0
r159 96 99 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=11.76 $Y2=0
r160 95 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r161 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r162 92 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=10.32 $Y2=0
r163 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=10.32
+ $Y2=0
r164 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r165 89 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.58 $Y=0
+ $X2=10.705 $Y2=0
r166 89 94 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=10.58 $Y=0
+ $X2=10.32 $Y2=0
r167 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r168 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r169 84 87 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.92
+ $Y2=0
r170 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r171 79 82 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r172 79 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r173 78 81 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r174 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r175 76 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.38 $Y=0
+ $X2=4.215 $Y2=0
r176 76 78 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.38 $Y=0 $X2=4.56
+ $Y2=0
r177 75 111 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r178 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r179 72 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=0
+ $X2=4.215 $Y2=0
r180 72 74 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=4.05 $Y=0 $X2=2.16
+ $Y2=0
r181 71 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r182 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r183 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r184 68 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r185 67 70 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r186 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r187 65 107 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r188 65 67 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r189 63 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r190 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r191 63 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r192 61 87 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=7.92
+ $Y2=0
r193 61 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=8.195
+ $Y2=0
r194 60 91 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=8.32 $Y=0 $X2=8.4
+ $Y2=0
r195 60 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.32 $Y=0 $X2=8.195
+ $Y2=0
r196 58 81 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6
+ $Y2=0
r197 58 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6.265
+ $Y2=0
r198 57 84 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.39 $Y=0 $X2=6.48
+ $Y2=0
r199 57 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.39 $Y=0 $X2=6.265
+ $Y2=0
r200 55 70 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r201 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.93
+ $Y2=0
r202 54 74 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.16
+ $Y2=0
r203 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=1.93
+ $Y2=0
r204 50 52 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=12.2 $Y=0.38
+ $X2=12.2 $Y2=0.77
r205 48 116 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.2 $Y=0.085
+ $X2=12.2 $Y2=0
r206 48 50 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=12.2 $Y=0.085
+ $X2=12.2 $Y2=0.38
r207 44 46 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=10.705 $Y=0.38
+ $X2=10.705 $Y2=0.835
r208 42 113 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.705 $Y=0.085
+ $X2=10.705 $Y2=0
r209 42 44 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=10.705 $Y=0.085
+ $X2=10.705 $Y2=0.38
r210 38 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.195 $Y=0.085
+ $X2=8.195 $Y2=0
r211 38 40 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=8.195 $Y=0.085
+ $X2=8.195 $Y2=0.505
r212 34 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.265 $Y=0.085
+ $X2=6.265 $Y2=0
r213 34 36 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=6.265 $Y=0.085
+ $X2=6.265 $Y2=0.415
r214 30 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0
r215 30 32 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0.545
r216 26 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0
r217 26 28 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0.4
r218 22 107 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r219 22 24 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.495
r220 7 52 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=12.02
+ $Y=0.655 $X2=12.24 $Y2=0.77
r221 7 50 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=12.02
+ $Y=0.655 $X2=12.24 $Y2=0.38
r222 6 46 182 $w=1.7e-07 $l=2.96648e-07 $layer=licon1_NDIFF $count=1 $X=10.525
+ $Y=0.655 $X2=10.745 $Y2=0.835
r223 6 44 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=10.525
+ $Y=0.655 $X2=10.745 $Y2=0.38
r224 5 40 182 $w=1.7e-07 $l=2.77399e-07 $layer=licon1_NDIFF $count=1 $X=7.885
+ $Y=0.49 $X2=8.155 $Y2=0.505
r225 4 36 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.16
+ $Y=0.27 $X2=6.305 $Y2=0.415
r226 3 32 182 $w=1.7e-07 $l=4.09145e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.235 $X2=4.215 $Y2=0.545
r227 2 28 182 $w=1.7e-07 $l=4.44916e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.93 $Y2=0.4
r228 1 24 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_917_47# 1 2 9 12 14 15
r26 14 15 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.745 $Y=0.395
+ $X2=5.58 $Y2=0.395
r27 12 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.89 $Y=0.35 $X2=5.58
+ $Y2=0.35
r28 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.725 $Y=0.435
+ $X2=4.89 $Y2=0.35
r29 7 9 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.725 $Y=0.435
+ $X2=4.725 $Y2=0.57
r30 2 14 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=5.605
+ $Y=0.235 $X2=5.745 $Y2=0.41
r31 1 9 182 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=1 $X=4.585
+ $Y=0.235 $X2=4.725 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBP_1%A_1705_54# 1 2 11
r17 8 11 35.4464 $w=3.28e-07 $l=1.015e-06 $layer=LI1_cond $X=8.665 $Y=0.43
+ $X2=9.68 $Y2=0.43
r18 2 11 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=9.54
+ $Y=0.27 $X2=9.68 $Y2=0.43
r19 1 8 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=8.525
+ $Y=0.27 $X2=8.665 $Y2=0.43
.ends

