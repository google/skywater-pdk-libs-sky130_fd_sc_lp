* File: sky130_fd_sc_lp__o2bb2a_lp.spice
* Created: Wed Sep  2 10:21:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2a_lp  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1009 A_116_48# N_A_86_22#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_86_22#_M1006_g A_116_48# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1010 A_274_48# N_A1_N_M1010_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_A_298_416#_M1011_d N_A2_N_M1011_g A_274_48# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_604_142#_M1012_d N_A_298_416#_M1012_g N_A_86_22#_M1012_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1449 PD=0.72 PS=1.53 NRD=5.712 NRS=17.136 M=1
+ R=2.8 SA=75000.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_B2_M1001_g N_A_604_142#_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.063 PD=0.7 PS=0.72 NRD=0 NRS=0 M=1 R=2.8 SA=75000.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_604_142#_M1003_d N_B1_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_86_22#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.28 AS=0.285 PD=1.56 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1007 N_A_298_416#_M1007_d N_A1_N_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.155 AS=0.28 PD=1.31 PS=1.56 NRD=5.8903 NRS=55.1403 M=1 R=4 SA=125001
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A2_N_M1004_g N_A_298_416#_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.27 AS=0.155 PD=1.54 PS=1.31 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1000 N_A_86_22#_M1000_d N_A_298_416#_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.27 PD=1.28 PS=1.54 NRD=0 NRS=51.2003 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1008 A_674_416# N_B2_M1008_g N_A_86_22#_M1000_d VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=16.7253 NRS=0 M=1 R=4 SA=125003 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g A_674_416# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=16.7253 M=1 R=4 SA=125003 SB=125000 A=0.25
+ P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__o2bb2a_lp.pxi.spice"
*
.ends
*
*
