* File: sky130_fd_sc_lp__dlymetal6s6s_1.pex.spice
* Created: Fri Aug 28 10:31:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A 3 7 9 12 13
c28 7 0 4.97211e-20 $X=0.475 $Y=2.045
r29 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.44
+ $X2=0.385 $Y2=1.605
r30 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.44
+ $X2=0.385 $Y2=1.275
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.44 $X2=0.385 $Y2=1.44
r32 9 13 5.98039 $w=4.48e-07 $l=2.25e-07 $layer=LI1_cond $X=0.325 $Y=1.665
+ $X2=0.325 $Y2=1.44
r33 7 15 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.475 $Y=2.045
+ $X2=0.475 $Y2=1.605
r34 3 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.475 $Y=0.865
+ $X2=0.475 $Y2=1.275
.ends

.subckt PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_27_131# 1 2 9 13 15 17 19 20 22 29
+ 33
c60 19 0 1.89796e-19 $X=0.805 $Y=1.605
r61 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.44
+ $X2=0.925 $Y2=1.605
r62 33 35 48.8344 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.925 $Y=1.44
+ $X2=0.925 $Y2=1.26
r63 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.44 $X2=0.925 $Y2=1.44
r64 30 32 19.9828 $w=2.32e-07 $l=3.8e-07 $layer=LI1_cond $X=0.865 $Y=1.06
+ $X2=0.865 $Y2=1.44
r65 27 29 7.16645 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=2.08
+ $X2=0.425 $Y2=2.08
r66 22 24 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=0.242 $Y=0.865
+ $X2=0.242 $Y2=1.06
r67 19 32 9.57122 $w=2.32e-07 $l=1.92678e-07 $layer=LI1_cond $X=0.805 $Y=1.605
+ $X2=0.865 $Y2=1.44
r68 19 20 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.805 $Y=1.605
+ $X2=0.805 $Y2=1.935
r69 17 20 6.9898 $w=2.25e-07 $l=1.4854e-07 $layer=LI1_cond $X=0.72 $Y=2.047
+ $X2=0.805 $Y2=1.935
r70 17 29 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=2.047
+ $X2=0.425 $Y2=2.047
r71 16 24 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.39 $Y=1.06
+ $X2=0.242 $Y2=1.06
r72 15 30 2.55969 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.72 $Y=1.06
+ $X2=0.865 $Y2=1.06
r73 15 16 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.72 $Y=1.06
+ $X2=0.39 $Y2=1.06
r74 13 36 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.965 $Y=2.465
+ $X2=0.965 $Y2=1.605
r75 9 35 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=0.965 $Y=0.655
+ $X2=0.965 $Y2=1.26
r76 2 27 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.06
r77 1 22 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.655 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_208_47# 1 2 9 13 17 20 25 26 28 29
+ 30 31 41
c64 26 0 1.89796e-19 $X=1.825 $Y=1.44
r65 41 43 36.1629 $w=2.88e-07 $l=9.1e-07 $layer=LI1_cond $X=1.205 $Y=2 $X2=1.205
+ $Y2=2.91
r66 28 41 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=1.205 $Y=1.98
+ $X2=1.205 $Y2=2
r67 28 29 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.205 $Y=1.98
+ $X2=1.205 $Y2=1.835
r68 26 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.44
+ $X2=1.825 $Y2=1.605
r69 26 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.44
+ $X2=1.825 $Y2=1.275
r70 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.44 $X2=1.825 $Y2=1.44
r71 23 31 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=1.46
+ $X2=1.265 $Y2=1.46
r72 23 25 18.8762 $w=2.88e-07 $l=4.75e-07 $layer=LI1_cond $X=1.35 $Y=1.46
+ $X2=1.825 $Y2=1.46
r73 21 31 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.265 $Y=1.605
+ $X2=1.265 $Y2=1.46
r74 21 29 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.265 $Y=1.605
+ $X2=1.265 $Y2=1.835
r75 20 31 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.265 $Y=1.315
+ $X2=1.265 $Y2=1.46
r76 20 30 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.265 $Y=1.315
+ $X2=1.265 $Y2=1.075
r77 15 30 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=1.217 $Y=0.943
+ $X2=1.217 $Y2=1.075
r78 15 17 22.7444 $w=2.63e-07 $l=5.23e-07 $layer=LI1_cond $X=1.217 $Y=0.943
+ $X2=1.217 $Y2=0.42
r79 13 39 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.915 $Y=2.045
+ $X2=1.915 $Y2=1.605
r80 9 38 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.915 $Y=0.865
+ $X2=1.915 $Y2=1.275
r81 2 43 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.835 $X2=1.18 $Y2=2.91
r82 2 41 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.835 $X2=1.18 $Y2=2
r83 1 17 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.04
+ $Y=0.235 $X2=1.18 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_315_131# 1 2 9 13 15 17 19 20 22 29
+ 33
c64 19 0 1.89796e-19 $X=2.245 $Y=1.605
r65 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.44
+ $X2=2.365 $Y2=1.605
r66 33 35 48.8344 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.365 $Y=1.44
+ $X2=2.365 $Y2=1.26
r67 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.365
+ $Y=1.44 $X2=2.365 $Y2=1.44
r68 30 32 19.9828 $w=2.32e-07 $l=3.8e-07 $layer=LI1_cond $X=2.305 $Y=1.06
+ $X2=2.305 $Y2=1.44
r69 27 29 6.24272 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=2.06
+ $X2=1.865 $Y2=2.06
r70 22 24 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=1.682 $Y=0.865
+ $X2=1.682 $Y2=1.06
r71 19 32 9.57122 $w=2.32e-07 $l=1.92678e-07 $layer=LI1_cond $X=2.245 $Y=1.605
+ $X2=2.305 $Y2=1.44
r72 19 20 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.245 $Y=1.605
+ $X2=2.245 $Y2=1.895
r73 17 20 7.24806 $w=2.65e-07 $l=1.69245e-07 $layer=LI1_cond $X=2.16 $Y=2.027
+ $X2=2.245 $Y2=1.895
r74 17 29 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=2.16 $Y=2.027
+ $X2=1.865 $Y2=2.027
r75 16 24 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.83 $Y=1.06
+ $X2=1.682 $Y2=1.06
r76 15 30 2.55969 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.16 $Y=1.06
+ $X2=2.305 $Y2=1.06
r77 15 16 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.16 $Y=1.06
+ $X2=1.83 $Y2=1.06
r78 13 36 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.405 $Y=2.465
+ $X2=2.405 $Y2=1.605
r79 9 35 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=2.405 $Y=0.655
+ $X2=2.405 $Y2=1.26
r80 2 27 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.835 $X2=1.7 $Y2=2.06
r81 1 22 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.575
+ $Y=0.655 $X2=1.7 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_496_47# 1 2 9 13 17 20 25 26 28 29
+ 30 31 41
c65 26 0 1.89796e-19 $X=3.265 $Y=1.44
r66 41 43 36.1629 $w=2.88e-07 $l=9.1e-07 $layer=LI1_cond $X=2.645 $Y=2 $X2=2.645
+ $Y2=2.91
r67 28 41 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=2.645 $Y=1.98
+ $X2=2.645 $Y2=2
r68 28 29 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.645 $Y=1.98
+ $X2=2.645 $Y2=1.835
r69 26 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.265 $Y=1.44
+ $X2=3.265 $Y2=1.605
r70 26 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.265 $Y=1.44
+ $X2=3.265 $Y2=1.275
r71 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.265
+ $Y=1.44 $X2=3.265 $Y2=1.44
r72 23 31 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=1.46
+ $X2=2.705 $Y2=1.46
r73 23 25 18.8762 $w=2.88e-07 $l=4.75e-07 $layer=LI1_cond $X=2.79 $Y=1.46
+ $X2=3.265 $Y2=1.46
r74 21 31 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.705 $Y=1.605
+ $X2=2.705 $Y2=1.46
r75 21 29 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.705 $Y=1.605
+ $X2=2.705 $Y2=1.835
r76 20 31 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.705 $Y=1.315
+ $X2=2.705 $Y2=1.46
r77 20 30 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.705 $Y=1.315
+ $X2=2.705 $Y2=1.075
r78 15 30 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=2.657 $Y=0.943
+ $X2=2.657 $Y2=1.075
r79 15 17 22.7444 $w=2.63e-07 $l=5.23e-07 $layer=LI1_cond $X=2.657 $Y=0.943
+ $X2=2.657 $Y2=0.42
r80 13 39 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.355 $Y=2.045
+ $X2=3.355 $Y2=1.605
r81 9 38 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.355 $Y=0.865
+ $X2=3.355 $Y2=1.275
r82 2 43 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2.91
r83 2 41 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2
r84 1 17 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.48
+ $Y=0.235 $X2=2.62 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_603_131# 1 2 9 13 15 17 19 20 22 29
+ 33
r64 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.805 $Y=1.44
+ $X2=3.805 $Y2=1.605
r65 33 35 48.8344 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.805 $Y=1.44
+ $X2=3.805 $Y2=1.26
r66 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.805
+ $Y=1.44 $X2=3.805 $Y2=1.44
r67 30 32 19.9828 $w=2.32e-07 $l=3.8e-07 $layer=LI1_cond $X=3.745 $Y=1.06
+ $X2=3.745 $Y2=1.44
r68 27 29 6.24272 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=2.06
+ $X2=3.305 $Y2=2.06
r69 22 24 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=3.122 $Y=0.865
+ $X2=3.122 $Y2=1.06
r70 19 32 9.57122 $w=2.32e-07 $l=1.92678e-07 $layer=LI1_cond $X=3.685 $Y=1.605
+ $X2=3.745 $Y2=1.44
r71 19 20 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.685 $Y=1.605
+ $X2=3.685 $Y2=1.895
r72 17 20 7.24806 $w=2.65e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.6 $Y=2.027
+ $X2=3.685 $Y2=1.895
r73 17 29 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=3.6 $Y=2.027
+ $X2=3.305 $Y2=2.027
r74 16 24 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.27 $Y=1.06
+ $X2=3.122 $Y2=1.06
r75 15 30 2.55969 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.6 $Y=1.06
+ $X2=3.745 $Y2=1.06
r76 15 16 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.6 $Y=1.06 $X2=3.27
+ $Y2=1.06
r77 13 36 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.845 $Y=2.465
+ $X2=3.845 $Y2=1.605
r78 9 35 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=3.845 $Y=0.655
+ $X2=3.845 $Y2=1.26
r79 2 27 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=1.835 $X2=3.14 $Y2=2.06
r80 1 22 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.655 $X2=3.14 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%VPWR 1 2 3 12 16 20 22 24 29 34 41 42
+ 45 48 51 58
r51 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 39 51 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.76 $Y=3.33
+ $X2=3.612 $Y2=3.33
r56 39 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.76 $Y=3.33 $X2=4.08
+ $Y2=3.33
r57 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 35 48 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.172 $Y2=3.33
r60 35 37 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=2.32 $Y=3.33 $X2=3.12
+ $Y2=3.33
r61 34 51 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.612 $Y2=3.33
r62 34 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 33 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.92 $Y2=3.33
r64 33 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 30 45 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.88 $Y=3.33
+ $X2=0.732 $Y2=3.33
r67 30 32 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.88 $Y=3.33 $X2=1.68
+ $Y2=3.33
r68 29 48 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.172 $Y2=3.33
r69 29 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 24 45 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.732 $Y2=3.33
r73 24 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 22 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 22 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.92 $Y2=3.33
r76 22 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 18 51 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.612 $Y=3.245
+ $X2=3.612 $Y2=3.33
r78 18 20 29.2994 $w=2.93e-07 $l=7.5e-07 $layer=LI1_cond $X=3.612 $Y=3.245
+ $X2=3.612 $Y2=2.495
r79 14 48 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.172 $Y=3.245
+ $X2=2.172 $Y2=3.33
r80 14 16 29.2994 $w=2.93e-07 $l=7.5e-07 $layer=LI1_cond $X=2.172 $Y=3.245
+ $X2=2.172 $Y2=2.495
r81 10 45 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.732 $Y=3.245
+ $X2=0.732 $Y2=3.33
r82 10 12 29.2994 $w=2.93e-07 $l=7.5e-07 $layer=LI1_cond $X=0.732 $Y=3.245
+ $X2=0.732 $Y2=2.495
r83 3 20 300 $w=1.7e-07 $l=7.53392e-07 $layer=licon1_PDIFF $count=2 $X=3.43
+ $Y=1.835 $X2=3.63 $Y2=2.495
r84 2 16 300 $w=1.7e-07 $l=7.53392e-07 $layer=licon1_PDIFF $count=2 $X=1.99
+ $Y=1.835 $X2=2.19 $Y2=2.495
r85 1 12 300 $w=1.7e-07 $l=7.53392e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.75 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%X 1 2 9 13 14 15 16 21 23 27 31
c47 27 0 4.97211e-20 $X=3.84 $Y=2.405
r48 27 31 1.20842 $w=1.7e-07 $l=1.255e-06 $layer=MET1_cond $X=3.84 $Y=2.405
+ $X2=2.585 $Y2=2.405
r49 21 25 35.5499 $w=2.93e-07 $l=9.1e-07 $layer=LI1_cond $X=4.087 $Y=2 $X2=4.087
+ $Y2=2.91
r50 21 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.06 $Y=2.035
+ $X2=4.06 $Y2=2.035
r51 16 27 0.0563365 $w=1.7e-07 $l=1.82e-07 $layer=MET1_cond $X=4.022 $Y=2.405
+ $X2=3.84 $Y2=2.405
r52 16 23 0.0840525 $w=7.3e-07 $l=2.85e-07 $layer=MET1_cond $X=4.022 $Y=2.32
+ $X2=4.022 $Y2=2.035
r53 16 31 0.178133 $w=1.7e-07 $l=1.85e-07 $layer=MET1_cond $X=2.4 $Y=2.405
+ $X2=2.585 $Y2=2.405
r54 14 15 48.1662 $w=1.73e-07 $l=7.6e-07 $layer=LI1_cond $X=4.147 $Y=1.835
+ $X2=4.147 $Y2=1.075
r55 13 21 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=4.087 $Y=1.982
+ $X2=4.087 $Y2=2
r56 13 14 7.6342 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=4.087 $Y=1.982
+ $X2=4.087 $Y2=1.835
r57 7 15 7.18642 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.1 $Y=0.94 $X2=4.1
+ $Y2=1.075
r58 7 9 22.1952 $w=2.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.1 $Y=0.94 $X2=4.1
+ $Y2=0.42
r59 2 25 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.835 $X2=4.06 $Y2=2.91
r60 2 21 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.835 $X2=4.06 $Y2=2
r61 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.92
+ $Y=0.235 $X2=4.06 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%VGND 1 2 3 12 16 20 22 24 29 34 41 42
+ 45 48 51 58
r61 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r62 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r63 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r64 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r65 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.63
+ $Y2=0
r66 39 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=4.08
+ $Y2=0
r67 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r68 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r69 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.19
+ $Y2=0
r70 35 37 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=3.12
+ $Y2=0
r71 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.63
+ $Y2=0
r72 34 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.12
+ $Y2=0
r73 33 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.92
+ $Y2=0
r74 33 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r75 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r76 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r77 30 32 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.68
+ $Y2=0
r78 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.19
+ $Y2=0
r79 29 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.68
+ $Y2=0
r80 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r81 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r82 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r83 24 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r84 22 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r85 22 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.92
+ $Y2=0
r86 22 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r87 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=0.085
+ $X2=3.63 $Y2=0
r88 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.63 $Y=0.085
+ $X2=3.63 $Y2=0.38
r89 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0
r90 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0.38
r91 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r92 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.38
r93 3 20 91 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_NDIFF $count=2 $X=3.43
+ $Y=0.655 $X2=3.63 $Y2=0.38
r94 2 16 91 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.655 $X2=2.19 $Y2=0.38
r95 1 12 91 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.655 $X2=0.75 $Y2=0.38
.ends

