* File: sky130_fd_sc_lp__a2bb2o_2.pxi.spice
* Created: Fri Aug 28 09:55:52 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2O_2%B1 N_B1_M1001_g N_B1_c_79_n N_B1_M1013_g B1 B1 B1
+ N_B1_c_81_n PM_SKY130_FD_SC_LP__A2BB2O_2%B1
x_PM_SKY130_FD_SC_LP__A2BB2O_2%B2 N_B2_M1008_g N_B2_M1010_g N_B2_c_107_n
+ N_B2_c_108_n B2 B2 B2 N_B2_c_105_n PM_SKY130_FD_SC_LP__A2BB2O_2%B2
x_PM_SKY130_FD_SC_LP__A2BB2O_2%A_260_341# N_A_260_341#_M1006_d
+ N_A_260_341#_M1005_s N_A_260_341#_M1002_g N_A_260_341#_M1011_g
+ N_A_260_341#_c_138_n N_A_260_341#_c_144_n N_A_260_341#_c_145_n
+ N_A_260_341#_c_139_n N_A_260_341#_c_140_n N_A_260_341#_c_153_p
+ N_A_260_341#_c_186_p N_A_260_341#_c_168_p N_A_260_341#_c_141_n
+ PM_SKY130_FD_SC_LP__A2BB2O_2%A_260_341#
x_PM_SKY130_FD_SC_LP__A2BB2O_2%A2_N N_A2_N_c_197_n N_A2_N_M1006_g N_A2_N_c_198_n
+ N_A2_N_M1005_g A2_N PM_SKY130_FD_SC_LP__A2BB2O_2%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2O_2%A1_N N_A1_N_M1009_g N_A1_N_M1007_g A1_N A1_N A1_N
+ N_A1_N_c_233_n PM_SKY130_FD_SC_LP__A2BB2O_2%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2O_2%A_218_131# N_A_218_131#_M1010_d
+ N_A_218_131#_M1002_d N_A_218_131#_M1004_g N_A_218_131#_M1000_g
+ N_A_218_131#_M1012_g N_A_218_131#_M1003_g N_A_218_131#_c_269_n
+ N_A_218_131#_c_275_n N_A_218_131#_c_276_n N_A_218_131#_c_277_n
+ N_A_218_131#_c_278_n N_A_218_131#_c_281_n N_A_218_131#_c_270_n
+ N_A_218_131#_c_271_n PM_SKY130_FD_SC_LP__A2BB2O_2%A_218_131#
x_PM_SKY130_FD_SC_LP__A2BB2O_2%A_27_481# N_A_27_481#_M1001_s N_A_27_481#_M1008_d
+ N_A_27_481#_c_358_n N_A_27_481#_c_359_n N_A_27_481#_c_360_n
+ PM_SKY130_FD_SC_LP__A2BB2O_2%A_27_481#
x_PM_SKY130_FD_SC_LP__A2BB2O_2%VPWR N_VPWR_M1001_d N_VPWR_M1009_d N_VPWR_M1003_d
+ N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n VPWR
+ N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n N_VPWR_c_389_n
+ N_VPWR_c_380_n PM_SKY130_FD_SC_LP__A2BB2O_2%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2O_2%X N_X_M1004_d N_X_M1000_s N_X_c_436_n N_X_c_433_n
+ X X X X N_X_c_434_n PM_SKY130_FD_SC_LP__A2BB2O_2%X
x_PM_SKY130_FD_SC_LP__A2BB2O_2%VGND N_VGND_M1013_s N_VGND_M1011_d N_VGND_M1007_d
+ N_VGND_M1012_s N_VGND_c_460_n N_VGND_c_461_n N_VGND_c_462_n N_VGND_c_463_n
+ N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n N_VGND_c_467_n N_VGND_c_468_n
+ VGND N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n
+ PM_SKY130_FD_SC_LP__A2BB2O_2%VGND
cc_1 VNB N_B1_M1001_g 0.00757866f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.725
cc_2 VNB N_B1_c_79_n 0.0211898f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.185
cc_3 VNB B1 0.0270415f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_c_81_n 0.0606548f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.35
cc_5 VNB N_B2_M1010_g 0.0346853f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.865
cc_6 VNB B2 0.0105905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B2_c_105_n 0.0122299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_260_341#_c_138_n 0.0224386f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.35
cc_9 VNB N_A_260_341#_c_139_n 0.00203992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_260_341#_c_140_n 0.0252903f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_11 VNB N_A_260_341#_c_141_n 0.0201641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_N_c_197_n 0.0204787f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.515
cc_13 VNB N_A2_N_c_198_n 0.0324413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_N_M1005_g 0.00795304f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.865
cc_15 VNB A2_N 0.00305282f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_A1_N_M1009_g 0.00494815f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.725
cc_17 VNB N_A1_N_M1007_g 0.019916f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.865
cc_18 VNB A1_N 0.00896326f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_A1_N_c_233_n 0.034195f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.35
cc_20 VNB N_A_218_131#_M1004_g 0.0274136f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_A_218_131#_M1012_g 0.0329094f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.35
cc_22 VNB N_A_218_131#_c_269_n 0.0093172f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.035
cc_23 VNB N_A_218_131#_c_270_n 0.00394643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_218_131#_c_271_n 0.0460144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_380_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_433_n 0.00460221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_434_n 0.00196553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_460_n 0.0485332f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.35
cc_29 VNB N_VGND_c_461_n 0.0326685f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.295
cc_30 VNB N_VGND_c_462_n 0.00484226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_463_n 0.0126166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_464_n 0.0143681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_465_n 0.0108943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_466_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_467_n 0.0309449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_468_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_469_n 0.0307367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_470_n 0.021138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_471_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_472_n 0.277486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_B1_M1001_g 0.0582542f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.725
cc_42 VPB B1 0.0330056f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_43 VPB N_B2_M1008_g 0.0211926f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.725
cc_44 VPB N_B2_c_107_n 0.0208011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_B2_c_108_n 0.0151579f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB B2 0.00641022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B2_c_105_n 0.00353249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_260_341#_M1002_g 0.0440668f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_49 VPB N_A_260_341#_c_138_n 0.00428159f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.35
cc_50 VPB N_A_260_341#_c_144_n 0.0240335f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.35
cc_51 VPB N_A_260_341#_c_145_n 0.0140136f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.295
cc_52 VPB N_A2_N_M1005_g 0.0226863f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=0.865
cc_53 VPB N_A1_N_M1009_g 0.0207063f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.725
cc_54 VPB A1_N 0.00252726f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_55 VPB N_A_218_131#_M1000_g 0.0208771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_218_131#_M1003_g 0.0252934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_218_131#_c_269_n 0.00256371f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.035
cc_58 VPB N_A_218_131#_c_275_n 0.0215695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_218_131#_c_276_n 0.00826133f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_218_131#_c_277_n 0.0115535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_218_131#_c_278_n 0.00136033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_218_131#_c_270_n 4.01188e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_218_131#_c_271_n 0.00546596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_27_481#_c_358_n 0.00929831f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_65 VPB N_A_27_481#_c_359_n 0.00215435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_27_481#_c_360_n 0.0317479f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.35
cc_67 VPB N_VPWR_c_381_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_382_n 0.0205687f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.35
cc_69 VPB N_VPWR_c_383_n 0.0125908f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.185
cc_70 VPB N_VPWR_c_384_n 0.0143681f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_385_n 0.0162474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_386_n 0.0582215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_387_n 0.0176396f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_388_n 0.00497946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_389_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_380_n 0.0713552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_X_c_434_n 0.00104585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 N_B1_M1001_g N_B2_M1008_g 0.0225661f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_79 N_B1_c_79_n N_B2_M1010_g 0.0488106f $X=0.655 $Y=1.185 $X2=0 $Y2=0
cc_80 N_B1_c_81_n N_B2_M1010_g 0.00556075f $X=0.475 $Y=1.35 $X2=0 $Y2=0
cc_81 B1 B2 0.0854577f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_B1_c_81_n B2 0.0238685f $X=0.475 $Y=1.35 $X2=0 $Y2=0
cc_83 N_B1_M1001_g N_B2_c_105_n 0.0390353f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_84 N_B1_c_79_n N_A_218_131#_c_281_n 8.9899e-19 $X=0.655 $Y=1.185 $X2=0 $Y2=0
cc_85 N_B1_M1001_g N_A_27_481#_c_358_n 0.0147164f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_86 B1 N_A_27_481#_c_358_n 0.00241154f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_87 N_B1_M1001_g N_A_27_481#_c_360_n 6.86005e-19 $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_88 B1 N_A_27_481#_c_360_n 0.0253259f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_B1_M1001_g N_VPWR_c_381_n 0.00723307f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_90 N_B1_M1001_g N_VPWR_c_385_n 0.00516525f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_91 N_B1_M1001_g N_VPWR_c_380_n 0.00550061f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_92 N_B1_c_79_n N_VGND_c_460_n 0.011853f $X=0.655 $Y=1.185 $X2=0 $Y2=0
cc_93 B1 N_VGND_c_460_n 0.010382f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B1_c_81_n N_VGND_c_460_n 0.00807585f $X=0.475 $Y=1.35 $X2=0 $Y2=0
cc_95 N_B1_c_79_n N_VGND_c_469_n 0.00332367f $X=0.655 $Y=1.185 $X2=0 $Y2=0
cc_96 N_B1_c_79_n N_VGND_c_472_n 0.00387424f $X=0.655 $Y=1.185 $X2=0 $Y2=0
cc_97 N_B2_M1008_g N_A_260_341#_M1002_g 0.0147267f $X=0.945 $Y=2.725 $X2=0 $Y2=0
cc_98 N_B2_c_107_n N_A_260_341#_M1002_g 0.0157138f $X=0.925 $Y=2.05 $X2=0 $Y2=0
cc_99 B2 N_A_260_341#_c_144_n 4.61115e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B2_c_105_n N_A_260_341#_c_144_n 0.0157138f $X=0.925 $Y=1.71 $X2=0 $Y2=0
cc_101 N_B2_c_105_n N_A_260_341#_c_140_n 0.0155021f $X=0.925 $Y=1.71 $X2=0 $Y2=0
cc_102 N_B2_M1010_g N_A_260_341#_c_141_n 0.0155021f $X=1.015 $Y=0.865 $X2=0
+ $Y2=0
cc_103 N_B2_M1010_g N_A_218_131#_c_269_n 0.00918679f $X=1.015 $Y=0.865 $X2=0
+ $Y2=0
cc_104 B2 N_A_218_131#_c_269_n 0.0661375f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B2_c_107_n N_A_218_131#_c_277_n 0.00115121f $X=0.925 $Y=2.05 $X2=0
+ $Y2=0
cc_106 B2 N_A_218_131#_c_277_n 0.0142716f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_107 N_B2_M1010_g N_A_218_131#_c_281_n 0.00678415f $X=1.015 $Y=0.865 $X2=0
+ $Y2=0
cc_108 N_B2_M1008_g N_A_27_481#_c_358_n 0.00992994f $X=0.945 $Y=2.725 $X2=0
+ $Y2=0
cc_109 N_B2_c_108_n N_A_27_481#_c_358_n 0.00388425f $X=0.925 $Y=2.215 $X2=0
+ $Y2=0
cc_110 B2 N_A_27_481#_c_358_n 0.0365262f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B2_M1008_g N_VPWR_c_381_n 0.00686186f $X=0.945 $Y=2.725 $X2=0 $Y2=0
cc_112 N_B2_M1008_g N_VPWR_c_386_n 0.00516525f $X=0.945 $Y=2.725 $X2=0 $Y2=0
cc_113 N_B2_M1008_g N_VPWR_c_380_n 0.0048725f $X=0.945 $Y=2.725 $X2=0 $Y2=0
cc_114 N_B2_M1010_g N_VGND_c_460_n 0.0017007f $X=1.015 $Y=0.865 $X2=0 $Y2=0
cc_115 B2 N_VGND_c_460_n 0.00258185f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_116 N_B2_M1010_g N_VGND_c_469_n 0.00385857f $X=1.015 $Y=0.865 $X2=0 $Y2=0
cc_117 N_B2_M1010_g N_VGND_c_472_n 0.0046122f $X=1.015 $Y=0.865 $X2=0 $Y2=0
cc_118 N_A_260_341#_c_139_n N_A2_N_c_197_n 0.00291412f $X=1.625 $Y=1.35
+ $X2=-0.19 $Y2=-0.245
cc_119 N_A_260_341#_c_153_p N_A2_N_c_197_n 0.0114145f $X=2.415 $Y=0.945
+ $X2=-0.19 $Y2=-0.245
cc_120 N_A_260_341#_c_141_n N_A2_N_c_197_n 0.00802982f $X=1.58 $Y=1.185
+ $X2=-0.19 $Y2=-0.245
cc_121 N_A_260_341#_c_145_n N_A2_N_c_198_n 0.00502377f $X=1.66 $Y=1.685 $X2=0
+ $Y2=0
cc_122 N_A_260_341#_c_139_n N_A2_N_c_198_n 9.76598e-19 $X=1.625 $Y=1.35 $X2=0
+ $Y2=0
cc_123 N_A_260_341#_c_140_n N_A2_N_c_198_n 0.0170668f $X=1.625 $Y=1.35 $X2=0
+ $Y2=0
cc_124 N_A_260_341#_c_153_p N_A2_N_c_198_n 0.0041066f $X=2.415 $Y=0.945 $X2=0
+ $Y2=0
cc_125 N_A_260_341#_c_138_n N_A2_N_M1005_g 0.0085324f $X=1.545 $Y=1.705 $X2=0
+ $Y2=0
cc_126 N_A_260_341#_c_145_n N_A2_N_M1005_g 0.0087335f $X=1.66 $Y=1.685 $X2=0
+ $Y2=0
cc_127 N_A_260_341#_c_139_n N_A2_N_M1005_g 9.33144e-19 $X=1.625 $Y=1.35 $X2=0
+ $Y2=0
cc_128 N_A_260_341#_c_145_n A2_N 0.0189686f $X=1.66 $Y=1.685 $X2=0 $Y2=0
cc_129 N_A_260_341#_c_139_n A2_N 0.0177975f $X=1.625 $Y=1.35 $X2=0 $Y2=0
cc_130 N_A_260_341#_c_140_n A2_N 0.00147595f $X=1.625 $Y=1.35 $X2=0 $Y2=0
cc_131 N_A_260_341#_c_153_p A2_N 0.0264625f $X=2.415 $Y=0.945 $X2=0 $Y2=0
cc_132 N_A_260_341#_c_145_n N_A1_N_M1009_g 4.22224e-19 $X=1.66 $Y=1.685 $X2=0
+ $Y2=0
cc_133 N_A_260_341#_c_145_n A1_N 0.0250367f $X=1.66 $Y=1.685 $X2=0 $Y2=0
cc_134 N_A_260_341#_c_168_p A1_N 0.00565531f $X=2.52 $Y=0.865 $X2=0 $Y2=0
cc_135 N_A_260_341#_M1002_g N_A_218_131#_c_269_n 0.00521521f $X=1.375 $Y=2.725
+ $X2=0 $Y2=0
cc_136 N_A_260_341#_c_144_n N_A_218_131#_c_269_n 0.00505292f $X=1.545 $Y=1.855
+ $X2=0 $Y2=0
cc_137 N_A_260_341#_c_145_n N_A_218_131#_c_269_n 0.0186378f $X=1.66 $Y=1.685
+ $X2=0 $Y2=0
cc_138 N_A_260_341#_c_139_n N_A_218_131#_c_269_n 0.045302f $X=1.625 $Y=1.35
+ $X2=0 $Y2=0
cc_139 N_A_260_341#_c_141_n N_A_218_131#_c_269_n 0.00559755f $X=1.58 $Y=1.185
+ $X2=0 $Y2=0
cc_140 N_A_260_341#_M1002_g N_A_218_131#_c_275_n 2.3258e-19 $X=1.375 $Y=2.725
+ $X2=0 $Y2=0
cc_141 N_A_260_341#_M1005_s N_A_218_131#_c_276_n 0.00725406f $X=1.985 $Y=1.835
+ $X2=0 $Y2=0
cc_142 N_A_260_341#_c_145_n N_A_218_131#_c_276_n 0.0287673f $X=1.66 $Y=1.685
+ $X2=0 $Y2=0
cc_143 N_A_260_341#_M1002_g N_A_218_131#_c_277_n 0.0257082f $X=1.375 $Y=2.725
+ $X2=0 $Y2=0
cc_144 N_A_260_341#_c_144_n N_A_218_131#_c_277_n 0.00540273f $X=1.545 $Y=1.855
+ $X2=0 $Y2=0
cc_145 N_A_260_341#_c_145_n N_A_218_131#_c_277_n 0.0217402f $X=1.66 $Y=1.685
+ $X2=0 $Y2=0
cc_146 N_A_260_341#_M1002_g N_A_27_481#_c_359_n 3.44761e-19 $X=1.375 $Y=2.725
+ $X2=0 $Y2=0
cc_147 N_A_260_341#_M1002_g N_VPWR_c_381_n 8.58002e-19 $X=1.375 $Y=2.725 $X2=0
+ $Y2=0
cc_148 N_A_260_341#_M1002_g N_VPWR_c_386_n 0.0053602f $X=1.375 $Y=2.725 $X2=0
+ $Y2=0
cc_149 N_A_260_341#_M1002_g N_VPWR_c_380_n 0.0113452f $X=1.375 $Y=2.725 $X2=0
+ $Y2=0
cc_150 N_A_260_341#_c_139_n N_VGND_M1011_d 6.76331e-19 $X=1.625 $Y=1.35 $X2=0
+ $Y2=0
cc_151 N_A_260_341#_c_153_p N_VGND_M1011_d 0.0139049f $X=2.415 $Y=0.945 $X2=0
+ $Y2=0
cc_152 N_A_260_341#_c_186_p N_VGND_M1011_d 0.00453446f $X=1.79 $Y=0.945 $X2=0
+ $Y2=0
cc_153 N_A_260_341#_c_140_n N_VGND_c_461_n 7.02585e-19 $X=1.625 $Y=1.35 $X2=0
+ $Y2=0
cc_154 N_A_260_341#_c_153_p N_VGND_c_461_n 0.0113023f $X=2.415 $Y=0.945 $X2=0
+ $Y2=0
cc_155 N_A_260_341#_c_186_p N_VGND_c_461_n 0.0150495f $X=1.79 $Y=0.945 $X2=0
+ $Y2=0
cc_156 N_A_260_341#_c_141_n N_VGND_c_461_n 0.00471351f $X=1.58 $Y=1.185 $X2=0
+ $Y2=0
cc_157 N_A_260_341#_c_168_p N_VGND_c_467_n 0.00299849f $X=2.52 $Y=0.865 $X2=0
+ $Y2=0
cc_158 N_A_260_341#_c_141_n N_VGND_c_469_n 0.00399858f $X=1.58 $Y=1.185 $X2=0
+ $Y2=0
cc_159 N_A_260_341#_c_153_p N_VGND_c_472_n 0.0161077f $X=2.415 $Y=0.945 $X2=0
+ $Y2=0
cc_160 N_A_260_341#_c_186_p N_VGND_c_472_n 0.0037891f $X=1.79 $Y=0.945 $X2=0
+ $Y2=0
cc_161 N_A_260_341#_c_168_p N_VGND_c_472_n 0.00581712f $X=2.52 $Y=0.865 $X2=0
+ $Y2=0
cc_162 N_A_260_341#_c_141_n N_VGND_c_472_n 0.0046122f $X=1.58 $Y=1.185 $X2=0
+ $Y2=0
cc_163 N_A2_N_M1005_g N_A1_N_M1009_g 0.0380668f $X=2.325 $Y=2.155 $X2=0 $Y2=0
cc_164 N_A2_N_c_197_n N_A1_N_M1007_g 0.0144665f $X=2.305 $Y=1.185 $X2=0 $Y2=0
cc_165 N_A2_N_c_198_n A1_N 0.0102418f $X=2.325 $Y=1.515 $X2=0 $Y2=0
cc_166 A2_N A1_N 0.0180858f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_167 N_A2_N_c_198_n N_A1_N_c_233_n 0.0466958f $X=2.325 $Y=1.515 $X2=0 $Y2=0
cc_168 A2_N N_A1_N_c_233_n 2.43808e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_169 N_A2_N_M1005_g N_A_218_131#_c_275_n 0.00349785f $X=2.325 $Y=2.155 $X2=0
+ $Y2=0
cc_170 N_A2_N_M1005_g N_A_218_131#_c_276_n 0.0169655f $X=2.325 $Y=2.155 $X2=0
+ $Y2=0
cc_171 N_A2_N_M1005_g N_A_218_131#_c_277_n 0.00346748f $X=2.325 $Y=2.155 $X2=0
+ $Y2=0
cc_172 N_A2_N_M1005_g N_VPWR_c_386_n 0.00312414f $X=2.325 $Y=2.155 $X2=0 $Y2=0
cc_173 N_A2_N_M1005_g N_VPWR_c_380_n 0.00410284f $X=2.325 $Y=2.155 $X2=0 $Y2=0
cc_174 N_A2_N_c_197_n N_VGND_c_461_n 0.00365985f $X=2.305 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A2_N_c_197_n N_VGND_c_467_n 0.00399858f $X=2.305 $Y=1.185 $X2=0 $Y2=0
cc_176 N_A2_N_c_197_n N_VGND_c_472_n 0.0046122f $X=2.305 $Y=1.185 $X2=0 $Y2=0
cc_177 N_A1_N_M1007_g N_A_218_131#_M1004_g 0.0147074f $X=2.735 $Y=0.865 $X2=0
+ $Y2=0
cc_178 A1_N N_A_218_131#_M1004_g 7.16385e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A1_N_c_233_n N_A_218_131#_M1004_g 0.00677471f $X=2.775 $Y=1.375 $X2=0
+ $Y2=0
cc_180 N_A1_N_M1009_g N_A_218_131#_M1000_g 0.0235087f $X=2.685 $Y=2.155 $X2=0
+ $Y2=0
cc_181 A1_N N_A_218_131#_M1000_g 0.00127576f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A1_N_M1009_g N_A_218_131#_c_276_n 0.011771f $X=2.685 $Y=2.155 $X2=0
+ $Y2=0
cc_183 A1_N N_A_218_131#_c_276_n 0.0162264f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A1_N_M1009_g N_A_218_131#_c_278_n 0.0045203f $X=2.685 $Y=2.155 $X2=0
+ $Y2=0
cc_185 A1_N N_A_218_131#_c_278_n 0.0355815f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A1_N_M1009_g N_A_218_131#_c_270_n 3.83794e-19 $X=2.685 $Y=2.155 $X2=0
+ $Y2=0
cc_187 A1_N N_A_218_131#_c_270_n 0.0267653f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A1_N_c_233_n N_A_218_131#_c_270_n 0.00130385f $X=2.775 $Y=1.375 $X2=0
+ $Y2=0
cc_189 N_A1_N_M1009_g N_A_218_131#_c_271_n 0.00375564f $X=2.685 $Y=2.155 $X2=0
+ $Y2=0
cc_190 A1_N N_A_218_131#_c_271_n 5.50855e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_191 N_A1_N_c_233_n N_A_218_131#_c_271_n 0.0124456f $X=2.775 $Y=1.375 $X2=0
+ $Y2=0
cc_192 A1_N N_VPWR_M1009_d 0.00324007f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_193 N_A1_N_M1009_g N_VPWR_c_386_n 0.00312414f $X=2.685 $Y=2.155 $X2=0 $Y2=0
cc_194 N_A1_N_M1009_g N_VPWR_c_380_n 0.00410284f $X=2.685 $Y=2.155 $X2=0 $Y2=0
cc_195 A1_N A_480_367# 0.00308225f $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_196 N_A1_N_M1007_g N_VGND_c_462_n 0.00571568f $X=2.735 $Y=0.865 $X2=0 $Y2=0
cc_197 N_A1_N_M1007_g N_VGND_c_467_n 0.00399858f $X=2.735 $Y=0.865 $X2=0 $Y2=0
cc_198 N_A1_N_M1007_g N_VGND_c_472_n 0.0046122f $X=2.735 $Y=0.865 $X2=0 $Y2=0
cc_199 N_A_218_131#_c_277_n N_A_27_481#_c_358_n 0.0111019f $X=1.755 $Y=2.385
+ $X2=0 $Y2=0
cc_200 N_A_218_131#_c_275_n N_A_27_481#_c_359_n 7.23808e-19 $X=1.59 $Y=2.55
+ $X2=0 $Y2=0
cc_201 N_A_218_131#_c_276_n N_VPWR_M1009_d 0.0115623f $X=3.04 $Y=2.385 $X2=0
+ $Y2=0
cc_202 N_A_218_131#_c_278_n N_VPWR_M1009_d 0.00470965f $X=3.125 $Y=2.3 $X2=0
+ $Y2=0
cc_203 N_A_218_131#_M1000_g N_VPWR_c_382_n 0.013421f $X=3.26 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_A_218_131#_M1003_g N_VPWR_c_382_n 0.00123574f $X=3.69 $Y=2.465 $X2=0
+ $Y2=0
cc_205 N_A_218_131#_c_276_n N_VPWR_c_382_n 0.0223659f $X=3.04 $Y=2.385 $X2=0
+ $Y2=0
cc_206 N_A_218_131#_M1003_g N_VPWR_c_384_n 0.0293047f $X=3.69 $Y=2.465 $X2=0
+ $Y2=0
cc_207 N_A_218_131#_c_275_n N_VPWR_c_386_n 0.0186437f $X=1.59 $Y=2.55 $X2=0
+ $Y2=0
cc_208 N_A_218_131#_M1000_g N_VPWR_c_387_n 0.00486043f $X=3.26 $Y=2.465 $X2=0
+ $Y2=0
cc_209 N_A_218_131#_M1003_g N_VPWR_c_387_n 0.00397139f $X=3.69 $Y=2.465 $X2=0
+ $Y2=0
cc_210 N_A_218_131#_M1000_g N_VPWR_c_380_n 0.00824727f $X=3.26 $Y=2.465 $X2=0
+ $Y2=0
cc_211 N_A_218_131#_M1003_g N_VPWR_c_380_n 0.00744526f $X=3.69 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_A_218_131#_c_275_n N_VPWR_c_380_n 0.0112813f $X=1.59 $Y=2.55 $X2=0
+ $Y2=0
cc_213 N_A_218_131#_c_276_n N_VPWR_c_380_n 0.0382965f $X=3.04 $Y=2.385 $X2=0
+ $Y2=0
cc_214 N_A_218_131#_c_276_n A_480_367# 0.00543298f $X=3.04 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A_218_131#_M1012_g N_X_c_436_n 0.0134355f $X=3.69 $Y=0.655 $X2=0 $Y2=0
cc_216 N_A_218_131#_M1004_g N_X_c_433_n 0.00107084f $X=3.26 $Y=0.655 $X2=0 $Y2=0
cc_217 N_A_218_131#_M1012_g N_X_c_433_n 0.00336016f $X=3.69 $Y=0.655 $X2=0 $Y2=0
cc_218 N_A_218_131#_c_270_n N_X_c_433_n 0.00186252f $X=3.315 $Y=1.505 $X2=0
+ $Y2=0
cc_219 N_A_218_131#_c_271_n N_X_c_433_n 0.00410025f $X=3.69 $Y=1.505 $X2=0 $Y2=0
cc_220 N_A_218_131#_M1003_g X 0.00309304f $X=3.69 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A_218_131#_c_270_n X 0.00102806f $X=3.315 $Y=1.505 $X2=0 $Y2=0
cc_222 N_A_218_131#_c_271_n X 0.0043964f $X=3.69 $Y=1.505 $X2=0 $Y2=0
cc_223 N_A_218_131#_M1003_g X 0.0200677f $X=3.69 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_218_131#_M1004_g N_X_c_434_n 0.00372485f $X=3.26 $Y=0.655 $X2=0 $Y2=0
cc_225 N_A_218_131#_M1000_g N_X_c_434_n 8.73872e-19 $X=3.26 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A_218_131#_M1012_g N_X_c_434_n 0.013532f $X=3.69 $Y=0.655 $X2=0 $Y2=0
cc_227 N_A_218_131#_M1003_g N_X_c_434_n 0.00863355f $X=3.69 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A_218_131#_c_278_n N_X_c_434_n 0.00530127f $X=3.125 $Y=2.3 $X2=0 $Y2=0
cc_229 N_A_218_131#_c_270_n N_X_c_434_n 0.023711f $X=3.315 $Y=1.505 $X2=0 $Y2=0
cc_230 N_A_218_131#_c_271_n N_X_c_434_n 0.0217574f $X=3.69 $Y=1.505 $X2=0 $Y2=0
cc_231 N_A_218_131#_c_281_n N_VGND_c_460_n 0.0109469f $X=1.23 $Y=0.85 $X2=0
+ $Y2=0
cc_232 N_A_218_131#_M1004_g N_VGND_c_462_n 0.00442088f $X=3.26 $Y=0.655 $X2=0
+ $Y2=0
cc_233 N_A_218_131#_c_270_n N_VGND_c_462_n 0.00378395f $X=3.315 $Y=1.505 $X2=0
+ $Y2=0
cc_234 N_A_218_131#_M1012_g N_VGND_c_464_n 0.020996f $X=3.69 $Y=0.655 $X2=0
+ $Y2=0
cc_235 N_A_218_131#_c_281_n N_VGND_c_469_n 0.00408946f $X=1.23 $Y=0.85 $X2=0
+ $Y2=0
cc_236 N_A_218_131#_M1004_g N_VGND_c_470_n 0.00585385f $X=3.26 $Y=0.655 $X2=0
+ $Y2=0
cc_237 N_A_218_131#_M1012_g N_VGND_c_470_n 0.00397139f $X=3.69 $Y=0.655 $X2=0
+ $Y2=0
cc_238 N_A_218_131#_M1004_g N_VGND_c_472_n 0.0119451f $X=3.26 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_A_218_131#_M1012_g N_VGND_c_472_n 0.00744526f $X=3.69 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_218_131#_c_281_n N_VGND_c_472_n 0.0084104f $X=1.23 $Y=0.85 $X2=0
+ $Y2=0
cc_241 N_A_27_481#_c_358_n N_VPWR_M1001_d 0.00214775f $X=1.055 $Y=2.47 $X2=-0.19
+ $Y2=1.655
cc_242 N_A_27_481#_c_358_n N_VPWR_c_381_n 0.0168196f $X=1.055 $Y=2.47 $X2=0
+ $Y2=0
cc_243 N_A_27_481#_c_359_n N_VPWR_c_381_n 0.0129072f $X=1.16 $Y=2.56 $X2=0 $Y2=0
cc_244 N_A_27_481#_c_360_n N_VPWR_c_381_n 0.0136686f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_245 N_A_27_481#_c_360_n N_VPWR_c_385_n 0.0192334f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_246 N_A_27_481#_c_359_n N_VPWR_c_386_n 0.0157099f $X=1.16 $Y=2.56 $X2=0 $Y2=0
cc_247 N_A_27_481#_c_358_n N_VPWR_c_380_n 0.0121906f $X=1.055 $Y=2.47 $X2=0
+ $Y2=0
cc_248 N_A_27_481#_c_359_n N_VPWR_c_380_n 0.00901551f $X=1.16 $Y=2.56 $X2=0
+ $Y2=0
cc_249 N_A_27_481#_c_360_n N_VPWR_c_380_n 0.0104232f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_250 N_VPWR_c_380_n N_X_M1000_s 0.00380103f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_251 N_VPWR_c_387_n X 0.0225053f $X=3.91 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_c_380_n X 0.0132777f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_253 N_VPWR_c_384_n N_X_c_434_n 0.0952254f $X=3.995 $Y=1.98 $X2=0 $Y2=0
cc_254 N_X_c_436_n N_VGND_c_464_n 0.0635511f $X=3.475 $Y=0.42 $X2=0 $Y2=0
cc_255 N_X_c_436_n N_VGND_c_470_n 0.0228601f $X=3.475 $Y=0.42 $X2=0 $Y2=0
cc_256 N_X_M1004_d N_VGND_c_472_n 0.00345315f $X=3.335 $Y=0.235 $X2=0 $Y2=0
cc_257 N_X_c_436_n N_VGND_c_472_n 0.0136664f $X=3.475 $Y=0.42 $X2=0 $Y2=0
