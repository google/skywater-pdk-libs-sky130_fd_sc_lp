* File: sky130_fd_sc_lp__xor2_1.pex.spice
* Created: Fri Aug 28 11:36:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XOR2_1%B 1 3 6 10 14 16 17 18 22 23 25 26 39 46
r88 39 46 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=0.27 $Y=1.725 $X2=0.27
+ $Y2=1.665
r89 34 36 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.8 $Y=1.51 $X2=1.82
+ $Y2=1.51
r90 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.46 $X2=0.29 $Y2=1.46
r91 26 39 2.55307 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=1.81 $X2=0.27
+ $Y2=1.725
r92 26 46 0.404912 $w=3.68e-07 $l=1.3e-08 $layer=LI1_cond $X=0.27 $Y=1.652
+ $X2=0.27 $Y2=1.665
r93 26 32 5.98024 $w=3.68e-07 $l=1.92e-07 $layer=LI1_cond $X=0.27 $Y=1.652
+ $X2=0.27 $Y2=1.46
r94 25 32 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.46
r95 23 36 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.03 $Y=1.51
+ $X2=1.82 $Y2=1.51
r96 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.51 $X2=2.03 $Y2=1.51
r97 20 22 13.2475 $w=1.78e-07 $l=2.15e-07 $layer=LI1_cond $X=2.025 $Y=1.725
+ $X2=2.025 $Y2=1.51
r98 19 26 5.55669 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.455 $Y=1.81
+ $X2=0.27 $Y2=1.81
r99 18 20 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.935 $Y=1.81
+ $X2=2.025 $Y2=1.725
r100 18 19 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=1.935 $Y=1.81
+ $X2=0.455 $Y2=1.81
r101 16 31 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.475 $Y=1.46
+ $X2=0.29 $Y2=1.46
r102 16 17 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.46
+ $X2=0.55 $Y2=1.46
r103 12 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=1.675
+ $X2=1.82 $Y2=1.51
r104 12 14 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.82 $Y=1.675
+ $X2=1.82 $Y2=2.465
r105 8 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=1.345
+ $X2=1.8 $Y2=1.51
r106 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.8 $Y=1.345 $X2=1.8
+ $Y2=0.765
r107 4 17 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.625
+ $X2=0.55 $Y2=1.46
r108 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.55 $Y=1.625
+ $X2=0.55 $Y2=2.465
r109 1 17 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.295
+ $X2=0.55 $Y2=1.46
r110 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.55 $Y=1.295
+ $X2=0.55 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_1%A 3 5 7 10 12 14 15 16 17 28
c51 28 0 1.28341e-19 $X=1.41 $Y=1.46
c52 10 0 3.61764e-20 $X=1.39 $Y=2.465
r53 27 28 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.39 $Y=1.46 $X2=1.41
+ $Y2=1.46
r54 25 27 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.34 $Y=1.46 $X2=1.39
+ $Y2=1.46
r55 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.34
+ $Y=1.46 $X2=1.34 $Y2=1.46
r56 23 25 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=0.98 $Y=1.46
+ $X2=1.34 $Y2=1.46
r57 21 23 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.94 $Y=1.46 $X2=0.98
+ $Y2=1.46
r58 17 26 11.3574 $w=3.43e-07 $l=3.4e-07 $layer=LI1_cond $X=1.68 $Y=1.382
+ $X2=1.34 $Y2=1.382
r59 16 26 4.67658 $w=3.43e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.382
+ $X2=1.34 $Y2=1.382
r60 15 16 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.382 $X2=1.2
+ $Y2=1.382
r61 12 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.46
r62 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=0.765
r63 8 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.625
+ $X2=1.39 $Y2=1.46
r64 8 10 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.39 $Y=1.625
+ $X2=1.39 $Y2=2.465
r65 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.295
+ $X2=0.98 $Y2=1.46
r66 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.98 $Y=1.295 $X2=0.98
+ $Y2=0.765
r67 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.625
+ $X2=0.94 $Y2=1.46
r68 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.94 $Y=1.625 $X2=0.94
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_1%A_42_367# 1 2 7 9 11 14 16 18 20 22 24 26 29
+ 30 31 32 35 37 42 48 49 52
c108 22 0 1.28341e-19 $X=0.73 $Y=0.87
r109 51 52 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=1.46
+ $X2=2.81 $Y2=1.46
r110 49 51 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.07 $Y=1.46
+ $X2=2.885 $Y2=1.46
r111 48 50 3.35395 $w=2.91e-07 $l=8e-08 $layer=LI1_cond $X=3.07 $Y=1.427
+ $X2=3.15 $Y2=1.427
r112 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.46 $X2=3.07 $Y2=1.46
r113 42 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.025 $Y=2.15
+ $X2=2.025 $Y2=2.32
r114 36 50 3.88217 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=3.15 $Y=1.625
+ $X2=3.15 $Y2=1.427
r115 36 37 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.15 $Y=1.625
+ $X2=3.15 $Y2=2.235
r116 35 48 15.0928 $w=2.91e-07 $l=4.47795e-07 $layer=LI1_cond $X=2.71 $Y=1.23
+ $X2=3.07 $Y2=1.427
r117 34 35 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=2.71 $Y=0.425
+ $X2=2.71 $Y2=1.23
r118 33 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=2.32
+ $X2=2.025 $Y2=2.32
r119 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.065 $Y=2.32
+ $X2=3.15 $Y2=2.235
r120 32 33 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.065 $Y=2.32
+ $X2=2.11 $Y2=2.32
r121 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.625 $Y=0.34
+ $X2=2.71 $Y2=0.425
r122 30 31 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.625 $Y=0.34
+ $X2=1.87 $Y2=0.34
r123 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.785 $Y=0.425
+ $X2=1.87 $Y2=0.34
r124 28 29 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.785 $Y=0.425
+ $X2=1.785 $Y2=0.87
r125 27 41 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.86 $Y=0.955
+ $X2=0.73 $Y2=0.955
r126 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.7 $Y=0.955
+ $X2=1.785 $Y2=0.87
r127 26 27 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.7 $Y=0.955
+ $X2=0.86 $Y2=0.955
r128 22 41 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.87
+ $X2=0.73 $Y2=0.955
r129 22 24 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=0.87
+ $X2=0.73 $Y2=0.5
r130 21 39 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.5 $Y=2.15
+ $X2=0.335 $Y2=2.15
r131 20 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.15
+ $X2=2.025 $Y2=2.15
r132 20 21 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.94 $Y=2.15
+ $X2=0.5 $Y2=2.15
r133 16 39 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.335 $Y=2.235
+ $X2=0.335 $Y2=2.15
r134 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.335 $Y=2.235
+ $X2=0.335 $Y2=2.91
r135 12 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.625
+ $X2=2.885 $Y2=1.46
r136 12 14 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.885 $Y=1.625
+ $X2=2.885 $Y2=2.465
r137 11 52 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.605 $Y=1.37
+ $X2=2.81 $Y2=1.37
r138 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.53 $Y=1.295
+ $X2=2.605 $Y2=1.37
r139 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.53 $Y=1.295
+ $X2=2.53 $Y2=0.765
r140 2 39 400 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=1.835 $X2=0.335 $Y2=2.15
r141 2 18 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=1.835 $X2=0.335 $Y2=2.91
r142 1 41 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.345 $X2=0.765 $Y2=0.955
r143 1 24 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.345 $X2=0.765 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_1%VPWR 1 2 9 12 13 14 20 26 27 30
r48 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 30 33 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.13 $Y=3.02 $X2=2.13
+ $Y2=3.33
r50 27 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 24 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.13 $Y2=3.33
r53 24 26 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 20 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=2.13 $Y2=3.33
r55 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 14 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 14 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 14 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 12 17 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=0.72
+ $Y2=3.33
r61 12 13 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.13
+ $Y2=3.33
r62 11 22 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 11 13 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.27 $Y=3.33 $X2=1.13
+ $Y2=3.33
r64 7 13 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=3.245
+ $X2=1.13 $Y2=3.33
r65 7 9 27.7821 $w=2.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.13 $Y=3.245
+ $X2=1.13 $Y2=2.57
r66 2 30 600 $w=1.7e-07 $l=1.29719e-06 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.835 $X2=2.13 $Y2=3.02
r67 1 9 300 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=2 $X=1.015
+ $Y=1.835 $X2=1.155 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_1%A_293_367# 1 2 7 10 14
c30 7 0 3.61764e-20 $X=2.935 $Y=2.66
r31 14 17 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.1 $Y=2.66 $X2=3.1
+ $Y2=2.76
r32 10 12 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.605 $Y=2.49
+ $X2=1.605 $Y2=2.66
r33 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=2.66
+ $X2=1.605 $Y2=2.66
r34 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=2.66 $X2=3.1
+ $Y2=2.66
r35 7 8 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=2.935 $Y=2.66
+ $X2=1.77 $Y2=2.66
r36 2 17 600 $w=1.7e-07 $l=9.92535e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.76
r37 1 10 300 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=2 $X=1.465
+ $Y=1.835 $X2=1.605 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_1%X 1 2 8 10 13
r32 13 19 1.11585 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.817 $X2=2.67
+ $Y2=1.817
r33 10 12 17.5996 $w=4.13e-07 $l=4.85e-07 $layer=LI1_cond $X=2.247 $Y=0.68
+ $X2=2.247 $Y2=1.165
r34 8 13 10.0427 $w=3.28e-07 $l=3.73617e-07 $layer=LI1_cond $X=2.37 $Y=1.57
+ $X2=2.64 $Y2=1.817
r35 8 12 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.37 $Y=1.57
+ $X2=2.37 $Y2=1.165
r36 2 19 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.835 $X2=2.67 $Y2=1.96
r37 1 10 91 $w=1.7e-07 $l=4.7199e-07 $layer=licon1_NDIFF $count=2 $X=1.875
+ $Y=0.345 $X2=2.205 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_1%VGND 1 2 3 10 12 16 18 20 22 24 29 41 45
r44 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 36 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r48 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r49 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 30 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=0 $X2=1.195
+ $Y2=0
r51 30 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.36 $Y=0 $X2=1.68
+ $Y2=0
r52 29 44 3.97515 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=3.162
+ $Y2=0
r53 29 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.64
+ $Y2=0
r54 28 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r55 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r56 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 25 38 4.0276 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r58 25 27 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r59 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.195
+ $Y2=0
r60 24 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r61 22 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r62 22 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r63 22 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 18 44 3.16801 $w=2.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=3.09 $Y=0.085
+ $X2=3.162 $Y2=0
r65 18 20 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=3.09 $Y=0.085
+ $X2=3.09 $Y2=0.49
r66 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0
r67 14 16 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0.575
r68 10 38 3.18462 $w=2.6e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.215 $Y2=0
r69 10 12 17.9515 $w=2.58e-07 $l=4.05e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.3 $Y2=0.49
r70 3 20 91 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_NDIFF $count=2 $X=2.605
+ $Y=0.345 $X2=3.05 $Y2=0.49
r71 2 16 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=1.055
+ $Y=0.345 $X2=1.195 $Y2=0.575
r72 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.345 $X2=0.335 $Y2=0.49
.ends

