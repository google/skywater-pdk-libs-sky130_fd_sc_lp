* File: sky130_fd_sc_lp__xor2_4.pex.spice
* Created: Fri Aug 28 11:36:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XOR2_4%A 3 7 11 15 19 23 27 30 34 38 42 46 50 54 58
+ 62 64 72 76 79 83 84 87 88 91 93 100 103 105 122
c250 76 0 1.71326e-19 $X=7.49 $Y=1.44
c251 3 0 1.414e-19 $X=0.475 $Y=0.655
r252 121 122 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.555 $Y=1.44
+ $X2=7.625 $Y2=1.44
r253 118 119 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.125 $Y=1.44
+ $X2=7.195 $Y2=1.44
r254 116 118 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=6.81 $Y=1.44
+ $X2=7.125 $Y2=1.44
r255 116 117 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.81
+ $Y=1.44 $X2=6.81 $Y2=1.44
r256 114 116 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.765 $Y=1.44
+ $X2=6.81 $Y2=1.44
r257 113 114 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.695 $Y=1.44
+ $X2=6.765 $Y2=1.44
r258 112 117 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=6.47 $Y=1.367
+ $X2=6.81 $Y2=1.367
r259 111 113 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=6.47 $Y=1.44
+ $X2=6.695 $Y2=1.44
r260 111 112 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.47
+ $Y=1.44 $X2=6.47 $Y2=1.44
r261 109 111 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.335 $Y=1.44
+ $X2=6.47 $Y2=1.44
r262 107 109 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.265 $Y=1.44
+ $X2=6.335 $Y2=1.44
r263 103 106 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.35
+ $X2=3.505 $Y2=1.515
r264 103 105 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.35
+ $X2=3.505 $Y2=1.185
r265 93 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.295
+ $X2=6.48 $Y2=1.295
r266 92 103 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.505
+ $Y=1.35 $X2=3.505 $Y2=1.35
r267 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=1.295
+ $X2=3.6 $Y2=1.295
r268 88 91 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=1.295
+ $X2=3.6 $Y2=1.295
r269 87 93 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.295
+ $X2=6.48 $Y2=1.295
r270 87 88 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=6.335 $Y=1.295
+ $X2=3.745 $Y2=1.295
r271 83 117 3.37133 $w=3.33e-07 $l=9.8e-08 $layer=LI1_cond $X=6.908 $Y=1.367
+ $X2=6.81 $Y2=1.367
r272 83 84 8.1966 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=6.908 $Y=1.367
+ $X2=7.075 $Y2=1.367
r273 77 121 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.49 $Y=1.44
+ $X2=7.555 $Y2=1.44
r274 77 119 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=7.49 $Y=1.44
+ $X2=7.195 $Y2=1.44
r275 76 84 25.5707 $w=1.78e-07 $l=4.15e-07 $layer=LI1_cond $X=7.49 $Y=1.445
+ $X2=7.075 $Y2=1.445
r276 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.49
+ $Y=1.44 $X2=7.49 $Y2=1.44
r277 73 79 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.555 $Y=1.16
+ $X2=1.407 $Y2=1.16
r278 72 92 4.50956 $w=3.43e-07 $l=1.35e-07 $layer=LI1_cond $X=3.512 $Y=1.16
+ $X2=3.512 $Y2=1.295
r279 72 73 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=3.34 $Y=1.16
+ $X2=1.555 $Y2=1.16
r280 71 100 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.245 $Y=1.44
+ $X2=1.335 $Y2=1.44
r281 71 98 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.245 $Y=1.44
+ $X2=0.905 $Y2=1.44
r282 70 71 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.245
+ $Y=1.44 $X2=1.245 $Y2=1.44
r283 67 98 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.565 $Y=1.44
+ $X2=0.905 $Y2=1.44
r284 67 95 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.565 $Y=1.44
+ $X2=0.475 $Y2=1.44
r285 66 70 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.565 $Y=1.4
+ $X2=1.245 $Y2=1.4
r286 66 67 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.565
+ $Y=1.44 $X2=0.565 $Y2=1.44
r287 64 79 9.37581 $w=2.93e-07 $l=2.4e-07 $layer=LI1_cond $X=1.407 $Y=1.4
+ $X2=1.407 $Y2=1.16
r288 64 70 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=1.26 $Y=1.4
+ $X2=1.245 $Y2=1.4
r289 60 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.625 $Y=1.605
+ $X2=7.625 $Y2=1.44
r290 60 62 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.625 $Y=1.605
+ $X2=7.625 $Y2=2.465
r291 56 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.555 $Y=1.275
+ $X2=7.555 $Y2=1.44
r292 56 58 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.555 $Y=1.275
+ $X2=7.555 $Y2=0.655
r293 52 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.195 $Y=1.605
+ $X2=7.195 $Y2=1.44
r294 52 54 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.195 $Y=1.605
+ $X2=7.195 $Y2=2.465
r295 48 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.125 $Y=1.275
+ $X2=7.125 $Y2=1.44
r296 48 50 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.125 $Y=1.275
+ $X2=7.125 $Y2=0.655
r297 44 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.765 $Y=1.605
+ $X2=6.765 $Y2=1.44
r298 44 46 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.765 $Y=1.605
+ $X2=6.765 $Y2=2.465
r299 40 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.275
+ $X2=6.695 $Y2=1.44
r300 40 42 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.695 $Y=1.275
+ $X2=6.695 $Y2=0.655
r301 36 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.605
+ $X2=6.335 $Y2=1.44
r302 36 38 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.335 $Y=1.605
+ $X2=6.335 $Y2=2.465
r303 32 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.265 $Y=1.275
+ $X2=6.265 $Y2=1.44
r304 32 34 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.265 $Y=1.275
+ $X2=6.265 $Y2=0.655
r305 30 106 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.515 $Y=2.465
+ $X2=3.515 $Y2=1.515
r306 27 105 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.485 $Y=0.655
+ $X2=3.485 $Y2=1.185
r307 21 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.605
+ $X2=1.335 $Y2=1.44
r308 21 23 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.335 $Y=1.605
+ $X2=1.335 $Y2=2.465
r309 17 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.275
+ $X2=1.335 $Y2=1.44
r310 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.335 $Y=1.275
+ $X2=1.335 $Y2=0.655
r311 13 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.605
+ $X2=0.905 $Y2=1.44
r312 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.905 $Y=1.605
+ $X2=0.905 $Y2=2.465
r313 9 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.275
+ $X2=0.905 $Y2=1.44
r314 9 11 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.905 $Y=1.275
+ $X2=0.905 $Y2=0.655
r315 5 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.605
+ $X2=0.475 $Y2=1.44
r316 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.475 $Y=1.605
+ $X2=0.475 $Y2=2.465
r317 1 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.275
+ $X2=0.475 $Y2=1.44
r318 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.475 $Y=1.275
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_4%B 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 70 71 73 74 79 93 94 113
c215 71 0 2.70796e-19 $X=9.435 $Y=1.44
r216 113 116 12.8421 $w=1.88e-07 $l=2.2e-07 $layer=LI1_cond $X=7.92 $Y=1.445
+ $X2=7.92 $Y2=1.665
r217 104 105 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=9.275 $Y=1.44
+ $X2=9.345 $Y2=1.44
r218 103 104 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=8.915 $Y=1.44
+ $X2=9.275 $Y2=1.44
r219 102 103 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.845 $Y=1.44
+ $X2=8.915 $Y2=1.44
r220 101 102 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=8.485 $Y=1.44
+ $X2=8.845 $Y2=1.44
r221 100 101 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.415 $Y=1.44
+ $X2=8.485 $Y2=1.44
r222 96 98 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.985 $Y=1.44
+ $X2=8.055 $Y2=1.44
r223 92 94 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.92 $Y=1.51
+ $X2=3.055 $Y2=1.51
r224 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.92
+ $Y=1.51 $X2=2.92 $Y2=1.51
r225 90 92 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.92 $Y2=1.51
r226 89 93 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.58 $Y=1.595
+ $X2=2.92 $Y2=1.595
r227 88 90 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=2.58 $Y=1.51
+ $X2=2.625 $Y2=1.51
r228 88 89 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.58
+ $Y=1.51 $X2=2.58 $Y2=1.51
r229 86 88 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.58 $Y2=1.51
r230 85 89 21.7684 $w=3.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.9 $Y=1.595
+ $X2=2.58 $Y2=1.595
r231 84 86 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=1.9 $Y=1.51
+ $X2=2.195 $Y2=1.51
r232 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.9
+ $Y=1.51 $X2=1.9 $Y2=1.51
r233 81 84 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.9 $Y2=1.51
r234 79 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.665
r235 76 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r236 74 76 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r237 73 79 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=1.665
+ $X2=7.92 $Y2=1.665
r238 73 74 6.17573 $w=1.4e-07 $l=4.99e-06 $layer=MET1_cond $X=7.775 $Y=1.665
+ $X2=2.785 $Y2=1.665
r239 71 105 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.435 $Y=1.44
+ $X2=9.345 $Y2=1.44
r240 70 71 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.435
+ $Y=1.44 $X2=9.435 $Y2=1.44
r241 68 100 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.075 $Y=1.44
+ $X2=8.415 $Y2=1.44
r242 68 98 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=8.075 $Y=1.44
+ $X2=8.055 $Y2=1.44
r243 67 70 83.798 $w=1.78e-07 $l=1.36e-06 $layer=LI1_cond $X=8.075 $Y=1.445
+ $X2=9.435 $Y2=1.445
r244 67 68 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.075
+ $Y=1.44 $X2=8.075 $Y2=1.44
r245 65 113 1.04402 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=8.015 $Y=1.445
+ $X2=7.92 $Y2=1.445
r246 65 67 3.69697 $w=1.78e-07 $l=6e-08 $layer=LI1_cond $X=8.015 $Y=1.445
+ $X2=8.075 $Y2=1.445
r247 61 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.345 $Y=1.605
+ $X2=9.345 $Y2=1.44
r248 61 63 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=9.345 $Y=1.605
+ $X2=9.345 $Y2=2.465
r249 57 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.275 $Y=1.275
+ $X2=9.275 $Y2=1.44
r250 57 59 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=9.275 $Y=1.275
+ $X2=9.275 $Y2=0.655
r251 53 103 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.915 $Y=1.605
+ $X2=8.915 $Y2=1.44
r252 53 55 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.915 $Y=1.605
+ $X2=8.915 $Y2=2.465
r253 49 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.845 $Y=1.275
+ $X2=8.845 $Y2=1.44
r254 49 51 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.845 $Y=1.275
+ $X2=8.845 $Y2=0.655
r255 45 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.485 $Y=1.605
+ $X2=8.485 $Y2=1.44
r256 45 47 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.485 $Y=1.605
+ $X2=8.485 $Y2=2.465
r257 41 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.415 $Y=1.275
+ $X2=8.415 $Y2=1.44
r258 41 43 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.415 $Y=1.275
+ $X2=8.415 $Y2=0.655
r259 37 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=1.605
+ $X2=8.055 $Y2=1.44
r260 37 39 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.055 $Y=1.605
+ $X2=8.055 $Y2=2.465
r261 33 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.985 $Y=1.275
+ $X2=7.985 $Y2=1.44
r262 33 35 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.985 $Y=1.275
+ $X2=7.985 $Y2=0.655
r263 29 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.675
+ $X2=3.055 $Y2=1.51
r264 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.055 $Y=1.675
+ $X2=3.055 $Y2=2.465
r265 25 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.345
+ $X2=3.055 $Y2=1.51
r266 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.055 $Y=1.345
+ $X2=3.055 $Y2=0.655
r267 21 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.675
+ $X2=2.625 $Y2=1.51
r268 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.625 $Y=1.675
+ $X2=2.625 $Y2=2.465
r269 17 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=1.51
r270 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=0.655
r271 13 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.675
+ $X2=2.195 $Y2=1.51
r272 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.195 $Y=1.675
+ $X2=2.195 $Y2=2.465
r273 9 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=1.51
r274 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=0.655
r275 5 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.675
+ $X2=1.765 $Y2=1.51
r276 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.765 $Y=1.675
+ $X2=1.765 $Y2=2.465
r277 1 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=1.51
r278 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_4%A_776_255# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 51 58 60 61 62 65 67 71 73 77 81 83 85 86 89 93 97 99 102 104 106 109 110
+ 111 112
c224 41 0 3.86629e-20 $X=4.845 $Y=0.655
c225 25 0 8.51568e-20 $X=3.985 $Y=0.655
r226 123 124 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.245 $Y=1.44
+ $X2=5.275 $Y2=1.44
r227 122 123 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=4.845 $Y=1.44
+ $X2=5.245 $Y2=1.44
r228 121 122 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.815 $Y=1.44
+ $X2=4.845 $Y2=1.44
r229 118 119 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.385 $Y=1.44
+ $X2=4.415 $Y2=1.44
r230 117 118 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=3.985 $Y=1.44
+ $X2=4.385 $Y2=1.44
r231 115 117 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.955 $Y=1.44
+ $X2=3.985 $Y2=1.44
r232 112 124 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.35 $Y=1.44
+ $X2=5.275 $Y2=1.44
r233 106 107 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=7.34 $Y=0.945
+ $X2=7.34 $Y2=1.1
r234 101 102 26.6342 $w=2.23e-07 $l=5.2e-07 $layer=LI1_cond $X=9.882 $Y=1.185
+ $X2=9.882 $Y2=1.705
r235 100 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.295 $Y=1.79
+ $X2=9.13 $Y2=1.79
r236 99 102 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=9.77 $Y=1.79
+ $X2=9.882 $Y2=1.705
r237 99 100 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=9.77 $Y=1.79
+ $X2=9.295 $Y2=1.79
r238 98 110 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.155 $Y=1.1
+ $X2=9.06 $Y2=1.1
r239 97 101 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=9.77 $Y=1.1
+ $X2=9.882 $Y2=1.185
r240 97 98 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=9.77 $Y=1.1
+ $X2=9.155 $Y2=1.1
r241 93 95 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=9.13 $Y=1.96
+ $X2=9.13 $Y2=2.65
r242 91 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.13 $Y=1.875
+ $X2=9.13 $Y2=1.79
r243 91 93 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=9.13 $Y=1.875
+ $X2=9.13 $Y2=1.96
r244 87 110 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.06 $Y=1.015
+ $X2=9.06 $Y2=1.1
r245 87 89 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=9.06 $Y=1.015
+ $X2=9.06 $Y2=0.42
r246 85 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.965 $Y=1.79
+ $X2=9.13 $Y2=1.79
r247 85 86 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.965 $Y=1.79
+ $X2=8.435 $Y2=1.79
r248 84 109 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.295 $Y=1.1
+ $X2=8.2 $Y2=1.1
r249 83 110 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.965 $Y=1.1
+ $X2=9.06 $Y2=1.1
r250 83 84 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.965 $Y=1.1
+ $X2=8.295 $Y2=1.1
r251 79 86 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.31 $Y=1.875
+ $X2=8.435 $Y2=1.79
r252 79 81 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=8.31 $Y=1.875
+ $X2=8.31 $Y2=1.96
r253 75 109 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.2 $Y=1.015
+ $X2=8.2 $Y2=1.1
r254 75 77 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=8.2 $Y=1.015
+ $X2=8.2 $Y2=0.42
r255 74 107 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.435 $Y=1.1 $X2=7.34
+ $Y2=1.1
r256 73 109 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.105 $Y=1.1
+ $X2=8.2 $Y2=1.1
r257 73 74 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.105 $Y=1.1
+ $X2=7.435 $Y2=1.1
r258 69 106 4.96172 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=7.34 $Y=0.86
+ $X2=7.34 $Y2=0.945
r259 69 71 25.6842 $w=1.88e-07 $l=4.4e-07 $layer=LI1_cond $X=7.34 $Y=0.86
+ $X2=7.34 $Y2=0.42
r260 68 104 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.575 $Y=0.945
+ $X2=6.48 $Y2=0.945
r261 67 106 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.245 $Y=0.945
+ $X2=7.34 $Y2=0.945
r262 67 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.245 $Y=0.945
+ $X2=6.575 $Y2=0.945
r263 63 104 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.48 $Y=0.86
+ $X2=6.48 $Y2=0.945
r264 63 65 25.6842 $w=1.88e-07 $l=4.4e-07 $layer=LI1_cond $X=6.48 $Y=0.86
+ $X2=6.48 $Y2=0.42
r265 61 104 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.385 $Y=0.945
+ $X2=6.48 $Y2=0.945
r266 61 62 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.385 $Y=0.945
+ $X2=6.135 $Y2=0.945
r267 59 62 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=5.98 $Y=1.03
+ $X2=6.135 $Y2=0.945
r268 59 60 12.0821 $w=3.08e-07 $l=3.25e-07 $layer=LI1_cond $X=5.98 $Y=1.03
+ $X2=5.98 $Y2=1.355
r269 58 112 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=5.74 $Y=1.44
+ $X2=5.35 $Y2=1.44
r270 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.74
+ $Y=1.44 $X2=5.74 $Y2=1.44
r271 54 121 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.61 $Y=1.44
+ $X2=4.815 $Y2=1.44
r272 54 119 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.61 $Y=1.44
+ $X2=4.415 $Y2=1.44
r273 53 57 69.6263 $w=1.78e-07 $l=1.13e-06 $layer=LI1_cond $X=4.61 $Y=1.445
+ $X2=5.74 $Y2=1.445
r274 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.61
+ $Y=1.44 $X2=4.61 $Y2=1.44
r275 51 60 7.45983 $w=1.8e-07 $l=1.94872e-07 $layer=LI1_cond $X=5.825 $Y=1.445
+ $X2=5.98 $Y2=1.355
r276 51 57 5.23737 $w=1.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.825 $Y=1.445
+ $X2=5.74 $Y2=1.445
r277 47 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.275 $Y=1.275
+ $X2=5.275 $Y2=1.44
r278 47 49 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.275 $Y=1.275
+ $X2=5.275 $Y2=0.655
r279 43 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=1.605
+ $X2=5.245 $Y2=1.44
r280 43 45 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.245 $Y=1.605
+ $X2=5.245 $Y2=2.465
r281 39 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.845 $Y=1.275
+ $X2=4.845 $Y2=1.44
r282 39 41 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=4.845 $Y=1.275
+ $X2=4.845 $Y2=0.655
r283 35 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=1.605
+ $X2=4.815 $Y2=1.44
r284 35 37 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.815 $Y=1.605
+ $X2=4.815 $Y2=2.465
r285 31 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.275
+ $X2=4.415 $Y2=1.44
r286 31 33 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=4.415 $Y=1.275
+ $X2=4.415 $Y2=0.655
r287 27 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.385 $Y=1.605
+ $X2=4.385 $Y2=1.44
r288 27 29 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.385 $Y=1.605
+ $X2=4.385 $Y2=2.465
r289 23 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.275
+ $X2=3.985 $Y2=1.44
r290 23 25 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.985 $Y=1.275
+ $X2=3.985 $Y2=0.655
r291 19 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.955 $Y=1.605
+ $X2=3.955 $Y2=1.44
r292 19 21 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.955 $Y=1.605
+ $X2=3.955 $Y2=2.465
r293 6 95 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=8.99
+ $Y=1.835 $X2=9.13 $Y2=2.65
r294 6 93 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=8.99
+ $Y=1.835 $X2=9.13 $Y2=1.96
r295 5 81 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=8.13
+ $Y=1.835 $X2=8.27 $Y2=1.96
r296 4 89 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.92
+ $Y=0.235 $X2=9.06 $Y2=0.42
r297 3 77 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.06
+ $Y=0.235 $X2=8.2 $Y2=0.42
r298 2 106 182 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_NDIFF $count=1 $X=7.2
+ $Y=0.235 $X2=7.34 $Y2=0.945
r299 2 71 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=7.2
+ $Y=0.235 $X2=7.34 $Y2=0.42
r300 1 104 182 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.235 $X2=6.48 $Y2=0.945
r301 1 65 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.235 $X2=6.48 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_4%A_27_367# 1 2 3 4 5 6 7 24 28 29 32 34 38 40
+ 44 46 48 49 50 54 56 58 65 67
r89 62 63 4.75232 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=2.03
+ $X2=1.125 $Y2=2.115
r90 61 62 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=1.125 $Y=1.98
+ $X2=1.125 $Y2=2.03
r91 58 61 11.0909 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=1.125 $Y=1.78
+ $X2=1.125 $Y2=1.98
r92 54 73 3.67598 $w=2.6e-07 $l=1.5e-07 $layer=LI1_cond $X=5.495 $Y=2.775
+ $X2=5.495 $Y2=2.925
r93 54 56 35.2382 $w=2.58e-07 $l=7.95e-07 $layer=LI1_cond $X=5.495 $Y=2.775
+ $X2=5.495 $Y2=1.98
r94 51 71 2.87089 $w=3e-07 $l=1e-07 $layer=LI1_cond $X=3.825 $Y=2.925 $X2=3.725
+ $Y2=2.925
r95 51 53 29.7714 $w=2.98e-07 $l=7.75e-07 $layer=LI1_cond $X=3.825 $Y=2.925
+ $X2=4.6 $Y2=2.925
r96 50 73 3.18585 $w=3e-07 $l=1.3e-07 $layer=LI1_cond $X=5.365 $Y=2.925
+ $X2=5.495 $Y2=2.925
r97 50 53 29.3873 $w=2.98e-07 $l=7.65e-07 $layer=LI1_cond $X=5.365 $Y=2.925
+ $X2=4.6 $Y2=2.925
r98 49 71 4.30634 $w=2e-07 $l=1.5e-07 $layer=LI1_cond $X=3.725 $Y=2.775
+ $X2=3.725 $Y2=2.925
r99 48 69 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=2.115
+ $X2=3.725 $Y2=2.03
r100 48 49 36.6 $w=1.98e-07 $l=6.6e-07 $layer=LI1_cond $X=3.725 $Y=2.115
+ $X2=3.725 $Y2=2.775
r101 47 67 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=2.95 $Y=2.03
+ $X2=2.847 $Y2=2.03
r102 46 69 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.625 $Y=2.03
+ $X2=3.725 $Y2=2.03
r103 46 47 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.625 $Y=2.03
+ $X2=2.95 $Y2=2.03
r104 42 67 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.847 $Y=2.115
+ $X2=2.847 $Y2=2.03
r105 42 44 19.7472 $w=2.03e-07 $l=3.65e-07 $layer=LI1_cond $X=2.847 $Y=2.115
+ $X2=2.847 $Y2=2.48
r106 41 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.075 $Y=2.03
+ $X2=1.98 $Y2=2.03
r107 40 67 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=2.745 $Y=2.03
+ $X2=2.847 $Y2=2.03
r108 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.745 $Y=2.03
+ $X2=2.075 $Y2=2.03
r109 36 65 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.115
+ $X2=1.98 $Y2=2.03
r110 36 38 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=1.98 $Y=2.115
+ $X2=1.98 $Y2=2.48
r111 35 62 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.225 $Y=2.03
+ $X2=1.125 $Y2=2.03
r112 34 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.885 $Y=2.03
+ $X2=1.98 $Y2=2.03
r113 34 35 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.885 $Y=2.03
+ $X2=1.225 $Y2=2.03
r114 32 63 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=1.12 $Y=2.44
+ $X2=1.12 $Y2=2.115
r115 28 58 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.025 $Y=1.78
+ $X2=1.125 $Y2=1.78
r116 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=1.78
+ $X2=0.355 $Y2=1.78
r117 24 26 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.225 $Y=1.98
+ $X2=0.225 $Y2=2.91
r118 22 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=1.865
+ $X2=0.355 $Y2=1.78
r119 22 24 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=0.225 $Y=1.865
+ $X2=0.225 $Y2=1.98
r120 7 73 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.32
+ $Y=1.835 $X2=5.46 $Y2=2.95
r121 7 56 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=5.32
+ $Y=1.835 $X2=5.46 $Y2=1.98
r122 6 53 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=1.835 $X2=4.6 $Y2=2.9
r123 5 71 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.59
+ $Y=1.835 $X2=3.73 $Y2=2.91
r124 5 69 300 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=2 $X=3.59
+ $Y=1.835 $X2=3.73 $Y2=2.11
r125 4 67 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.03
r126 4 44 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.48
r127 3 65 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.03
r128 3 38 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.48
r129 2 61 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=1.98
r130 2 32 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.44
r131 1 26 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r132 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_4%VPWR 1 2 3 4 5 6 21 27 31 33 37 41 45 48 49
+ 50 51 52 54 66 74 84 85 88 91 94 97
r139 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r140 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r141 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r142 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r143 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r144 82 85 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=9.84 $Y2=3.33
r145 82 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r146 81 84 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=9.84 $Y2=3.33
r147 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r148 79 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.575 $Y=3.33
+ $X2=7.41 $Y2=3.33
r149 79 81 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.575 $Y=3.33
+ $X2=7.92 $Y2=3.33
r150 78 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r151 78 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r152 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r153 75 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=3.33
+ $X2=6.55 $Y2=3.33
r154 75 77 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.715 $Y=3.33
+ $X2=6.96 $Y2=3.33
r155 74 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=3.33
+ $X2=7.41 $Y2=3.33
r156 74 77 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.245 $Y=3.33
+ $X2=6.96 $Y2=3.33
r157 73 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r158 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r159 70 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r160 69 72 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r161 69 70 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r162 67 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=3.33
+ $X2=3.285 $Y2=3.33
r163 67 69 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.45 $Y=3.33 $X2=3.6
+ $Y2=3.33
r164 66 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=3.33
+ $X2=6.55 $Y2=3.33
r165 66 72 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.385 $Y=3.33
+ $X2=6 $Y2=3.33
r166 65 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r167 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r168 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r169 62 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r170 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r171 59 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r172 59 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r173 57 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r174 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r175 54 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r176 54 56 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r177 52 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r178 52 70 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r179 50 64 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.16 $Y2=3.33
r180 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.41 $Y2=3.33
r181 48 61 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.2 $Y2=3.33
r182 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.55 $Y2=3.33
r183 47 64 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=2.16 $Y2=3.33
r184 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.55 $Y2=3.33
r185 43 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=3.245
+ $X2=7.41 $Y2=3.33
r186 43 45 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.41 $Y=3.245
+ $X2=7.41 $Y2=2.415
r187 39 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=3.245
+ $X2=6.55 $Y2=3.33
r188 39 41 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.55 $Y=3.245
+ $X2=6.55 $Y2=2.415
r189 35 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=3.245
+ $X2=3.285 $Y2=3.33
r190 35 37 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=3.285 $Y=3.245
+ $X2=3.285 $Y2=2.39
r191 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=3.33
+ $X2=2.41 $Y2=3.33
r192 33 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=3.285 $Y2=3.33
r193 33 34 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=2.575 $Y2=3.33
r194 29 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=3.245
+ $X2=2.41 $Y2=3.33
r195 29 31 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=2.41 $Y=3.245
+ $X2=2.41 $Y2=2.39
r196 25 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.55 $Y2=3.33
r197 25 27 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.55 $Y2=2.39
r198 21 24 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.69 $Y=2.12
+ $X2=0.69 $Y2=2.95
r199 19 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r200 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.95
r201 6 45 300 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_PDIFF $count=2 $X=7.27
+ $Y=1.835 $X2=7.41 $Y2=2.415
r202 5 41 300 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_PDIFF $count=2 $X=6.41
+ $Y=1.835 $X2=6.55 $Y2=2.415
r203 4 37 300 $w=1.7e-07 $l=6.27734e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=1.835 $X2=3.285 $Y2=2.39
r204 3 31 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.39
r205 2 27 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.39
r206 1 24 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.95
r207 1 21 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_4%X 1 2 3 4 5 6 19 26 28 31 33 35 37 41 43 49
+ 50 51 55
c83 33 0 8.51568e-20 $X=4.965 $Y=1.1
r84 51 55 3.49538 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=5.03 $Y=2.447
+ $X2=4.865 $Y2=2.447
r85 50 55 11.1586 $w=3.13e-07 $l=3.05e-07 $layer=LI1_cond $X=4.56 $Y=2.447
+ $X2=4.865 $Y2=2.447
r86 50 56 10.4269 $w=3.13e-07 $l=2.85e-07 $layer=LI1_cond $X=4.56 $Y=2.447
+ $X2=4.275 $Y2=2.447
r87 49 56 3.22764 $w=3.15e-07 $l=1.4e-07 $layer=LI1_cond $X=4.135 $Y=2.447
+ $X2=4.275 $Y2=2.447
r88 47 48 3.3328 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=1.1
+ $X2=4.145 $Y2=1.185
r89 46 47 6.53051 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=4.145 $Y=0.93
+ $X2=4.145 $Y2=1.1
r90 43 46 4.99392 $w=2.98e-07 $l=1.3e-07 $layer=LI1_cond $X=4.145 $Y=0.8
+ $X2=4.145 $Y2=0.93
r91 43 44 5.57628 $w=2.98e-07 $l=1.05e-07 $layer=LI1_cond $X=4.145 $Y=0.8
+ $X2=4.145 $Y2=0.695
r92 39 41 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=5.06 $Y=1.015
+ $X2=5.06 $Y2=0.42
r93 35 51 3.32591 $w=3.3e-07 $l=1.57e-07 $layer=LI1_cond $X=5.03 $Y=2.29
+ $X2=5.03 $Y2=2.447
r94 35 37 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.03 $Y=2.29
+ $X2=5.03 $Y2=1.96
r95 34 47 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.295 $Y=1.1 $X2=4.145
+ $Y2=1.1
r96 33 39 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.965 $Y=1.1
+ $X2=5.06 $Y2=1.015
r97 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.965 $Y=1.1
+ $X2=4.295 $Y2=1.1
r98 31 44 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=4.2 $Y=0.42 $X2=4.2
+ $Y2=0.695
r99 28 48 31.898 $w=2.78e-07 $l=7.75e-07 $layer=LI1_cond $X=4.135 $Y=1.96
+ $X2=4.135 $Y2=1.185
r100 26 49 3.61957 $w=2.8e-07 $l=1.57e-07 $layer=LI1_cond $X=4.135 $Y=2.29
+ $X2=4.135 $Y2=2.447
r101 26 28 13.5824 $w=2.78e-07 $l=3.3e-07 $layer=LI1_cond $X=4.135 $Y=2.29
+ $X2=4.135 $Y2=1.96
r102 21 24 45.4199 $w=2.08e-07 $l=8.6e-07 $layer=LI1_cond $X=1.98 $Y=0.8
+ $X2=2.84 $Y2=0.8
r103 19 43 2.82627 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=3.995 $Y=0.8
+ $X2=4.145 $Y2=0.8
r104 19 24 61 $w=2.08e-07 $l=1.155e-06 $layer=LI1_cond $X=3.995 $Y=0.8 $X2=2.84
+ $Y2=0.8
r105 6 37 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.89
+ $Y=1.835 $X2=5.03 $Y2=1.96
r106 5 49 600 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=1 $X=4.03
+ $Y=1.835 $X2=4.17 $Y2=2.44
r107 5 28 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.03
+ $Y=1.835 $X2=4.17 $Y2=1.96
r108 4 41 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.92
+ $Y=0.235 $X2=5.06 $Y2=0.42
r109 3 46 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.235 $X2=4.2 $Y2=0.93
r110 3 31 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.235 $X2=4.2 $Y2=0.42
r111 2 24 182 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.8
r112 1 21 182 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_4%A_1199_367# 1 2 3 4 5 18 22 23 26 28 31 34 38
+ 40 42 44 47 51
c60 28 0 9.94698e-20 $X=7.745 $Y=2.055
r61 42 53 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.595 $Y=2.905
+ $X2=9.595 $Y2=2.99
r62 42 44 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=9.595 $Y=2.905
+ $X2=9.595 $Y2=2.21
r63 41 51 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.795 $Y=2.99 $X2=8.7
+ $Y2=2.99
r64 40 53 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.465 $Y=2.99
+ $X2=9.595 $Y2=2.99
r65 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.465 $Y=2.99
+ $X2=8.795 $Y2=2.99
r66 36 51 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.7 $Y=2.905 $X2=8.7
+ $Y2=2.99
r67 36 38 40.5694 $w=1.88e-07 $l=6.95e-07 $layer=LI1_cond $X=8.7 $Y=2.905
+ $X2=8.7 $Y2=2.21
r68 35 49 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.935 $Y=2.99
+ $X2=7.84 $Y2=2.99
r69 34 51 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.605 $Y=2.99 $X2=8.7
+ $Y2=2.99
r70 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.605 $Y=2.99
+ $X2=7.935 $Y2=2.99
r71 31 49 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.84 $Y=2.905
+ $X2=7.84 $Y2=2.99
r72 31 33 40.5694 $w=1.88e-07 $l=6.95e-07 $layer=LI1_cond $X=7.84 $Y=2.905
+ $X2=7.84 $Y2=2.21
r73 30 33 4.08612 $w=1.88e-07 $l=7e-08 $layer=LI1_cond $X=7.84 $Y=2.14 $X2=7.84
+ $Y2=2.21
r74 29 47 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.075 $Y=2.055
+ $X2=6.98 $Y2=2.055
r75 28 30 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.745 $Y=2.055
+ $X2=7.84 $Y2=2.14
r76 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.745 $Y=2.055
+ $X2=7.075 $Y2=2.055
r77 24 47 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=2.14
+ $X2=6.98 $Y2=2.055
r78 24 26 44.9474 $w=1.88e-07 $l=7.7e-07 $layer=LI1_cond $X=6.98 $Y=2.14
+ $X2=6.98 $Y2=2.91
r79 22 47 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.885 $Y=2.055
+ $X2=6.98 $Y2=2.055
r80 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.885 $Y=2.055
+ $X2=6.215 $Y2=2.055
r81 18 20 30.5841 $w=2.58e-07 $l=6.9e-07 $layer=LI1_cond $X=6.085 $Y=2.22
+ $X2=6.085 $Y2=2.91
r82 16 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.085 $Y=2.14
+ $X2=6.215 $Y2=2.055
r83 16 18 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=6.085 $Y=2.14
+ $X2=6.085 $Y2=2.22
r84 5 53 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.42
+ $Y=1.835 $X2=9.56 $Y2=2.91
r85 5 44 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=9.42
+ $Y=1.835 $X2=9.56 $Y2=2.21
r86 4 51 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.56
+ $Y=1.835 $X2=8.7 $Y2=2.91
r87 4 38 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=8.56
+ $Y=1.835 $X2=8.7 $Y2=2.21
r88 3 49 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.7
+ $Y=1.835 $X2=7.84 $Y2=2.91
r89 3 33 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=7.7
+ $Y=1.835 $X2=7.84 $Y2=2.21
r90 2 47 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.835 $X2=6.98 $Y2=2.13
r91 2 26 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.835 $X2=6.98 $Y2=2.91
r92 1 20 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=5.995
+ $Y=1.835 $X2=6.12 $Y2=2.91
r93 1 18 400 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=1 $X=5.995
+ $Y=1.835 $X2=6.12 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_4%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 54 58 60 64 67 68 70 71 72 73 74 76 85 94 108 109 115 118 122 131 133 136
c172 46 0 3.86629e-20 $X=5.49 $Y=0.94
r173 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r174 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r175 130 131 11.2794 $w=7.73e-07 $l=1.65e-07 $layer=LI1_cond $X=6.05 $Y=0.302
+ $X2=6.215 $Y2=0.302
r176 127 130 0.771663 $w=7.73e-07 $l=5e-08 $layer=LI1_cond $X=6 $Y=0.302
+ $X2=6.05 $Y2=0.302
r177 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r178 125 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r179 124 127 7.40797 $w=7.73e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=0.302
+ $X2=6 $Y2=0.302
r180 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r181 121 124 0.462998 $w=7.73e-07 $l=3e-08 $layer=LI1_cond $X=5.49 $Y=0.302
+ $X2=5.52 $Y2=0.302
r182 121 122 11.2794 $w=7.73e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=0.302
+ $X2=5.325 $Y2=0.302
r183 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r184 115 116 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r185 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r186 109 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r187 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r188 106 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.655 $Y=0
+ $X2=9.49 $Y2=0
r189 106 108 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.655 $Y=0
+ $X2=9.84 $Y2=0
r190 105 137 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=9.36 $Y2=0
r191 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r192 102 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.4 $Y2=0
r193 102 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r194 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r195 99 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.075 $Y=0
+ $X2=6.91 $Y2=0
r196 99 101 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.075 $Y=0
+ $X2=7.44 $Y2=0
r197 98 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r198 98 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r199 97 131 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.48 $Y=0
+ $X2=6.215 $Y2=0
r200 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r201 94 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.91 $Y2=0
r202 94 97 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.48 $Y2=0
r203 92 122 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.04 $Y=0
+ $X2=5.325 $Y2=0
r204 90 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0
+ $X2=4.63 $Y2=0
r205 90 92 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=5.04
+ $Y2=0
r206 88 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r207 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r208 85 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.465 $Y=0
+ $X2=4.63 $Y2=0
r209 85 87 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.465 $Y=0
+ $X2=4.08 $Y2=0
r210 84 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r211 84 116 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=1.2
+ $Y2=0
r212 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r213 81 115 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.215 $Y=0 $X2=1.1
+ $Y2=0
r214 81 83 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=1.215 $Y=0
+ $X2=3.6 $Y2=0
r215 80 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r216 80 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r217 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r218 77 112 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r219 77 79 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r220 76 115 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.1
+ $Y2=0
r221 76 79 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0
+ $X2=0.72 $Y2=0
r222 74 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r223 74 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r224 74 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r225 72 104 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=8.465 $Y=0 $X2=8.4
+ $Y2=0
r226 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.465 $Y=0 $X2=8.63
+ $Y2=0
r227 70 101 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=0
+ $X2=7.44 $Y2=0
r228 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=0 $X2=7.77
+ $Y2=0
r229 69 104 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.935 $Y=0
+ $X2=8.4 $Y2=0
r230 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.935 $Y=0 $X2=7.77
+ $Y2=0
r231 67 83 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.605 $Y=0 $X2=3.6
+ $Y2=0
r232 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=0 $X2=3.77
+ $Y2=0
r233 66 87 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.935 $Y=0
+ $X2=4.08 $Y2=0
r234 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.935 $Y=0 $X2=3.77
+ $Y2=0
r235 62 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.49 $Y=0.085
+ $X2=9.49 $Y2=0
r236 62 64 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.49 $Y=0.085
+ $X2=9.49 $Y2=0.38
r237 61 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.63
+ $Y2=0
r238 60 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.325 $Y=0
+ $X2=9.49 $Y2=0
r239 60 61 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=9.325 $Y=0
+ $X2=8.795 $Y2=0
r240 56 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.63 $Y=0.085
+ $X2=8.63 $Y2=0
r241 56 58 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.63 $Y=0.085
+ $X2=8.63 $Y2=0.38
r242 52 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.77 $Y=0.085
+ $X2=7.77 $Y2=0
r243 52 54 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.77 $Y=0.085
+ $X2=7.77 $Y2=0.38
r244 48 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.91 $Y=0.085
+ $X2=6.91 $Y2=0
r245 48 50 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.91 $Y=0.085
+ $X2=6.91 $Y2=0.565
r246 44 121 5.76689 $w=3.3e-07 $l=3.88e-07 $layer=LI1_cond $X=5.49 $Y=0.69
+ $X2=5.49 $Y2=0.302
r247 44 46 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.49 $Y=0.69
+ $X2=5.49 $Y2=0.94
r248 40 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=0.085
+ $X2=4.63 $Y2=0
r249 40 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.63 $Y=0.085
+ $X2=4.63 $Y2=0.38
r250 36 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=0.085
+ $X2=3.77 $Y2=0
r251 36 38 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.77 $Y=0.085
+ $X2=3.77 $Y2=0.4
r252 32 115 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0
r253 32 34 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.4
r254 28 112 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r255 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r256 9 64 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.35
+ $Y=0.235 $X2=9.49 $Y2=0.38
r257 8 58 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.49
+ $Y=0.235 $X2=8.63 $Y2=0.38
r258 7 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.63
+ $Y=0.235 $X2=7.77 $Y2=0.38
r259 6 50 182 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_NDIFF $count=1 $X=6.77
+ $Y=0.235 $X2=6.91 $Y2=0.565
r260 5 130 182 $w=1.7e-07 $l=8.49117e-07 $layer=licon1_NDIFF $count=1 $X=5.35
+ $Y=0.235 $X2=6.05 $Y2=0.565
r261 5 121 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.35
+ $Y=0.235 $X2=5.49 $Y2=0.38
r262 5 46 182 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_NDIFF $count=1 $X=5.35
+ $Y=0.235 $X2=5.49 $Y2=0.94
r263 4 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.49
+ $Y=0.235 $X2=4.63 $Y2=0.38
r264 3 38 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.77 $Y2=0.4
r265 2 34 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.4
r266 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_4%A_110_47# 1 2 3 4 13 15 17 19 20 25
c46 13 0 1.414e-19 $X=0.705 $Y=0.735
r47 23 25 36.7074 $w=2.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.41 $Y=0.39
+ $X2=3.27 $Y2=0.39
r48 21 30 3.34549 $w=2.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.645 $Y=0.39
+ $X2=1.515 $Y2=0.39
r49 21 23 32.6526 $w=2.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.645 $Y=0.39
+ $X2=2.41 $Y2=0.39
r50 20 32 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.515 $Y=0.735
+ $X2=1.515 $Y2=0.82
r51 19 30 3.47416 $w=2.6e-07 $l=1.35e-07 $layer=LI1_cond $X=1.515 $Y=0.525
+ $X2=1.515 $Y2=0.39
r52 19 20 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.515 $Y=0.525
+ $X2=1.515 $Y2=0.735
r53 18 28 3.7077 $w=1.7e-07 $l=1.50167e-07 $layer=LI1_cond $X=0.815 $Y=0.82
+ $X2=0.705 $Y2=0.915
r54 17 32 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.385 $Y=0.82
+ $X2=1.515 $Y2=0.82
r55 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.385 $Y=0.82
+ $X2=0.815 $Y2=0.82
r56 13 28 3.25554 $w=2.2e-07 $l=1.8e-07 $layer=LI1_cond $X=0.705 $Y=0.735
+ $X2=0.705 $Y2=0.915
r57 13 15 16.5009 $w=2.18e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=0.735
+ $X2=0.705 $Y2=0.42
r58 4 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.38
r59 3 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.38
r60 2 32 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.74
r61 2 30 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.4
r62 1 28 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.93
r63 1 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

