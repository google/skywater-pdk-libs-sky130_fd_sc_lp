* File: sky130_fd_sc_lp__a21oi_2.pex.spice
* Created: Wed Sep  2 09:20:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21OI_2%A2 3 7 11 15 17 20 25 29 32
c70 32 0 8.34927e-20 $X=1.785 $Y=1.51
c71 20 0 8.8057e-20 $X=0.29 $Y=1.46
r72 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.51
+ $X2=1.785 $Y2=1.675
r73 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.51
+ $X2=1.785 $Y2=1.345
r74 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.785
+ $Y=1.51 $X2=1.785 $Y2=1.51
r75 25 39 1.15094 $w=3.18e-07 $l=3e-08 $layer=LI1_cond $X=1.697 $Y=1.665
+ $X2=1.697 $Y2=1.695
r76 25 33 5.94654 $w=3.18e-07 $l=1.55e-07 $layer=LI1_cond $X=1.697 $Y=1.665
+ $X2=1.697 $Y2=1.51
r77 21 29 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.29 $Y=1.46
+ $X2=0.475 $Y2=1.46
r78 20 23 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.29 $Y=1.46
+ $X2=0.29 $Y2=1.695
r79 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.46 $X2=0.29 $Y2=1.46
r80 18 23 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=1.695
+ $X2=0.29 $Y2=1.695
r81 17 39 4.06753 $w=1.8e-07 $l=1.72e-07 $layer=LI1_cond $X=1.525 $Y=1.695
+ $X2=1.697 $Y2=1.695
r82 17 18 65.9293 $w=1.78e-07 $l=1.07e-06 $layer=LI1_cond $X=1.525 $Y=1.695
+ $X2=0.455 $Y2=1.695
r83 15 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.805 $Y=2.465
+ $X2=1.805 $Y2=1.675
r84 11 34 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.765 $Y=0.655
+ $X2=1.765 $Y2=1.345
r85 5 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.625
+ $X2=0.475 $Y2=1.46
r86 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.475 $Y=1.625
+ $X2=0.475 $Y2=2.465
r87 1 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=1.46
r88 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_2%A1 1 3 6 8 10 13 15 16 24
c49 16 0 8.34927e-20 $X=1.2 $Y=1.295
c50 6 0 8.8057e-20 $X=0.905 $Y=2.465
r51 22 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=1.335 $Y2=1.35
r52 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.35 $X2=0.995 $Y2=1.35
r53 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.905 $Y=1.35
+ $X2=0.995 $Y2=1.35
r54 16 23 10.2718 $w=2.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.2 $Y=1.32
+ $X2=0.995 $Y2=1.32
r55 15 23 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=1.32
+ $X2=0.995 $Y2=1.32
r56 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.515
+ $X2=1.335 $Y2=1.35
r57 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.335 $Y=1.515
+ $X2=1.335 $Y2=2.465
r58 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.185
+ $X2=1.335 $Y2=1.35
r59 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.335 $Y=1.185
+ $X2=1.335 $Y2=0.655
r60 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.515
+ $X2=0.905 $Y2=1.35
r61 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.905 $Y=1.515
+ $X2=0.905 $Y2=2.465
r62 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=1.35
r63 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_2%B1 3 7 11 15 17 18 26
r49 24 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.325 $Y=1.51
+ $X2=2.665 $Y2=1.51
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.325
+ $Y=1.51 $X2=2.325 $Y2=1.51
r51 21 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.235 $Y=1.51
+ $X2=2.325 $Y2=1.51
r52 18 25 10.8364 $w=3.33e-07 $l=3.15e-07 $layer=LI1_cond $X=2.64 $Y=1.592
+ $X2=2.325 $Y2=1.592
r53 17 25 5.67621 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=2.325 $Y2=1.592
r54 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=1.675
+ $X2=2.665 $Y2=1.51
r55 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.665 $Y=1.675
+ $X2=2.665 $Y2=2.465
r56 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=1.345
+ $X2=2.665 $Y2=1.51
r57 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.665 $Y=1.345
+ $X2=2.665 $Y2=0.655
r58 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.675
+ $X2=2.235 $Y2=1.51
r59 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.235 $Y=1.675
+ $X2=2.235 $Y2=2.465
r60 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.345
+ $X2=2.235 $Y2=1.51
r61 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.235 $Y=1.345
+ $X2=2.235 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_2%A_27_367# 1 2 3 4 13 15 17 21 23 25 26 27 31
+ 36
r41 29 31 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=2.915 $Y=2.905
+ $X2=2.915 $Y2=2.435
r42 28 40 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.115 $Y=2.99
+ $X2=2.01 $Y2=2.99
r43 27 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.785 $Y=2.99
+ $X2=2.915 $Y2=2.905
r44 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.785 $Y=2.99
+ $X2=2.115 $Y2=2.99
r45 26 40 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=2.905
+ $X2=2.01 $Y2=2.99
r46 25 38 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=2.125
+ $X2=2.01 $Y2=2.04
r47 25 26 41.1948 $w=2.08e-07 $l=7.8e-07 $layer=LI1_cond $X=2.01 $Y=2.125
+ $X2=2.01 $Y2=2.905
r48 24 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.235 $Y=2.04
+ $X2=1.13 $Y2=2.04
r49 23 38 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.905 $Y=2.04
+ $X2=2.01 $Y2=2.04
r50 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.905 $Y=2.04
+ $X2=1.235 $Y2=2.04
r51 19 36 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=2.125
+ $X2=1.13 $Y2=2.04
r52 19 21 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.13 $Y=2.125
+ $X2=1.13 $Y2=2.495
r53 18 34 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.355 $Y=2.04
+ $X2=0.225 $Y2=2.04
r54 17 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.025 $Y=2.04
+ $X2=1.13 $Y2=2.04
r55 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=2.04
+ $X2=0.355 $Y2=2.04
r56 13 34 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=2.125
+ $X2=0.225 $Y2=2.04
r57 13 15 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=2.125
+ $X2=0.225 $Y2=2.495
r58 4 31 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=2.74
+ $Y=1.835 $X2=2.88 $Y2=2.435
r59 3 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.88
+ $Y=1.835 $X2=2.02 $Y2=2.91
r60 3 38 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=1.88
+ $Y=1.835 $X2=2.02 $Y2=2.12
r61 2 36 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.04
r62 2 21 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.495
r63 1 34 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.04
r64 1 15 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_2%VPWR 1 2 9 13 15 17 22 29 30 33 36
r45 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.57 $Y2=3.33
r48 27 29 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r52 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=3.33
+ $X2=1.57 $Y2=3.33
r54 22 25 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r58 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 15 30 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r60 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 15 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=3.245
+ $X2=1.57 $Y2=3.33
r63 11 13 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=1.57 $Y=3.245
+ $X2=1.57 $Y2=2.42
r64 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r65 7 9 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.42
r66 2 13 300 $w=1.7e-07 $l=6.6017e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=1.835 $X2=1.57 $Y2=2.42
r67 1 9 300 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_2%Y 1 2 3 10 16 18 20 23 28 29 33 34
r48 33 34 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.122 $Y=1.295
+ $X2=3.122 $Y2=1.665
r49 32 34 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=3.122 $Y=1.93
+ $X2=3.122 $Y2=1.665
r50 31 33 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=3.122 $Y=1.175
+ $X2=3.122 $Y2=1.295
r51 29 30 8.33171 $w=2.05e-07 $l=1.4e-07 $layer=LI1_cond $X=2.44 $Y=0.95
+ $X2=2.44 $Y2=1.09
r52 23 25 9.31762 $w=2.33e-07 $l=1.9e-07 $layer=LI1_cond $X=1.142 $Y=0.76
+ $X2=1.142 $Y2=0.95
r53 21 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=2.015
+ $X2=2.45 $Y2=2.015
r54 20 32 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=2.97 $Y=2.015
+ $X2=3.122 $Y2=1.93
r55 20 21 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.97 $Y=2.015
+ $X2=2.615 $Y2=2.015
r56 19 30 1.83547 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.545 $Y=1.09
+ $X2=2.44 $Y2=1.09
r57 18 31 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=2.97 $Y=1.09
+ $X2=3.122 $Y2=1.175
r58 18 19 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.97 $Y=1.09
+ $X2=2.545 $Y2=1.09
r59 14 29 4.9381 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.865 $X2=2.44
+ $Y2=0.95
r60 14 16 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=2.44 $Y=0.865
+ $X2=2.44 $Y2=0.42
r61 11 25 2.6346 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=1.26 $Y=0.95
+ $X2=1.142 $Y2=0.95
r62 10 29 1.83547 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.335 $Y=0.95
+ $X2=2.44 $Y2=0.95
r63 10 11 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=2.335 $Y=0.95
+ $X2=1.26 $Y2=0.95
r64 3 28 300 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=2 $X=2.31 $Y=1.835
+ $X2=2.45 $Y2=2.015
r65 2 16 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.31
+ $Y=0.235 $X2=2.45 $Y2=0.42
r66 1 23 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_2%VGND 1 2 3 10 12 16 20 23 24 26 27 28 41 42
r45 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 39 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r48 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r49 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r50 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r51 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 30 45 4.12789 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.177
+ $Y2=0
r53 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.72
+ $Y2=0
r54 28 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r55 28 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r56 28 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r57 26 38 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.64
+ $Y2=0
r58 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.88
+ $Y2=0
r59 25 41 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.12
+ $Y2=0
r60 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=2.88
+ $Y2=0
r61 23 35 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.68
+ $Y2=0
r62 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2
+ $Y2=0
r63 22 38 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.64
+ $Y2=0
r64 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2
+ $Y2=0
r65 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=0.085
+ $X2=2.88 $Y2=0
r66 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.88 $Y=0.085
+ $X2=2.88 $Y2=0.38
r67 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0
r68 14 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0.55
r69 10 45 3.08432 $w=2.6e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.177 $Y2=0
r70 10 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.38
r71 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.74
+ $Y=0.235 $X2=2.88 $Y2=0.38
r72 2 16 182 $w=1.7e-07 $l=3.86814e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=2 $Y2=0.55
r73 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_2%A_110_47# 1 2 9 11 12
r19 11 16 9.31762 $w=2.33e-07 $l=1.9e-07 $layer=LI1_cond $X=1.547 $Y=0.34
+ $X2=1.547 $Y2=0.53
r20 11 12 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.43 $Y=0.34
+ $X2=0.855 $Y2=0.34
r21 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.69 $Y=0.425
+ $X2=0.855 $Y2=0.34
r22 7 9 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=0.425 $X2=0.69
+ $Y2=0.43
r23 2 16 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.53
r24 1 9 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.43
.ends

