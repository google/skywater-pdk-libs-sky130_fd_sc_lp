* File: sky130_fd_sc_lp__or3b_lp.pxi.spice
* Created: Fri Aug 28 11:24:20 2020
* 
x_PM_SKY130_FD_SC_LP__OR3B_LP%C_N N_C_N_c_98_n N_C_N_M1002_g N_C_N_c_99_n
+ N_C_N_M1001_g N_C_N_c_100_n N_C_N_c_101_n N_C_N_M1014_g N_C_N_c_102_n
+ N_C_N_c_108_n C_N C_N N_C_N_c_104_n N_C_N_c_105_n
+ PM_SKY130_FD_SC_LP__OR3B_LP%C_N
x_PM_SKY130_FD_SC_LP__OR3B_LP%A_27_47# N_A_27_47#_M1002_s N_A_27_47#_M1001_s
+ N_A_27_47#_M1003_g N_A_27_47#_c_147_n N_A_27_47#_M1004_g N_A_27_47#_c_149_n
+ N_A_27_47#_M1010_g N_A_27_47#_c_151_n N_A_27_47#_c_152_n N_A_27_47#_c_153_n
+ N_A_27_47#_c_160_n N_A_27_47#_c_154_n N_A_27_47#_c_155_n N_A_27_47#_c_156_n
+ N_A_27_47#_c_161_n N_A_27_47#_c_157_n N_A_27_47#_c_158_n
+ PM_SKY130_FD_SC_LP__OR3B_LP%A_27_47#
x_PM_SKY130_FD_SC_LP__OR3B_LP%B N_B_M1009_g N_B_c_234_n N_B_M1006_g N_B_M1008_g
+ B B N_B_c_237_n N_B_c_238_n PM_SKY130_FD_SC_LP__OR3B_LP%B
x_PM_SKY130_FD_SC_LP__OR3B_LP%A N_A_c_293_n N_A_M1013_g N_A_M1012_g N_A_c_295_n
+ N_A_M1005_g A A N_A_c_297_n PM_SKY130_FD_SC_LP__OR3B_LP%A
x_PM_SKY130_FD_SC_LP__OR3B_LP%A_350_47# N_A_350_47#_M1004_d N_A_350_47#_M1006_d
+ N_A_350_47#_M1010_d N_A_350_47#_M1007_g N_A_350_47#_M1011_g
+ N_A_350_47#_M1000_g N_A_350_47#_c_341_n N_A_350_47#_c_354_n
+ N_A_350_47#_c_342_n N_A_350_47#_c_343_n N_A_350_47#_c_344_n
+ N_A_350_47#_c_345_n N_A_350_47#_c_346_n N_A_350_47#_c_391_n
+ N_A_350_47#_c_357_n N_A_350_47#_c_347_n N_A_350_47#_c_348_n
+ N_A_350_47#_c_349_n N_A_350_47#_c_359_n N_A_350_47#_c_350_n
+ N_A_350_47#_c_351_n N_A_350_47#_c_352_n PM_SKY130_FD_SC_LP__OR3B_LP%A_350_47#
x_PM_SKY130_FD_SC_LP__OR3B_LP%VPWR N_VPWR_M1001_d N_VPWR_M1012_d N_VPWR_c_478_n
+ N_VPWR_c_479_n N_VPWR_c_480_n N_VPWR_c_481_n VPWR N_VPWR_c_482_n
+ N_VPWR_c_477_n N_VPWR_c_484_n PM_SKY130_FD_SC_LP__OR3B_LP%VPWR
x_PM_SKY130_FD_SC_LP__OR3B_LP%A_263_373# N_A_263_373#_M1010_s
+ N_A_263_373#_M1008_s N_A_263_373#_c_524_n N_A_263_373#_c_525_n
+ N_A_263_373#_c_526_n N_A_263_373#_c_527_n
+ PM_SKY130_FD_SC_LP__OR3B_LP%A_263_373#
x_PM_SKY130_FD_SC_LP__OR3B_LP%X N_X_M1000_d N_X_M1011_d X X X X X X X X X
+ PM_SKY130_FD_SC_LP__OR3B_LP%X
x_PM_SKY130_FD_SC_LP__OR3B_LP%VGND N_VGND_M1014_d N_VGND_M1009_s N_VGND_M1005_d
+ N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n N_VGND_c_591_n N_VGND_c_592_n
+ N_VGND_c_593_n VGND N_VGND_c_594_n N_VGND_c_595_n N_VGND_c_596_n
+ N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n PM_SKY130_FD_SC_LP__OR3B_LP%VGND
cc_1 VNB N_C_N_c_98_n 0.0172366f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_2 VNB N_C_N_c_99_n 0.025655f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.668
cc_3 VNB N_C_N_c_100_n 0.0163702f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_4 VNB N_C_N_c_101_n 0.0137047f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_5 VNB N_C_N_c_102_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_6 VNB C_N 0.0112707f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_C_N_c_104_n 0.0158455f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.34
cc_8 VNB N_C_N_c_105_n 0.0166838f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.175
cc_9 VNB N_A_27_47#_M1003_g 0.0350089f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_10 VNB N_A_27_47#_c_147_n 0.0141374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1004_g 0.0373683f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_12 VNB N_A_27_47#_c_149_n 0.0121976f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_A_27_47#_M1010_g 0.0127056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_151_n 0.00620239f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.34
cc_15 VNB N_A_27_47#_c_152_n 0.00710603f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.34
cc_16 VNB N_A_27_47#_c_153_n 0.0227354f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_17 VNB N_A_27_47#_c_154_n 0.0104883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_155_n 0.0144053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_156_n 0.0141481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_157_n 0.0310373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_158_n 0.0382587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_M1009_g 0.0232158f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_23 VNB N_B_c_234_n 0.00299278f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.352
cc_24 VNB N_B_M1006_g 0.0253395f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_25 VNB B 0.0010685f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_26 VNB N_B_c_237_n 0.00241538f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_27 VNB N_B_c_238_n 0.022157f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.34
cc_28 VNB N_A_c_293_n 0.0181432f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_29 VNB N_A_M1012_g 0.011684f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.352
cc_30 VNB N_A_c_295_n 0.0156116f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.845
cc_31 VNB A 0.0119409f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_32 VNB N_A_c_297_n 0.049575f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_33 VNB N_A_350_47#_M1007_g 0.0246186f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_34 VNB N_A_350_47#_M1000_g 0.0286471f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_35 VNB N_A_350_47#_c_341_n 0.0196526f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.34
cc_36 VNB N_A_350_47#_c_342_n 0.00396917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_350_47#_c_343_n 0.00198372f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_38 VNB N_A_350_47#_c_344_n 0.00450354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_350_47#_c_345_n 0.0065387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_350_47#_c_346_n 8.58154e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_350_47#_c_347_n 2.06942e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_350_47#_c_348_n 0.00121962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_350_47#_c_349_n 0.0237817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_350_47#_c_350_n 0.00853836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_350_47#_c_351_n 0.00324766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_350_47#_c_352_n 0.0083159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VPWR_c_477_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB X 0.0161508f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.668
cc_49 VNB X 0.0452333f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.845
cc_50 VNB N_VGND_c_588_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_51 VNB N_VGND_c_589_n 0.0085253f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_52 VNB N_VGND_c_590_n 0.0213087f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_53 VNB N_VGND_c_591_n 0.0151056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_592_n 0.0258279f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.34
cc_55 VNB N_VGND_c_593_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.175
cc_56 VNB N_VGND_c_594_n 0.0266849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_595_n 0.0343386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_596_n 0.028795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_597_n 0.297317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_598_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_599_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VPB N_C_N_c_99_n 0.00108488f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.668
cc_63 VPB N_C_N_M1001_g 0.0376856f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_64 VPB N_C_N_c_108_n 0.0189991f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.845
cc_65 VPB C_N 0.00879429f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_66 VPB N_A_27_47#_M1010_g 0.0354808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_27_47#_c_160_n 0.0361574f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_c_161_n 0.013212f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_c_157_n 0.0175119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_B_c_234_n 0.0109094f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.352
cc_71 VPB N_B_M1008_g 0.0284829f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.805
cc_72 VPB B 0.0059346f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_73 VPB N_B_c_237_n 0.010711f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_74 VPB N_B_c_238_n 0.0331323f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.34
cc_75 VPB N_A_M1012_g 0.0388183f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.352
cc_76 VPB N_A_350_47#_M1011_g 0.0321176f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_77 VPB N_A_350_47#_c_354_n 0.0213398f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.175
cc_78 VPB N_A_350_47#_c_343_n 0.0155482f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.665
cc_79 VPB N_A_350_47#_c_346_n 0.00640958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_350_47#_c_357_n 0.00388006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_350_47#_c_349_n 0.00332148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_350_47#_c_359_n 0.00127447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_478_n 0.022459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_479_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.805
cc_85 VPB N_VPWR_c_480_n 0.0676588f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_86 VPB N_VPWR_c_481_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_482_n 0.0258985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_477_n 0.0732158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_484_n 0.0242279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_263_373#_c_524_n 0.0161454f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_91 VPB N_A_263_373#_c_525_n 0.0257134f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.805
cc_92 VPB N_A_263_373#_c_526_n 0.00488402f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.73
cc_93 VPB N_A_263_373#_c_527_n 0.00829285f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_94 VPB X 0.0216914f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.845
cc_95 VPB X 0.0142436f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB X 0.016179f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.805
cc_97 VPB X 0.0174462f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.805
cc_98 N_C_N_c_101_n N_A_27_47#_M1003_g 0.0181613f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_99 N_C_N_c_105_n N_A_27_47#_M1003_g 0.00139025f $X=0.597 $Y=1.175 $X2=0 $Y2=0
cc_100 N_C_N_c_98_n N_A_27_47#_c_153_n 0.00943525f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_101 N_C_N_c_101_n N_A_27_47#_c_153_n 0.00145474f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_102 N_C_N_c_102_n N_A_27_47#_c_153_n 0.00638389f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_103 N_C_N_M1001_g N_A_27_47#_c_160_n 0.0157367f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_104 N_C_N_c_100_n N_A_27_47#_c_154_n 0.0145084f $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_105 N_C_N_c_102_n N_A_27_47#_c_154_n 0.00357648f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_106 C_N N_A_27_47#_c_154_n 0.0294547f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_107 N_C_N_c_104_n N_A_27_47#_c_154_n 6.56795e-19 $X=0.61 $Y=1.34 $X2=0 $Y2=0
cc_108 N_C_N_c_105_n N_A_27_47#_c_154_n 0.00353992f $X=0.597 $Y=1.175 $X2=0
+ $Y2=0
cc_109 C_N N_A_27_47#_c_155_n 0.02113f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_110 N_C_N_c_104_n N_A_27_47#_c_155_n 3.10453e-19 $X=0.61 $Y=1.34 $X2=0 $Y2=0
cc_111 N_C_N_c_105_n N_A_27_47#_c_155_n 0.00171797f $X=0.597 $Y=1.175 $X2=0
+ $Y2=0
cc_112 N_C_N_c_102_n N_A_27_47#_c_156_n 0.00125708f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_113 N_C_N_c_105_n N_A_27_47#_c_156_n 0.00390346f $X=0.597 $Y=1.175 $X2=0
+ $Y2=0
cc_114 N_C_N_M1001_g N_A_27_47#_c_161_n 0.00470718f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_115 C_N N_A_27_47#_c_157_n 0.0487787f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_116 N_C_N_c_105_n N_A_27_47#_c_157_n 0.0255038f $X=0.597 $Y=1.175 $X2=0 $Y2=0
cc_117 C_N N_A_27_47#_c_158_n 0.00176218f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_118 N_C_N_c_104_n N_A_27_47#_c_158_n 0.0148239f $X=0.61 $Y=1.34 $X2=0 $Y2=0
cc_119 N_C_N_M1001_g N_VPWR_c_478_n 0.0249766f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_120 N_C_N_c_108_n N_VPWR_c_478_n 8.16152e-19 $X=0.597 $Y=1.845 $X2=0 $Y2=0
cc_121 C_N N_VPWR_c_478_n 0.0161922f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_122 N_C_N_M1001_g N_VPWR_c_477_n 0.014085f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_123 N_C_N_M1001_g N_VPWR_c_484_n 0.00769046f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_124 N_C_N_M1001_g N_A_263_373#_c_524_n 0.00619099f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_125 N_C_N_M1001_g N_A_263_373#_c_526_n 4.4929e-19 $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_126 N_C_N_c_98_n N_VGND_c_588_n 0.00231629f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_127 N_C_N_c_101_n N_VGND_c_588_n 0.0119457f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_128 N_C_N_c_98_n N_VGND_c_594_n 0.00549284f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_129 N_C_N_c_100_n N_VGND_c_594_n 4.87571e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_130 N_C_N_c_101_n N_VGND_c_594_n 0.00486043f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_131 N_C_N_c_98_n N_VGND_c_597_n 0.00712159f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_132 N_C_N_c_100_n N_VGND_c_597_n 6.51792e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_133 N_C_N_c_101_n N_VGND_c_597_n 0.00437711f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_134 N_A_27_47#_M1004_g N_B_M1009_g 0.0119375f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_149_n N_B_M1009_g 0.00578518f $X=1.725 $Y=1.545 $X2=0 $Y2=0
cc_136 N_A_27_47#_M1010_g N_B_c_234_n 0.00578518f $X=1.725 $Y=2.365 $X2=0 $Y2=0
cc_137 N_A_27_47#_M1010_g N_B_c_238_n 0.00146093f $X=1.725 $Y=2.365 $X2=0 $Y2=0
cc_138 N_A_27_47#_M1003_g N_A_350_47#_c_342_n 0.00460528f $X=1.285 $Y=0.445
+ $X2=0 $Y2=0
cc_139 N_A_27_47#_c_147_n N_A_350_47#_c_342_n 0.00425183f $X=1.6 $Y=1.195 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_M1004_g N_A_350_47#_c_342_n 0.0111796f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_c_151_n N_A_350_47#_c_342_n 0.00344961f $X=1.675 $Y=1.195
+ $X2=0 $Y2=0
cc_142 N_A_27_47#_c_152_n N_A_350_47#_c_342_n 0.00185319f $X=1.725 $Y=1.42 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_c_154_n N_A_350_47#_c_342_n 0.0130073f $X=1.015 $Y=0.91 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_c_155_n N_A_350_47#_c_342_n 0.0231179f $X=1.18 $Y=1.285 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_c_158_n N_A_350_47#_c_342_n 3.23682e-19 $X=1.36 $Y=1.285 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_c_149_n N_A_350_47#_c_343_n 0.00288768f $X=1.725 $Y=1.545
+ $X2=0 $Y2=0
cc_147 N_A_27_47#_M1010_g N_A_350_47#_c_343_n 0.0362226f $X=1.725 $Y=2.365 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_147_n N_A_350_47#_c_345_n 6.28633e-19 $X=1.6 $Y=1.195 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_149_n N_A_350_47#_c_345_n 0.0146628f $X=1.725 $Y=1.545 $X2=0
+ $Y2=0
cc_150 N_A_27_47#_c_152_n N_A_350_47#_c_345_n 0.00507611f $X=1.725 $Y=1.42 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_c_155_n N_A_350_47#_c_345_n 0.0100165f $X=1.18 $Y=1.285 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_158_n N_A_350_47#_c_345_n 8.43396e-19 $X=1.36 $Y=1.285 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_M1010_g N_A_350_47#_c_346_n 0.00137754f $X=1.725 $Y=2.365
+ $X2=0 $Y2=0
cc_154 N_A_27_47#_M1010_g N_A_350_47#_c_357_n 4.51726e-19 $X=1.725 $Y=2.365
+ $X2=0 $Y2=0
cc_155 N_A_27_47#_M1003_g N_A_350_47#_c_350_n 0.00362547f $X=1.285 $Y=0.445
+ $X2=0 $Y2=0
cc_156 N_A_27_47#_M1004_g N_A_350_47#_c_350_n 0.0112869f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_M1010_g N_VPWR_c_478_n 0.00221883f $X=1.725 $Y=2.365 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_c_161_n N_VPWR_c_478_n 0.0688031f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_159 N_A_27_47#_M1010_g N_VPWR_c_480_n 0.00132743f $X=1.725 $Y=2.365 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_160_n N_VPWR_c_477_n 0.0133547f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_160_n N_VPWR_c_484_n 0.0233806f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_147_n N_A_263_373#_c_524_n 0.0049538f $X=1.6 $Y=1.195 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_M1010_g N_A_263_373#_c_524_n 0.0246754f $X=1.725 $Y=2.365
+ $X2=0 $Y2=0
cc_164 N_A_27_47#_c_155_n N_A_263_373#_c_524_n 0.00226065f $X=1.18 $Y=1.285
+ $X2=0 $Y2=0
cc_165 N_A_27_47#_c_158_n N_A_263_373#_c_524_n 9.46444e-19 $X=1.36 $Y=1.285
+ $X2=0 $Y2=0
cc_166 N_A_27_47#_M1010_g N_A_263_373#_c_525_n 0.0171617f $X=1.725 $Y=2.365
+ $X2=0 $Y2=0
cc_167 N_A_27_47#_M1010_g N_A_263_373#_c_526_n 0.00264388f $X=1.725 $Y=2.365
+ $X2=0 $Y2=0
cc_168 N_A_27_47#_M1003_g N_VGND_c_588_n 0.0107313f $X=1.285 $Y=0.445 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_M1004_g N_VGND_c_588_n 0.00160329f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_153_n N_VGND_c_588_n 0.0127713f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_154_n N_VGND_c_588_n 0.0217339f $X=1.015 $Y=0.91 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_158_n N_VGND_c_588_n 7.11652e-19 $X=1.36 $Y=1.285 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_M1004_g N_VGND_c_589_n 0.00217641f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_M1004_g N_VGND_c_590_n 0.00552453f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_M1003_g N_VGND_c_592_n 0.00486043f $X=1.285 $Y=0.445 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1004_g N_VGND_c_592_n 0.00359964f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_153_n N_VGND_c_594_n 0.021137f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_178 N_A_27_47#_M1002_s N_VGND_c_597_n 0.00232985f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1003_g N_VGND_c_597_n 0.00491755f $X=1.285 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_M1004_g N_VGND_c_597_n 0.00670631f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_153_n N_VGND_c_597_n 0.0133547f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_154_n N_VGND_c_597_n 0.0183091f $X=1.015 $Y=0.91 $X2=0 $Y2=0
cc_183 N_B_M1006_g N_A_c_293_n 0.0167677f $X=2.615 $Y=1.135 $X2=-0.19 $Y2=-0.245
cc_184 B N_A_M1012_g 0.0272694f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_185 N_B_c_238_n N_A_M1012_g 0.0935916f $X=3.015 $Y=1.77 $X2=0 $Y2=0
cc_186 N_B_M1006_g A 0.00119796f $X=2.615 $Y=1.135 $X2=0 $Y2=0
cc_187 B A 0.0422525f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_188 N_B_c_238_n A 0.00192142f $X=3.015 $Y=1.77 $X2=0 $Y2=0
cc_189 N_B_M1006_g N_A_c_297_n 0.00392685f $X=2.615 $Y=1.135 $X2=0 $Y2=0
cc_190 B N_A_c_297_n 0.0016443f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_191 N_B_c_238_n N_A_c_297_n 0.00506941f $X=3.015 $Y=1.77 $X2=0 $Y2=0
cc_192 B N_A_350_47#_M1011_g 8.32612e-19 $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_193 N_B_M1009_g N_A_350_47#_c_342_n 0.00104629f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_194 N_B_M1009_g N_A_350_47#_c_343_n 0.0031805f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_195 N_B_c_238_n N_A_350_47#_c_343_n 7.04631e-19 $X=3.015 $Y=1.77 $X2=0 $Y2=0
cc_196 N_B_M1009_g N_A_350_47#_c_344_n 0.0144144f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_197 N_B_c_237_n N_A_350_47#_c_344_n 0.00109625f $X=2.54 $Y=1.77 $X2=0 $Y2=0
cc_198 N_B_M1009_g N_A_350_47#_c_346_n 7.46315e-19 $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_199 N_B_M1006_g N_A_350_47#_c_346_n 0.00566289f $X=2.615 $Y=1.135 $X2=0 $Y2=0
cc_200 N_B_M1008_g N_A_350_47#_c_346_n 0.00716964f $X=3.015 $Y=2.595 $X2=0 $Y2=0
cc_201 B N_A_350_47#_c_346_n 0.0360251f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_202 N_B_c_237_n N_A_350_47#_c_346_n 0.00525248f $X=2.54 $Y=1.77 $X2=0 $Y2=0
cc_203 N_B_c_238_n N_A_350_47#_c_346_n 0.0135989f $X=3.015 $Y=1.77 $X2=0 $Y2=0
cc_204 N_B_M1008_g N_A_350_47#_c_391_n 0.0185993f $X=3.015 $Y=2.595 $X2=0 $Y2=0
cc_205 B N_A_350_47#_c_391_n 0.0484768f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_206 N_B_c_238_n N_A_350_47#_c_391_n 0.00575703f $X=3.015 $Y=1.77 $X2=0 $Y2=0
cc_207 N_B_M1009_g N_A_350_47#_c_347_n 0.00120858f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_208 N_B_M1006_g N_A_350_47#_c_347_n 0.0110991f $X=2.615 $Y=1.135 $X2=0 $Y2=0
cc_209 B N_A_350_47#_c_348_n 0.0380091f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_210 B N_A_350_47#_c_349_n 0.00154299f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_211 N_B_M1006_g N_A_350_47#_c_351_n 0.0137334f $X=2.615 $Y=1.135 $X2=0 $Y2=0
cc_212 B N_A_350_47#_c_351_n 0.00111051f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_213 N_B_c_238_n N_A_350_47#_c_351_n 0.00517442f $X=3.015 $Y=1.77 $X2=0 $Y2=0
cc_214 N_B_M1006_g N_A_350_47#_c_352_n 0.00239739f $X=2.615 $Y=1.135 $X2=0 $Y2=0
cc_215 B N_VPWR_M1012_d 8.21888e-19 $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_216 N_B_M1008_g N_VPWR_c_479_n 0.00269982f $X=3.015 $Y=2.595 $X2=0 $Y2=0
cc_217 N_B_M1008_g N_VPWR_c_480_n 0.00939541f $X=3.015 $Y=2.595 $X2=0 $Y2=0
cc_218 N_B_M1008_g N_VPWR_c_477_n 0.0108803f $X=3.015 $Y=2.595 $X2=0 $Y2=0
cc_219 B N_A_263_373#_M1008_s 8.7279e-19 $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_220 N_B_M1008_g N_A_263_373#_c_527_n 0.00810934f $X=3.015 $Y=2.595 $X2=0
+ $Y2=0
cc_221 B A_628_419# 0.00141946f $X=3.515 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_222 N_B_M1009_g N_VGND_c_589_n 0.00905652f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_223 N_B_M1006_g N_VGND_c_589_n 0.00177558f $X=2.615 $Y=1.135 $X2=0 $Y2=0
cc_224 N_B_M1009_g N_VGND_c_590_n 0.00499358f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_225 N_B_M1006_g N_VGND_c_590_n 6.20616e-19 $X=2.615 $Y=1.135 $X2=0 $Y2=0
cc_226 N_B_M1009_g N_VGND_c_597_n 0.00147066f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_227 N_B_M1006_g N_VGND_c_597_n 0.00302011f $X=2.615 $Y=1.135 $X2=0 $Y2=0
cc_228 N_A_c_295_n N_A_350_47#_M1007_g 0.0142126f $X=3.515 $Y=1.035 $X2=0 $Y2=0
cc_229 A N_A_350_47#_M1007_g 0.00668888f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_230 N_A_M1012_g N_A_350_47#_M1011_g 0.0329931f $X=3.505 $Y=2.595 $X2=0 $Y2=0
cc_231 N_A_c_297_n N_A_350_47#_c_341_n 0.029047f $X=3.505 $Y=1.262 $X2=0 $Y2=0
cc_232 N_A_M1012_g N_A_350_47#_c_391_n 0.0174787f $X=3.505 $Y=2.595 $X2=0 $Y2=0
cc_233 N_A_c_293_n N_A_350_47#_c_347_n 0.00359743f $X=3.125 $Y=1.035 $X2=0 $Y2=0
cc_234 A N_A_350_47#_c_347_n 0.0231296f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_235 N_A_c_297_n N_A_350_47#_c_347_n 8.73072e-19 $X=3.505 $Y=1.262 $X2=0 $Y2=0
cc_236 N_A_M1012_g N_A_350_47#_c_348_n 2.27062e-19 $X=3.505 $Y=2.595 $X2=0 $Y2=0
cc_237 A N_A_350_47#_c_348_n 0.0148806f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_238 N_A_c_297_n N_A_350_47#_c_348_n 0.00189249f $X=3.505 $Y=1.262 $X2=0 $Y2=0
cc_239 N_A_M1012_g N_A_350_47#_c_349_n 0.0148344f $X=3.505 $Y=2.595 $X2=0 $Y2=0
cc_240 N_A_M1012_g N_A_350_47#_c_359_n 0.0042936f $X=3.505 $Y=2.595 $X2=0 $Y2=0
cc_241 A N_A_350_47#_c_351_n 0.0074554f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_242 N_A_c_297_n N_A_350_47#_c_351_n 0.00197368f $X=3.505 $Y=1.262 $X2=0 $Y2=0
cc_243 N_A_c_293_n N_A_350_47#_c_352_n 0.00718598f $X=3.125 $Y=1.035 $X2=0 $Y2=0
cc_244 N_A_c_295_n N_A_350_47#_c_352_n 0.00104143f $X=3.515 $Y=1.035 $X2=0 $Y2=0
cc_245 A N_A_350_47#_c_352_n 0.00362384f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_246 N_A_M1012_g N_VPWR_c_479_n 0.0139597f $X=3.505 $Y=2.595 $X2=0 $Y2=0
cc_247 N_A_M1012_g N_VPWR_c_480_n 0.008763f $X=3.505 $Y=2.595 $X2=0 $Y2=0
cc_248 N_A_M1012_g N_VPWR_c_477_n 0.00771816f $X=3.505 $Y=2.595 $X2=0 $Y2=0
cc_249 N_A_M1012_g N_A_263_373#_c_527_n 0.00166433f $X=3.505 $Y=2.595 $X2=0
+ $Y2=0
cc_250 N_A_M1012_g X 8.00949e-19 $X=3.505 $Y=2.595 $X2=0 $Y2=0
cc_251 N_A_c_293_n N_VGND_c_590_n 0.00277487f $X=3.125 $Y=1.035 $X2=0 $Y2=0
cc_252 N_A_c_293_n N_VGND_c_591_n 0.00159629f $X=3.125 $Y=1.035 $X2=0 $Y2=0
cc_253 N_A_c_295_n N_VGND_c_591_n 0.0104539f $X=3.515 $Y=1.035 $X2=0 $Y2=0
cc_254 A N_VGND_c_591_n 0.009847f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_255 N_A_c_293_n N_VGND_c_595_n 0.00463701f $X=3.125 $Y=1.035 $X2=0 $Y2=0
cc_256 N_A_c_295_n N_VGND_c_595_n 0.00402651f $X=3.515 $Y=1.035 $X2=0 $Y2=0
cc_257 N_A_c_293_n N_VGND_c_597_n 0.00503886f $X=3.125 $Y=1.035 $X2=0 $Y2=0
cc_258 N_A_c_295_n N_VGND_c_597_n 0.00423264f $X=3.515 $Y=1.035 $X2=0 $Y2=0
cc_259 N_A_350_47#_c_391_n N_VPWR_M1012_d 0.0101753f $X=3.895 $Y=2.415 $X2=0
+ $Y2=0
cc_260 N_A_350_47#_c_359_n N_VPWR_M1012_d 0.00272321f $X=3.98 $Y=2.33 $X2=0
+ $Y2=0
cc_261 N_A_350_47#_M1011_g N_VPWR_c_479_n 0.00790974f $X=4.145 $Y=2.595 $X2=0
+ $Y2=0
cc_262 N_A_350_47#_c_391_n N_VPWR_c_479_n 0.0206735f $X=3.895 $Y=2.415 $X2=0
+ $Y2=0
cc_263 N_A_350_47#_M1011_g N_VPWR_c_482_n 0.00938036f $X=4.145 $Y=2.595 $X2=0
+ $Y2=0
cc_264 N_A_350_47#_M1011_g N_VPWR_c_477_n 0.0161106f $X=4.145 $Y=2.595 $X2=0
+ $Y2=0
cc_265 N_A_350_47#_c_391_n N_VPWR_c_477_n 0.0272579f $X=3.895 $Y=2.415 $X2=0
+ $Y2=0
cc_266 N_A_350_47#_c_357_n N_VPWR_c_477_n 6.34548e-19 $X=2.63 $Y=2.415 $X2=0
+ $Y2=0
cc_267 N_A_350_47#_c_346_n N_A_263_373#_M1008_s 0.00299706f $X=2.545 $Y=2.33
+ $X2=0 $Y2=0
cc_268 N_A_350_47#_c_391_n N_A_263_373#_M1008_s 0.00562492f $X=3.895 $Y=2.415
+ $X2=0 $Y2=0
cc_269 N_A_350_47#_c_357_n N_A_263_373#_M1008_s 5.03301e-19 $X=2.63 $Y=2.415
+ $X2=0 $Y2=0
cc_270 N_A_350_47#_c_343_n N_A_263_373#_c_524_n 0.0573249f $X=1.99 $Y=2.01 $X2=0
+ $Y2=0
cc_271 N_A_350_47#_c_345_n N_A_263_373#_c_524_n 0.00485786f $X=2.155 $Y=1.41
+ $X2=0 $Y2=0
cc_272 N_A_350_47#_c_343_n N_A_263_373#_c_525_n 0.0219639f $X=1.99 $Y=2.01 $X2=0
+ $Y2=0
cc_273 N_A_350_47#_c_357_n N_A_263_373#_c_525_n 0.00498407f $X=2.63 $Y=2.415
+ $X2=0 $Y2=0
cc_274 N_A_350_47#_c_343_n N_A_263_373#_c_527_n 0.00153516f $X=1.99 $Y=2.01
+ $X2=0 $Y2=0
cc_275 N_A_350_47#_c_391_n N_A_263_373#_c_527_n 0.0162429f $X=3.895 $Y=2.415
+ $X2=0 $Y2=0
cc_276 N_A_350_47#_c_357_n N_A_263_373#_c_527_n 0.00355583f $X=2.63 $Y=2.415
+ $X2=0 $Y2=0
cc_277 N_A_350_47#_c_391_n A_628_419# 0.00388677f $X=3.895 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_278 N_A_350_47#_M1007_g X 0.00158012f $X=3.945 $Y=0.715 $X2=0 $Y2=0
cc_279 N_A_350_47#_M1000_g X 0.00727982f $X=4.305 $Y=0.715 $X2=0 $Y2=0
cc_280 N_A_350_47#_M1000_g X 0.0200527f $X=4.305 $Y=0.715 $X2=0 $Y2=0
cc_281 N_A_350_47#_c_348_n X 0.0425408f $X=4.06 $Y=1.39 $X2=0 $Y2=0
cc_282 N_A_350_47#_c_349_n X 0.0166809f $X=4.06 $Y=1.39 $X2=0 $Y2=0
cc_283 N_A_350_47#_c_359_n X 0.0072366f $X=3.98 $Y=2.33 $X2=0 $Y2=0
cc_284 N_A_350_47#_M1011_g X 0.00526614f $X=4.145 $Y=2.595 $X2=0 $Y2=0
cc_285 N_A_350_47#_c_341_n X 0.00308769f $X=4.125 $Y=1.375 $X2=0 $Y2=0
cc_286 N_A_350_47#_c_359_n X 0.0177357f $X=3.98 $Y=2.33 $X2=0 $Y2=0
cc_287 N_A_350_47#_M1011_g X 0.0122276f $X=4.145 $Y=2.595 $X2=0 $Y2=0
cc_288 N_A_350_47#_c_391_n X 0.013234f $X=3.895 $Y=2.415 $X2=0 $Y2=0
cc_289 N_A_350_47#_M1011_g X 0.00735125f $X=4.145 $Y=2.595 $X2=0 $Y2=0
cc_290 N_A_350_47#_c_345_n N_VGND_M1009_s 0.00248839f $X=2.155 $Y=1.41 $X2=0
+ $Y2=0
cc_291 N_A_350_47#_c_350_n N_VGND_c_588_n 0.0203482f $X=1.89 $Y=0.47 $X2=0 $Y2=0
cc_292 N_A_350_47#_c_342_n N_VGND_c_589_n 0.0187266f $X=1.61 $Y=1.325 $X2=0
+ $Y2=0
cc_293 N_A_350_47#_c_344_n N_VGND_c_589_n 0.00827348f $X=2.46 $Y=1.41 $X2=0
+ $Y2=0
cc_294 N_A_350_47#_c_345_n N_VGND_c_589_n 0.0214344f $X=2.155 $Y=1.41 $X2=0
+ $Y2=0
cc_295 N_A_350_47#_c_347_n N_VGND_c_589_n 0.0144251f $X=2.74 $Y=1.325 $X2=0
+ $Y2=0
cc_296 N_A_350_47#_c_350_n N_VGND_c_589_n 0.0124661f $X=1.89 $Y=0.47 $X2=0 $Y2=0
cc_297 N_A_350_47#_c_342_n N_VGND_c_590_n 0.006216f $X=1.61 $Y=1.325 $X2=0 $Y2=0
cc_298 N_A_350_47#_c_347_n N_VGND_c_590_n 0.00211705f $X=2.74 $Y=1.325 $X2=0
+ $Y2=0
cc_299 N_A_350_47#_c_350_n N_VGND_c_590_n 0.0324184f $X=1.89 $Y=0.47 $X2=0 $Y2=0
cc_300 N_A_350_47#_c_352_n N_VGND_c_590_n 0.0225473f $X=2.91 $Y=0.67 $X2=0 $Y2=0
cc_301 N_A_350_47#_M1007_g N_VGND_c_591_n 0.0109731f $X=3.945 $Y=0.715 $X2=0
+ $Y2=0
cc_302 N_A_350_47#_M1000_g N_VGND_c_591_n 0.00145557f $X=4.305 $Y=0.715 $X2=0
+ $Y2=0
cc_303 N_A_350_47#_c_352_n N_VGND_c_591_n 0.0119031f $X=2.91 $Y=0.67 $X2=0 $Y2=0
cc_304 N_A_350_47#_c_350_n N_VGND_c_592_n 0.0298581f $X=1.89 $Y=0.47 $X2=0 $Y2=0
cc_305 N_A_350_47#_c_352_n N_VGND_c_595_n 0.0114794f $X=2.91 $Y=0.67 $X2=0 $Y2=0
cc_306 N_A_350_47#_M1007_g N_VGND_c_596_n 0.00402651f $X=3.945 $Y=0.715 $X2=0
+ $Y2=0
cc_307 N_A_350_47#_M1000_g N_VGND_c_596_n 0.00463876f $X=4.305 $Y=0.715 $X2=0
+ $Y2=0
cc_308 N_A_350_47#_M1004_d N_VGND_c_597_n 0.00233022f $X=1.75 $Y=0.235 $X2=0
+ $Y2=0
cc_309 N_A_350_47#_M1007_g N_VGND_c_597_n 0.00423264f $X=3.945 $Y=0.715 $X2=0
+ $Y2=0
cc_310 N_A_350_47#_M1000_g N_VGND_c_597_n 0.00503886f $X=4.305 $Y=0.715 $X2=0
+ $Y2=0
cc_311 N_A_350_47#_c_350_n N_VGND_c_597_n 0.0195332f $X=1.89 $Y=0.47 $X2=0 $Y2=0
cc_312 N_A_350_47#_c_352_n N_VGND_c_597_n 0.013822f $X=2.91 $Y=0.67 $X2=0 $Y2=0
cc_313 N_A_350_47#_c_350_n A_272_47# 0.00437926f $X=1.89 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_314 N_A_350_47#_c_344_n A_466_185# 0.00225639f $X=2.46 $Y=1.41 $X2=-0.19
+ $Y2=-0.245
cc_315 N_A_350_47#_c_351_n A_466_185# 8.77578e-19 $X=2.74 $Y=1.41 $X2=-0.19
+ $Y2=-0.245
cc_316 N_VPWR_c_477_n N_A_263_373#_M1008_s 0.00232985f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_478_n N_A_263_373#_c_524_n 0.0467227f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_480_n N_A_263_373#_c_525_n 0.0581819f $X=3.605 $Y=3.33 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_477_n N_A_263_373#_c_525_n 0.035874f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_c_478_n N_A_263_373#_c_526_n 0.00968496f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_480_n N_A_263_373#_c_526_n 0.0222501f $X=3.605 $Y=3.33 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_477_n N_A_263_373#_c_526_n 0.0127687f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_480_n N_A_263_373#_c_527_n 0.0190464f $X=3.605 $Y=3.33 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_477_n N_A_263_373#_c_527_n 0.0123847f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_477_n A_628_419# 0.003486f $X=4.56 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_326 N_VPWR_c_477_n N_X_M1011_d 0.0023218f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_c_479_n X 0.0191282f $X=3.77 $Y=2.895 $X2=0 $Y2=0
cc_328 N_VPWR_c_482_n X 0.0234706f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_329 N_VPWR_c_477_n X 0.016409f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_330 X N_VGND_c_591_n 0.0138681f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_331 X N_VGND_c_596_n 0.0106031f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_332 X N_VGND_c_597_n 0.0113777f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_333 A_114_47# N_VGND_c_597_n 0.00303453f $X=0.57 $Y=0.235 $X2=4.56 $Y2=0
cc_334 N_VGND_c_597_n A_272_47# 0.00766269f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
cc_335 N_VGND_c_589_n A_466_185# 0.00238999f $X=2.235 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
