* File: sky130_fd_sc_lp__a22oi_lp.pxi.spice
* Created: Wed Sep  2 09:23:23 2020
* 
x_PM_SKY130_FD_SC_LP__A22OI_LP%B2 N_B2_M1004_g N_B2_M1005_g N_B2_c_58_n
+ N_B2_c_59_n B2 N_B2_c_61_n PM_SKY130_FD_SC_LP__A22OI_LP%B2
x_PM_SKY130_FD_SC_LP__A22OI_LP%B1 N_B1_M1007_g N_B1_M1002_g N_B1_c_95_n
+ N_B1_c_96_n B1 N_B1_c_98_n PM_SKY130_FD_SC_LP__A22OI_LP%B1
x_PM_SKY130_FD_SC_LP__A22OI_LP%A1 N_A1_M1000_g N_A1_M1006_g N_A1_c_139_n
+ N_A1_c_140_n A1 N_A1_c_141_n N_A1_c_142_n PM_SKY130_FD_SC_LP__A22OI_LP%A1
x_PM_SKY130_FD_SC_LP__A22OI_LP%A2 N_A2_M1003_g N_A2_M1001_g A2 N_A2_c_182_n
+ PM_SKY130_FD_SC_LP__A22OI_LP%A2
x_PM_SKY130_FD_SC_LP__A22OI_LP%A_64_409# N_A_64_409#_M1004_s N_A_64_409#_M1002_d
+ N_A_64_409#_M1001_d N_A_64_409#_c_206_n N_A_64_409#_c_207_n
+ N_A_64_409#_c_208_n N_A_64_409#_c_209_n N_A_64_409#_c_216_n
+ N_A_64_409#_c_210_n N_A_64_409#_c_211_n N_A_64_409#_c_212_n
+ PM_SKY130_FD_SC_LP__A22OI_LP%A_64_409#
x_PM_SKY130_FD_SC_LP__A22OI_LP%Y N_Y_M1007_d N_Y_M1004_d N_Y_c_259_n N_Y_c_263_n
+ N_Y_c_264_n N_Y_c_272_n N_Y_c_260_n Y Y Y N_Y_c_261_n Y
+ PM_SKY130_FD_SC_LP__A22OI_LP%Y
x_PM_SKY130_FD_SC_LP__A22OI_LP%VPWR N_VPWR_M1006_d N_VPWR_c_308_n N_VPWR_c_309_n
+ N_VPWR_c_310_n VPWR N_VPWR_c_311_n N_VPWR_c_307_n
+ PM_SKY130_FD_SC_LP__A22OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A22OI_LP%VGND N_VGND_M1005_s N_VGND_M1003_d N_VGND_c_337_n
+ N_VGND_c_338_n N_VGND_c_339_n VGND N_VGND_c_340_n N_VGND_c_341_n
+ N_VGND_c_342_n N_VGND_c_343_n PM_SKY130_FD_SC_LP__A22OI_LP%VGND
cc_1 VNB N_B2_M1005_g 0.0380115f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.445
cc_2 VNB N_B2_c_58_n 0.0256646f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.58
cc_3 VNB N_B2_c_59_n 0.00569481f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.745
cc_4 VNB B2 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_B2_c_61_n 0.0176374f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.24
cc_6 VNB N_B1_M1007_g 0.0323508f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=2.545
cc_7 VNB N_B1_c_95_n 0.023466f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.58
cc_8 VNB N_B1_c_96_n 0.00520696f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.745
cc_9 VNB B1 0.00170127f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_B1_c_98_n 0.0165176f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.24
cc_11 VNB N_A1_M1000_g 0.0381675f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=2.545
cc_12 VNB N_A1_c_139_n 0.0196784f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.58
cc_13 VNB N_A1_c_140_n 0.0043665f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.745
cc_14 VNB N_A1_c_141_n 0.0195118f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.24
cc_15 VNB N_A1_c_142_n 0.0111701f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.24
cc_16 VNB N_A2_M1003_g 0.030049f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=2.545
cc_17 VNB N_A2_M1001_g 0.0121064f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.445
cc_18 VNB A2 0.0289245f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.24
cc_19 VNB N_A2_c_182_n 0.0792177f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.745
cc_20 VNB N_Y_c_259_n 0.0324589f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.445
cc_21 VNB N_Y_c_260_n 0.00100281f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.24
cc_22 VNB N_Y_c_261_n 0.0115469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB Y 0.0386937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_307_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_337_n 0.0145548f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.24
cc_26 VNB N_VGND_c_338_n 0.014353f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.58
cc_27 VNB N_VGND_c_339_n 0.0212949f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_28 VNB N_VGND_c_340_n 0.0138531f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.24
cc_29 VNB N_VGND_c_341_n 0.0439035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_342_n 0.00510584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_343_n 0.174741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_B2_M1004_g 0.0392136f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=2.545
cc_33 VPB N_B2_c_59_n 0.00908871f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.745
cc_34 VPB B2 7.56276e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_35 VPB N_B1_M1002_g 0.0337718f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.445
cc_36 VPB N_B1_c_96_n 0.00845676f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.745
cc_37 VPB B1 7.45264e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_38 VPB N_A1_M1006_g 0.0336115f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.445
cc_39 VPB N_A1_c_140_n 0.00731246f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.745
cc_40 VPB N_A1_c_142_n 0.0021248f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.24
cc_41 VPB N_A2_M1001_g 0.0521038f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.445
cc_42 VPB N_A_64_409#_c_206_n 0.0236858f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.745
cc_43 VPB N_A_64_409#_c_207_n 0.00202865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_64_409#_c_208_n 0.00938685f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.24
cc_45 VPB N_A_64_409#_c_209_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.24
cc_46 VPB N_A_64_409#_c_210_n 0.0194859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_64_409#_c_211_n 0.00819087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_64_409#_c_212_n 0.0391242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_Y_c_263_n 0.0160414f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.24
cc_50 VPB N_Y_c_264_n 0.0155696f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.075
cc_51 VPB Y 0.0141649f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_308_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.445
cc_53 VPB N_VPWR_c_309_n 0.0487587f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.24
cc_54 VPB N_VPWR_c_310_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.075
cc_55 VPB N_VPWR_c_311_n 0.0194022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_307_n 0.0618284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 N_B2_M1005_g N_B1_M1007_g 0.0523413f $X=0.78 $Y=0.445 $X2=0 $Y2=0
cc_58 N_B2_M1004_g N_B1_M1002_g 0.0355146f $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_59 N_B2_c_58_n N_B1_c_95_n 0.0135694f $X=0.69 $Y=1.58 $X2=0 $Y2=0
cc_60 N_B2_c_59_n N_B1_c_96_n 0.0135694f $X=0.69 $Y=1.745 $X2=0 $Y2=0
cc_61 B2 B1 0.0423335f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_B2_c_61_n B1 0.00232658f $X=0.69 $Y=1.24 $X2=0 $Y2=0
cc_63 B2 N_B1_c_98_n 0.00232658f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_64 N_B2_c_61_n N_B1_c_98_n 0.0135694f $X=0.69 $Y=1.24 $X2=0 $Y2=0
cc_65 N_B2_M1004_g N_A_64_409#_c_206_n 0.0127599f $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_66 N_B2_M1004_g N_A_64_409#_c_207_n 0.0164477f $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_67 N_B2_M1004_g N_A_64_409#_c_208_n 9.65935e-19 $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_68 N_B2_M1004_g N_A_64_409#_c_216_n 7.1089e-19 $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_69 N_B2_M1005_g N_Y_c_259_n 0.0135656f $X=0.78 $Y=0.445 $X2=0 $Y2=0
cc_70 B2 N_Y_c_259_n 0.0245051f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_B2_c_61_n N_Y_c_259_n 0.00123061f $X=0.69 $Y=1.24 $X2=0 $Y2=0
cc_72 N_B2_M1004_g N_Y_c_263_n 0.0217809f $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_73 N_B2_c_59_n N_Y_c_263_n 5.43485e-19 $X=0.69 $Y=1.745 $X2=0 $Y2=0
cc_74 B2 N_Y_c_263_n 0.0242891f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_75 N_B2_M1004_g N_Y_c_272_n 0.0160162f $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_76 N_B2_M1005_g N_Y_c_260_n 0.00168185f $X=0.78 $Y=0.445 $X2=0 $Y2=0
cc_77 N_B2_M1004_g Y 0.00607662f $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_78 N_B2_M1005_g Y 0.00516327f $X=0.78 $Y=0.445 $X2=0 $Y2=0
cc_79 B2 Y 0.0491281f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B2_c_61_n Y 0.0149783f $X=0.69 $Y=1.24 $X2=0 $Y2=0
cc_81 N_B2_M1004_g N_VPWR_c_309_n 0.00546179f $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_82 N_B2_M1004_g N_VPWR_c_307_n 0.00814996f $X=0.73 $Y=2.545 $X2=0 $Y2=0
cc_83 N_B2_M1005_g N_VGND_c_337_n 0.0113946f $X=0.78 $Y=0.445 $X2=0 $Y2=0
cc_84 N_B2_M1005_g N_VGND_c_341_n 0.00364083f $X=0.78 $Y=0.445 $X2=0 $Y2=0
cc_85 N_B2_M1005_g N_VGND_c_343_n 0.00429664f $X=0.78 $Y=0.445 $X2=0 $Y2=0
cc_86 N_B1_M1007_g N_A1_M1000_g 0.0226843f $X=1.17 $Y=0.445 $X2=0 $Y2=0
cc_87 N_B1_M1002_g N_A1_M1006_g 0.0217656f $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_88 N_B1_c_95_n N_A1_c_139_n 0.0117589f $X=1.23 $Y=1.58 $X2=0 $Y2=0
cc_89 N_B1_c_96_n N_A1_c_140_n 0.0117589f $X=1.23 $Y=1.745 $X2=0 $Y2=0
cc_90 B1 N_A1_c_141_n 7.5249e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B1_c_98_n N_A1_c_141_n 0.0117589f $X=1.23 $Y=1.24 $X2=0 $Y2=0
cc_92 B1 N_A1_c_142_n 0.0514906f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_93 N_B1_c_98_n N_A1_c_142_n 0.00410596f $X=1.23 $Y=1.24 $X2=0 $Y2=0
cc_94 N_B1_M1002_g N_A_64_409#_c_206_n 7.1089e-19 $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_95 N_B1_M1002_g N_A_64_409#_c_207_n 0.0164696f $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_96 N_B1_M1002_g N_A_64_409#_c_209_n 8.05528e-19 $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_97 N_B1_M1002_g N_A_64_409#_c_216_n 0.0139941f $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_98 N_B1_M1002_g N_A_64_409#_c_211_n 0.00471192f $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_99 B1 N_A_64_409#_c_211_n 0.00278552f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B1_M1007_g N_Y_c_259_n 0.0114869f $X=1.17 $Y=0.445 $X2=0 $Y2=0
cc_101 B1 N_Y_c_259_n 0.0259012f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B1_c_98_n N_Y_c_259_n 0.00134249f $X=1.23 $Y=1.24 $X2=0 $Y2=0
cc_103 N_B1_M1002_g N_Y_c_263_n 0.00471192f $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_104 N_B1_c_96_n N_Y_c_263_n 5.35995e-19 $X=1.23 $Y=1.745 $X2=0 $Y2=0
cc_105 B1 N_Y_c_263_n 0.00790183f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B1_M1002_g N_Y_c_272_n 0.010704f $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_107 N_B1_M1007_g N_Y_c_260_n 0.0090314f $X=1.17 $Y=0.445 $X2=0 $Y2=0
cc_108 N_B1_M1002_g N_VPWR_c_308_n 8.74508e-19 $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_109 N_B1_M1002_g N_VPWR_c_309_n 0.00546179f $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_110 N_B1_M1002_g N_VPWR_c_307_n 0.00742485f $X=1.26 $Y=2.545 $X2=0 $Y2=0
cc_111 N_B1_M1007_g N_VGND_c_337_n 0.00202904f $X=1.17 $Y=0.445 $X2=0 $Y2=0
cc_112 N_B1_M1007_g N_VGND_c_341_n 0.00426341f $X=1.17 $Y=0.445 $X2=0 $Y2=0
cc_113 N_B1_M1007_g N_VGND_c_343_n 0.00630672f $X=1.17 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A1_M1000_g N_A2_M1003_g 0.0282532f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A1_M1006_g N_A2_M1001_g 0.0321554f $X=1.79 $Y=2.545 $X2=0 $Y2=0
cc_116 N_A1_c_139_n N_A2_M1001_g 0.0180257f $X=1.8 $Y=1.58 $X2=0 $Y2=0
cc_117 N_A1_M1000_g A2 9.95563e-19 $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_118 N_A1_c_141_n A2 4.74837e-19 $X=1.8 $Y=1.24 $X2=0 $Y2=0
cc_119 N_A1_c_142_n A2 0.0188721f $X=1.8 $Y=1.24 $X2=0 $Y2=0
cc_120 N_A1_c_141_n N_A2_c_182_n 0.0180257f $X=1.8 $Y=1.24 $X2=0 $Y2=0
cc_121 N_A1_c_142_n N_A2_c_182_n 0.00337014f $X=1.8 $Y=1.24 $X2=0 $Y2=0
cc_122 N_A1_M1006_g N_A_64_409#_c_209_n 0.00336125f $X=1.79 $Y=2.545 $X2=0 $Y2=0
cc_123 N_A1_M1006_g N_A_64_409#_c_216_n 0.0140379f $X=1.79 $Y=2.545 $X2=0 $Y2=0
cc_124 N_A1_M1006_g N_A_64_409#_c_210_n 0.0179194f $X=1.79 $Y=2.545 $X2=0 $Y2=0
cc_125 N_A1_c_140_n N_A_64_409#_c_210_n 0.00128924f $X=1.8 $Y=1.745 $X2=0 $Y2=0
cc_126 N_A1_c_142_n N_A_64_409#_c_210_n 0.0200417f $X=1.8 $Y=1.24 $X2=0 $Y2=0
cc_127 N_A1_M1006_g N_A_64_409#_c_211_n 0.00216835f $X=1.79 $Y=2.545 $X2=0 $Y2=0
cc_128 N_A1_c_140_n N_A_64_409#_c_211_n 8.1248e-19 $X=1.8 $Y=1.745 $X2=0 $Y2=0
cc_129 N_A1_c_142_n N_A_64_409#_c_211_n 0.00992419f $X=1.8 $Y=1.24 $X2=0 $Y2=0
cc_130 N_A1_M1006_g N_A_64_409#_c_212_n 9.45905e-19 $X=1.79 $Y=2.545 $X2=0 $Y2=0
cc_131 N_A1_M1000_g N_Y_c_259_n 0.00540896f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A1_M1000_g N_Y_c_260_n 0.0125935f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_133 N_A1_M1006_g N_VPWR_c_308_n 0.0189228f $X=1.79 $Y=2.545 $X2=0 $Y2=0
cc_134 N_A1_M1006_g N_VPWR_c_309_n 0.00767656f $X=1.79 $Y=2.545 $X2=0 $Y2=0
cc_135 N_A1_M1006_g N_VPWR_c_307_n 0.0134103f $X=1.79 $Y=2.545 $X2=0 $Y2=0
cc_136 N_A1_M1000_g N_VGND_c_339_n 0.00285442f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A1_M1000_g N_VGND_c_341_n 0.00585385f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_138 N_A1_M1000_g N_VGND_c_343_n 0.0116195f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A2_M1001_g N_A_64_409#_c_216_n 8.87218e-19 $X=2.33 $Y=2.545 $X2=0 $Y2=0
cc_140 N_A2_M1001_g N_A_64_409#_c_210_n 0.0261403f $X=2.33 $Y=2.545 $X2=0 $Y2=0
cc_141 A2 N_A_64_409#_c_210_n 0.0193135f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_142 N_A2_c_182_n N_A_64_409#_c_210_n 0.00470735f $X=2.495 $Y=1.02 $X2=0 $Y2=0
cc_143 N_A2_M1001_g N_A_64_409#_c_212_n 0.017771f $X=2.33 $Y=2.545 $X2=0 $Y2=0
cc_144 N_A2_M1001_g N_VPWR_c_308_n 0.0191596f $X=2.33 $Y=2.545 $X2=0 $Y2=0
cc_145 N_A2_M1001_g N_VPWR_c_311_n 0.00804781f $X=2.33 $Y=2.545 $X2=0 $Y2=0
cc_146 N_A2_M1001_g N_VPWR_c_307_n 0.0147099f $X=2.33 $Y=2.545 $X2=0 $Y2=0
cc_147 N_A2_M1003_g N_VGND_c_339_n 0.0162023f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_148 A2 N_VGND_c_339_n 0.027017f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A2_c_182_n N_VGND_c_339_n 0.00815362f $X=2.495 $Y=1.02 $X2=0 $Y2=0
cc_150 N_A2_M1003_g N_VGND_c_341_n 0.00486043f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_151 N_A2_M1003_g N_VGND_c_343_n 0.00870566f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_152 A2 N_VGND_c_343_n 0.00480119f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_153 N_A_64_409#_c_207_n N_Y_M1004_d 0.00180746f $X=1.36 $Y=2.98 $X2=0 $Y2=0
cc_154 N_A_64_409#_M1004_s N_Y_c_263_n 0.0024137f $X=0.32 $Y=2.045 $X2=0 $Y2=0
cc_155 N_A_64_409#_c_206_n N_Y_c_263_n 0.0174952f $X=0.465 $Y=2.44 $X2=0 $Y2=0
cc_156 N_A_64_409#_c_211_n N_Y_c_263_n 0.0126166f $X=1.69 $Y=2.01 $X2=0 $Y2=0
cc_157 N_A_64_409#_M1004_s N_Y_c_264_n 3.52625e-19 $X=0.32 $Y=2.045 $X2=0 $Y2=0
cc_158 N_A_64_409#_c_206_n N_Y_c_264_n 0.00386824f $X=0.465 $Y=2.44 $X2=0 $Y2=0
cc_159 N_A_64_409#_c_206_n N_Y_c_272_n 0.0289919f $X=0.465 $Y=2.44 $X2=0 $Y2=0
cc_160 N_A_64_409#_c_207_n N_Y_c_272_n 0.0152054f $X=1.36 $Y=2.98 $X2=0 $Y2=0
cc_161 N_A_64_409#_c_216_n N_Y_c_272_n 0.0407863f $X=1.525 $Y=2.19 $X2=0 $Y2=0
cc_162 N_A_64_409#_c_210_n N_VPWR_M1006_d 0.00191634f $X=2.43 $Y=2.01 $X2=-0.19
+ $Y2=1.655
cc_163 N_A_64_409#_c_209_n N_VPWR_c_308_n 0.0119061f $X=1.525 $Y=2.895 $X2=0
+ $Y2=0
cc_164 N_A_64_409#_c_216_n N_VPWR_c_308_n 0.0408193f $X=1.525 $Y=2.19 $X2=0
+ $Y2=0
cc_165 N_A_64_409#_c_210_n N_VPWR_c_308_n 0.0164036f $X=2.43 $Y=2.01 $X2=0 $Y2=0
cc_166 N_A_64_409#_c_212_n N_VPWR_c_308_n 0.0500655f $X=2.595 $Y=2.19 $X2=0
+ $Y2=0
cc_167 N_A_64_409#_c_207_n N_VPWR_c_309_n 0.0429009f $X=1.36 $Y=2.98 $X2=0 $Y2=0
cc_168 N_A_64_409#_c_208_n N_VPWR_c_309_n 0.0221635f $X=0.63 $Y=2.98 $X2=0 $Y2=0
cc_169 N_A_64_409#_c_209_n N_VPWR_c_309_n 0.0220769f $X=1.525 $Y=2.895 $X2=0
+ $Y2=0
cc_170 N_A_64_409#_c_212_n N_VPWR_c_311_n 0.0220321f $X=2.595 $Y=2.19 $X2=0
+ $Y2=0
cc_171 N_A_64_409#_c_207_n N_VPWR_c_307_n 0.0252115f $X=1.36 $Y=2.98 $X2=0 $Y2=0
cc_172 N_A_64_409#_c_208_n N_VPWR_c_307_n 0.0126536f $X=0.63 $Y=2.98 $X2=0 $Y2=0
cc_173 N_A_64_409#_c_209_n N_VPWR_c_307_n 0.0125384f $X=1.525 $Y=2.895 $X2=0
+ $Y2=0
cc_174 N_A_64_409#_c_212_n N_VPWR_c_307_n 0.0125808f $X=2.595 $Y=2.19 $X2=0
+ $Y2=0
cc_175 N_Y_c_259_n N_VGND_c_337_n 0.0222461f $X=1.22 $Y=0.81 $X2=0 $Y2=0
cc_176 N_Y_c_260_n N_VGND_c_337_n 0.00887059f $X=1.385 $Y=0.47 $X2=0 $Y2=0
cc_177 N_Y_c_259_n N_VGND_c_340_n 8.21074e-19 $X=1.22 $Y=0.81 $X2=0 $Y2=0
cc_178 N_Y_c_261_n N_VGND_c_340_n 0.00373548f $X=0.235 $Y=0.895 $X2=0 $Y2=0
cc_179 N_Y_c_259_n N_VGND_c_341_n 0.00697632f $X=1.22 $Y=0.81 $X2=0 $Y2=0
cc_180 N_Y_c_260_n N_VGND_c_341_n 0.0196636f $X=1.385 $Y=0.47 $X2=0 $Y2=0
cc_181 N_Y_M1007_d N_VGND_c_343_n 0.00614092f $X=1.245 $Y=0.235 $X2=0 $Y2=0
cc_182 N_Y_c_259_n N_VGND_c_343_n 0.0146112f $X=1.22 $Y=0.81 $X2=0 $Y2=0
cc_183 N_Y_c_260_n N_VGND_c_343_n 0.0125545f $X=1.385 $Y=0.47 $X2=0 $Y2=0
cc_184 N_Y_c_261_n N_VGND_c_343_n 0.0062458f $X=0.235 $Y=0.895 $X2=0 $Y2=0
cc_185 N_VGND_c_343_n A_171_47# 0.0031085f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_186 N_VGND_c_343_n A_357_47# 0.0180084f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
