* File: sky130_fd_sc_lp__sleep_sergate_plv_21.pxi.spice
* Created: Wed Sep  2 10:38:12 2020
* 
x_PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_21%SLEEP N_SLEEP_c_42_n N_SLEEP_c_43_n
+ N_SLEEP_M1002_g N_SLEEP_c_44_n N_SLEEP_c_45_n N_SLEEP_M1000_g N_SLEEP_c_46_n
+ N_SLEEP_c_47_n N_SLEEP_M1001_g N_SLEEP_c_48_n SLEEP SLEEP SLEEP SLEEP SLEEP
+ N_SLEEP_c_41_n PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_21%SLEEP
x_PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_21%VPWR N_VPWR_M1000_s N_VPWR_M1001_s
+ VPWR N_VPWR_c_104_n N_VPWR_c_105_n N_VPWR_c_106_n N_VPWR_c_107_n
+ N_VPWR_c_108_n N_VPWR_c_109_n N_VPWR_c_110_n N_VPWR_c_103_n
+ PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_21%VPWR
x_PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_21%VIRTPWR N_VIRTPWR_M1000_d
+ N_VIRTPWR_M1002_d N_VIRTPWR_c_206_n N_VIRTPWR_c_207_n VIRTPWR
+ N_VIRTPWR_c_208_n N_VIRTPWR_c_209_n N_VIRTPWR_c_210_n N_VIRTPWR_c_211_n
+ N_VIRTPWR_c_212_n N_VIRTPWR_c_213_n N_VIRTPWR_c_214_n N_VIRTPWR_c_201_n
+ N_VIRTPWR_c_216_n N_VIRTPWR_c_202_n N_VIRTPWR_c_203_n N_VIRTPWR_c_204_n
+ VIRTPWR N_VIRTPWR_c_205_n PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_21%VIRTPWR
cc_1 noxref_1 SLEEP 0.0459532f $X=-0.19 $Y=-0.002 $X2=8.315 $Y2=0.84
cc_2 noxref_1 N_SLEEP_c_41_n 0.028932f $X=-0.19 $Y=-0.002 $X2=8.42 $Y2=1.535
cc_3 noxref_1 N_VPWR_c_103_n 0.618373f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_4 noxref_1 VIRTPWR 0.105802f $X=-0.19 $Y=-0.002 $X2=4.555 $Y2=2.325
cc_5 noxref_1 N_VIRTPWR_c_201_n 0.0836651f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_6 noxref_1 N_VIRTPWR_c_202_n 0.0786895f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_7 noxref_1 N_VIRTPWR_c_203_n 0.0386646f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_8 noxref_1 N_VIRTPWR_c_204_n 0.0386646f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_9 noxref_1 N_VIRTPWR_c_205_n 0.0386646f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_10 VPB N_SLEEP_c_42_n 0.0188377f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.25
cc_11 VPB N_SLEEP_c_43_n 0.0317437f $X=-0.19 $Y=1.655 $X2=8.13 $Y2=2.755
cc_12 VPB N_SLEEP_c_44_n 0.0423621f $X=-0.19 $Y=1.655 $X2=8.205 $Y2=1.895
cc_13 VPB N_SLEEP_c_45_n 0.0139468f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.895
cc_14 VPB N_SLEEP_c_46_n 0.0149312f $X=-0.19 $Y=1.655 $X2=8.13 $Y2=2.325
cc_15 VPB N_SLEEP_c_47_n 0.0125894f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.325
cc_16 VPB N_SLEEP_c_48_n 0.0161409f $X=-0.19 $Y=1.655 $X2=8.205 $Y2=2.68
cc_17 VPB SLEEP 0.0360919f $X=-0.19 $Y=1.655 $X2=8.315 $Y2=0.84
cc_18 VPB N_SLEEP_c_41_n 0.0304926f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=1.535
cc_19 VPB N_VPWR_c_104_n 0.0994951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_20 VPB N_VPWR_c_105_n 0.00214921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_21 VPB N_VPWR_c_106_n 0.0155703f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_107_n 0.00821471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_23 VPB N_VPWR_c_108_n 0.00821471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_109_n 0.00821471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 VPB N_VPWR_c_110_n 0.00821471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_VPWR_c_103_n 0.115514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_VIRTPWR_c_206_n 0.0130323f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.895
cc_28 VPB N_VIRTPWR_c_207_n 0.0357155f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.325
cc_29 VPB N_VIRTPWR_c_208_n 0.15875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VIRTPWR_c_209_n 0.00789876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VIRTPWR_c_210_n 0.00789876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VIRTPWR_c_211_n 0.00789876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VIRTPWR_c_212_n 0.00815152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VIRTPWR_c_213_n 0.00214921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_VIRTPWR_c_214_n 0.0329627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VIRTPWR_c_201_n 0.0405705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VIRTPWR_c_216_n 0.0130323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VIRTPWR_c_202_n 0.0404102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 N_SLEEP_c_44_n N_VPWR_c_104_n 0.0112707f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_40 SLEEP N_VPWR_c_104_n 0.0112305f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_41 N_SLEEP_c_41_n N_VPWR_c_104_n 0.0049252f $X=8.42 $Y=1.535 $X2=0 $Y2=0
cc_42 N_SLEEP_c_43_n N_VPWR_c_105_n 0.010275f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_43 N_SLEEP_c_46_n N_VPWR_c_105_n 0.0102402f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_44 N_SLEEP_c_48_n N_VPWR_c_105_n 0.00197123f $X=8.205 $Y=2.68 $X2=0 $Y2=0
cc_45 SLEEP N_VPWR_c_105_n 0.0107074f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_46 N_SLEEP_c_43_n N_VPWR_c_106_n 0.00303147f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_47 N_SLEEP_c_44_n N_VPWR_c_106_n 0.00419339f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_48 N_SLEEP_c_46_n N_VPWR_c_106_n 0.00352159f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_49 N_SLEEP_c_44_n N_VPWR_c_107_n 0.00101546f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_50 N_SLEEP_c_46_n N_VPWR_c_107_n 0.00101546f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_51 N_SLEEP_c_44_n N_VPWR_c_108_n 0.00101546f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_52 N_SLEEP_c_46_n N_VPWR_c_108_n 0.00101546f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_53 N_SLEEP_c_44_n N_VPWR_c_109_n 0.00101546f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_54 N_SLEEP_c_46_n N_VPWR_c_109_n 0.00101546f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_55 N_SLEEP_c_44_n N_VPWR_c_110_n 0.0034209f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_56 N_SLEEP_c_46_n N_VPWR_c_110_n 0.00285945f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_57 SLEEP N_VPWR_c_110_n 0.0204982f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_58 N_SLEEP_c_41_n N_VPWR_c_110_n 2.24623e-19 $X=8.42 $Y=1.535 $X2=0 $Y2=0
cc_59 N_SLEEP_c_42_n N_VPWR_c_103_n 0.00351535f $X=0.905 $Y=2.25 $X2=0 $Y2=0
cc_60 N_SLEEP_c_43_n N_VPWR_c_103_n 0.00708282f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_61 N_SLEEP_c_44_n N_VPWR_c_103_n 0.00542344f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_62 N_SLEEP_c_45_n N_VPWR_c_103_n 0.00314945f $X=0.98 $Y=1.895 $X2=0 $Y2=0
cc_63 N_SLEEP_c_46_n N_VPWR_c_103_n 0.00225492f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_64 N_SLEEP_c_47_n N_VPWR_c_103_n 0.00269623f $X=0.98 $Y=2.325 $X2=0 $Y2=0
cc_65 N_SLEEP_c_48_n N_VPWR_c_103_n 0.00108676f $X=8.205 $Y=2.68 $X2=0 $Y2=0
cc_66 SLEEP N_VPWR_c_103_n 0.0998334f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_67 N_SLEEP_c_41_n N_VPWR_c_103_n 0.00592277f $X=8.42 $Y=1.535 $X2=0 $Y2=0
cc_68 N_SLEEP_c_43_n N_VIRTPWR_c_206_n 0.0158929f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_69 N_SLEEP_c_43_n N_VIRTPWR_c_207_n 0.00259154f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_70 N_SLEEP_c_43_n N_VIRTPWR_c_209_n 0.00539584f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_71 N_SLEEP_c_44_n N_VIRTPWR_c_209_n 0.00101539f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_72 N_SLEEP_c_46_n N_VIRTPWR_c_209_n 0.00101539f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_73 N_SLEEP_c_43_n N_VIRTPWR_c_210_n 0.00539584f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_74 N_SLEEP_c_44_n N_VIRTPWR_c_210_n 0.00101539f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_75 N_SLEEP_c_46_n N_VIRTPWR_c_210_n 0.00101539f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_76 N_SLEEP_c_43_n N_VIRTPWR_c_211_n 0.00539584f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_77 N_SLEEP_c_44_n N_VIRTPWR_c_211_n 0.00101539f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_78 N_SLEEP_c_46_n N_VIRTPWR_c_211_n 0.00101539f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_79 N_SLEEP_c_43_n N_VIRTPWR_c_212_n 0.00539734f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_80 N_SLEEP_c_44_n N_VIRTPWR_c_212_n 0.00101545f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_81 N_SLEEP_c_46_n N_VIRTPWR_c_212_n 0.00101545f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_82 N_SLEEP_c_42_n N_VIRTPWR_c_213_n 0.00374504f $X=0.905 $Y=2.25 $X2=0 $Y2=0
cc_83 N_SLEEP_c_44_n N_VIRTPWR_c_213_n 0.0113049f $X=8.205 $Y=1.895 $X2=0 $Y2=0
cc_84 N_SLEEP_c_46_n N_VIRTPWR_c_213_n 0.0102402f $X=8.13 $Y=2.325 $X2=0 $Y2=0
cc_85 SLEEP N_VIRTPWR_c_213_n 0.0115213f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_86 N_SLEEP_c_43_n N_VIRTPWR_c_214_n 0.00439978f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_87 SLEEP N_VIRTPWR_c_214_n 0.017839f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_88 N_SLEEP_c_43_n N_VIRTPWR_c_201_n 0.00379335f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_89 SLEEP N_VIRTPWR_c_201_n 0.0126174f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_90 N_SLEEP_c_43_n N_VIRTPWR_c_202_n 0.00224979f $X=8.13 $Y=2.755 $X2=0 $Y2=0
cc_91 N_VPWR_c_106_n N_VIRTPWR_M1000_d 3.18208e-19 $X=1.545 $Y=1.68 $X2=-0.19
+ $Y2=-0.002
cc_92 N_VPWR_c_110_n N_VIRTPWR_M1000_d 2.87889e-19 $X=7.775 $Y=1.68 $X2=-0.19
+ $Y2=-0.002
cc_93 N_VPWR_c_105_n N_VIRTPWR_c_206_n 0.262559f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_94 N_VPWR_c_106_n N_VIRTPWR_c_206_n 0.00580238f $X=1.545 $Y=1.68 $X2=0 $Y2=0
cc_95 N_VPWR_c_103_n N_VIRTPWR_c_206_n 0.00611837f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_96 N_VPWR_c_103_n VIRTPWR 0.224849f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_97 N_VPWR_c_107_n N_VIRTPWR_c_208_n 0.00708574f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_98 N_VPWR_c_108_n N_VIRTPWR_c_208_n 0.00708574f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_99 N_VPWR_c_109_n N_VIRTPWR_c_208_n 0.00708574f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_100 N_VPWR_c_110_n N_VIRTPWR_c_208_n 0.00580238f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_101 N_VPWR_c_103_n N_VIRTPWR_c_208_n 0.0186573f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_102 N_VPWR_M1001_s N_VIRTPWR_c_209_n 2.87738e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_103 N_VPWR_c_104_n N_VIRTPWR_c_209_n 0.0389016f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_104 N_VPWR_c_105_n N_VIRTPWR_c_209_n 0.0346616f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_105 N_VPWR_c_106_n N_VIRTPWR_c_209_n 0.0970367f $X=1.545 $Y=1.68 $X2=0 $Y2=0
cc_106 N_VPWR_c_107_n N_VIRTPWR_c_209_n 0.0970367f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_107 N_VPWR_c_103_n N_VIRTPWR_c_209_n 0.219944f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_108 N_VPWR_M1001_s N_VIRTPWR_c_210_n 2.87738e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_109 N_VPWR_c_104_n N_VIRTPWR_c_210_n 0.0389016f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_110 N_VPWR_c_105_n N_VIRTPWR_c_210_n 0.0346616f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_111 N_VPWR_c_107_n N_VIRTPWR_c_210_n 0.0970367f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_112 N_VPWR_c_108_n N_VIRTPWR_c_210_n 0.0970367f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_113 N_VPWR_c_103_n N_VIRTPWR_c_210_n 0.219944f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_114 N_VPWR_M1001_s N_VIRTPWR_c_211_n 2.87738e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_115 N_VPWR_c_104_n N_VIRTPWR_c_211_n 0.0389016f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_116 N_VPWR_c_105_n N_VIRTPWR_c_211_n 0.0346616f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_117 N_VPWR_c_108_n N_VIRTPWR_c_211_n 0.0970367f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_118 N_VPWR_c_109_n N_VIRTPWR_c_211_n 0.0970367f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_119 N_VPWR_c_103_n N_VIRTPWR_c_211_n 0.219944f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_120 N_VPWR_M1001_s N_VIRTPWR_c_212_n 2.8786e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_121 N_VPWR_c_104_n N_VIRTPWR_c_212_n 0.0400253f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_122 N_VPWR_c_105_n N_VIRTPWR_c_212_n 0.0356496f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_123 N_VPWR_c_109_n N_VIRTPWR_c_212_n 0.0970546f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_124 N_VPWR_c_110_n N_VIRTPWR_c_212_n 0.0970546f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_125 N_VPWR_c_103_n N_VIRTPWR_c_212_n 0.225341f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_126 N_VPWR_c_104_n N_VIRTPWR_c_213_n 0.251237f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_127 N_VPWR_c_105_n N_VIRTPWR_c_213_n 0.251237f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_128 N_VPWR_c_106_n N_VIRTPWR_c_213_n 0.0377876f $X=1.545 $Y=1.68 $X2=0 $Y2=0
cc_129 N_VPWR_c_107_n N_VIRTPWR_c_213_n 0.0358966f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_130 N_VPWR_c_108_n N_VIRTPWR_c_213_n 0.0358966f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_131 N_VPWR_c_109_n N_VIRTPWR_c_213_n 0.0358966f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_132 N_VPWR_c_110_n N_VIRTPWR_c_213_n 0.0393669f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_133 N_VPWR_c_103_n N_VIRTPWR_c_213_n 0.0173287f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_134 N_VPWR_c_105_n N_VIRTPWR_c_201_n 0.00290716f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_135 N_VPWR_c_110_n N_VIRTPWR_c_201_n 0.026124f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_136 N_VPWR_c_103_n N_VIRTPWR_c_201_n 0.227442f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_137 N_VPWR_c_103_n N_VIRTPWR_c_216_n 0.00787277f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_138 N_VPWR_c_105_n N_VIRTPWR_c_202_n 0.00285709f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_139 N_VPWR_c_106_n N_VIRTPWR_c_202_n 0.026124f $X=1.545 $Y=1.68 $X2=0 $Y2=0
cc_140 N_VPWR_c_103_n N_VIRTPWR_c_202_n 0.212348f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_141 N_VPWR_c_105_n N_VIRTPWR_c_203_n 0.0012824f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_142 N_VPWR_c_107_n N_VIRTPWR_c_203_n 0.0229031f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_143 N_VPWR_c_103_n N_VIRTPWR_c_203_n 0.0980574f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_144 N_VPWR_c_105_n N_VIRTPWR_c_204_n 0.0012824f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_145 N_VPWR_c_108_n N_VIRTPWR_c_204_n 0.0229031f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_146 N_VPWR_c_103_n N_VIRTPWR_c_204_n 0.0980574f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_147 N_VPWR_c_105_n N_VIRTPWR_c_205_n 0.0012824f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_148 N_VPWR_c_109_n N_VIRTPWR_c_205_n 0.0229031f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_149 N_VPWR_c_103_n N_VIRTPWR_c_205_n 0.0980574f $X=7.775 $Y=1.68 $X2=0 $Y2=0
