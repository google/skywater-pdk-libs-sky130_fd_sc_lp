# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__nor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.185000 1.160000 1.515000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.670000 1.345000 1.870000 1.605000 ;
        RECT 1.670000 1.605000 3.745000 1.785000 ;
        RECT 2.940000 1.285000 3.745000 1.605000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.040000 1.210000 2.760000 1.435000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.117200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 0.255000 1.175000 0.840000 ;
        RECT 0.965000 0.840000 2.980000 1.015000 ;
        RECT 1.330000 1.015000 2.980000 1.040000 ;
        RECT 1.330000 1.040000 1.500000 1.965000 ;
        RECT 1.330000 1.965000 2.505000 2.295000 ;
        RECT 1.845000 0.255000 2.085000 0.840000 ;
        RECT 2.755000 0.255000 2.980000 0.840000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.140000  1.685000 1.160000 1.855000 ;
      RECT 0.140000  1.855000 0.410000 3.075000 ;
      RECT 0.465000  0.085000 0.795000 1.015000 ;
      RECT 0.580000  2.025000 0.820000 2.815000 ;
      RECT 0.580000  2.815000 1.245000 3.245000 ;
      RECT 0.990000  1.855000 1.160000 2.465000 ;
      RECT 0.990000  2.465000 2.845000 2.645000 ;
      RECT 1.345000  0.085000 1.675000 0.670000 ;
      RECT 1.415000  2.645000 1.605000 3.075000 ;
      RECT 1.775000  2.815000 3.315000 3.075000 ;
      RECT 2.255000  0.085000 2.585000 0.670000 ;
      RECT 2.675000  1.955000 3.745000 2.125000 ;
      RECT 2.675000  2.125000 2.845000 2.465000 ;
      RECT 3.015000  2.295000 3.315000 2.815000 ;
      RECT 3.150000  0.085000 3.445000 1.095000 ;
      RECT 3.485000  2.125000 3.745000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__nor3_2
END LIBRARY
