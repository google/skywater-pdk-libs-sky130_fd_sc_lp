* File: sky130_fd_sc_lp__nor4b_lp.pxi.spice
* Created: Wed Sep  2 10:11:16 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4B_LP%D_N N_D_N_c_86_n N_D_N_M1013_g N_D_N_c_87_n
+ N_D_N_M1009_g N_D_N_c_88_n N_D_N_c_89_n N_D_N_M1006_g N_D_N_c_95_n
+ N_D_N_c_90_n D_N D_N N_D_N_c_92_n N_D_N_c_93_n
+ PM_SKY130_FD_SC_LP__NOR4B_LP%D_N
x_PM_SKY130_FD_SC_LP__NOR4B_LP%A_31_409# N_A_31_409#_M1009_s N_A_31_409#_M1013_s
+ N_A_31_409#_c_138_n N_A_31_409#_M1011_g N_A_31_409#_c_148_n
+ N_A_31_409#_c_149_n N_A_31_409#_M1010_g N_A_31_409#_c_151_n
+ N_A_31_409#_c_152_n N_A_31_409#_M1008_g N_A_31_409#_c_153_n
+ N_A_31_409#_c_141_n N_A_31_409#_c_154_n N_A_31_409#_c_155_n
+ N_A_31_409#_c_142_n N_A_31_409#_c_143_n N_A_31_409#_c_144_n
+ N_A_31_409#_c_145_n N_A_31_409#_c_146_n PM_SKY130_FD_SC_LP__NOR4B_LP%A_31_409#
x_PM_SKY130_FD_SC_LP__NOR4B_LP%C N_C_M1003_g N_C_c_222_n N_C_c_223_n N_C_M1005_g
+ N_C_M1014_g C C C C N_C_c_225_n N_C_c_226_n PM_SKY130_FD_SC_LP__NOR4B_LP%C
x_PM_SKY130_FD_SC_LP__NOR4B_LP%B N_B_c_271_n N_B_M1000_g N_B_c_272_n N_B_c_273_n
+ N_B_c_274_n N_B_M1012_g N_B_M1004_g N_B_c_275_n N_B_c_276_n N_B_c_277_n
+ N_B_c_282_n B B B B N_B_c_278_n N_B_c_279_n PM_SKY130_FD_SC_LP__NOR4B_LP%B
x_PM_SKY130_FD_SC_LP__NOR4B_LP%A N_A_c_332_n N_A_M1007_g N_A_c_338_n N_A_M1001_g
+ N_A_M1002_g N_A_c_333_n N_A_c_334_n N_A_c_335_n A A N_A_c_337_n
+ PM_SKY130_FD_SC_LP__NOR4B_LP%A
x_PM_SKY130_FD_SC_LP__NOR4B_LP%VPWR N_VPWR_M1013_d N_VPWR_M1001_d N_VPWR_c_370_n
+ N_VPWR_c_371_n N_VPWR_c_372_n VPWR N_VPWR_c_373_n N_VPWR_c_374_n
+ N_VPWR_c_369_n PM_SKY130_FD_SC_LP__NOR4B_LP%VPWR
x_PM_SKY130_FD_SC_LP__NOR4B_LP%Y N_Y_M1010_d N_Y_M1012_d N_Y_M1008_s N_Y_c_404_n
+ N_Y_c_405_n N_Y_c_406_n Y Y Y Y Y Y Y N_Y_c_408_n
+ PM_SKY130_FD_SC_LP__NOR4B_LP%Y
x_PM_SKY130_FD_SC_LP__NOR4B_LP%VGND N_VGND_M1006_d N_VGND_M1005_d N_VGND_M1002_d
+ N_VGND_c_466_n N_VGND_c_467_n N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n
+ N_VGND_c_471_n VGND N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n
+ N_VGND_c_475_n PM_SKY130_FD_SC_LP__NOR4B_LP%VGND
cc_1 VNB N_D_N_c_86_n 0.0220255f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.658
cc_2 VNB N_D_N_c_87_n 0.0175316f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.78
cc_3 VNB N_D_N_c_88_n 0.0171406f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.855
cc_4 VNB N_D_N_c_89_n 0.0138865f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.78
cc_5 VNB N_D_N_c_90_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.855
cc_6 VNB D_N 0.00478821f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_D_N_c_92_n 0.0188288f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.34
cc_8 VNB N_D_N_c_93_n 0.0177994f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.175
cc_9 VNB N_A_31_409#_c_138_n 0.0206189f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.495
cc_10 VNB N_A_31_409#_M1011_g 0.034433f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.175
cc_11 VNB N_A_31_409#_M1010_g 0.0528215f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.845
cc_12 VNB N_A_31_409#_c_141_n 0.0285332f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.295
cc_13 VNB N_A_31_409#_c_142_n 0.0108515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_31_409#_c_143_n 0.0021381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_31_409#_c_144_n 0.0268475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_31_409#_c_145_n 0.0150782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_31_409#_c_146_n 0.0312812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C_M1003_g 0.0305029f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.845
cc_19 VNB N_C_c_222_n 0.00900967f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.545
cc_20 VNB N_C_c_223_n 0.00709894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C_M1005_g 0.0413679f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.495
cc_22 VNB N_C_c_225_n 0.0568188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_c_226_n 0.00974444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_271_n 0.0149554f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.362
cc_25 VNB N_B_c_272_n 0.0102086f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.545
cc_26 VNB N_B_c_273_n 0.00879346f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.545
cc_27 VNB N_B_c_274_n 0.0137589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_275_n 0.00437176f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.495
cc_29 VNB N_B_c_276_n 0.0218753f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.845
cc_30 VNB N_B_c_277_n 0.019964f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.855
cc_31 VNB N_B_c_278_n 0.0173748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_c_279_n 0.00188741f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.665
cc_33 VNB N_A_c_332_n 0.0372957f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.362
cc_34 VNB N_A_c_333_n 0.0258162f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.78
cc_35 VNB N_A_c_334_n 0.0192733f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.495
cc_36 VNB N_A_c_335_n 0.00443853f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.845
cc_37 VNB A 0.0440991f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_38 VNB N_A_c_337_n 0.0343734f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.295
cc_39 VNB N_VPWR_c_369_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_404_n 0.0293526f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.93
cc_41 VNB N_Y_c_405_n 0.00129592f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.855
cc_42 VNB N_Y_c_406_n 0.00635637f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.495
cc_43 VNB Y 0.00846983f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_44 VNB N_Y_c_408_n 0.00651903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_466_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.855
cc_46 VNB N_VGND_c_467_n 0.00422339f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.495
cc_47 VNB N_VGND_c_468_n 0.0121802f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.855
cc_48 VNB N_VGND_c_469_n 0.0250343f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_49 VNB N_VGND_c_470_n 0.0330554f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.34
cc_50 VNB N_VGND_c_471_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.34
cc_51 VNB N_VGND_c_472_n 0.0307725f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.295
cc_52 VNB N_VGND_c_473_n 0.0386751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_474_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_475_n 0.290396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VPB N_D_N_M1013_g 0.038348f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.545
cc_56 VPB N_D_N_c_95_n 0.0176732f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.845
cc_57 VPB D_N 0.00266092f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_58 VPB N_A_31_409#_c_138_n 0.0105549f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=0.495
cc_59 VPB N_A_31_409#_c_148_n 0.0137758f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.855
cc_60 VPB N_A_31_409#_c_149_n 0.0355825f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.78
cc_61 VPB N_A_31_409#_M1010_g 0.00723352f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.845
cc_62 VPB N_A_31_409#_c_151_n 0.0484887f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_63 VPB N_A_31_409#_c_152_n 0.0248509f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_31_409#_c_153_n 0.00666874f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.34
cc_65 VPB N_A_31_409#_c_154_n 0.0118411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_31_409#_c_155_n 0.035517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_31_409#_c_146_n 0.0173555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_C_M1014_g 0.0360647f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.855
cc_69 VPB N_C_c_225_n 0.0010012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_C_c_226_n 0.00348261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_B_M1004_g 0.0253187f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.855
cc_72 VPB N_B_c_277_n 0.00452214f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=0.855
cc_73 VPB N_B_c_282_n 0.013931f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_74 VPB N_B_c_279_n 0.00171813f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.665
cc_75 VPB N_A_c_338_n 0.0407652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_c_335_n 0.00978284f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.845
cc_77 VPB A 0.0173577f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_78 VPB N_VPWR_c_370_n 0.0292045f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.175
cc_79 VPB N_VPWR_c_371_n 0.0159821f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.495
cc_80 VPB N_VPWR_c_372_n 0.0470929f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.845
cc_81 VPB N_VPWR_c_373_n 0.0875541f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.34
cc_82 VPB N_VPWR_c_374_n 0.0250488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_369_n 0.108421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB Y 0.045421f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_85 N_D_N_c_86_n N_A_31_409#_c_138_n 0.0121713f $X=0.627 $Y=1.658 $X2=0 $Y2=0
cc_86 N_D_N_c_89_n N_A_31_409#_M1011_g 0.018891f $X=1.005 $Y=0.78 $X2=0 $Y2=0
cc_87 N_D_N_c_93_n N_A_31_409#_M1011_g 0.00283511f $X=0.627 $Y=1.175 $X2=0 $Y2=0
cc_88 N_D_N_M1013_g N_A_31_409#_c_149_n 0.00420194f $X=0.565 $Y=2.545 $X2=0
+ $Y2=0
cc_89 N_D_N_c_95_n N_A_31_409#_c_149_n 0.0121713f $X=0.627 $Y=1.845 $X2=0 $Y2=0
cc_90 N_D_N_c_87_n N_A_31_409#_c_141_n 0.011359f $X=0.645 $Y=0.78 $X2=0 $Y2=0
cc_91 N_D_N_c_89_n N_A_31_409#_c_141_n 0.00170023f $X=1.005 $Y=0.78 $X2=0 $Y2=0
cc_92 N_D_N_c_90_n N_A_31_409#_c_141_n 0.00311141f $X=0.645 $Y=0.855 $X2=0 $Y2=0
cc_93 N_D_N_M1013_g N_A_31_409#_c_154_n 0.00451956f $X=0.565 $Y=2.545 $X2=0
+ $Y2=0
cc_94 N_D_N_M1013_g N_A_31_409#_c_155_n 0.015872f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_95 N_D_N_c_88_n N_A_31_409#_c_142_n 0.0171046f $X=0.93 $Y=0.855 $X2=0 $Y2=0
cc_96 N_D_N_c_90_n N_A_31_409#_c_142_n 0.00407103f $X=0.645 $Y=0.855 $X2=0 $Y2=0
cc_97 D_N N_A_31_409#_c_142_n 0.0178482f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_98 N_D_N_c_92_n N_A_31_409#_c_142_n 2.90584e-19 $X=0.65 $Y=1.34 $X2=0 $Y2=0
cc_99 N_D_N_c_93_n N_A_31_409#_c_142_n 0.00373203f $X=0.627 $Y=1.175 $X2=0 $Y2=0
cc_100 D_N N_A_31_409#_c_143_n 0.0438819f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_101 N_D_N_c_92_n N_A_31_409#_c_143_n 8.21899e-19 $X=0.65 $Y=1.34 $X2=0 $Y2=0
cc_102 N_D_N_c_93_n N_A_31_409#_c_143_n 0.00392528f $X=0.627 $Y=1.175 $X2=0
+ $Y2=0
cc_103 N_D_N_c_88_n N_A_31_409#_c_144_n 0.0013606f $X=0.93 $Y=0.855 $X2=0 $Y2=0
cc_104 D_N N_A_31_409#_c_144_n 0.00428486f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_105 N_D_N_c_92_n N_A_31_409#_c_144_n 0.0121713f $X=0.65 $Y=1.34 $X2=0 $Y2=0
cc_106 N_D_N_c_90_n N_A_31_409#_c_145_n 0.00254537f $X=0.645 $Y=0.855 $X2=0
+ $Y2=0
cc_107 D_N N_A_31_409#_c_145_n 0.0091809f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_108 N_D_N_c_92_n N_A_31_409#_c_145_n 0.00285405f $X=0.65 $Y=1.34 $X2=0 $Y2=0
cc_109 N_D_N_c_93_n N_A_31_409#_c_145_n 0.00192368f $X=0.627 $Y=1.175 $X2=0
+ $Y2=0
cc_110 D_N N_A_31_409#_c_146_n 0.0483739f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_111 N_D_N_c_92_n N_A_31_409#_c_146_n 0.020953f $X=0.65 $Y=1.34 $X2=0 $Y2=0
cc_112 N_D_N_c_93_n N_A_31_409#_c_146_n 0.00400465f $X=0.627 $Y=1.175 $X2=0
+ $Y2=0
cc_113 N_D_N_M1013_g N_VPWR_c_370_n 0.0249766f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_114 N_D_N_c_95_n N_VPWR_c_370_n 9.71359e-19 $X=0.627 $Y=1.845 $X2=0 $Y2=0
cc_115 D_N N_VPWR_c_370_n 0.0143035f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_116 N_D_N_M1013_g N_VPWR_c_374_n 0.00769046f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_117 N_D_N_M1013_g N_VPWR_c_369_n 0.014097f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_118 N_D_N_c_87_n N_VGND_c_466_n 0.00189426f $X=0.645 $Y=0.78 $X2=0 $Y2=0
cc_119 N_D_N_c_89_n N_VGND_c_466_n 0.0106297f $X=1.005 $Y=0.78 $X2=0 $Y2=0
cc_120 N_D_N_c_87_n N_VGND_c_472_n 0.00502664f $X=0.645 $Y=0.78 $X2=0 $Y2=0
cc_121 N_D_N_c_88_n N_VGND_c_472_n 4.57848e-19 $X=0.93 $Y=0.855 $X2=0 $Y2=0
cc_122 N_D_N_c_89_n N_VGND_c_472_n 0.00445056f $X=1.005 $Y=0.78 $X2=0 $Y2=0
cc_123 N_D_N_c_87_n N_VGND_c_475_n 0.00635263f $X=0.645 $Y=0.78 $X2=0 $Y2=0
cc_124 N_D_N_c_88_n N_VGND_c_475_n 6.33118e-19 $X=0.93 $Y=0.855 $X2=0 $Y2=0
cc_125 N_D_N_c_89_n N_VGND_c_475_n 0.00417935f $X=1.005 $Y=0.78 $X2=0 $Y2=0
cc_126 N_A_31_409#_M1010_g N_C_M1003_g 0.0375457f $X=1.825 $Y=0.495 $X2=0 $Y2=0
cc_127 N_A_31_409#_c_151_n N_C_c_223_n 0.0121119f $X=2.435 $Y=1.86 $X2=0 $Y2=0
cc_128 N_A_31_409#_c_151_n N_C_M1014_g 0.0778064f $X=2.435 $Y=1.86 $X2=0 $Y2=0
cc_129 N_A_31_409#_M1010_g N_C_c_225_n 0.00214073f $X=1.825 $Y=0.495 $X2=0 $Y2=0
cc_130 N_A_31_409#_c_151_n N_C_c_225_n 0.00803981f $X=2.435 $Y=1.86 $X2=0 $Y2=0
cc_131 N_A_31_409#_M1010_g N_C_c_226_n 0.00121299f $X=1.825 $Y=0.495 $X2=0 $Y2=0
cc_132 N_A_31_409#_c_151_n N_C_c_226_n 0.00780042f $X=2.435 $Y=1.86 $X2=0 $Y2=0
cc_133 N_A_31_409#_c_152_n N_C_c_226_n 0.0339935f $X=2.56 $Y=1.935 $X2=0 $Y2=0
cc_134 N_A_31_409#_c_154_n N_VPWR_c_370_n 0.0684934f $X=0.3 $Y=2.19 $X2=0 $Y2=0
cc_135 N_A_31_409#_c_152_n N_VPWR_c_373_n 0.00703646f $X=2.56 $Y=1.935 $X2=0
+ $Y2=0
cc_136 N_A_31_409#_c_155_n N_VPWR_c_374_n 0.0220321f $X=0.3 $Y=2.9 $X2=0 $Y2=0
cc_137 N_A_31_409#_c_152_n N_VPWR_c_369_n 0.0118134f $X=2.56 $Y=1.935 $X2=0
+ $Y2=0
cc_138 N_A_31_409#_c_155_n N_VPWR_c_369_n 0.0125808f $X=0.3 $Y=2.9 $X2=0 $Y2=0
cc_139 N_A_31_409#_M1011_g Y 0.0064397f $X=1.435 $Y=0.495 $X2=0 $Y2=0
cc_140 N_A_31_409#_c_148_n Y 0.0138667f $X=1.75 $Y=1.86 $X2=0 $Y2=0
cc_141 N_A_31_409#_M1010_g Y 0.0283359f $X=1.825 $Y=0.495 $X2=0 $Y2=0
cc_142 N_A_31_409#_c_151_n Y 0.0284074f $X=2.435 $Y=1.86 $X2=0 $Y2=0
cc_143 N_A_31_409#_c_152_n Y 0.0316177f $X=2.56 $Y=1.935 $X2=0 $Y2=0
cc_144 N_A_31_409#_c_153_n Y 0.00588934f $X=1.825 $Y=1.86 $X2=0 $Y2=0
cc_145 N_A_31_409#_c_143_n Y 0.0647237f $X=1.22 $Y=1.34 $X2=0 $Y2=0
cc_146 N_A_31_409#_M1011_g N_Y_c_408_n 0.00679776f $X=1.435 $Y=0.495 $X2=0 $Y2=0
cc_147 N_A_31_409#_M1010_g N_Y_c_408_n 0.0221824f $X=1.825 $Y=0.495 $X2=0 $Y2=0
cc_148 N_A_31_409#_c_142_n N_Y_c_408_n 0.0145092f $X=1.055 $Y=0.91 $X2=0 $Y2=0
cc_149 N_A_31_409#_c_143_n N_Y_c_408_n 0.00319463f $X=1.22 $Y=1.34 $X2=0 $Y2=0
cc_150 N_A_31_409#_M1011_g N_VGND_c_466_n 0.00960025f $X=1.435 $Y=0.495 $X2=0
+ $Y2=0
cc_151 N_A_31_409#_M1010_g N_VGND_c_466_n 0.00148359f $X=1.825 $Y=0.495 $X2=0
+ $Y2=0
cc_152 N_A_31_409#_c_141_n N_VGND_c_466_n 0.0130451f $X=0.43 $Y=0.495 $X2=0
+ $Y2=0
cc_153 N_A_31_409#_c_142_n N_VGND_c_466_n 0.0226848f $X=1.055 $Y=0.91 $X2=0
+ $Y2=0
cc_154 N_A_31_409#_c_144_n N_VGND_c_466_n 8.8109e-19 $X=1.22 $Y=1.34 $X2=0 $Y2=0
cc_155 N_A_31_409#_M1011_g N_VGND_c_470_n 0.00445056f $X=1.435 $Y=0.495 $X2=0
+ $Y2=0
cc_156 N_A_31_409#_M1010_g N_VGND_c_470_n 0.00352123f $X=1.825 $Y=0.495 $X2=0
+ $Y2=0
cc_157 N_A_31_409#_c_141_n N_VGND_c_472_n 0.0307973f $X=0.43 $Y=0.495 $X2=0
+ $Y2=0
cc_158 N_A_31_409#_M1011_g N_VGND_c_475_n 0.00802306f $X=1.435 $Y=0.495 $X2=0
+ $Y2=0
cc_159 N_A_31_409#_M1010_g N_VGND_c_475_n 0.00496368f $X=1.825 $Y=0.495 $X2=0
+ $Y2=0
cc_160 N_A_31_409#_c_141_n N_VGND_c_475_n 0.0176109f $X=0.43 $Y=0.495 $X2=0
+ $Y2=0
cc_161 N_A_31_409#_c_142_n N_VGND_c_475_n 0.0147838f $X=1.055 $Y=0.91 $X2=0
+ $Y2=0
cc_162 N_C_M1005_g N_B_c_271_n 0.0187739f $X=2.615 $Y=0.495 $X2=-0.19 $Y2=-0.245
cc_163 N_C_c_225_n N_B_c_273_n 0.00220278f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_164 N_C_c_226_n N_B_c_273_n 7.52211e-19 $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_165 N_C_c_225_n N_B_c_277_n 0.0437589f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_166 N_C_M1014_g N_B_c_282_n 0.0437589f $X=3.05 $Y=2.545 $X2=0 $Y2=0
cc_167 N_C_c_225_n N_B_c_278_n 0.0109285f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_168 N_C_c_226_n N_B_c_278_n 0.0111753f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_169 N_C_c_225_n N_B_c_279_n 0.00185191f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_170 N_C_c_226_n N_B_c_279_n 0.133576f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_171 N_C_M1014_g N_VPWR_c_373_n 0.00595064f $X=3.05 $Y=2.545 $X2=0 $Y2=0
cc_172 N_C_c_226_n N_VPWR_c_373_n 0.0192058f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_173 N_C_M1014_g N_VPWR_c_369_n 0.00758588f $X=3.05 $Y=2.545 $X2=0 $Y2=0
cc_174 N_C_c_226_n N_VPWR_c_369_n 0.0226334f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_175 N_C_c_222_n N_Y_c_404_n 0.00101607f $X=2.54 $Y=1.29 $X2=0 $Y2=0
cc_176 N_C_M1005_g N_Y_c_404_n 0.0153478f $X=2.615 $Y=0.495 $X2=0 $Y2=0
cc_177 N_C_c_225_n N_Y_c_404_n 0.00278281f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_178 N_C_c_226_n N_Y_c_404_n 0.0542952f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_179 N_C_M1003_g Y 0.00487176f $X=2.255 $Y=0.495 $X2=0 $Y2=0
cc_180 N_C_c_222_n Y 0.00264064f $X=2.54 $Y=1.29 $X2=0 $Y2=0
cc_181 N_C_c_223_n Y 0.00634336f $X=2.33 $Y=1.29 $X2=0 $Y2=0
cc_182 N_C_M1005_g Y 0.00464914f $X=2.615 $Y=0.495 $X2=0 $Y2=0
cc_183 N_C_c_225_n Y 0.00170895f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_184 N_C_c_226_n Y 0.141227f $X=2.705 $Y=1.38 $X2=0 $Y2=0
cc_185 N_C_M1003_g N_Y_c_408_n 0.0200398f $X=2.255 $Y=0.495 $X2=0 $Y2=0
cc_186 N_C_M1005_g N_Y_c_408_n 0.00532076f $X=2.615 $Y=0.495 $X2=0 $Y2=0
cc_187 N_C_c_226_n A_537_409# 0.00175001f $X=2.705 $Y=1.38 $X2=-0.19 $Y2=-0.245
cc_188 N_C_c_226_n A_635_409# 0.00757755f $X=2.705 $Y=1.38 $X2=-0.19 $Y2=-0.245
cc_189 N_C_M1003_g N_VGND_c_467_n 0.00157055f $X=2.255 $Y=0.495 $X2=0 $Y2=0
cc_190 N_C_M1005_g N_VGND_c_467_n 0.0106801f $X=2.615 $Y=0.495 $X2=0 $Y2=0
cc_191 N_C_M1003_g N_VGND_c_470_n 0.00338359f $X=2.255 $Y=0.495 $X2=0 $Y2=0
cc_192 N_C_M1005_g N_VGND_c_470_n 0.00445056f $X=2.615 $Y=0.495 $X2=0 $Y2=0
cc_193 N_C_M1003_g N_VGND_c_475_n 0.00481888f $X=2.255 $Y=0.495 $X2=0 $Y2=0
cc_194 N_C_M1005_g N_VGND_c_475_n 0.00796275f $X=2.615 $Y=0.495 $X2=0 $Y2=0
cc_195 N_B_c_274_n N_A_c_332_n 0.00965821f $X=3.49 $Y=0.78 $X2=-0.19 $Y2=-0.245
cc_196 N_B_M1004_g N_A_c_338_n 0.048393f $X=3.54 $Y=2.545 $X2=0 $Y2=0
cc_197 N_B_c_279_n N_A_c_338_n 0.0110482f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_198 N_B_c_275_n N_A_c_333_n 0.00965821f $X=3.49 $Y=0.855 $X2=0 $Y2=0
cc_199 N_B_c_277_n N_A_c_334_n 0.0119579f $X=3.58 $Y=1.72 $X2=0 $Y2=0
cc_200 N_B_c_282_n N_A_c_335_n 0.0119579f $X=3.58 $Y=1.885 $X2=0 $Y2=0
cc_201 N_B_c_279_n N_A_c_335_n 7.06261e-19 $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_202 N_B_c_276_n A 0.00417519f $X=3.58 $Y=1.215 $X2=0 $Y2=0
cc_203 N_B_c_278_n A 0.00374749f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_204 N_B_c_279_n A 0.0392993f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_205 N_B_c_276_n N_A_c_337_n 0.00591472f $X=3.58 $Y=1.215 $X2=0 $Y2=0
cc_206 N_B_c_278_n N_A_c_337_n 0.0119579f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_207 N_B_c_279_n N_A_c_337_n 6.93166e-19 $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_208 N_B_M1004_g N_VPWR_c_372_n 0.00212315f $X=3.54 $Y=2.545 $X2=0 $Y2=0
cc_209 N_B_c_279_n N_VPWR_c_372_n 0.0308427f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_210 N_B_M1004_g N_VPWR_c_373_n 0.00596257f $X=3.54 $Y=2.545 $X2=0 $Y2=0
cc_211 N_B_c_279_n N_VPWR_c_373_n 0.00914393f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_212 N_B_M1004_g N_VPWR_c_369_n 0.00771107f $X=3.54 $Y=2.545 $X2=0 $Y2=0
cc_213 N_B_c_279_n N_VPWR_c_369_n 0.0101955f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_214 N_B_c_272_n N_Y_c_404_n 0.0136522f $X=3.415 $Y=0.855 $X2=0 $Y2=0
cc_215 N_B_c_273_n N_Y_c_404_n 0.0102838f $X=3.205 $Y=0.855 $X2=0 $Y2=0
cc_216 N_B_c_275_n N_Y_c_404_n 0.00685914f $X=3.49 $Y=0.855 $X2=0 $Y2=0
cc_217 N_B_c_276_n N_Y_c_404_n 0.00695939f $X=3.58 $Y=1.215 $X2=0 $Y2=0
cc_218 N_B_c_278_n N_Y_c_404_n 0.00112623f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_219 N_B_c_279_n N_Y_c_404_n 0.0233855f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_220 N_B_c_274_n N_Y_c_405_n 0.00124703f $X=3.49 $Y=0.78 $X2=0 $Y2=0
cc_221 N_B_c_275_n N_Y_c_405_n 0.00430014f $X=3.49 $Y=0.855 $X2=0 $Y2=0
cc_222 N_B_c_271_n N_Y_c_406_n 0.0016682f $X=3.13 $Y=0.78 $X2=0 $Y2=0
cc_223 N_B_c_274_n N_Y_c_406_n 0.00897601f $X=3.49 $Y=0.78 $X2=0 $Y2=0
cc_224 N_B_c_278_n N_Y_c_406_n 2.12718e-19 $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_225 N_B_c_279_n N_Y_c_406_n 0.00132174f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_226 N_B_c_279_n A_733_409# 0.0116484f $X=3.58 $Y=1.38 $X2=-0.19 $Y2=-0.245
cc_227 N_B_c_271_n N_VGND_c_467_n 0.00844158f $X=3.13 $Y=0.78 $X2=0 $Y2=0
cc_228 N_B_c_271_n N_VGND_c_473_n 0.0053602f $X=3.13 $Y=0.78 $X2=0 $Y2=0
cc_229 N_B_c_272_n N_VGND_c_473_n 4.57848e-19 $X=3.415 $Y=0.855 $X2=0 $Y2=0
cc_230 N_B_c_274_n N_VGND_c_473_n 0.00502664f $X=3.49 $Y=0.78 $X2=0 $Y2=0
cc_231 N_B_c_271_n N_VGND_c_475_n 0.0103357f $X=3.13 $Y=0.78 $X2=0 $Y2=0
cc_232 N_B_c_272_n N_VGND_c_475_n 6.33118e-19 $X=3.415 $Y=0.855 $X2=0 $Y2=0
cc_233 N_B_c_274_n N_VGND_c_475_n 0.00942073f $X=3.49 $Y=0.78 $X2=0 $Y2=0
cc_234 N_A_c_338_n N_VPWR_c_372_n 0.0262314f $X=4.11 $Y=1.94 $X2=0 $Y2=0
cc_235 N_A_c_334_n N_VPWR_c_372_n 6.15125e-19 $X=4.17 $Y=1.575 $X2=0 $Y2=0
cc_236 A N_VPWR_c_372_n 0.0235749f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_237 N_A_c_338_n N_VPWR_c_373_n 0.00802402f $X=4.11 $Y=1.94 $X2=0 $Y2=0
cc_238 N_A_c_338_n N_VPWR_c_369_n 0.0144019f $X=4.11 $Y=1.94 $X2=0 $Y2=0
cc_239 N_A_c_333_n N_Y_c_404_n 0.00187706f $X=4.1 $Y=0.975 $X2=0 $Y2=0
cc_240 A N_Y_c_404_n 0.00878526f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_241 N_A_c_337_n N_Y_c_404_n 2.70936e-19 $X=4.19 $Y=1.07 $X2=0 $Y2=0
cc_242 N_A_c_332_n N_Y_c_405_n 0.00302883f $X=3.92 $Y=0.825 $X2=0 $Y2=0
cc_243 N_A_c_332_n N_Y_c_406_n 0.0106507f $X=3.92 $Y=0.825 $X2=0 $Y2=0
cc_244 N_A_c_332_n N_VGND_c_469_n 0.0161795f $X=3.92 $Y=0.825 $X2=0 $Y2=0
cc_245 A N_VGND_c_469_n 0.0291689f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_246 N_A_c_332_n N_VGND_c_473_n 0.00947719f $X=3.92 $Y=0.825 $X2=0 $Y2=0
cc_247 N_A_c_332_n N_VGND_c_475_n 0.0173835f $X=3.92 $Y=0.825 $X2=0 $Y2=0
cc_248 N_A_c_333_n N_VGND_c_475_n 7.74273e-19 $X=4.1 $Y=0.975 $X2=0 $Y2=0
cc_249 N_VPWR_c_370_n Y 0.0395659f $X=0.83 $Y=2.19 $X2=0 $Y2=0
cc_250 N_VPWR_c_373_n Y 0.0524562f $X=4.21 $Y=3.33 $X2=0 $Y2=0
cc_251 N_VPWR_c_369_n Y 0.0301033f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_252 N_Y_c_408_n N_VGND_c_466_n 0.00563913f $X=1.955 $Y=1.035 $X2=0 $Y2=0
cc_253 N_Y_c_404_n N_VGND_c_467_n 0.0234047f $X=3.54 $Y=0.95 $X2=0 $Y2=0
cc_254 N_Y_c_406_n N_VGND_c_467_n 0.0131248f $X=3.705 $Y=0.495 $X2=0 $Y2=0
cc_255 N_Y_c_408_n N_VGND_c_467_n 0.00684781f $X=1.955 $Y=1.035 $X2=0 $Y2=0
cc_256 N_Y_c_406_n N_VGND_c_469_n 0.0153904f $X=3.705 $Y=0.495 $X2=0 $Y2=0
cc_257 N_Y_c_408_n N_VGND_c_470_n 0.0372012f $X=1.955 $Y=1.035 $X2=0 $Y2=0
cc_258 N_Y_c_406_n N_VGND_c_473_n 0.0216454f $X=3.705 $Y=0.495 $X2=0 $Y2=0
cc_259 N_Y_c_406_n N_VGND_c_475_n 0.012407f $X=3.705 $Y=0.495 $X2=0 $Y2=0
cc_260 N_Y_c_408_n N_VGND_c_475_n 0.0272627f $X=1.955 $Y=1.035 $X2=0 $Y2=0
cc_261 N_Y_c_408_n A_302_57# 0.00179402f $X=1.955 $Y=1.035 $X2=-0.19 $Y2=-0.245
