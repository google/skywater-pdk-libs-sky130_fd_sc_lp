* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
X0 a_884_131# CIN a_978_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_978_419# B a_1050_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 COUT a_328_131# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR a_328_131# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 COUT a_328_131# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 SUM a_884_131# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR A a_604_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VGND B a_37_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR CIN a_604_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 COUT a_328_131# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR a_328_131# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_37_131# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_37_131# CIN a_328_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_440# CIN a_328_131# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VGND CIN a_604_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND A a_604_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_978_131# B a_1050_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR B a_27_440# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_604_419# a_328_131# a_884_131# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_414_131# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_884_131# SUM VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_884_131# CIN a_978_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 SUM a_884_131# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_328_131# B a_445_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 VGND a_328_131# COUT VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_604_419# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 a_27_440# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_1050_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 VPWR a_884_131# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 SUM a_884_131# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_328_131# B a_414_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_604_131# a_328_131# a_884_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VGND a_884_131# SUM VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 a_604_131# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1050_131# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 COUT a_328_131# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 SUM a_884_131# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 VGND a_328_131# COUT VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 VPWR a_884_131# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 a_445_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
