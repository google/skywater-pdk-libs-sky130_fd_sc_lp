* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_lp A0 A1 S VGND VNB VPB VPWR X
M1000 a_123_527# a_84_29# X VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1001 a_84_29# A1 a_281_527# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.008e+11p ps=1.32e+06u
M1002 VGND a_84_29# a_114_55# VNB nshort w=420000u l=150000u
+  ad=3.087e+11p pd=3.15e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_516_55# A1 a_84_29# VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=2.121e+11p ps=1.85e+06u
M1004 a_702_527# S VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=4.305e+11p ps=3.73e+06u
M1005 a_307_55# a_200_367# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1006 a_84_29# A0 a_307_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_200_367# S a_702_527# VPB phighvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1008 VGND S a_516_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_114_55# a_84_29# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1010 a_281_527# a_200_367# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_445_527# A0 a_84_29# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1012 VPWR S a_445_527# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_704_55# S VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1014 a_200_367# S a_704_55# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1015 VPWR a_84_29# a_123_527# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
