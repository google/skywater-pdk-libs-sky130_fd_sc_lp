* File: sky130_fd_sc_lp__a21o_lp.pex.spice
* Created: Wed Sep  2 09:20:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21O_LP%A2 3 7 9 10 14 15
r28 14 17 68.5216 $w=4.8e-07 $l=5.05e-07 $layer=POLY_cond $X=0.46 $Y=1.275
+ $X2=0.46 $Y2=1.78
r29 14 16 45.9721 $w=4.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.46 $Y=1.275
+ $X2=0.46 $Y2=1.11
r30 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.275 $X2=0.385 $Y2=1.275
r31 9 10 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r32 9 15 0.542326 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.275
r33 7 16 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.625 $Y=0.495
+ $X2=0.625 $Y2=1.11
r34 3 17 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.575 $Y=2.545
+ $X2=0.575 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_LP%A1 3 5 7 11 12 13 17 18
r39 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.105
+ $Y=1.29 $X2=1.105 $Y2=1.29
r40 12 13 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.127 $Y=1.295
+ $X2=1.127 $Y2=1.665
r41 12 18 0.153659 $w=3.73e-07 $l=5e-09 $layer=LI1_cond $X=1.127 $Y=1.295
+ $X2=1.127 $Y2=1.29
r42 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.105 $Y=1.63
+ $X2=1.105 $Y2=1.29
r43 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.125
+ $X2=1.105 $Y2=1.29
r44 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.795
+ $X2=1.105 $Y2=1.63
r45 5 7 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.105 $Y=1.795
+ $X2=1.105 $Y2=2.545
r46 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.015 $Y=0.495
+ $X2=1.015 $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_LP%B1 3 7 11 17 20 21 22 26
r51 21 22 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.675 $Y=1.29
+ $X2=1.675 $Y2=1.665
r52 21 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.675
+ $Y=1.29 $X2=1.675 $Y2=1.29
r53 19 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.675 $Y=1.63
+ $X2=1.675 $Y2=1.29
r54 19 20 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.63
+ $X2=1.675 $Y2=1.795
r55 16 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.675 $Y=1.275
+ $X2=1.675 $Y2=1.29
r56 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.675 $Y=1.2
+ $X2=1.945 $Y2=1.2
r57 13 16 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.585 $Y=1.2 $X2=1.675
+ $Y2=1.2
r58 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.945 $Y=1.125
+ $X2=1.945 $Y2=1.2
r59 9 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.945 $Y=1.125
+ $X2=1.945 $Y2=0.495
r60 7 20 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.635 $Y=2.545
+ $X2=1.635 $Y2=1.795
r61 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.585 $Y=1.125
+ $X2=1.585 $Y2=1.2
r62 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.585 $Y=1.125
+ $X2=1.585 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_LP%A_218_57# 1 2 7 9 10 12 13 15 19 21 22 25 30
+ 31 32
r72 35 37 16.8879 $w=6.08e-07 $l=5.05e-07 $layer=LI1_cond $X=2.325 $Y=0.98
+ $X2=2.325 $Y2=1.485
r73 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.465
+ $Y=0.98 $X2=2.465 $Y2=0.98
r74 32 35 2.35294 $w=6.08e-07 $l=1.2e-07 $layer=LI1_cond $X=2.325 $Y=0.86
+ $X2=2.325 $Y2=0.98
r75 31 37 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.105 $Y=2.025
+ $X2=2.105 $Y2=1.485
r76 30 31 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=1.962 $Y=2.19
+ $X2=1.962 $Y2=2.025
r77 23 30 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=1.962 $Y=2.252
+ $X2=1.962 $Y2=2.19
r78 23 25 17.0343 $w=4.53e-07 $l=6.48e-07 $layer=LI1_cond $X=1.962 $Y=2.252
+ $X2=1.962 $Y2=2.9
r79 21 32 8.42348 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=2.02 $Y=0.86
+ $X2=2.325 $Y2=0.86
r80 21 22 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.02 $Y=0.86
+ $X2=1.535 $Y2=0.86
r81 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.37 $Y=0.775
+ $X2=1.535 $Y2=0.86
r82 17 19 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.37 $Y=0.775
+ $X2=1.37 $Y2=0.495
r83 13 36 57.5495 $w=5.93e-07 $l=5.94559e-07 $layer=POLY_cond $X=2.815 $Y=1.485
+ $X2=2.62 $Y2=0.98
r84 13 15 247.211 $w=2.5e-07 $l=9.95e-07 $layer=POLY_cond $X=2.815 $Y=1.485
+ $X2=2.815 $Y2=2.48
r85 10 36 29.5333 $w=2.96e-07 $l=2.26164e-07 $layer=POLY_cond $X=2.765 $Y=0.815
+ $X2=2.62 $Y2=0.98
r86 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.765 $Y=0.815
+ $X2=2.765 $Y2=0.495
r87 7 36 29.5333 $w=2.96e-07 $l=3.16938e-07 $layer=POLY_cond $X=2.375 $Y=0.815
+ $X2=2.62 $Y2=0.98
r88 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.375 $Y=0.815
+ $X2=2.375 $Y2=0.495
r89 2 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.76
+ $Y=2.045 $X2=1.9 $Y2=2.19
r90 2 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.76
+ $Y=2.045 $X2=1.9 $Y2=2.9
r91 1 19 182 $w=1.7e-07 $l=3.70405e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.285 $X2=1.37 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_LP%A_33_409# 1 2 9 13 14 17
r30 17 19 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.37 $Y=2.19 $X2=1.37
+ $Y2=2.9
r31 15 17 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.37 $Y=2.145
+ $X2=1.37 $Y2=2.19
r32 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.205 $Y=2.06
+ $X2=1.37 $Y2=2.145
r33 13 14 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.205 $Y=2.06
+ $X2=0.475 $Y2=2.06
r34 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.31 $Y=2.19 $X2=0.31
+ $Y2=2.9
r35 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.31 $Y=2.145
+ $X2=0.475 $Y2=2.06
r36 7 9 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.31 $Y=2.145 $X2=0.31
+ $Y2=2.19
r37 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.23
+ $Y=2.045 $X2=1.37 $Y2=2.9
r38 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.23
+ $Y=2.045 $X2=1.37 $Y2=2.19
r39 1 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.045 $X2=0.31 $Y2=2.9
r40 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.045 $X2=0.31 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_LP%VPWR 1 2 11 15 20 21 22 32 33 36
r37 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 26 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r43 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.84 $Y2=3.33
r45 24 26 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 22 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 20 29 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.55 $Y2=3.33
r50 19 32 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.715 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=3.33
+ $X2=2.55 $Y2=3.33
r52 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.55 $Y=2.125
+ $X2=2.55 $Y2=2.835
r53 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=3.245
+ $X2=2.55 $Y2=3.33
r54 13 18 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.55 $Y=3.245
+ $X2=2.55 $Y2=2.835
r55 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=3.245 $X2=0.84
+ $Y2=3.33
r56 9 11 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.84 $Y=3.245
+ $X2=0.84 $Y2=2.49
r57 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=1.98 $X2=2.55 $Y2=2.835
r58 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=1.98 $X2=2.55 $Y2=2.125
r59 1 11 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=0.7
+ $Y=2.045 $X2=0.84 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_LP%X 1 2 9 13 14 15 16 23
r18 16 33 3.73456 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.03 $Y=1.665
+ $X2=3.03 $Y2=1.78
r19 16 21 2.6801 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=3.03 $Y=1.665 $X2=3.03
+ $Y2=1.565
r20 15 21 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.03 $Y=1.295
+ $X2=3.03 $Y2=1.565
r21 14 15 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.03 $Y=0.925
+ $X2=3.03 $Y2=1.295
r22 13 14 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.03 $Y=0.555
+ $X2=3.03 $Y2=0.925
r23 13 23 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=3.03 $Y=0.555 $X2=3.03
+ $Y2=0.495
r24 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.08 $Y=2.125 $X2=3.08
+ $Y2=2.835
r25 9 33 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.08 $Y=2.125
+ $X2=3.08 $Y2=1.78
r26 2 11 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.98 $X2=3.08 $Y2=2.835
r27 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.98 $X2=3.08 $Y2=2.125
r28 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.84
+ $Y=0.285 $X2=2.98 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_LP%VGND 1 2 7 9 13 15 17 27 28 34
r38 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r40 28 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r41 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.16
+ $Y2=0
r43 25 27 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=3.12
+ $Y2=0
r44 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r45 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r46 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 18 31 4.50939 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.287
+ $Y2=0
r48 18 20 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.72
+ $Y2=0
r49 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=2.16
+ $Y2=0
r50 17 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=1.68
+ $Y2=0
r51 15 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r52 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r53 15 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r54 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r55 11 13 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.43
r56 7 31 3.25678 $w=3.3e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.41 $Y=0.085
+ $X2=0.287 $Y2=0
r57 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.41 $Y=0.085 $X2=0.41
+ $Y2=0.495
r58 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.285 $X2=2.16 $Y2=0.43
r59 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.265
+ $Y=0.285 $X2=0.41 $Y2=0.495
.ends

