* File: sky130_fd_sc_lp__invkapwr_4.pex.spice
* Created: Fri Aug 28 10:39:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INVKAPWR_4%A 3 7 11 15 19 23 27 31 35 39 41 42 43 44
+ 45 69 70
r92 69 71 12.0818 $w=3.79e-07 $l=9.5e-08 $layer=POLY_cond $X=2.7 $Y=1.485
+ $X2=2.795 $Y2=1.485
r93 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7
+ $Y=1.46 $X2=2.7 $Y2=1.46
r94 67 69 42.6042 $w=3.79e-07 $l=3.35e-07 $layer=POLY_cond $X=2.365 $Y=1.485
+ $X2=2.7 $Y2=1.485
r95 65 67 0.635884 $w=3.79e-07 $l=5e-09 $layer=POLY_cond $X=2.36 $Y=1.485
+ $X2=2.365 $Y2=1.485
r96 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.36
+ $Y=1.46 $X2=2.36 $Y2=1.46
r97 63 65 54.0501 $w=3.79e-07 $l=4.25e-07 $layer=POLY_cond $X=1.935 $Y=1.485
+ $X2=2.36 $Y2=1.485
r98 61 63 32.4301 $w=3.79e-07 $l=2.55e-07 $layer=POLY_cond $X=1.68 $Y=1.485
+ $X2=1.935 $Y2=1.485
r99 59 61 22.2559 $w=3.79e-07 $l=1.75e-07 $layer=POLY_cond $X=1.505 $Y=1.485
+ $X2=1.68 $Y2=1.485
r100 57 59 20.9842 $w=3.79e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.485
+ $X2=1.505 $Y2=1.485
r101 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.34
+ $Y=1.46 $X2=1.34 $Y2=1.46
r102 55 57 33.7018 $w=3.79e-07 $l=2.65e-07 $layer=POLY_cond $X=1.075 $Y=1.485
+ $X2=1.34 $Y2=1.485
r103 53 55 9.53826 $w=3.79e-07 $l=7.5e-08 $layer=POLY_cond $X=1 $Y=1.485
+ $X2=1.075 $Y2=1.485
r104 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.46
+ $X2=1 $Y2=1.46
r105 51 53 45.1478 $w=3.79e-07 $l=3.55e-07 $layer=POLY_cond $X=0.645 $Y=1.485
+ $X2=1 $Y2=1.485
r106 45 70 2.06408 $w=3.33e-07 $l=6e-08 $layer=LI1_cond $X=2.64 $Y=1.377 $X2=2.7
+ $Y2=1.377
r107 45 66 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=2.64 $Y=1.377
+ $X2=2.36 $Y2=1.377
r108 44 66 6.88026 $w=3.33e-07 $l=2e-07 $layer=LI1_cond $X=2.16 $Y=1.377
+ $X2=2.36 $Y2=1.377
r109 43 44 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.377
+ $X2=2.16 $Y2=1.377
r110 43 58 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=1.68 $Y=1.377
+ $X2=1.34 $Y2=1.377
r111 43 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.46 $X2=1.68 $Y2=1.46
r112 42 58 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.377
+ $X2=1.34 $Y2=1.377
r113 42 54 6.88026 $w=3.33e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=1.377 $X2=1
+ $Y2=1.377
r114 41 54 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=0.72 $Y=1.377 $X2=1
+ $Y2=1.377
r115 37 71 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.795 $Y=1.675
+ $X2=2.795 $Y2=1.485
r116 37 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.795 $Y=1.675
+ $X2=2.795 $Y2=2.465
r117 33 67 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.365 $Y=1.675
+ $X2=2.365 $Y2=1.485
r118 33 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.365 $Y=1.675
+ $X2=2.365 $Y2=2.465
r119 29 67 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.365 $Y=1.295
+ $X2=2.365 $Y2=1.485
r120 29 31 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=2.365 $Y=1.295
+ $X2=2.365 $Y2=0.56
r121 25 63 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.935 $Y=1.675
+ $X2=1.935 $Y2=1.485
r122 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.935 $Y=1.675
+ $X2=1.935 $Y2=2.465
r123 21 63 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.935 $Y=1.295
+ $X2=1.935 $Y2=1.485
r124 21 23 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.935 $Y=1.295
+ $X2=1.935 $Y2=0.56
r125 17 59 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.505 $Y=1.675
+ $X2=1.505 $Y2=1.485
r126 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.505 $Y=1.675
+ $X2=1.505 $Y2=2.465
r127 13 59 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.505 $Y=1.295
+ $X2=1.505 $Y2=1.485
r128 13 15 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.505 $Y=1.295
+ $X2=1.505 $Y2=0.56
r129 9 55 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.075 $Y=1.675
+ $X2=1.075 $Y2=1.485
r130 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.075 $Y=1.675
+ $X2=1.075 $Y2=2.465
r131 5 55 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.075 $Y=1.295
+ $X2=1.075 $Y2=1.485
r132 5 7 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.075 $Y=1.295
+ $X2=1.075 $Y2=0.56
r133 1 51 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.645 $Y=1.675
+ $X2=0.645 $Y2=1.485
r134 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.645 $Y=1.675
+ $X2=0.645 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_4%KAPWR 1 2 3 4 13 16 24 32 40 44 52
r45 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=2.81
+ $X2=3.015 $Y2=2.81
r46 40 43 26.6644 $w=2.53e-07 $l=5.9e-07 $layer=LI1_cond $X=3.007 $Y=2.22
+ $X2=3.007 $Y2=2.81
r47 36 44 0.503471 $w=2.55e-07 $l=8.7e-07 $layer=MET1_cond $X=2.145 $Y=2.817
+ $X2=3.015 $Y2=2.817
r48 36 52 0.266203 $w=2.55e-07 $l=4.6e-07 $layer=MET1_cond $X=2.145 $Y=2.817
+ $X2=1.685 $Y2=2.817
r49 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.145 $Y=2.81
+ $X2=2.145 $Y2=2.81
r50 32 35 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=2.15 $Y=2.22
+ $X2=2.15 $Y2=2.81
r51 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.295 $Y=2.81
+ $X2=1.295 $Y2=2.81
r52 24 27 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=1.29 $Y=2.22
+ $X2=1.29 $Y2=2.81
r53 20 28 0.500577 $w=2.55e-07 $l=8.65e-07 $layer=MET1_cond $X=0.43 $Y=2.817
+ $X2=1.295 $Y2=2.817
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.43 $Y=2.81
+ $X2=0.43 $Y2=2.81
r55 16 19 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=0.43 $Y=2.22
+ $X2=0.43 $Y2=2.81
r56 13 52 0.00289351 $w=2.55e-07 $l=5e-09 $layer=MET1_cond $X=1.68 $Y=2.817
+ $X2=1.685 $Y2=2.817
r57 13 28 0.2228 $w=2.55e-07 $l=3.85e-07 $layer=MET1_cond $X=1.68 $Y=2.817
+ $X2=1.295 $Y2=2.817
r58 4 43 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.835 $X2=3.01 $Y2=2.91
r59 4 40 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.835 $X2=3.01 $Y2=2.22
r60 3 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.15 $Y2=2.91
r61 3 32 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.15 $Y2=2.22
r62 2 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=1.835 $X2=1.29 $Y2=2.91
r63 2 24 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=1.835 $X2=1.29 $Y2=2.22
r64 1 19 400 $w=1.7e-07 $l=1.13815e-06 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.835 $X2=0.43 $Y2=2.91
r65 1 16 400 $w=1.7e-07 $l=4.45281e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.835 $X2=0.43 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_4%Y 1 2 3 4 5 17 18 19 20 21 24 28 32 34 38
+ 42 46 50 54 55 56 58 60 61 62 63 70 71 76
r116 71 76 2.99754 $w=1.83e-07 $l=5e-08 $layer=LI1_cond $X=3.127 $Y=1.715
+ $X2=3.127 $Y2=1.665
r117 63 71 3.28106 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.127 $Y=1.8
+ $X2=3.127 $Y2=1.715
r118 63 76 1.07912 $w=1.83e-07 $l=1.8e-08 $layer=LI1_cond $X=3.127 $Y=1.647
+ $X2=3.127 $Y2=1.665
r119 62 63 21.1027 $w=1.83e-07 $l=3.52e-07 $layer=LI1_cond $X=3.127 $Y=1.295
+ $X2=3.127 $Y2=1.647
r120 62 70 15.2875 $w=1.83e-07 $l=2.55e-07 $layer=LI1_cond $X=3.127 $Y=1.295
+ $X2=3.127 $Y2=1.04
r121 61 70 3.55727 $w=1.85e-07 $l=1e-07 $layer=LI1_cond $X=3.127 $Y=0.94
+ $X2=3.127 $Y2=1.04
r122 59 63 17.9392 $w=2.03e-07 $l=3.25e-07 $layer=LI1_cond $X=2.71 $Y=1.8
+ $X2=3.035 $Y2=1.8
r123 59 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=1.8 $X2=2.58
+ $Y2=1.8
r124 57 61 24.9971 $w=3.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.275 $Y=0.94
+ $X2=3.035 $Y2=0.94
r125 57 58 6.29182 $w=2e-07 $l=1.28e-07 $layer=LI1_cond $X=2.275 $Y=0.94
+ $X2=2.147 $Y2=0.94
r126 50 52 39.0058 $w=2.58e-07 $l=8.8e-07 $layer=LI1_cond $X=2.58 $Y=2 $X2=2.58
+ $Y2=2.88
r127 48 60 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=1.885
+ $X2=2.58 $Y2=1.8
r128 48 50 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=2.58 $Y=1.885
+ $X2=2.58 $Y2=2
r129 44 58 0.484182 $w=2.55e-07 $l=1e-07 $layer=LI1_cond $X=2.147 $Y=0.84
+ $X2=2.147 $Y2=0.94
r130 44 46 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=2.147 $Y=0.84
+ $X2=2.147 $Y2=0.56
r131 43 56 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.85 $Y=1.8
+ $X2=1.722 $Y2=1.8
r132 42 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.45 $Y=1.8 $X2=2.58
+ $Y2=1.8
r133 42 43 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.45 $Y=1.8 $X2=1.85
+ $Y2=1.8
r134 38 40 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=1.722 $Y=2
+ $X2=1.722 $Y2=2.88
r135 36 56 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.722 $Y=1.885
+ $X2=1.722 $Y2=1.8
r136 36 38 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=1.722 $Y=1.885
+ $X2=1.722 $Y2=2
r137 35 55 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.42 $Y=0.94 $X2=1.29
+ $Y2=0.94
r138 34 58 6.29182 $w=2e-07 $l=1.27e-07 $layer=LI1_cond $X=2.02 $Y=0.94
+ $X2=2.147 $Y2=0.94
r139 34 35 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=2.02 $Y=0.94 $X2=1.42
+ $Y2=0.94
r140 30 55 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=1.29 $Y=0.84 $X2=1.29
+ $Y2=0.94
r141 30 32 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=1.29 $Y=0.84
+ $X2=1.29 $Y2=0.56
r142 29 54 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.99 $Y=1.8
+ $X2=0.862 $Y2=1.8
r143 28 56 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.595 $Y=1.8
+ $X2=1.722 $Y2=1.8
r144 28 29 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.595 $Y=1.8
+ $X2=0.99 $Y2=1.8
r145 24 26 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=0.862 $Y=2
+ $X2=0.862 $Y2=2.88
r146 22 54 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.862 $Y=1.885
+ $X2=0.862 $Y2=1.8
r147 22 24 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=0.862 $Y=1.885
+ $X2=0.862 $Y2=2
r148 20 54 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.735 $Y=1.8
+ $X2=0.862 $Y2=1.8
r149 20 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.735 $Y=1.8
+ $X2=0.4 $Y2=1.8
r150 18 55 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.16 $Y=0.94 $X2=1.29
+ $Y2=0.94
r151 18 19 42.1455 $w=1.98e-07 $l=7.6e-07 $layer=LI1_cond $X=1.16 $Y=0.94
+ $X2=0.4 $Y2=0.94
r152 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.315 $Y=1.715
+ $X2=0.4 $Y2=1.8
r153 16 19 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.315 $Y=1.04
+ $X2=0.4 $Y2=0.94
r154 16 17 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.315 $Y=1.04
+ $X2=0.315 $Y2=1.715
r155 5 52 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.835 $X2=2.58 $Y2=2.88
r156 5 50 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.835 $X2=2.58 $Y2=2
r157 4 40 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.835 $X2=1.72 $Y2=2.88
r158 4 38 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.835 $X2=1.72 $Y2=2
r159 3 26 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.835 $X2=0.86 $Y2=2.88
r160 3 24 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.835 $X2=0.86 $Y2=2
r161 2 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.01
+ $Y=0.35 $X2=2.15 $Y2=0.56
r162 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.15
+ $Y=0.35 $X2=1.29 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_4%VGND 1 2 3 14 18 22 24 26 31 38 39 42 45
+ 48
r34 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 39 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r37 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r38 36 48 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.595
+ $Y2=0
r39 36 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=3.12
+ $Y2=0
r40 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 32 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.72
+ $Y2=0
r43 32 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.16
+ $Y2=0
r44 31 48 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.595
+ $Y2=0
r45 31 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.16
+ $Y2=0
r46 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r47 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r48 27 42 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.842
+ $Y2=0
r49 27 29 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r50 26 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.59 $Y=0 $X2=1.72
+ $Y2=0
r51 26 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.59 $Y=0 $X2=1.2
+ $Y2=0
r52 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r53 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 24 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 20 48 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0
r56 20 22 16.1342 $w=2.98e-07 $l=4.2e-07 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0.505
r57 16 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0
r58 16 18 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0.505
r59 12 42 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0
r60 12 14 16.4077 $w=2.93e-07 $l=4.2e-07 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0.505
r61 3 22 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.35 $X2=2.58 $Y2=0.505
r62 2 18 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.58
+ $Y=0.35 $X2=1.72 $Y2=0.505
r63 1 14 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.735
+ $Y=0.35 $X2=0.86 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_4%VPWR 1 8 14
r38 5 14 0.00453869 $w=3.36e-06 $l=1.22e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.208
r39 5 8 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 4 8 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=3.12
+ $Y2=3.33
r41 4 5 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 1 14 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=3.207
+ $X2=1.68 $Y2=3.208
.ends

