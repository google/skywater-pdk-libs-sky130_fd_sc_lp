* File: sky130_fd_sc_lp__einvp_m.pxi.spice
* Created: Wed Sep  2 09:52:56 2020
* 
x_PM_SKY130_FD_SC_LP__EINVP_M%TE N_TE_c_40_n N_TE_M1001_g N_TE_c_48_n
+ N_TE_M1005_g N_TE_c_42_n N_TE_c_43_n N_TE_M1004_g N_TE_c_44_n N_TE_c_49_n TE
+ TE N_TE_c_46_n PM_SKY130_FD_SC_LP__EINVP_M%TE
x_PM_SKY130_FD_SC_LP__EINVP_M%A_42_129# N_A_42_129#_M1001_s N_A_42_129#_M1005_s
+ N_A_42_129#_M1000_g N_A_42_129#_c_99_n N_A_42_129#_c_93_n N_A_42_129#_c_100_n
+ N_A_42_129#_c_94_n N_A_42_129#_c_95_n N_A_42_129#_c_96_n N_A_42_129#_c_97_n
+ PM_SKY130_FD_SC_LP__EINVP_M%A_42_129#
x_PM_SKY130_FD_SC_LP__EINVP_M%A N_A_M1003_g N_A_M1002_g A N_A_c_140_n
+ N_A_c_141_n PM_SKY130_FD_SC_LP__EINVP_M%A
x_PM_SKY130_FD_SC_LP__EINVP_M%VPWR N_VPWR_M1005_d N_VPWR_c_164_n N_VPWR_c_165_n
+ N_VPWR_c_166_n VPWR N_VPWR_c_167_n N_VPWR_c_163_n
+ PM_SKY130_FD_SC_LP__EINVP_M%VPWR
x_PM_SKY130_FD_SC_LP__EINVP_M%Z N_Z_M1003_d N_Z_M1002_d Z Z Z Z Z Z
+ PM_SKY130_FD_SC_LP__EINVP_M%Z
x_PM_SKY130_FD_SC_LP__EINVP_M%VGND N_VGND_M1001_d N_VGND_c_207_n N_VGND_c_202_n
+ N_VGND_c_203_n N_VGND_c_204_n VGND N_VGND_c_205_n N_VGND_c_206_n
+ PM_SKY130_FD_SC_LP__EINVP_M%VGND
cc_1 VNB N_TE_c_40_n 0.0258556f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=2.415
cc_2 VNB N_TE_M1001_g 0.0138411f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.855
cc_3 VNB N_TE_c_42_n 0.0178492f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.46
cc_4 VNB N_TE_c_43_n 0.0161561f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=0.535
cc_5 VNB N_TE_c_44_n 0.0177263f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.25
cc_6 VNB TE 0.0265935f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_7 VNB N_TE_c_46_n 0.0399868f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.37
cc_8 VNB N_A_42_129#_c_93_n 0.0273234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_42_129#_c_94_n 0.00416241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_42_129#_c_95_n 0.00504264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_42_129#_c_96_n 0.00232623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_42_129#_c_97_n 0.0164931f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.37
cc_13 VNB N_A_M1003_g 0.0506113f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.535
cc_14 VNB N_A_c_140_n 0.0440338f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.46
cc_15 VNB N_A_c_141_n 0.0200747f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.46
cc_16 VNB N_VPWR_c_163_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=2.49
cc_17 VNB Z 0.0348805f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.565
cc_18 VNB N_VGND_c_202_n 0.00835621f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.885
cc_19 VNB N_VGND_c_203_n 0.0277324f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.46
cc_20 VNB N_VGND_c_204_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=0.535
cc_21 VNB N_VGND_c_205_n 0.0226012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_206_n 0.14388f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.49
cc_23 VPB N_TE_c_40_n 0.0483378f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=2.415
cc_24 VPB N_TE_c_48_n 0.019498f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.565
cc_25 VPB N_TE_c_49_n 0.0266064f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.49
cc_26 VPB N_A_42_129#_M1000_g 0.035645f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.885
cc_27 VPB N_A_42_129#_c_99_n 0.0190735f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=0.855
cc_28 VPB N_A_42_129#_c_100_n 0.0524634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_A_42_129#_c_94_n 0.00824485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_A_42_129#_c_95_n 0.0021011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_A_42_129#_c_96_n 0.00295858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_42_129#_c_97_n 0.0279257f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.37
cc_33 VPB N_A_M1003_g 0.0755289f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.535
cc_34 VPB N_VPWR_c_164_n 0.00494119f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.855
cc_35 VPB N_VPWR_c_165_n 0.0229334f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.885
cc_36 VPB N_VPWR_c_166_n 0.00401177f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=0.46
cc_37 VPB N_VPWR_c_167_n 0.0307105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_163_n 0.0493669f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=2.49
cc_39 VPB Z 0.0527368f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.565
cc_40 N_TE_c_40_n N_A_42_129#_M1000_g 0.00570558f $X=0.46 $Y=2.415 $X2=0 $Y2=0
cc_41 N_TE_c_49_n N_A_42_129#_M1000_g 0.0226793f $X=0.63 $Y=2.49 $X2=0 $Y2=0
cc_42 N_TE_c_40_n N_A_42_129#_c_93_n 0.0144185f $X=0.46 $Y=2.415 $X2=0 $Y2=0
cc_43 N_TE_M1001_g N_A_42_129#_c_93_n 0.00737703f $X=0.55 $Y=0.855 $X2=0 $Y2=0
cc_44 N_TE_c_43_n N_A_42_129#_c_93_n 6.9098e-19 $X=1.06 $Y=0.535 $X2=0 $Y2=0
cc_45 N_TE_c_44_n N_A_42_129#_c_93_n 0.0119707f $X=0.55 $Y=1.25 $X2=0 $Y2=0
cc_46 TE N_A_42_129#_c_93_n 0.0226266f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_47 N_TE_c_40_n N_A_42_129#_c_100_n 0.0297507f $X=0.46 $Y=2.415 $X2=0 $Y2=0
cc_48 N_TE_c_48_n N_A_42_129#_c_100_n 0.00472061f $X=0.63 $Y=2.565 $X2=0 $Y2=0
cc_49 N_TE_c_49_n N_A_42_129#_c_100_n 0.0102133f $X=0.63 $Y=2.49 $X2=0 $Y2=0
cc_50 N_TE_c_40_n N_A_42_129#_c_94_n 0.00317005f $X=0.46 $Y=2.415 $X2=0 $Y2=0
cc_51 N_TE_c_44_n N_A_42_129#_c_94_n 0.00357807f $X=0.55 $Y=1.25 $X2=0 $Y2=0
cc_52 N_TE_c_40_n N_A_42_129#_c_95_n 0.00637328f $X=0.46 $Y=2.415 $X2=0 $Y2=0
cc_53 N_TE_c_40_n N_A_42_129#_c_96_n 0.00143165f $X=0.46 $Y=2.415 $X2=0 $Y2=0
cc_54 N_TE_c_43_n N_A_42_129#_c_96_n 2.00878e-19 $X=1.06 $Y=0.535 $X2=0 $Y2=0
cc_55 N_TE_c_40_n N_A_42_129#_c_97_n 0.0342622f $X=0.46 $Y=2.415 $X2=0 $Y2=0
cc_56 N_TE_c_43_n N_A_42_129#_c_97_n 0.00529345f $X=1.06 $Y=0.535 $X2=0 $Y2=0
cc_57 N_TE_c_43_n N_A_M1003_g 0.0247998f $X=1.06 $Y=0.535 $X2=0 $Y2=0
cc_58 N_TE_c_44_n N_A_M1003_g 0.00284316f $X=0.55 $Y=1.25 $X2=0 $Y2=0
cc_59 N_TE_c_42_n N_A_c_140_n 0.0247998f $X=0.985 $Y=0.46 $X2=0 $Y2=0
cc_60 N_TE_c_46_n N_A_c_140_n 0.00320788f $X=0.805 $Y=0.37 $X2=0 $Y2=0
cc_61 N_TE_c_42_n N_A_c_141_n 8.4183e-19 $X=0.985 $Y=0.46 $X2=0 $Y2=0
cc_62 N_TE_c_48_n N_VPWR_c_164_n 0.00288714f $X=0.63 $Y=2.565 $X2=0 $Y2=0
cc_63 N_TE_c_48_n N_VPWR_c_165_n 0.00585385f $X=0.63 $Y=2.565 $X2=0 $Y2=0
cc_64 N_TE_c_49_n N_VPWR_c_165_n 9.47564e-19 $X=0.63 $Y=2.49 $X2=0 $Y2=0
cc_65 N_TE_c_48_n N_VPWR_c_163_n 0.0118545f $X=0.63 $Y=2.565 $X2=0 $Y2=0
cc_66 N_TE_c_49_n N_VPWR_c_163_n 8.53344e-19 $X=0.63 $Y=2.49 $X2=0 $Y2=0
cc_67 N_TE_c_43_n Z 0.00104353f $X=1.06 $Y=0.535 $X2=0 $Y2=0
cc_68 N_TE_c_42_n N_VGND_c_207_n 0.00277855f $X=0.985 $Y=0.46 $X2=0 $Y2=0
cc_69 N_TE_c_43_n N_VGND_c_207_n 0.00685999f $X=1.06 $Y=0.535 $X2=0 $Y2=0
cc_70 TE N_VGND_c_207_n 0.00919486f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_71 N_TE_c_46_n N_VGND_c_207_n 4.91325e-19 $X=0.805 $Y=0.37 $X2=0 $Y2=0
cc_72 N_TE_M1001_g N_VGND_c_202_n 9.0767e-19 $X=0.55 $Y=0.855 $X2=0 $Y2=0
cc_73 N_TE_c_42_n N_VGND_c_202_n 0.00779128f $X=0.985 $Y=0.46 $X2=0 $Y2=0
cc_74 N_TE_c_43_n N_VGND_c_202_n 0.00618273f $X=1.06 $Y=0.535 $X2=0 $Y2=0
cc_75 TE N_VGND_c_202_n 0.0263926f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_76 N_TE_c_46_n N_VGND_c_202_n 0.00210454f $X=0.805 $Y=0.37 $X2=0 $Y2=0
cc_77 N_TE_c_42_n N_VGND_c_203_n 0.00512312f $X=0.985 $Y=0.46 $X2=0 $Y2=0
cc_78 TE N_VGND_c_203_n 0.036111f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_79 N_TE_c_46_n N_VGND_c_203_n 0.00649036f $X=0.805 $Y=0.37 $X2=0 $Y2=0
cc_80 N_TE_c_42_n N_VGND_c_206_n 0.00540455f $X=0.985 $Y=0.46 $X2=0 $Y2=0
cc_81 TE N_VGND_c_206_n 0.0229022f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_82 N_TE_c_46_n N_VGND_c_206_n 0.00896615f $X=0.805 $Y=0.37 $X2=0 $Y2=0
cc_83 N_A_42_129#_c_99_n N_A_M1003_g 0.0721907f $X=0.955 $Y=2.205 $X2=0 $Y2=0
cc_84 N_A_42_129#_c_96_n N_A_M1003_g 0.00200334f $X=0.94 $Y=1.7 $X2=0 $Y2=0
cc_85 N_A_42_129#_c_97_n N_A_M1003_g 0.0265267f $X=0.94 $Y=1.7 $X2=0 $Y2=0
cc_86 N_A_42_129#_M1000_g N_VPWR_c_164_n 0.00288714f $X=1.06 $Y=2.885 $X2=0
+ $Y2=0
cc_87 N_A_42_129#_c_99_n N_VPWR_c_164_n 0.00298806f $X=0.955 $Y=2.205 $X2=0
+ $Y2=0
cc_88 N_A_42_129#_c_96_n N_VPWR_c_164_n 0.00269513f $X=0.94 $Y=1.7 $X2=0 $Y2=0
cc_89 N_A_42_129#_c_100_n N_VPWR_c_165_n 0.0151286f $X=0.415 $Y=2.82 $X2=0 $Y2=0
cc_90 N_A_42_129#_M1000_g N_VPWR_c_167_n 0.00585385f $X=1.06 $Y=2.885 $X2=0
+ $Y2=0
cc_91 N_A_42_129#_M1005_s N_VPWR_c_163_n 0.00265135f $X=0.29 $Y=2.675 $X2=0
+ $Y2=0
cc_92 N_A_42_129#_M1000_g N_VPWR_c_163_n 0.0105559f $X=1.06 $Y=2.885 $X2=0 $Y2=0
cc_93 N_A_42_129#_c_100_n N_VPWR_c_163_n 0.0128913f $X=0.415 $Y=2.82 $X2=0 $Y2=0
cc_94 N_A_42_129#_c_99_n Z 0.0037681f $X=0.955 $Y=2.205 $X2=0 $Y2=0
cc_95 N_A_42_129#_c_96_n Z 0.0225526f $X=0.94 $Y=1.7 $X2=0 $Y2=0
cc_96 N_A_42_129#_c_97_n Z 0.00164221f $X=0.94 $Y=1.7 $X2=0 $Y2=0
cc_97 N_A_42_129#_c_94_n N_VGND_c_207_n 0.00567928f $X=0.855 $Y=1.62 $X2=0 $Y2=0
cc_98 N_A_42_129#_c_96_n N_VGND_c_207_n 0.00482889f $X=0.94 $Y=1.7 $X2=0 $Y2=0
cc_99 N_A_42_129#_c_97_n N_VGND_c_207_n 0.00260049f $X=0.94 $Y=1.7 $X2=0 $Y2=0
cc_100 N_A_M1003_g N_VPWR_c_167_n 0.00553654f $X=1.42 $Y=0.855 $X2=0 $Y2=0
cc_101 N_A_M1003_g N_VPWR_c_163_n 0.0109726f $X=1.42 $Y=0.855 $X2=0 $Y2=0
cc_102 N_A_M1003_g Z 0.0765969f $X=1.42 $Y=0.855 $X2=0 $Y2=0
cc_103 N_A_c_140_n Z 9.48991e-19 $X=1.51 $Y=0.37 $X2=0 $Y2=0
cc_104 N_A_c_141_n Z 0.0213231f $X=1.51 $Y=0.37 $X2=0 $Y2=0
cc_105 N_A_M1003_g N_VGND_c_202_n 5.13034e-19 $X=1.42 $Y=0.855 $X2=0 $Y2=0
cc_106 N_A_c_140_n N_VGND_c_202_n 0.0027488f $X=1.51 $Y=0.37 $X2=0 $Y2=0
cc_107 N_A_c_141_n N_VGND_c_202_n 0.0287939f $X=1.51 $Y=0.37 $X2=0 $Y2=0
cc_108 N_A_c_140_n N_VGND_c_205_n 0.00634027f $X=1.51 $Y=0.37 $X2=0 $Y2=0
cc_109 N_A_c_141_n N_VGND_c_205_n 0.0241449f $X=1.51 $Y=0.37 $X2=0 $Y2=0
cc_110 N_A_c_140_n N_VGND_c_206_n 0.00878401f $X=1.51 $Y=0.37 $X2=0 $Y2=0
cc_111 N_A_c_141_n N_VGND_c_206_n 0.0149444f $X=1.51 $Y=0.37 $X2=0 $Y2=0
cc_112 N_VPWR_c_163_n A_227_535# 0.00899413f $X=1.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_113 N_VPWR_c_163_n N_Z_M1002_d 0.00235821f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_114 N_VPWR_c_167_n Z 0.010662f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_115 N_VPWR_c_163_n Z 0.0115728f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_116 Z N_VGND_c_206_n 0.00197725f $X=1.595 $Y=0.84 $X2=0 $Y2=0
