# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a221o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a221o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 1.185000 3.955000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.190000 1.185000 3.205000 1.515000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.295000 1.195000 6.135000 1.525000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.630000 1.405000 7.525000 1.620000 ;
        RECT 6.640000 1.620000 7.525000 1.750000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.465000 1.195000 5.125000 1.525000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.060000 1.660000 1.230000 ;
        RECT 0.110000 1.230000 0.335000 1.755000 ;
        RECT 0.110000 1.755000 1.660000 1.925000 ;
        RECT 0.610000 0.255000 0.800000 1.045000 ;
        RECT 0.610000 1.045000 1.660000 1.060000 ;
        RECT 0.610000 1.925000 0.790000 3.075000 ;
        RECT 1.470000 0.255000 1.660000 1.045000 ;
        RECT 1.470000 1.925000 1.660000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.110000  0.085000 0.440000 0.890000 ;
      RECT 0.110000  2.095000 0.440000 3.245000 ;
      RECT 0.505000  1.400000 2.020000 1.585000 ;
      RECT 0.970000  0.085000 1.300000 0.875000 ;
      RECT 0.970000  2.095000 1.300000 3.245000 ;
      RECT 1.830000  0.085000 2.160000 1.015000 ;
      RECT 1.830000  2.045000 2.160000 3.245000 ;
      RECT 1.850000  1.585000 2.020000 1.690000 ;
      RECT 1.850000  1.690000 4.295000 1.705000 ;
      RECT 1.850000  1.705000 4.830000 1.875000 ;
      RECT 2.330000  0.255000 2.520000 0.845000 ;
      RECT 2.330000  0.845000 3.955000 1.015000 ;
      RECT 2.330000  2.045000 4.315000 2.215000 ;
      RECT 2.330000  2.215000 3.380000 2.225000 ;
      RECT 2.330000  2.225000 2.520000 3.075000 ;
      RECT 2.690000  0.085000 3.020000 0.675000 ;
      RECT 2.690000  2.395000 3.020000 3.245000 ;
      RECT 3.190000  2.225000 3.380000 3.065000 ;
      RECT 3.210000  0.255000 4.365000 0.425000 ;
      RECT 3.210000  0.425000 3.530000 0.675000 ;
      RECT 3.550000  2.385000 3.880000 3.245000 ;
      RECT 3.700000  0.595000 3.955000 0.845000 ;
      RECT 4.070000  2.215000 4.315000 2.445000 ;
      RECT 4.070000  2.445000 5.620000 2.615000 ;
      RECT 4.070000  2.785000 6.120000 2.895000 ;
      RECT 4.070000  2.895000 6.980000 3.065000 ;
      RECT 4.125000  0.425000 4.365000 0.855000 ;
      RECT 4.125000  0.855000 5.235000 1.025000 ;
      RECT 4.125000  1.025000 4.295000 1.690000 ;
      RECT 4.500000  1.875000 4.830000 2.275000 ;
      RECT 4.535000  0.085000 4.795000 0.685000 ;
      RECT 4.965000  0.255000 6.120000 0.515000 ;
      RECT 4.965000  0.515000 5.235000 0.855000 ;
      RECT 5.360000  1.705000 6.470000 1.875000 ;
      RECT 5.360000  1.875000 5.620000 2.445000 ;
      RECT 5.405000  0.685000 6.570000 1.015000 ;
      RECT 5.790000  2.055000 6.120000 2.785000 ;
      RECT 6.290000  1.875000 6.470000 2.725000 ;
      RECT 6.310000  0.255000 6.570000 0.685000 ;
      RECT 6.370000  1.015000 6.570000 1.065000 ;
      RECT 6.370000  1.065000 7.500000 1.235000 ;
      RECT 6.650000  1.920000 6.980000 2.895000 ;
      RECT 6.740000  0.085000 7.070000 0.895000 ;
      RECT 7.240000  0.255000 7.500000 1.065000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__a221o_4
END LIBRARY
