* File: sky130_fd_sc_lp__dfrtn_1.pex.spice
* Created: Wed Sep  2 09:43:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFRTN_1%D 3 6 8 9 10 15 17
c44 10 0 1.04924e-19 $X=1.2 $Y=1.295
r45 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.3
+ $X2=1.085 $Y2=1.465
r46 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.3
+ $X2=1.085 $Y2=1.135
r47 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.3 $X2=1.085 $Y2=1.3
r48 10 16 5.40943 $w=2.43e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.272
+ $X2=1.085 $Y2=1.272
r49 9 16 17.169 $w=2.43e-07 $l=3.65e-07 $layer=LI1_cond $X=0.72 $Y=1.272
+ $X2=1.085 $Y2=1.272
r50 8 9 22.5785 $w=2.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.272 $X2=0.72
+ $Y2=1.272
r51 6 18 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=1.135 $Y=2.525
+ $X2=1.135 $Y2=1.465
r52 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.995 $Y=0.815
+ $X2=0.995 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%A_294_35# 1 2 9 12 16 20 21 24 27 31 32 33
+ 35 37 39 40 42 43 44 46 49 50 52 56 57 59 62 71
c196 62 0 7.41338e-20 $X=1.635 $Y=0.505
c197 59 0 1.17612e-20 $X=5.745 $Y=0.345
c198 44 0 4.89731e-20 $X=5.14 $Y=0.34
c199 40 0 1.44421e-19 $X=4.245 $Y=0.675
c200 16 0 1.88823e-19 $X=5.42 $Y=2.655
c201 12 0 1.75901e-19 $X=2.16 $Y=2.525
r202 57 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.47 $Y=1.645
+ $X2=5.47 $Y2=1.81
r203 56 58 11.8551 $w=2.83e-07 $l=2.75e-07 $layer=LI1_cond $X=5.47 $Y=1.645
+ $X2=5.745 $Y2=1.645
r204 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.47
+ $Y=1.645 $X2=5.47 $Y2=1.645
r205 50 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.21 $Y=0.35
+ $X2=6.21 $Y2=0.515
r206 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.21
+ $Y=0.35 $X2=6.21 $Y2=0.35
r207 47 59 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=0.345
+ $X2=5.745 $Y2=0.345
r208 47 49 23.4141 $w=1.78e-07 $l=3.8e-07 $layer=LI1_cond $X=5.83 $Y=0.345
+ $X2=6.21 $Y2=0.345
r209 46 58 3.71884 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.745 $Y=1.48
+ $X2=5.745 $Y2=1.645
r210 45 59 1.44715 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.745 $Y=0.435
+ $X2=5.745 $Y2=0.345
r211 45 46 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=5.745 $Y=0.435
+ $X2=5.745 $Y2=1.48
r212 43 59 5.04255 $w=1.75e-07 $l=8.74643e-08 $layer=LI1_cond $X=5.66 $Y=0.34
+ $X2=5.745 $Y2=0.345
r213 43 44 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.66 $Y=0.34
+ $X2=5.14 $Y2=0.34
r214 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.055 $Y=0.425
+ $X2=5.14 $Y2=0.34
r215 41 42 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.055 $Y=0.425
+ $X2=5.055 $Y2=0.585
r216 40 54 8.64067 $w=3.02e-07 $l=1.83916e-07 $layer=LI1_cond $X=4.245 $Y=0.675
+ $X2=4.08 $Y2=0.715
r217 39 42 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.97 $Y=0.675
+ $X2=5.055 $Y2=0.585
r218 39 40 44.6717 $w=1.78e-07 $l=7.25e-07 $layer=LI1_cond $X=4.97 $Y=0.675
+ $X2=4.245 $Y2=0.675
r219 35 37 104.747 $w=1.78e-07 $l=1.7e-06 $layer=LI1_cond $X=2.335 $Y=2.01
+ $X2=4.035 $Y2=2.01
r220 34 52 1.54918 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.335 $Y=0.795
+ $X2=2.245 $Y2=0.795
r221 33 54 8.97739 $w=3.02e-07 $l=2.0106e-07 $layer=LI1_cond $X=3.915 $Y=0.795
+ $X2=4.08 $Y2=0.715
r222 33 34 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=3.915 $Y=0.795
+ $X2=2.335 $Y2=0.795
r223 32 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.91
+ $X2=2.25 $Y2=2.075
r224 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.91 $X2=2.25 $Y2=1.91
r225 29 35 6.81649 $w=1.8e-07 $l=1.27279e-07 $layer=LI1_cond $X=2.245 $Y=1.92
+ $X2=2.335 $Y2=2.01
r226 29 31 0.616162 $w=1.78e-07 $l=1e-08 $layer=LI1_cond $X=2.245 $Y=1.92
+ $X2=2.245 $Y2=1.91
r227 28 52 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0.88
+ $X2=2.245 $Y2=0.795
r228 28 31 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=2.245 $Y=0.88
+ $X2=2.245 $Y2=1.91
r229 27 52 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0.71
+ $X2=2.245 $Y2=0.795
r230 26 27 14.1717 $w=1.78e-07 $l=2.3e-07 $layer=LI1_cond $X=2.245 $Y=0.48
+ $X2=2.245 $Y2=0.71
r231 24 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=0.34
+ $X2=1.635 $Y2=0.505
r232 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=0.34 $X2=1.635 $Y2=0.34
r233 21 26 6.92652 $w=2.25e-07 $l=1.51456e-07 $layer=LI1_cond $X=2.155 $Y=0.367
+ $X2=2.245 $Y2=0.48
r234 21 23 26.6342 $w=2.23e-07 $l=5.2e-07 $layer=LI1_cond $X=2.155 $Y=0.367
+ $X2=1.635 $Y2=0.367
r235 20 71 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.3 $Y=0.835
+ $X2=6.3 $Y2=0.515
r236 16 68 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=5.42 $Y=2.655
+ $X2=5.42 $Y2=1.81
r237 12 65 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.16 $Y=2.525
+ $X2=2.16 $Y2=2.075
r238 9 62 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.675 $Y=0.825
+ $X2=1.675 $Y2=0.505
r239 2 37 600 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.835 $X2=4.035 $Y2=2.015
r240 1 54 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.545 $X2=4.08 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%A_501_229# 1 2 9 12 14 19 22 24 28 30 35 36
+ 41 44
c105 41 0 1.76463e-19 $X=5.205 $Y=2.36
c106 36 0 8.90097e-20 $X=5.395 $Y=1.07
c107 24 0 1.16419e-19 $X=2.67 $Y=1.135
c108 12 0 1.12518e-19 $X=2.7 $Y=2.525
r109 38 41 4.75325 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=5.115 $Y=2.35
+ $X2=5.205 $Y2=2.35
r110 34 36 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.115 $Y=1.07
+ $X2=5.395 $Y2=1.07
r111 34 35 5.41468 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=5.115 $Y=1.07
+ $X2=5.025 $Y2=1.07
r112 30 32 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.42 $Y=1.02
+ $X2=4.42 $Y2=1.135
r113 28 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.31
+ $X2=2.67 $Y2=1.475
r114 28 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.31
+ $X2=2.67 $Y2=1.145
r115 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.31 $X2=2.67 $Y2=1.31
r116 24 27 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.67 $Y=1.135
+ $X2=2.67 $Y2=1.31
r117 20 36 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.395 $Y=0.935
+ $X2=5.395 $Y2=1.07
r118 20 22 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.395 $Y=0.935
+ $X2=5.395 $Y2=0.76
r119 19 38 1.64051 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=5.115 $Y=2.245
+ $X2=5.115 $Y2=2.35
r120 18 34 3.11056 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=5.115 $Y=1.205
+ $X2=5.115 $Y2=1.07
r121 18 19 64.0808 $w=1.78e-07 $l=1.04e-06 $layer=LI1_cond $X=5.115 $Y=1.205
+ $X2=5.115 $Y2=2.245
r122 17 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.505 $Y=1.02
+ $X2=4.42 $Y2=1.02
r123 17 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.505 $Y=1.02
+ $X2=5.025 $Y2=1.02
r124 15 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=1.135
+ $X2=2.67 $Y2=1.135
r125 14 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.335 $Y=1.135
+ $X2=4.42 $Y2=1.135
r126 14 15 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=4.335 $Y=1.135
+ $X2=2.835 $Y2=1.135
r127 12 45 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.7 $Y=2.525
+ $X2=2.7 $Y2=1.475
r128 9 44 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.625 $Y=0.825
+ $X2=2.625 $Y2=1.145
r129 2 41 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=5.065
+ $Y=2.235 $X2=5.205 $Y2=2.36
r130 1 22 182 $w=1.7e-07 $l=5.65442e-07 $layer=licon1_NDIFF $count=1 $X=5.095
+ $Y=0.325 $X2=5.395 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%RESET_B 4 5 6 9 13 16 20 21 23 27 32 33 34
+ 37 40 41 42 43 48 51 54 55 57 58 60 61 76
c201 32 0 1.4009e-19 $X=0.515 $Y=2.005
c202 20 0 1.8083e-19 $X=3.29 $Y=2.525
r203 60 63 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.65
+ $X2=3.21 $Y2=1.815
r204 60 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.65
+ $X2=3.21 $Y2=1.485
r205 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.21
+ $Y=1.65 $X2=3.21 $Y2=1.65
r206 58 76 1.80775 $w=2.53e-07 $l=4e-08 $layer=LI1_cond $X=7.21 $Y=1.707
+ $X2=7.17 $Y2=1.707
r207 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.21
+ $Y=1.745 $X2=7.21 $Y2=1.745
r208 55 65 5.92651 $w=5.53e-07 $l=2.75e-07 $layer=LI1_cond $X=0.515 $Y=1.842
+ $X2=0.24 $Y2=1.842
r209 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.515
+ $Y=1.65 $X2=0.515 $Y2=1.65
r210 51 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.665
r211 49 76 9.49071 $w=2.53e-07 $l=2.1e-07 $layer=LI1_cond $X=6.96 $Y=1.707
+ $X2=7.17 $Y2=1.707
r212 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.665
+ $X2=6.96 $Y2=1.665
r213 46 61 34.172 $w=1.83e-07 $l=5.7e-07 $layer=LI1_cond $X=2.64 $Y=1.657
+ $X2=3.21 $Y2=1.657
r214 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r215 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r216 42 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=1.665
+ $X2=6.96 $Y2=1.665
r217 42 43 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=6.815 $Y=1.665
+ $X2=2.785 $Y2=1.665
r218 41 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=1.665
+ $X2=0.24 $Y2=1.665
r219 40 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.495 $Y=1.665
+ $X2=2.64 $Y2=1.665
r220 40 41 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=2.495 $Y=1.665
+ $X2=0.385 $Y2=1.665
r221 37 57 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.21 $Y=2.085
+ $X2=7.21 $Y2=1.745
r222 36 57 40.0117 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.21 $Y=1.58
+ $X2=7.21 $Y2=1.745
r223 32 54 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.515 $Y=2.005
+ $X2=0.515 $Y2=1.65
r224 32 33 40.0117 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=2.005
+ $X2=0.515 $Y2=2.17
r225 30 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.485
+ $X2=0.53 $Y2=1.65
r226 27 36 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=7.25 $Y=0.835
+ $X2=7.25 $Y2=1.58
r227 21 37 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.21 $Y=2.25
+ $X2=7.21 $Y2=2.085
r228 21 23 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=7.21 $Y=2.25
+ $X2=7.21 $Y2=2.865
r229 20 34 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.29 $Y=2.525
+ $X2=3.29 $Y2=2.24
r230 18 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.29 $Y=3.075
+ $X2=3.29 $Y2=2.525
r231 16 34 45.2492 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=3.205 $Y=2.08
+ $X2=3.205 $Y2=2.24
r232 16 63 47.7863 $w=3.2e-07 $l=2.65e-07 $layer=POLY_cond $X=3.205 $Y=2.08
+ $X2=3.205 $Y2=1.815
r233 13 62 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.12 $Y=0.825
+ $X2=3.12 $Y2=1.485
r234 9 30 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.635 $Y=0.815
+ $X2=0.635 $Y2=1.485
r235 5 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.215 $Y=3.15
+ $X2=3.29 $Y2=3.075
r236 5 6 1366.52 $w=1.5e-07 $l=2.665e-06 $layer=POLY_cond $X=3.215 $Y=3.15
+ $X2=0.55 $Y2=3.15
r237 4 33 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=0.475 $Y=2.525
+ $X2=0.475 $Y2=2.17
r238 2 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=3.075
+ $X2=0.55 $Y2=3.15
r239 2 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.475 $Y=3.075
+ $X2=0.475 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%A_306_277# 1 2 9 11 12 14 16 17 18 20 21 22
+ 23 25 29 32 34 35 40 43 44 46 49 50 53 54 55 57 58 59 62 64 65 69 70 76 81 82
+ 87 90 93
c272 93 0 1.33575e-19 $X=6.047 $Y=2.165
c273 82 0 7.10242e-20 $X=6.085 $Y=2.33
c274 44 0 1.88823e-19 $X=5.2 $Y=2.71
c275 43 0 8.90097e-20 $X=4.31 $Y=1.115
c276 35 0 1.45194e-19 $X=5.685 $Y=1.195
c277 32 0 1.59204e-19 $X=5.61 $Y=0.645
c278 29 0 1.76463e-19 $X=4.31 $Y=2.28
c279 23 0 4.89731e-20 $X=4.31 $Y=1.04
c280 14 0 1.16419e-19 $X=2.115 $Y=1.11
c281 12 0 2.28752e-19 $X=1.68 $Y=1.46
c282 9 0 4.78183e-20 $X=1.605 $Y=2.525
r283 84 85 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.085 $Y=2.515
+ $X2=6.085 $Y2=2.6
r284 82 94 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=6.047 $Y=2.33
+ $X2=6.047 $Y2=2.495
r285 82 93 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=6.047 $Y=2.33
+ $X2=6.047 $Y2=2.165
r286 81 84 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=6.085 $Y=2.33
+ $X2=6.085 $Y2=2.515
r287 81 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.085
+ $Y=2.33 $X2=6.085 $Y2=2.33
r288 76 78 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.285 $Y=2.71
+ $X2=5.285 $Y2=2.85
r289 74 90 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=4.19 $Y=2.925
+ $X2=4.31 $Y2=2.925
r290 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.19
+ $Y=2.925 $X2=4.19 $Y2=2.925
r291 70 73 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.19 $Y=2.71
+ $X2=4.19 $Y2=2.925
r292 69 87 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.76 $Y=2.405
+ $X2=8.675 $Y2=2.49
r293 68 69 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=8.76 $Y=1.4
+ $X2=8.76 $Y2=2.405
r294 64 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.675 $Y=1.315
+ $X2=8.76 $Y2=1.4
r295 64 65 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=8.675 $Y=1.315
+ $X2=8.475 $Y2=1.315
r296 60 65 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=8.345 $Y=1.23
+ $X2=8.475 $Y2=1.315
r297 60 62 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=8.345 $Y=1.23
+ $X2=8.345 $Y2=1.105
r298 58 87 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.505 $Y=2.49
+ $X2=8.675 $Y2=2.49
r299 58 59 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.505 $Y=2.49
+ $X2=7.975 $Y2=2.49
r300 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.89 $Y=2.575
+ $X2=7.975 $Y2=2.49
r301 56 57 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.89 $Y=2.575
+ $X2=7.89 $Y2=2.895
r302 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.805 $Y=2.98
+ $X2=7.89 $Y2=2.895
r303 54 55 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=7.805 $Y=2.98
+ $X2=7.26 $Y2=2.98
r304 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.175 $Y=2.895
+ $X2=7.26 $Y2=2.98
r305 52 53 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.175 $Y=2.6
+ $X2=7.175 $Y2=2.895
r306 51 84 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.25 $Y=2.515
+ $X2=6.085 $Y2=2.515
r307 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.09 $Y=2.515
+ $X2=7.175 $Y2=2.6
r308 50 51 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=7.09 $Y=2.515
+ $X2=6.25 $Y2=2.515
r309 49 85 5.85086 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=6.082 $Y=2.765
+ $X2=6.082 $Y2=2.6
r310 47 78 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.37 $Y=2.85
+ $X2=5.285 $Y2=2.85
r311 46 49 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=5.92 $Y=2.85
+ $X2=6.082 $Y2=2.765
r312 46 47 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.92 $Y=2.85
+ $X2=5.37 $Y2=2.85
r313 45 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=2.71
+ $X2=4.19 $Y2=2.71
r314 44 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.2 $Y=2.71
+ $X2=5.285 $Y2=2.71
r315 44 45 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.2 $Y=2.71
+ $X2=4.355 $Y2=2.71
r316 40 94 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.07 $Y=2.865
+ $X2=6.07 $Y2=2.495
r317 36 93 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=5.92 $Y=1.27
+ $X2=5.92 $Y2=2.165
r318 34 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.845 $Y=1.195
+ $X2=5.92 $Y2=1.27
r319 34 35 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=5.845 $Y=1.195
+ $X2=5.685 $Y2=1.195
r320 30 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.61 $Y=1.12
+ $X2=5.685 $Y2=1.195
r321 30 32 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=5.61 $Y=1.12
+ $X2=5.61 $Y2=0.645
r322 27 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.31 $Y=2.76
+ $X2=4.31 $Y2=2.925
r323 27 29 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.31 $Y=2.76
+ $X2=4.31 $Y2=2.28
r324 26 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.31 $Y=1.19
+ $X2=4.31 $Y2=1.115
r325 26 29 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=4.31 $Y=1.19
+ $X2=4.31 $Y2=2.28
r326 23 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.31 $Y=1.04
+ $X2=4.31 $Y2=1.115
r327 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.31 $Y=1.04
+ $X2=4.31 $Y2=0.755
r328 21 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.235 $Y=1.115
+ $X2=4.31 $Y2=1.115
r329 21 22 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=4.235 $Y=1.115
+ $X2=3.86 $Y2=1.115
r330 20 22 28.3559 $w=1.5e-07 $l=1.45753e-07 $layer=POLY_cond $X=3.747 $Y=1.04
+ $X2=3.86 $Y2=1.115
r331 19 20 223.888 $w=2.25e-07 $l=7.85e-07 $layer=POLY_cond $X=3.747 $Y=0.255
+ $X2=3.747 $Y2=1.04
r332 17 19 28.3559 $w=1.5e-07 $l=1.4472e-07 $layer=POLY_cond $X=3.635 $Y=0.18
+ $X2=3.747 $Y2=0.255
r333 17 18 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=3.635 $Y=0.18
+ $X2=2.19 $Y2=0.18
r334 14 42 98.0041 $w=1.74e-07 $l=3.67083e-07 $layer=POLY_cond $X=2.115 $Y=1.11
+ $X2=2.08 $Y2=1.46
r335 14 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.115 $Y=1.11
+ $X2=2.115 $Y2=0.825
r336 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.115 $Y=0.255
+ $X2=2.19 $Y2=0.18
r337 13 16 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.115 $Y=0.255
+ $X2=2.115 $Y2=0.825
r338 11 42 6.34751 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.97 $Y=1.46
+ $X2=2.08 $Y2=1.46
r339 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.97 $Y=1.46
+ $X2=1.68 $Y2=1.46
r340 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.605 $Y=1.535
+ $X2=1.68 $Y2=1.46
r341 7 9 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=1.605 $Y=1.535
+ $X2=1.605 $Y2=2.525
r342 2 87 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.53
+ $Y=2.425 $X2=8.67 $Y2=2.57
r343 1 62 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=8.255
+ $Y=0.895 $X2=8.38 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%A_336_463# 1 2 3 12 16 20 22 24 28 31 40
c95 24 0 1.8083e-19 $X=4.675 $Y=2.355
c96 20 0 1.12518e-19 $X=1.89 $Y=0.84
c97 16 0 1.56182e-19 $X=5.02 $Y=0.645
r98 40 41 4.46296 $w=3.24e-07 $l=3e-08 $layer=POLY_cond $X=4.99 $Y=1.44 $X2=5.02
+ $Y2=1.44
r99 31 33 6.75433 $w=2.89e-07 $l=1.6e-07 $layer=LI1_cond $X=1.887 $Y=2.355
+ $X2=1.887 $Y2=2.515
r100 29 40 34.216 $w=3.24e-07 $l=2.3e-07 $layer=POLY_cond $X=4.76 $Y=1.44
+ $X2=4.99 $Y2=1.44
r101 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.76
+ $Y=1.44 $X2=4.76 $Y2=1.44
r102 26 28 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.76 $Y=2.27
+ $X2=4.76 $Y2=1.44
r103 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.675 $Y=2.355
+ $X2=4.76 $Y2=2.27
r104 24 25 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=4.675 $Y=2.355
+ $X2=3.645 $Y2=2.355
r105 23 31 3.84173 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.04 $Y=2.355
+ $X2=1.887 $Y2=2.355
r106 22 37 5.85368 $w=3.13e-07 $l=1.6e-07 $layer=LI1_cond $X=3.487 $Y=2.355
+ $X2=3.487 $Y2=2.515
r107 22 25 4.34843 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=3.487 $Y=2.355
+ $X2=3.645 $Y2=2.355
r108 22 23 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=3.33 $Y=2.355
+ $X2=2.04 $Y2=2.355
r109 18 31 13.1235 $w=2.89e-07 $l=2.73971e-07 $layer=LI1_cond $X=1.895 $Y=2.085
+ $X2=1.887 $Y2=2.355
r110 18 20 76.7121 $w=1.78e-07 $l=1.245e-06 $layer=LI1_cond $X=1.895 $Y=2.085
+ $X2=1.895 $Y2=0.84
r111 14 41 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.02 $Y=1.275
+ $X2=5.02 $Y2=1.44
r112 14 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=5.02 $Y=1.275
+ $X2=5.02 $Y2=0.645
r113 10 40 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.99 $Y=1.605
+ $X2=4.99 $Y2=1.44
r114 10 12 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=4.99 $Y=1.605
+ $X2=4.99 $Y2=2.655
r115 3 37 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=2.315 $X2=3.505 $Y2=2.515
r116 2 33 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=2.315 $X2=1.9 $Y2=2.515
r117 1 20 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.615 $X2=1.89 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%A_1287_276# 1 2 9 13 17 18 21 22 24 25 28 32
+ 34
c94 21 0 1.33575e-19 $X=6.6 $Y=1.545
r95 30 34 3.70735 $w=2.5e-07 $l=1.33918e-07 $layer=LI1_cond $X=7.825 $Y=1.23
+ $X2=7.727 $Y2=1.315
r96 30 32 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=7.825 $Y=1.23
+ $X2=7.825 $Y2=0.825
r97 26 34 3.70735 $w=2.5e-07 $l=2.15346e-07 $layer=LI1_cond $X=7.55 $Y=1.4
+ $X2=7.727 $Y2=1.315
r98 26 28 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=7.55 $Y=1.4
+ $X2=7.55 $Y2=2.55
r99 24 34 2.76166 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=7.465 $Y=1.315
+ $X2=7.727 $Y2=1.315
r100 24 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=7.465 $Y=1.315
+ $X2=6.685 $Y2=1.315
r101 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.6
+ $Y=1.545 $X2=6.6 $Y2=1.545
r102 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.6 $Y=1.4
+ $X2=6.685 $Y2=1.315
r103 19 21 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.6 $Y=1.4 $X2=6.6
+ $Y2=1.545
r104 17 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.6 $Y=1.885
+ $X2=6.6 $Y2=1.545
r105 17 18 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.6 $Y=1.885
+ $X2=6.6 $Y2=2.05
r106 16 22 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.6 $Y=1.38
+ $X2=6.6 $Y2=1.545
r107 13 16 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.66 $Y=0.835
+ $X2=6.66 $Y2=1.38
r108 9 18 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=6.61 $Y=2.865
+ $X2=6.61 $Y2=2.05
r109 2 28 600 $w=1.7e-07 $l=3.13129e-07 $layer=licon1_PDIFF $count=1 $X=7.285
+ $Y=2.655 $X2=7.55 $Y2=2.55
r110 1 32 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.625 $X2=7.825 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%CLK_N 3 7 9 11 18
r38 18 21 82.2934 $w=5.15e-07 $l=5.05e-07 $layer=POLY_cond $X=8.412 $Y=1.71
+ $X2=8.412 $Y2=2.215
r39 18 20 46.971 $w=5.15e-07 $l=1.65e-07 $layer=POLY_cond $X=8.412 $Y=1.71
+ $X2=8.412 $Y2=1.545
r40 11 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.32
+ $Y=1.71 $X2=8.32 $Y2=1.71
r41 9 11 7.41754 $w=6.43e-07 $l=4e-07 $layer=LI1_cond $X=7.92 $Y=1.892 $X2=8.32
+ $Y2=1.892
r42 7 20 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.595 $Y=1.105
+ $X2=8.595 $Y2=1.545
r43 3 21 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.455 $Y=2.745
+ $X2=8.455 $Y2=2.215
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%A_1099_447# 1 2 7 9 12 15 16 19 20 21 24 26
+ 28 32 34 37 41 44 45 48 49 51 54 56 60
c161 54 0 1.45194e-19 $X=5.63 $Y=2.03
c162 44 0 1.59204e-19 $X=6.085 $Y=1.905
r163 54 55 29.8441 $w=1.86e-07 $l=4.55e-07 $layer=LI1_cond $X=5.63 $Y=2.03
+ $X2=6.085 $Y2=2.03
r164 52 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.195 $Y=0.35
+ $X2=8.36 $Y2=0.35
r165 52 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.195 $Y=0.35
+ $X2=8.105 $Y2=0.35
r166 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.195
+ $Y=0.35 $X2=8.195 $Y2=0.35
r167 49 51 36.1099 $w=2.23e-07 $l=7.05e-07 $layer=LI1_cond $X=7.49 $Y=0.377
+ $X2=8.195 $Y2=0.377
r168 47 49 6.92652 $w=2.25e-07 $l=1.51456e-07 $layer=LI1_cond $X=7.4 $Y=0.49
+ $X2=7.49 $Y2=0.377
r169 47 48 24.0303 $w=1.78e-07 $l=3.9e-07 $layer=LI1_cond $X=7.4 $Y=0.49 $X2=7.4
+ $Y2=0.88
r170 46 56 1.6787 $w=1.8e-07 $l=1.13e-07 $layer=LI1_cond $X=6.225 $Y=0.97
+ $X2=6.112 $Y2=0.97
r171 45 48 6.81649 $w=1.8e-07 $l=1.27279e-07 $layer=LI1_cond $X=7.31 $Y=0.97
+ $X2=7.4 $Y2=0.88
r172 45 46 66.8535 $w=1.78e-07 $l=1.085e-06 $layer=LI1_cond $X=7.31 $Y=0.97
+ $X2=6.225 $Y2=0.97
r173 44 55 1.25915 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.085 $Y=1.905
+ $X2=6.085 $Y2=2.03
r174 43 56 4.77889 $w=1.97e-07 $l=1.02616e-07 $layer=LI1_cond $X=6.085 $Y=1.06
+ $X2=6.112 $Y2=0.97
r175 43 44 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=6.085 $Y=1.06
+ $X2=6.085 $Y2=1.905
r176 39 56 4.77889 $w=1.97e-07 $l=9e-08 $layer=LI1_cond $X=6.112 $Y=0.88
+ $X2=6.112 $Y2=0.97
r177 39 41 5.63417 $w=2.23e-07 $l=1.1e-07 $layer=LI1_cond $X=6.112 $Y=0.88
+ $X2=6.112 $Y2=0.77
r178 35 54 0.915649 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=5.63 $Y=2.155
+ $X2=5.63 $Y2=2.03
r179 35 37 16.3283 $w=1.78e-07 $l=2.65e-07 $layer=LI1_cond $X=5.63 $Y=2.155
+ $X2=5.63 $Y2=2.42
r180 31 32 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=7.87 $Y=1.23
+ $X2=8.105 $Y2=1.23
r181 29 31 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=7.61 $Y=1.23
+ $X2=7.87 $Y2=1.23
r182 26 34 20.4101 $w=1.5e-07 $l=8.87412e-08 $layer=POLY_cond $X=9.56 $Y=0.765
+ $X2=9.53 $Y2=0.84
r183 26 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.56 $Y=0.765
+ $X2=9.56 $Y2=0.445
r184 22 34 20.4101 $w=1.5e-07 $l=8.87412e-08 $layer=POLY_cond $X=9.5 $Y=0.915
+ $X2=9.53 $Y2=0.84
r185 22 24 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=9.5 $Y=0.915
+ $X2=9.5 $Y2=2.155
r186 20 34 5.30422 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=9.425 $Y=0.84
+ $X2=9.53 $Y2=0.84
r187 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.425 $Y=0.84
+ $X2=9.145 $Y2=0.84
r188 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.07 $Y=0.765
+ $X2=9.145 $Y2=0.84
r189 18 19 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=9.07 $Y=0.515
+ $X2=9.07 $Y2=0.765
r190 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.995 $Y=0.44
+ $X2=9.07 $Y2=0.515
r191 16 60 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.995 $Y=0.44
+ $X2=8.36 $Y2=0.44
r192 15 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.105 $Y=1.155
+ $X2=8.105 $Y2=1.23
r193 14 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.105 $Y=0.515
+ $X2=8.105 $Y2=0.35
r194 14 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=8.105 $Y=0.515
+ $X2=8.105 $Y2=1.155
r195 10 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.87 $Y=1.305
+ $X2=7.87 $Y2=1.23
r196 10 12 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=7.87 $Y=1.305
+ $X2=7.87 $Y2=2.635
r197 7 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.61 $Y=1.155
+ $X2=7.61 $Y2=1.23
r198 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.61 $Y=1.155
+ $X2=7.61 $Y2=0.835
r199 2 37 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=5.495
+ $Y=2.235 $X2=5.635 $Y2=2.42
r200 1 41 182 $w=1.7e-07 $l=6.13209e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.325 $X2=6.085 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%A_1832_367# 1 2 9 13 17 20 23 24 26 30
r61 28 30 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=9.345 $Y=0.445
+ $X2=9.47 $Y2=0.445
r62 24 34 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.972 $Y=1.51
+ $X2=9.972 $Y2=1.675
r63 24 33 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.972 $Y=1.51
+ $X2=9.972 $Y2=1.345
r64 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.95
+ $Y=1.51 $X2=9.95 $Y2=1.51
r65 21 26 0.260482 $w=3.3e-07 $l=4.37493e-07 $layer=LI1_cond $X=9.555 $Y=1.51
+ $X2=9.12 $Y2=1.505
r66 21 23 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=9.555 $Y=1.51
+ $X2=9.95 $Y2=1.51
r67 20 26 6.62118 $w=2.42e-07 $l=4.22493e-07 $layer=LI1_cond $X=9.47 $Y=1.345
+ $X2=9.12 $Y2=1.505
r68 19 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.47 $Y=0.61
+ $X2=9.47 $Y2=0.445
r69 19 20 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=9.47 $Y=0.61
+ $X2=9.47 $Y2=1.345
r70 15 26 6.62118 $w=2.42e-07 $l=2.35775e-07 $layer=LI1_cond $X=9.277 $Y=1.675
+ $X2=9.12 $Y2=1.505
r71 15 17 11.1586 $w=3.13e-07 $l=3.05e-07 $layer=LI1_cond $X=9.277 $Y=1.675
+ $X2=9.277 $Y2=1.98
r72 13 34 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.085 $Y=2.465
+ $X2=10.085 $Y2=1.675
r73 9 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=10.085 $Y=0.655
+ $X2=10.085 $Y2=1.345
r74 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=9.16
+ $Y=1.835 $X2=9.285 $Y2=1.98
r75 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.22
+ $Y=0.235 $X2=9.345 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%A_27_463# 1 2 3 10 13 16 24 26 27
c59 24 0 1.97962e-19 $X=1.55 $Y=0.815
c60 13 0 1.75901e-19 $X=1.362 $Y=2.29
c61 10 0 4.78183e-20 $X=1.16 $Y=2.375
r62 26 27 11.2298 $w=4.03e-07 $l=2.55e-07 $layer=LI1_cond $X=1.397 $Y=1.565
+ $X2=1.397 $Y2=1.82
r63 22 24 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.315 $Y=0.815
+ $X2=1.55 $Y2=0.815
r64 16 19 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.285 $Y=2.375
+ $X2=0.285 $Y2=2.525
r65 14 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=0.98
+ $X2=1.55 $Y2=0.815
r66 14 26 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.55 $Y=0.98
+ $X2=1.55 $Y2=1.565
r67 13 27 13.374 $w=4.03e-07 $l=4.7e-07 $layer=LI1_cond $X=1.362 $Y=2.29
+ $X2=1.362 $Y2=1.82
r68 11 16 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.47 $Y=2.375
+ $X2=0.285 $Y2=2.375
r69 10 30 5.5488 $w=4.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.362 $Y=2.375
+ $X2=1.362 $Y2=2.57
r70 10 13 2.41871 $w=4.03e-07 $l=8.5e-08 $layer=LI1_cond $X=1.362 $Y=2.375
+ $X2=1.362 $Y2=2.29
r71 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.16 $Y=2.375
+ $X2=0.47 $Y2=2.375
r72 3 30 600 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=1.21
+ $Y=2.315 $X2=1.35 $Y2=2.57
r73 2 19 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.315 $X2=0.26 $Y2=2.525
r74 1 22 182 $w=1.7e-07 $l=3.33879e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.605 $X2=1.315 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%VPWR 1 2 3 4 5 6 23 27 29 33 37 41 46 47 49
+ 50 51 53 74 83 84 87 90 93 100
c113 84 0 7.10242e-20 $X=10.32 $Y=3.33
r114 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r115 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 93 96 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.69 $Y=3.06
+ $X2=4.69 $Y2=3.33
r117 91 97 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r119 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 84 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r121 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r122 81 100 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=9.975 $Y=3.33
+ $X2=9.79 $Y2=3.33
r123 81 83 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.975 $Y=3.33
+ $X2=10.32 $Y2=3.33
r124 80 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r125 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r126 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r127 76 79 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33 $X2=9.36
+ $Y2=3.33
r128 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r129 74 100 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.79 $Y2=3.33
r130 74 79 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.36 $Y2=3.33
r131 73 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r132 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r133 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 69 72 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r135 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r136 67 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r137 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r138 64 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r139 63 66 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r140 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r141 61 96 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.69 $Y2=3.33
r142 61 63 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=5.04 $Y2=3.33
r143 60 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r144 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r145 57 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r146 57 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 56 59 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r148 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r149 54 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.805 $Y2=3.33
r150 54 56 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.2 $Y2=3.33
r151 53 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=2.995 $Y2=3.33
r152 53 59 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=2.64 $Y2=3.33
r153 51 67 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=6.48 $Y2=3.33
r154 51 64 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r155 49 72 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.145 $Y=3.33
+ $X2=7.92 $Y2=3.33
r156 49 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.145 $Y=3.33
+ $X2=8.24 $Y2=3.33
r157 48 76 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=8.335 $Y=3.33
+ $X2=8.4 $Y2=3.33
r158 48 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.335 $Y=3.33
+ $X2=8.24 $Y2=3.33
r159 46 66 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r160 46 47 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.72 $Y=3.33 $X2=6.82
+ $Y2=3.33
r161 45 69 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=6.92 $Y=3.33 $X2=6.96
+ $Y2=3.33
r162 45 47 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.92 $Y=3.33 $X2=6.82
+ $Y2=3.33
r163 41 44 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=9.79 $Y=1.98
+ $X2=9.79 $Y2=2.46
r164 39 100 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.79 $Y=3.245
+ $X2=9.79 $Y2=3.33
r165 39 44 24.4505 $w=3.68e-07 $l=7.85e-07 $layer=LI1_cond $X=9.79 $Y=3.245
+ $X2=9.79 $Y2=2.46
r166 35 50 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.24 $Y=3.245
+ $X2=8.24 $Y2=3.33
r167 35 37 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=8.24 $Y=3.245
+ $X2=8.24 $Y2=2.92
r168 31 47 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=3.245
+ $X2=6.82 $Y2=3.33
r169 31 33 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=6.82 $Y=3.245
+ $X2=6.82 $Y2=2.95
r170 30 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=3.33
+ $X2=2.995 $Y2=3.33
r171 29 96 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.69 $Y2=3.33
r172 29 30 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=3.16 $Y2=3.33
r173 25 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=3.33
r174 25 27 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=2.705
r175 21 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.33
r176 21 23 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=2.725
r177 6 44 300 $w=1.7e-07 $l=7.58288e-07 $layer=licon1_PDIFF $count=2 $X=9.575
+ $Y=1.835 $X2=9.87 $Y2=2.46
r178 6 41 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=9.575
+ $Y=1.835 $X2=9.77 $Y2=1.98
r179 5 37 600 $w=1.7e-07 $l=6.2534e-07 $layer=licon1_PDIFF $count=1 $X=7.945
+ $Y=2.425 $X2=8.24 $Y2=2.92
r180 4 33 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=6.685
+ $Y=2.655 $X2=6.825 $Y2=2.95
r181 3 93 600 $w=1.7e-07 $l=1.24318e-06 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.96 $X2=4.69 $Y2=3.06
r182 2 27 600 $w=1.7e-07 $l=4.8775e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=2.315 $X2=2.995 $Y2=2.705
r183 1 23 600 $w=1.7e-07 $l=5.22159e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.315 $X2=0.805 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%Q 1 2 7 8 9 10 11 12 13 25 31 41
r18 23 31 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=10.315 $Y=0.93
+ $X2=10.315 $Y2=0.925
r19 13 48 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=10.31 $Y=2.775
+ $X2=10.31 $Y2=2.91
r20 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.31 $Y=2.405
+ $X2=10.31 $Y2=2.775
r21 11 41 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=10.31 $Y=1.98
+ $X2=10.31 $Y2=2.01
r22 11 53 5.12956 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=10.31 $Y=1.98
+ $X2=10.31 $Y2=1.845
r23 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=10.31 $Y=2.065
+ $X2=10.31 $Y2=2.405
r24 11 41 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=10.31 $Y=2.065
+ $X2=10.31 $Y2=2.01
r25 10 53 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.34 $Y=1.665
+ $X2=10.34 $Y2=1.845
r26 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.34 $Y=1.295
+ $X2=10.34 $Y2=1.665
r27 9 51 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=10.34 $Y=1.295
+ $X2=10.34 $Y2=1.09
r28 8 51 4.63652 $w=3.18e-07 $l=1.2e-07 $layer=LI1_cond $X=10.315 $Y=0.97
+ $X2=10.315 $Y2=1.09
r29 8 23 1.44055 $w=3.18e-07 $l=4e-08 $layer=LI1_cond $X=10.315 $Y=0.97
+ $X2=10.315 $Y2=0.93
r30 8 31 1.44055 $w=3.18e-07 $l=4e-08 $layer=LI1_cond $X=10.315 $Y=0.885
+ $X2=10.315 $Y2=0.925
r31 7 8 11.8846 $w=3.18e-07 $l=3.3e-07 $layer=LI1_cond $X=10.315 $Y=0.555
+ $X2=10.315 $Y2=0.885
r32 7 25 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=10.315 $Y=0.555
+ $X2=10.315 $Y2=0.42
r33 2 48 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.835 $X2=10.3 $Y2=2.91
r34 2 41 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.835 $X2=10.3 $Y2=2.01
r35 1 25 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=10.16
+ $Y=0.235 $X2=10.3 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTN_1%VGND 1 2 3 4 5 6 19 21 25 29 32 35 40 41 43
+ 44 48 57 61 76 82 83 90 96 99
r129 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r130 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r131 90 93 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.635 $Y=0
+ $X2=4.635 $Y2=0.32
r132 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r133 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r134 83 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r135 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r136 80 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.985 $Y=0 $X2=9.855
+ $Y2=0
r137 80 82 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=10.32 $Y2=0
r138 79 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r139 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r140 76 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.725 $Y=0 $X2=9.855
+ $Y2=0
r141 76 78 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.725 $Y=0
+ $X2=9.36 $Y2=0
r142 75 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r143 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r144 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r145 72 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r146 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r147 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r148 69 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.12 $Y=0 $X2=6.955
+ $Y2=0
r149 69 71 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.12 $Y=0 $X2=7.44
+ $Y2=0
r150 68 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r151 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r152 65 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r153 64 67 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r154 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r155 62 90 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=4.635
+ $Y2=0
r156 62 64 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r157 61 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.79 $Y=0 $X2=6.955
+ $Y2=0
r158 61 67 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.79 $Y=0 $X2=6.48
+ $Y2=0
r159 60 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r160 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r161 57 90 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.635
+ $Y2=0
r162 57 59 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.08
+ $Y2=0
r163 56 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r164 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r165 53 56 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.72 $Y=0 $X2=3.12
+ $Y2=0
r166 53 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r167 52 55 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=3.12
+ $Y2=0
r168 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r169 50 86 4.49701 $w=1.7e-07 $l=2.93e-07 $layer=LI1_cond $X=0.585 $Y=0
+ $X2=0.292 $Y2=0
r170 50 52 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.585 $Y=0
+ $X2=0.72 $Y2=0
r171 48 68 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=6.48
+ $Y2=0
r172 48 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.04 $Y2=0
r173 43 74 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.76 $Y=0 $X2=8.4
+ $Y2=0
r174 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=0 $X2=8.845
+ $Y2=0
r175 42 78 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.93 $Y=0 $X2=9.36
+ $Y2=0
r176 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.93 $Y=0 $X2=8.845
+ $Y2=0
r177 40 55 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.12
+ $Y2=0
r178 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.415
+ $Y2=0
r179 39 59 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=4.08
+ $Y2=0
r180 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=3.415
+ $Y2=0
r181 35 37 24.157 $w=2.58e-07 $l=5.45e-07 $layer=LI1_cond $X=9.855 $Y=0.38
+ $X2=9.855 $Y2=0.925
r182 33 99 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.855 $Y=0.085
+ $X2=9.855 $Y2=0
r183 33 35 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=9.855 $Y=0.085
+ $X2=9.855 $Y2=0.38
r184 32 47 10.9542 $w=2.84e-07 $l=4.08044e-07 $layer=LI1_cond $X=8.845 $Y=0.89
+ $X2=9.1 $Y2=1.19
r185 31 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.845 $Y=0.085
+ $X2=8.845 $Y2=0
r186 31 32 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=8.845 $Y=0.085
+ $X2=8.845 $Y2=0.89
r187 27 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0.085
+ $X2=6.955 $Y2=0
r188 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=6.955 $Y=0.085
+ $X2=6.955 $Y2=0.615
r189 23 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=0.085
+ $X2=3.415 $Y2=0
r190 23 25 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.415 $Y=0.085
+ $X2=3.415 $Y2=0.455
r191 19 86 3.26916 $w=3.3e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.42 $Y=0.085
+ $X2=0.292 $Y2=0
r192 19 21 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=0.42 $Y=0.085
+ $X2=0.42 $Y2=0.815
r193 6 37 182 $w=1.7e-07 $l=7.98906e-07 $layer=licon1_NDIFF $count=1 $X=9.635
+ $Y=0.235 $X2=9.87 $Y2=0.925
r194 6 35 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=9.635
+ $Y=0.235 $X2=9.835 $Y2=0.38
r195 5 47 182 $w=1.7e-07 $l=5.44702e-07 $layer=licon1_NDIFF $count=1 $X=8.67
+ $Y=0.895 $X2=9.1 $Y2=1.155
r196 4 29 182 $w=1.7e-07 $l=2.24944e-07 $layer=licon1_NDIFF $count=1 $X=6.735
+ $Y=0.625 $X2=6.955 $Y2=0.615
r197 3 93 182 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.545 $X2=4.635 $Y2=0.32
r198 2 25 182 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.615 $X2=3.415 $Y2=0.455
r199 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.295
+ $Y=0.605 $X2=0.42 $Y2=0.815
.ends

