* File: sky130_fd_sc_lp__sdfbbn_2.pxi.spice
* Created: Fri Aug 28 11:27:21 2020
* 
x_PM_SKY130_FD_SC_LP__SDFBBN_2%SCD N_SCD_c_350_n N_SCD_M1013_g N_SCD_c_355_n
+ N_SCD_M1048_g N_SCD_c_357_n N_SCD_c_358_n SCD N_SCD_c_352_n N_SCD_c_353_n
+ PM_SKY130_FD_SC_LP__SDFBBN_2%SCD
x_PM_SKY130_FD_SC_LP__SDFBBN_2%D N_D_M1019_g N_D_M1051_g N_D_c_387_n N_D_c_388_n
+ N_D_c_389_n D D D N_D_c_391_n PM_SKY130_FD_SC_LP__SDFBBN_2%D
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_407_93# N_A_407_93#_M1016_d N_A_407_93#_M1028_d
+ N_A_407_93#_M1004_g N_A_407_93#_c_439_n N_A_407_93#_M1015_g
+ N_A_407_93#_c_435_n N_A_407_93#_c_436_n N_A_407_93#_c_437_n
+ N_A_407_93#_c_442_n N_A_407_93#_c_443_n N_A_407_93#_c_444_n
+ N_A_407_93#_c_438_n PM_SKY130_FD_SC_LP__SDFBBN_2%A_407_93#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%SCE N_SCE_M1036_g N_SCE_c_504_n N_SCE_c_505_n
+ N_SCE_c_506_n N_SCE_M1050_g N_SCE_M1016_g N_SCE_M1028_g N_SCE_c_515_n
+ N_SCE_c_509_n SCE N_SCE_c_511_n PM_SKY130_FD_SC_LP__SDFBBN_2%SCE
x_PM_SKY130_FD_SC_LP__SDFBBN_2%CLK_N N_CLK_N_M1049_g N_CLK_N_M1025_g
+ N_CLK_N_c_578_n N_CLK_N_c_579_n CLK_N CLK_N N_CLK_N_c_581_n
+ PM_SKY130_FD_SC_LP__SDFBBN_2%CLK_N
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_840_95# N_A_840_95#_M1049_d N_A_840_95#_M1025_d
+ N_A_840_95#_M1010_g N_A_840_95#_M1008_g N_A_840_95#_c_612_n
+ N_A_840_95#_c_613_n N_A_840_95#_c_631_n N_A_840_95#_c_632_n
+ N_A_840_95#_M1042_g N_A_840_95#_M1044_g N_A_840_95#_M1022_g
+ N_A_840_95#_c_634_n N_A_840_95#_M1009_g N_A_840_95#_c_615_n
+ N_A_840_95#_c_616_n N_A_840_95#_c_637_n N_A_840_95#_c_617_n
+ N_A_840_95#_c_618_n N_A_840_95#_c_619_n N_A_840_95#_c_620_n
+ N_A_840_95#_c_656_p N_A_840_95#_c_817_p N_A_840_95#_c_621_n
+ N_A_840_95#_c_622_n N_A_840_95#_c_623_n N_A_840_95#_c_624_n
+ N_A_840_95#_c_625_n N_A_840_95#_c_626_n N_A_840_95#_c_639_n
+ N_A_840_95#_c_640_n N_A_840_95#_c_641_n N_A_840_95#_c_642_n
+ N_A_840_95#_c_643_n N_A_840_95#_c_627_n N_A_840_95#_c_628_n
+ N_A_840_95#_c_629_n PM_SKY130_FD_SC_LP__SDFBBN_2%A_840_95#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_1423_401# N_A_1423_401#_M1029_d
+ N_A_1423_401#_M1043_d N_A_1423_401#_M1018_g N_A_1423_401#_M1017_g
+ N_A_1423_401#_M1046_g N_A_1423_401#_M1039_g N_A_1423_401#_c_832_n
+ N_A_1423_401#_c_833_n N_A_1423_401#_c_834_n N_A_1423_401#_c_843_n
+ N_A_1423_401#_c_844_n N_A_1423_401#_c_845_n N_A_1423_401#_c_835_n
+ N_A_1423_401#_c_836_n N_A_1423_401#_c_837_n N_A_1423_401#_c_838_n
+ N_A_1423_401#_c_848_n PM_SKY130_FD_SC_LP__SDFBBN_2%A_1423_401#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%SET_B N_SET_B_c_954_n N_SET_B_M1021_g
+ N_SET_B_M1043_g N_SET_B_M1030_g N_SET_B_c_965_n N_SET_B_c_966_n
+ N_SET_B_M1023_g N_SET_B_c_967_n SET_B N_SET_B_c_956_n N_SET_B_c_957_n
+ N_SET_B_c_958_n N_SET_B_c_959_n N_SET_B_c_960_n N_SET_B_c_961_n
+ N_SET_B_c_962_n N_SET_B_c_963_n PM_SKY130_FD_SC_LP__SDFBBN_2%SET_B
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_1273_137# N_A_1273_137#_M1011_d
+ N_A_1273_137#_M1042_d N_A_1273_137#_M1029_g N_A_1273_137#_M1033_g
+ N_A_1273_137#_c_1087_n N_A_1273_137#_c_1095_n N_A_1273_137#_c_1096_n
+ N_A_1273_137#_c_1097_n N_A_1273_137#_c_1088_n N_A_1273_137#_c_1089_n
+ N_A_1273_137#_c_1098_n N_A_1273_137#_c_1090_n N_A_1273_137#_c_1091_n
+ N_A_1273_137#_c_1100_n N_A_1273_137#_c_1092_n
+ PM_SKY130_FD_SC_LP__SDFBBN_2%A_1273_137#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_978_67# N_A_978_67#_M1010_s N_A_978_67#_M1008_s
+ N_A_978_67#_c_1206_n N_A_978_67#_c_1207_n N_A_978_67#_M1011_g
+ N_A_978_67#_c_1209_n N_A_978_67#_M1045_g N_A_978_67#_c_1211_n
+ N_A_978_67#_c_1212_n N_A_978_67#_M1020_g N_A_978_67#_c_1214_n
+ N_A_978_67#_c_1215_n N_A_978_67#_c_1198_n N_A_978_67#_c_1199_n
+ N_A_978_67#_c_1200_n N_A_978_67#_c_1201_n N_A_978_67#_M1007_g
+ N_A_978_67#_c_1217_n N_A_978_67#_c_1202_n N_A_978_67#_c_1219_n
+ N_A_978_67#_c_1203_n N_A_978_67#_c_1204_n N_A_978_67#_c_1205_n
+ PM_SKY130_FD_SC_LP__SDFBBN_2%A_978_67#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_2415_137# N_A_2415_137#_M1047_d
+ N_A_2415_137#_M1023_d N_A_2415_137#_c_1329_n N_A_2415_137#_M1037_g
+ N_A_2415_137#_M1035_g N_A_2415_137#_M1001_g N_A_2415_137#_M1012_g
+ N_A_2415_137#_c_1332_n N_A_2415_137#_M1024_g N_A_2415_137#_M1041_g
+ N_A_2415_137#_c_1335_n N_A_2415_137#_c_1336_n N_A_2415_137#_c_1337_n
+ N_A_2415_137#_c_1338_n N_A_2415_137#_c_1339_n N_A_2415_137#_c_1353_n
+ N_A_2415_137#_c_1354_n N_A_2415_137#_M1038_g N_A_2415_137#_c_1355_n
+ N_A_2415_137#_M1006_g N_A_2415_137#_c_1341_n N_A_2415_137#_c_1342_n
+ N_A_2415_137#_c_1343_n N_A_2415_137#_c_1356_n N_A_2415_137#_c_1397_p
+ N_A_2415_137#_c_1412_p N_A_2415_137#_c_1344_n N_A_2415_137#_c_1358_n
+ N_A_2415_137#_c_1345_n N_A_2415_137#_c_1360_n N_A_2415_137#_c_1361_n
+ N_A_2415_137#_c_1362_n N_A_2415_137#_c_1392_n N_A_2415_137#_c_1409_p
+ N_A_2415_137#_c_1418_p N_A_2415_137#_c_1346_n N_A_2415_137#_c_1347_n
+ N_A_2415_137#_c_1348_n PM_SKY130_FD_SC_LP__SDFBBN_2%A_2415_137#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_2211_428# N_A_2211_428#_M1022_d
+ N_A_2211_428#_M1020_d N_A_2211_428#_M1047_g N_A_2211_428#_M1000_g
+ N_A_2211_428#_c_1563_n N_A_2211_428#_c_1536_n N_A_2211_428#_c_1542_n
+ N_A_2211_428#_c_1537_n N_A_2211_428#_c_1538_n N_A_2211_428#_c_1539_n
+ N_A_2211_428#_c_1540_n PM_SKY130_FD_SC_LP__SDFBBN_2%A_2211_428#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_1840_21# N_A_1840_21#_M1032_s
+ N_A_1840_21#_M1040_s N_A_1840_21#_M1014_g N_A_1840_21#_M1005_g
+ N_A_1840_21#_c_1627_n N_A_1840_21#_c_1628_n N_A_1840_21#_M1031_g
+ N_A_1840_21#_M1026_g N_A_1840_21#_c_1630_n N_A_1840_21#_c_1631_n
+ N_A_1840_21#_c_1632_n N_A_1840_21#_c_1633_n N_A_1840_21#_c_1634_n
+ N_A_1840_21#_c_1639_n N_A_1840_21#_c_1640_n N_A_1840_21#_c_1635_n
+ PM_SKY130_FD_SC_LP__SDFBBN_2%A_1840_21#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%RESET_B N_RESET_B_c_1735_n N_RESET_B_M1040_g
+ N_RESET_B_M1032_g RESET_B N_RESET_B_c_1737_n
+ PM_SKY130_FD_SC_LP__SDFBBN_2%RESET_B
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_3289_47# N_A_3289_47#_M1038_s
+ N_A_3289_47#_M1006_s N_A_3289_47#_c_1773_n N_A_3289_47#_M1003_g
+ N_A_3289_47#_M1002_g N_A_3289_47#_c_1775_n N_A_3289_47#_c_1776_n
+ N_A_3289_47#_M1027_g N_A_3289_47#_M1034_g N_A_3289_47#_c_1778_n
+ N_A_3289_47#_c_1779_n N_A_3289_47#_c_1780_n N_A_3289_47#_c_1781_n
+ N_A_3289_47#_c_1782_n N_A_3289_47#_c_1783_n
+ PM_SKY130_FD_SC_LP__SDFBBN_2%A_3289_47#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_56_481# N_A_56_481#_M1048_s N_A_56_481#_M1015_d
+ N_A_56_481#_c_1839_n N_A_56_481#_c_1840_n N_A_56_481#_c_1841_n
+ N_A_56_481#_c_1842_n N_A_56_481#_c_1843_n N_A_56_481#_c_1844_n
+ N_A_56_481#_c_1845_n PM_SKY130_FD_SC_LP__SDFBBN_2%A_56_481#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%VPWR N_VPWR_M1048_d N_VPWR_M1028_s N_VPWR_M1025_s
+ N_VPWR_M1008_d N_VPWR_M1018_d N_VPWR_M1005_d N_VPWR_M1035_d N_VPWR_M1026_d
+ N_VPWR_M1040_d N_VPWR_M1024_d N_VPWR_M1006_d N_VPWR_M1034_s N_VPWR_c_1890_n
+ N_VPWR_c_1891_n N_VPWR_c_1892_n N_VPWR_c_1893_n N_VPWR_c_1894_n
+ N_VPWR_c_1895_n N_VPWR_c_1896_n N_VPWR_c_1897_n N_VPWR_c_1898_n
+ N_VPWR_c_1899_n N_VPWR_c_1900_n N_VPWR_c_1901_n N_VPWR_c_1902_n
+ N_VPWR_c_1903_n N_VPWR_c_1904_n N_VPWR_c_1905_n N_VPWR_c_1906_n
+ N_VPWR_c_1907_n N_VPWR_c_1908_n N_VPWR_c_1909_n N_VPWR_c_1910_n
+ N_VPWR_c_1911_n N_VPWR_c_1912_n VPWR N_VPWR_c_1913_n N_VPWR_c_1914_n
+ N_VPWR_c_1915_n N_VPWR_c_1916_n N_VPWR_c_1917_n N_VPWR_c_1918_n
+ N_VPWR_c_1919_n N_VPWR_c_1920_n N_VPWR_c_1921_n N_VPWR_c_1922_n
+ N_VPWR_c_1923_n N_VPWR_c_1924_n N_VPWR_c_1925_n N_VPWR_c_1889_n
+ PM_SKY130_FD_SC_LP__SDFBBN_2%VPWR
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_202_119# N_A_202_119#_M1036_d
+ N_A_202_119#_M1011_s N_A_202_119#_M1051_d N_A_202_119#_M1042_s
+ N_A_202_119#_c_2083_n N_A_202_119#_c_2084_n N_A_202_119#_c_2085_n
+ N_A_202_119#_c_2089_n N_A_202_119#_c_2086_n N_A_202_119#_c_2091_n
+ N_A_202_119#_c_2092_n N_A_202_119#_c_2093_n N_A_202_119#_c_2094_n
+ N_A_202_119#_c_2147_n N_A_202_119#_c_2148_n N_A_202_119#_c_2087_n
+ N_A_202_119#_c_2096_n N_A_202_119#_c_2088_n N_A_202_119#_c_2097_n
+ N_A_202_119#_c_2098_n PM_SKY130_FD_SC_LP__SDFBBN_2%A_202_119#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%Q_N N_Q_N_M1012_s N_Q_N_M1001_s N_Q_N_c_2231_n
+ N_Q_N_c_2232_n Q_N Q_N Q_N Q_N N_Q_N_c_2233_n PM_SKY130_FD_SC_LP__SDFBBN_2%Q_N
x_PM_SKY130_FD_SC_LP__SDFBBN_2%Q N_Q_M1003_d N_Q_M1002_d Q Q Q Q Q Q Q
+ N_Q_c_2270_n PM_SKY130_FD_SC_LP__SDFBBN_2%Q
x_PM_SKY130_FD_SC_LP__SDFBBN_2%VGND N_VGND_M1013_s N_VGND_M1004_d N_VGND_M1049_s
+ N_VGND_M1010_d N_VGND_M1017_d N_VGND_M1046_s N_VGND_M1037_d N_VGND_M1032_d
+ N_VGND_M1041_d N_VGND_M1038_d N_VGND_M1027_s N_VGND_c_2290_n N_VGND_c_2291_n
+ N_VGND_c_2292_n N_VGND_c_2293_n N_VGND_c_2294_n N_VGND_c_2295_n
+ N_VGND_c_2296_n N_VGND_c_2297_n N_VGND_c_2298_n N_VGND_c_2299_n
+ N_VGND_c_2300_n N_VGND_c_2301_n N_VGND_c_2302_n N_VGND_c_2303_n
+ N_VGND_c_2304_n N_VGND_c_2305_n N_VGND_c_2306_n N_VGND_c_2307_n
+ N_VGND_c_2308_n VGND N_VGND_c_2309_n N_VGND_c_2310_n N_VGND_c_2311_n
+ N_VGND_c_2312_n N_VGND_c_2313_n N_VGND_c_2314_n N_VGND_c_2315_n
+ N_VGND_c_2316_n N_VGND_c_2317_n N_VGND_c_2318_n N_VGND_c_2319_n
+ N_VGND_c_2320_n N_VGND_c_2321_n N_VGND_c_2322_n
+ PM_SKY130_FD_SC_LP__SDFBBN_2%VGND
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_1670_93# N_A_1670_93#_M1021_d
+ N_A_1670_93#_M1014_d N_A_1670_93#_c_2482_n N_A_1670_93#_c_2483_n
+ N_A_1670_93#_c_2481_n PM_SKY130_FD_SC_LP__SDFBBN_2%A_1670_93#
x_PM_SKY130_FD_SC_LP__SDFBBN_2%A_2574_119# N_A_2574_119#_M1030_d
+ N_A_2574_119#_M1031_d N_A_2574_119#_c_2507_n N_A_2574_119#_c_2508_n
+ N_A_2574_119#_c_2509_n PM_SKY130_FD_SC_LP__SDFBBN_2%A_2574_119#
cc_1 VNB N_SCD_c_350_n 0.0212702f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.685
cc_2 VNB N_SCD_M1013_g 0.0281566f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.805
cc_3 VNB N_SCD_c_352_n 0.0242818f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_4 VNB N_SCD_c_353_n 0.0190682f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_5 VNB N_D_c_387_n 0.0147994f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.275
cc_6 VNB N_D_c_388_n 0.0259253f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.725
cc_7 VNB N_D_c_389_n 0.00194589f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.725
cc_8 VNB D 7.03048e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_D_c_391_n 0.0197348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_407_93#_M1004_g 0.0203203f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.275
cc_11 VNB N_A_407_93#_c_435_n 0.0332208f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_A_407_93#_c_436_n 0.00241733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_407_93#_c_437_n 0.016727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_407_93#_c_438_n 0.019454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_M1036_g 0.0307843f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.805
cc_16 VNB N_SCE_c_504_n 0.017547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_SCE_c_505_n 0.143145f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.885
cc_18 VNB N_SCE_c_506_n 0.0125534f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.125
cc_19 VNB N_SCE_M1016_g 0.0299592f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.2
cc_20 VNB N_SCE_M1028_g 0.0071187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_SCE_c_509_n 0.0228881f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.55
cc_22 VNB SCE 0.00354856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_SCE_c_511_n 0.0180407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_CLK_N_M1049_g 0.0271407f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.215
cc_25 VNB N_CLK_N_c_578_n 0.0276616f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.725
cc_26 VNB N_CLK_N_c_579_n 0.00327296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB CLK_N 0.00348574f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.885
cc_28 VNB N_CLK_N_c_581_n 0.0186137f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_A_840_95#_M1010_g 0.0210246f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.725
cc_30 VNB N_A_840_95#_c_612_n 0.106824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_840_95#_c_613_n 0.0127422f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.2
cc_32 VNB N_A_840_95#_M1044_g 0.0415173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_840_95#_c_615_n 0.0883737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_840_95#_c_616_n 0.0275393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_840_95#_c_617_n 0.0291997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_840_95#_c_618_n 0.00325837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_840_95#_c_619_n 0.00326772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_840_95#_c_620_n 0.0395447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_840_95#_c_621_n 5.73082e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_840_95#_c_622_n 0.0335298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_840_95#_c_623_n 0.00317033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_840_95#_c_624_n 0.0165345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_840_95#_c_625_n 0.00767352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_840_95#_c_626_n 0.00346876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_840_95#_c_627_n 0.00379887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_840_95#_c_628_n 0.0241541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_840_95#_c_629_n 0.0186391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1423_401#_M1017_g 0.0514723f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.885
cc_49 VNB N_A_1423_401#_M1046_g 0.0223961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1423_401#_c_832_n 0.00174989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1423_401#_c_833_n 0.00190422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1423_401#_c_834_n 2.39447e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1423_401#_c_835_n 0.0010669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1423_401#_c_836_n 0.00149185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1423_401#_c_837_n 0.0293337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1423_401#_c_838_n 0.0299437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_SET_B_c_954_n 0.0200796f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.415
cc_58 VNB N_SET_B_M1043_g 0.00620931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_SET_B_c_956_n 0.0395482f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_60 VNB N_SET_B_c_957_n 0.00258354f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.215
cc_61 VNB N_SET_B_c_958_n 0.00183115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_SET_B_c_959_n 0.00567914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_SET_B_c_960_n 0.0358053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_SET_B_c_961_n 0.00588303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_SET_B_c_962_n 0.0253305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_SET_B_c_963_n 0.0162541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1273_137#_M1029_g 0.0262315f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.275
cc_68 VNB N_A_1273_137#_c_1087_n 0.0122872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1273_137#_c_1088_n 0.0116565f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.55
cc_70 VNB N_A_1273_137#_c_1089_n 0.00368511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1273_137#_c_1090_n 0.00146693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1273_137#_c_1091_n 0.0225964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1273_137#_c_1092_n 0.00553839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_978_67#_M1011_g 0.0410057f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.725
cc_75 VNB N_A_978_67#_c_1198_n 0.0142017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_978_67#_c_1199_n 0.0273057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_978_67#_c_1200_n 0.00826908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_978_67#_c_1201_n 0.0155461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_978_67#_c_1202_n 0.00545727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_978_67#_c_1203_n 0.00875881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_978_67#_c_1204_n 0.0334719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_978_67#_c_1205_n 0.0103785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2415_137#_c_1329_n 0.0152179f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=1.885
cc_84 VNB N_A_2415_137#_M1001_g 9.39904e-19 $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_85 VNB N_A_2415_137#_M1012_g 0.0240097f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_86 VNB N_A_2415_137#_c_1332_n 0.0116657f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.55
cc_87 VNB N_A_2415_137#_M1024_g 0.00957381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_2415_137#_M1041_g 0.0231592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2415_137#_c_1335_n 0.016058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2415_137#_c_1336_n 0.0195662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2415_137#_c_1337_n 0.0119732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2415_137#_c_1338_n 0.0345071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2415_137#_c_1339_n 0.0118257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2415_137#_M1038_g 0.0228988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2415_137#_c_1341_n 0.023523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2415_137#_c_1342_n 0.0024675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2415_137#_c_1343_n 0.00650699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2415_137#_c_1344_n 0.00294146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2415_137#_c_1345_n 2.14969e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2415_137#_c_1346_n 0.00269692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2415_137#_c_1347_n 0.0156068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2415_137#_c_1348_n 0.0290506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2211_428#_M1047_g 0.0238237f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=2.275
cc_104 VNB N_A_2211_428#_c_1536_n 0.0032813f $X=-0.19 $Y=-0.245 $X2=0.42
+ $Y2=1.38
cc_105 VNB N_A_2211_428#_c_1537_n 0.00286394f $X=-0.19 $Y=-0.245 $X2=0.42
+ $Y2=1.215
cc_106 VNB N_A_2211_428#_c_1538_n 0.0109104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2211_428#_c_1539_n 0.00128675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2211_428#_c_1540_n 0.0221677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1840_21#_M1014_g 0.0189173f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.725
cc_110 VNB N_A_1840_21#_M1005_g 0.0210906f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.885
cc_111 VNB N_A_1840_21#_c_1627_n 0.347173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1840_21#_c_1628_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.2
cc_113 VNB N_A_1840_21#_M1031_g 0.0113441f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.38
cc_114 VNB N_A_1840_21#_c_1630_n 0.0112574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1840_21#_c_1631_n 0.00989567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_1840_21#_c_1632_n 0.0293833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_1840_21#_c_1633_n 0.00412838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_1840_21#_c_1634_n 0.0362938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_1840_21#_c_1635_n 0.00833607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_RESET_B_c_1735_n 0.0261817f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.415
cc_121 VNB N_RESET_B_M1032_g 0.028832f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.885
cc_122 VNB N_RESET_B_c_1737_n 0.00435583f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.885
cc_123 VNB N_A_3289_47#_c_1773_n 0.0173121f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=1.885
cc_124 VNB N_A_3289_47#_M1002_g 0.007943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_3289_47#_c_1775_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.2
cc_126 VNB N_A_3289_47#_c_1776_n 0.0210934f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.2
cc_127 VNB N_A_3289_47#_M1034_g 0.0243375f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_128 VNB N_A_3289_47#_c_1778_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0.42
+ $Y2=1.215
cc_129 VNB N_A_3289_47#_c_1779_n 0.0096277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_3289_47#_c_1780_n 0.00367207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_3289_47#_c_1781_n 0.00682262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_3289_47#_c_1782_n 0.00723502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_3289_47#_c_1783_n 0.0434731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VPWR_c_1889_n 0.760753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_202_119#_c_2083_n 0.0024095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_202_119#_c_2084_n 0.00565537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_202_119#_c_2085_n 0.00279572f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_138 VNB N_A_202_119#_c_2086_n 0.00708087f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.55
cc_139 VNB N_A_202_119#_c_2087_n 0.00487337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_202_119#_c_2088_n 0.0138662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_Q_N_c_2231_n 0.0012299f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.275
cc_142 VNB N_Q_N_c_2232_n 0.00446691f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.885
cc_143 VNB N_Q_N_c_2233_n 0.00244613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2290_n 0.0138117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2291_n 0.042535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2292_n 0.0143756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2293_n 0.0318548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2294_n 0.0249838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2295_n 0.0158928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2296_n 0.0117815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2297_n 0.0190236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2298_n 0.0258886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2299_n 0.0177711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2300_n 0.0078123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2301_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2302_n 0.0469148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2303_n 0.0285324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2304_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2305_n 0.05269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2306_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2307_n 0.0560233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2308_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2309_n 0.0498314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2310_n 0.0375823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2311_n 0.0566772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2312_n 0.0590607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2313_n 0.0194324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2314_n 0.020631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2315_n 0.0188675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2316_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2317_n 0.00445561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2318_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2319_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2320_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2321_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2322_n 0.915222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_A_1670_93#_c_2481_n 0.00300559f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=2.2
cc_178 VNB N_A_2574_119#_c_2507_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=1.885
cc_179 VNB N_A_2574_119#_c_2508_n 0.00743815f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=2.725
cc_180 VNB N_A_2574_119#_c_2509_n 0.0079228f $X=-0.19 $Y=-0.245 $X2=0.42
+ $Y2=1.885
cc_181 VPB N_SCD_c_350_n 0.0025809f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.685
cc_182 VPB N_SCD_c_355_n 0.0195441f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.125
cc_183 VPB N_SCD_M1048_g 0.0226257f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.725
cc_184 VPB N_SCD_c_357_n 0.0254319f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_185 VPB N_SCD_c_358_n 0.0162564f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.2
cc_186 VPB N_SCD_c_353_n 0.0126687f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_187 VPB N_D_M1051_g 0.0440745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_D_c_389_n 0.0159846f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.725
cc_189 VPB D 0.00295819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_407_93#_c_439_n 0.0388306f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.725
cc_191 VPB N_A_407_93#_M1015_g 0.0437333f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_192 VPB N_A_407_93#_c_437_n 0.00966614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_407_93#_c_442_n 0.0102432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_407_93#_c_443_n 0.00171359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_407_93#_c_444_n 0.00469707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_407_93#_c_438_n 0.00343808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_SCE_c_504_n 0.00320899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_SCE_M1050_g 0.0384073f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.725
cc_199 VPB N_SCE_M1028_g 0.0308345f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_SCE_c_515_n 0.018044f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_201 VPB SCE 0.00260879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_CLK_N_M1025_g 0.0350059f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.885
cc_203 VPB N_CLK_N_c_579_n 0.0160906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB CLK_N 0.00195539f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_205 VPB N_A_840_95#_M1008_g 0.0457462f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.2
cc_206 VPB N_A_840_95#_c_631_n 0.067643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_840_95#_c_632_n 0.0128077f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_208 VPB N_A_840_95#_M1042_g 0.0326987f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_209 VPB N_A_840_95#_c_634_n 0.0158937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_840_95#_c_615_n 0.0292414f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_840_95#_c_616_n 6.74914e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_840_95#_c_637_n 0.0389698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_840_95#_c_618_n 0.0217055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_840_95#_c_639_n 0.00655786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_840_95#_c_640_n 0.00873071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_840_95#_c_641_n 0.00448393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_840_95#_c_642_n 0.00481627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_840_95#_c_643_n 0.0512358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_840_95#_c_627_n 0.00458909f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_840_95#_c_628_n 0.00700152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_1423_401#_M1018_g 0.0216519f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.275
cc_222 VPB N_A_1423_401#_M1017_g 0.0117162f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_223 VPB N_A_1423_401#_M1039_g 0.0242843f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_224 VPB N_A_1423_401#_c_834_n 0.00147176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1423_401#_c_843_n 0.00929405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_1423_401#_c_844_n 0.0138281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_1423_401#_c_845_n 0.00465681f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_1423_401#_c_836_n 0.00182751f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_1423_401#_c_837_n 0.0215349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_1423_401#_c_848_n 0.0634801f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_SET_B_M1043_g 0.0252397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_SET_B_c_965_n 0.0209982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_SET_B_c_966_n 0.0168474f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_234 VPB N_SET_B_c_967_n 0.0255792f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_235 VPB N_SET_B_c_959_n 0.00367426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_SET_B_c_962_n 0.00640607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_1273_137#_M1033_g 0.0170284f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_238 VPB N_A_1273_137#_c_1087_n 0.00443004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_1273_137#_c_1095_n 0.00461787f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.38
cc_240 VPB N_A_1273_137#_c_1096_n 0.015353f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.215
cc_241 VPB N_A_1273_137#_c_1097_n 0.00359115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_1273_137#_c_1098_n 0.0144494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1273_137#_c_1091_n 0.0106555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_1273_137#_c_1100_n 0.00346726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_1273_137#_c_1092_n 0.00587883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_978_67#_c_1206_n 0.0145514f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.885
cc_247 VPB N_A_978_67#_c_1207_n 0.0192593f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.125
cc_248 VPB N_A_978_67#_M1011_g 0.0069578f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.725
cc_249 VPB N_A_978_67#_c_1209_n 0.0362207f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_250 VPB N_A_978_67#_M1045_g 0.0445319f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_251 VPB N_A_978_67#_c_1211_n 0.340116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_978_67#_c_1212_n 0.0103267f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.38
cc_253 VPB N_A_978_67#_M1020_g 0.0105781f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.55
cc_254 VPB N_A_978_67#_c_1214_n 0.0268866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_978_67#_c_1215_n 0.00830324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_A_978_67#_c_1198_n 0.0167653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_978_67#_c_1217_n 0.004984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_978_67#_c_1202_n 0.00432795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_978_67#_c_1219_n 0.0147408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_978_67#_c_1204_n 0.00963969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_2415_137#_M1035_g 0.0292174f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.2
cc_262 VPB N_A_2415_137#_M1001_g 0.0213395f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_263 VPB N_A_2415_137#_M1024_g 0.0224184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_2415_137#_c_1337_n 0.00392557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_2415_137#_c_1353_n 0.0348193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_2415_137#_c_1354_n 0.013871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_2415_137#_c_1355_n 0.0184002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_2415_137#_c_1356_n 0.00799352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_2415_137#_c_1344_n 0.00448058f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_2415_137#_c_1358_n 0.0137396f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_2415_137#_c_1345_n 0.00137162f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_2415_137#_c_1360_n 0.00998514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_2415_137#_c_1361_n 0.0328285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_A_2415_137#_c_1362_n 0.0024362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_2415_137#_c_1347_n 0.0182928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_2211_428#_M1000_g 0.0356112f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_277 VPB N_A_2211_428#_c_1542_n 0.00370572f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.38
cc_278 VPB N_A_2211_428#_c_1537_n 0.00426347f $X=-0.19 $Y=1.655 $X2=0.42
+ $Y2=1.215
cc_279 VPB N_A_2211_428#_c_1539_n 0.00119081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_A_2211_428#_c_1540_n 0.0169045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_A_1840_21#_M1005_g 0.027016f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_282 VPB N_A_1840_21#_M1026_g 0.0236185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_A_1840_21#_c_1634_n 0.0464258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_1840_21#_c_1639_n 0.00410537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_A_1840_21#_c_1640_n 0.00722656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_RESET_B_c_1735_n 0.00653147f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.415
cc_287 VPB N_RESET_B_M1040_g 0.0236418f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.215
cc_288 VPB N_RESET_B_c_1737_n 0.00310576f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.885
cc_289 VPB N_A_3289_47#_M1002_g 0.0230937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_290 VPB N_A_3289_47#_M1034_g 0.0265102f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_291 VPB N_A_3289_47#_c_1780_n 0.0135419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB N_A_56_481#_c_1839_n 0.0338707f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.275
cc_293 VPB N_A_56_481#_c_1840_n 0.0239417f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.725
cc_294 VPB N_A_56_481#_c_1841_n 0.00843023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_295 VPB N_A_56_481#_c_1842_n 0.00154399f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.2
cc_296 VPB N_A_56_481#_c_1843_n 0.00732312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_A_56_481#_c_1844_n 0.00134745f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.2
cc_298 VPB N_A_56_481#_c_1845_n 0.00896469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_1890_n 0.00415775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_1891_n 0.0265465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_1892_n 0.0236959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_1893_n 0.00639252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_1894_n 0.018998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_1895_n 0.0252893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_1896_n 0.00808769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_1897_n 0.016554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_1898_n 0.0161915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_1899_n 0.0309629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_1900_n 0.022221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_1901_n 0.0106521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_1902_n 0.062339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_1903_n 0.0236202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_1904_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_1905_n 0.0397935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_1906_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_1907_n 0.0188705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_1908_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_1909_n 0.0667219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_1910_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_1911_n 0.0327958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_321 VPB N_VPWR_c_1912_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_1913_n 0.0354234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_1914_n 0.0770723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_1915_n 0.0276855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_1916_n 0.02253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_1917_n 0.0166909f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_1918_n 0.0221759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_1919_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_1920_n 0.00455177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_1921_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_1922_n 0.00510817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_1923_n 0.00510817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_1924_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_1925_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_1889_n 0.182633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_336 VPB N_A_202_119#_c_2089_n 0.00463885f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.38
cc_337 VPB N_A_202_119#_c_2086_n 0.00515096f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.55
cc_338 VPB N_A_202_119#_c_2091_n 0.0564993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_339 VPB N_A_202_119#_c_2092_n 0.00697344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_340 VPB N_A_202_119#_c_2093_n 0.0256866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_341 VPB N_A_202_119#_c_2094_n 0.00326464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_342 VPB N_A_202_119#_c_2087_n 0.00786784f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_343 VPB N_A_202_119#_c_2096_n 0.013071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_344 VPB N_A_202_119#_c_2097_n 0.0091443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_345 VPB N_A_202_119#_c_2098_n 0.00945764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_346 VPB Q_N 0.00158315f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.2
cc_347 VPB N_Q_N_c_2233_n 7.87357e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_348 N_SCD_M1013_g N_SCE_M1036_g 0.0187336f $X=0.545 $Y=0.805 $X2=0 $Y2=0
cc_349 N_SCD_c_350_n N_SCE_c_504_n 0.0187336f $X=0.42 $Y=1.685 $X2=0 $Y2=0
cc_350 N_SCD_c_355_n N_SCE_M1050_g 0.0072044f $X=0.545 $Y=2.125 $X2=0 $Y2=0
cc_351 N_SCD_c_358_n N_SCE_M1050_g 0.0248986f $X=0.64 $Y=2.2 $X2=0 $Y2=0
cc_352 N_SCD_c_357_n N_SCE_c_515_n 0.0187336f $X=0.42 $Y=1.885 $X2=0 $Y2=0
cc_353 N_SCD_c_352_n SCE 0.00250463f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_354 N_SCD_c_353_n SCE 0.0295869f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_355 N_SCD_c_352_n N_SCE_c_511_n 0.0187336f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_356 N_SCD_c_353_n N_SCE_c_511_n 0.00228677f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_357 N_SCD_M1048_g N_A_56_481#_c_1839_n 0.0126781f $X=0.64 $Y=2.725 $X2=0
+ $Y2=0
cc_358 N_SCD_c_358_n N_A_56_481#_c_1839_n 0.00422291f $X=0.64 $Y=2.2 $X2=0 $Y2=0
cc_359 N_SCD_c_355_n N_A_56_481#_c_1840_n 0.00240509f $X=0.545 $Y=2.125 $X2=0
+ $Y2=0
cc_360 N_SCD_c_358_n N_A_56_481#_c_1840_n 0.00976765f $X=0.64 $Y=2.2 $X2=0 $Y2=0
cc_361 N_SCD_c_355_n N_A_56_481#_c_1841_n 0.00503383f $X=0.545 $Y=2.125 $X2=0
+ $Y2=0
cc_362 N_SCD_c_357_n N_A_56_481#_c_1841_n 0.00560551f $X=0.42 $Y=1.885 $X2=0
+ $Y2=0
cc_363 N_SCD_c_358_n N_A_56_481#_c_1841_n 0.00328627f $X=0.64 $Y=2.2 $X2=0 $Y2=0
cc_364 N_SCD_c_353_n N_A_56_481#_c_1841_n 0.0242556f $X=0.385 $Y=1.38 $X2=0
+ $Y2=0
cc_365 N_SCD_M1048_g N_VPWR_c_1890_n 0.00606558f $X=0.64 $Y=2.725 $X2=0 $Y2=0
cc_366 N_SCD_M1048_g N_VPWR_c_1903_n 0.00502664f $X=0.64 $Y=2.725 $X2=0 $Y2=0
cc_367 N_SCD_M1048_g N_VPWR_c_1889_n 0.010292f $X=0.64 $Y=2.725 $X2=0 $Y2=0
cc_368 N_SCD_M1013_g N_A_202_119#_c_2083_n 0.00114555f $X=0.545 $Y=0.805 $X2=0
+ $Y2=0
cc_369 N_SCD_M1013_g N_A_202_119#_c_2085_n 4.65148e-19 $X=0.545 $Y=0.805 $X2=0
+ $Y2=0
cc_370 N_SCD_M1013_g N_VGND_c_2291_n 0.0140065f $X=0.545 $Y=0.805 $X2=0 $Y2=0
cc_371 N_SCD_c_352_n N_VGND_c_2291_n 0.00667323f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_372 N_SCD_c_353_n N_VGND_c_2291_n 0.0279841f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_373 N_SCD_M1013_g N_VGND_c_2309_n 0.0035863f $X=0.545 $Y=0.805 $X2=0 $Y2=0
cc_374 N_SCD_M1013_g N_VGND_c_2322_n 0.00401353f $X=0.545 $Y=0.805 $X2=0 $Y2=0
cc_375 N_D_c_387_n N_A_407_93#_M1004_g 0.0166356f $X=1.63 $Y=1.125 $X2=0 $Y2=0
cc_376 D N_A_407_93#_M1004_g 0.00129718f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_377 N_D_c_391_n N_A_407_93#_M1004_g 0.0055196f $X=1.63 $Y=1.29 $X2=0 $Y2=0
cc_378 N_D_M1051_g N_A_407_93#_c_439_n 0.0302494f $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_379 N_D_c_389_n N_A_407_93#_c_439_n 0.00329761f $X=1.63 $Y=1.795 $X2=0 $Y2=0
cc_380 N_D_c_388_n N_A_407_93#_c_435_n 0.0055196f $X=1.63 $Y=1.63 $X2=0 $Y2=0
cc_381 N_D_c_388_n N_A_407_93#_c_437_n 0.00329761f $X=1.63 $Y=1.63 $X2=0 $Y2=0
cc_382 N_D_c_387_n N_SCE_M1036_g 0.0098253f $X=1.63 $Y=1.125 $X2=0 $Y2=0
cc_383 D N_SCE_M1036_g 5.45014e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_384 N_D_c_388_n N_SCE_c_504_n 0.025404f $X=1.63 $Y=1.63 $X2=0 $Y2=0
cc_385 N_D_c_387_n N_SCE_c_505_n 0.00895556f $X=1.63 $Y=1.125 $X2=0 $Y2=0
cc_386 N_D_M1051_g N_SCE_M1050_g 0.025404f $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_387 N_D_c_389_n N_SCE_c_515_n 0.025404f $X=1.63 $Y=1.795 $X2=0 $Y2=0
cc_388 D SCE 0.0445848f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_389 N_D_c_391_n SCE 0.00487283f $X=1.63 $Y=1.29 $X2=0 $Y2=0
cc_390 D N_SCE_c_511_n 5.88162e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_391 N_D_c_391_n N_SCE_c_511_n 0.025404f $X=1.63 $Y=1.29 $X2=0 $Y2=0
cc_392 N_D_M1051_g N_A_56_481#_c_1840_n 0.00357016f $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_393 N_D_M1051_g N_A_56_481#_c_1842_n 0.0120522f $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_394 N_D_M1051_g N_A_56_481#_c_1843_n 0.0124379f $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_395 N_D_M1051_g N_A_56_481#_c_1844_n 0.00127595f $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_396 N_D_M1051_g N_A_56_481#_c_1845_n 8.88533e-19 $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_397 N_D_M1051_g N_VPWR_c_1890_n 0.00135656f $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_398 N_D_M1051_g N_VPWR_c_1905_n 0.0032772f $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_399 N_D_M1051_g N_VPWR_c_1889_n 0.00504385f $X=1.54 $Y=2.725 $X2=0 $Y2=0
cc_400 N_D_c_387_n N_A_202_119#_c_2083_n 0.00429145f $X=1.63 $Y=1.125 $X2=0
+ $Y2=0
cc_401 D N_A_202_119#_c_2083_n 0.0166259f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_402 N_D_c_387_n N_A_202_119#_c_2084_n 0.0108591f $X=1.63 $Y=1.125 $X2=0 $Y2=0
cc_403 D N_A_202_119#_c_2084_n 0.0175193f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_404 N_D_c_391_n N_A_202_119#_c_2084_n 5.58334e-19 $X=1.63 $Y=1.29 $X2=0 $Y2=0
cc_405 N_D_M1051_g N_A_202_119#_c_2089_n 0.00386482f $X=1.54 $Y=2.725 $X2=0
+ $Y2=0
cc_406 N_D_M1051_g N_A_202_119#_c_2086_n 0.00399208f $X=1.54 $Y=2.725 $X2=0
+ $Y2=0
cc_407 N_D_c_387_n N_A_202_119#_c_2086_n 0.00224486f $X=1.63 $Y=1.125 $X2=0
+ $Y2=0
cc_408 D N_A_202_119#_c_2086_n 0.0710291f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_409 N_D_c_391_n N_A_202_119#_c_2086_n 0.00665717f $X=1.63 $Y=1.29 $X2=0 $Y2=0
cc_410 N_D_M1051_g N_A_202_119#_c_2096_n 0.00248814f $X=1.54 $Y=2.725 $X2=0
+ $Y2=0
cc_411 N_D_c_389_n N_A_202_119#_c_2096_n 0.00107601f $X=1.63 $Y=1.795 $X2=0
+ $Y2=0
cc_412 D N_A_202_119#_c_2096_n 0.00990081f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_413 D A_323_119# 0.00306091f $X=1.595 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_414 N_A_407_93#_M1004_g N_SCE_c_505_n 0.00934409f $X=2.11 $Y=0.805 $X2=0
+ $Y2=0
cc_415 N_A_407_93#_M1004_g N_SCE_M1016_g 0.00891539f $X=2.11 $Y=0.805 $X2=0
+ $Y2=0
cc_416 N_A_407_93#_c_438_n N_SCE_M1016_g 0.0130137f $X=3.11 $Y=0.805 $X2=0 $Y2=0
cc_417 N_A_407_93#_c_439_n N_SCE_M1028_g 0.00411971f $X=2.11 $Y=2.005 $X2=0
+ $Y2=0
cc_418 N_A_407_93#_c_435_n N_SCE_M1028_g 0.0165637f $X=2.415 $Y=1.335 $X2=0
+ $Y2=0
cc_419 N_A_407_93#_c_436_n N_SCE_M1028_g 3.29189e-19 $X=2.415 $Y=1.35 $X2=0
+ $Y2=0
cc_420 N_A_407_93#_c_444_n N_SCE_M1028_g 0.0126698f $X=3.195 $Y=1.515 $X2=0
+ $Y2=0
cc_421 N_A_407_93#_c_438_n N_SCE_M1028_g 0.0112913f $X=3.11 $Y=0.805 $X2=0 $Y2=0
cc_422 N_A_407_93#_c_435_n N_SCE_c_509_n 0.00303664f $X=2.415 $Y=1.335 $X2=0
+ $Y2=0
cc_423 N_A_407_93#_c_436_n N_SCE_c_509_n 2.17594e-19 $X=2.415 $Y=1.35 $X2=0
+ $Y2=0
cc_424 N_A_407_93#_c_442_n N_SCE_c_509_n 0.00495325f $X=2.945 $Y=1.685 $X2=0
+ $Y2=0
cc_425 N_A_407_93#_c_438_n N_SCE_c_509_n 0.015419f $X=3.11 $Y=0.805 $X2=0 $Y2=0
cc_426 N_A_407_93#_c_438_n N_CLK_N_M1049_g 0.00540093f $X=3.11 $Y=0.805 $X2=0
+ $Y2=0
cc_427 N_A_407_93#_c_444_n N_CLK_N_M1025_g 0.00195235f $X=3.195 $Y=1.515 $X2=0
+ $Y2=0
cc_428 N_A_407_93#_c_444_n N_CLK_N_c_578_n 0.00523611f $X=3.195 $Y=1.515 $X2=0
+ $Y2=0
cc_429 N_A_407_93#_c_444_n CLK_N 0.0112768f $X=3.195 $Y=1.515 $X2=0 $Y2=0
cc_430 N_A_407_93#_c_438_n CLK_N 0.0167329f $X=3.11 $Y=0.805 $X2=0 $Y2=0
cc_431 N_A_407_93#_c_438_n N_CLK_N_c_581_n 0.00785852f $X=3.11 $Y=0.805 $X2=0
+ $Y2=0
cc_432 N_A_407_93#_M1015_g N_A_56_481#_c_1842_n 8.96477e-19 $X=2.11 $Y=2.725
+ $X2=0 $Y2=0
cc_433 N_A_407_93#_M1015_g N_A_56_481#_c_1843_n 0.0119851f $X=2.11 $Y=2.725
+ $X2=0 $Y2=0
cc_434 N_A_407_93#_M1015_g N_A_56_481#_c_1845_n 0.00787022f $X=2.11 $Y=2.725
+ $X2=0 $Y2=0
cc_435 N_A_407_93#_c_442_n N_VPWR_M1028_s 0.00303482f $X=2.945 $Y=1.685 $X2=0
+ $Y2=0
cc_436 N_A_407_93#_M1015_g N_VPWR_c_1891_n 0.00299758f $X=2.11 $Y=2.725 $X2=0
+ $Y2=0
cc_437 N_A_407_93#_M1015_g N_VPWR_c_1905_n 0.00327695f $X=2.11 $Y=2.725 $X2=0
+ $Y2=0
cc_438 N_A_407_93#_M1015_g N_VPWR_c_1889_n 0.00599582f $X=2.11 $Y=2.725 $X2=0
+ $Y2=0
cc_439 N_A_407_93#_M1004_g N_A_202_119#_c_2084_n 0.0054637f $X=2.11 $Y=0.805
+ $X2=0 $Y2=0
cc_440 N_A_407_93#_M1015_g N_A_202_119#_c_2089_n 0.00719918f $X=2.11 $Y=2.725
+ $X2=0 $Y2=0
cc_441 N_A_407_93#_M1004_g N_A_202_119#_c_2086_n 0.0152679f $X=2.11 $Y=0.805
+ $X2=0 $Y2=0
cc_442 N_A_407_93#_c_439_n N_A_202_119#_c_2086_n 0.0106442f $X=2.11 $Y=2.005
+ $X2=0 $Y2=0
cc_443 N_A_407_93#_M1015_g N_A_202_119#_c_2086_n 0.00153923f $X=2.11 $Y=2.725
+ $X2=0 $Y2=0
cc_444 N_A_407_93#_c_435_n N_A_202_119#_c_2086_n 0.00622804f $X=2.415 $Y=1.335
+ $X2=0 $Y2=0
cc_445 N_A_407_93#_c_436_n N_A_202_119#_c_2086_n 0.0226636f $X=2.415 $Y=1.35
+ $X2=0 $Y2=0
cc_446 N_A_407_93#_c_437_n N_A_202_119#_c_2086_n 0.00323037f $X=2.415 $Y=1.35
+ $X2=0 $Y2=0
cc_447 N_A_407_93#_c_443_n N_A_202_119#_c_2086_n 0.0259744f $X=2.58 $Y=1.685
+ $X2=0 $Y2=0
cc_448 N_A_407_93#_M1028_d N_A_202_119#_c_2091_n 0.00301164f $X=3.14 $Y=1.535
+ $X2=0 $Y2=0
cc_449 N_A_407_93#_c_439_n N_A_202_119#_c_2091_n 0.0098017f $X=2.11 $Y=2.005
+ $X2=0 $Y2=0
cc_450 N_A_407_93#_M1015_g N_A_202_119#_c_2091_n 0.00717659f $X=2.11 $Y=2.725
+ $X2=0 $Y2=0
cc_451 N_A_407_93#_c_442_n N_A_202_119#_c_2091_n 0.0263425f $X=2.945 $Y=1.685
+ $X2=0 $Y2=0
cc_452 N_A_407_93#_c_443_n N_A_202_119#_c_2091_n 0.0194875f $X=2.58 $Y=1.685
+ $X2=0 $Y2=0
cc_453 N_A_407_93#_c_444_n N_A_202_119#_c_2091_n 0.0302691f $X=3.195 $Y=1.515
+ $X2=0 $Y2=0
cc_454 N_A_407_93#_M1015_g N_A_202_119#_c_2096_n 0.00987918f $X=2.11 $Y=2.725
+ $X2=0 $Y2=0
cc_455 N_A_407_93#_M1004_g N_VGND_c_2292_n 0.00533347f $X=2.11 $Y=0.805 $X2=0
+ $Y2=0
cc_456 N_A_407_93#_c_435_n N_VGND_c_2292_n 0.00196592f $X=2.415 $Y=1.335 $X2=0
+ $Y2=0
cc_457 N_A_407_93#_c_436_n N_VGND_c_2292_n 0.0211246f $X=2.415 $Y=1.35 $X2=0
+ $Y2=0
cc_458 N_A_407_93#_c_442_n N_VGND_c_2292_n 0.00289626f $X=2.945 $Y=1.685 $X2=0
+ $Y2=0
cc_459 N_A_407_93#_c_438_n N_VGND_c_2292_n 0.0228902f $X=3.11 $Y=0.805 $X2=0
+ $Y2=0
cc_460 N_A_407_93#_c_438_n N_VGND_c_2293_n 0.0244052f $X=3.11 $Y=0.805 $X2=0
+ $Y2=0
cc_461 N_A_407_93#_c_438_n N_VGND_c_2303_n 0.0114264f $X=3.11 $Y=0.805 $X2=0
+ $Y2=0
cc_462 N_A_407_93#_M1004_g N_VGND_c_2322_n 2.50464e-19 $X=2.11 $Y=0.805 $X2=0
+ $Y2=0
cc_463 N_A_407_93#_c_438_n N_VGND_c_2322_n 0.0156679f $X=3.11 $Y=0.805 $X2=0
+ $Y2=0
cc_464 N_SCE_M1050_g N_A_56_481#_c_1839_n 0.00112038f $X=1.15 $Y=2.725 $X2=0
+ $Y2=0
cc_465 N_SCE_M1050_g N_A_56_481#_c_1840_n 0.0146379f $X=1.15 $Y=2.725 $X2=0
+ $Y2=0
cc_466 N_SCE_c_515_n N_A_56_481#_c_1840_n 0.00612316f $X=1.042 $Y=1.885 $X2=0
+ $Y2=0
cc_467 SCE N_A_56_481#_c_1840_n 0.0318981f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_468 N_SCE_M1050_g N_A_56_481#_c_1842_n 0.00724504f $X=1.15 $Y=2.725 $X2=0
+ $Y2=0
cc_469 N_SCE_M1050_g N_A_56_481#_c_1844_n 0.00132979f $X=1.15 $Y=2.725 $X2=0
+ $Y2=0
cc_470 N_SCE_M1050_g N_VPWR_c_1890_n 0.0146125f $X=1.15 $Y=2.725 $X2=0 $Y2=0
cc_471 N_SCE_M1028_g N_VPWR_c_1891_n 0.00175888f $X=3.065 $Y=1.855 $X2=0 $Y2=0
cc_472 N_SCE_M1050_g N_VPWR_c_1905_n 0.00445056f $X=1.15 $Y=2.725 $X2=0 $Y2=0
cc_473 N_SCE_M1050_g N_VPWR_c_1889_n 0.00804604f $X=1.15 $Y=2.725 $X2=0 $Y2=0
cc_474 N_SCE_M1036_g N_A_202_119#_c_2083_n 0.00754356f $X=0.935 $Y=0.805 $X2=0
+ $Y2=0
cc_475 SCE N_A_202_119#_c_2083_n 0.0277811f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_476 N_SCE_c_511_n N_A_202_119#_c_2083_n 0.00576357f $X=1.06 $Y=1.38 $X2=0
+ $Y2=0
cc_477 N_SCE_c_505_n N_A_202_119#_c_2084_n 0.0136254f $X=2.82 $Y=0.18 $X2=0
+ $Y2=0
cc_478 N_SCE_M1036_g N_A_202_119#_c_2085_n 0.00579034f $X=0.935 $Y=0.805 $X2=0
+ $Y2=0
cc_479 N_SCE_c_505_n N_A_202_119#_c_2085_n 0.00468683f $X=2.82 $Y=0.18 $X2=0
+ $Y2=0
cc_480 N_SCE_M1016_g N_A_202_119#_c_2086_n 9.4274e-19 $X=2.895 $Y=0.805 $X2=0
+ $Y2=0
cc_481 SCE N_A_202_119#_c_2086_n 0.00276129f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_482 N_SCE_M1028_g N_A_202_119#_c_2091_n 0.0165516f $X=3.065 $Y=1.855 $X2=0
+ $Y2=0
cc_483 N_SCE_M1036_g N_VGND_c_2291_n 0.00161317f $X=0.935 $Y=0.805 $X2=0 $Y2=0
cc_484 N_SCE_c_506_n N_VGND_c_2291_n 0.0102374f $X=1.01 $Y=0.18 $X2=0 $Y2=0
cc_485 N_SCE_c_505_n N_VGND_c_2292_n 0.0258022f $X=2.82 $Y=0.18 $X2=0 $Y2=0
cc_486 N_SCE_M1016_g N_VGND_c_2292_n 0.0154689f $X=2.895 $Y=0.805 $X2=0 $Y2=0
cc_487 N_SCE_c_505_n N_VGND_c_2293_n 0.00889775f $X=2.82 $Y=0.18 $X2=0 $Y2=0
cc_488 N_SCE_M1016_g N_VGND_c_2293_n 4.9575e-19 $X=2.895 $Y=0.805 $X2=0 $Y2=0
cc_489 N_SCE_c_505_n N_VGND_c_2303_n 0.0117032f $X=2.82 $Y=0.18 $X2=0 $Y2=0
cc_490 N_SCE_c_506_n N_VGND_c_2309_n 0.0379972f $X=1.01 $Y=0.18 $X2=0 $Y2=0
cc_491 N_SCE_c_505_n N_VGND_c_2322_n 0.0568351f $X=2.82 $Y=0.18 $X2=0 $Y2=0
cc_492 N_SCE_c_506_n N_VGND_c_2322_n 0.0107139f $X=1.01 $Y=0.18 $X2=0 $Y2=0
cc_493 N_CLK_N_M1049_g N_A_840_95#_c_615_n 0.0354317f $X=4.125 $Y=0.685 $X2=0
+ $Y2=0
cc_494 CLK_N N_A_840_95#_c_615_n 6.97921e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_495 N_CLK_N_M1049_g N_A_840_95#_c_617_n 0.0128402f $X=4.125 $Y=0.685 $X2=0
+ $Y2=0
cc_496 CLK_N N_A_840_95#_c_617_n 0.00609632f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_497 N_CLK_N_M1025_g N_A_840_95#_c_618_n 0.00451904f $X=4.125 $Y=2.375 $X2=0
+ $Y2=0
cc_498 CLK_N N_A_840_95#_c_618_n 0.0387551f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_499 N_CLK_N_c_581_n N_A_840_95#_c_618_n 0.0143071f $X=4.035 $Y=1.275 $X2=0
+ $Y2=0
cc_500 N_CLK_N_M1049_g N_A_978_67#_c_1205_n 0.00302314f $X=4.125 $Y=0.685 $X2=0
+ $Y2=0
cc_501 N_CLK_N_M1025_g N_VPWR_c_1892_n 0.00870221f $X=4.125 $Y=2.375 $X2=0 $Y2=0
cc_502 N_CLK_N_M1025_g N_VPWR_c_1913_n 0.00114147f $X=4.125 $Y=2.375 $X2=0 $Y2=0
cc_503 N_CLK_N_M1025_g N_VPWR_c_1889_n 7.94274e-19 $X=4.125 $Y=2.375 $X2=0 $Y2=0
cc_504 N_CLK_N_M1025_g N_A_202_119#_c_2091_n 0.0126218f $X=4.125 $Y=2.375 $X2=0
+ $Y2=0
cc_505 N_CLK_N_c_579_n N_A_202_119#_c_2091_n 0.00114681f $X=4.035 $Y=1.78 $X2=0
+ $Y2=0
cc_506 CLK_N N_A_202_119#_c_2091_n 0.0194334f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_507 N_CLK_N_M1025_g N_A_202_119#_c_2092_n 0.0279702f $X=4.125 $Y=2.375 $X2=0
+ $Y2=0
cc_508 N_CLK_N_M1049_g N_VGND_c_2293_n 0.0135661f $X=4.125 $Y=0.685 $X2=0 $Y2=0
cc_509 CLK_N N_VGND_c_2293_n 0.00987215f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_510 N_CLK_N_c_581_n N_VGND_c_2293_n 9.46932e-19 $X=4.035 $Y=1.275 $X2=0 $Y2=0
cc_511 N_CLK_N_M1049_g N_VGND_c_2310_n 0.00481548f $X=4.125 $Y=0.685 $X2=0 $Y2=0
cc_512 N_CLK_N_M1049_g N_VGND_c_2322_n 0.00512916f $X=4.125 $Y=0.685 $X2=0 $Y2=0
cc_513 N_A_840_95#_M1044_g N_A_1423_401#_M1017_g 0.0156934f $X=6.72 $Y=0.895
+ $X2=0 $Y2=0
cc_514 N_A_840_95#_c_619_n N_A_1423_401#_M1017_g 0.00555586f $X=6.855 $Y=1.38
+ $X2=0 $Y2=0
cc_515 N_A_840_95#_c_620_n N_A_1423_401#_M1017_g 0.0185604f $X=6.855 $Y=1.38
+ $X2=0 $Y2=0
cc_516 N_A_840_95#_c_656_p N_A_1423_401#_M1017_g 0.0160804f $X=7.975 $Y=0.915
+ $X2=0 $Y2=0
cc_517 N_A_840_95#_c_621_n N_A_1423_401#_M1017_g 0.00417932f $X=8.06 $Y=0.83
+ $X2=0 $Y2=0
cc_518 N_A_840_95#_c_624_n N_A_1423_401#_M1046_g 0.00549154f $X=9.94 $Y=1.095
+ $X2=0 $Y2=0
cc_519 N_A_840_95#_c_625_n N_A_1423_401#_M1046_g 0.0157659f $X=10.68 $Y=1.18
+ $X2=0 $Y2=0
cc_520 N_A_840_95#_c_627_n N_A_1423_401#_M1046_g 0.0185365f $X=10.9 $Y=1.18
+ $X2=0 $Y2=0
cc_521 N_A_840_95#_c_628_n N_A_1423_401#_M1046_g 0.0206552f $X=10.955 $Y=1.51
+ $X2=0 $Y2=0
cc_522 N_A_840_95#_c_629_n N_A_1423_401#_M1046_g 0.0314322f $X=10.955 $Y=1.345
+ $X2=0 $Y2=0
cc_523 N_A_840_95#_c_624_n N_A_1423_401#_c_832_n 0.00130895f $X=9.94 $Y=1.095
+ $X2=0 $Y2=0
cc_524 N_A_840_95#_c_626_n N_A_1423_401#_c_832_n 0.00482664f $X=10.025 $Y=1.18
+ $X2=0 $Y2=0
cc_525 N_A_840_95#_c_626_n N_A_1423_401#_c_833_n 7.13716e-19 $X=10.025 $Y=1.18
+ $X2=0 $Y2=0
cc_526 N_A_840_95#_c_627_n N_A_1423_401#_c_836_n 0.020617f $X=10.9 $Y=1.18 $X2=0
+ $Y2=0
cc_527 N_A_840_95#_c_628_n N_A_1423_401#_c_836_n 2.03767e-19 $X=10.955 $Y=1.51
+ $X2=0 $Y2=0
cc_528 N_A_840_95#_c_625_n N_A_1423_401#_c_837_n 0.00594544f $X=10.68 $Y=1.18
+ $X2=0 $Y2=0
cc_529 N_A_840_95#_c_639_n N_A_1423_401#_c_837_n 0.0182409f $X=10.765 $Y=2.895
+ $X2=0 $Y2=0
cc_530 N_A_840_95#_c_625_n N_A_1423_401#_c_838_n 0.0282853f $X=10.68 $Y=1.18
+ $X2=0 $Y2=0
cc_531 N_A_840_95#_c_626_n N_A_1423_401#_c_838_n 0.0106774f $X=10.025 $Y=1.18
+ $X2=0 $Y2=0
cc_532 N_A_840_95#_c_621_n N_SET_B_c_954_n 0.00811663f $X=8.06 $Y=0.83 $X2=-0.19
+ $Y2=-0.245
cc_533 N_A_840_95#_c_622_n N_SET_B_c_954_n 0.0127235f $X=9.855 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_534 N_A_840_95#_c_625_n N_SET_B_c_956_n 0.0301202f $X=10.68 $Y=1.18 $X2=0
+ $Y2=0
cc_535 N_A_840_95#_c_626_n N_SET_B_c_956_n 0.0116448f $X=10.025 $Y=1.18 $X2=0
+ $Y2=0
cc_536 N_A_840_95#_c_642_n N_SET_B_c_956_n 0.0128513f $X=11.855 $Y=1.865 $X2=0
+ $Y2=0
cc_537 N_A_840_95#_c_627_n N_SET_B_c_956_n 0.0483284f $X=10.9 $Y=1.18 $X2=0
+ $Y2=0
cc_538 N_A_840_95#_c_642_n N_SET_B_c_959_n 0.0024876f $X=11.855 $Y=1.865 $X2=0
+ $Y2=0
cc_539 N_A_840_95#_c_656_p N_SET_B_c_960_n 0.00143579f $X=7.975 $Y=0.915 $X2=0
+ $Y2=0
cc_540 N_A_840_95#_c_622_n N_A_1273_137#_M1029_g 0.00850531f $X=9.855 $Y=0.35
+ $X2=0 $Y2=0
cc_541 N_A_840_95#_c_612_n N_A_1273_137#_c_1087_n 0.00255267f $X=6.645 $Y=0.185
+ $X2=0 $Y2=0
cc_542 N_A_840_95#_M1044_g N_A_1273_137#_c_1087_n 0.00403954f $X=6.72 $Y=0.895
+ $X2=0 $Y2=0
cc_543 N_A_840_95#_c_619_n N_A_1273_137#_c_1087_n 0.0335198f $X=6.855 $Y=1.38
+ $X2=0 $Y2=0
cc_544 N_A_840_95#_M1042_g N_A_1273_137#_c_1095_n 0.00300307f $X=6.29 $Y=2.525
+ $X2=0 $Y2=0
cc_545 N_A_840_95#_c_619_n N_A_1273_137#_c_1096_n 0.00545723f $X=6.855 $Y=1.38
+ $X2=0 $Y2=0
cc_546 N_A_840_95#_c_620_n N_A_1273_137#_c_1096_n 0.00250947f $X=6.855 $Y=1.38
+ $X2=0 $Y2=0
cc_547 N_A_840_95#_c_656_p N_A_1273_137#_c_1088_n 0.0174843f $X=7.975 $Y=0.915
+ $X2=0 $Y2=0
cc_548 N_A_840_95#_c_619_n N_A_1273_137#_c_1089_n 0.00544029f $X=6.855 $Y=1.38
+ $X2=0 $Y2=0
cc_549 N_A_840_95#_c_620_n N_A_1273_137#_c_1089_n 5.41887e-19 $X=6.855 $Y=1.38
+ $X2=0 $Y2=0
cc_550 N_A_840_95#_c_656_p N_A_1273_137#_c_1089_n 0.00556785f $X=7.975 $Y=0.915
+ $X2=0 $Y2=0
cc_551 N_A_840_95#_M1042_g N_A_1273_137#_c_1100_n 5.58607e-19 $X=6.29 $Y=2.525
+ $X2=0 $Y2=0
cc_552 N_A_840_95#_c_656_p N_A_1273_137#_c_1092_n 0.00651005f $X=7.975 $Y=0.915
+ $X2=0 $Y2=0
cc_553 N_A_840_95#_M1008_g N_A_978_67#_c_1207_n 0.0194911f $X=5.31 $Y=2.665
+ $X2=0 $Y2=0
cc_554 N_A_840_95#_c_612_n N_A_978_67#_M1011_g 0.00720713f $X=6.645 $Y=0.185
+ $X2=0 $Y2=0
cc_555 N_A_840_95#_M1044_g N_A_978_67#_M1011_g 0.0235545f $X=6.72 $Y=0.895 $X2=0
+ $Y2=0
cc_556 N_A_840_95#_c_619_n N_A_978_67#_c_1209_n 5.11372e-19 $X=6.855 $Y=1.38
+ $X2=0 $Y2=0
cc_557 N_A_840_95#_c_620_n N_A_978_67#_c_1209_n 0.0133875f $X=6.855 $Y=1.38
+ $X2=0 $Y2=0
cc_558 N_A_840_95#_M1042_g N_A_978_67#_M1045_g 0.0141284f $X=6.29 $Y=2.525 $X2=0
+ $Y2=0
cc_559 N_A_840_95#_c_634_n N_A_978_67#_c_1211_n 0.0100806f $X=11.49 $Y=2.455
+ $X2=0 $Y2=0
cc_560 N_A_840_95#_c_641_n N_A_978_67#_c_1211_n 0.00332103f $X=10.85 $Y=2.98
+ $X2=0 $Y2=0
cc_561 N_A_840_95#_c_631_n N_A_978_67#_c_1212_n 0.0141284f $X=6.215 $Y=3.135
+ $X2=0 $Y2=0
cc_562 N_A_840_95#_c_637_n N_A_978_67#_M1020_g 0.0100806f $X=11.855 $Y=2.305
+ $X2=0 $Y2=0
cc_563 N_A_840_95#_c_640_n N_A_978_67#_M1020_g 0.0151989f $X=11.69 $Y=2.98 $X2=0
+ $Y2=0
cc_564 N_A_840_95#_c_643_n N_A_978_67#_M1020_g 0.00228806f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_565 N_A_840_95#_c_637_n N_A_978_67#_c_1214_n 0.00380864f $X=11.855 $Y=2.305
+ $X2=0 $Y2=0
cc_566 N_A_840_95#_c_639_n N_A_978_67#_c_1215_n 0.00676641f $X=10.765 $Y=2.895
+ $X2=0 $Y2=0
cc_567 N_A_840_95#_c_627_n N_A_978_67#_c_1215_n 0.00129252f $X=10.9 $Y=1.18
+ $X2=0 $Y2=0
cc_568 N_A_840_95#_c_628_n N_A_978_67#_c_1215_n 0.0117932f $X=10.955 $Y=1.51
+ $X2=0 $Y2=0
cc_569 N_A_840_95#_c_639_n N_A_978_67#_c_1198_n 0.00128999f $X=10.765 $Y=2.895
+ $X2=0 $Y2=0
cc_570 N_A_840_95#_c_642_n N_A_978_67#_c_1198_n 0.00123584f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_571 N_A_840_95#_c_643_n N_A_978_67#_c_1198_n 0.0219192f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_572 N_A_840_95#_c_642_n N_A_978_67#_c_1199_n 0.00108175f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_573 N_A_840_95#_c_643_n N_A_978_67#_c_1199_n 0.00825636f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_574 N_A_840_95#_c_627_n N_A_978_67#_c_1200_n 4.92054e-19 $X=10.9 $Y=1.18
+ $X2=0 $Y2=0
cc_575 N_A_840_95#_c_628_n N_A_978_67#_c_1200_n 0.0206946f $X=10.955 $Y=1.51
+ $X2=0 $Y2=0
cc_576 N_A_840_95#_c_629_n N_A_978_67#_c_1200_n 0.0018943f $X=10.955 $Y=1.345
+ $X2=0 $Y2=0
cc_577 N_A_840_95#_c_629_n N_A_978_67#_c_1201_n 0.00782077f $X=10.955 $Y=1.345
+ $X2=0 $Y2=0
cc_578 N_A_840_95#_M1042_g N_A_978_67#_c_1217_n 0.0106605f $X=6.29 $Y=2.525
+ $X2=0 $Y2=0
cc_579 N_A_840_95#_M1008_g N_A_978_67#_c_1202_n 0.0103432f $X=5.31 $Y=2.665
+ $X2=0 $Y2=0
cc_580 N_A_840_95#_c_615_n N_A_978_67#_c_1202_n 0.0544652f $X=5.235 $Y=1.34
+ $X2=0 $Y2=0
cc_581 N_A_840_95#_c_617_n N_A_978_67#_c_1202_n 0.0233671f $X=4.597 $Y=1.177
+ $X2=0 $Y2=0
cc_582 N_A_840_95#_c_618_n N_A_978_67#_c_1202_n 0.0726225f $X=4.51 $Y=2.2 $X2=0
+ $Y2=0
cc_583 N_A_840_95#_M1008_g N_A_978_67#_c_1219_n 0.0169887f $X=5.31 $Y=2.665
+ $X2=0 $Y2=0
cc_584 N_A_840_95#_c_615_n N_A_978_67#_c_1219_n 0.001444f $X=5.235 $Y=1.34 $X2=0
+ $Y2=0
cc_585 N_A_840_95#_c_616_n N_A_978_67#_c_1203_n 0.00216685f $X=5.31 $Y=1.34
+ $X2=0 $Y2=0
cc_586 N_A_840_95#_c_616_n N_A_978_67#_c_1204_n 0.0194911f $X=5.31 $Y=1.34 $X2=0
+ $Y2=0
cc_587 N_A_840_95#_M1010_g N_A_978_67#_c_1205_n 0.0189513f $X=5.31 $Y=0.545
+ $X2=0 $Y2=0
cc_588 N_A_840_95#_c_615_n N_A_978_67#_c_1205_n 0.00338038f $X=5.235 $Y=1.34
+ $X2=0 $Y2=0
cc_589 N_A_840_95#_c_617_n N_A_978_67#_c_1205_n 0.0194867f $X=4.597 $Y=1.177
+ $X2=0 $Y2=0
cc_590 N_A_840_95#_c_634_n N_A_2415_137#_M1035_g 0.00576977f $X=11.49 $Y=2.455
+ $X2=0 $Y2=0
cc_591 N_A_840_95#_c_640_n N_A_2415_137#_M1035_g 0.00254833f $X=11.69 $Y=2.98
+ $X2=0 $Y2=0
cc_592 N_A_840_95#_c_642_n N_A_2415_137#_M1035_g 0.00718751f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_593 N_A_840_95#_c_643_n N_A_2415_137#_M1035_g 0.00963765f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_594 N_A_840_95#_c_642_n N_A_2415_137#_c_1360_n 0.0209133f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_595 N_A_840_95#_c_643_n N_A_2415_137#_c_1360_n 0.00114936f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_596 N_A_840_95#_c_642_n N_A_2415_137#_c_1347_n 0.00266035f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_597 N_A_840_95#_c_643_n N_A_2415_137#_c_1347_n 0.0365551f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_598 N_A_840_95#_c_640_n N_A_2211_428#_M1020_d 0.00267852f $X=11.69 $Y=2.98
+ $X2=0 $Y2=0
cc_599 N_A_840_95#_c_634_n N_A_2211_428#_c_1542_n 0.00812282f $X=11.49 $Y=2.455
+ $X2=0 $Y2=0
cc_600 N_A_840_95#_c_637_n N_A_2211_428#_c_1542_n 0.0059583f $X=11.855 $Y=2.305
+ $X2=0 $Y2=0
cc_601 N_A_840_95#_c_639_n N_A_2211_428#_c_1542_n 0.0229716f $X=10.765 $Y=2.895
+ $X2=0 $Y2=0
cc_602 N_A_840_95#_c_640_n N_A_2211_428#_c_1542_n 0.0229954f $X=11.69 $Y=2.98
+ $X2=0 $Y2=0
cc_603 N_A_840_95#_c_627_n N_A_2211_428#_c_1542_n 0.00360382f $X=10.9 $Y=1.18
+ $X2=0 $Y2=0
cc_604 N_A_840_95#_c_639_n N_A_2211_428#_c_1537_n 0.0164529f $X=10.765 $Y=2.895
+ $X2=0 $Y2=0
cc_605 N_A_840_95#_c_642_n N_A_2211_428#_c_1537_n 0.0632549f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_606 N_A_840_95#_c_643_n N_A_2211_428#_c_1537_n 0.00370725f $X=11.855 $Y=1.865
+ $X2=0 $Y2=0
cc_607 N_A_840_95#_c_628_n N_A_2211_428#_c_1537_n 0.00171813f $X=10.955 $Y=1.51
+ $X2=0 $Y2=0
cc_608 N_A_840_95#_c_627_n N_A_2211_428#_c_1538_n 0.0369977f $X=10.9 $Y=1.18
+ $X2=0 $Y2=0
cc_609 N_A_840_95#_c_629_n N_A_2211_428#_c_1538_n 0.0151351f $X=10.955 $Y=1.345
+ $X2=0 $Y2=0
cc_610 N_A_840_95#_c_622_n N_A_1840_21#_M1014_g 0.0129324f $X=9.855 $Y=0.35
+ $X2=0 $Y2=0
cc_611 N_A_840_95#_c_624_n N_A_1840_21#_M1014_g 0.00772074f $X=9.94 $Y=1.095
+ $X2=0 $Y2=0
cc_612 N_A_840_95#_c_626_n N_A_1840_21#_M1014_g 0.00138732f $X=10.025 $Y=1.18
+ $X2=0 $Y2=0
cc_613 N_A_840_95#_c_622_n N_A_1840_21#_c_1627_n 0.0138767f $X=9.855 $Y=0.35
+ $X2=0 $Y2=0
cc_614 N_A_840_95#_c_629_n N_A_1840_21#_c_1627_n 0.0104164f $X=10.955 $Y=1.345
+ $X2=0 $Y2=0
cc_615 N_A_840_95#_c_626_n N_A_1840_21#_c_1630_n 0.00119064f $X=10.025 $Y=1.18
+ $X2=0 $Y2=0
cc_616 N_A_840_95#_M1008_g N_VPWR_c_1893_n 0.00453604f $X=5.31 $Y=2.665 $X2=0
+ $Y2=0
cc_617 N_A_840_95#_c_631_n N_VPWR_c_1893_n 0.0185374f $X=6.215 $Y=3.135 $X2=0
+ $Y2=0
cc_618 N_A_840_95#_c_632_n N_VPWR_c_1893_n 0.00406034f $X=5.385 $Y=3.135 $X2=0
+ $Y2=0
cc_619 N_A_840_95#_M1042_g N_VPWR_c_1893_n 0.00802773f $X=6.29 $Y=2.525 $X2=0
+ $Y2=0
cc_620 N_A_840_95#_c_640_n N_VPWR_c_1896_n 0.00542215f $X=11.69 $Y=2.98 $X2=0
+ $Y2=0
cc_621 N_A_840_95#_c_642_n N_VPWR_c_1896_n 0.0120603f $X=11.855 $Y=1.865 $X2=0
+ $Y2=0
cc_622 N_A_840_95#_c_631_n N_VPWR_c_1909_n 0.0203807f $X=6.215 $Y=3.135 $X2=0
+ $Y2=0
cc_623 N_A_840_95#_c_632_n N_VPWR_c_1913_n 0.00473366f $X=5.385 $Y=3.135 $X2=0
+ $Y2=0
cc_624 N_A_840_95#_c_634_n N_VPWR_c_1914_n 0.00392127f $X=11.49 $Y=2.455 $X2=0
+ $Y2=0
cc_625 N_A_840_95#_c_640_n N_VPWR_c_1914_n 0.0722692f $X=11.69 $Y=2.98 $X2=0
+ $Y2=0
cc_626 N_A_840_95#_c_641_n N_VPWR_c_1914_n 0.0114245f $X=10.85 $Y=2.98 $X2=0
+ $Y2=0
cc_627 N_A_840_95#_c_631_n N_VPWR_c_1889_n 0.023764f $X=6.215 $Y=3.135 $X2=0
+ $Y2=0
cc_628 N_A_840_95#_c_632_n N_VPWR_c_1889_n 0.00585401f $X=5.385 $Y=3.135 $X2=0
+ $Y2=0
cc_629 N_A_840_95#_c_634_n N_VPWR_c_1889_n 0.00542671f $X=11.49 $Y=2.455 $X2=0
+ $Y2=0
cc_630 N_A_840_95#_c_640_n N_VPWR_c_1889_n 0.0431301f $X=11.69 $Y=2.98 $X2=0
+ $Y2=0
cc_631 N_A_840_95#_c_641_n N_VPWR_c_1889_n 0.00589433f $X=10.85 $Y=2.98 $X2=0
+ $Y2=0
cc_632 N_A_840_95#_c_618_n N_A_202_119#_c_2091_n 0.00748703f $X=4.51 $Y=2.2
+ $X2=0 $Y2=0
cc_633 N_A_840_95#_c_618_n N_A_202_119#_c_2092_n 0.0204508f $X=4.51 $Y=2.2 $X2=0
+ $Y2=0
cc_634 N_A_840_95#_M1008_g N_A_202_119#_c_2093_n 0.00433764f $X=5.31 $Y=2.665
+ $X2=0 $Y2=0
cc_635 N_A_840_95#_c_618_n N_A_202_119#_c_2093_n 0.0259156f $X=4.51 $Y=2.2 $X2=0
+ $Y2=0
cc_636 N_A_840_95#_c_618_n N_A_202_119#_c_2147_n 0.0134166f $X=4.51 $Y=2.2 $X2=0
+ $Y2=0
cc_637 N_A_840_95#_c_615_n N_A_202_119#_c_2148_n 5.28327e-19 $X=5.235 $Y=1.34
+ $X2=0 $Y2=0
cc_638 N_A_840_95#_c_618_n N_A_202_119#_c_2148_n 0.0115264f $X=4.51 $Y=2.2 $X2=0
+ $Y2=0
cc_639 N_A_840_95#_M1008_g N_A_202_119#_c_2087_n 0.00629886f $X=5.31 $Y=2.665
+ $X2=0 $Y2=0
cc_640 N_A_840_95#_M1042_g N_A_202_119#_c_2087_n 0.00338222f $X=6.29 $Y=2.525
+ $X2=0 $Y2=0
cc_641 N_A_840_95#_c_616_n N_A_202_119#_c_2087_n 0.00463241f $X=5.31 $Y=1.34
+ $X2=0 $Y2=0
cc_642 N_A_840_95#_M1010_g N_A_202_119#_c_2088_n 0.00979493f $X=5.31 $Y=0.545
+ $X2=0 $Y2=0
cc_643 N_A_840_95#_c_612_n N_A_202_119#_c_2088_n 0.00577498f $X=6.645 $Y=0.185
+ $X2=0 $Y2=0
cc_644 N_A_840_95#_M1008_g N_A_202_119#_c_2097_n 0.0159394f $X=5.31 $Y=2.665
+ $X2=0 $Y2=0
cc_645 N_A_840_95#_c_631_n N_A_202_119#_c_2097_n 0.00568785f $X=6.215 $Y=3.135
+ $X2=0 $Y2=0
cc_646 N_A_840_95#_M1008_g N_A_202_119#_c_2098_n 0.00500765f $X=5.31 $Y=2.665
+ $X2=0 $Y2=0
cc_647 N_A_840_95#_c_631_n N_A_202_119#_c_2098_n 0.00431984f $X=6.215 $Y=3.135
+ $X2=0 $Y2=0
cc_648 N_A_840_95#_M1042_g N_A_202_119#_c_2098_n 0.0067875f $X=6.29 $Y=2.525
+ $X2=0 $Y2=0
cc_649 N_A_840_95#_c_639_n A_2116_379# 0.0197069f $X=10.765 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_650 N_A_840_95#_c_641_n A_2116_379# 0.00404611f $X=10.85 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_651 N_A_840_95#_c_640_n A_2313_506# 0.00269361f $X=11.69 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_652 N_A_840_95#_c_642_n A_2313_506# 0.013752f $X=11.855 $Y=1.865 $X2=-0.19
+ $Y2=-0.245
cc_653 N_A_840_95#_c_656_p N_VGND_M1017_d 0.0269007f $X=7.975 $Y=0.915 $X2=0
+ $Y2=0
cc_654 N_A_840_95#_c_621_n N_VGND_M1017_d 0.00718615f $X=8.06 $Y=0.83 $X2=0
+ $Y2=0
cc_655 N_A_840_95#_c_625_n N_VGND_M1046_s 0.00495367f $X=10.68 $Y=1.18 $X2=0
+ $Y2=0
cc_656 N_A_840_95#_c_617_n N_VGND_c_2293_n 0.0187201f $X=4.597 $Y=1.177 $X2=0
+ $Y2=0
cc_657 N_A_840_95#_M1010_g N_VGND_c_2294_n 0.00736357f $X=5.31 $Y=0.545 $X2=0
+ $Y2=0
cc_658 N_A_840_95#_c_612_n N_VGND_c_2294_n 0.0197174f $X=6.645 $Y=0.185 $X2=0
+ $Y2=0
cc_659 N_A_840_95#_c_613_n N_VGND_c_2294_n 0.00332703f $X=5.385 $Y=0.185 $X2=0
+ $Y2=0
cc_660 N_A_840_95#_c_612_n N_VGND_c_2295_n 0.00887494f $X=6.645 $Y=0.185 $X2=0
+ $Y2=0
cc_661 N_A_840_95#_c_656_p N_VGND_c_2295_n 0.0248838f $X=7.975 $Y=0.915 $X2=0
+ $Y2=0
cc_662 N_A_840_95#_c_621_n N_VGND_c_2295_n 0.0157982f $X=8.06 $Y=0.83 $X2=0
+ $Y2=0
cc_663 N_A_840_95#_c_623_n N_VGND_c_2295_n 0.0144408f $X=8.145 $Y=0.35 $X2=0
+ $Y2=0
cc_664 N_A_840_95#_c_622_n N_VGND_c_2296_n 0.0141601f $X=9.855 $Y=0.35 $X2=0
+ $Y2=0
cc_665 N_A_840_95#_c_624_n N_VGND_c_2296_n 0.0352568f $X=9.94 $Y=1.095 $X2=0
+ $Y2=0
cc_666 N_A_840_95#_c_625_n N_VGND_c_2296_n 0.0135261f $X=10.68 $Y=1.18 $X2=0
+ $Y2=0
cc_667 N_A_840_95#_c_629_n N_VGND_c_2296_n 0.00212381f $X=10.955 $Y=1.345 $X2=0
+ $Y2=0
cc_668 N_A_840_95#_c_612_n N_VGND_c_2305_n 0.0336803f $X=6.645 $Y=0.185 $X2=0
+ $Y2=0
cc_669 N_A_840_95#_c_613_n N_VGND_c_2310_n 0.00559147f $X=5.385 $Y=0.185 $X2=0
+ $Y2=0
cc_670 N_A_840_95#_c_617_n N_VGND_c_2310_n 0.0128629f $X=4.597 $Y=1.177 $X2=0
+ $Y2=0
cc_671 N_A_840_95#_c_622_n N_VGND_c_2311_n 0.114649f $X=9.855 $Y=0.35 $X2=0
+ $Y2=0
cc_672 N_A_840_95#_c_623_n N_VGND_c_2311_n 0.0114622f $X=8.145 $Y=0.35 $X2=0
+ $Y2=0
cc_673 N_A_840_95#_c_612_n N_VGND_c_2322_n 0.0457019f $X=6.645 $Y=0.185 $X2=0
+ $Y2=0
cc_674 N_A_840_95#_c_613_n N_VGND_c_2322_n 0.0109933f $X=5.385 $Y=0.185 $X2=0
+ $Y2=0
cc_675 N_A_840_95#_c_617_n N_VGND_c_2322_n 0.0143408f $X=4.597 $Y=1.177 $X2=0
+ $Y2=0
cc_676 N_A_840_95#_c_656_p N_VGND_c_2322_n 0.0250258f $X=7.975 $Y=0.915 $X2=0
+ $Y2=0
cc_677 N_A_840_95#_c_817_p N_VGND_c_2322_n 0.00680238f $X=6.945 $Y=0.915 $X2=0
+ $Y2=0
cc_678 N_A_840_95#_c_622_n N_VGND_c_2322_n 0.0670691f $X=9.855 $Y=0.35 $X2=0
+ $Y2=0
cc_679 N_A_840_95#_c_623_n N_VGND_c_2322_n 0.00657784f $X=8.145 $Y=0.35 $X2=0
+ $Y2=0
cc_680 N_A_840_95#_c_629_n N_VGND_c_2322_n 9.39239e-19 $X=10.955 $Y=1.345 $X2=0
+ $Y2=0
cc_681 N_A_840_95#_c_619_n A_1359_137# 0.00136016f $X=6.855 $Y=1.38 $X2=-0.19
+ $Y2=-0.245
cc_682 N_A_840_95#_c_656_p A_1359_137# 0.0123613f $X=7.975 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_683 N_A_840_95#_c_817_p A_1359_137# 0.00217934f $X=6.945 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_684 N_A_840_95#_c_622_n N_A_1670_93#_c_2482_n 0.0407794f $X=9.855 $Y=0.35
+ $X2=0 $Y2=0
cc_685 N_A_840_95#_c_622_n N_A_1670_93#_c_2483_n 0.0190834f $X=9.855 $Y=0.35
+ $X2=0 $Y2=0
cc_686 N_A_840_95#_c_622_n N_A_1670_93#_c_2481_n 0.0207318f $X=9.855 $Y=0.35
+ $X2=0 $Y2=0
cc_687 N_A_840_95#_c_624_n N_A_1670_93#_c_2481_n 0.0198001f $X=9.94 $Y=1.095
+ $X2=0 $Y2=0
cc_688 N_A_840_95#_c_625_n A_2116_119# 0.00196198f $X=10.68 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_689 N_A_840_95#_c_627_n A_2116_119# 0.00939045f $X=10.9 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_690 N_A_1423_401#_c_843_n N_SET_B_M1043_g 0.00106169f $X=7.565 $Y=1.99 $X2=0
+ $Y2=0
cc_691 N_A_1423_401#_c_844_n N_SET_B_M1043_g 0.0163532f $X=8.525 $Y=2.415 $X2=0
+ $Y2=0
cc_692 N_A_1423_401#_c_845_n N_SET_B_M1043_g 0.00885321f $X=9.245 $Y=2.415 $X2=0
+ $Y2=0
cc_693 N_A_1423_401#_c_848_n N_SET_B_M1043_g 0.0073047f $X=7.335 $Y=1.99 $X2=0
+ $Y2=0
cc_694 N_A_1423_401#_M1029_d N_SET_B_c_956_n 0.00192085f $X=8.8 $Y=0.465 $X2=0
+ $Y2=0
cc_695 N_A_1423_401#_M1046_g N_SET_B_c_956_n 0.00621779f $X=10.505 $Y=0.915
+ $X2=0 $Y2=0
cc_696 N_A_1423_401#_c_832_n N_SET_B_c_956_n 0.0172349f $X=9.16 $Y=1.095 $X2=0
+ $Y2=0
cc_697 N_A_1423_401#_c_833_n N_SET_B_c_956_n 0.0185608f $X=9.245 $Y=1.445 $X2=0
+ $Y2=0
cc_698 N_A_1423_401#_c_837_n N_SET_B_c_956_n 0.00677778f $X=10.335 $Y=1.57 $X2=0
+ $Y2=0
cc_699 N_A_1423_401#_c_838_n N_SET_B_c_956_n 0.0384134f $X=10.17 $Y=1.575 $X2=0
+ $Y2=0
cc_700 N_A_1423_401#_c_832_n N_SET_B_c_957_n 0.00125044f $X=9.16 $Y=1.095 $X2=0
+ $Y2=0
cc_701 N_A_1423_401#_c_833_n N_SET_B_c_957_n 8.65672e-19 $X=9.245 $Y=1.445 $X2=0
+ $Y2=0
cc_702 N_A_1423_401#_M1017_g N_SET_B_c_960_n 0.0066645f $X=7.335 $Y=0.895 $X2=0
+ $Y2=0
cc_703 N_A_1423_401#_c_832_n N_SET_B_c_961_n 0.001634f $X=9.16 $Y=1.095 $X2=0
+ $Y2=0
cc_704 N_A_1423_401#_c_833_n N_SET_B_c_961_n 0.00280898f $X=9.245 $Y=1.445 $X2=0
+ $Y2=0
cc_705 N_A_1423_401#_c_832_n N_A_1273_137#_M1029_g 0.00374836f $X=9.16 $Y=1.095
+ $X2=0 $Y2=0
cc_706 N_A_1423_401#_c_833_n N_A_1273_137#_M1029_g 0.00111894f $X=9.245 $Y=1.445
+ $X2=0 $Y2=0
cc_707 N_A_1423_401#_c_834_n N_A_1273_137#_M1033_g 0.00360061f $X=9.245 $Y=2.075
+ $X2=0 $Y2=0
cc_708 N_A_1423_401#_c_845_n N_A_1273_137#_M1033_g 0.0208571f $X=9.245 $Y=2.415
+ $X2=0 $Y2=0
cc_709 N_A_1423_401#_M1017_g N_A_1273_137#_c_1087_n 0.00120048f $X=7.335
+ $Y=0.895 $X2=0 $Y2=0
cc_710 N_A_1423_401#_M1018_g N_A_1273_137#_c_1095_n 0.00252509f $X=7.19 $Y=2.525
+ $X2=0 $Y2=0
cc_711 N_A_1423_401#_M1018_g N_A_1273_137#_c_1096_n 0.0107584f $X=7.19 $Y=2.525
+ $X2=0 $Y2=0
cc_712 N_A_1423_401#_c_843_n N_A_1273_137#_c_1096_n 0.0131692f $X=7.565 $Y=1.99
+ $X2=0 $Y2=0
cc_713 N_A_1423_401#_c_848_n N_A_1273_137#_c_1096_n 0.00416615f $X=7.335 $Y=1.99
+ $X2=0 $Y2=0
cc_714 N_A_1423_401#_M1017_g N_A_1273_137#_c_1097_n 0.00644982f $X=7.335
+ $Y=0.895 $X2=0 $Y2=0
cc_715 N_A_1423_401#_c_843_n N_A_1273_137#_c_1097_n 0.0162251f $X=7.565 $Y=1.99
+ $X2=0 $Y2=0
cc_716 N_A_1423_401#_c_848_n N_A_1273_137#_c_1097_n 0.0107091f $X=7.335 $Y=1.99
+ $X2=0 $Y2=0
cc_717 N_A_1423_401#_M1017_g N_A_1273_137#_c_1088_n 0.0127532f $X=7.335 $Y=0.895
+ $X2=0 $Y2=0
cc_718 N_A_1423_401#_c_843_n N_A_1273_137#_c_1088_n 0.0131135f $X=7.565 $Y=1.99
+ $X2=0 $Y2=0
cc_719 N_A_1423_401#_c_844_n N_A_1273_137#_c_1088_n 0.00684551f $X=8.525
+ $Y=2.415 $X2=0 $Y2=0
cc_720 N_A_1423_401#_c_848_n N_A_1273_137#_c_1088_n 0.00559748f $X=7.335 $Y=1.99
+ $X2=0 $Y2=0
cc_721 N_A_1423_401#_M1017_g N_A_1273_137#_c_1089_n 0.00358564f $X=7.335
+ $Y=0.895 $X2=0 $Y2=0
cc_722 N_A_1423_401#_M1043_d N_A_1273_137#_c_1098_n 0.00139513f $X=8.41 $Y=1.895
+ $X2=0 $Y2=0
cc_723 N_A_1423_401#_c_834_n N_A_1273_137#_c_1098_n 0.0129673f $X=9.245 $Y=2.075
+ $X2=0 $Y2=0
cc_724 N_A_1423_401#_c_844_n N_A_1273_137#_c_1098_n 0.0461463f $X=8.525 $Y=2.415
+ $X2=0 $Y2=0
cc_725 N_A_1423_401#_c_845_n N_A_1273_137#_c_1098_n 0.0197787f $X=9.245 $Y=2.415
+ $X2=0 $Y2=0
cc_726 N_A_1423_401#_c_832_n N_A_1273_137#_c_1090_n 0.0082847f $X=9.16 $Y=1.095
+ $X2=0 $Y2=0
cc_727 N_A_1423_401#_c_833_n N_A_1273_137#_c_1090_n 0.00279404f $X=9.245
+ $Y=1.445 $X2=0 $Y2=0
cc_728 N_A_1423_401#_c_834_n N_A_1273_137#_c_1090_n 0.00773912f $X=9.245
+ $Y=2.075 $X2=0 $Y2=0
cc_729 N_A_1423_401#_c_835_n N_A_1273_137#_c_1090_n 0.0135641f $X=9.245 $Y=1.53
+ $X2=0 $Y2=0
cc_730 N_A_1423_401#_c_832_n N_A_1273_137#_c_1091_n 0.00102285f $X=9.16 $Y=1.095
+ $X2=0 $Y2=0
cc_731 N_A_1423_401#_c_833_n N_A_1273_137#_c_1091_n 2.24878e-19 $X=9.245
+ $Y=1.445 $X2=0 $Y2=0
cc_732 N_A_1423_401#_c_834_n N_A_1273_137#_c_1091_n 0.00114398f $X=9.245
+ $Y=2.075 $X2=0 $Y2=0
cc_733 N_A_1423_401#_c_845_n N_A_1273_137#_c_1091_n 8.48333e-19 $X=9.245
+ $Y=2.415 $X2=0 $Y2=0
cc_734 N_A_1423_401#_c_835_n N_A_1273_137#_c_1091_n 0.00111656f $X=9.245 $Y=1.53
+ $X2=0 $Y2=0
cc_735 N_A_1423_401#_M1017_g N_A_1273_137#_c_1092_n 0.00335664f $X=7.335
+ $Y=0.895 $X2=0 $Y2=0
cc_736 N_A_1423_401#_c_843_n N_A_1273_137#_c_1092_n 0.0048158f $X=7.565 $Y=1.99
+ $X2=0 $Y2=0
cc_737 N_A_1423_401#_c_844_n N_A_1273_137#_c_1092_n 0.0130131f $X=8.525 $Y=2.415
+ $X2=0 $Y2=0
cc_738 N_A_1423_401#_c_848_n N_A_1273_137#_c_1092_n 7.76342e-19 $X=7.335 $Y=1.99
+ $X2=0 $Y2=0
cc_739 N_A_1423_401#_M1017_g N_A_978_67#_c_1209_n 0.00302047f $X=7.335 $Y=0.895
+ $X2=0 $Y2=0
cc_740 N_A_1423_401#_c_848_n N_A_978_67#_M1045_g 0.0498329f $X=7.335 $Y=1.99
+ $X2=0 $Y2=0
cc_741 N_A_1423_401#_M1018_g N_A_978_67#_c_1211_n 0.0104164f $X=7.19 $Y=2.525
+ $X2=0 $Y2=0
cc_742 N_A_1423_401#_M1039_g N_A_978_67#_c_1211_n 0.0104164f $X=10.505 $Y=2.315
+ $X2=0 $Y2=0
cc_743 N_A_1423_401#_c_845_n N_A_978_67#_c_1211_n 0.011757f $X=9.245 $Y=2.415
+ $X2=0 $Y2=0
cc_744 N_A_1423_401#_M1039_g N_A_978_67#_c_1215_n 0.0273224f $X=10.505 $Y=2.315
+ $X2=0 $Y2=0
cc_745 N_A_1423_401#_c_832_n N_A_1840_21#_M1014_g 0.00742347f $X=9.16 $Y=1.095
+ $X2=0 $Y2=0
cc_746 N_A_1423_401#_c_833_n N_A_1840_21#_M1005_g 0.0054016f $X=9.245 $Y=1.445
+ $X2=0 $Y2=0
cc_747 N_A_1423_401#_c_834_n N_A_1840_21#_M1005_g 0.0176872f $X=9.245 $Y=2.075
+ $X2=0 $Y2=0
cc_748 N_A_1423_401#_c_845_n N_A_1840_21#_M1005_g 0.0199619f $X=9.245 $Y=2.415
+ $X2=0 $Y2=0
cc_749 N_A_1423_401#_c_835_n N_A_1840_21#_M1005_g 0.00242835f $X=9.245 $Y=1.53
+ $X2=0 $Y2=0
cc_750 N_A_1423_401#_c_838_n N_A_1840_21#_M1005_g 0.00709967f $X=10.17 $Y=1.575
+ $X2=0 $Y2=0
cc_751 N_A_1423_401#_M1046_g N_A_1840_21#_c_1627_n 0.0103107f $X=10.505 $Y=0.915
+ $X2=0 $Y2=0
cc_752 N_A_1423_401#_c_832_n N_A_1840_21#_c_1630_n 0.00179995f $X=9.16 $Y=1.095
+ $X2=0 $Y2=0
cc_753 N_A_1423_401#_c_833_n N_A_1840_21#_c_1630_n 0.00393763f $X=9.245 $Y=1.445
+ $X2=0 $Y2=0
cc_754 N_A_1423_401#_c_844_n N_VPWR_M1018_d 0.00582972f $X=8.525 $Y=2.415 $X2=0
+ $Y2=0
cc_755 N_A_1423_401#_M1018_g N_VPWR_c_1894_n 0.00956232f $X=7.19 $Y=2.525 $X2=0
+ $Y2=0
cc_756 N_A_1423_401#_c_844_n N_VPWR_c_1894_n 0.0209859f $X=8.525 $Y=2.415 $X2=0
+ $Y2=0
cc_757 N_A_1423_401#_c_845_n N_VPWR_c_1894_n 0.0208698f $X=9.245 $Y=2.415 $X2=0
+ $Y2=0
cc_758 N_A_1423_401#_M1039_g N_VPWR_c_1895_n 0.0237369f $X=10.505 $Y=2.315 $X2=0
+ $Y2=0
cc_759 N_A_1423_401#_c_834_n N_VPWR_c_1895_n 0.0141919f $X=9.245 $Y=2.075 $X2=0
+ $Y2=0
cc_760 N_A_1423_401#_c_845_n N_VPWR_c_1895_n 0.0534686f $X=9.245 $Y=2.415 $X2=0
+ $Y2=0
cc_761 N_A_1423_401#_c_838_n N_VPWR_c_1895_n 0.0186383f $X=10.17 $Y=1.575 $X2=0
+ $Y2=0
cc_762 N_A_1423_401#_c_845_n N_VPWR_c_1911_n 0.0178647f $X=9.245 $Y=2.415 $X2=0
+ $Y2=0
cc_763 N_A_1423_401#_M1018_g N_VPWR_c_1889_n 9.39239e-19 $X=7.19 $Y=2.525 $X2=0
+ $Y2=0
cc_764 N_A_1423_401#_M1039_g N_VPWR_c_1889_n 9.39239e-19 $X=10.505 $Y=2.315
+ $X2=0 $Y2=0
cc_765 N_A_1423_401#_c_845_n N_VPWR_c_1889_n 0.0220065f $X=9.245 $Y=2.415 $X2=0
+ $Y2=0
cc_766 N_A_1423_401#_c_834_n A_1796_379# 0.00210186f $X=9.245 $Y=2.075 $X2=-0.19
+ $Y2=-0.245
cc_767 N_A_1423_401#_c_845_n A_1796_379# 0.00559173f $X=9.245 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_768 N_A_1423_401#_M1017_g N_VGND_c_2295_n 0.00399502f $X=7.335 $Y=0.895 $X2=0
+ $Y2=0
cc_769 N_A_1423_401#_M1046_g N_VGND_c_2296_n 0.0115035f $X=10.505 $Y=0.915 $X2=0
+ $Y2=0
cc_770 N_A_1423_401#_M1017_g N_VGND_c_2305_n 0.00385058f $X=7.335 $Y=0.895 $X2=0
+ $Y2=0
cc_771 N_A_1423_401#_M1017_g N_VGND_c_2322_n 0.00453162f $X=7.335 $Y=0.895 $X2=0
+ $Y2=0
cc_772 N_A_1423_401#_M1046_g N_VGND_c_2322_n 7.88961e-19 $X=10.505 $Y=0.915
+ $X2=0 $Y2=0
cc_773 N_A_1423_401#_M1029_d N_A_1670_93#_c_2482_n 0.00627361f $X=8.8 $Y=0.465
+ $X2=0 $Y2=0
cc_774 N_A_1423_401#_c_832_n N_A_1670_93#_c_2482_n 0.0257513f $X=9.16 $Y=1.095
+ $X2=0 $Y2=0
cc_775 N_A_1423_401#_c_838_n N_A_1670_93#_c_2481_n 0.00396532f $X=10.17 $Y=1.575
+ $X2=0 $Y2=0
cc_776 N_SET_B_c_954_n N_A_1273_137#_M1029_g 0.0206637f $X=8.275 $Y=1.215 $X2=0
+ $Y2=0
cc_777 N_SET_B_c_956_n N_A_1273_137#_M1029_g 0.00584289f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_778 N_SET_B_c_957_n N_A_1273_137#_M1029_g 0.00141383f $X=8.545 $Y=1.295 $X2=0
+ $Y2=0
cc_779 N_SET_B_c_960_n N_A_1273_137#_M1029_g 0.0210216f $X=8.275 $Y=1.38 $X2=0
+ $Y2=0
cc_780 N_SET_B_c_961_n N_A_1273_137#_M1029_g 0.00279424f $X=8.275 $Y=1.38 $X2=0
+ $Y2=0
cc_781 N_SET_B_M1043_g N_A_1273_137#_M1033_g 0.0205992f $X=8.335 $Y=2.315 $X2=0
+ $Y2=0
cc_782 N_SET_B_M1043_g N_A_1273_137#_c_1098_n 0.0120637f $X=8.335 $Y=2.315 $X2=0
+ $Y2=0
cc_783 N_SET_B_c_956_n N_A_1273_137#_c_1098_n 0.00560714f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_784 N_SET_B_c_957_n N_A_1273_137#_c_1098_n 0.0025993f $X=8.545 $Y=1.295 $X2=0
+ $Y2=0
cc_785 N_SET_B_c_960_n N_A_1273_137#_c_1098_n 0.00536011f $X=8.275 $Y=1.38 $X2=0
+ $Y2=0
cc_786 N_SET_B_c_961_n N_A_1273_137#_c_1098_n 0.0223937f $X=8.275 $Y=1.38 $X2=0
+ $Y2=0
cc_787 N_SET_B_M1043_g N_A_1273_137#_c_1090_n 0.00102711f $X=8.335 $Y=2.315
+ $X2=0 $Y2=0
cc_788 N_SET_B_c_956_n N_A_1273_137#_c_1090_n 0.00881073f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_789 N_SET_B_c_961_n N_A_1273_137#_c_1090_n 0.00996286f $X=8.275 $Y=1.38 $X2=0
+ $Y2=0
cc_790 N_SET_B_M1043_g N_A_1273_137#_c_1091_n 0.0101643f $X=8.335 $Y=2.315 $X2=0
+ $Y2=0
cc_791 N_SET_B_M1043_g N_A_1273_137#_c_1092_n 0.00611099f $X=8.335 $Y=2.315
+ $X2=0 $Y2=0
cc_792 N_SET_B_c_960_n N_A_1273_137#_c_1092_n 8.75061e-19 $X=8.275 $Y=1.38 $X2=0
+ $Y2=0
cc_793 N_SET_B_c_961_n N_A_1273_137#_c_1092_n 0.00498982f $X=8.275 $Y=1.38 $X2=0
+ $Y2=0
cc_794 N_SET_B_M1043_g N_A_978_67#_c_1211_n 0.0103107f $X=8.335 $Y=2.315 $X2=0
+ $Y2=0
cc_795 N_SET_B_c_956_n N_A_978_67#_c_1214_n 0.00306946f $X=12.575 $Y=1.295 $X2=0
+ $Y2=0
cc_796 N_SET_B_c_956_n N_A_978_67#_c_1199_n 0.0113366f $X=12.575 $Y=1.295 $X2=0
+ $Y2=0
cc_797 N_SET_B_c_956_n N_A_978_67#_c_1200_n 5.46722e-19 $X=12.575 $Y=1.295 $X2=0
+ $Y2=0
cc_798 N_SET_B_c_956_n N_A_978_67#_c_1201_n 0.00307148f $X=12.575 $Y=1.295 $X2=0
+ $Y2=0
cc_799 N_SET_B_c_956_n N_A_2415_137#_c_1329_n 0.00314005f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_800 N_SET_B_c_958_n N_A_2415_137#_c_1329_n 6.53386e-19 $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_801 N_SET_B_c_959_n N_A_2415_137#_c_1329_n 0.00172105f $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_802 N_SET_B_c_963_n N_A_2415_137#_c_1329_n 0.0159102f $X=12.785 $Y=1.345
+ $X2=0 $Y2=0
cc_803 N_SET_B_c_966_n N_A_2415_137#_M1035_g 0.00975519f $X=13.065 $Y=2.18 $X2=0
+ $Y2=0
cc_804 N_SET_B_c_956_n N_A_2415_137#_c_1341_n 0.0106156f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_805 N_SET_B_c_958_n N_A_2415_137#_c_1341_n 6.81397e-19 $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_806 N_SET_B_c_959_n N_A_2415_137#_c_1341_n 0.00892458f $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_807 N_SET_B_c_962_n N_A_2415_137#_c_1341_n 0.0169861f $X=12.785 $Y=1.51 $X2=0
+ $Y2=0
cc_808 N_SET_B_c_963_n N_A_2415_137#_c_1341_n 0.00131804f $X=12.785 $Y=1.345
+ $X2=0 $Y2=0
cc_809 N_SET_B_c_966_n N_A_2415_137#_c_1356_n 0.00885285f $X=13.065 $Y=2.18
+ $X2=0 $Y2=0
cc_810 N_SET_B_c_967_n N_A_2415_137#_c_1356_n 0.0148444f $X=13.065 $Y=2.105
+ $X2=0 $Y2=0
cc_811 N_SET_B_c_959_n N_A_2415_137#_c_1356_n 0.0164459f $X=12.72 $Y=1.295 $X2=0
+ $Y2=0
cc_812 N_SET_B_c_962_n N_A_2415_137#_c_1356_n 8.94052e-19 $X=12.785 $Y=1.51
+ $X2=0 $Y2=0
cc_813 N_SET_B_c_965_n N_A_2415_137#_c_1360_n 0.00108547f $X=12.875 $Y=2.03
+ $X2=0 $Y2=0
cc_814 N_SET_B_c_956_n N_A_2415_137#_c_1360_n 0.00901802f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_815 N_SET_B_c_965_n N_A_2415_137#_c_1361_n 0.0124944f $X=12.875 $Y=2.03 $X2=0
+ $Y2=0
cc_816 N_SET_B_c_966_n N_A_2415_137#_c_1361_n 0.00273172f $X=13.065 $Y=2.18
+ $X2=0 $Y2=0
cc_817 N_SET_B_c_966_n N_A_2415_137#_c_1362_n 0.0102105f $X=13.065 $Y=2.18 $X2=0
+ $Y2=0
cc_818 N_SET_B_c_967_n N_A_2415_137#_c_1362_n 0.00175167f $X=13.065 $Y=2.105
+ $X2=0 $Y2=0
cc_819 N_SET_B_c_966_n N_A_2415_137#_c_1392_n 0.0070004f $X=13.065 $Y=2.18 $X2=0
+ $Y2=0
cc_820 N_SET_B_c_965_n N_A_2415_137#_c_1347_n 0.00872223f $X=12.875 $Y=2.03
+ $X2=0 $Y2=0
cc_821 N_SET_B_c_956_n N_A_2211_428#_M1022_d 0.00729998f $X=12.575 $Y=1.295
+ $X2=-0.19 $Y2=-0.245
cc_822 N_SET_B_c_962_n N_A_2211_428#_M1047_g 0.00300062f $X=12.785 $Y=1.51 $X2=0
+ $Y2=0
cc_823 N_SET_B_c_963_n N_A_2211_428#_M1047_g 0.0187382f $X=12.785 $Y=1.345 $X2=0
+ $Y2=0
cc_824 N_SET_B_c_965_n N_A_2211_428#_M1000_g 0.00758145f $X=12.875 $Y=2.03 $X2=0
+ $Y2=0
cc_825 N_SET_B_c_967_n N_A_2211_428#_M1000_g 0.0220163f $X=13.065 $Y=2.105 $X2=0
+ $Y2=0
cc_826 N_SET_B_c_956_n N_A_2211_428#_c_1563_n 0.0383524f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_827 N_SET_B_c_958_n N_A_2211_428#_c_1563_n 0.00335616f $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_828 N_SET_B_c_959_n N_A_2211_428#_c_1563_n 0.0147976f $X=12.72 $Y=1.295 $X2=0
+ $Y2=0
cc_829 N_SET_B_c_962_n N_A_2211_428#_c_1563_n 6.51766e-19 $X=12.785 $Y=1.51
+ $X2=0 $Y2=0
cc_830 N_SET_B_c_963_n N_A_2211_428#_c_1563_n 0.0114057f $X=12.785 $Y=1.345
+ $X2=0 $Y2=0
cc_831 N_SET_B_c_958_n N_A_2211_428#_c_1536_n 0.00136221f $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_832 N_SET_B_c_959_n N_A_2211_428#_c_1536_n 0.0193707f $X=12.72 $Y=1.295 $X2=0
+ $Y2=0
cc_833 N_SET_B_c_962_n N_A_2211_428#_c_1536_n 8.23359e-19 $X=12.785 $Y=1.51
+ $X2=0 $Y2=0
cc_834 N_SET_B_c_963_n N_A_2211_428#_c_1536_n 0.0040614f $X=12.785 $Y=1.345
+ $X2=0 $Y2=0
cc_835 N_SET_B_c_956_n N_A_2211_428#_c_1537_n 0.0147792f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_836 N_SET_B_c_956_n N_A_2211_428#_c_1538_n 0.0238597f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_837 N_SET_B_c_967_n N_A_2211_428#_c_1539_n 2.64677e-19 $X=13.065 $Y=2.105
+ $X2=0 $Y2=0
cc_838 N_SET_B_c_959_n N_A_2211_428#_c_1539_n 0.0244811f $X=12.72 $Y=1.295 $X2=0
+ $Y2=0
cc_839 N_SET_B_c_962_n N_A_2211_428#_c_1539_n 0.00197133f $X=12.785 $Y=1.51
+ $X2=0 $Y2=0
cc_840 N_SET_B_c_959_n N_A_2211_428#_c_1540_n 3.74311e-19 $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_841 N_SET_B_c_962_n N_A_2211_428#_c_1540_n 0.0202901f $X=12.785 $Y=1.51 $X2=0
+ $Y2=0
cc_842 N_SET_B_c_956_n N_A_1840_21#_M1005_g 8.79627e-19 $X=12.575 $Y=1.295 $X2=0
+ $Y2=0
cc_843 N_SET_B_c_963_n N_A_1840_21#_c_1627_n 0.0100396f $X=12.785 $Y=1.345 $X2=0
+ $Y2=0
cc_844 N_SET_B_c_956_n N_A_1840_21#_c_1630_n 0.00207442f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_845 N_SET_B_M1043_g N_VPWR_c_1894_n 0.00937708f $X=8.335 $Y=2.315 $X2=0 $Y2=0
cc_846 N_SET_B_c_966_n N_VPWR_c_1896_n 0.00645378f $X=13.065 $Y=2.18 $X2=0 $Y2=0
cc_847 N_SET_B_c_967_n N_VPWR_c_1896_n 7.96395e-19 $X=13.065 $Y=2.105 $X2=0
+ $Y2=0
cc_848 N_SET_B_c_966_n N_VPWR_c_1915_n 0.00549284f $X=13.065 $Y=2.18 $X2=0 $Y2=0
cc_849 N_SET_B_M1043_g N_VPWR_c_1889_n 7.88961e-19 $X=8.335 $Y=2.315 $X2=0 $Y2=0
cc_850 N_SET_B_c_966_n N_VPWR_c_1889_n 0.0113256f $X=13.065 $Y=2.18 $X2=0 $Y2=0
cc_851 N_SET_B_c_956_n N_VGND_M1037_d 0.00293216f $X=12.575 $Y=1.295 $X2=0 $Y2=0
cc_852 N_SET_B_c_958_n N_VGND_M1037_d 0.00153626f $X=12.72 $Y=1.295 $X2=0 $Y2=0
cc_853 N_SET_B_c_959_n N_VGND_M1037_d 0.00122482f $X=12.72 $Y=1.295 $X2=0 $Y2=0
cc_854 N_SET_B_c_954_n N_VGND_c_2295_n 8.31682e-19 $X=8.275 $Y=1.215 $X2=0 $Y2=0
cc_855 N_SET_B_c_956_n N_VGND_c_2296_n 0.00156661f $X=12.575 $Y=1.295 $X2=0
+ $Y2=0
cc_856 N_SET_B_c_963_n N_VGND_c_2297_n 0.00415562f $X=12.785 $Y=1.345 $X2=0
+ $Y2=0
cc_857 N_SET_B_c_954_n N_VGND_c_2311_n 7.85522e-19 $X=8.275 $Y=1.215 $X2=0 $Y2=0
cc_858 N_SET_B_c_963_n N_VGND_c_2322_n 9.39239e-19 $X=12.785 $Y=1.345 $X2=0
+ $Y2=0
cc_859 N_SET_B_c_956_n N_A_1670_93#_c_2482_n 0.00565957f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_860 N_SET_B_c_954_n N_A_1670_93#_c_2483_n 0.004849f $X=8.275 $Y=1.215 $X2=0
+ $Y2=0
cc_861 N_SET_B_c_956_n N_A_1670_93#_c_2483_n 0.00500868f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_862 N_SET_B_c_957_n N_A_1670_93#_c_2483_n 0.00669705f $X=8.545 $Y=1.295 $X2=0
+ $Y2=0
cc_863 N_SET_B_c_960_n N_A_1670_93#_c_2483_n 4.60607e-19 $X=8.275 $Y=1.38 $X2=0
+ $Y2=0
cc_864 N_SET_B_c_961_n N_A_1670_93#_c_2483_n 0.0104851f $X=8.275 $Y=1.38 $X2=0
+ $Y2=0
cc_865 N_SET_B_c_956_n N_A_1670_93#_c_2481_n 0.00823565f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_866 N_SET_B_c_956_n A_2367_163# 0.00201638f $X=12.575 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_867 N_SET_B_c_959_n N_A_2574_119#_M1030_d 7.21505e-19 $X=12.72 $Y=1.295
+ $X2=-0.19 $Y2=-0.245
cc_868 N_SET_B_c_963_n N_A_2574_119#_c_2509_n 0.00175602f $X=12.785 $Y=1.345
+ $X2=0 $Y2=0
cc_869 N_A_1273_137#_c_1087_n N_A_978_67#_M1011_g 0.0089045f $X=6.505 $Y=0.895
+ $X2=0 $Y2=0
cc_870 N_A_1273_137#_c_1087_n N_A_978_67#_c_1209_n 0.0155037f $X=6.505 $Y=0.895
+ $X2=0 $Y2=0
cc_871 N_A_1273_137#_c_1097_n N_A_978_67#_c_1209_n 0.00212164f $X=7.21 $Y=2.075
+ $X2=0 $Y2=0
cc_872 N_A_1273_137#_c_1100_n N_A_978_67#_c_1209_n 0.00573373f $X=6.585 $Y=2.16
+ $X2=0 $Y2=0
cc_873 N_A_1273_137#_c_1087_n N_A_978_67#_M1045_g 0.00308693f $X=6.505 $Y=0.895
+ $X2=0 $Y2=0
cc_874 N_A_1273_137#_c_1095_n N_A_978_67#_M1045_g 0.0109527f $X=6.585 $Y=2.525
+ $X2=0 $Y2=0
cc_875 N_A_1273_137#_c_1096_n N_A_978_67#_M1045_g 0.0114503f $X=7.125 $Y=2.16
+ $X2=0 $Y2=0
cc_876 N_A_1273_137#_c_1097_n N_A_978_67#_M1045_g 2.61615e-19 $X=7.21 $Y=2.075
+ $X2=0 $Y2=0
cc_877 N_A_1273_137#_c_1100_n N_A_978_67#_M1045_g 0.00384477f $X=6.585 $Y=2.16
+ $X2=0 $Y2=0
cc_878 N_A_1273_137#_M1033_g N_A_978_67#_c_1211_n 0.00969257f $X=8.905 $Y=2.315
+ $X2=0 $Y2=0
cc_879 N_A_1273_137#_M1029_g N_A_1840_21#_M1014_g 0.0285258f $X=8.725 $Y=0.785
+ $X2=0 $Y2=0
cc_880 N_A_1273_137#_M1029_g N_A_1840_21#_M1005_g 0.00193673f $X=8.725 $Y=0.785
+ $X2=0 $Y2=0
cc_881 N_A_1273_137#_c_1090_n N_A_1840_21#_M1005_g 3.70013e-19 $X=8.815 $Y=1.57
+ $X2=0 $Y2=0
cc_882 N_A_1273_137#_c_1091_n N_A_1840_21#_M1005_g 0.0781564f $X=8.815 $Y=1.57
+ $X2=0 $Y2=0
cc_883 N_A_1273_137#_c_1092_n N_VPWR_M1018_d 3.24744e-19 $X=7.92 $Y=1.56 $X2=0
+ $Y2=0
cc_884 N_A_1273_137#_M1033_g N_VPWR_c_1894_n 6.05222e-19 $X=8.905 $Y=2.315 $X2=0
+ $Y2=0
cc_885 N_A_1273_137#_c_1095_n N_VPWR_c_1909_n 0.00750623f $X=6.585 $Y=2.525
+ $X2=0 $Y2=0
cc_886 N_A_1273_137#_M1033_g N_VPWR_c_1889_n 9.39239e-19 $X=8.905 $Y=2.315 $X2=0
+ $Y2=0
cc_887 N_A_1273_137#_c_1095_n N_VPWR_c_1889_n 0.0102775f $X=6.585 $Y=2.525 $X2=0
+ $Y2=0
cc_888 N_A_1273_137#_c_1095_n N_A_202_119#_c_2087_n 0.00357659f $X=6.585
+ $Y=2.525 $X2=0 $Y2=0
cc_889 N_A_1273_137#_c_1100_n N_A_202_119#_c_2087_n 0.0135583f $X=6.585 $Y=2.16
+ $X2=0 $Y2=0
cc_890 N_A_1273_137#_c_1087_n N_A_202_119#_c_2088_n 0.0827729f $X=6.505 $Y=0.895
+ $X2=0 $Y2=0
cc_891 N_A_1273_137#_c_1095_n N_A_202_119#_c_2098_n 0.0186607f $X=6.585 $Y=2.525
+ $X2=0 $Y2=0
cc_892 N_A_1273_137#_c_1087_n N_VGND_c_2305_n 0.00319683f $X=6.505 $Y=0.895
+ $X2=0 $Y2=0
cc_893 N_A_1273_137#_M1029_g N_VGND_c_2311_n 7.85522e-19 $X=8.725 $Y=0.785 $X2=0
+ $Y2=0
cc_894 N_A_1273_137#_c_1087_n N_VGND_c_2322_n 0.00432875f $X=6.505 $Y=0.895
+ $X2=0 $Y2=0
cc_895 N_A_1273_137#_M1029_g N_A_1670_93#_c_2482_n 0.0109394f $X=8.725 $Y=0.785
+ $X2=0 $Y2=0
cc_896 N_A_1273_137#_c_1090_n N_A_1670_93#_c_2482_n 0.00113312f $X=8.815 $Y=1.57
+ $X2=0 $Y2=0
cc_897 N_A_1273_137#_M1029_g N_A_1670_93#_c_2483_n 0.00425749f $X=8.725 $Y=0.785
+ $X2=0 $Y2=0
cc_898 N_A_1273_137#_M1029_g N_A_1670_93#_c_2481_n 4.80356e-19 $X=8.725 $Y=0.785
+ $X2=0 $Y2=0
cc_899 N_A_978_67#_c_1201_n N_A_2415_137#_c_1329_n 0.021922f $X=11.76 $Y=1.31
+ $X2=0 $Y2=0
cc_900 N_A_978_67#_c_1199_n N_A_2415_137#_c_1341_n 0.021922f $X=11.685 $Y=1.385
+ $X2=0 $Y2=0
cc_901 N_A_978_67#_c_1201_n N_A_2211_428#_c_1563_n 0.00952769f $X=11.76 $Y=1.31
+ $X2=0 $Y2=0
cc_902 N_A_978_67#_M1020_g N_A_2211_428#_c_1542_n 0.0102077f $X=10.98 $Y=2.56
+ $X2=0 $Y2=0
cc_903 N_A_978_67#_c_1214_n N_A_2211_428#_c_1542_n 0.00997989f $X=11.33 $Y=1.99
+ $X2=0 $Y2=0
cc_904 N_A_978_67#_M1020_g N_A_2211_428#_c_1537_n 5.56793e-19 $X=10.98 $Y=2.56
+ $X2=0 $Y2=0
cc_905 N_A_978_67#_c_1214_n N_A_2211_428#_c_1537_n 0.0101706f $X=11.33 $Y=1.99
+ $X2=0 $Y2=0
cc_906 N_A_978_67#_c_1198_n N_A_2211_428#_c_1537_n 0.0197994f $X=11.405 $Y=1.915
+ $X2=0 $Y2=0
cc_907 N_A_978_67#_c_1200_n N_A_2211_428#_c_1537_n 0.0088094f $X=11.48 $Y=1.385
+ $X2=0 $Y2=0
cc_908 N_A_978_67#_c_1201_n N_A_2211_428#_c_1537_n 9.23128e-19 $X=11.76 $Y=1.31
+ $X2=0 $Y2=0
cc_909 N_A_978_67#_c_1200_n N_A_2211_428#_c_1538_n 0.00580376f $X=11.48 $Y=1.385
+ $X2=0 $Y2=0
cc_910 N_A_978_67#_c_1201_n N_A_2211_428#_c_1538_n 0.00652056f $X=11.76 $Y=1.31
+ $X2=0 $Y2=0
cc_911 N_A_978_67#_c_1211_n N_A_1840_21#_M1005_g 0.00988558f $X=10.905 $Y=3.15
+ $X2=0 $Y2=0
cc_912 N_A_978_67#_c_1201_n N_A_1840_21#_c_1627_n 0.0042225f $X=11.76 $Y=1.31
+ $X2=0 $Y2=0
cc_913 N_A_978_67#_c_1211_n N_VPWR_c_1894_n 0.0256338f $X=10.905 $Y=3.15 $X2=0
+ $Y2=0
cc_914 N_A_978_67#_c_1211_n N_VPWR_c_1895_n 0.0261591f $X=10.905 $Y=3.15 $X2=0
+ $Y2=0
cc_915 N_A_978_67#_c_1212_n N_VPWR_c_1909_n 0.0440016f $X=6.875 $Y=3.15 $X2=0
+ $Y2=0
cc_916 N_A_978_67#_c_1211_n N_VPWR_c_1911_n 0.0341141f $X=10.905 $Y=3.15 $X2=0
+ $Y2=0
cc_917 N_A_978_67#_c_1211_n N_VPWR_c_1914_n 0.0381055f $X=10.905 $Y=3.15 $X2=0
+ $Y2=0
cc_918 N_A_978_67#_c_1211_n N_VPWR_c_1889_n 0.149421f $X=10.905 $Y=3.15 $X2=0
+ $Y2=0
cc_919 N_A_978_67#_c_1212_n N_VPWR_c_1889_n 0.00968212f $X=6.875 $Y=3.15 $X2=0
+ $Y2=0
cc_920 N_A_978_67#_M1008_s N_A_202_119#_c_2093_n 0.0053174f $X=4.905 $Y=1.835
+ $X2=0 $Y2=0
cc_921 N_A_978_67#_M1008_s N_A_202_119#_c_2147_n 0.0120156f $X=4.905 $Y=1.835
+ $X2=0 $Y2=0
cc_922 N_A_978_67#_M1008_s N_A_202_119#_c_2148_n 0.00419556f $X=4.905 $Y=1.835
+ $X2=0 $Y2=0
cc_923 N_A_978_67#_c_1202_n N_A_202_119#_c_2148_n 0.0147539f $X=5.075 $Y=1.815
+ $X2=0 $Y2=0
cc_924 N_A_978_67#_c_1206_n N_A_202_119#_c_2087_n 0.00834753f $X=6.215 $Y=1.87
+ $X2=0 $Y2=0
cc_925 N_A_978_67#_c_1207_n N_A_202_119#_c_2087_n 9.50286e-19 $X=5.945 $Y=1.87
+ $X2=0 $Y2=0
cc_926 N_A_978_67#_M1011_g N_A_202_119#_c_2087_n 0.0137378f $X=6.29 $Y=0.895
+ $X2=0 $Y2=0
cc_927 N_A_978_67#_M1045_g N_A_202_119#_c_2087_n 4.839e-19 $X=6.8 $Y=2.525 $X2=0
+ $Y2=0
cc_928 N_A_978_67#_c_1217_n N_A_202_119#_c_2087_n 0.00270391f $X=6.29 $Y=1.87
+ $X2=0 $Y2=0
cc_929 N_A_978_67#_c_1219_n N_A_202_119#_c_2087_n 0.0125169f $X=5.615 $Y=1.9
+ $X2=0 $Y2=0
cc_930 N_A_978_67#_c_1203_n N_A_202_119#_c_2087_n 0.0353525f $X=5.78 $Y=1.48
+ $X2=0 $Y2=0
cc_931 N_A_978_67#_c_1204_n N_A_202_119#_c_2087_n 0.0032415f $X=5.78 $Y=1.48
+ $X2=0 $Y2=0
cc_932 N_A_978_67#_c_1206_n N_A_202_119#_c_2088_n 8.10252e-19 $X=6.215 $Y=1.87
+ $X2=0 $Y2=0
cc_933 N_A_978_67#_M1011_g N_A_202_119#_c_2088_n 0.00653517f $X=6.29 $Y=0.895
+ $X2=0 $Y2=0
cc_934 N_A_978_67#_c_1204_n N_A_202_119#_c_2088_n 0.00151867f $X=5.78 $Y=1.48
+ $X2=0 $Y2=0
cc_935 N_A_978_67#_c_1207_n N_A_202_119#_c_2097_n 0.00232728f $X=5.945 $Y=1.87
+ $X2=0 $Y2=0
cc_936 N_A_978_67#_c_1202_n N_A_202_119#_c_2097_n 0.0015858f $X=5.075 $Y=1.815
+ $X2=0 $Y2=0
cc_937 N_A_978_67#_c_1219_n N_A_202_119#_c_2097_n 0.0311744f $X=5.615 $Y=1.9
+ $X2=0 $Y2=0
cc_938 N_A_978_67#_c_1206_n N_A_202_119#_c_2098_n 0.00498028f $X=6.215 $Y=1.87
+ $X2=0 $Y2=0
cc_939 N_A_978_67#_c_1207_n N_A_202_119#_c_2098_n 0.00137355f $X=5.945 $Y=1.87
+ $X2=0 $Y2=0
cc_940 N_A_978_67#_M1011_g N_VGND_c_2294_n 0.00312944f $X=6.29 $Y=0.895 $X2=0
+ $Y2=0
cc_941 N_A_978_67#_c_1203_n N_VGND_c_2294_n 0.00345613f $X=5.78 $Y=1.48 $X2=0
+ $Y2=0
cc_942 N_A_978_67#_c_1204_n N_VGND_c_2294_n 6.04595e-19 $X=5.78 $Y=1.48 $X2=0
+ $Y2=0
cc_943 N_A_978_67#_c_1205_n N_VGND_c_2294_n 0.0180054f $X=5.035 $Y=0.545 $X2=0
+ $Y2=0
cc_944 N_A_978_67#_c_1205_n N_VGND_c_2310_n 0.0169023f $X=5.035 $Y=0.545 $X2=0
+ $Y2=0
cc_945 N_A_978_67#_M1011_g N_VGND_c_2322_n 9.58071e-19 $X=6.29 $Y=0.895 $X2=0
+ $Y2=0
cc_946 N_A_978_67#_c_1201_n N_VGND_c_2322_n 9.72468e-19 $X=11.76 $Y=1.31 $X2=0
+ $Y2=0
cc_947 N_A_978_67#_c_1205_n N_VGND_c_2322_n 0.0123275f $X=5.035 $Y=0.545 $X2=0
+ $Y2=0
cc_948 N_A_2415_137#_c_1344_n N_A_2211_428#_M1047_g 0.00230031f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_949 N_A_2415_137#_c_1397_p N_A_2211_428#_M1000_g 0.011778f $X=13.665 $Y=2.475
+ $X2=0 $Y2=0
cc_950 N_A_2415_137#_c_1362_n N_A_2211_428#_M1000_g 0.00595172f $X=13.28
+ $Y=2.205 $X2=0 $Y2=0
cc_951 N_A_2415_137#_c_1392_n N_A_2211_428#_M1000_g 0.0100578f $X=13.28 $Y=2.475
+ $X2=0 $Y2=0
cc_952 N_A_2415_137#_c_1329_n N_A_2211_428#_c_1563_n 0.0107445f $X=12.15 $Y=1.31
+ $X2=0 $Y2=0
cc_953 N_A_2415_137#_c_1341_n N_A_2211_428#_c_1563_n 0.0034285f $X=12.305
+ $Y=1.385 $X2=0 $Y2=0
cc_954 N_A_2415_137#_c_1344_n N_A_2211_428#_c_1536_n 0.0113598f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_955 N_A_2415_137#_c_1341_n N_A_2211_428#_c_1537_n 6.08269e-19 $X=12.305
+ $Y=1.385 $X2=0 $Y2=0
cc_956 N_A_2415_137#_c_1397_p N_A_2211_428#_c_1539_n 0.0010066f $X=13.665
+ $Y=2.475 $X2=0 $Y2=0
cc_957 N_A_2415_137#_c_1344_n N_A_2211_428#_c_1539_n 0.0238515f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_958 N_A_2415_137#_c_1362_n N_A_2211_428#_c_1539_n 0.0161408f $X=13.28
+ $Y=2.205 $X2=0 $Y2=0
cc_959 N_A_2415_137#_c_1344_n N_A_2211_428#_c_1540_n 0.0114194f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_960 N_A_2415_137#_c_1362_n N_A_2211_428#_c_1540_n 0.00587513f $X=13.28
+ $Y=2.205 $X2=0 $Y2=0
cc_961 N_A_2415_137#_c_1409_p N_A_2211_428#_c_1540_n 0.00293878f $X=13.657
+ $Y=1.165 $X2=0 $Y2=0
cc_962 N_A_2415_137#_c_1358_n N_A_1840_21#_M1040_s 0.00274313f $X=15.135
+ $Y=2.475 $X2=0 $Y2=0
cc_963 N_A_2415_137#_c_1329_n N_A_1840_21#_c_1627_n 0.0042225f $X=12.15 $Y=1.31
+ $X2=0 $Y2=0
cc_964 N_A_2415_137#_c_1412_p N_A_1840_21#_M1031_g 0.00655523f $X=13.645
+ $Y=0.815 $X2=0 $Y2=0
cc_965 N_A_2415_137#_c_1409_p N_A_1840_21#_M1031_g 0.00240289f $X=13.657
+ $Y=1.165 $X2=0 $Y2=0
cc_966 N_A_2415_137#_c_1344_n N_A_1840_21#_M1026_g 0.0111794f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_967 N_A_2415_137#_c_1358_n N_A_1840_21#_M1026_g 0.0140219f $X=15.135 $Y=2.475
+ $X2=0 $Y2=0
cc_968 N_A_2415_137#_c_1362_n N_A_1840_21#_M1026_g 3.09787e-19 $X=13.28 $Y=2.205
+ $X2=0 $Y2=0
cc_969 N_A_2415_137#_c_1392_n N_A_1840_21#_M1026_g 0.00180922f $X=13.28 $Y=2.475
+ $X2=0 $Y2=0
cc_970 N_A_2415_137#_c_1418_p N_A_1840_21#_M1026_g 0.00274355f $X=13.75 $Y=2.475
+ $X2=0 $Y2=0
cc_971 N_A_2415_137#_c_1344_n N_A_1840_21#_c_1631_n 0.0017618f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_972 N_A_2415_137#_c_1409_p N_A_1840_21#_c_1631_n 0.00235737f $X=13.657
+ $Y=1.165 $X2=0 $Y2=0
cc_973 N_A_2415_137#_M1012_g N_A_1840_21#_c_1632_n 2.97301e-19 $X=15.36 $Y=0.685
+ $X2=0 $Y2=0
cc_974 N_A_2415_137#_c_1412_p N_A_1840_21#_c_1632_n 0.00507539f $X=13.645
+ $Y=0.815 $X2=0 $Y2=0
cc_975 N_A_2415_137#_c_1409_p N_A_1840_21#_c_1632_n 0.0137627f $X=13.657
+ $Y=1.165 $X2=0 $Y2=0
cc_976 N_A_2415_137#_c_1344_n N_A_1840_21#_c_1633_n 0.0548532f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_977 N_A_2415_137#_c_1344_n N_A_1840_21#_c_1634_n 0.0153812f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_978 N_A_2415_137#_c_1358_n N_A_1840_21#_c_1634_n 0.00151208f $X=15.135
+ $Y=2.475 $X2=0 $Y2=0
cc_979 N_A_2415_137#_c_1344_n N_A_1840_21#_c_1639_n 0.0189019f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_980 N_A_2415_137#_c_1358_n N_A_1840_21#_c_1639_n 0.0259973f $X=15.135
+ $Y=2.475 $X2=0 $Y2=0
cc_981 N_A_2415_137#_M1001_g N_A_1840_21#_c_1640_n 2.21268e-19 $X=15.355
+ $Y=2.465 $X2=0 $Y2=0
cc_982 N_A_2415_137#_c_1358_n N_A_1840_21#_c_1640_n 0.0287848f $X=15.135
+ $Y=2.475 $X2=0 $Y2=0
cc_983 N_A_2415_137#_c_1345_n N_A_1840_21#_c_1640_n 0.0114001f $X=15.22 $Y=2.39
+ $X2=0 $Y2=0
cc_984 N_A_2415_137#_c_1344_n N_A_1840_21#_c_1635_n 0.00302954f $X=13.75 $Y=2.39
+ $X2=0 $Y2=0
cc_985 N_A_2415_137#_M1001_g N_RESET_B_c_1735_n 0.0289957f $X=15.355 $Y=2.465
+ $X2=-0.19 $Y2=-0.245
cc_986 N_A_2415_137#_c_1345_n N_RESET_B_c_1735_n 0.0101664f $X=15.22 $Y=2.39
+ $X2=-0.19 $Y2=-0.245
cc_987 N_A_2415_137#_c_1346_n N_RESET_B_c_1735_n 8.40516e-19 $X=15.33 $Y=1.47
+ $X2=-0.19 $Y2=-0.245
cc_988 N_A_2415_137#_c_1348_n N_RESET_B_c_1735_n 0.00725117f $X=15.33 $Y=1.38
+ $X2=-0.19 $Y2=-0.245
cc_989 N_A_2415_137#_c_1358_n N_RESET_B_M1040_g 0.0153965f $X=15.135 $Y=2.475
+ $X2=0 $Y2=0
cc_990 N_A_2415_137#_M1012_g N_RESET_B_M1032_g 0.0156028f $X=15.36 $Y=0.685
+ $X2=0 $Y2=0
cc_991 N_A_2415_137#_c_1346_n N_RESET_B_M1032_g 0.00173926f $X=15.33 $Y=1.47
+ $X2=0 $Y2=0
cc_992 N_A_2415_137#_c_1348_n N_RESET_B_M1032_g 0.00999942f $X=15.33 $Y=1.38
+ $X2=0 $Y2=0
cc_993 N_A_2415_137#_c_1358_n N_RESET_B_c_1737_n 0.00314888f $X=15.135 $Y=2.475
+ $X2=0 $Y2=0
cc_994 N_A_2415_137#_c_1345_n N_RESET_B_c_1737_n 0.00923197f $X=15.22 $Y=2.39
+ $X2=0 $Y2=0
cc_995 N_A_2415_137#_c_1346_n N_RESET_B_c_1737_n 0.0192671f $X=15.33 $Y=1.47
+ $X2=0 $Y2=0
cc_996 N_A_2415_137#_c_1348_n N_RESET_B_c_1737_n 3.45351e-19 $X=15.33 $Y=1.38
+ $X2=0 $Y2=0
cc_997 N_A_2415_137#_M1038_g N_A_3289_47#_c_1773_n 0.0148332f $X=16.805 $Y=0.445
+ $X2=0 $Y2=0
cc_998 N_A_2415_137#_c_1353_n N_A_3289_47#_M1002_g 0.0160189f $X=16.73 $Y=1.83
+ $X2=0 $Y2=0
cc_999 N_A_2415_137#_M1041_g N_A_3289_47#_c_1779_n 2.82754e-19 $X=15.79 $Y=0.685
+ $X2=0 $Y2=0
cc_1000 N_A_2415_137#_c_1336_n N_A_3289_47#_c_1779_n 0.00401296f $X=16.325
+ $Y=1.305 $X2=0 $Y2=0
cc_1001 N_A_2415_137#_c_1338_n N_A_3289_47#_c_1779_n 0.0222048f $X=16.73 $Y=0.87
+ $X2=0 $Y2=0
cc_1002 N_A_2415_137#_M1038_g N_A_3289_47#_c_1779_n 0.00858557f $X=16.805
+ $Y=0.445 $X2=0 $Y2=0
cc_1003 N_A_2415_137#_M1024_g N_A_3289_47#_c_1780_n 0.00110512f $X=15.785
+ $Y=2.465 $X2=0 $Y2=0
cc_1004 N_A_2415_137#_c_1337_n N_A_3289_47#_c_1780_n 0.00457381f $X=16.325
+ $Y=1.755 $X2=0 $Y2=0
cc_1005 N_A_2415_137#_c_1353_n N_A_3289_47#_c_1780_n 0.0237048f $X=16.73 $Y=1.83
+ $X2=0 $Y2=0
cc_1006 N_A_2415_137#_c_1355_n N_A_3289_47#_c_1780_n 0.00997626f $X=16.805
+ $Y=1.905 $X2=0 $Y2=0
cc_1007 N_A_2415_137#_c_1338_n N_A_3289_47#_c_1781_n 0.00512525f $X=16.73
+ $Y=0.87 $X2=0 $Y2=0
cc_1008 N_A_2415_137#_c_1353_n N_A_3289_47#_c_1781_n 0.00512525f $X=16.73
+ $Y=1.83 $X2=0 $Y2=0
cc_1009 N_A_2415_137#_c_1336_n N_A_3289_47#_c_1782_n 0.00727134f $X=16.325
+ $Y=1.305 $X2=0 $Y2=0
cc_1010 N_A_2415_137#_c_1336_n N_A_3289_47#_c_1783_n 0.00520866f $X=16.325
+ $Y=1.305 $X2=0 $Y2=0
cc_1011 N_A_2415_137#_c_1356_n N_VPWR_M1035_d 0.00231921f $X=13.115 $Y=2.205
+ $X2=0 $Y2=0
cc_1012 N_A_2415_137#_c_1358_n N_VPWR_M1026_d 0.00505472f $X=15.135 $Y=2.475
+ $X2=0 $Y2=0
cc_1013 N_A_2415_137#_c_1358_n N_VPWR_M1040_d 0.00843932f $X=15.135 $Y=2.475
+ $X2=0 $Y2=0
cc_1014 N_A_2415_137#_c_1345_n N_VPWR_M1040_d 0.00647076f $X=15.22 $Y=2.39 $X2=0
+ $Y2=0
cc_1015 N_A_2415_137#_M1035_g N_VPWR_c_1896_n 0.00718839f $X=12.335 $Y=2.74
+ $X2=0 $Y2=0
cc_1016 N_A_2415_137#_c_1356_n N_VPWR_c_1896_n 0.0193616f $X=13.115 $Y=2.205
+ $X2=0 $Y2=0
cc_1017 N_A_2415_137#_c_1358_n N_VPWR_c_1897_n 0.0203541f $X=15.135 $Y=2.475
+ $X2=0 $Y2=0
cc_1018 N_A_2415_137#_c_1392_n N_VPWR_c_1897_n 0.0102962f $X=13.28 $Y=2.475
+ $X2=0 $Y2=0
cc_1019 N_A_2415_137#_M1001_g N_VPWR_c_1898_n 0.00918181f $X=15.355 $Y=2.465
+ $X2=0 $Y2=0
cc_1020 N_A_2415_137#_M1024_g N_VPWR_c_1898_n 5.02705e-19 $X=15.785 $Y=2.465
+ $X2=0 $Y2=0
cc_1021 N_A_2415_137#_c_1358_n N_VPWR_c_1898_n 0.021106f $X=15.135 $Y=2.475
+ $X2=0 $Y2=0
cc_1022 N_A_2415_137#_M1024_g N_VPWR_c_1899_n 0.0105759f $X=15.785 $Y=2.465
+ $X2=0 $Y2=0
cc_1023 N_A_2415_137#_c_1335_n N_VPWR_c_1899_n 0.00708393f $X=16.25 $Y=1.38
+ $X2=0 $Y2=0
cc_1024 N_A_2415_137#_c_1354_n N_VPWR_c_1899_n 0.00105805f $X=16.4 $Y=1.83 $X2=0
+ $Y2=0
cc_1025 N_A_2415_137#_c_1355_n N_VPWR_c_1899_n 0.0040956f $X=16.805 $Y=1.905
+ $X2=0 $Y2=0
cc_1026 N_A_2415_137#_c_1353_n N_VPWR_c_1900_n 0.00801714f $X=16.73 $Y=1.83
+ $X2=0 $Y2=0
cc_1027 N_A_2415_137#_M1035_g N_VPWR_c_1914_n 0.00570944f $X=12.335 $Y=2.74
+ $X2=0 $Y2=0
cc_1028 N_A_2415_137#_c_1392_n N_VPWR_c_1915_n 0.0177952f $X=13.28 $Y=2.475
+ $X2=0 $Y2=0
cc_1029 N_A_2415_137#_M1001_g N_VPWR_c_1917_n 0.00486043f $X=15.355 $Y=2.465
+ $X2=0 $Y2=0
cc_1030 N_A_2415_137#_M1024_g N_VPWR_c_1917_n 0.00504158f $X=15.785 $Y=2.465
+ $X2=0 $Y2=0
cc_1031 N_A_2415_137#_c_1355_n N_VPWR_c_1918_n 0.00360349f $X=16.805 $Y=1.905
+ $X2=0 $Y2=0
cc_1032 N_A_2415_137#_M1023_d N_VPWR_c_1889_n 0.00223819f $X=13.14 $Y=2.255
+ $X2=0 $Y2=0
cc_1033 N_A_2415_137#_M1035_g N_VPWR_c_1889_n 0.00542671f $X=12.335 $Y=2.74
+ $X2=0 $Y2=0
cc_1034 N_A_2415_137#_M1001_g N_VPWR_c_1889_n 0.00824727f $X=15.355 $Y=2.465
+ $X2=0 $Y2=0
cc_1035 N_A_2415_137#_M1024_g N_VPWR_c_1889_n 0.0100635f $X=15.785 $Y=2.465
+ $X2=0 $Y2=0
cc_1036 N_A_2415_137#_c_1355_n N_VPWR_c_1889_n 0.00446563f $X=16.805 $Y=1.905
+ $X2=0 $Y2=0
cc_1037 N_A_2415_137#_c_1397_p N_VPWR_c_1889_n 0.00716124f $X=13.665 $Y=2.475
+ $X2=0 $Y2=0
cc_1038 N_A_2415_137#_c_1358_n N_VPWR_c_1889_n 0.0310731f $X=15.135 $Y=2.475
+ $X2=0 $Y2=0
cc_1039 N_A_2415_137#_c_1392_n N_VPWR_c_1889_n 0.0123247f $X=13.28 $Y=2.475
+ $X2=0 $Y2=0
cc_1040 N_A_2415_137#_c_1418_p N_VPWR_c_1889_n 0.00689755f $X=13.75 $Y=2.475
+ $X2=0 $Y2=0
cc_1041 N_A_2415_137#_c_1397_p A_2714_451# 0.00211059f $X=13.665 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1042 N_A_2415_137#_c_1344_n A_2714_451# 9.95692e-19 $X=13.75 $Y=2.39
+ $X2=-0.19 $Y2=-0.245
cc_1043 N_A_2415_137#_c_1418_p A_2714_451# 0.0019409f $X=13.75 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1044 N_A_2415_137#_M1012_g N_Q_N_c_2231_n 0.00914485f $X=15.36 $Y=0.685 $X2=0
+ $Y2=0
cc_1045 N_A_2415_137#_M1041_g N_Q_N_c_2231_n 0.0106208f $X=15.79 $Y=0.685 $X2=0
+ $Y2=0
cc_1046 N_A_2415_137#_c_1336_n N_Q_N_c_2231_n 6.66365e-19 $X=16.325 $Y=1.305
+ $X2=0 $Y2=0
cc_1047 N_A_2415_137#_M1012_g N_Q_N_c_2232_n 0.00331259f $X=15.36 $Y=0.685 $X2=0
+ $Y2=0
cc_1048 N_A_2415_137#_c_1332_n N_Q_N_c_2232_n 0.00284666f $X=15.71 $Y=1.38 $X2=0
+ $Y2=0
cc_1049 N_A_2415_137#_M1041_g N_Q_N_c_2232_n 0.00238778f $X=15.79 $Y=0.685 $X2=0
+ $Y2=0
cc_1050 N_A_2415_137#_M1001_g Q_N 7.35776e-19 $X=15.355 $Y=2.465 $X2=0 $Y2=0
cc_1051 N_A_2415_137#_c_1332_n Q_N 0.00351777f $X=15.71 $Y=1.38 $X2=0 $Y2=0
cc_1052 N_A_2415_137#_M1024_g Q_N 0.00194945f $X=15.785 $Y=2.465 $X2=0 $Y2=0
cc_1053 N_A_2415_137#_c_1354_n Q_N 6.82447e-19 $X=16.4 $Y=1.83 $X2=0 $Y2=0
cc_1054 N_A_2415_137#_c_1345_n Q_N 0.019322f $X=15.22 $Y=2.39 $X2=0 $Y2=0
cc_1055 N_A_2415_137#_c_1348_n Q_N 4.30792e-19 $X=15.33 $Y=1.38 $X2=0 $Y2=0
cc_1056 N_A_2415_137#_M1024_g Q_N 0.0161105f $X=15.785 $Y=2.465 $X2=0 $Y2=0
cc_1057 N_A_2415_137#_M1001_g N_Q_N_c_2233_n 9.02127e-19 $X=15.355 $Y=2.465
+ $X2=0 $Y2=0
cc_1058 N_A_2415_137#_M1012_g N_Q_N_c_2233_n 0.00271801f $X=15.36 $Y=0.685 $X2=0
+ $Y2=0
cc_1059 N_A_2415_137#_c_1332_n N_Q_N_c_2233_n 0.00714577f $X=15.71 $Y=1.38 $X2=0
+ $Y2=0
cc_1060 N_A_2415_137#_M1024_g N_Q_N_c_2233_n 0.0102282f $X=15.785 $Y=2.465 $X2=0
+ $Y2=0
cc_1061 N_A_2415_137#_M1041_g N_Q_N_c_2233_n 0.00531894f $X=15.79 $Y=0.685 $X2=0
+ $Y2=0
cc_1062 N_A_2415_137#_c_1337_n N_Q_N_c_2233_n 6.82447e-19 $X=16.325 $Y=1.755
+ $X2=0 $Y2=0
cc_1063 N_A_2415_137#_c_1342_n N_Q_N_c_2233_n 0.00476979f $X=15.787 $Y=1.38
+ $X2=0 $Y2=0
cc_1064 N_A_2415_137#_c_1345_n N_Q_N_c_2233_n 0.00622568f $X=15.22 $Y=2.39 $X2=0
+ $Y2=0
cc_1065 N_A_2415_137#_c_1346_n N_Q_N_c_2233_n 0.0228669f $X=15.33 $Y=1.47 $X2=0
+ $Y2=0
cc_1066 N_A_2415_137#_c_1348_n N_Q_N_c_2233_n 0.00113483f $X=15.33 $Y=1.38 $X2=0
+ $Y2=0
cc_1067 N_A_2415_137#_c_1353_n N_Q_c_2270_n 4.66768e-19 $X=16.73 $Y=1.83 $X2=0
+ $Y2=0
cc_1068 N_A_2415_137#_M1012_g N_VGND_c_2298_n 0.0055345f $X=15.36 $Y=0.685 $X2=0
+ $Y2=0
cc_1069 N_A_2415_137#_c_1346_n N_VGND_c_2298_n 0.00771837f $X=15.33 $Y=1.47
+ $X2=0 $Y2=0
cc_1070 N_A_2415_137#_c_1348_n N_VGND_c_2298_n 0.00148357f $X=15.33 $Y=1.38
+ $X2=0 $Y2=0
cc_1071 N_A_2415_137#_M1041_g N_VGND_c_2299_n 0.0100682f $X=15.79 $Y=0.685 $X2=0
+ $Y2=0
cc_1072 N_A_2415_137#_c_1335_n N_VGND_c_2299_n 0.00833665f $X=16.25 $Y=1.38
+ $X2=0 $Y2=0
cc_1073 N_A_2415_137#_c_1339_n N_VGND_c_2299_n 0.00367244f $X=16.4 $Y=0.87 $X2=0
+ $Y2=0
cc_1074 N_A_2415_137#_M1038_g N_VGND_c_2299_n 0.00389969f $X=16.805 $Y=0.445
+ $X2=0 $Y2=0
cc_1075 N_A_2415_137#_M1038_g N_VGND_c_2300_n 0.00787301f $X=16.805 $Y=0.445
+ $X2=0 $Y2=0
cc_1076 N_A_2415_137#_M1012_g N_VGND_c_2313_n 0.00520813f $X=15.36 $Y=0.685
+ $X2=0 $Y2=0
cc_1077 N_A_2415_137#_M1041_g N_VGND_c_2313_n 0.00484947f $X=15.79 $Y=0.685
+ $X2=0 $Y2=0
cc_1078 N_A_2415_137#_M1038_g N_VGND_c_2314_n 0.00550269f $X=16.805 $Y=0.445
+ $X2=0 $Y2=0
cc_1079 N_A_2415_137#_c_1329_n N_VGND_c_2322_n 9.72468e-19 $X=12.15 $Y=1.31
+ $X2=0 $Y2=0
cc_1080 N_A_2415_137#_M1012_g N_VGND_c_2322_n 0.0107404f $X=15.36 $Y=0.685 $X2=0
+ $Y2=0
cc_1081 N_A_2415_137#_M1041_g N_VGND_c_2322_n 0.00988247f $X=15.79 $Y=0.685
+ $X2=0 $Y2=0
cc_1082 N_A_2415_137#_c_1339_n N_VGND_c_2322_n 0.00447465f $X=16.4 $Y=0.87 $X2=0
+ $Y2=0
cc_1083 N_A_2415_137#_M1038_g N_VGND_c_2322_n 0.0115948f $X=16.805 $Y=0.445
+ $X2=0 $Y2=0
cc_1084 N_A_2415_137#_M1047_d N_A_2574_119#_c_2507_n 0.00240753f $X=13.46
+ $Y=0.595 $X2=0 $Y2=0
cc_1085 N_A_2415_137#_c_1412_p N_A_2574_119#_c_2507_n 0.018109f $X=13.645
+ $Y=0.815 $X2=0 $Y2=0
cc_1086 N_A_2415_137#_c_1409_p N_A_2574_119#_c_2507_n 6.83881e-19 $X=13.657
+ $Y=1.165 $X2=0 $Y2=0
cc_1087 N_A_2211_428#_M1047_g N_A_1840_21#_c_1627_n 0.00881852f $X=13.385
+ $Y=0.915 $X2=0 $Y2=0
cc_1088 N_A_2211_428#_c_1563_n N_A_1840_21#_c_1627_n 0.00982857f $X=13.13
+ $Y=0.915 $X2=0 $Y2=0
cc_1089 N_A_2211_428#_c_1538_n N_A_1840_21#_c_1627_n 0.00665063f $X=11.465
+ $Y=0.74 $X2=0 $Y2=0
cc_1090 N_A_2211_428#_M1047_g N_A_1840_21#_M1031_g 0.0125982f $X=13.385 $Y=0.915
+ $X2=0 $Y2=0
cc_1091 N_A_2211_428#_M1000_g N_A_1840_21#_M1026_g 0.0455532f $X=13.495 $Y=2.675
+ $X2=0 $Y2=0
cc_1092 N_A_2211_428#_c_1539_n N_A_1840_21#_c_1634_n 2.79993e-19 $X=13.325
+ $Y=1.625 $X2=0 $Y2=0
cc_1093 N_A_2211_428#_c_1540_n N_A_1840_21#_c_1634_n 0.0455532f $X=13.325
+ $Y=1.625 $X2=0 $Y2=0
cc_1094 N_A_2211_428#_M1047_g N_A_1840_21#_c_1635_n 0.00719057f $X=13.385
+ $Y=0.915 $X2=0 $Y2=0
cc_1095 N_A_2211_428#_M1000_g N_VPWR_c_1897_n 0.00215642f $X=13.495 $Y=2.675
+ $X2=0 $Y2=0
cc_1096 N_A_2211_428#_M1000_g N_VPWR_c_1915_n 0.00549284f $X=13.495 $Y=2.675
+ $X2=0 $Y2=0
cc_1097 N_A_2211_428#_M1000_g N_VPWR_c_1889_n 0.00606697f $X=13.495 $Y=2.675
+ $X2=0 $Y2=0
cc_1098 N_A_2211_428#_c_1563_n N_VGND_M1037_d 0.00893372f $X=13.13 $Y=0.915
+ $X2=0 $Y2=0
cc_1099 N_A_2211_428#_c_1563_n N_VGND_c_2297_n 0.0239225f $X=13.13 $Y=0.915
+ $X2=0 $Y2=0
cc_1100 N_A_2211_428#_c_1538_n N_VGND_c_2307_n 0.00755126f $X=11.465 $Y=0.74
+ $X2=0 $Y2=0
cc_1101 N_A_2211_428#_c_1563_n N_VGND_c_2322_n 0.0303859f $X=13.13 $Y=0.915
+ $X2=0 $Y2=0
cc_1102 N_A_2211_428#_c_1538_n N_VGND_c_2322_n 0.00910022f $X=11.465 $Y=0.74
+ $X2=0 $Y2=0
cc_1103 N_A_2211_428#_c_1563_n A_2367_163# 0.002809f $X=13.13 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_1104 N_A_2211_428#_c_1563_n N_A_2574_119#_M1030_d 0.0121238f $X=13.13
+ $Y=0.915 $X2=-0.19 $Y2=-0.245
cc_1105 N_A_2211_428#_c_1536_n N_A_2574_119#_M1030_d 0.00425707f $X=13.215
+ $Y=1.46 $X2=-0.19 $Y2=-0.245
cc_1106 N_A_2211_428#_M1047_g N_A_2574_119#_c_2507_n 0.00376655f $X=13.385
+ $Y=0.915 $X2=0 $Y2=0
cc_1107 N_A_2211_428#_M1047_g N_A_2574_119#_c_2509_n 0.0040979f $X=13.385
+ $Y=0.915 $X2=0 $Y2=0
cc_1108 N_A_2211_428#_c_1563_n N_A_2574_119#_c_2509_n 0.024484f $X=13.13
+ $Y=0.915 $X2=0 $Y2=0
cc_1109 N_A_1840_21#_c_1632_n N_RESET_B_c_1735_n 0.00140661f $X=14.177 $Y=1.165
+ $X2=-0.19 $Y2=-0.245
cc_1110 N_A_1840_21#_c_1633_n N_RESET_B_c_1735_n 4.51847e-19 $X=14.175 $Y=1.54
+ $X2=-0.19 $Y2=-0.245
cc_1111 N_A_1840_21#_c_1634_n N_RESET_B_c_1735_n 0.0155674f $X=14.175 $Y=1.54
+ $X2=-0.19 $Y2=-0.245
cc_1112 N_A_1840_21#_c_1640_n N_RESET_B_c_1735_n 8.80366e-19 $X=14.63 $Y=2.125
+ $X2=-0.19 $Y2=-0.245
cc_1113 N_A_1840_21#_c_1635_n N_RESET_B_c_1735_n 3.25854e-19 $X=14.075 $Y=1.375
+ $X2=-0.19 $Y2=-0.245
cc_1114 N_A_1840_21#_c_1633_n N_RESET_B_M1040_g 0.00101375f $X=14.175 $Y=1.54
+ $X2=0 $Y2=0
cc_1115 N_A_1840_21#_c_1634_n N_RESET_B_M1040_g 0.00901722f $X=14.175 $Y=1.54
+ $X2=0 $Y2=0
cc_1116 N_A_1840_21#_c_1640_n N_RESET_B_M1040_g 0.00420437f $X=14.63 $Y=2.125
+ $X2=0 $Y2=0
cc_1117 N_A_1840_21#_c_1632_n N_RESET_B_M1032_g 0.00900047f $X=14.177 $Y=1.165
+ $X2=0 $Y2=0
cc_1118 N_A_1840_21#_c_1633_n N_RESET_B_M1032_g 0.00501084f $X=14.175 $Y=1.54
+ $X2=0 $Y2=0
cc_1119 N_A_1840_21#_c_1632_n N_RESET_B_c_1737_n 0.0222728f $X=14.177 $Y=1.165
+ $X2=0 $Y2=0
cc_1120 N_A_1840_21#_c_1633_n N_RESET_B_c_1737_n 0.0328683f $X=14.175 $Y=1.54
+ $X2=0 $Y2=0
cc_1121 N_A_1840_21#_c_1634_n N_RESET_B_c_1737_n 0.00296355f $X=14.175 $Y=1.54
+ $X2=0 $Y2=0
cc_1122 N_A_1840_21#_c_1640_n N_RESET_B_c_1737_n 0.0189127f $X=14.63 $Y=2.125
+ $X2=0 $Y2=0
cc_1123 N_A_1840_21#_M1005_g N_VPWR_c_1895_n 0.0221195f $X=9.295 $Y=2.315 $X2=0
+ $Y2=0
cc_1124 N_A_1840_21#_M1026_g N_VPWR_c_1897_n 0.0121417f $X=13.885 $Y=2.675 $X2=0
+ $Y2=0
cc_1125 N_A_1840_21#_M1026_g N_VPWR_c_1915_n 0.00486043f $X=13.885 $Y=2.675
+ $X2=0 $Y2=0
cc_1126 N_A_1840_21#_M1005_g N_VPWR_c_1889_n 9.39239e-19 $X=9.295 $Y=2.315 $X2=0
+ $Y2=0
cc_1127 N_A_1840_21#_M1026_g N_VPWR_c_1889_n 0.00439071f $X=13.885 $Y=2.675
+ $X2=0 $Y2=0
cc_1128 N_A_1840_21#_c_1627_n N_VGND_c_2296_n 0.021158f $X=13.785 $Y=0.18 $X2=0
+ $Y2=0
cc_1129 N_A_1840_21#_c_1627_n N_VGND_c_2297_n 0.0252872f $X=13.785 $Y=0.18 $X2=0
+ $Y2=0
cc_1130 N_A_1840_21#_c_1632_n N_VGND_c_2298_n 0.0185826f $X=14.177 $Y=1.165
+ $X2=0 $Y2=0
cc_1131 N_A_1840_21#_c_1627_n N_VGND_c_2307_n 0.0626184f $X=13.785 $Y=0.18 $X2=0
+ $Y2=0
cc_1132 N_A_1840_21#_c_1628_n N_VGND_c_2311_n 0.0239302f $X=9.35 $Y=0.18 $X2=0
+ $Y2=0
cc_1133 N_A_1840_21#_c_1627_n N_VGND_c_2312_n 0.0305321f $X=13.785 $Y=0.18 $X2=0
+ $Y2=0
cc_1134 N_A_1840_21#_c_1632_n N_VGND_c_2312_n 0.0060842f $X=14.177 $Y=1.165
+ $X2=0 $Y2=0
cc_1135 N_A_1840_21#_c_1627_n N_VGND_c_2322_n 0.12791f $X=13.785 $Y=0.18 $X2=0
+ $Y2=0
cc_1136 N_A_1840_21#_c_1628_n N_VGND_c_2322_n 0.00600134f $X=9.35 $Y=0.18 $X2=0
+ $Y2=0
cc_1137 N_A_1840_21#_c_1632_n N_VGND_c_2322_n 0.00962445f $X=14.177 $Y=1.165
+ $X2=0 $Y2=0
cc_1138 N_A_1840_21#_M1014_g N_A_1670_93#_c_2482_n 0.0100481f $X=9.275 $Y=0.785
+ $X2=0 $Y2=0
cc_1139 N_A_1840_21#_M1014_g N_A_1670_93#_c_2483_n 8.90911e-19 $X=9.275 $Y=0.785
+ $X2=0 $Y2=0
cc_1140 N_A_1840_21#_M1014_g N_A_1670_93#_c_2481_n 0.00225586f $X=9.275 $Y=0.785
+ $X2=0 $Y2=0
cc_1141 N_A_1840_21#_c_1632_n N_A_2574_119#_M1031_d 0.00232419f $X=14.177
+ $Y=1.165 $X2=0 $Y2=0
cc_1142 N_A_1840_21#_c_1627_n N_A_2574_119#_c_2507_n 0.00779334f $X=13.785
+ $Y=0.18 $X2=0 $Y2=0
cc_1143 N_A_1840_21#_M1031_g N_A_2574_119#_c_2507_n 0.0152481f $X=13.86 $Y=0.675
+ $X2=0 $Y2=0
cc_1144 N_A_1840_21#_c_1632_n N_A_2574_119#_c_2508_n 0.0290521f $X=14.177
+ $Y=1.165 $X2=0 $Y2=0
cc_1145 N_A_1840_21#_c_1634_n N_A_2574_119#_c_2508_n 0.00152709f $X=14.175
+ $Y=1.54 $X2=0 $Y2=0
cc_1146 N_A_1840_21#_c_1627_n N_A_2574_119#_c_2509_n 0.00788421f $X=13.785
+ $Y=0.18 $X2=0 $Y2=0
cc_1147 N_A_1840_21#_M1031_g N_A_2574_119#_c_2509_n 0.00146115f $X=13.86
+ $Y=0.675 $X2=0 $Y2=0
cc_1148 N_RESET_B_M1040_g N_VPWR_c_1916_n 0.00312414f $X=14.845 $Y=2.155 $X2=0
+ $Y2=0
cc_1149 N_RESET_B_M1040_g N_VPWR_c_1889_n 0.00410284f $X=14.845 $Y=2.155 $X2=0
+ $Y2=0
cc_1150 N_RESET_B_M1032_g N_VGND_c_2298_n 0.00546601f $X=14.85 $Y=0.895 $X2=0
+ $Y2=0
cc_1151 N_RESET_B_M1032_g N_VGND_c_2312_n 0.00370937f $X=14.85 $Y=0.895 $X2=0
+ $Y2=0
cc_1152 N_RESET_B_M1032_g N_VGND_c_2322_n 0.00453162f $X=14.85 $Y=0.895 $X2=0
+ $Y2=0
cc_1153 N_RESET_B_M1032_g N_A_2574_119#_c_2508_n 0.00301278f $X=14.85 $Y=0.895
+ $X2=0 $Y2=0
cc_1154 N_A_3289_47#_c_1780_n N_VPWR_c_1899_n 0.05409f $X=16.59 $Y=2.125 $X2=0
+ $Y2=0
cc_1155 N_A_3289_47#_M1002_g N_VPWR_c_1900_n 0.0057288f $X=17.315 $Y=2.465 $X2=0
+ $Y2=0
cc_1156 N_A_3289_47#_c_1780_n N_VPWR_c_1900_n 0.0365448f $X=16.59 $Y=2.125 $X2=0
+ $Y2=0
cc_1157 N_A_3289_47#_c_1781_n N_VPWR_c_1900_n 0.0137074f $X=17.1 $Y=1.35 $X2=0
+ $Y2=0
cc_1158 N_A_3289_47#_c_1783_n N_VPWR_c_1900_n 0.00536034f $X=17.39 $Y=1.35 $X2=0
+ $Y2=0
cc_1159 N_A_3289_47#_M1034_g N_VPWR_c_1902_n 0.00858314f $X=17.745 $Y=2.465
+ $X2=0 $Y2=0
cc_1160 N_A_3289_47#_c_1780_n N_VPWR_c_1918_n 0.00589611f $X=16.59 $Y=2.125
+ $X2=0 $Y2=0
cc_1161 N_A_3289_47#_M1002_g N_VPWR_c_1919_n 0.00549284f $X=17.315 $Y=2.465
+ $X2=0 $Y2=0
cc_1162 N_A_3289_47#_M1034_g N_VPWR_c_1919_n 0.00549284f $X=17.745 $Y=2.465
+ $X2=0 $Y2=0
cc_1163 N_A_3289_47#_M1002_g N_VPWR_c_1889_n 0.0110929f $X=17.315 $Y=2.465 $X2=0
+ $Y2=0
cc_1164 N_A_3289_47#_M1034_g N_VPWR_c_1889_n 0.0107443f $X=17.745 $Y=2.465 $X2=0
+ $Y2=0
cc_1165 N_A_3289_47#_c_1780_n N_VPWR_c_1889_n 0.00952683f $X=16.59 $Y=2.125
+ $X2=0 $Y2=0
cc_1166 N_A_3289_47#_c_1779_n N_Q_N_c_2233_n 0.00170366f $X=16.59 $Y=0.445 $X2=0
+ $Y2=0
cc_1167 N_A_3289_47#_c_1780_n N_Q_N_c_2233_n 0.0079232f $X=16.59 $Y=2.125 $X2=0
+ $Y2=0
cc_1168 N_A_3289_47#_c_1782_n N_Q_N_c_2233_n 0.00941547f $X=16.59 $Y=1.35 $X2=0
+ $Y2=0
cc_1169 N_A_3289_47#_c_1773_n N_Q_c_2270_n 0.0143929f $X=17.315 $Y=1.185 $X2=0
+ $Y2=0
cc_1170 N_A_3289_47#_M1002_g N_Q_c_2270_n 0.025152f $X=17.315 $Y=2.465 $X2=0
+ $Y2=0
cc_1171 N_A_3289_47#_c_1775_n N_Q_c_2270_n 0.00874467f $X=17.67 $Y=1.26 $X2=0
+ $Y2=0
cc_1172 N_A_3289_47#_c_1776_n N_Q_c_2270_n 0.0157454f $X=17.745 $Y=1.185 $X2=0
+ $Y2=0
cc_1173 N_A_3289_47#_M1034_g N_Q_c_2270_n 0.0422869f $X=17.745 $Y=2.465 $X2=0
+ $Y2=0
cc_1174 N_A_3289_47#_c_1778_n N_Q_c_2270_n 0.00651517f $X=17.745 $Y=1.26 $X2=0
+ $Y2=0
cc_1175 N_A_3289_47#_c_1779_n N_Q_c_2270_n 0.00538817f $X=16.59 $Y=0.445 $X2=0
+ $Y2=0
cc_1176 N_A_3289_47#_c_1780_n N_Q_c_2270_n 0.00875623f $X=16.59 $Y=2.125 $X2=0
+ $Y2=0
cc_1177 N_A_3289_47#_c_1781_n N_Q_c_2270_n 0.0250026f $X=17.1 $Y=1.35 $X2=0
+ $Y2=0
cc_1178 N_A_3289_47#_c_1783_n N_Q_c_2270_n 0.00764151f $X=17.39 $Y=1.35 $X2=0
+ $Y2=0
cc_1179 N_A_3289_47#_c_1779_n N_VGND_c_2299_n 0.0541506f $X=16.59 $Y=0.445 $X2=0
+ $Y2=0
cc_1180 N_A_3289_47#_c_1773_n N_VGND_c_2300_n 0.00330886f $X=17.315 $Y=1.185
+ $X2=0 $Y2=0
cc_1181 N_A_3289_47#_c_1779_n N_VGND_c_2300_n 0.0390339f $X=16.59 $Y=0.445 $X2=0
+ $Y2=0
cc_1182 N_A_3289_47#_c_1781_n N_VGND_c_2300_n 0.0195835f $X=17.1 $Y=1.35 $X2=0
+ $Y2=0
cc_1183 N_A_3289_47#_c_1783_n N_VGND_c_2300_n 0.0057457f $X=17.39 $Y=1.35 $X2=0
+ $Y2=0
cc_1184 N_A_3289_47#_c_1776_n N_VGND_c_2302_n 0.00800849f $X=17.745 $Y=1.185
+ $X2=0 $Y2=0
cc_1185 N_A_3289_47#_c_1779_n N_VGND_c_2314_n 0.0167325f $X=16.59 $Y=0.445 $X2=0
+ $Y2=0
cc_1186 N_A_3289_47#_c_1773_n N_VGND_c_2315_n 0.00549284f $X=17.315 $Y=1.185
+ $X2=0 $Y2=0
cc_1187 N_A_3289_47#_c_1776_n N_VGND_c_2315_n 0.00549284f $X=17.745 $Y=1.185
+ $X2=0 $Y2=0
cc_1188 N_A_3289_47#_M1038_s N_VGND_c_2322_n 0.00234843f $X=16.445 $Y=0.235
+ $X2=0 $Y2=0
cc_1189 N_A_3289_47#_c_1773_n N_VGND_c_2322_n 0.00999943f $X=17.315 $Y=1.185
+ $X2=0 $Y2=0
cc_1190 N_A_3289_47#_c_1776_n N_VGND_c_2322_n 0.0107443f $X=17.745 $Y=1.185
+ $X2=0 $Y2=0
cc_1191 N_A_3289_47#_c_1779_n N_VGND_c_2322_n 0.0123752f $X=16.59 $Y=0.445 $X2=0
+ $Y2=0
cc_1192 N_A_56_481#_c_1839_n N_VPWR_c_1890_n 0.0240561f $X=0.425 $Y=2.55 $X2=0
+ $Y2=0
cc_1193 N_A_56_481#_c_1840_n N_VPWR_c_1890_n 0.0233617f $X=1.3 $Y=2.15 $X2=0
+ $Y2=0
cc_1194 N_A_56_481#_c_1842_n N_VPWR_c_1890_n 0.0312336f $X=1.385 $Y=2.895 $X2=0
+ $Y2=0
cc_1195 N_A_56_481#_c_1844_n N_VPWR_c_1890_n 0.0124177f $X=1.47 $Y=2.98 $X2=0
+ $Y2=0
cc_1196 N_A_56_481#_c_1843_n N_VPWR_c_1891_n 0.0121618f $X=2.16 $Y=2.98 $X2=0
+ $Y2=0
cc_1197 N_A_56_481#_c_1845_n N_VPWR_c_1891_n 0.0316534f $X=2.325 $Y=2.55 $X2=0
+ $Y2=0
cc_1198 N_A_56_481#_c_1839_n N_VPWR_c_1903_n 0.0220321f $X=0.425 $Y=2.55 $X2=0
+ $Y2=0
cc_1199 N_A_56_481#_c_1843_n N_VPWR_c_1905_n 0.0631546f $X=2.16 $Y=2.98 $X2=0
+ $Y2=0
cc_1200 N_A_56_481#_c_1844_n N_VPWR_c_1905_n 0.0114448f $X=1.47 $Y=2.98 $X2=0
+ $Y2=0
cc_1201 N_A_56_481#_c_1839_n N_VPWR_c_1889_n 0.0125808f $X=0.425 $Y=2.55 $X2=0
+ $Y2=0
cc_1202 N_A_56_481#_c_1843_n N_VPWR_c_1889_n 0.0371942f $X=2.16 $Y=2.98 $X2=0
+ $Y2=0
cc_1203 N_A_56_481#_c_1844_n N_VPWR_c_1889_n 0.00655481f $X=1.47 $Y=2.98 $X2=0
+ $Y2=0
cc_1204 N_A_56_481#_c_1842_n A_245_481# 0.00427037f $X=1.385 $Y=2.895 $X2=-0.19
+ $Y2=1.655
cc_1205 N_A_56_481#_c_1844_n A_245_481# 0.00135713f $X=1.47 $Y=2.98 $X2=-0.19
+ $Y2=1.655
cc_1206 N_A_56_481#_c_1843_n N_A_202_119#_M1051_d 0.00382665f $X=2.16 $Y=2.98
+ $X2=0 $Y2=0
cc_1207 N_A_56_481#_c_1840_n N_A_202_119#_c_2089_n 0.00237012f $X=1.3 $Y=2.15
+ $X2=0 $Y2=0
cc_1208 N_A_56_481#_c_1842_n N_A_202_119#_c_2089_n 0.022259f $X=1.385 $Y=2.895
+ $X2=0 $Y2=0
cc_1209 N_A_56_481#_c_1843_n N_A_202_119#_c_2089_n 0.0222237f $X=2.16 $Y=2.98
+ $X2=0 $Y2=0
cc_1210 N_A_56_481#_c_1845_n N_A_202_119#_c_2089_n 0.0125869f $X=2.325 $Y=2.55
+ $X2=0 $Y2=0
cc_1211 N_A_56_481#_c_1845_n N_A_202_119#_c_2091_n 0.026401f $X=2.325 $Y=2.55
+ $X2=0 $Y2=0
cc_1212 N_A_56_481#_c_1840_n N_A_202_119#_c_2096_n 0.0119486f $X=1.3 $Y=2.15
+ $X2=0 $Y2=0
cc_1213 N_VPWR_M1028_s N_A_202_119#_c_2091_n 0.00454204f $X=2.74 $Y=1.535 $X2=0
+ $Y2=0
cc_1214 N_VPWR_M1025_s N_A_202_119#_c_2091_n 0.00767446f $X=3.68 $Y=2.055 $X2=0
+ $Y2=0
cc_1215 N_VPWR_c_1891_n N_A_202_119#_c_2091_n 0.0223859f $X=2.885 $Y=2.59 $X2=0
+ $Y2=0
cc_1216 N_VPWR_c_1892_n N_A_202_119#_c_2091_n 0.0194396f $X=3.81 $Y=2.55 $X2=0
+ $Y2=0
cc_1217 N_VPWR_c_1892_n N_A_202_119#_c_2092_n 0.0358359f $X=3.81 $Y=2.55 $X2=0
+ $Y2=0
cc_1218 N_VPWR_c_1893_n N_A_202_119#_c_2093_n 0.00962064f $X=5.525 $Y=2.84 $X2=0
+ $Y2=0
cc_1219 N_VPWR_c_1913_n N_A_202_119#_c_2093_n 0.057793f $X=5.36 $Y=3.33 $X2=0
+ $Y2=0
cc_1220 N_VPWR_c_1889_n N_A_202_119#_c_2093_n 0.03516f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1221 N_VPWR_c_1892_n N_A_202_119#_c_2094_n 0.0141601f $X=3.81 $Y=2.55 $X2=0
+ $Y2=0
cc_1222 N_VPWR_c_1913_n N_A_202_119#_c_2094_n 0.0114622f $X=5.36 $Y=3.33 $X2=0
+ $Y2=0
cc_1223 N_VPWR_c_1889_n N_A_202_119#_c_2094_n 0.00657784f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1224 N_VPWR_M1008_d N_A_202_119#_c_2097_n 0.00284423f $X=5.385 $Y=2.345 $X2=0
+ $Y2=0
cc_1225 N_VPWR_c_1893_n N_A_202_119#_c_2097_n 0.0205112f $X=5.525 $Y=2.84 $X2=0
+ $Y2=0
cc_1226 N_VPWR_c_1889_n N_A_202_119#_c_2097_n 0.0132566f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1227 N_VPWR_c_1893_n N_A_202_119#_c_2098_n 0.00551243f $X=5.525 $Y=2.84 $X2=0
+ $Y2=0
cc_1228 N_VPWR_c_1909_n N_A_202_119#_c_2098_n 0.00729963f $X=7.955 $Y=3.33 $X2=0
+ $Y2=0
cc_1229 N_VPWR_c_1889_n N_A_202_119#_c_2098_n 0.00891423f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1230 N_VPWR_c_1889_n A_2714_451# 0.00326794f $X=18 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1231 N_VPWR_c_1889_n N_Q_N_M1001_s 0.00415099f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1232 N_VPWR_c_1899_n Q_N 0.0897723f $X=16.03 $Y=1.98 $X2=0 $Y2=0
cc_1233 N_VPWR_c_1917_n Q_N 0.0163333f $X=15.945 $Y=3.33 $X2=0 $Y2=0
cc_1234 N_VPWR_c_1889_n Q_N 0.0104297f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1235 N_VPWR_c_1889_n N_Q_M1002_d 0.00223819f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1236 N_VPWR_c_1900_n N_Q_c_2270_n 0.0455296f $X=17.1 $Y=1.98 $X2=0 $Y2=0
cc_1237 N_VPWR_c_1902_n N_Q_c_2270_n 0.0455296f $X=17.96 $Y=1.98 $X2=0 $Y2=0
cc_1238 N_VPWR_c_1919_n N_Q_c_2270_n 0.0177952f $X=17.875 $Y=3.33 $X2=0 $Y2=0
cc_1239 N_VPWR_c_1889_n N_Q_c_2270_n 0.0123247f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1240 N_A_202_119#_c_2083_n N_VGND_c_2291_n 0.0128148f $X=1.15 $Y=0.805 $X2=0
+ $Y2=0
cc_1241 N_A_202_119#_c_2085_n N_VGND_c_2291_n 0.00573253f $X=1.315 $Y=0.545
+ $X2=0 $Y2=0
cc_1242 N_A_202_119#_c_2084_n N_VGND_c_2292_n 0.013629f $X=1.975 $Y=0.545 $X2=0
+ $Y2=0
cc_1243 N_A_202_119#_c_2086_n N_VGND_c_2292_n 0.0265199f $X=2.06 $Y=2.035 $X2=0
+ $Y2=0
cc_1244 N_A_202_119#_c_2088_n N_VGND_c_2294_n 0.00817197f $X=6.075 $Y=0.895
+ $X2=0 $Y2=0
cc_1245 N_A_202_119#_c_2088_n N_VGND_c_2305_n 0.00609437f $X=6.075 $Y=0.895
+ $X2=0 $Y2=0
cc_1246 N_A_202_119#_c_2084_n N_VGND_c_2309_n 0.023626f $X=1.975 $Y=0.545 $X2=0
+ $Y2=0
cc_1247 N_A_202_119#_c_2085_n N_VGND_c_2309_n 0.00998302f $X=1.315 $Y=0.545
+ $X2=0 $Y2=0
cc_1248 N_A_202_119#_c_2084_n N_VGND_c_2322_n 0.0240741f $X=1.975 $Y=0.545 $X2=0
+ $Y2=0
cc_1249 N_A_202_119#_c_2085_n N_VGND_c_2322_n 0.00990635f $X=1.315 $Y=0.545
+ $X2=0 $Y2=0
cc_1250 N_A_202_119#_c_2088_n N_VGND_c_2322_n 0.00833638f $X=6.075 $Y=0.895
+ $X2=0 $Y2=0
cc_1251 N_A_202_119#_c_2084_n A_323_119# 0.00815797f $X=1.975 $Y=0.545 $X2=-0.19
+ $Y2=-0.245
cc_1252 N_A_202_119#_c_2086_n A_323_119# 0.00462203f $X=2.06 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_1253 N_Q_N_c_2231_n N_VGND_c_2298_n 0.0318617f $X=15.575 $Y=0.43 $X2=0 $Y2=0
cc_1254 N_Q_N_c_2231_n N_VGND_c_2299_n 0.0628727f $X=15.575 $Y=0.43 $X2=0 $Y2=0
cc_1255 N_Q_N_c_2231_n N_VGND_c_2313_n 0.0193942f $X=15.575 $Y=0.43 $X2=0 $Y2=0
cc_1256 N_Q_N_c_2231_n N_VGND_c_2322_n 0.0133019f $X=15.575 $Y=0.43 $X2=0 $Y2=0
cc_1257 N_Q_c_2270_n N_VGND_c_2302_n 0.0304763f $X=17.53 $Y=0.43 $X2=0 $Y2=0
cc_1258 N_Q_c_2270_n N_VGND_c_2315_n 0.0177952f $X=17.53 $Y=0.43 $X2=0 $Y2=0
cc_1259 N_Q_M1003_d N_VGND_c_2322_n 0.00223819f $X=17.39 $Y=0.235 $X2=0 $Y2=0
cc_1260 N_Q_c_2270_n N_VGND_c_2322_n 0.0123247f $X=17.53 $Y=0.43 $X2=0 $Y2=0
cc_1261 N_VGND_c_2312_n N_A_2574_119#_c_2507_n 0.0606913f $X=14.98 $Y=0 $X2=0
+ $Y2=0
cc_1262 N_VGND_c_2322_n N_A_2574_119#_c_2507_n 0.0342536f $X=18 $Y=0 $X2=0 $Y2=0
cc_1263 N_VGND_c_2297_n N_A_2574_119#_c_2509_n 0.0203686f $X=12.5 $Y=0.485 $X2=0
+ $Y2=0
cc_1264 N_VGND_c_2312_n N_A_2574_119#_c_2509_n 0.0211946f $X=14.98 $Y=0 $X2=0
+ $Y2=0
cc_1265 N_VGND_c_2322_n N_A_2574_119#_c_2509_n 0.0111959f $X=18 $Y=0 $X2=0 $Y2=0
