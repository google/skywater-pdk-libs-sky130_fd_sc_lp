* File: sky130_fd_sc_lp__a2111o_1.pex.spice
* Created: Fri Aug 28 09:45:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111O_1%A_105_239# 1 2 3 12 14 16 20 21 22 23 24 25
+ 28 34 36 40 42
c81 36 0 1.21937e-19 $X=2.53 $Y=1.08
r82 43 45 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.6 $Y=1.36 $X2=0.64
+ $Y2=1.36
r83 38 40 9.68655 $w=7.08e-07 $l=5.75e-07 $layer=LI1_cond $X=2.885 $Y=0.995
+ $X2=2.885 $Y2=0.42
r84 37 42 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.86 $Y=1.08
+ $X2=1.745 $Y2=1.08
r85 36 38 80.387 $w=5.9e-08 $l=3.95221e-07 $layer=LI1_cond $X=2.53 $Y=1.08
+ $X2=2.885 $Y2=0.995
r86 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.53 $Y=1.08
+ $X2=1.86 $Y2=1.08
r87 32 42 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=0.995
+ $X2=1.745 $Y2=1.08
r88 32 34 28.8111 $w=2.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.745 $Y=0.995
+ $X2=1.745 $Y2=0.42
r89 28 30 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=1.335 $Y=2.095
+ $X2=1.335 $Y2=2.91
r90 26 28 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.335 $Y=2.09
+ $X2=1.335 $Y2=2.095
r91 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=2.005
+ $X2=1.335 $Y2=2.09
r92 24 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.17 $Y=2.005
+ $X2=0.905 $Y2=2.005
r93 22 42 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.63 $Y=1.08
+ $X2=1.745 $Y2=1.08
r94 22 23 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.63 $Y=1.08
+ $X2=0.905 $Y2=1.08
r95 21 45 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.795 $Y=1.36
+ $X2=0.64 $Y2=1.36
r96 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.795
+ $Y=1.36 $X2=0.795 $Y2=1.36
r97 18 25 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=0.797 $Y=1.92
+ $X2=0.905 $Y2=2.005
r98 18 20 30.0171 $w=2.13e-07 $l=5.6e-07 $layer=LI1_cond $X=0.797 $Y=1.92
+ $X2=0.797 $Y2=1.36
r99 17 23 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=0.797 $Y=1.165
+ $X2=0.905 $Y2=1.08
r100 17 20 10.4524 $w=2.13e-07 $l=1.95e-07 $layer=LI1_cond $X=0.797 $Y=1.165
+ $X2=0.797 $Y2=1.36
r101 14 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=1.195
+ $X2=0.64 $Y2=1.36
r102 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.64 $Y=1.195
+ $X2=0.64 $Y2=0.665
r103 10 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.525
+ $X2=0.6 $Y2=1.36
r104 10 12 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=0.6 $Y=1.525 $X2=0.6
+ $Y2=2.465
r105 3 30 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.21
+ $Y=1.835 $X2=1.335 $Y2=2.91
r106 3 28 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=1.21
+ $Y=1.835 $X2=1.335 $Y2=2.095
r107 2 40 45.5 $w=1.7e-07 $l=6.01166e-07 $layer=licon1_NDIFF $count=4 $X=2.555
+ $Y=0.245 $X2=3.075 $Y2=0.42
r108 1 34 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.585
+ $Y=0.245 $X2=1.725 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_1%D1 3 7 9 10 14
c36 3 0 6.66526e-21 $X=1.51 $Y=0.665
r37 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.46 $Y=1.51
+ $X2=1.46 $Y2=1.675
r38 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.46 $Y=1.51
+ $X2=1.46 $Y2=1.345
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.46
+ $Y=1.51 $X2=1.46 $Y2=1.51
r40 10 15 6.10934 $w=4.13e-07 $l=2.2e-07 $layer=LI1_cond $X=1.68 $Y=1.542
+ $X2=1.46 $Y2=1.542
r41 9 15 7.22012 $w=4.13e-07 $l=2.6e-07 $layer=LI1_cond $X=1.2 $Y=1.542 $X2=1.46
+ $Y2=1.542
r42 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.55 $Y=2.465
+ $X2=1.55 $Y2=1.675
r43 3 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.51 $Y=0.665
+ $X2=1.51 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_1%C1 3 7 9 10 11 12 18 19
c39 19 0 6.66526e-21 $X=2.03 $Y=1.51
c40 7 0 1.96363e-19 $X=1.94 $Y=2.465
c41 3 0 7.72595e-21 $X=1.94 $Y=0.665
r42 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=1.51
+ $X2=2.03 $Y2=1.675
r43 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=1.51
+ $X2=2.03 $Y2=1.345
r44 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.51 $X2=2.03 $Y2=1.51
r45 11 12 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.105 $Y=2.405
+ $X2=2.105 $Y2=2.775
r46 10 11 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=2.105 $Y2=2.405
r47 9 10 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.105 $Y=1.665
+ $X2=2.105 $Y2=2.035
r48 9 19 5.58215 $w=3.18e-07 $l=1.55e-07 $layer=LI1_cond $X=2.105 $Y=1.665
+ $X2=2.105 $Y2=1.51
r49 7 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.94 $Y=2.465
+ $X2=1.94 $Y2=1.675
r50 3 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.94 $Y=0.665
+ $X2=1.94 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_1%B1 3 7 9 12 13
c36 13 0 7.12504e-20 $X=2.6 $Y=1.51
r37 12 15 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.51 $X2=2.6
+ $Y2=1.675
r38 12 14 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.51 $X2=2.6
+ $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.6
+ $Y=1.51 $X2=2.6 $Y2=1.51
r40 9 13 4.63971 $w=3.83e-07 $l=1.55e-07 $layer=LI1_cond $X=2.627 $Y=1.665
+ $X2=2.627 $Y2=1.51
r41 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.48 $Y=2.465
+ $X2=2.48 $Y2=1.675
r42 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.48 $Y=0.665
+ $X2=2.48 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_1%A1 3 7 8 10 17 19
c37 17 0 1.60131e-19 $X=3.2 $Y=1.375
r38 17 20 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.185 $Y=1.375
+ $X2=3.185 $Y2=1.54
r39 17 19 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.185 $Y=1.375
+ $X2=3.185 $Y2=1.21
r40 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.375 $X2=3.2 $Y2=1.375
r41 10 18 8.69875 $w=5.48e-07 $l=4e-07 $layer=LI1_cond $X=3.6 $Y=1.485 $X2=3.2
+ $Y2=1.485
r42 8 18 1.73975 $w=5.48e-07 $l=8e-08 $layer=LI1_cond $X=3.12 $Y=1.485 $X2=3.2
+ $Y2=1.485
r43 7 19 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.29 $Y=0.665
+ $X2=3.29 $Y2=1.21
r44 3 20 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.25 $Y=2.465
+ $X2=3.25 $Y2=1.54
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_1%A2 1 3 6 8 9 16
c24 8 0 1.60131e-19 $X=4.08 $Y=1.295
c25 1 0 1.21937e-19 $X=3.65 $Y=1.21
r26 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.375 $X2=3.95 $Y2=1.375
r27 14 16 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.68 $Y=1.375
+ $X2=3.95 $Y2=1.375
r28 12 14 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.65 $Y=1.375 $X2=3.68
+ $Y2=1.375
r29 9 17 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.05 $Y=1.665
+ $X2=4.05 $Y2=1.375
r30 8 17 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=4.05 $Y=1.295 $X2=4.05
+ $Y2=1.375
r31 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.54
+ $X2=3.68 $Y2=1.375
r32 4 6 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.68 $Y=1.54 $X2=3.68
+ $Y2=2.465
r33 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.21
+ $X2=3.65 $Y2=1.375
r34 1 3 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.65 $Y=1.21 $X2=3.65
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_1%X 1 2 7 8 9 10 11 12 13 23 33
r17 33 45 5.98103 $w=3.93e-07 $l=2.05e-07 $layer=LI1_cond $X=0.282 $Y=1.98
+ $X2=0.282 $Y2=1.775
r18 13 41 3.93873 $w=3.93e-07 $l=1.35e-07 $layer=LI1_cond $X=0.282 $Y=2.775
+ $X2=0.282 $Y2=2.91
r19 12 13 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.282 $Y=2.405
+ $X2=0.282 $Y2=2.775
r20 11 12 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.282 $Y=2.035
+ $X2=0.282 $Y2=2.405
r21 11 33 1.60467 $w=3.93e-07 $l=5.5e-08 $layer=LI1_cond $X=0.282 $Y=2.035
+ $X2=0.282 $Y2=1.98
r22 10 45 3.03487 $w=4.33e-07 $l=1.1e-07 $layer=LI1_cond $X=0.302 $Y=1.665
+ $X2=0.302 $Y2=1.775
r23 10 21 2.83474 $w=4.33e-07 $l=1.07e-07 $layer=LI1_cond $X=0.302 $Y=1.665
+ $X2=0.302 $Y2=1.558
r24 9 21 6.96764 $w=4.33e-07 $l=2.63e-07 $layer=LI1_cond $X=0.302 $Y=1.295
+ $X2=0.302 $Y2=1.558
r25 8 9 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.302 $Y=0.925
+ $X2=0.302 $Y2=1.295
r26 7 8 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.302 $Y=0.555
+ $X2=0.302 $Y2=0.925
r27 7 23 3.57655 $w=4.33e-07 $l=1.35e-07 $layer=LI1_cond $X=0.302 $Y=0.555
+ $X2=0.302 $Y2=0.42
r28 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.835 $X2=0.385 $Y2=2.91
r29 2 33 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.835 $X2=0.385 $Y2=1.98
r30 1 23 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=0.3
+ $Y=0.245 $X2=0.425 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_1%VPWR 1 2 11 15 18 19 20 30 31 34
r48 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r51 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 24 27 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r56 22 24 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 20 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 20 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 18 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.3 $Y=3.33 $X2=3.12
+ $Y2=3.33
r60 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=3.33
+ $X2=3.465 $Y2=3.33
r61 17 30 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=3.465 $Y2=3.33
r63 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=3.245
+ $X2=3.465 $Y2=3.33
r64 13 15 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3.465 $Y=3.245
+ $X2=3.465 $Y2=2.375
r65 9 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r66 9 11 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.365
r67 2 15 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=3.325
+ $Y=1.835 $X2=3.465 $Y2=2.375
r68 1 11 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=0.675
+ $Y=1.835 $X2=0.815 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_1%A_511_367# 1 2 7 9 11 13 15
c24 7 0 1.32838e-19 $X=2.83 $Y=2.1
r25 13 20 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=2.1 $X2=3.93
+ $Y2=2.015
r26 13 15 16.6218 $w=2.58e-07 $l=3.75e-07 $layer=LI1_cond $X=3.93 $Y=2.1
+ $X2=3.93 $Y2=2.475
r27 12 18 7.82736 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=3.13 $Y=2.015 $X2=2.83
+ $Y2=2.015
r28 11 20 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.8 $Y=2.015 $X2=3.93
+ $Y2=2.015
r29 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.8 $Y=2.015
+ $X2=3.13 $Y2=2.015
r30 7 18 2.21775 $w=6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.83 $Y=2.1 $X2=2.83
+ $Y2=2.015
r31 7 9 7.47549 $w=5.98e-07 $l=3.75e-07 $layer=LI1_cond $X=2.83 $Y=2.1 $X2=2.83
+ $Y2=2.475
r32 2 20 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=1.835 $X2=3.895 $Y2=2.015
r33 2 15 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=3.755
+ $Y=1.835 $X2=3.895 $Y2=2.475
r34 1 18 300 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=2 $X=2.555
+ $Y=1.835 $X2=3.035 $Y2=2.015
r35 1 9 150 $w=1.7e-07 $l=8.4664e-07 $layer=licon1_PDIFF $count=4 $X=2.555
+ $Y=1.835 $X2=3.035 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_1%VGND 1 2 3 14 18 20 21 22 23 25 39 42 50
r48 43 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r49 42 47 5.74739 $w=7.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=1.075
+ $Y2=0.37
r50 42 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r53 36 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r54 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r56 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r57 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r58 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.195
+ $Y2=0
r59 30 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.64
+ $Y2=0
r60 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r61 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r62 26 42 9.95332 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=1.46 $Y=0 $X2=1.075
+ $Y2=0
r63 26 28 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.46 $Y=0 $X2=1.68
+ $Y2=0
r64 25 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.195
+ $Y2=0
r65 25 28 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=1.68
+ $Y2=0
r66 23 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r67 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r68 23 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r69 21 35 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.6 $Y2=0
r70 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.865
+ $Y2=0
r71 20 38 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=4.03 $Y=0 $X2=4.08
+ $Y2=0
r72 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.03 $Y=0 $X2=3.865
+ $Y2=0
r73 16 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=0.085
+ $X2=3.865 $Y2=0
r74 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.865 $Y=0.085
+ $X2=3.865 $Y2=0.39
r75 12 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0
r76 12 14 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0.37
r77 3 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.725
+ $Y=0.245 $X2=3.865 $Y2=0.39
r78 2 14 91 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=2 $X=2.015
+ $Y=0.245 $X2=2.195 $Y2=0.37
r79 1 47 45.5 $w=1.7e-07 $l=6.39453e-07 $layer=licon1_NDIFF $count=4 $X=0.715
+ $Y=0.245 $X2=1.295 $Y2=0.37
.ends

