* File: sky130_fd_sc_lp__o31a_4.pex.spice
* Created: Wed Sep  2 10:24:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31A_4%A_101_23# 1 2 3 12 16 20 24 28 32 36 40 42 51
+ 55 58 59 60 64 68 70 72 83
c129 58 0 8.21834e-20 $X=3.13 $Y=1.16
r130 80 81 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.665 $Y=1.49
+ $X2=1.87 $Y2=1.49
r131 79 80 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.44 $Y=1.49
+ $X2=1.665 $Y2=1.49
r132 78 79 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.235 $Y=1.49
+ $X2=1.44 $Y2=1.49
r133 77 78 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.01 $Y=1.49
+ $X2=1.235 $Y2=1.49
r134 76 77 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.805 $Y=1.49
+ $X2=1.01 $Y2=1.49
r135 62 64 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.295 $Y=1.075
+ $X2=3.295 $Y2=0.69
r136 61 70 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.835 $Y=2.375
+ $X2=2.74 $Y2=2.375
r137 60 72 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.99 $Y=2.375
+ $X2=4.125 $Y2=2.375
r138 60 61 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=3.99 $Y=2.375
+ $X2=2.835 $Y2=2.375
r139 58 62 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.13 $Y=1.16
+ $X2=3.295 $Y2=1.075
r140 58 59 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.13 $Y=1.16
+ $X2=2.835 $Y2=1.16
r141 53 70 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=2.29
+ $X2=2.74 $Y2=2.375
r142 53 55 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=2.74 $Y=2.29
+ $X2=2.74 $Y2=1.98
r143 52 68 4.60183 $w=1.95e-07 $l=8.74643e-08 $layer=LI1_cond $X=2.74 $Y=1.575
+ $X2=2.735 $Y2=1.49
r144 52 55 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=2.74 $Y=1.575
+ $X2=2.74 $Y2=1.98
r145 51 68 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=1.405
+ $X2=2.735 $Y2=1.49
r146 50 59 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.735 $Y=1.245
+ $X2=2.835 $Y2=1.16
r147 50 51 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.735 $Y=1.245
+ $X2=2.735 $Y2=1.405
r148 49 83 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=2.03 $Y=1.49
+ $X2=2.095 $Y2=1.49
r149 49 81 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.03 $Y=1.49
+ $X2=1.87 $Y2=1.49
r150 48 49 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.03
+ $Y=1.49 $X2=2.03 $Y2=1.49
r151 45 76 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.67 $Y=1.49
+ $X2=0.805 $Y2=1.49
r152 45 73 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.67 $Y=1.49 $X2=0.58
+ $Y2=1.49
r153 44 48 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.67 $Y=1.49
+ $X2=2.03 $Y2=1.49
r154 44 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.67
+ $Y=1.49 $X2=0.67 $Y2=1.49
r155 42 68 1.84097 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.635 $Y=1.49
+ $X2=2.735 $Y2=1.49
r156 42 48 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.635 $Y=1.49
+ $X2=2.03 $Y2=1.49
r157 38 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.655
+ $X2=2.095 $Y2=1.49
r158 38 40 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.095 $Y=1.655
+ $X2=2.095 $Y2=2.465
r159 34 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.325
+ $X2=1.87 $Y2=1.49
r160 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.87 $Y=1.325
+ $X2=1.87 $Y2=0.665
r161 30 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.655
+ $X2=1.665 $Y2=1.49
r162 30 32 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.665 $Y=1.655
+ $X2=1.665 $Y2=2.465
r163 26 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.44 $Y=1.325
+ $X2=1.44 $Y2=1.49
r164 26 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.44 $Y=1.325
+ $X2=1.44 $Y2=0.665
r165 22 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.235 $Y=1.655
+ $X2=1.235 $Y2=1.49
r166 22 24 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.235 $Y=1.655
+ $X2=1.235 $Y2=2.465
r167 18 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.325
+ $X2=1.01 $Y2=1.49
r168 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.01 $Y=1.325
+ $X2=1.01 $Y2=0.665
r169 14 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.805 $Y=1.655
+ $X2=0.805 $Y2=1.49
r170 14 16 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.805 $Y=1.655
+ $X2=0.805 $Y2=2.465
r171 10 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.325
+ $X2=0.58 $Y2=1.49
r172 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.58 $Y=1.325
+ $X2=0.58 $Y2=0.665
r173 3 72 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=4.015
+ $Y=1.835 $X2=4.155 $Y2=2.455
r174 2 70 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=2.6
+ $Y=1.835 $X2=2.74 $Y2=2.425
r175 2 55 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.6
+ $Y=1.835 $X2=2.74 $Y2=1.98
r176 1 64 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=3.155
+ $Y=0.325 $X2=3.295 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%B1 3 5 6 9 13 17 19 20 26 27
c59 27 0 1.77905e-19 $X=3.17 $Y=1.51
c60 26 0 9.93349e-20 $X=3.17 $Y=1.51
r61 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.51 $X2=3.17 $Y2=1.51
r62 24 26 16.3083 $w=2.66e-07 $l=9e-08 $layer=POLY_cond $X=3.08 $Y=1.51 $X2=3.17
+ $Y2=1.51
r63 23 24 22.6504 $w=2.66e-07 $l=1.25e-07 $layer=POLY_cond $X=2.955 $Y=1.51
+ $X2=3.08 $Y2=1.51
r64 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.17 $Y=1.665
+ $X2=3.17 $Y2=2.035
r65 19 27 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.17 $Y=1.665
+ $X2=3.17 $Y2=1.51
r66 15 26 61.609 $w=2.66e-07 $l=4.14367e-07 $layer=POLY_cond $X=3.51 $Y=1.345
+ $X2=3.17 $Y2=1.51
r67 15 17 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.51 $Y=1.345 $X2=3.51
+ $Y2=0.745
r68 11 24 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=1.345
+ $X2=3.08 $Y2=1.51
r69 11 13 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.08 $Y=1.345 $X2=3.08
+ $Y2=0.745
r70 7 23 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.675
+ $X2=2.955 $Y2=1.51
r71 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.955 $Y=1.675
+ $X2=2.955 $Y2=2.465
r72 5 23 22.6819 $w=2.66e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.88 $Y=1.42
+ $X2=2.955 $Y2=1.51
r73 5 6 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.88 $Y=1.42 $X2=2.6
+ $Y2=1.42
r74 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.525 $Y=1.495
+ $X2=2.6 $Y2=1.42
r75 1 3 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.525 $Y=1.495
+ $X2=2.525 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%A3 3 7 11 15 17 18 19 28
c52 28 0 1.77905e-19 $X=4.37 $Y=1.51
c53 15 0 3.21372e-20 $X=4.37 $Y=2.465
c54 3 0 8.21834e-20 $X=3.94 $Y=0.745
r55 26 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.03 $Y=1.51
+ $X2=4.37 $Y2=1.51
r56 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.51 $X2=4.03 $Y2=1.51
r57 23 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.94 $Y=1.51 $X2=4.03
+ $Y2=1.51
r58 18 19 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.56 $Y2=1.587
r59 18 27 1.77299 $w=3.23e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.587 $X2=4.03
+ $Y2=1.587
r60 17 27 15.2477 $w=3.23e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.587
+ $X2=4.03 $Y2=1.587
r61 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.675
+ $X2=4.37 $Y2=1.51
r62 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.37 $Y=1.675
+ $X2=4.37 $Y2=2.465
r63 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.345
+ $X2=4.37 $Y2=1.51
r64 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.37 $Y=1.345 $X2=4.37
+ $Y2=0.745
r65 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.94 $Y=1.675
+ $X2=3.94 $Y2=1.51
r66 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.94 $Y=1.675 $X2=3.94
+ $Y2=2.465
r67 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.94 $Y=1.345
+ $X2=3.94 $Y2=1.51
r68 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.94 $Y=1.345 $X2=3.94
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%A2 3 7 11 15 17 21 22 24 28 29 36 41
c76 36 0 3.21372e-20 $X=5.027 $Y=1.705
c77 28 0 1.71625e-19 $X=4.935 $Y=1.51
r78 36 41 1.29853 $w=3.53e-07 $l=4e-08 $layer=LI1_cond $X=5.027 $Y=1.705
+ $X2=5.027 $Y2=1.665
r79 28 31 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.912 $Y=1.51
+ $X2=4.912 $Y2=1.675
r80 28 30 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.912 $Y=1.51
+ $X2=4.912 $Y2=1.345
r81 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.51 $X2=4.935 $Y2=1.51
r82 24 36 2.57906 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.027 $Y=1.79
+ $X2=5.027 $Y2=1.705
r83 24 41 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=5.027 $Y=1.642
+ $X2=5.027 $Y2=1.665
r84 24 29 4.28514 $w=3.53e-07 $l=1.32e-07 $layer=LI1_cond $X=5.027 $Y=1.642
+ $X2=5.027 $Y2=1.51
r85 22 32 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=6.43 $Y=1.46
+ $X2=6.245 $Y2=1.46
r86 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.43
+ $Y=1.46 $X2=6.43 $Y2=1.46
r87 19 21 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.43 $Y=1.705
+ $X2=6.43 $Y2=1.46
r88 18 24 5.40086 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=5.205 $Y=1.79
+ $X2=5.027 $Y2=1.79
r89 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.265 $Y=1.79
+ $X2=6.43 $Y2=1.705
r90 17 18 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=6.265 $Y=1.79
+ $X2=5.205 $Y2=1.79
r91 13 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.625
+ $X2=6.245 $Y2=1.46
r92 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.245 $Y=1.625
+ $X2=6.245 $Y2=2.465
r93 9 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.295
+ $X2=6.245 $Y2=1.46
r94 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.245 $Y=1.295
+ $X2=6.245 $Y2=0.745
r95 7 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.8 $Y=2.465 $X2=4.8
+ $Y2=1.675
r96 3 30 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.8 $Y=0.745 $X2=4.8
+ $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%A1 1 3 6 8 10 13 15 16 24
c54 16 0 1.71625e-19 $X=6 $Y=1.295
r55 22 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.725 $Y=1.44
+ $X2=5.815 $Y2=1.44
r56 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.725
+ $Y=1.44 $X2=5.725 $Y2=1.44
r57 19 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.385 $Y=1.44
+ $X2=5.725 $Y2=1.44
r58 16 23 9.75144 $w=3.23e-07 $l=2.75e-07 $layer=LI1_cond $X=6 $Y=1.372
+ $X2=5.725 $Y2=1.372
r59 15 23 7.26926 $w=3.23e-07 $l=2.05e-07 $layer=LI1_cond $X=5.52 $Y=1.372
+ $X2=5.725 $Y2=1.372
r60 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.605
+ $X2=5.815 $Y2=1.44
r61 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.815 $Y=1.605
+ $X2=5.815 $Y2=2.465
r62 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.275
+ $X2=5.815 $Y2=1.44
r63 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.815 $Y=1.275
+ $X2=5.815 $Y2=0.745
r64 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.605
+ $X2=5.385 $Y2=1.44
r65 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.385 $Y=1.605
+ $X2=5.385 $Y2=2.465
r66 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.275
+ $X2=5.385 $Y2=1.44
r67 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.385 $Y=1.275
+ $X2=5.385 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%VPWR 1 2 3 4 5 18 24 28 32 38 40 45 47 48 49
+ 50 51 60 65 74 77 81
r101 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r102 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 72 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r105 71 72 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r106 69 72 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r107 68 71 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r108 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r109 66 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.17 $Y2=3.33
r110 66 68 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.6 $Y2=3.33
r111 65 80 4.13127 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=6.365 $Y=3.33
+ $X2=6.542 $Y2=3.33
r112 65 71 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.365 $Y=3.33
+ $X2=6 $Y2=3.33
r113 64 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 64 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r116 61 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.31 $Y2=3.33
r117 61 63 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 60 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=3.33
+ $X2=3.17 $Y2=3.33
r119 60 63 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.005 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 59 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r121 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 55 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r124 51 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r125 51 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 49 58 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.45 $Y2=3.33
r128 47 54 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.24 $Y2=3.33
r129 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.59 $Y2=3.33
r130 46 58 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.59 $Y2=3.33
r132 45 80 3.08095 $w=2.6e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.495 $Y=3.245
+ $X2=6.542 $Y2=3.33
r133 44 45 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=6.495 $Y=2.665
+ $X2=6.495 $Y2=3.245
r134 40 44 6.84978 $w=2.3e-07 $l=1.78466e-07 $layer=LI1_cond $X=6.365 $Y=2.55
+ $X2=6.495 $Y2=2.665
r135 40 42 38.3313 $w=2.28e-07 $l=7.65e-07 $layer=LI1_cond $X=6.365 $Y=2.55
+ $X2=5.6 $Y2=2.55
r136 36 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=3.245
+ $X2=3.17 $Y2=3.33
r137 36 38 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.17 $Y=3.245
+ $X2=3.17 $Y2=2.75
r138 32 35 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=2.31 $Y=1.98
+ $X2=2.31 $Y2=2.95
r139 30 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=3.245
+ $X2=2.31 $Y2=3.33
r140 30 35 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.31 $Y=3.245
+ $X2=2.31 $Y2=2.95
r141 29 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=1.45 $Y2=3.33
r142 28 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=2.31 $Y2=3.33
r143 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=1.615 $Y2=3.33
r144 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.45 $Y=2.18
+ $X2=1.45 $Y2=2.95
r145 22 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=3.245
+ $X2=1.45 $Y2=3.33
r146 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.45 $Y=3.245
+ $X2=1.45 $Y2=2.95
r147 18 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.59 $Y=2.18
+ $X2=0.59 $Y2=2.95
r148 16 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.59 $Y=3.245
+ $X2=0.59 $Y2=3.33
r149 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.59 $Y=3.245
+ $X2=0.59 $Y2=2.95
r150 5 42 600 $w=1.7e-07 $l=7.91912e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.56
r151 4 38 600 $w=1.7e-07 $l=9.8251e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.835 $X2=3.17 $Y2=2.75
r152 3 35 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.17
+ $Y=1.835 $X2=2.31 $Y2=2.95
r153 3 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.17
+ $Y=1.835 $X2=2.31 $Y2=1.98
r154 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.31
+ $Y=1.835 $X2=1.45 $Y2=2.95
r155 2 24 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.31
+ $Y=1.835 $X2=1.45 $Y2=2.18
r156 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.465
+ $Y=1.835 $X2=0.59 $Y2=2.95
r157 1 18 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.465
+ $Y=1.835 $X2=0.59 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%X 1 2 3 4 13 15 16 19 21 25 29 33 37 42 43 44
+ 45 49 51
r58 49 51 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=0.21 $Y=1.225 $X2=0.21
+ $Y2=1.295
r59 44 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.21 $Y=1.14 $X2=0.21
+ $Y2=1.225
r60 44 45 16.7335 $w=2.48e-07 $l=3.63e-07 $layer=LI1_cond $X=0.21 $Y=1.302
+ $X2=0.21 $Y2=1.665
r61 44 51 0.322684 $w=2.48e-07 $l=7e-09 $layer=LI1_cond $X=0.21 $Y=1.302
+ $X2=0.21 $Y2=1.295
r62 41 45 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.21 $Y=1.755 $X2=0.21
+ $Y2=1.665
r63 37 39 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=1.885 $Y=1.98
+ $X2=1.885 $Y2=2.91
r64 35 37 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=1.885 $Y=1.925
+ $X2=1.885 $Y2=1.98
r65 31 33 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=1.655 $Y=1.055
+ $X2=1.655 $Y2=0.42
r66 30 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.115 $Y=1.84
+ $X2=1.02 $Y2=1.84
r67 29 35 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.795 $Y=1.84
+ $X2=1.885 $Y2=1.925
r68 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.795 $Y=1.84
+ $X2=1.115 $Y2=1.84
r69 25 27 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.02 $Y=1.98
+ $X2=1.02 $Y2=2.91
r70 23 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.02 $Y=1.925
+ $X2=1.02 $Y2=1.84
r71 23 25 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.02 $Y=1.925
+ $X2=1.02 $Y2=1.98
r72 22 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.89 $Y=1.14
+ $X2=0.795 $Y2=1.14
r73 21 31 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.56 $Y=1.14
+ $X2=1.655 $Y2=1.055
r74 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.56 $Y=1.14
+ $X2=0.89 $Y2=1.14
r75 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=1.055
+ $X2=0.795 $Y2=1.14
r76 17 19 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=0.795 $Y=1.055
+ $X2=0.795 $Y2=0.42
r77 16 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.335 $Y=1.84
+ $X2=0.21 $Y2=1.755
r78 15 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.925 $Y=1.84
+ $X2=1.02 $Y2=1.84
r79 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.925 $Y=1.84
+ $X2=0.335 $Y2=1.84
r80 14 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.335 $Y=1.14
+ $X2=0.21 $Y2=1.14
r81 13 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.7 $Y=1.14 $X2=0.795
+ $Y2=1.14
r82 13 14 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.7 $Y=1.14
+ $X2=0.335 $Y2=1.14
r83 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.835 $X2=1.88 $Y2=2.91
r84 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.835 $X2=1.88 $Y2=1.98
r85 3 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.88
+ $Y=1.835 $X2=1.02 $Y2=2.91
r86 3 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.88
+ $Y=1.835 $X2=1.02 $Y2=1.98
r87 2 33 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.245 $X2=1.655 $Y2=0.42
r88 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.655
+ $Y=0.245 $X2=0.795 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%A_720_367# 1 2 3 10 16 20 23
c43 10 0 9.93349e-20 $X=4.43 $Y=2.02
r44 18 23 7.22005 $w=2.1e-07 $l=1.88892e-07 $layer=LI1_cond $X=4.75 $Y=2.155
+ $X2=4.59 $Y2=2.092
r45 18 20 89.5762 $w=2.18e-07 $l=1.71e-06 $layer=LI1_cond $X=4.75 $Y=2.155
+ $X2=6.46 $Y2=2.155
r46 14 23 0.120199 $w=3.2e-07 $l=1.73e-07 $layer=LI1_cond $X=4.59 $Y=2.265
+ $X2=4.59 $Y2=2.092
r47 14 16 23.2289 $w=3.18e-07 $l=6.45e-07 $layer=LI1_cond $X=4.59 $Y=2.265
+ $X2=4.59 $Y2=2.91
r48 10 23 7.22005 $w=2.1e-07 $l=1.92666e-07 $layer=LI1_cond $X=4.43 $Y=2.02
+ $X2=4.59 $Y2=2.092
r49 10 12 39.0955 $w=1.98e-07 $l=7.05e-07 $layer=LI1_cond $X=4.43 $Y=2.02
+ $X2=3.725 $Y2=2.02
r50 3 20 600 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.16
r51 2 23 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=4.445
+ $Y=1.835 $X2=4.585 $Y2=2.005
r52 2 16 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.445
+ $Y=1.835 $X2=4.585 $Y2=2.91
r53 1 12 600 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=3.6
+ $Y=1.835 $X2=3.725 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%A_975_367# 1 2 7 9 13
r19 11 16 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=5.255 $Y=2.955
+ $X2=5.09 $Y2=2.955
r20 11 13 37.2143 $w=2.38e-07 $l=7.75e-07 $layer=LI1_cond $X=5.255 $Y=2.955
+ $X2=6.03 $Y2=2.955
r21 7 16 2.96416 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=5.09 $Y=2.835 $X2=5.09
+ $Y2=2.955
r22 7 9 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=5.09 $Y=2.835 $X2=5.09
+ $Y2=2.545
r23 2 13 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=1.835 $X2=6.03 $Y2=2.95
r24 1 16 600 $w=1.7e-07 $l=1.21776e-06 $layer=licon1_PDIFF $count=1 $X=4.875
+ $Y=1.835 $X2=5.09 $Y2=2.95
r25 1 9 600 $w=1.7e-07 $l=8.10401e-07 $layer=licon1_PDIFF $count=1 $X=4.875
+ $Y=1.835 $X2=5.09 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 43 45
+ 50 55 63 68 75 76 82 85 88 91 94
r100 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r101 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r102 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r103 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r104 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r105 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r106 76 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r107 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r108 73 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6.03
+ $Y2=0
r109 73 75 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.195 $Y=0
+ $X2=6.48 $Y2=0
r110 72 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r111 72 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r112 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r113 69 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.255 $Y=0 $X2=5.09
+ $Y2=0
r114 69 71 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.255 $Y=0
+ $X2=5.52 $Y2=0
r115 68 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=6.03
+ $Y2=0
r116 68 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=5.52
+ $Y2=0
r117 67 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r118 67 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r119 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r120 64 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.155
+ $Y2=0
r121 64 66 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.56
+ $Y2=0
r122 63 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=0 $X2=5.09
+ $Y2=0
r123 63 66 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.925 $Y=0
+ $X2=4.56 $Y2=0
r124 62 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r125 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r126 59 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r127 58 61 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r128 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r129 56 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.085
+ $Y2=0
r130 56 58 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.64
+ $Y2=0
r131 55 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=4.155
+ $Y2=0
r132 55 61 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=3.6
+ $Y2=0
r133 54 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r134 54 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r135 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r136 51 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.225
+ $Y2=0
r137 51 53 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.68
+ $Y2=0
r138 50 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=2.085
+ $Y2=0
r139 50 53 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r140 49 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r141 49 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r142 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r143 46 79 4.57341 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.265
+ $Y2=0
r144 46 48 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.72
+ $Y2=0
r145 45 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=1.225
+ $Y2=0
r146 45 48 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=0.72
+ $Y2=0
r147 43 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r148 43 59 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.64
+ $Y2=0
r149 39 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0
r150 39 41 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0.47
r151 35 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=0.085
+ $X2=5.09 $Y2=0
r152 35 37 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.09 $Y=0.085
+ $X2=5.09 $Y2=0.565
r153 31 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=0.085
+ $X2=4.155 $Y2=0
r154 31 33 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.155 $Y=0.085
+ $X2=4.155 $Y2=0.45
r155 27 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.085 $Y2=0
r156 27 29 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.085 $Y2=0.39
r157 23 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0
r158 23 25 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0.37
r159 19 79 3.19276 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.365 $Y=0.085
+ $X2=0.265 $Y2=0
r160 19 21 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.365 $Y=0.085
+ $X2=0.365 $Y2=0.39
r161 6 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.89
+ $Y=0.325 $X2=6.03 $Y2=0.47
r162 5 37 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.325 $X2=5.09 $Y2=0.565
r163 4 33 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.015
+ $Y=0.325 $X2=4.155 $Y2=0.45
r164 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.245 $X2=2.085 $Y2=0.39
r165 2 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.245 $X2=1.225 $Y2=0.37
r166 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.24
+ $Y=0.245 $X2=0.365 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_4%A_528_65# 1 2 3 4 5 18 20 21 26 27 30 32 36
+ 38 42 46 48
r79 46 47 7.17647 $w=2.38e-07 $l=1.4e-07 $layer=LI1_cond $X=4.62 $Y=1.02
+ $X2=4.62 $Y2=1.16
r80 44 46 3.33193 $w=2.38e-07 $l=6.5e-08 $layer=LI1_cond $X=4.62 $Y=0.955
+ $X2=4.62 $Y2=1.02
r81 40 42 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=6.495 $Y=0.87
+ $X2=6.495 $Y2=0.47
r82 39 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.695 $Y=0.955
+ $X2=5.565 $Y2=0.955
r83 38 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.365 $Y=0.955
+ $X2=6.495 $Y2=0.87
r84 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.365 $Y=0.955
+ $X2=5.695 $Y2=0.955
r85 34 48 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0.87
+ $X2=5.565 $Y2=0.955
r86 34 36 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=5.565 $Y=0.87
+ $X2=5.565 $Y2=0.47
r87 33 44 2.70854 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.75 $Y=0.955
+ $X2=4.62 $Y2=0.955
r88 32 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.435 $Y=0.955
+ $X2=5.565 $Y2=0.955
r89 32 33 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.435 $Y=0.955
+ $X2=4.75 $Y2=0.955
r90 28 44 4.09839 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=0.87 $X2=4.62
+ $Y2=0.955
r91 28 30 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=4.62 $Y=0.87 $X2=4.62
+ $Y2=0.47
r92 26 47 2.70854 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.49 $Y=1.16 $X2=4.62
+ $Y2=1.16
r93 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.49 $Y=1.16
+ $X2=3.82 $Y2=1.16
r94 23 27 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.725 $Y=1.075
+ $X2=3.82 $Y2=1.16
r95 23 25 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=3.725 $Y=1.075
+ $X2=3.725 $Y2=0.47
r96 22 25 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=3.725 $Y=0.435
+ $X2=3.725 $Y2=0.47
r97 20 22 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=3.63 $Y=0.345
+ $X2=3.725 $Y2=0.435
r98 20 21 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.63 $Y=0.345
+ $X2=2.95 $Y2=0.345
r99 16 21 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.785 $Y=0.435
+ $X2=2.95 $Y2=0.345
r100 16 18 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.785 $Y=0.435
+ $X2=2.785 $Y2=0.45
r101 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.32
+ $Y=0.325 $X2=6.46 $Y2=0.47
r102 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.46
+ $Y=0.325 $X2=5.6 $Y2=0.47
r103 3 46 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.325 $X2=4.585 $Y2=1.02
r104 3 30 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.325 $X2=4.585 $Y2=0.47
r105 2 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.585
+ $Y=0.325 $X2=3.725 $Y2=0.47
r106 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.64
+ $Y=0.325 $X2=2.785 $Y2=0.45
.ends

