* File: sky130_fd_sc_lp__or2_1.spice
* Created: Wed Sep  2 10:28:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2_1.pex.spice"
.subckt sky130_fd_sc_lp__or2_1  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1001 N_A_76_367#_M1001_d N_B_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_76_367#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.105 AS=0.0588 PD=0.883333 PS=0.7 NRD=55.704 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_76_367#_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.21 PD=2.21 PS=1.76667 NRD=0 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 A_159_367# N_B_M1003_g N_A_76_367#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1113 PD=0.66 PS=1.37 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_159_367# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.125475 AS=0.0504 PD=0.9625 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_76_367#_M1004_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.376425 PD=3.05 PS=2.8875 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__or2_1.pxi.spice"
*
.ends
*
*
