* File: sky130_fd_sc_lp__and4_1.pxi.spice
* Created: Fri Aug 28 10:07:30 2020
* 
x_PM_SKY130_FD_SC_LP__AND4_1%A N_A_c_61_n N_A_M1001_g N_A_M1008_g N_A_c_64_n A A
+ A N_A_c_66_n PM_SKY130_FD_SC_LP__AND4_1%A
x_PM_SKY130_FD_SC_LP__AND4_1%B N_B_M1002_g N_B_M1003_g N_B_c_91_n N_B_c_92_n B B
+ N_B_c_94_n PM_SKY130_FD_SC_LP__AND4_1%B
x_PM_SKY130_FD_SC_LP__AND4_1%C N_C_M1006_g N_C_M1009_g N_C_c_125_n N_C_c_126_n C
+ C N_C_c_128_n PM_SKY130_FD_SC_LP__AND4_1%C
x_PM_SKY130_FD_SC_LP__AND4_1%D N_D_M1000_g N_D_M1004_g D N_D_c_154_n N_D_c_155_n
+ PM_SKY130_FD_SC_LP__AND4_1%D
x_PM_SKY130_FD_SC_LP__AND4_1%A_40_47# N_A_40_47#_M1001_s N_A_40_47#_M1008_d
+ N_A_40_47#_M1009_d N_A_40_47#_c_187_n N_A_40_47#_M1005_g N_A_40_47#_M1007_g
+ N_A_40_47#_c_189_n N_A_40_47#_c_190_n N_A_40_47#_c_204_n N_A_40_47#_c_191_n
+ N_A_40_47#_c_225_n N_A_40_47#_c_192_n N_A_40_47#_c_193_n N_A_40_47#_c_194_n
+ PM_SKY130_FD_SC_LP__AND4_1%A_40_47#
x_PM_SKY130_FD_SC_LP__AND4_1%VPWR N_VPWR_M1008_s N_VPWR_M1003_d N_VPWR_M1004_d
+ N_VPWR_c_256_n N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_259_n N_VPWR_c_260_n
+ VPWR N_VPWR_c_261_n N_VPWR_c_262_n N_VPWR_c_255_n N_VPWR_c_264_n
+ N_VPWR_c_265_n PM_SKY130_FD_SC_LP__AND4_1%VPWR
x_PM_SKY130_FD_SC_LP__AND4_1%X N_X_M1005_d N_X_M1007_d X X X X X X X N_X_c_285_n
+ PM_SKY130_FD_SC_LP__AND4_1%X
x_PM_SKY130_FD_SC_LP__AND4_1%VGND N_VGND_M1000_d N_VGND_c_304_n N_VGND_c_305_n
+ N_VGND_c_306_n VGND N_VGND_c_307_n N_VGND_c_308_n
+ PM_SKY130_FD_SC_LP__AND4_1%VGND
cc_1 VNB N_A_c_61_n 0.0265032f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.325
cc_2 VNB N_A_M1001_g 0.0278941f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.445
cc_3 VNB N_A_M1008_g 0.00964471f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.045
cc_4 VNB N_A_c_64_n 0.0228007f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_5 VNB A 0.0376049f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A_c_66_n 0.0227329f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.005
cc_7 VNB N_B_M1002_g 0.0204084f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.84
cc_8 VNB N_B_M1003_g 0.0113085f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.51
cc_9 VNB N_B_c_91_n 0.0223959f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_10 VNB N_B_c_92_n 0.0159374f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_11 VNB B 0.0107449f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_12 VNB N_B_c_94_n 0.0160705f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.005
cc_13 VNB N_C_M1006_g 0.0210347f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.84
cc_14 VNB N_C_M1009_g 0.0106714f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.51
cc_15 VNB N_C_c_125_n 0.020874f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_16 VNB N_C_c_126_n 0.0152587f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_17 VNB C 0.0113493f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_C_c_128_n 0.0153273f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.005
cc_19 VNB N_D_M1000_g 0.0506145f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.84
cc_20 VNB N_D_c_154_n 0.0279968f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_21 VNB N_D_c_155_n 0.0041508f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_A_40_47#_c_187_n 0.0207621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_40_47#_M1007_g 0.00782237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_40_47#_c_189_n 0.0145038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_40_47#_c_190_n 0.0186074f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.925
cc_26 VNB N_A_40_47#_c_191_n 0.00169411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_40_47#_c_192_n 0.00203855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_40_47#_c_193_n 0.00452698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_40_47#_c_194_n 0.0418722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_255_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB X 0.0339647f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.045
cc_32 VNB N_X_c_285_n 0.0417885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_304_n 0.00907274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_305_n 0.0677042f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.51
cc_35 VNB N_VGND_c_306_n 0.00519006f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_36 VNB N_VGND_c_307_n 0.0232649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_308_n 0.190912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_M1008_g 0.0300234f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_39 VPB A 0.00998109f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_40 VPB N_B_M1003_g 0.0245309f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.51
cc_41 VPB N_C_M1009_g 0.0246027f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.51
cc_42 VPB N_D_M1004_g 0.0263431f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.51
cc_43 VPB N_D_c_154_n 0.0066872f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_44 VPB N_D_c_155_n 0.00231123f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_45 VPB N_A_40_47#_M1007_g 0.025789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_40_47#_c_191_n 0.0199744f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_40_47#_c_192_n 0.00200322f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_40_47#_c_193_n 0.00684442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_256_n 0.0136263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_257_n 0.0677515f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_51 VPB N_VPWR_c_258_n 0.0203024f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_52 VPB N_VPWR_c_259_n 0.0508781f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=1.005
cc_53 VPB N_VPWR_c_260_n 0.0314529f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=0.925
cc_54 VPB N_VPWR_c_261_n 0.0331904f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.295
cc_55 VPB N_VPWR_c_262_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_255_n 0.116087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_264_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_265_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB X 0.0570103f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_60 N_A_M1001_g N_B_M1002_g 0.0110772f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_61 N_A_c_64_n N_B_M1003_g 0.0169449f $X=0.43 $Y=1.51 $X2=0 $Y2=0
cc_62 N_A_c_61_n N_B_c_91_n 0.0110772f $X=0.43 $Y=1.325 $X2=0 $Y2=0
cc_63 N_A_c_64_n N_B_c_92_n 0.0110772f $X=0.43 $Y=1.51 $X2=0 $Y2=0
cc_64 N_A_c_66_n N_B_c_94_n 0.0110772f $X=0.41 $Y=1.005 $X2=0 $Y2=0
cc_65 N_A_M1001_g N_A_40_47#_c_189_n 0.0155343f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_66 A N_A_40_47#_c_189_n 0.0256069f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A_c_66_n N_A_40_47#_c_189_n 0.00124355f $X=0.41 $Y=1.005 $X2=0 $Y2=0
cc_68 N_A_M1001_g N_A_40_47#_c_190_n 0.0109022f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_69 A N_A_40_47#_c_190_n 0.0666689f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_70 N_A_M1008_g N_A_40_47#_c_204_n 3.20853e-19 $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_71 N_A_M1008_g N_A_40_47#_c_193_n 0.00340199f $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_72 A N_A_40_47#_c_193_n 0.0081314f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_73 N_A_M1008_g N_VPWR_c_257_n 0.0103484f $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_74 N_A_c_64_n N_VPWR_c_257_n 8.96548e-19 $X=0.43 $Y=1.51 $X2=0 $Y2=0
cc_75 A N_VPWR_c_257_n 0.0274352f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_76 N_A_M1008_g N_VPWR_c_259_n 5.18118e-19 $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_77 N_A_M1001_g N_VGND_c_305_n 0.00363059f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_78 N_A_M1001_g N_VGND_c_308_n 0.00664499f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_79 A N_VGND_c_308_n 0.00374268f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 N_B_M1002_g N_C_M1006_g 0.0236812f $X=1.02 $Y=0.445 $X2=0 $Y2=0
cc_81 N_B_M1003_g N_C_M1009_g 0.0182893f $X=1.08 $Y=2.045 $X2=0 $Y2=0
cc_82 N_B_c_91_n N_C_c_125_n 0.0138608f $X=1.11 $Y=1.31 $X2=0 $Y2=0
cc_83 N_B_c_92_n N_C_c_126_n 0.0138608f $X=1.11 $Y=1.475 $X2=0 $Y2=0
cc_84 B C 0.0525778f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_85 N_B_c_94_n C 6.90662e-19 $X=1.11 $Y=0.97 $X2=0 $Y2=0
cc_86 B N_C_c_128_n 0.00398963f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_87 N_B_c_94_n N_C_c_128_n 0.0138608f $X=1.11 $Y=0.97 $X2=0 $Y2=0
cc_88 N_B_M1002_g N_A_40_47#_c_189_n 0.0098343f $X=1.02 $Y=0.445 $X2=0 $Y2=0
cc_89 N_B_M1002_g N_A_40_47#_c_190_n 0.009746f $X=1.02 $Y=0.445 $X2=0 $Y2=0
cc_90 N_B_M1003_g N_A_40_47#_c_190_n 0.00390272f $X=1.08 $Y=2.045 $X2=0 $Y2=0
cc_91 B N_A_40_47#_c_190_n 0.0461304f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_92 N_B_M1003_g N_A_40_47#_c_204_n 0.00228049f $X=1.08 $Y=2.045 $X2=0 $Y2=0
cc_93 N_B_M1003_g N_A_40_47#_c_191_n 0.0162292f $X=1.08 $Y=2.045 $X2=0 $Y2=0
cc_94 N_B_c_92_n N_A_40_47#_c_191_n 0.00265612f $X=1.11 $Y=1.475 $X2=0 $Y2=0
cc_95 B N_A_40_47#_c_191_n 0.0241324f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_96 N_B_c_92_n N_A_40_47#_c_193_n 6.98672e-19 $X=1.11 $Y=1.475 $X2=0 $Y2=0
cc_97 N_B_M1003_g N_VPWR_c_257_n 6.08258e-19 $X=1.08 $Y=2.045 $X2=0 $Y2=0
cc_98 N_B_M1003_g N_VPWR_c_259_n 0.00837765f $X=1.08 $Y=2.045 $X2=0 $Y2=0
cc_99 N_B_M1002_g N_VGND_c_305_n 0.00585385f $X=1.02 $Y=0.445 $X2=0 $Y2=0
cc_100 N_B_M1002_g N_VGND_c_308_n 0.00933411f $X=1.02 $Y=0.445 $X2=0 $Y2=0
cc_101 B N_VGND_c_308_n 0.0116688f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_102 N_C_M1006_g N_D_M1000_g 0.0234218f $X=1.56 $Y=0.445 $X2=0 $Y2=0
cc_103 C N_D_M1000_g 0.00946194f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_104 N_C_c_128_n N_D_M1000_g 0.0200737f $X=1.65 $Y=0.97 $X2=0 $Y2=0
cc_105 N_C_M1009_g N_D_c_154_n 0.0233804f $X=1.67 $Y=2.045 $X2=0 $Y2=0
cc_106 N_C_c_125_n N_D_c_154_n 0.0200737f $X=1.65 $Y=1.31 $X2=0 $Y2=0
cc_107 N_C_M1009_g N_D_c_155_n 0.00123666f $X=1.67 $Y=2.045 $X2=0 $Y2=0
cc_108 C N_D_c_155_n 0.00906388f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_109 N_C_M1009_g N_A_40_47#_c_191_n 0.022828f $X=1.67 $Y=2.045 $X2=0 $Y2=0
cc_110 N_C_c_126_n N_A_40_47#_c_191_n 0.0023409f $X=1.65 $Y=1.475 $X2=0 $Y2=0
cc_111 C N_A_40_47#_c_191_n 0.0241536f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_112 N_C_M1009_g N_VPWR_c_259_n 0.00759874f $X=1.67 $Y=2.045 $X2=0 $Y2=0
cc_113 C N_VGND_c_304_n 0.00926981f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_114 N_C_M1006_g N_VGND_c_305_n 0.00585385f $X=1.56 $Y=0.445 $X2=0 $Y2=0
cc_115 N_C_M1006_g N_VGND_c_308_n 0.0079575f $X=1.56 $Y=0.445 $X2=0 $Y2=0
cc_116 C N_VGND_c_308_n 0.0108752f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_117 N_D_M1000_g N_A_40_47#_c_187_n 0.0249968f $X=2.1 $Y=0.445 $X2=0 $Y2=0
cc_118 N_D_M1004_g N_A_40_47#_M1007_g 0.00971282f $X=2.1 $Y=2.045 $X2=0 $Y2=0
cc_119 N_D_c_154_n N_A_40_47#_M1007_g 0.0034065f $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_120 N_D_c_155_n N_A_40_47#_M1007_g 3.70865e-19 $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_121 N_D_c_154_n N_A_40_47#_c_191_n 0.00403636f $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_122 N_D_c_155_n N_A_40_47#_c_191_n 0.00802582f $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_123 N_D_M1004_g N_A_40_47#_c_225_n 0.0151221f $X=2.1 $Y=2.045 $X2=0 $Y2=0
cc_124 N_D_c_154_n N_A_40_47#_c_225_n 9.14836e-19 $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_125 N_D_c_155_n N_A_40_47#_c_225_n 0.0234099f $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_126 N_D_M1000_g N_A_40_47#_c_192_n 9.24595e-19 $X=2.1 $Y=0.445 $X2=0 $Y2=0
cc_127 N_D_M1004_g N_A_40_47#_c_192_n 0.00359606f $X=2.1 $Y=2.045 $X2=0 $Y2=0
cc_128 N_D_c_154_n N_A_40_47#_c_192_n 0.001934f $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_129 N_D_c_155_n N_A_40_47#_c_192_n 0.0272622f $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_130 N_D_c_154_n N_A_40_47#_c_194_n 0.0105027f $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_131 N_D_c_155_n N_A_40_47#_c_194_n 6.12358e-19 $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_132 N_D_M1004_g N_VPWR_c_260_n 0.00165223f $X=2.1 $Y=2.045 $X2=0 $Y2=0
cc_133 N_D_M1000_g N_VGND_c_304_n 0.020599f $X=2.1 $Y=0.445 $X2=0 $Y2=0
cc_134 N_D_c_154_n N_VGND_c_304_n 7.51726e-19 $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_135 N_D_c_155_n N_VGND_c_304_n 0.00532205f $X=2.19 $Y=1.51 $X2=0 $Y2=0
cc_136 N_D_M1000_g N_VGND_c_305_n 0.00585385f $X=2.1 $Y=0.445 $X2=0 $Y2=0
cc_137 N_D_M1000_g N_VGND_c_308_n 0.0114913f $X=2.1 $Y=0.445 $X2=0 $Y2=0
cc_138 N_A_40_47#_c_225_n N_VPWR_M1004_d 0.0258559f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_139 N_A_40_47#_c_192_n N_VPWR_M1004_d 0.00171986f $X=2.73 $Y=1.35 $X2=0 $Y2=0
cc_140 N_A_40_47#_c_191_n N_VPWR_c_259_n 0.0353109f $X=1.63 $Y=1.74 $X2=0 $Y2=0
cc_141 N_A_40_47#_M1007_g N_VPWR_c_260_n 0.0166953f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_40_47#_c_225_n N_VPWR_c_260_n 0.0237955f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_143 N_A_40_47#_M1007_g N_VPWR_c_262_n 0.00486043f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_40_47#_M1007_g N_VPWR_c_255_n 0.00917987f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_40_47#_c_187_n X 0.00443904f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_146 N_A_40_47#_c_192_n X 0.053229f $X=2.73 $Y=1.35 $X2=0 $Y2=0
cc_147 N_A_40_47#_c_194_n X 0.0191032f $X=2.885 $Y=1.35 $X2=0 $Y2=0
cc_148 N_A_40_47#_c_187_n N_X_c_285_n 0.011917f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_149 N_A_40_47#_c_192_n N_X_c_285_n 0.00982092f $X=2.73 $Y=1.35 $X2=0 $Y2=0
cc_150 N_A_40_47#_c_194_n N_X_c_285_n 0.00686342f $X=2.885 $Y=1.35 $X2=0 $Y2=0
cc_151 N_A_40_47#_c_189_n A_123_47# 0.00675385f $X=0.665 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_40_47#_c_190_n A_123_47# 5.88103e-19 $X=0.75 $Y=1.655 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A_40_47#_c_187_n N_VGND_c_304_n 0.00355091f $X=2.64 $Y=1.185 $X2=0
+ $Y2=0
cc_154 N_A_40_47#_c_189_n N_VGND_c_305_n 0.0358839f $X=0.665 $Y=0.445 $X2=0
+ $Y2=0
cc_155 N_A_40_47#_c_187_n N_VGND_c_307_n 0.0054895f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_156 N_A_40_47#_M1001_s N_VGND_c_308_n 0.0021695f $X=0.2 $Y=0.235 $X2=0 $Y2=0
cc_157 N_A_40_47#_c_187_n N_VGND_c_308_n 0.0111296f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_158 N_A_40_47#_c_189_n N_VGND_c_308_n 0.0248237f $X=0.665 $Y=0.445 $X2=0
+ $Y2=0
cc_159 N_VPWR_c_255_n N_X_M1007_d 0.00371702f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_c_262_n X 0.018528f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_161 N_VPWR_c_255_n X 0.0104192f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_162 N_X_c_285_n N_VGND_c_307_n 0.0393268f $X=2.855 $Y=0.385 $X2=0 $Y2=0
cc_163 N_X_M1005_d N_VGND_c_308_n 0.00215158f $X=2.715 $Y=0.235 $X2=0 $Y2=0
cc_164 N_X_c_285_n N_VGND_c_308_n 0.0224827f $X=2.855 $Y=0.385 $X2=0 $Y2=0
cc_165 A_123_47# N_VGND_c_308_n 0.00648821f $X=0.615 $Y=0.235 $X2=0.812
+ $Y2=2.045
cc_166 A_219_47# N_VGND_c_308_n 0.00956873f $X=1.095 $Y=0.235 $X2=3.12 $Y2=0
cc_167 A_327_47# N_VGND_c_308_n 0.0112904f $X=1.635 $Y=0.235 $X2=3.12 $Y2=0
