* File: sky130_fd_sc_lp__o311a_0.pex.spice
* Created: Fri Aug 28 11:13:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311A_0%A_96_161# 1 2 3 12 13 16 18 20 22 23 24 27
+ 28 30 31 34 36 39 42 44 48 50
c106 42 0 1.12907e-19 $X=3.35 $Y=2.55
c107 34 0 1.65606e-19 $X=2.405 $Y=2.55
r108 45 48 4.29547 $w=3.28e-07 $l=1.23e-07 $layer=LI1_cond $X=3.197 $Y=0.485
+ $X2=3.32 $Y2=0.485
r109 40 50 3.77418 $w=2.45e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.377 $Y=2.215
+ $X2=3.302 $Y2=2.13
r110 40 42 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=3.377 $Y=2.215
+ $X2=3.377 $Y2=2.55
r111 39 50 3.77418 $w=2.45e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.197 $Y=2.045
+ $X2=3.302 $Y2=2.13
r112 38 45 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=3.197 $Y=0.65
+ $X2=3.197 $Y2=0.485
r113 38 39 74.7748 $w=2.13e-07 $l=1.395e-06 $layer=LI1_cond $X=3.197 $Y=0.65
+ $X2=3.197 $Y2=2.045
r114 37 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=2.13
+ $X2=2.405 $Y2=2.13
r115 36 50 2.68609 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.09 $Y=2.13
+ $X2=3.302 $Y2=2.13
r116 36 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.09 $Y=2.13
+ $X2=2.57 $Y2=2.13
r117 32 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=2.215
+ $X2=2.405 $Y2=2.13
r118 32 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.405 $Y=2.215
+ $X2=2.405 $Y2=2.55
r119 30 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=2.13
+ $X2=2.405 $Y2=2.13
r120 30 31 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=2.24 $Y=2.13
+ $X2=0.855 $Y2=2.13
r121 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.645
+ $Y=1.71 $X2=0.645 $Y2=1.71
r122 25 31 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=0.702 $Y=2.045
+ $X2=0.855 $Y2=2.13
r123 25 27 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=0.702 $Y=2.045
+ $X2=0.702 $Y2=1.71
r124 23 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.645 $Y=2.05
+ $X2=0.645 $Y2=1.71
r125 23 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=2.05
+ $X2=0.645 $Y2=2.215
r126 22 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=1.545
+ $X2=0.645 $Y2=1.71
r127 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.915 $Y=0.805
+ $X2=0.915 $Y2=0.485
r128 16 24 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.735 $Y=2.725
+ $X2=0.735 $Y2=2.215
r129 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.84 $Y=0.88
+ $X2=0.915 $Y2=0.805
r130 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.84 $Y=0.88
+ $X2=0.63 $Y2=0.88
r131 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.555 $Y=0.955
+ $X2=0.63 $Y2=0.88
r132 10 22 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.555 $Y=0.955
+ $X2=0.555 $Y2=1.545
r133 3 42 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.21
+ $Y=2.405 $X2=3.35 $Y2=2.55
r134 2 34 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.25
+ $Y=2.405 $X2=2.405 $Y2=2.55
r135 1 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.18
+ $Y=0.275 $X2=3.32 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_0%A1 5 7 9 11 12 13 16 18 19 20 25 27
r57 19 20 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.192 $Y=1.295
+ $X2=1.192 $Y2=1.665
r58 19 27 4.40336 $w=3.33e-07 $l=1.28e-07 $layer=LI1_cond $X=1.192 $Y=1.295
+ $X2=1.192 $Y2=1.167
r59 19 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.185
+ $Y=1.36 $X2=1.185 $Y2=1.36
r60 18 27 8.81313 $w=3.35e-07 $l=2.42e-07 $layer=LI1_cond $X=1.192 $Y=0.925
+ $X2=1.192 $Y2=1.167
r61 14 16 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.275 $Y=0.88
+ $X2=1.385 $Y2=0.88
r62 12 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.185 $Y=1.7
+ $X2=1.185 $Y2=1.36
r63 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.7
+ $X2=1.185 $Y2=1.865
r64 11 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.195
+ $X2=1.185 $Y2=1.36
r65 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.385 $Y=0.805
+ $X2=1.385 $Y2=0.88
r66 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.385 $Y=0.805
+ $X2=1.385 $Y2=0.485
r67 5 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.275 $Y=2.725
+ $X2=1.275 $Y2=1.865
r68 1 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.275 $Y=0.955
+ $X2=1.275 $Y2=0.88
r69 1 11 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.275 $Y=0.955
+ $X2=1.275 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_0%A2 1 3 7 11 12 13 17
c46 12 0 1.10727e-19 $X=1.68 $Y=1.295
r47 12 13 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=1.295
+ $X2=1.69 $Y2=1.665
r48 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.725
+ $Y=1.36 $X2=1.725 $Y2=1.36
r49 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.725 $Y=1.7
+ $X2=1.725 $Y2=1.36
r50 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.195
+ $X2=1.725 $Y2=1.36
r51 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.815 $Y=0.485
+ $X2=1.815 $Y2=1.195
r52 1 11 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.865
+ $X2=1.725 $Y2=1.7
r53 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.725 $Y=1.865
+ $X2=1.725 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_0%A3 3 7 11 12 13 14 18 19
c44 3 0 1.10727e-19 $X=2.175 $Y=2.725
r45 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.265
+ $Y=1.245 $X2=2.265 $Y2=1.245
r46 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.185 $Y=1.295
+ $X2=2.185 $Y2=1.665
r47 13 19 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.185 $Y=1.295
+ $X2=2.185 $Y2=1.245
r48 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.265 $Y=1.585
+ $X2=2.265 $Y2=1.245
r49 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.585
+ $X2=2.265 $Y2=1.75
r50 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.08
+ $X2=2.265 $Y2=1.245
r51 7 10 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=2.315 $Y=0.485
+ $X2=2.315 $Y2=1.08
r52 3 12 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=2.175 $Y=2.725
+ $X2=2.175 $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_0%B1 3 7 9 12 13 17
c46 3 0 1.12907e-19 $X=2.635 $Y=2.725
r47 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.835
+ $Y=1.36 $X2=2.835 $Y2=1.36
r48 13 18 8.78738 $w=3.98e-07 $l=3.05e-07 $layer=LI1_cond $X=2.72 $Y=1.665
+ $X2=2.72 $Y2=1.36
r49 12 18 1.87272 $w=3.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.72 $Y=1.295
+ $X2=2.72 $Y2=1.36
r50 11 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.195
+ $X2=2.835 $Y2=1.36
r51 9 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.835 $Y=1.7
+ $X2=2.835 $Y2=1.36
r52 7 11 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.745 $Y=0.485
+ $X2=2.745 $Y2=1.195
r53 1 9 83.1686 $w=2.55e-07 $l=5.3066e-07 $layer=POLY_cond $X=2.635 $Y=2.14
+ $X2=2.835 $Y2=1.7
r54 1 3 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=2.635 $Y=2.14
+ $X2=2.635 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_0%C1 1 3 6 8 9 10 11 13 16 17 18 19 24
c44 6 0 1.65606e-19 $X=3.135 $Y=2.725
r45 18 19 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.615 $Y=1.295
+ $X2=3.615 $Y2=1.665
r46 17 18 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.615 $Y=0.925
+ $X2=3.615 $Y2=1.295
r47 17 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.005 $X2=3.57 $Y2=1.005
r48 15 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.57 $Y=1.345
+ $X2=3.57 $Y2=1.005
r49 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.345
+ $X2=3.57 $Y2=1.51
r50 14 24 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=3.57 $Y=0.955 $X2=3.57
+ $Y2=1.005
r51 13 16 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=3.48 $Y=2.105
+ $X2=3.48 $Y2=1.51
r52 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.405 $Y=2.18
+ $X2=3.48 $Y2=2.105
r53 10 11 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.405 $Y=2.18
+ $X2=3.21 $Y2=2.18
r54 8 14 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.405 $Y=0.88
+ $X2=3.57 $Y2=0.955
r55 8 9 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=3.405 $Y=0.88
+ $X2=3.18 $Y2=0.88
r56 4 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.135 $Y=2.255
+ $X2=3.21 $Y2=2.18
r57 4 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.135 $Y=2.255 $X2=3.135
+ $Y2=2.725
r58 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.105 $Y=0.805
+ $X2=3.18 $Y2=0.88
r59 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.105 $Y=0.805
+ $X2=3.105 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_0%X 1 2 9 11 12 13 14 15 16 17 26 40
r22 40 41 3.34382 $w=5.83e-07 $l=2e-08 $layer=LI1_cond $X=0.377 $Y=2.405
+ $X2=0.377 $Y2=2.385
r23 17 44 4.6003 $w=5.83e-07 $l=2.25e-07 $layer=LI1_cond $X=0.377 $Y=2.775
+ $X2=0.377 $Y2=2.55
r24 16 44 2.31037 $w=5.83e-07 $l=1.13e-07 $layer=LI1_cond $X=0.377 $Y=2.437
+ $X2=0.377 $Y2=2.55
r25 16 40 0.654265 $w=5.83e-07 $l=3.2e-08 $layer=LI1_cond $X=0.377 $Y=2.437
+ $X2=0.377 $Y2=2.405
r26 16 41 1.28917 $w=2.93e-07 $l=3.3e-08 $layer=LI1_cond $X=0.232 $Y=2.352
+ $X2=0.232 $Y2=2.385
r27 15 16 12.3839 $w=2.93e-07 $l=3.17e-07 $layer=LI1_cond $X=0.232 $Y=2.035
+ $X2=0.232 $Y2=2.352
r28 14 15 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.232 $Y=1.665
+ $X2=0.232 $Y2=2.035
r29 13 14 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.232 $Y=1.295
+ $X2=0.232 $Y2=1.665
r30 12 13 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.232 $Y=0.925
+ $X2=0.232 $Y2=1.295
r31 12 26 10.7431 $w=2.93e-07 $l=2.75e-07 $layer=LI1_cond $X=0.232 $Y=0.925
+ $X2=0.232 $Y2=0.65
r32 11 26 3.60803 $w=2.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.232 $Y=0.485
+ $X2=0.232 $Y2=0.65
r33 7 11 3.2363 $w=3.3e-07 $l=1.48e-07 $layer=LI1_cond $X=0.38 $Y=0.485
+ $X2=0.232 $Y2=0.485
r34 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.38 $Y=0.485 $X2=0.7
+ $Y2=0.485
r35 2 44 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.395
+ $Y=2.405 $X2=0.52 $Y2=2.55
r36 1 9 91 $w=1.7e-07 $l=5.60245e-07 $layer=licon1_NDIFF $count=2 $X=0.235
+ $Y=0.275 $X2=0.7 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_0%VPWR 1 2 9 13 16 17 19 20 21 34 35
r38 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r39 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r40 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 21 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 21 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 19 31 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.74 $Y=3.33 $X2=2.64
+ $Y2=3.33
r48 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.905 $Y2=3.33
r49 18 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.07 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=3.33
+ $X2=2.905 $Y2=3.33
r51 16 24 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.84 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.84 $Y=3.33
+ $X2=1.005 $Y2=3.33
r53 15 28 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.17 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=3.33
+ $X2=1.005 $Y2=3.33
r55 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=3.33
r56 11 13 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=2.56
r57 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.005 $Y=3.245
+ $X2=1.005 $Y2=3.33
r58 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.005 $Y=3.245
+ $X2=1.005 $Y2=2.55
r59 2 13 300 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=2 $X=2.71
+ $Y=2.405 $X2=2.905 $Y2=2.56
r60 1 9 300 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=2 $X=0.81
+ $Y=2.405 $X2=1.005 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_0%VGND 1 2 9 13 15 17 22 29 30 33 36
r47 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 30 37 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r50 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.03
+ $Y2=0
r52 27 29 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.195 $Y=0 $X2=3.6
+ $Y2=0
r53 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=1.15
+ $Y2=0
r56 23 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=1.68
+ $Y2=0
r57 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.03
+ $Y2=0
r58 22 25 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.68
+ $Y2=0
r59 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r60 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.15
+ $Y2=0
r62 17 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r63 15 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r64 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r65 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0
r66 11 13 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0.465
r67 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085 $X2=1.15
+ $Y2=0
r68 7 9 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=1.15 $Y=0.085 $X2=1.15
+ $Y2=0.485
r69 2 13 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.275 $X2=2.03 $Y2=0.465
r70 1 9 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.275 $X2=1.15 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_0%A_292_55# 1 2 9 11 12 15
r33 13 15 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.53 $Y=0.74
+ $X2=2.53 $Y2=0.485
r34 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.365 $Y=0.825
+ $X2=2.53 $Y2=0.74
r35 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.365 $Y=0.825
+ $X2=1.695 $Y2=0.825
r36 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.6 $Y=0.74
+ $X2=1.695 $Y2=0.825
r37 7 9 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=1.6 $Y=0.74 $X2=1.6
+ $Y2=0.485
r38 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.275 $X2=2.53 $Y2=0.485
r39 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.46
+ $Y=0.275 $X2=1.6 $Y2=0.485
.ends

