* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
X0 VGND a_27_465# a_196_465# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_614_93# a_486_119# a_857_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND D a_400_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1855_47# a_1158_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_400_119# a_196_465# a_486_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_486_119# a_196_465# a_572_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_857_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 Q a_1855_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR D a_400_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR a_486_119# a_614_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_614_93# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_27_465# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1086_47# a_196_465# a_1158_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 a_486_119# a_27_465# a_572_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_572_463# a_614_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VPWR SET_B a_1158_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 Q a_1855_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_1339_91# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_1158_47# a_1309_65# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_1855_47# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_1095_425# a_1309_65# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VPWR a_1158_47# a_1309_65# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_1855_47# a_1158_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_1267_91# a_1309_65# a_1339_91# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_1158_47# a_27_465# a_988_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 VGND a_486_119# a_1086_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 VPWR a_486_119# a_988_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 a_1095_425# a_196_465# a_1158_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 VPWR a_27_465# a_196_465# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_400_119# a_27_465# a_486_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_1158_47# a_27_465# a_1267_91# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_572_119# a_614_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VPWR a_1855_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 a_27_465# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
