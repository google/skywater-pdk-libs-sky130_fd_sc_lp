* File: sky130_fd_sc_lp__dfxtp_lp.pxi.spice
* Created: Wed Sep  2 09:45:28 2020
* 
x_PM_SKY130_FD_SC_LP__DFXTP_LP%CLK N_CLK_M1026_g N_CLK_M1003_g N_CLK_M1020_g
+ N_CLK_c_195_n N_CLK_c_199_n CLK CLK N_CLK_c_197_n
+ PM_SKY130_FD_SC_LP__DFXTP_LP%CLK
x_PM_SKY130_FD_SC_LP__DFXTP_LP%D N_D_M1011_g N_D_c_237_n N_D_c_238_n N_D_M1022_g
+ N_D_c_240_n N_D_M1004_g D D N_D_c_242_n N_D_c_243_n
+ PM_SKY130_FD_SC_LP__DFXTP_LP%D
x_PM_SKY130_FD_SC_LP__DFXTP_LP%A_263_409# N_A_263_409#_M1000_d
+ N_A_263_409#_M1019_d N_A_263_409#_c_297_n N_A_263_409#_M1010_g
+ N_A_263_409#_c_280_n N_A_263_409#_M1024_g N_A_263_409#_M1006_g
+ N_A_263_409#_c_298_n N_A_263_409#_M1023_g N_A_263_409#_c_282_n
+ N_A_263_409#_c_283_n N_A_263_409#_c_284_n N_A_263_409#_c_302_n
+ N_A_263_409#_c_285_n N_A_263_409#_c_304_n N_A_263_409#_c_317_n
+ N_A_263_409#_c_286_n N_A_263_409#_c_287_n N_A_263_409#_c_288_n
+ N_A_263_409#_c_289_n N_A_263_409#_c_290_n N_A_263_409#_c_347_p
+ N_A_263_409#_c_343_p N_A_263_409#_c_371_p N_A_263_409#_c_291_n
+ N_A_263_409#_c_292_n N_A_263_409#_c_341_p N_A_263_409#_c_306_n
+ N_A_263_409#_c_307_n N_A_263_409#_c_293_n N_A_263_409#_c_308_n
+ N_A_263_409#_c_294_n N_A_263_409#_c_295_n N_A_263_409#_c_296_n
+ PM_SKY130_FD_SC_LP__DFXTP_LP%A_263_409#
x_PM_SKY130_FD_SC_LP__DFXTP_LP%A_1005_99# N_A_1005_99#_M1018_d
+ N_A_1005_99#_M1015_d N_A_1005_99#_c_472_n N_A_1005_99#_M1029_g
+ N_A_1005_99#_M1016_g N_A_1005_99#_c_474_n N_A_1005_99#_c_475_n
+ N_A_1005_99#_c_509_p N_A_1005_99#_c_518_p N_A_1005_99#_c_481_n
+ N_A_1005_99#_c_482_n N_A_1005_99#_c_476_n N_A_1005_99#_c_477_n
+ N_A_1005_99#_c_484_n N_A_1005_99#_c_478_n
+ PM_SKY130_FD_SC_LP__DFXTP_LP%A_1005_99#
x_PM_SKY130_FD_SC_LP__DFXTP_LP%A_747_79# N_A_747_79#_M1013_d N_A_747_79#_M1010_d
+ N_A_747_79#_M1015_g N_A_747_79#_M1021_g N_A_747_79#_c_578_n
+ N_A_747_79#_M1018_g N_A_747_79#_c_580_n N_A_747_79#_c_581_n
+ N_A_747_79#_c_589_n N_A_747_79#_c_590_n N_A_747_79#_c_582_n
+ N_A_747_79#_c_618_n N_A_747_79#_c_621_n N_A_747_79#_c_583_n
+ N_A_747_79#_c_584_n N_A_747_79#_c_585_n N_A_747_79#_c_594_n
+ N_A_747_79#_c_586_n PM_SKY130_FD_SC_LP__DFXTP_LP%A_747_79#
x_PM_SKY130_FD_SC_LP__DFXTP_LP%A_27_57# N_A_27_57#_M1026_s N_A_27_57#_M1003_s
+ N_A_27_57#_M1019_g N_A_27_57#_c_701_n N_A_27_57#_M1028_g N_A_27_57#_c_702_n
+ N_A_27_57#_M1000_g N_A_27_57#_c_703_n N_A_27_57#_c_704_n N_A_27_57#_c_705_n
+ N_A_27_57#_c_706_n N_A_27_57#_c_723_n N_A_27_57#_c_724_n N_A_27_57#_c_707_n
+ N_A_27_57#_c_708_n N_A_27_57#_M1013_g N_A_27_57#_c_710_n N_A_27_57#_M1007_g
+ N_A_27_57#_c_726_n N_A_27_57#_M1008_g N_A_27_57#_c_711_n N_A_27_57#_M1001_g
+ N_A_27_57#_c_712_n N_A_27_57#_c_713_n N_A_27_57#_c_714_n N_A_27_57#_c_729_n
+ N_A_27_57#_c_715_n N_A_27_57#_c_730_n N_A_27_57#_c_716_n N_A_27_57#_c_717_n
+ N_A_27_57#_c_731_n N_A_27_57#_c_718_n N_A_27_57#_c_719_n N_A_27_57#_c_720_n
+ PM_SKY130_FD_SC_LP__DFXTP_LP%A_27_57#
x_PM_SKY130_FD_SC_LP__DFXTP_LP%A_1583_285# N_A_1583_285#_M1014_d
+ N_A_1583_285#_M1017_d N_A_1583_285#_M1005_g N_A_1583_285#_M1002_g
+ N_A_1583_285#_M1009_g N_A_1583_285#_c_878_n N_A_1583_285#_M1027_g
+ N_A_1583_285#_M1025_g N_A_1583_285#_c_880_n N_A_1583_285#_c_881_n
+ N_A_1583_285#_c_882_n N_A_1583_285#_c_893_n N_A_1583_285#_c_894_n
+ N_A_1583_285#_c_883_n N_A_1583_285#_c_896_n N_A_1583_285#_c_884_n
+ N_A_1583_285#_c_885_n N_A_1583_285#_c_886_n N_A_1583_285#_c_887_n
+ PM_SKY130_FD_SC_LP__DFXTP_LP%A_1583_285#
x_PM_SKY130_FD_SC_LP__DFXTP_LP%A_1429_383# N_A_1429_383#_M1006_d
+ N_A_1429_383#_M1008_d N_A_1429_383#_c_987_n N_A_1429_383#_M1012_g
+ N_A_1429_383#_M1017_g N_A_1429_383#_c_989_n N_A_1429_383#_M1014_g
+ N_A_1429_383#_c_990_n N_A_1429_383#_c_991_n N_A_1429_383#_c_1002_n
+ N_A_1429_383#_c_992_n N_A_1429_383#_c_993_n N_A_1429_383#_c_994_n
+ N_A_1429_383#_c_995_n N_A_1429_383#_c_1001_n N_A_1429_383#_c_996_n
+ N_A_1429_383#_c_997_n N_A_1429_383#_c_998_n
+ PM_SKY130_FD_SC_LP__DFXTP_LP%A_1429_383#
x_PM_SKY130_FD_SC_LP__DFXTP_LP%VPWR N_VPWR_M1003_d N_VPWR_M1022_s N_VPWR_M1016_d
+ N_VPWR_M1005_d N_VPWR_M1027_s N_VPWR_c_1082_n N_VPWR_c_1083_n N_VPWR_c_1084_n
+ N_VPWR_c_1085_n N_VPWR_c_1086_n N_VPWR_c_1087_n N_VPWR_c_1088_n
+ N_VPWR_c_1089_n N_VPWR_c_1090_n N_VPWR_c_1091_n N_VPWR_c_1092_n VPWR
+ N_VPWR_c_1093_n N_VPWR_c_1094_n N_VPWR_c_1095_n N_VPWR_c_1081_n
+ N_VPWR_c_1097_n N_VPWR_c_1098_n PM_SKY130_FD_SC_LP__DFXTP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DFXTP_LP%A_629_125# N_A_629_125#_M1004_d
+ N_A_629_125#_M1022_d N_A_629_125#_c_1173_n N_A_629_125#_c_1174_n
+ N_A_629_125#_c_1185_n N_A_629_125#_c_1187_n N_A_629_125#_c_1175_n
+ N_A_629_125#_c_1177_n PM_SKY130_FD_SC_LP__DFXTP_LP%A_629_125#
x_PM_SKY130_FD_SC_LP__DFXTP_LP%Q N_Q_M1025_d N_Q_M1027_d N_Q_c_1219_n Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DFXTP_LP%Q
x_PM_SKY130_FD_SC_LP__DFXTP_LP%VGND N_VGND_M1020_d N_VGND_M1011_s N_VGND_M1029_d
+ N_VGND_M1002_d N_VGND_M1009_s N_VGND_c_1235_n N_VGND_c_1236_n N_VGND_c_1237_n
+ N_VGND_c_1238_n N_VGND_c_1239_n N_VGND_c_1240_n N_VGND_c_1241_n
+ N_VGND_c_1242_n N_VGND_c_1243_n N_VGND_c_1244_n N_VGND_c_1245_n VGND
+ N_VGND_c_1246_n N_VGND_c_1247_n N_VGND_c_1248_n N_VGND_c_1249_n
+ N_VGND_c_1250_n N_VGND_c_1251_n PM_SKY130_FD_SC_LP__DFXTP_LP%VGND
cc_1 VNB N_CLK_M1026_g 0.0401047f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.495
cc_2 VNB N_CLK_M1020_g 0.0311126f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.495
cc_3 VNB N_CLK_c_195_n 0.0200671f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.325
cc_4 VNB CLK 0.00355077f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_CLK_c_197_n 0.0262488f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.34
cc_6 VNB N_D_c_237_n 0.0137423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_D_c_238_n 0.0130666f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.545
cc_8 VNB N_D_M1022_g 0.00489859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_D_c_240_n 0.018249f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.495
cc_10 VNB D 0.0075588f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.325
cc_11 VNB N_D_c_242_n 0.0298543f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_D_c_243_n 0.0161112f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_13 VNB N_A_263_409#_c_280_n 0.0186468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_263_409#_M1006_g 0.020198f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.845
cc_15 VNB N_A_263_409#_c_282_n 0.0322051f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.34
cc_16 VNB N_A_263_409#_c_283_n 0.0137588f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.295
cc_17 VNB N_A_263_409#_c_284_n 0.00876374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_263_409#_c_285_n 0.0146787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_263_409#_c_286_n 0.00379913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_263_409#_c_287_n 0.00273328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_263_409#_c_288_n 0.0412288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_263_409#_c_289_n 0.0298899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_263_409#_c_290_n 0.0035809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_263_409#_c_291_n 0.00580575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_263_409#_c_292_n 0.00794802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_263_409#_c_293_n 0.00869099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_263_409#_c_294_n 0.0028787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_263_409#_c_295_n 0.0350401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_263_409#_c_296_n 0.0246096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_1005_99#_c_472_n 0.0170623f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.545
cc_31 VNB N_A_1005_99#_M1016_g 0.002789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1005_99#_c_474_n 0.00214839f $X=-0.19 $Y=-0.245 $X2=0.597
+ $Y2=1.658
cc_33 VNB N_A_1005_99#_c_475_n 0.0463968f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.845
cc_34 VNB N_A_1005_99#_c_476_n 0.00235241f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.665
cc_35 VNB N_A_1005_99#_c_477_n 0.00835771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1005_99#_c_478_n 0.00246454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_747_79#_M1021_g 0.019397f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.325
cc_38 VNB N_A_747_79#_c_578_n 0.0163505f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.325
cc_39 VNB N_A_747_79#_M1018_g 0.0175204f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_40 VNB N_A_747_79#_c_580_n 0.0110756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_747_79#_c_581_n 0.00475669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_747_79#_c_582_n 0.00349723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_747_79#_c_583_n 0.00826115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_747_79#_c_584_n 0.00385312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_747_79#_c_585_n 0.00347665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_747_79#_c_586_n 0.0525283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_57#_c_701_n 0.0138897f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.495
cc_48 VNB N_A_27_57#_c_702_n 0.0142205f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.175
cc_49 VNB N_A_27_57#_c_703_n 0.0153367f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.845
cc_50 VNB N_A_27_57#_c_704_n 0.0187753f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_51 VNB N_A_27_57#_c_705_n 0.046708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_57#_c_706_n 0.0297998f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.34
cc_53 VNB N_A_27_57#_c_707_n 0.101455f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.295
cc_54 VNB N_A_27_57#_c_708_n 0.0108465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_57#_M1013_g 0.0241653f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.665
cc_56 VNB N_A_27_57#_c_710_n 0.320335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_57#_c_711_n 0.0197745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_27_57#_c_712_n 0.0337213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_27_57#_c_713_n 0.0085541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_57#_c_714_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_27_57#_c_715_n 0.0241735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_27_57#_c_716_n 0.0139302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_27_57#_c_717_n 0.0132078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_27_57#_c_718_n 0.0308667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_27_57#_c_719_n 0.00322439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_27_57#_c_720_n 0.0301745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1583_285#_M1002_g 0.0502818f $X=-0.19 $Y=-0.245 $X2=0.597
+ $Y2=1.325
cc_68 VNB N_A_1583_285#_M1009_g 0.0233224f $X=-0.19 $Y=-0.245 $X2=0.597
+ $Y2=1.845
cc_69 VNB N_A_1583_285#_c_878_n 0.0687563f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_70 VNB N_A_1583_285#_M1025_g 0.025778f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.295
cc_71 VNB N_A_1583_285#_c_880_n 0.0299455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1583_285#_c_881_n 0.00314316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1583_285#_c_882_n 0.0217309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1583_285#_c_883_n 0.00147606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1583_285#_c_884_n 0.0180161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1583_285#_c_885_n 0.0129399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1583_285#_c_886_n 0.00154761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1583_285#_c_887_n 0.0088611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1429_383#_c_987_n 0.0158609f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.545
cc_80 VNB N_A_1429_383#_M1017_g 0.00539552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1429_383#_c_989_n 0.0187347f $X=-0.19 $Y=-0.245 $X2=0.665
+ $Y2=1.175
cc_82 VNB N_A_1429_383#_c_990_n 0.0277629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1429_383#_c_991_n 0.0159273f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.34
cc_84 VNB N_A_1429_383#_c_992_n 0.0109858f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.665
cc_85 VNB N_A_1429_383#_c_993_n 0.0015015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1429_383#_c_994_n 0.00191479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1429_383#_c_995_n 0.0100051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1429_383#_c_996_n 0.00132384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1429_383#_c_997_n 0.00135938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1429_383#_c_998_n 0.0323368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VPWR_c_1081_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_629_125#_c_1173_n 0.00606688f $X=-0.19 $Y=-0.245 $X2=0.845
+ $Y2=1.175
cc_93 VNB N_A_629_125#_c_1174_n 0.00794022f $X=-0.19 $Y=-0.245 $X2=0.597
+ $Y2=1.325
cc_94 VNB N_A_629_125#_c_1175_n 0.00323625f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_95 VNB Q 0.0507138f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.325
cc_96 VNB Q 0.00190626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1235_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_98 VNB N_VGND_c_1236_n 0.0135924f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.34
cc_99 VNB N_VGND_c_1237_n 0.0148052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1238_n 0.00761282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1239_n 0.018831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1240_n 0.0279894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1241_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1242_n 0.0549356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1243_n 0.00465705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1244_n 0.0312589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1245_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1246_n 0.0268803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1247_n 0.0991336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1248_n 0.0284113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1249_n 0.561577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1250_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1251_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VPB N_CLK_M1003_g 0.0333343f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.545
cc_115 VPB N_CLK_c_199_n 0.0178939f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.845
cc_116 VPB CLK 0.00332822f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_117 VPB N_D_M1022_g 0.0334668f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_263_409#_c_297_n 0.0153912f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.545
cc_119 VPB N_A_263_409#_c_298_n 0.0226933f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_120 VPB N_A_263_409#_c_282_n 0.0132369f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.34
cc_121 VPB N_A_263_409#_c_283_n 0.0133424f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.295
cc_122 VPB N_A_263_409#_c_284_n 0.008289f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_263_409#_c_302_n 0.0192203f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.665
cc_124 VPB N_A_263_409#_c_285_n 6.21236e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_263_409#_c_304_n 0.0321037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_263_409#_c_286_n 0.00504514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_263_409#_c_306_n 0.0150331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_263_409#_c_307_n 0.00447808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_263_409#_c_308_n 0.00314937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_1005_99#_M1016_g 0.0280963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_1005_99#_c_474_n 0.00569789f $X=-0.19 $Y=1.655 $X2=0.597
+ $Y2=1.658
cc_132 VPB N_A_1005_99#_c_481_n 0.00771539f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.34
cc_133 VPB N_A_1005_99#_c_482_n 0.0183005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_1005_99#_c_477_n 6.57884e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_1005_99#_c_484_n 0.00336798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_747_79#_M1015_g 0.0345403f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.175
cc_137 VPB N_A_747_79#_c_581_n 0.00406359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_747_79#_c_589_n 0.00553273f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.665
cc_139 VPB N_A_747_79#_c_590_n 0.0104471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_747_79#_c_582_n 0.00312116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_747_79#_c_584_n 0.00187626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_747_79#_c_585_n 0.00200047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_747_79#_c_594_n 0.00214867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_747_79#_c_586_n 0.0155786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_27_57#_M1019_g 0.0431597f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.175
cc_146 VPB N_A_27_57#_c_705_n 0.104069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_27_57#_c_723_n 0.188308f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.34
cc_148 VPB N_A_27_57#_c_724_n 0.0117286f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.34
cc_149 VPB N_A_27_57#_M1007_g 0.0339985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_27_57#_c_726_n 0.181435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_27_57#_M1008_g 0.0278573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_27_57#_c_712_n 0.00263085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_27_57#_c_729_n 0.0124845f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_27_57#_c_730_n 0.0390561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_27_57#_c_731_n 0.0166056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_27_57#_c_718_n 0.0177642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_1583_285#_M1005_g 0.0256808f $X=-0.19 $Y=1.655 $X2=0.845
+ $Y2=1.175
cc_158 VPB N_A_1583_285#_c_878_n 0.0194947f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_159 VPB N_A_1583_285#_M1027_g 0.0405981f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_1583_285#_c_880_n 0.0201029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_1583_285#_c_882_n 0.0166473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_1583_285#_c_893_n 0.00384933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_1583_285#_c_894_n 0.00111311f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_1583_285#_c_883_n 0.0122877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_1583_285#_c_896_n 0.0144339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_1583_285#_c_885_n 0.0155455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_1429_383#_M1017_g 0.0392545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_1429_383#_c_994_n 0.00248067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_1429_383#_c_1001_n 0.00259127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1082_n 0.00962351f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_171 VPB N_VPWR_c_1083_n 0.026784f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.34
cc_172 VPB N_VPWR_c_1084_n 0.0156306f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.34
cc_173 VPB N_VPWR_c_1085_n 0.0140465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1086_n 0.0254412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1087_n 0.0214312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1088_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1089_n 0.0847316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1090_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1091_n 0.035777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1092_n 0.00598038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1093_n 0.0392121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1094_n 0.0734295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1095_n 0.0197141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1081_n 0.131068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1097_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1098_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_629_125#_c_1175_n 0.00231859f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.21
cc_188 VPB N_A_629_125#_c_1177_n 0.00348922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_Q_c_1219_n 0.0496579f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.175
cc_190 VPB Q 0.00566171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 N_CLK_M1003_g N_A_263_409#_c_306_n 2.75279e-19 $X=0.66 $Y=2.545 $X2=0
+ $Y2=0
cc_192 N_CLK_c_199_n N_A_27_57#_M1019_g 0.0142859f $X=0.597 $Y=1.845 $X2=0 $Y2=0
cc_193 N_CLK_M1020_g N_A_27_57#_c_701_n 0.0124312f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_194 N_CLK_M1020_g N_A_27_57#_c_704_n 0.0148988f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_195 CLK N_A_27_57#_c_712_n 0.00640943f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_196 N_CLK_c_197_n N_A_27_57#_c_712_n 0.0142859f $X=0.62 $Y=1.34 $X2=0 $Y2=0
cc_197 N_CLK_M1026_g N_A_27_57#_c_715_n 0.01276f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_198 N_CLK_M1020_g N_A_27_57#_c_715_n 0.00193397f $X=0.845 $Y=0.495 $X2=0
+ $Y2=0
cc_199 N_CLK_M1003_g N_A_27_57#_c_730_n 0.0143689f $X=0.66 $Y=2.545 $X2=0 $Y2=0
cc_200 N_CLK_M1026_g N_A_27_57#_c_716_n 0.0086968f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_201 N_CLK_M1020_g N_A_27_57#_c_716_n 0.0132282f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_202 N_CLK_c_195_n N_A_27_57#_c_716_n 2.06137e-19 $X=0.665 $Y=1.325 $X2=0
+ $Y2=0
cc_203 CLK N_A_27_57#_c_716_n 0.0282577f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_204 N_CLK_M1026_g N_A_27_57#_c_717_n 0.00513266f $X=0.485 $Y=0.495 $X2=0
+ $Y2=0
cc_205 N_CLK_M1003_g N_A_27_57#_c_731_n 0.00462174f $X=0.66 $Y=2.545 $X2=0 $Y2=0
cc_206 N_CLK_c_199_n N_A_27_57#_c_731_n 0.00281522f $X=0.597 $Y=1.845 $X2=0
+ $Y2=0
cc_207 CLK N_A_27_57#_c_731_n 0.00867382f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_208 N_CLK_M1026_g N_A_27_57#_c_718_n 0.0209089f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_209 N_CLK_M1003_g N_A_27_57#_c_718_n 0.00427061f $X=0.66 $Y=2.545 $X2=0 $Y2=0
cc_210 CLK N_A_27_57#_c_718_n 0.0486798f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_211 N_CLK_M1020_g N_A_27_57#_c_719_n 0.00178879f $X=0.845 $Y=0.495 $X2=0
+ $Y2=0
cc_212 CLK N_A_27_57#_c_719_n 0.0149817f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_213 N_CLK_c_195_n N_A_27_57#_c_720_n 0.0148988f $X=0.665 $Y=1.325 $X2=0 $Y2=0
cc_214 CLK N_A_27_57#_c_720_n 0.00320817f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_215 N_CLK_c_197_n N_A_27_57#_c_720_n 0.00690315f $X=0.62 $Y=1.34 $X2=0 $Y2=0
cc_216 N_CLK_M1003_g N_VPWR_c_1082_n 0.0237294f $X=0.66 $Y=2.545 $X2=0 $Y2=0
cc_217 N_CLK_c_195_n N_VPWR_c_1082_n 0.00255475f $X=0.665 $Y=1.325 $X2=0 $Y2=0
cc_218 CLK N_VPWR_c_1082_n 0.00634012f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_219 N_CLK_M1003_g N_VPWR_c_1087_n 0.00769046f $X=0.66 $Y=2.545 $X2=0 $Y2=0
cc_220 N_CLK_M1003_g N_VPWR_c_1081_n 0.014145f $X=0.66 $Y=2.545 $X2=0 $Y2=0
cc_221 N_CLK_M1026_g N_VGND_c_1235_n 0.00189426f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_222 N_CLK_M1020_g N_VGND_c_1235_n 0.0106455f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_223 N_CLK_M1026_g N_VGND_c_1246_n 0.00502664f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_224 N_CLK_M1020_g N_VGND_c_1246_n 0.00445056f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_225 N_CLK_M1026_g N_VGND_c_1249_n 0.00627191f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_226 N_CLK_M1020_g N_VGND_c_1249_n 0.0041956f $X=0.845 $Y=0.495 $X2=0 $Y2=0
cc_227 N_D_c_238_n N_A_263_409#_c_282_n 0.0224727f $X=3.05 $Y=1.445 $X2=0 $Y2=0
cc_228 N_D_M1022_g N_A_263_409#_c_283_n 0.0140606f $X=3.05 $Y=2.205 $X2=0 $Y2=0
cc_229 D N_A_263_409#_c_285_n 0.0232511f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_230 N_D_c_237_n N_A_263_409#_c_304_n 0.00533043f $X=2.925 $Y=1.245 $X2=0
+ $Y2=0
cc_231 N_D_M1022_g N_A_263_409#_c_304_n 0.00618396f $X=3.05 $Y=2.205 $X2=0 $Y2=0
cc_232 D N_A_263_409#_c_304_n 0.0519007f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_233 N_D_c_242_n N_A_263_409#_c_304_n 0.00793591f $X=2.55 $Y=1.245 $X2=0 $Y2=0
cc_234 N_D_c_238_n N_A_263_409#_c_317_n 0.0150388f $X=3.05 $Y=1.445 $X2=0 $Y2=0
cc_235 N_D_M1022_g N_A_263_409#_c_317_n 0.0304437f $X=3.05 $Y=2.205 $X2=0 $Y2=0
cc_236 D N_A_263_409#_c_317_n 0.0215211f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_237 N_D_c_242_n N_A_263_409#_c_317_n 2.04324e-19 $X=2.55 $Y=1.245 $X2=0 $Y2=0
cc_238 N_D_c_238_n N_A_263_409#_c_286_n 0.00688747f $X=3.05 $Y=1.445 $X2=0 $Y2=0
cc_239 N_D_M1022_g N_A_263_409#_c_286_n 0.00545839f $X=3.05 $Y=2.205 $X2=0 $Y2=0
cc_240 D N_A_27_57#_c_705_n 0.0148604f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_241 N_D_c_242_n N_A_27_57#_c_705_n 0.0181297f $X=2.55 $Y=1.245 $X2=0 $Y2=0
cc_242 N_D_c_243_n N_A_27_57#_c_705_n 0.00686713f $X=2.55 $Y=1.17 $X2=0 $Y2=0
cc_243 N_D_c_243_n N_A_27_57#_c_706_n 0.00797257f $X=2.55 $Y=1.17 $X2=0 $Y2=0
cc_244 N_D_M1022_g N_A_27_57#_c_723_n 0.0151223f $X=3.05 $Y=2.205 $X2=0 $Y2=0
cc_245 N_D_c_240_n N_A_27_57#_c_707_n 0.00907339f $X=3.07 $Y=1.17 $X2=0 $Y2=0
cc_246 N_D_c_243_n N_A_27_57#_c_707_n 0.00894529f $X=2.55 $Y=1.17 $X2=0 $Y2=0
cc_247 N_D_c_240_n N_A_27_57#_M1013_g 0.00819347f $X=3.07 $Y=1.17 $X2=0 $Y2=0
cc_248 D N_A_27_57#_c_713_n 0.00267488f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_249 N_D_M1022_g N_VPWR_c_1083_n 0.0198996f $X=3.05 $Y=2.205 $X2=0 $Y2=0
cc_250 N_D_M1022_g N_VPWR_c_1081_n 0.00158331f $X=3.05 $Y=2.205 $X2=0 $Y2=0
cc_251 N_D_c_240_n N_A_629_125#_c_1173_n 0.00352454f $X=3.07 $Y=1.17 $X2=0 $Y2=0
cc_252 N_D_c_238_n N_A_629_125#_c_1175_n 2.22996e-19 $X=3.05 $Y=1.445 $X2=0
+ $Y2=0
cc_253 N_D_M1022_g N_A_629_125#_c_1175_n 0.00232626f $X=3.05 $Y=2.205 $X2=0
+ $Y2=0
cc_254 N_D_c_240_n N_A_629_125#_c_1175_n 0.00308228f $X=3.07 $Y=1.17 $X2=0 $Y2=0
cc_255 N_D_M1022_g N_A_629_125#_c_1177_n 0.0179112f $X=3.05 $Y=2.205 $X2=0 $Y2=0
cc_256 N_D_c_240_n N_VGND_c_1236_n 0.00150476f $X=3.07 $Y=1.17 $X2=0 $Y2=0
cc_257 D N_VGND_c_1236_n 0.0239126f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_258 N_D_c_242_n N_VGND_c_1236_n 0.00399301f $X=2.55 $Y=1.245 $X2=0 $Y2=0
cc_259 N_D_c_243_n N_VGND_c_1236_n 0.0114207f $X=2.55 $Y=1.17 $X2=0 $Y2=0
cc_260 N_D_c_240_n N_VGND_c_1249_n 9.49986e-19 $X=3.07 $Y=1.17 $X2=0 $Y2=0
cc_261 N_D_c_243_n N_VGND_c_1249_n 7.97988e-19 $X=2.55 $Y=1.17 $X2=0 $Y2=0
cc_262 N_A_263_409#_c_280_n N_A_1005_99#_c_472_n 0.0102575f $X=4.435 $Y=1.155
+ $X2=0 $Y2=0
cc_263 N_A_263_409#_c_287_n N_A_1005_99#_c_472_n 0.00451739f $X=4.62 $Y=1.32
+ $X2=0 $Y2=0
cc_264 N_A_263_409#_c_289_n N_A_1005_99#_c_472_n 0.00974601f $X=5.97 $Y=0.54
+ $X2=0 $Y2=0
cc_265 N_A_263_409#_c_287_n N_A_1005_99#_c_475_n 2.97114e-19 $X=4.62 $Y=1.32
+ $X2=0 $Y2=0
cc_266 N_A_263_409#_c_288_n N_A_1005_99#_c_475_n 0.0179067f $X=4.62 $Y=1.32
+ $X2=0 $Y2=0
cc_267 N_A_263_409#_c_298_n N_A_1005_99#_c_482_n 0.00887905f $X=7.55 $Y=1.91
+ $X2=0 $Y2=0
cc_268 N_A_263_409#_c_284_n N_A_1005_99#_c_482_n 0.0054989f $X=7.55 $Y=1.785
+ $X2=0 $Y2=0
cc_269 N_A_263_409#_c_292_n N_A_1005_99#_c_482_n 0.0235112f $X=7.345 $Y=1.3
+ $X2=0 $Y2=0
cc_270 N_A_263_409#_c_294_n N_A_1005_99#_c_482_n 0.0217892f $X=7.5 $Y=1.3 $X2=0
+ $Y2=0
cc_271 N_A_263_409#_c_295_n N_A_1005_99#_c_482_n 8.54265e-19 $X=7.51 $Y=1.38
+ $X2=0 $Y2=0
cc_272 N_A_263_409#_M1006_g N_A_1005_99#_c_476_n 0.0101368f $X=7.5 $Y=0.835
+ $X2=0 $Y2=0
cc_273 N_A_263_409#_c_294_n N_A_1005_99#_c_476_n 0.0125273f $X=7.5 $Y=1.3 $X2=0
+ $Y2=0
cc_274 N_A_263_409#_c_295_n N_A_1005_99#_c_476_n 0.00127654f $X=7.51 $Y=1.38
+ $X2=0 $Y2=0
cc_275 N_A_263_409#_M1006_g N_A_1005_99#_c_477_n 0.00556462f $X=7.5 $Y=0.835
+ $X2=0 $Y2=0
cc_276 N_A_263_409#_c_294_n N_A_1005_99#_c_477_n 0.0236428f $X=7.5 $Y=1.3 $X2=0
+ $Y2=0
cc_277 N_A_263_409#_c_295_n N_A_1005_99#_c_477_n 0.0066343f $X=7.51 $Y=1.38
+ $X2=0 $Y2=0
cc_278 N_A_263_409#_c_284_n N_A_1005_99#_c_484_n 8.75045e-19 $X=7.55 $Y=1.785
+ $X2=0 $Y2=0
cc_279 N_A_263_409#_c_292_n N_A_1005_99#_c_484_n 0.00870019f $X=7.345 $Y=1.3
+ $X2=0 $Y2=0
cc_280 N_A_263_409#_c_341_p N_A_1005_99#_c_484_n 0.00970825f $X=6.68 $Y=1.3
+ $X2=0 $Y2=0
cc_281 N_A_263_409#_M1006_g N_A_1005_99#_c_478_n 0.00629944f $X=7.5 $Y=0.835
+ $X2=0 $Y2=0
cc_282 N_A_263_409#_c_343_p N_A_1005_99#_c_478_n 0.00634968f $X=6.51 $Y=0.95
+ $X2=0 $Y2=0
cc_283 N_A_263_409#_c_292_n N_A_1005_99#_c_478_n 0.015102f $X=7.345 $Y=1.3 $X2=0
+ $Y2=0
cc_284 N_A_263_409#_c_294_n N_A_1005_99#_c_478_n 0.00515087f $X=7.5 $Y=1.3 $X2=0
+ $Y2=0
cc_285 N_A_263_409#_c_295_n N_A_1005_99#_c_478_n 4.34354e-19 $X=7.51 $Y=1.38
+ $X2=0 $Y2=0
cc_286 N_A_263_409#_c_347_p N_A_747_79#_M1021_g 0.00449073f $X=6.055 $Y=0.865
+ $X2=0 $Y2=0
cc_287 N_A_263_409#_c_343_p N_A_747_79#_M1021_g 0.00766482f $X=6.51 $Y=0.95
+ $X2=0 $Y2=0
cc_288 N_A_263_409#_c_291_n N_A_747_79#_M1021_g 0.00625598f $X=6.595 $Y=1.215
+ $X2=0 $Y2=0
cc_289 N_A_263_409#_c_292_n N_A_747_79#_c_578_n 0.0246314f $X=7.345 $Y=1.3 $X2=0
+ $Y2=0
cc_290 N_A_263_409#_c_295_n N_A_747_79#_c_578_n 0.00978597f $X=7.51 $Y=1.38
+ $X2=0 $Y2=0
cc_291 N_A_263_409#_M1006_g N_A_747_79#_M1018_g 0.015494f $X=7.5 $Y=0.835 $X2=0
+ $Y2=0
cc_292 N_A_263_409#_c_343_p N_A_747_79#_M1018_g 4.84883e-19 $X=6.51 $Y=0.95
+ $X2=0 $Y2=0
cc_293 N_A_263_409#_c_291_n N_A_747_79#_M1018_g 9.62666e-19 $X=6.595 $Y=1.215
+ $X2=0 $Y2=0
cc_294 N_A_263_409#_c_280_n N_A_747_79#_c_580_n 0.00222855f $X=4.435 $Y=1.155
+ $X2=0 $Y2=0
cc_295 N_A_263_409#_c_282_n N_A_747_79#_c_580_n 6.80129e-19 $X=3.87 $Y=1.365
+ $X2=0 $Y2=0
cc_296 N_A_263_409#_c_283_n N_A_747_79#_c_580_n 0.00480855f $X=3.87 $Y=1.185
+ $X2=0 $Y2=0
cc_297 N_A_263_409#_c_290_n N_A_747_79#_c_580_n 0.0151147f $X=4.715 $Y=0.54
+ $X2=0 $Y2=0
cc_298 N_A_263_409#_c_280_n N_A_747_79#_c_581_n 0.0076778f $X=4.435 $Y=1.155
+ $X2=0 $Y2=0
cc_299 N_A_263_409#_c_283_n N_A_747_79#_c_581_n 0.00605665f $X=3.87 $Y=1.185
+ $X2=0 $Y2=0
cc_300 N_A_263_409#_c_287_n N_A_747_79#_c_581_n 0.0301712f $X=4.62 $Y=1.32 $X2=0
+ $Y2=0
cc_301 N_A_263_409#_c_288_n N_A_747_79#_c_581_n 0.00150778f $X=4.62 $Y=1.32
+ $X2=0 $Y2=0
cc_302 N_A_263_409#_c_296_n N_A_747_79#_c_581_n 0.0146442f $X=4.36 $Y=1.32 $X2=0
+ $Y2=0
cc_303 N_A_263_409#_c_297_n N_A_747_79#_c_589_n 0.00942938f $X=3.995 $Y=1.7
+ $X2=0 $Y2=0
cc_304 N_A_263_409#_c_287_n N_A_747_79#_c_590_n 0.0132822f $X=4.62 $Y=1.32 $X2=0
+ $Y2=0
cc_305 N_A_263_409#_c_288_n N_A_747_79#_c_590_n 0.00290452f $X=4.62 $Y=1.32
+ $X2=0 $Y2=0
cc_306 N_A_263_409#_c_287_n N_A_747_79#_c_582_n 0.0356951f $X=4.62 $Y=1.32 $X2=0
+ $Y2=0
cc_307 N_A_263_409#_c_288_n N_A_747_79#_c_582_n 0.00231241f $X=4.62 $Y=1.32
+ $X2=0 $Y2=0
cc_308 N_A_263_409#_c_289_n N_A_747_79#_c_618_n 0.0485251f $X=5.97 $Y=0.54 $X2=0
+ $Y2=0
cc_309 N_A_263_409#_c_347_p N_A_747_79#_c_618_n 0.00464226f $X=6.055 $Y=0.865
+ $X2=0 $Y2=0
cc_310 N_A_263_409#_c_371_p N_A_747_79#_c_618_n 0.00953072f $X=6.14 $Y=0.95
+ $X2=0 $Y2=0
cc_311 N_A_263_409#_c_287_n N_A_747_79#_c_621_n 0.0133519f $X=4.62 $Y=1.32 $X2=0
+ $Y2=0
cc_312 N_A_263_409#_c_289_n N_A_747_79#_c_621_n 0.0104568f $X=5.97 $Y=0.54 $X2=0
+ $Y2=0
cc_313 N_A_263_409#_c_371_p N_A_747_79#_c_583_n 0.00465883f $X=6.14 $Y=0.95
+ $X2=0 $Y2=0
cc_314 N_A_263_409#_c_289_n N_A_747_79#_c_585_n 0.00597822f $X=5.97 $Y=0.54
+ $X2=0 $Y2=0
cc_315 N_A_263_409#_c_343_p N_A_747_79#_c_585_n 0.0133878f $X=6.51 $Y=0.95 $X2=0
+ $Y2=0
cc_316 N_A_263_409#_c_371_p N_A_747_79#_c_585_n 0.0133845f $X=6.14 $Y=0.95 $X2=0
+ $Y2=0
cc_317 N_A_263_409#_c_341_p N_A_747_79#_c_585_n 0.0137025f $X=6.68 $Y=1.3 $X2=0
+ $Y2=0
cc_318 N_A_263_409#_c_283_n N_A_747_79#_c_594_n 0.00182271f $X=3.87 $Y=1.185
+ $X2=0 $Y2=0
cc_319 N_A_263_409#_c_288_n N_A_747_79#_c_594_n 0.00679264f $X=4.62 $Y=1.32
+ $X2=0 $Y2=0
cc_320 N_A_263_409#_c_296_n N_A_747_79#_c_594_n 4.95198e-19 $X=4.36 $Y=1.32
+ $X2=0 $Y2=0
cc_321 N_A_263_409#_c_343_p N_A_747_79#_c_586_n 0.0118769f $X=6.51 $Y=0.95 $X2=0
+ $Y2=0
cc_322 N_A_263_409#_c_371_p N_A_747_79#_c_586_n 0.00322409f $X=6.14 $Y=0.95
+ $X2=0 $Y2=0
cc_323 N_A_263_409#_c_292_n N_A_747_79#_c_586_n 0.00720465f $X=7.345 $Y=1.3
+ $X2=0 $Y2=0
cc_324 N_A_263_409#_c_341_p N_A_747_79#_c_586_n 0.00976376f $X=6.68 $Y=1.3 $X2=0
+ $Y2=0
cc_325 N_A_263_409#_c_294_n N_A_747_79#_c_586_n 0.0010437f $X=7.5 $Y=1.3 $X2=0
+ $Y2=0
cc_326 N_A_263_409#_c_295_n N_A_747_79#_c_586_n 0.00434048f $X=7.51 $Y=1.38
+ $X2=0 $Y2=0
cc_327 N_A_263_409#_c_302_n N_A_27_57#_M1019_g 0.013572f $X=1.455 $Y=2.9 $X2=0
+ $Y2=0
cc_328 N_A_263_409#_c_306_n N_A_27_57#_M1019_g 0.00575263f $X=1.455 $Y=2.19
+ $X2=0 $Y2=0
cc_329 N_A_263_409#_c_307_n N_A_27_57#_M1019_g 0.00343701f $X=1.567 $Y=2.025
+ $X2=0 $Y2=0
cc_330 N_A_263_409#_c_293_n N_A_27_57#_c_701_n 0.00173624f $X=1.85 $Y=0.495
+ $X2=0 $Y2=0
cc_331 N_A_263_409#_c_285_n N_A_27_57#_c_702_n 0.00135522f $X=1.76 $Y=1.68 $X2=0
+ $Y2=0
cc_332 N_A_263_409#_c_293_n N_A_27_57#_c_702_n 0.00880202f $X=1.85 $Y=0.495
+ $X2=0 $Y2=0
cc_333 N_A_263_409#_c_285_n N_A_27_57#_c_703_n 0.00905619f $X=1.76 $Y=1.68 $X2=0
+ $Y2=0
cc_334 N_A_263_409#_c_293_n N_A_27_57#_c_703_n 0.00602847f $X=1.85 $Y=0.495
+ $X2=0 $Y2=0
cc_335 N_A_263_409#_c_285_n N_A_27_57#_c_704_n 0.00469391f $X=1.76 $Y=1.68 $X2=0
+ $Y2=0
cc_336 N_A_263_409#_c_285_n N_A_27_57#_c_705_n 0.0121249f $X=1.76 $Y=1.68 $X2=0
+ $Y2=0
cc_337 N_A_263_409#_c_304_n N_A_27_57#_c_705_n 0.0195329f $X=2.935 $Y=1.765
+ $X2=0 $Y2=0
cc_338 N_A_263_409#_c_307_n N_A_27_57#_c_705_n 0.0360451f $X=1.567 $Y=2.025
+ $X2=0 $Y2=0
cc_339 N_A_263_409#_c_285_n N_A_27_57#_c_706_n 4.41971e-19 $X=1.76 $Y=1.68 $X2=0
+ $Y2=0
cc_340 N_A_263_409#_c_293_n N_A_27_57#_c_706_n 0.00452666f $X=1.85 $Y=0.495
+ $X2=0 $Y2=0
cc_341 N_A_263_409#_c_297_n N_A_27_57#_c_723_n 0.0151223f $X=3.995 $Y=1.7 $X2=0
+ $Y2=0
cc_342 N_A_263_409#_c_280_n N_A_27_57#_M1013_g 0.00333634f $X=4.435 $Y=1.155
+ $X2=0 $Y2=0
cc_343 N_A_263_409#_c_282_n N_A_27_57#_M1013_g 0.0079605f $X=3.87 $Y=1.365 $X2=0
+ $Y2=0
cc_344 N_A_263_409#_c_280_n N_A_27_57#_c_710_n 0.00907339f $X=4.435 $Y=1.155
+ $X2=0 $Y2=0
cc_345 N_A_263_409#_M1006_g N_A_27_57#_c_710_n 0.00861067f $X=7.5 $Y=0.835 $X2=0
+ $Y2=0
cc_346 N_A_263_409#_c_289_n N_A_27_57#_c_710_n 0.0274132f $X=5.97 $Y=0.54 $X2=0
+ $Y2=0
cc_347 N_A_263_409#_c_290_n N_A_27_57#_c_710_n 0.00421105f $X=4.715 $Y=0.54
+ $X2=0 $Y2=0
cc_348 N_A_263_409#_c_343_p N_A_27_57#_c_710_n 0.00484557f $X=6.51 $Y=0.95 $X2=0
+ $Y2=0
cc_349 N_A_263_409#_c_297_n N_A_27_57#_M1007_g 0.0214795f $X=3.995 $Y=1.7 $X2=0
+ $Y2=0
cc_350 N_A_263_409#_c_288_n N_A_27_57#_M1007_g 0.0122814f $X=4.62 $Y=1.32 $X2=0
+ $Y2=0
cc_351 N_A_263_409#_c_298_n N_A_27_57#_M1008_g 0.0258902f $X=7.55 $Y=1.91 $X2=0
+ $Y2=0
cc_352 N_A_263_409#_c_292_n N_A_27_57#_M1008_g 8.49446e-19 $X=7.345 $Y=1.3 $X2=0
+ $Y2=0
cc_353 N_A_263_409#_M1006_g N_A_27_57#_c_711_n 0.00799181f $X=7.5 $Y=0.835 $X2=0
+ $Y2=0
cc_354 N_A_263_409#_c_285_n N_A_27_57#_c_712_n 0.00360583f $X=1.76 $Y=1.68 $X2=0
+ $Y2=0
cc_355 N_A_263_409#_c_306_n N_A_27_57#_c_712_n 0.00116963f $X=1.455 $Y=2.19
+ $X2=0 $Y2=0
cc_356 N_A_263_409#_c_308_n N_A_27_57#_c_712_n 0.00431424f $X=1.76 $Y=1.765
+ $X2=0 $Y2=0
cc_357 N_A_263_409#_c_285_n N_A_27_57#_c_719_n 0.0484938f $X=1.76 $Y=1.68 $X2=0
+ $Y2=0
cc_358 N_A_263_409#_c_306_n N_A_27_57#_c_719_n 0.00754636f $X=1.455 $Y=2.19
+ $X2=0 $Y2=0
cc_359 N_A_263_409#_c_285_n N_A_27_57#_c_720_n 0.00459798f $X=1.76 $Y=1.68 $X2=0
+ $Y2=0
cc_360 N_A_263_409#_c_284_n N_A_1583_285#_M1005_g 0.046031f $X=7.55 $Y=1.785
+ $X2=0 $Y2=0
cc_361 N_A_263_409#_c_295_n N_A_1583_285#_M1002_g 0.00222721f $X=7.51 $Y=1.38
+ $X2=0 $Y2=0
cc_362 N_A_263_409#_c_295_n N_A_1583_285#_c_880_n 0.046031f $X=7.51 $Y=1.38
+ $X2=0 $Y2=0
cc_363 N_A_263_409#_c_298_n N_A_1429_383#_c_1002_n 0.0182875f $X=7.55 $Y=1.91
+ $X2=0 $Y2=0
cc_364 N_A_263_409#_M1006_g N_A_1429_383#_c_992_n 0.00419527f $X=7.5 $Y=0.835
+ $X2=0 $Y2=0
cc_365 N_A_263_409#_M1006_g N_A_1429_383#_c_993_n 2.30093e-19 $X=7.5 $Y=0.835
+ $X2=0 $Y2=0
cc_366 N_A_263_409#_c_298_n N_A_1429_383#_c_1001_n 0.0164162f $X=7.55 $Y=1.91
+ $X2=0 $Y2=0
cc_367 N_A_263_409#_M1006_g N_A_1429_383#_c_996_n 3.33074e-19 $X=7.5 $Y=0.835
+ $X2=0 $Y2=0
cc_368 N_A_263_409#_c_304_n N_VPWR_M1022_s 0.00482813f $X=2.935 $Y=1.765 $X2=0
+ $Y2=0
cc_369 N_A_263_409#_c_306_n N_VPWR_c_1082_n 0.0713253f $X=1.455 $Y=2.19 $X2=0
+ $Y2=0
cc_370 N_A_263_409#_c_304_n N_VPWR_c_1083_n 0.0255507f $X=2.935 $Y=1.765 $X2=0
+ $Y2=0
cc_371 N_A_263_409#_c_298_n N_VPWR_c_1089_n 0.00884004f $X=7.55 $Y=1.91 $X2=0
+ $Y2=0
cc_372 N_A_263_409#_c_302_n N_VPWR_c_1093_n 0.0372026f $X=1.455 $Y=2.9 $X2=0
+ $Y2=0
cc_373 N_A_263_409#_c_297_n N_VPWR_c_1081_n 0.00158331f $X=3.995 $Y=1.7 $X2=0
+ $Y2=0
cc_374 N_A_263_409#_c_298_n N_VPWR_c_1081_n 0.00885833f $X=7.55 $Y=1.91 $X2=0
+ $Y2=0
cc_375 N_A_263_409#_c_302_n N_VPWR_c_1081_n 0.0212868f $X=1.455 $Y=2.9 $X2=0
+ $Y2=0
cc_376 N_A_263_409#_c_282_n N_A_629_125#_c_1174_n 0.00705704f $X=3.87 $Y=1.365
+ $X2=0 $Y2=0
cc_377 N_A_263_409#_c_286_n N_A_629_125#_c_1174_n 0.00824215f $X=3.55 $Y=1.38
+ $X2=0 $Y2=0
cc_378 N_A_263_409#_c_282_n N_A_629_125#_c_1185_n 0.00353588f $X=3.87 $Y=1.365
+ $X2=0 $Y2=0
cc_379 N_A_263_409#_c_286_n N_A_629_125#_c_1185_n 0.0267255f $X=3.55 $Y=1.38
+ $X2=0 $Y2=0
cc_380 N_A_263_409#_c_297_n N_A_629_125#_c_1187_n 0.0132322f $X=3.995 $Y=1.7
+ $X2=0 $Y2=0
cc_381 N_A_263_409#_c_282_n N_A_629_125#_c_1187_n 0.00723375f $X=3.87 $Y=1.365
+ $X2=0 $Y2=0
cc_382 N_A_263_409#_c_286_n N_A_629_125#_c_1187_n 0.00208456f $X=3.55 $Y=1.38
+ $X2=0 $Y2=0
cc_383 N_A_263_409#_c_297_n N_A_629_125#_c_1175_n 6.89899e-19 $X=3.995 $Y=1.7
+ $X2=0 $Y2=0
cc_384 N_A_263_409#_c_282_n N_A_629_125#_c_1175_n 0.00834945f $X=3.87 $Y=1.365
+ $X2=0 $Y2=0
cc_385 N_A_263_409#_c_283_n N_A_629_125#_c_1175_n 0.0148058f $X=3.87 $Y=1.185
+ $X2=0 $Y2=0
cc_386 N_A_263_409#_c_286_n N_A_629_125#_c_1175_n 0.0234047f $X=3.55 $Y=1.38
+ $X2=0 $Y2=0
cc_387 N_A_263_409#_c_297_n N_A_629_125#_c_1177_n 0.0108879f $X=3.995 $Y=1.7
+ $X2=0 $Y2=0
cc_388 N_A_263_409#_c_282_n N_A_629_125#_c_1177_n 0.00542395f $X=3.87 $Y=1.365
+ $X2=0 $Y2=0
cc_389 N_A_263_409#_c_317_n N_A_629_125#_c_1177_n 0.00947413f $X=3.105 $Y=1.38
+ $X2=0 $Y2=0
cc_390 N_A_263_409#_c_286_n N_A_629_125#_c_1177_n 0.0264859f $X=3.55 $Y=1.38
+ $X2=0 $Y2=0
cc_391 N_A_263_409#_c_347_p N_VGND_M1029_d 0.0129752f $X=6.055 $Y=0.865 $X2=0
+ $Y2=0
cc_392 N_A_263_409#_c_343_p N_VGND_M1029_d 0.0120452f $X=6.51 $Y=0.95 $X2=0
+ $Y2=0
cc_393 N_A_263_409#_c_371_p N_VGND_M1029_d 0.00511516f $X=6.14 $Y=0.95 $X2=0
+ $Y2=0
cc_394 N_A_263_409#_c_291_n N_VGND_M1029_d 3.434e-19 $X=6.595 $Y=1.215 $X2=0
+ $Y2=0
cc_395 N_A_263_409#_c_293_n N_VGND_c_1235_n 0.0129849f $X=1.85 $Y=0.495 $X2=0
+ $Y2=0
cc_396 N_A_263_409#_c_285_n N_VGND_c_1236_n 0.0107001f $X=1.76 $Y=1.68 $X2=0
+ $Y2=0
cc_397 N_A_263_409#_c_293_n N_VGND_c_1236_n 0.0297074f $X=1.85 $Y=0.495 $X2=0
+ $Y2=0
cc_398 N_A_263_409#_c_289_n N_VGND_c_1237_n 0.0139106f $X=5.97 $Y=0.54 $X2=0
+ $Y2=0
cc_399 N_A_263_409#_c_347_p N_VGND_c_1237_n 0.00426607f $X=6.055 $Y=0.865 $X2=0
+ $Y2=0
cc_400 N_A_263_409#_c_343_p N_VGND_c_1237_n 0.0194844f $X=6.51 $Y=0.95 $X2=0
+ $Y2=0
cc_401 N_A_263_409#_c_293_n N_VGND_c_1240_n 0.0223445f $X=1.85 $Y=0.495 $X2=0
+ $Y2=0
cc_402 N_A_263_409#_c_289_n N_VGND_c_1247_n 0.0407503f $X=5.97 $Y=0.54 $X2=0
+ $Y2=0
cc_403 N_A_263_409#_c_290_n N_VGND_c_1247_n 0.00593614f $X=4.715 $Y=0.54 $X2=0
+ $Y2=0
cc_404 N_A_263_409#_c_280_n N_VGND_c_1249_n 9.49986e-19 $X=4.435 $Y=1.155 $X2=0
+ $Y2=0
cc_405 N_A_263_409#_M1006_g N_VGND_c_1249_n 9.49986e-19 $X=7.5 $Y=0.835 $X2=0
+ $Y2=0
cc_406 N_A_263_409#_c_289_n N_VGND_c_1249_n 0.0412635f $X=5.97 $Y=0.54 $X2=0
+ $Y2=0
cc_407 N_A_263_409#_c_290_n N_VGND_c_1249_n 0.00579697f $X=4.715 $Y=0.54 $X2=0
+ $Y2=0
cc_408 N_A_263_409#_c_343_p N_VGND_c_1249_n 0.00375058f $X=6.51 $Y=0.95 $X2=0
+ $Y2=0
cc_409 N_A_263_409#_c_293_n N_VGND_c_1249_n 0.0128543f $X=1.85 $Y=0.495 $X2=0
+ $Y2=0
cc_410 N_A_263_409#_c_287_n A_902_125# 0.00736423f $X=4.62 $Y=1.32 $X2=-0.19
+ $Y2=-0.245
cc_411 N_A_1005_99#_c_509_p N_A_747_79#_M1015_g 0.0293391f $X=6.51 $Y=1.81 $X2=0
+ $Y2=0
cc_412 N_A_1005_99#_c_481_n N_A_747_79#_M1015_g 0.00948544f $X=6.675 $Y=2.31
+ $X2=0 $Y2=0
cc_413 N_A_1005_99#_c_484_n N_A_747_79#_M1015_g 0.00129799f $X=6.675 $Y=1.85
+ $X2=0 $Y2=0
cc_414 N_A_1005_99#_c_478_n N_A_747_79#_M1021_g 0.0015701f $X=7.28 $Y=0.82 $X2=0
+ $Y2=0
cc_415 N_A_1005_99#_c_482_n N_A_747_79#_c_578_n 0.00117883f $X=7.835 $Y=1.81
+ $X2=0 $Y2=0
cc_416 N_A_1005_99#_c_484_n N_A_747_79#_c_578_n 4.5407e-19 $X=6.675 $Y=1.85
+ $X2=0 $Y2=0
cc_417 N_A_1005_99#_c_478_n N_A_747_79#_M1018_g 0.00797242f $X=7.28 $Y=0.82
+ $X2=0 $Y2=0
cc_418 N_A_1005_99#_M1016_g N_A_747_79#_c_590_n 0.00219551f $X=5.26 $Y=2.205
+ $X2=0 $Y2=0
cc_419 N_A_1005_99#_c_474_n N_A_747_79#_c_590_n 0.0030505f $X=5.34 $Y=1.32 $X2=0
+ $Y2=0
cc_420 N_A_1005_99#_c_518_p N_A_747_79#_c_590_n 0.0108661f $X=5.44 $Y=1.81 $X2=0
+ $Y2=0
cc_421 N_A_1005_99#_c_472_n N_A_747_79#_c_582_n 0.00576906f $X=5.1 $Y=1.155
+ $X2=0 $Y2=0
cc_422 N_A_1005_99#_M1016_g N_A_747_79#_c_582_n 0.00477737f $X=5.26 $Y=2.205
+ $X2=0 $Y2=0
cc_423 N_A_1005_99#_c_474_n N_A_747_79#_c_582_n 0.0353639f $X=5.34 $Y=1.32 $X2=0
+ $Y2=0
cc_424 N_A_1005_99#_c_475_n N_A_747_79#_c_582_n 0.00863992f $X=5.34 $Y=1.32
+ $X2=0 $Y2=0
cc_425 N_A_1005_99#_c_472_n N_A_747_79#_c_618_n 0.0117747f $X=5.1 $Y=1.155 $X2=0
+ $Y2=0
cc_426 N_A_1005_99#_c_474_n N_A_747_79#_c_618_n 0.0145086f $X=5.34 $Y=1.32 $X2=0
+ $Y2=0
cc_427 N_A_1005_99#_c_475_n N_A_747_79#_c_618_n 0.00572137f $X=5.34 $Y=1.32
+ $X2=0 $Y2=0
cc_428 N_A_1005_99#_c_472_n N_A_747_79#_c_621_n 0.00312875f $X=5.1 $Y=1.155
+ $X2=0 $Y2=0
cc_429 N_A_1005_99#_c_472_n N_A_747_79#_c_583_n 0.00294159f $X=5.1 $Y=1.155
+ $X2=0 $Y2=0
cc_430 N_A_1005_99#_c_474_n N_A_747_79#_c_583_n 0.00411602f $X=5.34 $Y=1.32
+ $X2=0 $Y2=0
cc_431 N_A_1005_99#_c_475_n N_A_747_79#_c_583_n 0.00155567f $X=5.34 $Y=1.32
+ $X2=0 $Y2=0
cc_432 N_A_1005_99#_M1016_g N_A_747_79#_c_584_n 2.56218e-19 $X=5.26 $Y=2.205
+ $X2=0 $Y2=0
cc_433 N_A_1005_99#_c_474_n N_A_747_79#_c_584_n 0.0260618f $X=5.34 $Y=1.32 $X2=0
+ $Y2=0
cc_434 N_A_1005_99#_c_475_n N_A_747_79#_c_584_n 0.00310022f $X=5.34 $Y=1.32
+ $X2=0 $Y2=0
cc_435 N_A_1005_99#_c_509_p N_A_747_79#_c_584_n 0.0135574f $X=6.51 $Y=1.81 $X2=0
+ $Y2=0
cc_436 N_A_1005_99#_c_509_p N_A_747_79#_c_585_n 0.0366925f $X=6.51 $Y=1.81 $X2=0
+ $Y2=0
cc_437 N_A_1005_99#_M1016_g N_A_747_79#_c_586_n 7.83211e-19 $X=5.26 $Y=2.205
+ $X2=0 $Y2=0
cc_438 N_A_1005_99#_c_474_n N_A_747_79#_c_586_n 2.92333e-19 $X=5.34 $Y=1.32
+ $X2=0 $Y2=0
cc_439 N_A_1005_99#_c_475_n N_A_747_79#_c_586_n 0.00508482f $X=5.34 $Y=1.32
+ $X2=0 $Y2=0
cc_440 N_A_1005_99#_c_509_p N_A_747_79#_c_586_n 0.00443747f $X=6.51 $Y=1.81
+ $X2=0 $Y2=0
cc_441 N_A_1005_99#_c_484_n N_A_747_79#_c_586_n 0.00758618f $X=6.675 $Y=1.85
+ $X2=0 $Y2=0
cc_442 N_A_1005_99#_c_472_n N_A_27_57#_c_710_n 0.00754956f $X=5.1 $Y=1.155 $X2=0
+ $Y2=0
cc_443 N_A_1005_99#_c_476_n N_A_27_57#_c_710_n 0.0021325f $X=7.835 $Y=0.95 $X2=0
+ $Y2=0
cc_444 N_A_1005_99#_c_478_n N_A_27_57#_c_710_n 0.00567968f $X=7.28 $Y=0.82 $X2=0
+ $Y2=0
cc_445 N_A_1005_99#_M1016_g N_A_27_57#_M1007_g 0.0435492f $X=5.26 $Y=2.205 $X2=0
+ $Y2=0
cc_446 N_A_1005_99#_c_518_p N_A_27_57#_M1007_g 3.05276e-19 $X=5.44 $Y=1.81 $X2=0
+ $Y2=0
cc_447 N_A_1005_99#_M1016_g N_A_27_57#_c_726_n 0.0149942f $X=5.26 $Y=2.205 $X2=0
+ $Y2=0
cc_448 N_A_1005_99#_c_481_n N_A_27_57#_c_726_n 0.00677547f $X=6.675 $Y=2.31
+ $X2=0 $Y2=0
cc_449 N_A_1005_99#_c_481_n N_A_27_57#_M1008_g 0.00919221f $X=6.675 $Y=2.31
+ $X2=0 $Y2=0
cc_450 N_A_1005_99#_c_482_n N_A_27_57#_M1008_g 0.0179442f $X=7.835 $Y=1.81 $X2=0
+ $Y2=0
cc_451 N_A_1005_99#_c_476_n N_A_27_57#_c_711_n 0.00236111f $X=7.835 $Y=0.95
+ $X2=0 $Y2=0
cc_452 N_A_1005_99#_c_478_n N_A_27_57#_c_711_n 7.80328e-19 $X=7.28 $Y=0.82 $X2=0
+ $Y2=0
cc_453 N_A_1005_99#_c_482_n N_A_1583_285#_M1005_g 0.00527609f $X=7.835 $Y=1.81
+ $X2=0 $Y2=0
cc_454 N_A_1005_99#_c_476_n N_A_1583_285#_M1002_g 6.53643e-19 $X=7.835 $Y=0.95
+ $X2=0 $Y2=0
cc_455 N_A_1005_99#_c_477_n N_A_1583_285#_M1002_g 0.00148416f $X=7.92 $Y=1.725
+ $X2=0 $Y2=0
cc_456 N_A_1005_99#_c_482_n N_A_1583_285#_c_880_n 0.00101517f $X=7.835 $Y=1.81
+ $X2=0 $Y2=0
cc_457 N_A_1005_99#_c_477_n N_A_1583_285#_c_880_n 0.00999844f $X=7.92 $Y=1.725
+ $X2=0 $Y2=0
cc_458 N_A_1005_99#_c_476_n N_A_1429_383#_M1006_d 0.00880095f $X=7.835 $Y=0.95
+ $X2=-0.19 $Y2=-0.245
cc_459 N_A_1005_99#_c_482_n N_A_1429_383#_c_1002_n 0.0347598f $X=7.835 $Y=1.81
+ $X2=0 $Y2=0
cc_460 N_A_1005_99#_c_476_n N_A_1429_383#_c_992_n 0.0230612f $X=7.835 $Y=0.95
+ $X2=0 $Y2=0
cc_461 N_A_1005_99#_c_478_n N_A_1429_383#_c_992_n 0.00520519f $X=7.28 $Y=0.82
+ $X2=0 $Y2=0
cc_462 N_A_1005_99#_c_476_n N_A_1429_383#_c_993_n 0.0100715f $X=7.835 $Y=0.95
+ $X2=0 $Y2=0
cc_463 N_A_1005_99#_c_482_n N_A_1429_383#_c_994_n 0.0128523f $X=7.835 $Y=1.81
+ $X2=0 $Y2=0
cc_464 N_A_1005_99#_c_477_n N_A_1429_383#_c_994_n 0.0381585f $X=7.92 $Y=1.725
+ $X2=0 $Y2=0
cc_465 N_A_1005_99#_c_481_n N_A_1429_383#_c_1001_n 0.0179092f $X=6.675 $Y=2.31
+ $X2=0 $Y2=0
cc_466 N_A_1005_99#_c_482_n N_A_1429_383#_c_1001_n 0.0208609f $X=7.835 $Y=1.81
+ $X2=0 $Y2=0
cc_467 N_A_1005_99#_c_476_n N_A_1429_383#_c_996_n 0.00354742f $X=7.835 $Y=0.95
+ $X2=0 $Y2=0
cc_468 N_A_1005_99#_c_477_n N_A_1429_383#_c_996_n 0.0105068f $X=7.92 $Y=1.725
+ $X2=0 $Y2=0
cc_469 N_A_1005_99#_c_509_p N_VPWR_M1016_d 0.0350509f $X=6.51 $Y=1.81 $X2=0
+ $Y2=0
cc_470 N_A_1005_99#_M1016_g N_VPWR_c_1084_n 0.0240515f $X=5.26 $Y=2.205 $X2=0
+ $Y2=0
cc_471 N_A_1005_99#_c_509_p N_VPWR_c_1084_n 0.0192545f $X=6.51 $Y=1.81 $X2=0
+ $Y2=0
cc_472 N_A_1005_99#_c_518_p N_VPWR_c_1084_n 0.00193953f $X=5.44 $Y=1.81 $X2=0
+ $Y2=0
cc_473 N_A_1005_99#_c_481_n N_VPWR_c_1089_n 0.012377f $X=6.675 $Y=2.31 $X2=0
+ $Y2=0
cc_474 N_A_1005_99#_M1016_g N_VPWR_c_1081_n 0.00143131f $X=5.26 $Y=2.205 $X2=0
+ $Y2=0
cc_475 N_A_1005_99#_c_481_n N_VPWR_c_1081_n 0.0104642f $X=6.675 $Y=2.31 $X2=0
+ $Y2=0
cc_476 N_A_1005_99#_c_478_n N_VGND_c_1237_n 0.00148716f $X=7.28 $Y=0.82 $X2=0
+ $Y2=0
cc_477 N_A_1005_99#_c_478_n N_VGND_c_1242_n 0.00674486f $X=7.28 $Y=0.82 $X2=0
+ $Y2=0
cc_478 N_A_1005_99#_c_478_n N_VGND_c_1249_n 0.00863043f $X=7.28 $Y=0.82 $X2=0
+ $Y2=0
cc_479 N_A_747_79#_c_589_n N_A_27_57#_c_723_n 0.00651605f $X=4.34 $Y=2.28 $X2=0
+ $Y2=0
cc_480 N_A_747_79#_c_580_n N_A_27_57#_M1013_g 0.00440785f $X=4.175 $Y=0.53 $X2=0
+ $Y2=0
cc_481 N_A_747_79#_c_581_n N_A_27_57#_M1013_g 0.0013645f $X=4.26 $Y=1.685 $X2=0
+ $Y2=0
cc_482 N_A_747_79#_M1021_g N_A_27_57#_c_710_n 0.00891853f $X=6.7 $Y=0.835 $X2=0
+ $Y2=0
cc_483 N_A_747_79#_M1018_g N_A_27_57#_c_710_n 0.00897576f $X=7.06 $Y=0.835 $X2=0
+ $Y2=0
cc_484 N_A_747_79#_c_580_n N_A_27_57#_c_710_n 0.0117828f $X=4.175 $Y=0.53 $X2=0
+ $Y2=0
cc_485 N_A_747_79#_c_589_n N_A_27_57#_M1007_g 0.00810551f $X=4.34 $Y=2.28 $X2=0
+ $Y2=0
cc_486 N_A_747_79#_c_590_n N_A_27_57#_M1007_g 0.0184753f $X=4.895 $Y=1.77 $X2=0
+ $Y2=0
cc_487 N_A_747_79#_M1015_g N_A_27_57#_c_726_n 0.0151223f $X=6.33 $Y=2.205 $X2=0
+ $Y2=0
cc_488 N_A_747_79#_M1015_g N_A_27_57#_M1008_g 0.0205686f $X=6.33 $Y=2.205 $X2=0
+ $Y2=0
cc_489 N_A_747_79#_c_578_n N_A_27_57#_M1008_g 0.00624767f $X=6.985 $Y=1.29 $X2=0
+ $Y2=0
cc_490 N_A_747_79#_M1015_g N_VPWR_c_1084_n 0.0207515f $X=6.33 $Y=2.205 $X2=0
+ $Y2=0
cc_491 N_A_747_79#_c_589_n N_VPWR_c_1094_n 0.0102491f $X=4.34 $Y=2.28 $X2=0
+ $Y2=0
cc_492 N_A_747_79#_M1015_g N_VPWR_c_1081_n 0.00158331f $X=6.33 $Y=2.205 $X2=0
+ $Y2=0
cc_493 N_A_747_79#_c_589_n N_VPWR_c_1081_n 0.0100074f $X=4.34 $Y=2.28 $X2=0
+ $Y2=0
cc_494 N_A_747_79#_c_580_n N_A_629_125#_c_1173_n 0.0129833f $X=4.175 $Y=0.53
+ $X2=0 $Y2=0
cc_495 N_A_747_79#_c_581_n N_A_629_125#_c_1173_n 0.00315686f $X=4.26 $Y=1.685
+ $X2=0 $Y2=0
cc_496 N_A_747_79#_c_580_n N_A_629_125#_c_1174_n 0.0198497f $X=4.175 $Y=0.53
+ $X2=0 $Y2=0
cc_497 N_A_747_79#_c_581_n N_A_629_125#_c_1174_n 0.0135567f $X=4.26 $Y=1.685
+ $X2=0 $Y2=0
cc_498 N_A_747_79#_c_581_n N_A_629_125#_c_1175_n 0.044454f $X=4.26 $Y=1.685
+ $X2=0 $Y2=0
cc_499 N_A_747_79#_c_594_n N_A_629_125#_c_1175_n 0.00208615f $X=4.34 $Y=1.85
+ $X2=0 $Y2=0
cc_500 N_A_747_79#_c_589_n N_A_629_125#_c_1177_n 0.0141953f $X=4.34 $Y=2.28
+ $X2=0 $Y2=0
cc_501 N_A_747_79#_c_590_n A_962_371# 0.00993389f $X=4.895 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_502 N_A_747_79#_c_618_n N_VGND_M1029_d 0.0183712f $X=5.62 $Y=0.89 $X2=0 $Y2=0
cc_503 N_A_747_79#_c_583_n N_VGND_M1029_d 0.00266904f $X=5.705 $Y=1.215 $X2=0
+ $Y2=0
cc_504 N_A_747_79#_M1021_g N_VGND_c_1237_n 0.00615937f $X=6.7 $Y=0.835 $X2=0
+ $Y2=0
cc_505 N_A_747_79#_c_586_n N_VGND_c_1237_n 2.19889e-19 $X=6.775 $Y=1.38 $X2=0
+ $Y2=0
cc_506 N_A_747_79#_c_580_n N_VGND_c_1247_n 0.0245567f $X=4.175 $Y=0.53 $X2=0
+ $Y2=0
cc_507 N_A_747_79#_M1021_g N_VGND_c_1249_n 9.49986e-19 $X=6.7 $Y=0.835 $X2=0
+ $Y2=0
cc_508 N_A_747_79#_M1018_g N_VGND_c_1249_n 9.49986e-19 $X=7.06 $Y=0.835 $X2=0
+ $Y2=0
cc_509 N_A_747_79#_c_580_n N_VGND_c_1249_n 0.0200405f $X=4.175 $Y=0.53 $X2=0
+ $Y2=0
cc_510 N_A_747_79#_c_582_n A_902_125# 6.41675e-19 $X=4.98 $Y=1.685 $X2=-0.19
+ $Y2=-0.245
cc_511 N_A_747_79#_c_621_n A_902_125# 0.00238044f $X=5.065 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_512 N_A_27_57#_c_710_n N_A_1583_285#_M1002_g 0.0420758f $X=7.98 $Y=0.18 $X2=0
+ $Y2=0
cc_513 N_A_27_57#_c_711_n N_A_1583_285#_c_880_n 0.00524353f $X=8.055 $Y=0.255
+ $X2=0 $Y2=0
cc_514 N_A_27_57#_c_710_n N_A_1429_383#_c_992_n 0.00488144f $X=7.98 $Y=0.18
+ $X2=0 $Y2=0
cc_515 N_A_27_57#_c_711_n N_A_1429_383#_c_992_n 0.0155163f $X=8.055 $Y=0.255
+ $X2=0 $Y2=0
cc_516 N_A_27_57#_c_711_n N_A_1429_383#_c_993_n 0.00231161f $X=8.055 $Y=0.255
+ $X2=0 $Y2=0
cc_517 N_A_27_57#_M1008_g N_A_1429_383#_c_1001_n 0.0158007f $X=7.02 $Y=2.415
+ $X2=0 $Y2=0
cc_518 N_A_27_57#_M1019_g N_VPWR_c_1082_n 0.0245357f $X=1.19 $Y=2.545 $X2=0
+ $Y2=0
cc_519 N_A_27_57#_c_731_n N_VPWR_c_1082_n 0.0702172f $X=0.395 $Y=2.19 $X2=0
+ $Y2=0
cc_520 N_A_27_57#_c_705_n N_VPWR_c_1083_n 0.0305318f $X=2.07 $Y=3.075 $X2=0
+ $Y2=0
cc_521 N_A_27_57#_c_723_n N_VPWR_c_1083_n 0.0260211f $X=4.56 $Y=3.15 $X2=0 $Y2=0
cc_522 N_A_27_57#_M1007_g N_VPWR_c_1084_n 0.00955426f $X=4.685 $Y=2.355 $X2=0
+ $Y2=0
cc_523 N_A_27_57#_c_726_n N_VPWR_c_1084_n 0.0258253f $X=6.895 $Y=3.15 $X2=0
+ $Y2=0
cc_524 N_A_27_57#_c_730_n N_VPWR_c_1087_n 0.0304602f $X=0.395 $Y=2.9 $X2=0 $Y2=0
cc_525 N_A_27_57#_c_726_n N_VPWR_c_1089_n 0.0478909f $X=6.895 $Y=3.15 $X2=0
+ $Y2=0
cc_526 N_A_27_57#_M1019_g N_VPWR_c_1093_n 0.00769046f $X=1.19 $Y=2.545 $X2=0
+ $Y2=0
cc_527 N_A_27_57#_c_724_n N_VPWR_c_1093_n 0.0200932f $X=2.145 $Y=3.15 $X2=0
+ $Y2=0
cc_528 N_A_27_57#_c_723_n N_VPWR_c_1094_n 0.0816539f $X=4.56 $Y=3.15 $X2=0 $Y2=0
cc_529 N_A_27_57#_M1019_g N_VPWR_c_1081_n 0.0139316f $X=1.19 $Y=2.545 $X2=0
+ $Y2=0
cc_530 N_A_27_57#_c_723_n N_VPWR_c_1081_n 0.0842662f $X=4.56 $Y=3.15 $X2=0 $Y2=0
cc_531 N_A_27_57#_c_724_n N_VPWR_c_1081_n 0.0111576f $X=2.145 $Y=3.15 $X2=0
+ $Y2=0
cc_532 N_A_27_57#_c_726_n N_VPWR_c_1081_n 0.0928089f $X=6.895 $Y=3.15 $X2=0
+ $Y2=0
cc_533 N_A_27_57#_c_729_n N_VPWR_c_1081_n 0.0154456f $X=4.685 $Y=3.15 $X2=0
+ $Y2=0
cc_534 N_A_27_57#_c_730_n N_VPWR_c_1081_n 0.0174175f $X=0.395 $Y=2.9 $X2=0 $Y2=0
cc_535 N_A_27_57#_c_707_n N_A_629_125#_c_1173_n 0.0068262f $X=3.585 $Y=0.18
+ $X2=0 $Y2=0
cc_536 N_A_27_57#_M1013_g N_A_629_125#_c_1173_n 0.0051503f $X=3.66 $Y=0.605
+ $X2=0 $Y2=0
cc_537 N_A_27_57#_M1013_g N_A_629_125#_c_1174_n 0.0101104f $X=3.66 $Y=0.605
+ $X2=0 $Y2=0
cc_538 N_A_27_57#_c_723_n N_A_629_125#_c_1177_n 0.00653589f $X=4.56 $Y=3.15
+ $X2=0 $Y2=0
cc_539 N_A_27_57#_c_701_n N_VGND_c_1235_n 0.0105779f $X=1.275 $Y=0.78 $X2=0
+ $Y2=0
cc_540 N_A_27_57#_c_702_n N_VGND_c_1235_n 0.00188833f $X=1.635 $Y=0.78 $X2=0
+ $Y2=0
cc_541 N_A_27_57#_c_715_n N_VGND_c_1235_n 0.0127138f $X=0.27 $Y=0.495 $X2=0
+ $Y2=0
cc_542 N_A_27_57#_c_716_n N_VGND_c_1235_n 0.0171154f $X=1.165 $Y=0.91 $X2=0
+ $Y2=0
cc_543 N_A_27_57#_c_719_n N_VGND_c_1235_n 0.00316485f $X=1.33 $Y=0.99 $X2=0
+ $Y2=0
cc_544 N_A_27_57#_c_702_n N_VGND_c_1236_n 5.89795e-19 $X=1.635 $Y=0.78 $X2=0
+ $Y2=0
cc_545 N_A_27_57#_c_705_n N_VGND_c_1236_n 6.88645e-19 $X=2.07 $Y=3.075 $X2=0
+ $Y2=0
cc_546 N_A_27_57#_c_706_n N_VGND_c_1236_n 0.010994f $X=2.135 $Y=0.78 $X2=0 $Y2=0
cc_547 N_A_27_57#_c_707_n N_VGND_c_1236_n 0.024104f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_548 N_A_27_57#_c_710_n N_VGND_c_1237_n 0.0210695f $X=7.98 $Y=0.18 $X2=0 $Y2=0
cc_549 N_A_27_57#_c_710_n N_VGND_c_1238_n 0.00297089f $X=7.98 $Y=0.18 $X2=0
+ $Y2=0
cc_550 N_A_27_57#_c_701_n N_VGND_c_1240_n 0.00445056f $X=1.275 $Y=0.78 $X2=0
+ $Y2=0
cc_551 N_A_27_57#_c_702_n N_VGND_c_1240_n 0.00488765f $X=1.635 $Y=0.78 $X2=0
+ $Y2=0
cc_552 N_A_27_57#_c_704_n N_VGND_c_1240_n 5.84324e-19 $X=1.71 $Y=0.855 $X2=0
+ $Y2=0
cc_553 N_A_27_57#_c_708_n N_VGND_c_1240_n 0.0077661f $X=2.21 $Y=0.18 $X2=0 $Y2=0
cc_554 N_A_27_57#_c_710_n N_VGND_c_1242_n 0.0460214f $X=7.98 $Y=0.18 $X2=0 $Y2=0
cc_555 N_A_27_57#_c_715_n N_VGND_c_1246_n 0.0220321f $X=0.27 $Y=0.495 $X2=0
+ $Y2=0
cc_556 N_A_27_57#_c_707_n N_VGND_c_1247_n 0.099357f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_557 N_A_27_57#_c_701_n N_VGND_c_1249_n 0.0041935f $X=1.275 $Y=0.78 $X2=0
+ $Y2=0
cc_558 N_A_27_57#_c_702_n N_VGND_c_1249_n 0.00915117f $X=1.635 $Y=0.78 $X2=0
+ $Y2=0
cc_559 N_A_27_57#_c_704_n N_VGND_c_1249_n 7.93839e-19 $X=1.71 $Y=0.855 $X2=0
+ $Y2=0
cc_560 N_A_27_57#_c_707_n N_VGND_c_1249_n 0.0413034f $X=3.585 $Y=0.18 $X2=0
+ $Y2=0
cc_561 N_A_27_57#_c_708_n N_VGND_c_1249_n 0.0106372f $X=2.21 $Y=0.18 $X2=0 $Y2=0
cc_562 N_A_27_57#_c_710_n N_VGND_c_1249_n 0.124042f $X=7.98 $Y=0.18 $X2=0 $Y2=0
cc_563 N_A_27_57#_c_714_n N_VGND_c_1249_n 0.00835521f $X=3.66 $Y=0.18 $X2=0
+ $Y2=0
cc_564 N_A_27_57#_c_715_n N_VGND_c_1249_n 0.0125808f $X=0.27 $Y=0.495 $X2=0
+ $Y2=0
cc_565 N_A_27_57#_c_716_n N_VGND_c_1249_n 0.0152176f $X=1.165 $Y=0.91 $X2=0
+ $Y2=0
cc_566 N_A_27_57#_c_719_n N_VGND_c_1249_n 0.00947285f $X=1.33 $Y=0.99 $X2=0
+ $Y2=0
cc_567 N_A_1583_285#_M1002_g N_A_1429_383#_c_987_n 0.0182326f $X=8.415 $Y=0.585
+ $X2=0 $Y2=0
cc_568 N_A_1583_285#_c_887_n N_A_1429_383#_c_987_n 0.00100061f $X=9.63 $Y=0.54
+ $X2=0 $Y2=0
cc_569 N_A_1583_285#_c_881_n N_A_1429_383#_M1017_g 0.00121712f $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_570 N_A_1583_285#_c_882_n N_A_1429_383#_M1017_g 0.0106274f $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_571 N_A_1583_285#_c_893_n N_A_1429_383#_M1017_g 0.0259581f $X=9.39 $Y=1.84
+ $X2=0 $Y2=0
cc_572 N_A_1583_285#_c_883_n N_A_1429_383#_M1017_g 0.0070341f $X=9.555 $Y=1.925
+ $X2=0 $Y2=0
cc_573 N_A_1583_285#_c_896_n N_A_1429_383#_M1017_g 0.0219f $X=9.555 $Y=2.06
+ $X2=0 $Y2=0
cc_574 N_A_1583_285#_c_884_n N_A_1429_383#_M1017_g 3.13142e-19 $X=9.63 $Y=1.585
+ $X2=0 $Y2=0
cc_575 N_A_1583_285#_c_884_n N_A_1429_383#_c_989_n 0.00539816f $X=9.63 $Y=1.585
+ $X2=0 $Y2=0
cc_576 N_A_1583_285#_c_887_n N_A_1429_383#_c_989_n 0.00687218f $X=9.63 $Y=0.54
+ $X2=0 $Y2=0
cc_577 N_A_1583_285#_c_882_n N_A_1429_383#_c_990_n 0.00236081f $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_578 N_A_1583_285#_c_884_n N_A_1429_383#_c_990_n 0.00996954f $X=9.63 $Y=1.585
+ $X2=0 $Y2=0
cc_579 N_A_1583_285#_c_887_n N_A_1429_383#_c_990_n 0.00134873f $X=9.63 $Y=0.54
+ $X2=0 $Y2=0
cc_580 N_A_1583_285#_c_881_n N_A_1429_383#_c_991_n 5.22586e-19 $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_581 N_A_1583_285#_c_882_n N_A_1429_383#_c_991_n 0.00971337f $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_582 N_A_1583_285#_c_893_n N_A_1429_383#_c_991_n 0.00125287f $X=9.39 $Y=1.84
+ $X2=0 $Y2=0
cc_583 N_A_1583_285#_M1005_g N_A_1429_383#_c_1002_n 0.0278862f $X=8.04 $Y=2.415
+ $X2=0 $Y2=0
cc_584 N_A_1583_285#_M1002_g N_A_1429_383#_c_992_n 0.00637637f $X=8.415 $Y=0.585
+ $X2=0 $Y2=0
cc_585 N_A_1583_285#_M1002_g N_A_1429_383#_c_993_n 0.00680161f $X=8.415 $Y=0.585
+ $X2=0 $Y2=0
cc_586 N_A_1583_285#_M1005_g N_A_1429_383#_c_994_n 0.00796362f $X=8.04 $Y=2.415
+ $X2=0 $Y2=0
cc_587 N_A_1583_285#_M1002_g N_A_1429_383#_c_994_n 0.0139331f $X=8.415 $Y=0.585
+ $X2=0 $Y2=0
cc_588 N_A_1583_285#_c_880_n N_A_1429_383#_c_994_n 0.0218529f $X=8.49 $Y=1.59
+ $X2=0 $Y2=0
cc_589 N_A_1583_285#_c_881_n N_A_1429_383#_c_994_n 0.0223622f $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_590 N_A_1583_285#_c_894_n N_A_1429_383#_c_994_n 0.0137557f $X=8.845 $Y=1.84
+ $X2=0 $Y2=0
cc_591 N_A_1583_285#_M1002_g N_A_1429_383#_c_995_n 0.0164609f $X=8.415 $Y=0.585
+ $X2=0 $Y2=0
cc_592 N_A_1583_285#_c_881_n N_A_1429_383#_c_995_n 0.017448f $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_593 N_A_1583_285#_c_882_n N_A_1429_383#_c_995_n 0.00332462f $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_594 N_A_1583_285#_c_893_n N_A_1429_383#_c_995_n 0.00662936f $X=9.39 $Y=1.84
+ $X2=0 $Y2=0
cc_595 N_A_1583_285#_M1005_g N_A_1429_383#_c_1001_n 0.00298041f $X=8.04 $Y=2.415
+ $X2=0 $Y2=0
cc_596 N_A_1583_285#_M1002_g N_A_1429_383#_c_996_n 0.00320991f $X=8.415 $Y=0.585
+ $X2=0 $Y2=0
cc_597 N_A_1583_285#_M1002_g N_A_1429_383#_c_997_n 0.00165544f $X=8.415 $Y=0.585
+ $X2=0 $Y2=0
cc_598 N_A_1583_285#_c_881_n N_A_1429_383#_c_997_n 0.00941545f $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_599 N_A_1583_285#_c_882_n N_A_1429_383#_c_997_n 6.05775e-19 $X=8.68 $Y=1.59
+ $X2=0 $Y2=0
cc_600 N_A_1583_285#_c_893_n N_A_1429_383#_c_997_n 0.0225956f $X=9.39 $Y=1.84
+ $X2=0 $Y2=0
cc_601 N_A_1583_285#_c_884_n N_A_1429_383#_c_997_n 0.0487486f $X=9.63 $Y=1.585
+ $X2=0 $Y2=0
cc_602 N_A_1583_285#_c_887_n N_A_1429_383#_c_997_n 0.00639351f $X=9.63 $Y=0.54
+ $X2=0 $Y2=0
cc_603 N_A_1583_285#_M1002_g N_A_1429_383#_c_998_n 0.00769862f $X=8.415 $Y=0.585
+ $X2=0 $Y2=0
cc_604 N_A_1583_285#_c_878_n N_A_1429_383#_c_998_n 0.00527205f $X=10.495
+ $Y=1.755 $X2=0 $Y2=0
cc_605 N_A_1583_285#_c_893_n N_VPWR_M1005_d 0.0064535f $X=9.39 $Y=1.84 $X2=0
+ $Y2=0
cc_606 N_A_1583_285#_c_894_n N_VPWR_M1005_d 0.0035555f $X=8.845 $Y=1.84 $X2=0
+ $Y2=0
cc_607 N_A_1583_285#_M1005_g N_VPWR_c_1085_n 0.0260302f $X=8.04 $Y=2.415 $X2=0
+ $Y2=0
cc_608 N_A_1583_285#_c_882_n N_VPWR_c_1085_n 0.00163568f $X=8.68 $Y=1.59 $X2=0
+ $Y2=0
cc_609 N_A_1583_285#_c_893_n N_VPWR_c_1085_n 0.00144617f $X=9.39 $Y=1.84 $X2=0
+ $Y2=0
cc_610 N_A_1583_285#_c_894_n N_VPWR_c_1085_n 0.0260939f $X=8.845 $Y=1.84 $X2=0
+ $Y2=0
cc_611 N_A_1583_285#_c_896_n N_VPWR_c_1085_n 0.0147614f $X=9.555 $Y=2.06 $X2=0
+ $Y2=0
cc_612 N_A_1583_285#_c_878_n N_VPWR_c_1086_n 0.00217959f $X=10.495 $Y=1.755
+ $X2=0 $Y2=0
cc_613 N_A_1583_285#_M1027_g N_VPWR_c_1086_n 0.0264343f $X=10.495 $Y=2.48 $X2=0
+ $Y2=0
cc_614 N_A_1583_285#_c_896_n N_VPWR_c_1086_n 0.0497626f $X=9.555 $Y=2.06 $X2=0
+ $Y2=0
cc_615 N_A_1583_285#_c_885_n N_VPWR_c_1086_n 0.025146f $X=10.085 $Y=1.67 $X2=0
+ $Y2=0
cc_616 N_A_1583_285#_M1005_g N_VPWR_c_1089_n 0.00908496f $X=8.04 $Y=2.415 $X2=0
+ $Y2=0
cc_617 N_A_1583_285#_c_896_n N_VPWR_c_1091_n 0.0123893f $X=9.555 $Y=2.06 $X2=0
+ $Y2=0
cc_618 N_A_1583_285#_M1027_g N_VPWR_c_1095_n 0.00687065f $X=10.495 $Y=2.48 $X2=0
+ $Y2=0
cc_619 N_A_1583_285#_M1005_g N_VPWR_c_1081_n 0.00885833f $X=8.04 $Y=2.415 $X2=0
+ $Y2=0
cc_620 N_A_1583_285#_M1027_g N_VPWR_c_1081_n 0.013111f $X=10.495 $Y=2.48 $X2=0
+ $Y2=0
cc_621 N_A_1583_285#_c_896_n N_VPWR_c_1081_n 0.0117798f $X=9.555 $Y=2.06 $X2=0
+ $Y2=0
cc_622 N_A_1583_285#_M1027_g N_Q_c_1219_n 0.0308063f $X=10.495 $Y=2.48 $X2=0
+ $Y2=0
cc_623 N_A_1583_285#_M1009_g Q 0.00221352f $X=10.195 $Y=0.67 $X2=0 $Y2=0
cc_624 N_A_1583_285#_c_878_n Q 0.0198246f $X=10.495 $Y=1.755 $X2=0 $Y2=0
cc_625 N_A_1583_285#_M1025_g Q 0.0164455f $X=10.555 $Y=0.67 $X2=0 $Y2=0
cc_626 N_A_1583_285#_c_885_n Q 0.0129505f $X=10.085 $Y=1.67 $X2=0 $Y2=0
cc_627 N_A_1583_285#_c_886_n Q 0.0358876f $X=10.25 $Y=1.25 $X2=0 $Y2=0
cc_628 N_A_1583_285#_c_878_n Q 0.00537765f $X=10.495 $Y=1.755 $X2=0 $Y2=0
cc_629 N_A_1583_285#_M1027_g Q 0.00156333f $X=10.495 $Y=2.48 $X2=0 $Y2=0
cc_630 N_A_1583_285#_M1002_g N_VGND_c_1238_n 0.00324809f $X=8.415 $Y=0.585 $X2=0
+ $Y2=0
cc_631 N_A_1583_285#_c_887_n N_VGND_c_1238_n 0.0124042f $X=9.63 $Y=0.54 $X2=0
+ $Y2=0
cc_632 N_A_1583_285#_M1009_g N_VGND_c_1239_n 0.0133811f $X=10.195 $Y=0.67 $X2=0
+ $Y2=0
cc_633 N_A_1583_285#_c_878_n N_VGND_c_1239_n 2.63397e-19 $X=10.495 $Y=1.755
+ $X2=0 $Y2=0
cc_634 N_A_1583_285#_M1025_g N_VGND_c_1239_n 0.00180169f $X=10.555 $Y=0.67 $X2=0
+ $Y2=0
cc_635 N_A_1583_285#_c_884_n N_VGND_c_1239_n 0.0128109f $X=9.63 $Y=1.585 $X2=0
+ $Y2=0
cc_636 N_A_1583_285#_c_886_n N_VGND_c_1239_n 0.00473449f $X=10.25 $Y=1.25 $X2=0
+ $Y2=0
cc_637 N_A_1583_285#_c_887_n N_VGND_c_1239_n 0.0293233f $X=9.63 $Y=0.54 $X2=0
+ $Y2=0
cc_638 N_A_1583_285#_M1002_g N_VGND_c_1242_n 0.0044062f $X=8.415 $Y=0.585 $X2=0
+ $Y2=0
cc_639 N_A_1583_285#_c_887_n N_VGND_c_1244_n 0.0191167f $X=9.63 $Y=0.54 $X2=0
+ $Y2=0
cc_640 N_A_1583_285#_M1009_g N_VGND_c_1248_n 0.00426961f $X=10.195 $Y=0.67 $X2=0
+ $Y2=0
cc_641 N_A_1583_285#_M1025_g N_VGND_c_1248_n 0.00482473f $X=10.555 $Y=0.67 $X2=0
+ $Y2=0
cc_642 N_A_1583_285#_M1002_g N_VGND_c_1249_n 0.00544287f $X=8.415 $Y=0.585 $X2=0
+ $Y2=0
cc_643 N_A_1583_285#_M1009_g N_VGND_c_1249_n 0.00434697f $X=10.195 $Y=0.67 $X2=0
+ $Y2=0
cc_644 N_A_1583_285#_M1025_g N_VGND_c_1249_n 0.00517496f $X=10.555 $Y=0.67 $X2=0
+ $Y2=0
cc_645 N_A_1583_285#_c_887_n N_VGND_c_1249_n 0.0164682f $X=9.63 $Y=0.54 $X2=0
+ $Y2=0
cc_646 N_A_1429_383#_c_1002_n N_VPWR_M1005_d 0.00899303f $X=8.185 $Y=2.16 $X2=0
+ $Y2=0
cc_647 N_A_1429_383#_c_994_n N_VPWR_M1005_d 0.0058633f $X=8.27 $Y=2.075 $X2=0
+ $Y2=0
cc_648 N_A_1429_383#_M1017_g N_VPWR_c_1085_n 0.024203f $X=9.21 $Y=2.415 $X2=0
+ $Y2=0
cc_649 N_A_1429_383#_c_1002_n N_VPWR_c_1085_n 0.0114239f $X=8.185 $Y=2.16 $X2=0
+ $Y2=0
cc_650 N_A_1429_383#_c_1001_n N_VPWR_c_1089_n 0.0122551f $X=7.285 $Y=2.24 $X2=0
+ $Y2=0
cc_651 N_A_1429_383#_M1017_g N_VPWR_c_1091_n 0.00908496f $X=9.21 $Y=2.415 $X2=0
+ $Y2=0
cc_652 N_A_1429_383#_M1017_g N_VPWR_c_1081_n 0.00885833f $X=9.21 $Y=2.415 $X2=0
+ $Y2=0
cc_653 N_A_1429_383#_c_1001_n N_VPWR_c_1081_n 0.0116403f $X=7.285 $Y=2.24 $X2=0
+ $Y2=0
cc_654 N_A_1429_383#_c_1002_n A_1535_383# 0.00618217f $X=8.185 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_655 N_A_1429_383#_c_987_n N_VGND_c_1238_n 0.0117341f $X=8.845 $Y=0.905 $X2=0
+ $Y2=0
cc_656 N_A_1429_383#_c_989_n N_VGND_c_1238_n 0.00202084f $X=9.205 $Y=0.905 $X2=0
+ $Y2=0
cc_657 N_A_1429_383#_c_992_n N_VGND_c_1238_n 0.0134127f $X=8.185 $Y=0.52 $X2=0
+ $Y2=0
cc_658 N_A_1429_383#_c_993_n N_VGND_c_1238_n 0.00469993f $X=8.27 $Y=0.995 $X2=0
+ $Y2=0
cc_659 N_A_1429_383#_c_995_n N_VGND_c_1238_n 0.0199133f $X=9.055 $Y=1.08 $X2=0
+ $Y2=0
cc_660 N_A_1429_383#_c_989_n N_VGND_c_1239_n 0.00296068f $X=9.205 $Y=0.905 $X2=0
+ $Y2=0
cc_661 N_A_1429_383#_c_992_n N_VGND_c_1242_n 0.0280653f $X=8.185 $Y=0.52 $X2=0
+ $Y2=0
cc_662 N_A_1429_383#_c_987_n N_VGND_c_1244_n 0.00379792f $X=8.845 $Y=0.905 $X2=0
+ $Y2=0
cc_663 N_A_1429_383#_c_989_n N_VGND_c_1244_n 0.00429444f $X=9.205 $Y=0.905 $X2=0
+ $Y2=0
cc_664 N_A_1429_383#_c_987_n N_VGND_c_1249_n 0.00457201f $X=8.845 $Y=0.905 $X2=0
+ $Y2=0
cc_665 N_A_1429_383#_c_989_n N_VGND_c_1249_n 0.00544287f $X=9.205 $Y=0.905 $X2=0
+ $Y2=0
cc_666 N_A_1429_383#_c_992_n N_VGND_c_1249_n 0.0225369f $X=8.185 $Y=0.52 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_1083_n N_A_629_125#_c_1177_n 0.0150944f $X=2.705 $Y=2.195 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_1094_n N_A_629_125#_c_1177_n 0.00714332f $X=5.36 $Y=3.33 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_1081_n N_A_629_125#_c_1177_n 0.00891647f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_1086_n N_Q_c_1219_n 0.0685263f $X=10.23 $Y=2.125 $X2=0 $Y2=0
cc_671 N_VPWR_c_1095_n N_Q_c_1219_n 0.0158357f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_672 N_VPWR_c_1081_n N_Q_c_1219_n 0.0121432f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_673 N_A_629_125#_c_1173_n N_VGND_c_1236_n 0.0110928f $X=3.365 $Y=0.705 $X2=0
+ $Y2=0
cc_674 N_A_629_125#_c_1173_n N_VGND_c_1247_n 0.013258f $X=3.365 $Y=0.705 $X2=0
+ $Y2=0
cc_675 N_A_629_125#_c_1173_n N_VGND_c_1249_n 0.0106015f $X=3.365 $Y=0.705 $X2=0
+ $Y2=0
cc_676 Q N_VGND_c_1239_n 0.015392f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_677 Q N_VGND_c_1248_n 0.0109624f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_678 Q N_VGND_c_1249_n 0.0117517f $X=10.715 $Y=0.47 $X2=0 $Y2=0
