* File: sky130_fd_sc_lp__xnor3_lp.spice
* Created: Wed Sep  2 10:40:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xnor3_lp.pex.spice"
.subckt sky130_fd_sc_lp__xnor3_lp  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 A_114_109# N_A_M1004_g N_A_27_109#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_M1018_g A_114_109# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1020 A_272_109# N_A_27_109#_M1020_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_A_265_409#_M1015_d N_A_27_109#_M1015_g A_272_109# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 A_570_101# N_B_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1021 N_A_647_367#_M1021_d N_B_M1021_g A_570_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.1533 AS=0.0504 PD=1.57 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1008 N_A_265_409#_M1008_d N_A_647_367#_M1008_g N_A_803_81#_M1008_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0756 AS=0.411 PD=0.78 PS=2.85 NRD=0 NRS=263.868 M=1 R=2.8
+ SA=75000.6 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1026 N_A_763_347#_M1026_d N_B_M1026_g N_A_265_409#_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.09485 AS=0.0756 PD=1 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1023 N_A_27_109#_M1023_d N_A_647_367#_M1023_g N_A_763_347#_M1026_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.09485 PD=0.7 PS=1 NRD=0 NRS=48.804 M=1 R=2.8
+ SA=75000.8 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_803_81#_M1025_d N_B_M1025_g N_A_27_109#_M1023_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0714 AS=0.0588 PD=0.76 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_1348_111#_M1002_d N_A_1318_85#_M1002_g N_A_803_81#_M1025_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0714 PD=0.7 PS=0.76 NRD=0 NRS=17.136 M=1 R=2.8
+ SA=75001.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_763_347#_M1005_d N_C_M1005_g N_A_1348_111#_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 A_1634_89# N_C_M1017_g N_A_1318_85#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0870625 AS=0.1197 PD=0.96 PS=1.41 NRD=43.5 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_C_M1009_g A_1634_89# VNB NSHORT L=0.15 W=0.42 AD=0.10605
+ AS=0.0870625 PD=0.925 PS=0.96 NRD=64.284 NRS=43.5 M=1 R=2.8 SA=75000.4
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1001 A_1860_132# N_A_1348_111#_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.10605 PD=0.63 PS=0.925 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_X_M1019_d N_A_1348_111#_M1019_g A_1860_132# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_A_M1024_g N_A_27_109#_M1024_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1010 N_A_265_409#_M1010_d N_A_27_109#_M1010_g N_VPWR_M1024_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1003 N_A_647_367#_M1003_d N_B_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.3853 PD=2.57 PS=2.87 NRD=0 NRS=16.7253 M=1 R=4 SA=125000
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1011 N_A_265_409#_M1011_d N_A_647_367#_M1011_g N_A_763_347#_M1011_s VPB
+ PHIGHVT L=0.25 W=1 AD=0.305 AS=0.3911 PD=1.61 PS=2.91 NRD=0 NRS=16.7253 M=1
+ R=4 SA=125000 SB=125003 A=0.25 P=2.5 MULT=1
MM1014 N_A_803_81#_M1014_d N_B_M1014_g N_A_265_409#_M1011_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.305 PD=1.28 PS=1.61 NRD=0 NRS=65.01 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1006 N_A_27_109#_M1006_d N_A_647_367#_M1006_g N_A_803_81#_M1014_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1016 N_A_763_347#_M1016_d N_B_M1016_g N_A_27_109#_M1006_d VPB PHIGHVT L=0.25
+ W=1 AD=0.186125 AS=0.14 PD=1.43 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1007 N_A_1348_111#_M1007_d N_A_1318_85#_M1007_g N_A_763_347#_M1016_d VPB
+ PHIGHVT L=0.25 W=1 AD=0.14 AS=0.186125 PD=1.28 PS=1.43 NRD=0 NRS=16.7253 M=1
+ R=4 SA=125003 SB=125001 A=0.25 P=2.5 MULT=1
MM1022 N_A_803_81#_M1022_d N_C_M1022_g N_A_1348_111#_M1007_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_A_1318_85#_M1000_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1013 N_X_M1013_d N_A_1348_111#_M1013_g N_VPWR_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX27_noxref VNB VPB NWDIODE A=20.0571 P=24.99
c_99 VNB 0 1.41873e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__xnor3_lp.pxi.spice"
*
.ends
*
*
