* File: sky130_fd_sc_lp__o221a_lp.spice
* Created: Fri Aug 28 11:07:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o221a_lp  VNB VPB A1 A2 B2 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* B2	B2
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 A_114_47# N_A_84_21#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_84_21#_M1009_g A_114_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_A_272_47#_M1003_d N_A1_M1003_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_272_47#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1797 AS=0.0588 PD=1.76 PS=0.7 NRD=24.276 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1007 N_A_272_47#_M1007_d N_B2_M1007_g N_A_490_141#_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0839125 AS=0.1176 PD=0.875 PS=1.4 NRD=24.276 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1011 N_A_490_141#_M1011_d N_B1_M1011_g N_A_272_47#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0839125 PD=0.7 PS=0.875 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_84_21#_M1012_d N_C1_M1012_g N_A_490_141#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_84_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.25 W=1
+ AD=0.1925 AS=0.285 PD=1.385 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1005 A_270_419# N_A1_M1005_g N_VPWR_M1000_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.1925 PD=1.24 PS=1.385 NRD=12.7853 NRS=20.685 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1001 N_A_84_21#_M1001_d N_A2_M1001_g A_270_419# VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.12 PD=1.32 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1008 A_482_419# N_B2_M1008_g N_A_84_21#_M1001_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.16 PD=1.24 PS=1.32 NRD=12.7853 NRS=7.8603 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g A_482_419# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1010 N_A_84_21#_M1010_d N_C1_M1010_g N_VPWR_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=8.7655 P=13.13
c_92 VPB 0 1.41911e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o221a_lp.pxi.spice"
*
.ends
*
*
