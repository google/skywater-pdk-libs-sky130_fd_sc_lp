* NGSPICE file created from sky130_fd_sc_lp__o2bb2ai_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o2bb2ai_m A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_110_535# A2_N a_116_81# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_410_78# B1 VGND VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.289e+11p ps=2.77e+06u
M1002 a_390_535# B2 Y VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1003 a_410_78# a_110_535# Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 VPWR A2_N a_110_535# VPB phighvt w=420000u l=150000u
+  ad=3.864e+11p pd=4.36e+06u as=1.176e+11p ps=1.4e+06u
M1005 VPWR B1 a_390_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_116_81# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_110_535# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_110_535# A1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B2 a_410_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

