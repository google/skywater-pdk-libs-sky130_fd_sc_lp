* File: sky130_fd_sc_lp__dfrtp_2.spice
* Created: Wed Sep  2 09:43:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfrtp_2.pex.spice"
.subckt sky130_fd_sc_lp__dfrtp_2  VNB VPB CLK D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_CLK_M1009_g N_A_27_101#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.09555 AS=0.1113 PD=0.875 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1021 N_A_196_464#_M1021_d N_A_27_101#_M1021_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1512 AS=0.09555 PD=1.56 PS=0.875 NRD=27.132 NRS=49.992 M=1 R=2.8
+ SA=75000.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1032 A_483_78# N_RESET_B_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.42
+ AD=0.08995 AS=0.1197 PD=0.985 PS=1.41 NRD=45.468 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_318_535#_M1002_d N_D_M1002_g A_483_78# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.08995 PD=0.7 PS=0.985 NRD=0 NRS=45.468 M=1 R=2.8 SA=75000.5
+ SB=75004.9 A=0.063 P=1.14 MULT=1
MM1004 N_A_573_535#_M1004_d N_A_27_101#_M1004_g N_A_318_535#_M1002_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1155 AS=0.0588 PD=0.97 PS=0.7 NRD=77.136 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1023 A_811_119# N_A_196_464#_M1023_g N_A_573_535#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1155 PD=0.63 PS=0.97 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1014 A_883_119# N_A_709_411#_M1014_g A_811_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0852 AS=0.0441 PD=0.87 PS=0.63 NRD=42.24 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_RESET_B_M1027_g A_883_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.159045 AS=0.0852 PD=1.03415 PS=0.87 NRD=34.284 NRS=42.24 M=1 R=2.8
+ SA=75002.2 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1017 N_A_709_411#_M1017_d N_A_573_535#_M1017_g N_VGND_M1027_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1456 AS=0.242355 PD=1.095 PS=1.57585 NRD=0 NRS=50.616 M=1
+ R=4.26667 SA=75002.1 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1020 N_A_1252_451#_M1020_d N_A_196_464#_M1020_g N_A_709_411#_M1017_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.180589 AS=0.1456 PD=1.44906 PS=1.095 NRD=17.808
+ NRS=32.808 M=1 R=4.26667 SA=75002.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1012 A_1399_125# N_A_27_101#_M1012_g N_A_1252_451#_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.118511 PD=0.81 PS=0.950943 NRD=39.996 NRS=27.132 M=1
+ R=2.8 SA=75003.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_1399_473#_M1024_g A_1399_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75004.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1028 A_1593_125# N_RESET_B_M1028_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75004.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_1399_473#_M1018_d N_A_1252_451#_M1018_g A_1593_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75005
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_1252_451#_M1013_g N_A_1836_47#_M1013_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0987 AS=0.1113 PD=0.853333 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1022 N_Q_M1022_d N_A_1836_47#_M1022_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1974 PD=1.12 PS=1.70667 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1025 N_Q_M1022_d N_A_1836_47#_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_CLK_M1003_g N_A_27_101#_M1003_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1019 N_A_196_464#_M1019_d N_A_27_101#_M1019_g N_VPWR_M1003_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_RESET_B_M1001_g N_A_318_535#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1026 N_A_318_535#_M1026_d N_D_M1026_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_573_535#_M1010_d N_A_196_464#_M1010_g N_A_318_535#_M1026_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=18.7544 NRS=0 M=1
+ R=2.8 SA=75001.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 A_667_535# N_A_27_101#_M1006_g N_A_573_535#_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_709_411#_M1008_g A_667_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=11.7215 NRS=23.443 M=1 R=2.8
+ SA=75001.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_A_573_535#_M1011_d N_RESET_B_M1011_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.06405 PD=1.37 PS=0.725 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_709_411#_M1007_d N_A_573_535#_M1007_g N_VPWR_M1007_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.4998 PD=1.12 PS=2.87 NRD=0 NRS=72.693 M=1 R=5.6
+ SA=75000.5 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1030 N_A_1252_451#_M1030_d N_A_27_101#_M1030_g N_A_709_411#_M1007_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1792 AS=0.1176 PD=1.62 PS=1.12 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.9 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1015 A_1357_535# N_A_196_464#_M1015_g N_A_1252_451#_M1030_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0896 PD=0.63 PS=0.81 NRD=23.443 NRS=74.2493 M=1 R=2.8
+ SA=75001.5 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_1399_473#_M1005_g A_1357_535# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.21 AS=0.0441 PD=1.42 PS=0.63 NRD=39.8531 NRS=23.443 M=1 R=2.8
+ SA=75001.8 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1031 N_A_1399_473#_M1031_d N_RESET_B_M1031_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.21 PD=0.7 PS=1.42 NRD=0 NRS=4.6886 M=1 R=2.8 SA=75003
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_VPWR_M1016_d N_A_1252_451#_M1016_g N_A_1399_473#_M1031_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75003.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_1252_451#_M1000_g N_A_1836_47#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.132952 AS=0.1696 PD=1.09137 PS=1.81 NRD=13.0808 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1029 N_Q_M1029_d N_A_1836_47#_M1029_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.261748 PD=1.54 PS=2.14863 NRD=0 NRS=4.1567 M=1 R=8.4 SA=75000.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1033 N_Q_M1029_d N_A_1836_47#_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=21.2983 P=26.57
c_129 VNB 0 1.88632e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dfrtp_2.pxi.spice"
*
.ends
*
*
