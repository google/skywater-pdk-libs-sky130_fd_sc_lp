* File: sky130_fd_sc_lp__sdfsbp_1.pxi.spice
* Created: Fri Aug 28 11:29:09 2020
* 
x_PM_SKY130_FD_SC_LP__SDFSBP_1%SCE N_SCE_c_285_n N_SCE_c_286_n N_SCE_c_287_n
+ N_SCE_M1022_g N_SCE_c_288_n N_SCE_M1013_g N_SCE_M1034_g N_SCE_M1006_g
+ N_SCE_c_295_n N_SCE_c_290_n N_SCE_c_291_n SCE N_SCE_c_298_n N_SCE_c_299_n
+ PM_SKY130_FD_SC_LP__SDFSBP_1%SCE
x_PM_SKY130_FD_SC_LP__SDFSBP_1%D N_D_M1039_g N_D_c_378_n N_D_M1014_g D D D
+ N_D_c_383_n N_D_c_380_n PM_SKY130_FD_SC_LP__SDFSBP_1%D
x_PM_SKY130_FD_SC_LP__SDFSBP_1%A_34_481# N_A_34_481#_M1013_s N_A_34_481#_M1022_s
+ N_A_34_481#_M1032_g N_A_34_481#_c_423_n N_A_34_481#_M1008_g
+ N_A_34_481#_c_425_n N_A_34_481#_c_426_n N_A_34_481#_c_427_n
+ N_A_34_481#_c_428_n N_A_34_481#_c_429_n N_A_34_481#_c_430_n
+ N_A_34_481#_c_431_n PM_SKY130_FD_SC_LP__SDFSBP_1%A_34_481#
x_PM_SKY130_FD_SC_LP__SDFSBP_1%SCD N_SCD_M1011_g N_SCD_c_492_n N_SCD_M1036_g SCD
+ SCD SCD N_SCD_c_495_n N_SCD_c_496_n PM_SKY130_FD_SC_LP__SDFSBP_1%SCD
x_PM_SKY130_FD_SC_LP__SDFSBP_1%CLK N_CLK_c_534_n N_CLK_M1009_g N_CLK_M1023_g CLK
+ CLK CLK PM_SKY130_FD_SC_LP__SDFSBP_1%CLK
x_PM_SKY130_FD_SC_LP__SDFSBP_1%A_901_441# N_A_901_441#_M1026_d
+ N_A_901_441#_M1017_d N_A_901_441#_M1018_g N_A_901_441#_M1025_g
+ N_A_901_441#_c_575_n N_A_901_441#_M1038_g N_A_901_441#_M1012_g
+ N_A_901_441#_c_576_n N_A_901_441#_c_577_n N_A_901_441#_c_578_n
+ N_A_901_441#_c_579_n N_A_901_441#_c_580_n N_A_901_441#_c_595_n
+ N_A_901_441#_c_581_n N_A_901_441#_c_582_n N_A_901_441#_c_583_n
+ N_A_901_441#_c_597_n N_A_901_441#_c_607_p N_A_901_441#_c_584_n
+ N_A_901_441#_c_612_p N_A_901_441#_c_585_n N_A_901_441#_c_586_n
+ N_A_901_441#_c_587_n PM_SKY130_FD_SC_LP__SDFSBP_1%A_901_441#
x_PM_SKY130_FD_SC_LP__SDFSBP_1%A_1274_401# N_A_1274_401#_M1005_s
+ N_A_1274_401#_M1004_d N_A_1274_401#_M1031_g N_A_1274_401#_M1015_g
+ N_A_1274_401#_c_745_n N_A_1274_401#_c_738_n N_A_1274_401#_c_746_n
+ N_A_1274_401#_c_747_n N_A_1274_401#_c_739_n N_A_1274_401#_c_740_n
+ N_A_1274_401#_c_741_n N_A_1274_401#_c_766_n N_A_1274_401#_c_748_n
+ N_A_1274_401#_c_749_n N_A_1274_401#_c_742_n N_A_1274_401#_c_751_n
+ PM_SKY130_FD_SC_LP__SDFSBP_1%A_1274_401#
x_PM_SKY130_FD_SC_LP__SDFSBP_1%A_1146_463# N_A_1146_463#_M1024_d
+ N_A_1146_463#_M1018_d N_A_1146_463#_M1004_g N_A_1146_463#_c_868_n
+ N_A_1146_463#_c_869_n N_A_1146_463#_M1005_g N_A_1146_463#_c_870_n
+ N_A_1146_463#_M1019_g N_A_1146_463#_c_871_n N_A_1146_463#_M1029_g
+ N_A_1146_463#_c_872_n N_A_1146_463#_c_873_n N_A_1146_463#_c_887_n
+ N_A_1146_463#_c_904_n N_A_1146_463#_c_874_n N_A_1146_463#_c_875_n
+ N_A_1146_463#_c_876_n N_A_1146_463#_c_877_n N_A_1146_463#_c_878_n
+ N_A_1146_463#_c_879_n N_A_1146_463#_c_880_n N_A_1146_463#_c_881_n
+ N_A_1146_463#_c_882_n N_A_1146_463#_c_889_n N_A_1146_463#_c_927_n
+ PM_SKY130_FD_SC_LP__SDFSBP_1%A_1146_463#
x_PM_SKY130_FD_SC_LP__SDFSBP_1%SET_B N_SET_B_c_1012_n N_SET_B_M1010_g
+ N_SET_B_c_1014_n N_SET_B_M1041_g N_SET_B_M1028_g N_SET_B_c_1009_n
+ N_SET_B_c_1010_n N_SET_B_M1003_g N_SET_B_c_1017_n N_SET_B_c_1018_n
+ N_SET_B_c_1019_n SET_B N_SET_B_c_1021_n N_SET_B_c_1022_n N_SET_B_c_1011_n
+ PM_SKY130_FD_SC_LP__SDFSBP_1%SET_B
x_PM_SKY130_FD_SC_LP__SDFSBP_1%A_640_481# N_A_640_481#_M1023_d
+ N_A_640_481#_M1009_d N_A_640_481#_c_1124_n N_A_640_481#_c_1125_n
+ N_A_640_481#_M1017_g N_A_640_481#_c_1139_n N_A_640_481#_c_1140_n
+ N_A_640_481#_M1026_g N_A_640_481#_c_1128_n N_A_640_481#_c_1129_n
+ N_A_640_481#_M1024_g N_A_640_481#_c_1131_n N_A_640_481#_M1000_g
+ N_A_640_481#_c_1142_n N_A_640_481#_M1040_g N_A_640_481#_M1030_g
+ N_A_640_481#_c_1133_n N_A_640_481#_c_1134_n N_A_640_481#_c_1144_n
+ N_A_640_481#_c_1231_p N_A_640_481#_c_1135_n N_A_640_481#_c_1145_n
+ N_A_640_481#_c_1146_n N_A_640_481#_c_1136_n N_A_640_481#_c_1137_n
+ PM_SKY130_FD_SC_LP__SDFSBP_1%A_640_481#
x_PM_SKY130_FD_SC_LP__SDFSBP_1%A_2067_92# N_A_2067_92#_M1033_s
+ N_A_2067_92#_M1016_s N_A_2067_92#_M1035_g N_A_2067_92#_M1001_g
+ N_A_2067_92#_c_1261_n N_A_2067_92#_c_1262_n N_A_2067_92#_c_1263_n
+ N_A_2067_92#_c_1264_n N_A_2067_92#_c_1270_n N_A_2067_92#_c_1265_n
+ N_A_2067_92#_c_1272_n PM_SKY130_FD_SC_LP__SDFSBP_1%A_2067_92#
x_PM_SKY130_FD_SC_LP__SDFSBP_1%A_1920_119# N_A_1920_119#_M1038_d
+ N_A_1920_119#_M1040_d N_A_1920_119#_M1003_d N_A_1920_119#_M1033_g
+ N_A_1920_119#_c_1341_n N_A_1920_119#_c_1342_n N_A_1920_119#_M1016_g
+ N_A_1920_119#_c_1360_n N_A_1920_119#_M1002_g N_A_1920_119#_c_1344_n
+ N_A_1920_119#_c_1345_n N_A_1920_119#_c_1361_n N_A_1920_119#_M1037_g
+ N_A_1920_119#_M1007_g N_A_1920_119#_M1021_g N_A_1920_119#_c_1346_n
+ N_A_1920_119#_c_1376_n N_A_1920_119#_c_1347_n N_A_1920_119#_c_1365_n
+ N_A_1920_119#_c_1366_n N_A_1920_119#_c_1367_n N_A_1920_119#_c_1368_n
+ N_A_1920_119#_c_1369_n N_A_1920_119#_c_1348_n N_A_1920_119#_c_1371_n
+ N_A_1920_119#_c_1349_n N_A_1920_119#_c_1350_n N_A_1920_119#_c_1351_n
+ N_A_1920_119#_c_1352_n N_A_1920_119#_c_1353_n N_A_1920_119#_c_1354_n
+ N_A_1920_119#_c_1374_n N_A_1920_119#_c_1441_p N_A_1920_119#_c_1355_n
+ N_A_1920_119#_c_1375_n N_A_1920_119#_c_1356_n
+ PM_SKY130_FD_SC_LP__SDFSBP_1%A_1920_119#
x_PM_SKY130_FD_SC_LP__SDFSBP_1%A_2582_150# N_A_2582_150#_M1002_d
+ N_A_2582_150#_M1037_d N_A_2582_150#_c_1545_n N_A_2582_150#_c_1546_n
+ N_A_2582_150#_M1020_g N_A_2582_150#_M1027_g N_A_2582_150#_c_1548_n
+ N_A_2582_150#_c_1549_n N_A_2582_150#_c_1550_n N_A_2582_150#_c_1551_n
+ N_A_2582_150#_c_1554_n N_A_2582_150#_c_1552_n N_A_2582_150#_c_1556_n
+ PM_SKY130_FD_SC_LP__SDFSBP_1%A_2582_150#
x_PM_SKY130_FD_SC_LP__SDFSBP_1%VPWR N_VPWR_M1022_d N_VPWR_M1011_d N_VPWR_M1017_s
+ N_VPWR_M1031_d N_VPWR_M1010_d N_VPWR_M1001_d N_VPWR_M1016_d N_VPWR_M1027_d
+ N_VPWR_c_1609_n N_VPWR_c_1610_n N_VPWR_c_1611_n N_VPWR_c_1612_n
+ N_VPWR_c_1613_n N_VPWR_c_1614_n N_VPWR_c_1615_n N_VPWR_c_1616_n
+ N_VPWR_c_1617_n N_VPWR_c_1618_n N_VPWR_c_1619_n N_VPWR_c_1620_n
+ N_VPWR_c_1621_n VPWR N_VPWR_c_1622_n N_VPWR_c_1623_n N_VPWR_c_1624_n
+ N_VPWR_c_1625_n N_VPWR_c_1626_n N_VPWR_c_1627_n N_VPWR_c_1608_n
+ N_VPWR_c_1629_n N_VPWR_c_1630_n N_VPWR_c_1631_n N_VPWR_c_1632_n
+ N_VPWR_c_1633_n PM_SKY130_FD_SC_LP__SDFSBP_1%VPWR
x_PM_SKY130_FD_SC_LP__SDFSBP_1%A_275_481# N_A_275_481#_M1014_d
+ N_A_275_481#_M1024_s N_A_275_481#_M1039_d N_A_275_481#_M1018_s
+ N_A_275_481#_c_1770_n N_A_275_481#_c_1785_n N_A_275_481#_c_1771_n
+ N_A_275_481#_c_1772_n N_A_275_481#_c_1806_n N_A_275_481#_c_1776_n
+ N_A_275_481#_c_1777_n N_A_275_481#_c_1778_n N_A_275_481#_c_1773_n
+ N_A_275_481#_c_1788_n N_A_275_481#_c_1816_n N_A_275_481#_c_1779_n
+ N_A_275_481#_c_1780_n N_A_275_481#_c_1774_n
+ PM_SKY130_FD_SC_LP__SDFSBP_1%A_275_481#
x_PM_SKY130_FD_SC_LP__SDFSBP_1%Q N_Q_M1020_s N_Q_M1027_s Q Q Q Q Q N_Q_c_1898_n
+ PM_SKY130_FD_SC_LP__SDFSBP_1%Q
x_PM_SKY130_FD_SC_LP__SDFSBP_1%Q_N N_Q_N_M1021_d N_Q_N_M1007_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N Q_N PM_SKY130_FD_SC_LP__SDFSBP_1%Q_N
x_PM_SKY130_FD_SC_LP__SDFSBP_1%VGND N_VGND_M1013_d N_VGND_M1036_d N_VGND_M1026_s
+ N_VGND_M1015_d N_VGND_M1041_d N_VGND_M1028_d N_VGND_M1033_d N_VGND_M1020_d
+ N_VGND_c_1931_n N_VGND_c_1932_n N_VGND_c_1933_n N_VGND_c_1934_n
+ N_VGND_c_1935_n N_VGND_c_1936_n N_VGND_c_1937_n N_VGND_c_1938_n
+ N_VGND_c_1939_n N_VGND_c_1940_n N_VGND_c_1941_n N_VGND_c_1942_n
+ N_VGND_c_1943_n N_VGND_c_1944_n N_VGND_c_1945_n N_VGND_c_1946_n
+ N_VGND_c_1947_n N_VGND_c_1948_n VGND N_VGND_c_1949_n N_VGND_c_1950_n
+ N_VGND_c_1951_n N_VGND_c_1952_n N_VGND_c_1953_n N_VGND_c_1954_n
+ N_VGND_c_1955_n N_VGND_c_1956_n PM_SKY130_FD_SC_LP__SDFSBP_1%VGND
cc_1 VNB N_SCE_c_285_n 0.0458062f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.915
cc_2 VNB N_SCE_c_286_n 0.0270247f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.84
cc_3 VNB N_SCE_c_287_n 0.0109511f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=0.84
cc_4 VNB N_SCE_c_288_n 0.019598f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.765
cc_5 VNB N_SCE_M1006_g 0.0308306f $X=-0.19 $Y=-0.245 $X2=2.315 $Y2=0.445
cc_6 VNB N_SCE_c_290_n 0.00152356f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_7 VNB N_SCE_c_291_n 0.0515753f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_8 VNB N_D_c_378_n 0.0184213f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.245
cc_9 VNB D 0.0323544f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.445
cc_10 VNB N_D_c_380_n 0.0363633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_34_481#_M1032_g 0.0336969f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.765
cc_12 VNB N_A_34_481#_c_423_n 0.0318282f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.445
cc_13 VNB N_A_34_481#_M1008_g 0.0108967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_34_481#_c_425_n 0.0474204f $X=-0.19 $Y=-0.245 $X2=2.315 $Y2=0.445
cc_15 VNB N_A_34_481#_c_426_n 0.0140785f $X=-0.19 $Y=-0.245 $X2=2.315 $Y2=0.445
cc_16 VNB N_A_34_481#_c_427_n 0.028422f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_17 VNB N_A_34_481#_c_428_n 0.0144057f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.21
cc_18 VNB N_A_34_481#_c_429_n 0.00443619f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_19 VNB N_A_34_481#_c_430_n 0.019059f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=2.08
cc_20 VNB N_A_34_481#_c_431_n 0.0135197f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.08
cc_21 VNB N_SCD_M1036_g 0.05676f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.765
cc_22 VNB SCD 0.00466122f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.445
cc_23 VNB N_CLK_c_534_n 0.0906264f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.915
cc_24 VNB N_CLK_M1023_g 0.0250855f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.725
cc_25 VNB CLK 0.0106855f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.765
cc_26 VNB N_A_901_441#_M1025_g 0.0275385f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.725
cc_27 VNB N_A_901_441#_c_575_n 0.0161471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_901_441#_c_576_n 0.0521398f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.21
cc_29 VNB N_A_901_441#_c_577_n 0.00747833f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=2.125
cc_30 VNB N_A_901_441#_c_578_n 0.0261734f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.16
cc_31 VNB N_A_901_441#_c_579_n 0.00966289f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_32 VNB N_A_901_441#_c_580_n 0.0296954f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_33 VNB N_A_901_441#_c_581_n 0.0223734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_901_441#_c_582_n 0.0341531f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.08
cc_35 VNB N_A_901_441#_c_583_n 0.00273757f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.08
cc_36 VNB N_A_901_441#_c_584_n 4.80011e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_901_441#_c_585_n 0.00555509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_901_441#_c_586_n 0.00748171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_901_441#_c_587_n 9.99738e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1274_401#_M1015_g 0.0414397f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.725
cc_41 VNB N_A_1274_401#_c_738_n 0.00215173f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_42 VNB N_A_1274_401#_c_739_n 0.00159693f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_43 VNB N_A_1274_401#_c_740_n 0.0141772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1274_401#_c_741_n 0.00314317f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_45 VNB N_A_1274_401#_c_742_n 0.00362627f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.08
cc_46 VNB N_A_1146_463#_M1004_g 0.0273134f $X=-0.19 $Y=-0.245 $X2=0.755
+ $Y2=0.765
cc_47 VNB N_A_1146_463#_c_868_n 0.0318112f $X=-0.19 $Y=-0.245 $X2=0.755
+ $Y2=0.445
cc_48 VNB N_A_1146_463#_c_869_n 0.0160009f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.725
cc_49 VNB N_A_1146_463#_c_870_n 0.0198132f $X=-0.19 $Y=-0.245 $X2=2.315
+ $Y2=0.995
cc_50 VNB N_A_1146_463#_c_871_n 0.0181597f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_51 VNB N_A_1146_463#_c_872_n 0.0129593f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=2.125
cc_52 VNB N_A_1146_463#_c_873_n 0.0319086f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_53 VNB N_A_1146_463#_c_874_n 0.0191758f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.08
cc_54 VNB N_A_1146_463#_c_875_n 0.0056084f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.08
cc_55 VNB N_A_1146_463#_c_876_n 0.00139438f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=2.105
cc_56 VNB N_A_1146_463#_c_877_n 0.052521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1146_463#_c_878_n 0.0128609f $X=-0.19 $Y=-0.245 $X2=0.935
+ $Y2=2.105
cc_58 VNB N_A_1146_463#_c_879_n 0.00448617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1146_463#_c_880_n 8.28295e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1146_463#_c_881_n 0.00257089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1146_463#_c_882_n 0.0028204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_SET_B_M1041_g 0.0477156f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.765
cc_63 VNB N_SET_B_M1028_g 0.0202204f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.725
cc_64 VNB N_SET_B_c_1009_n 0.0374443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_SET_B_c_1010_n 0.00747509f $X=-0.19 $Y=-0.245 $X2=2.315 $Y2=0.995
cc_66 VNB N_SET_B_c_1011_n 0.0231757f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.08
cc_67 VNB N_A_640_481#_c_1124_n 0.0335459f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.725
cc_68 VNB N_A_640_481#_c_1125_n 0.0196048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_640_481#_M1017_g 0.00486961f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.245
cc_70 VNB N_A_640_481#_M1026_g 0.0161285f $X=-0.19 $Y=-0.245 $X2=2.315 $Y2=0.445
cc_71 VNB N_A_640_481#_c_1128_n 0.0709025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_640_481#_c_1129_n 0.0125016f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_73 VNB N_A_640_481#_M1024_g 0.0396722f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.21
cc_74 VNB N_A_640_481#_c_1131_n 0.328873f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.16
cc_75 VNB N_A_640_481#_M1030_g 0.0355085f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.08
cc_76 VNB N_A_640_481#_c_1133_n 0.0409981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_640_481#_c_1134_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_640_481#_c_1135_n 0.0232176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_640_481#_c_1136_n 0.00710829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_640_481#_c_1137_n 0.0257416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_2067_92#_M1035_g 0.0427304f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.765
cc_82 VNB N_A_2067_92#_c_1261_n 0.00420943f $X=-0.19 $Y=-0.245 $X2=2.315
+ $Y2=0.995
cc_83 VNB N_A_2067_92#_c_1262_n 0.00646271f $X=-0.19 $Y=-0.245 $X2=2.315
+ $Y2=0.445
cc_84 VNB N_A_2067_92#_c_1263_n 0.0229676f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_85 VNB N_A_2067_92#_c_1264_n 0.0114804f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=2.125
cc_86 VNB N_A_2067_92#_c_1265_n 0.00618256f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_87 VNB N_A_1920_119#_M1033_g 0.0469979f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.245
cc_88 VNB N_A_1920_119#_c_1341_n 0.012623f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.725
cc_89 VNB N_A_1920_119#_c_1342_n 0.00209167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1920_119#_M1002_g 0.034379f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.16
cc_91 VNB N_A_1920_119#_c_1344_n 0.0292861f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_92 VNB N_A_1920_119#_c_1345_n 0.0108925f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_93 VNB N_A_1920_119#_c_1346_n 0.0158104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1920_119#_c_1347_n 0.0049629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1920_119#_c_1348_n 0.00897668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1920_119#_c_1349_n 0.0136972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1920_119#_c_1350_n 0.00601058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1920_119#_c_1351_n 0.00331826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1920_119#_c_1352_n 0.00528053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1920_119#_c_1353_n 9.68688e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1920_119#_c_1354_n 0.0317953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1920_119#_c_1355_n 0.0733976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1920_119#_c_1356_n 0.021038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2582_150#_c_1545_n 0.0330666f $X=-0.19 $Y=-0.245 $X2=0.755
+ $Y2=0.765
cc_105 VNB N_A_2582_150#_c_1546_n 0.0190088f $X=-0.19 $Y=-0.245 $X2=0.755
+ $Y2=0.445
cc_106 VNB N_A_2582_150#_M1027_g 0.00861335f $X=-0.19 $Y=-0.245 $X2=2.315
+ $Y2=0.995
cc_107 VNB N_A_2582_150#_c_1548_n 0.0049727f $X=-0.19 $Y=-0.245 $X2=2.315
+ $Y2=0.445
cc_108 VNB N_A_2582_150#_c_1549_n 0.0109021f $X=-0.19 $Y=-0.245 $X2=2.29
+ $Y2=0.995
cc_109 VNB N_A_2582_150#_c_1550_n 0.0104789f $X=-0.19 $Y=-0.245 $X2=0.935
+ $Y2=2.21
cc_110 VNB N_A_2582_150#_c_1551_n 0.00340522f $X=-0.19 $Y=-0.245 $X2=2.25
+ $Y2=2.125
cc_111 VNB N_A_2582_150#_c_1552_n 0.0415955f $X=-0.19 $Y=-0.245 $X2=0.29
+ $Y2=2.08
cc_112 VNB N_VPWR_c_1608_n 0.641339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_275_481#_c_1770_n 0.00436961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_275_481#_c_1771_n 0.00945716f $X=-0.19 $Y=-0.245 $X2=2.29
+ $Y2=0.995
cc_115 VNB N_A_275_481#_c_1772_n 0.0122203f $X=-0.19 $Y=-0.245 $X2=2.25
+ $Y2=2.125
cc_116 VNB N_A_275_481#_c_1773_n 0.00994243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_275_481#_c_1774_n 0.00713377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_Q_c_1898_n 0.00788785f $X=-0.19 $Y=-0.245 $X2=2.315 $Y2=0.445
cc_119 VNB Q_N 0.0570191f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.725
cc_120 VNB N_VGND_c_1931_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.16
cc_121 VNB N_VGND_c_1932_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1933_n 0.0110269f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.08
cc_123 VNB N_VGND_c_1934_n 0.0216655f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=2.08
cc_124 VNB N_VGND_c_1935_n 0.0194558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1936_n 0.0302705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1937_n 0.0442513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1938_n 0.010023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1939_n 0.0221938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1940_n 0.00436868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1941_n 0.0409845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1942_n 0.00436274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1943_n 0.0295069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1944_n 0.00461634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1945_n 0.0580412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1946_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1947_n 0.0510728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1948_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1949_n 0.0537103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1950_n 0.0238029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1951_n 0.0521376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1952_n 0.0191001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1953_n 0.769324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1954_n 0.00266338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1955_n 0.0106753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_1956_n 0.00631708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VPB N_SCE_c_285_n 0.0164004f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.915
cc_147 VPB N_SCE_M1022_g 0.0216094f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.725
cc_148 VPB N_SCE_M1034_g 0.017757f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.725
cc_149 VPB N_SCE_c_295_n 0.029818f $X=-0.19 $Y=1.655 $X2=2.125 $Y2=2.21
cc_150 VPB N_SCE_c_290_n 0.00616961f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_151 VPB N_SCE_c_291_n 0.00690798f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_152 VPB N_SCE_c_298_n 0.0706652f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.08
cc_153 VPB N_SCE_c_299_n 0.00260306f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.105
cc_154 VPB N_D_M1039_g 0.0302745f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.84
cc_155 VPB D 0.0170954f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=0.445
cc_156 VPB N_D_c_383_n 0.0313853f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=0.995
cc_157 VPB N_A_34_481#_M1008_g 0.0521799f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_34_481#_c_428_n 0.0648823f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.21
cc_159 VPB N_SCD_M1011_g 0.0245242f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.84
cc_160 VPB N_SCD_c_492_n 0.00696162f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.725
cc_161 VPB N_SCD_M1036_g 0.013332f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=0.765
cc_162 VPB SCD 0.00375957f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=0.445
cc_163 VPB N_SCD_c_495_n 0.0128038f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_164 VPB N_SCD_c_496_n 0.0392018f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=0.995
cc_165 VPB N_CLK_c_534_n 0.00275643f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=0.915
cc_166 VPB N_CLK_M1009_g 0.0642226f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.84
cc_167 VPB CLK 0.0125741f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=0.765
cc_168 VPB N_A_901_441#_M1018_g 0.0283941f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=0.765
cc_169 VPB N_A_901_441#_M1012_g 0.0464654f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_170 VPB N_A_901_441#_c_576_n 0.0584987f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.21
cc_171 VPB N_A_901_441#_c_577_n 0.0142394f $X=-0.19 $Y=1.655 $X2=2.25 $Y2=2.125
cc_172 VPB N_A_901_441#_c_578_n 0.0154457f $X=-0.19 $Y=1.655 $X2=2.25 $Y2=1.16
cc_173 VPB N_A_901_441#_c_579_n 0.00350479f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_174 VPB N_A_901_441#_c_580_n 0.0104032f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_175 VPB N_A_901_441#_c_595_n 0.0080662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_901_441#_c_583_n 0.00293772f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.08
cc_177 VPB N_A_901_441#_c_597_n 0.0139277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_901_441#_c_584_n 0.00367374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_901_441#_c_587_n 0.00468504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_1274_401#_M1031_g 0.0187323f $X=-0.19 $Y=1.655 $X2=0.755
+ $Y2=0.765
cc_181 VPB N_A_1274_401#_M1015_g 0.011408f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.725
cc_182 VPB N_A_1274_401#_c_745_n 0.0118339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_1274_401#_c_746_n 0.0076873f $X=-0.19 $Y=1.655 $X2=2.25 $Y2=2.125
cc_184 VPB N_A_1274_401#_c_747_n 0.0104643f $X=-0.19 $Y=1.655 $X2=2.25 $Y2=1.16
cc_185 VPB N_A_1274_401#_c_748_n 0.00705287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_1274_401#_c_749_n 0.00224442f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=2.08
cc_187 VPB N_A_1274_401#_c_742_n 0.00417159f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.08
cc_188 VPB N_A_1274_401#_c_751_n 0.0427821f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.105
cc_189 VPB N_A_1146_463#_M1004_g 0.0435082f $X=-0.19 $Y=1.655 $X2=0.755
+ $Y2=0.765
cc_190 VPB N_A_1146_463#_c_870_n 8.04604e-19 $X=-0.19 $Y=1.655 $X2=2.315
+ $Y2=0.995
cc_191 VPB N_A_1146_463#_M1019_g 0.0254638f $X=-0.19 $Y=1.655 $X2=2.315
+ $Y2=0.445
cc_192 VPB N_A_1146_463#_c_873_n 0.0132814f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_193 VPB N_A_1146_463#_c_887_n 0.00321931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_1146_463#_c_882_n 0.0018805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_1146_463#_c_889_n 0.00481975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_SET_B_c_1012_n 0.0190382f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=0.915
cc_197 VPB N_SET_B_M1010_g 0.0250843f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.84
cc_198 VPB N_SET_B_c_1014_n 0.0588736f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.245
cc_199 VPB N_SET_B_M1041_g 0.00885389f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=0.765
cc_200 VPB N_SET_B_M1003_g 0.0293687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_SET_B_c_1017_n 0.021105f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.21
cc_202 VPB N_SET_B_c_1018_n 0.00326753f $X=-0.19 $Y=1.655 $X2=2.25 $Y2=2.125
cc_203 VPB N_SET_B_c_1019_n 0.0033743f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_204 VPB SET_B 0.00464402f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_205 VPB N_SET_B_c_1021_n 0.0386189f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.08
cc_206 VPB N_SET_B_c_1022_n 0.0128223f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.08
cc_207 VPB N_SET_B_c_1011_n 0.0129875f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.08
cc_208 VPB N_A_640_481#_M1017_g 0.0523731f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.245
cc_209 VPB N_A_640_481#_c_1139_n 0.106382f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.725
cc_210 VPB N_A_640_481#_c_1140_n 0.0125039f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.725
cc_211 VPB N_A_640_481#_M1000_g 0.0348934f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_212 VPB N_A_640_481#_c_1142_n 0.254826f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_640_481#_M1040_g 0.0245335f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.08
cc_214 VPB N_A_640_481#_c_1144_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_640_481#_c_1145_n 0.0186213f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_640_481#_c_1146_n 0.00532581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_640_481#_c_1136_n 0.0220009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_2067_92#_M1001_g 0.0451249f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.725
cc_219 VPB N_A_2067_92#_c_1261_n 0.00456285f $X=-0.19 $Y=1.655 $X2=2.315
+ $Y2=0.995
cc_220 VPB N_A_2067_92#_c_1262_n 0.00212064f $X=-0.19 $Y=1.655 $X2=2.315
+ $Y2=0.445
cc_221 VPB N_A_2067_92#_c_1263_n 0.0247656f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_222 VPB N_A_2067_92#_c_1270_n 0.0162368f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_223 VPB N_A_2067_92#_c_1265_n 0.014945f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_224 VPB N_A_2067_92#_c_1272_n 0.00420999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1920_119#_c_1341_n 0.0190844f $X=-0.19 $Y=1.655 $X2=0.94
+ $Y2=2.725
cc_226 VPB N_A_1920_119#_c_1342_n 0.0070161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_1920_119#_M1016_g 0.0238177f $X=-0.19 $Y=1.655 $X2=2.315
+ $Y2=0.445
cc_228 VPB N_A_1920_119#_c_1360_n 0.0414424f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_229 VPB N_A_1920_119#_c_1361_n 0.0173918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_1920_119#_M1007_g 0.0228386f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=2.08
cc_231 VPB N_A_1920_119#_c_1346_n 0.0108638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_1920_119#_c_1347_n 0.00388752f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_1920_119#_c_1365_n 0.0117281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_1920_119#_c_1366_n 0.00655825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_1920_119#_c_1367_n 0.00641481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_1920_119#_c_1368_n 0.0266397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_1920_119#_c_1369_n 0.00477129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_1920_119#_c_1348_n 0.00979629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_1920_119#_c_1371_n 0.00335887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_1920_119#_c_1353_n 0.00138473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_1920_119#_c_1354_n 0.00795285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_1920_119#_c_1374_n 0.016727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1920_119#_c_1375_n 0.0266133f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_2582_150#_M1027_g 0.0231525f $X=-0.19 $Y=1.655 $X2=2.315
+ $Y2=0.995
cc_245 VPB N_A_2582_150#_c_1554_n 0.020213f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_246 VPB N_A_2582_150#_c_1552_n 0.0256853f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=2.08
cc_247 VPB N_A_2582_150#_c_1556_n 0.00683501f $X=-0.19 $Y=1.655 $X2=0.51
+ $Y2=2.08
cc_248 VPB N_VPWR_c_1609_n 0.00177638f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_249 VPB N_VPWR_c_1610_n 0.00727945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1611_n 0.013013f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.08
cc_251 VPB N_VPWR_c_1612_n 0.0146292f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.08
cc_252 VPB N_VPWR_c_1613_n 0.00481217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1614_n 0.0614402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1615_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1616_n 0.0159261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1617_n 0.0216781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1618_n 0.0397179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1619_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1620_n 0.0367709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1621_n 0.00362723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1622_n 0.0168658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1623_n 0.0421485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1624_n 0.0291278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1625_n 0.00668967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1626_n 0.0457681f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1627_n 0.0217301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1608_n 0.133661f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1629_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1630_n 0.00631736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1631_n 0.0155187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1632_n 0.0107599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1633_n 0.0301066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_275_481#_c_1772_n 0.00584059f $X=-0.19 $Y=1.655 $X2=2.25
+ $Y2=2.125
cc_274 VPB N_A_275_481#_c_1776_n 0.0062913f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.16
cc_275 VPB N_A_275_481#_c_1777_n 0.00121439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_275_481#_c_1778_n 0.0184258f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_277 VPB N_A_275_481#_c_1779_n 0.0118797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_A_275_481#_c_1780_n 0.0116921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_275_481#_c_1774_n 0.00543208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_Q_c_1898_n 0.0207985f $X=-0.19 $Y=1.655 $X2=2.315 $Y2=0.445
cc_281 VPB Q_N 0.0102592f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.725
cc_282 VPB Q_N 0.0586979f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=0.445
cc_283 N_SCE_M1034_g N_D_M1039_g 0.0396024f $X=0.94 $Y=2.725 $X2=0 $Y2=0
cc_284 N_SCE_c_295_n N_D_M1039_g 0.0150935f $X=2.125 $Y=2.21 $X2=0 $Y2=0
cc_285 N_SCE_M1006_g N_D_c_378_n 0.00572266f $X=2.315 $Y=0.445 $X2=0 $Y2=0
cc_286 N_SCE_c_286_n D 0.00380975f $X=0.68 $Y=0.84 $X2=0 $Y2=0
cc_287 N_SCE_M1006_g D 0.00124039f $X=2.315 $Y=0.445 $X2=0 $Y2=0
cc_288 N_SCE_c_295_n D 0.0515434f $X=2.125 $Y=2.21 $X2=0 $Y2=0
cc_289 N_SCE_c_290_n D 0.0582266f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_290 N_SCE_c_291_n D 0.0063706f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_291 N_SCE_c_298_n D 2.46634e-19 $X=0.94 $Y=2.08 $X2=0 $Y2=0
cc_292 N_SCE_c_299_n D 0.00239721f $X=0.935 $Y=2.105 $X2=0 $Y2=0
cc_293 N_SCE_c_295_n N_D_c_383_n 0.0044058f $X=2.125 $Y=2.21 $X2=0 $Y2=0
cc_294 N_SCE_c_298_n N_D_c_383_n 0.0396024f $X=0.94 $Y=2.08 $X2=0 $Y2=0
cc_295 N_SCE_c_299_n N_D_c_383_n 0.00104852f $X=0.935 $Y=2.105 $X2=0 $Y2=0
cc_296 N_SCE_M1006_g N_D_c_380_n 0.00793805f $X=2.315 $Y=0.445 $X2=0 $Y2=0
cc_297 N_SCE_c_291_n N_D_c_380_n 0.00630029f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_298 N_SCE_c_288_n N_A_34_481#_M1032_g 0.019748f $X=0.755 $Y=0.765 $X2=0 $Y2=0
cc_299 N_SCE_c_295_n N_A_34_481#_c_423_n 7.74269e-19 $X=2.125 $Y=2.21 $X2=0
+ $Y2=0
cc_300 N_SCE_c_290_n N_A_34_481#_c_423_n 4.5648e-19 $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_301 N_SCE_c_291_n N_A_34_481#_c_423_n 0.0225971f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_302 N_SCE_c_295_n N_A_34_481#_M1008_g 0.0115587f $X=2.125 $Y=2.21 $X2=0 $Y2=0
cc_303 N_SCE_c_290_n N_A_34_481#_M1008_g 0.0069447f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_304 N_SCE_c_285_n N_A_34_481#_c_425_n 0.0181643f $X=0.29 $Y=1.915 $X2=0 $Y2=0
cc_305 N_SCE_c_286_n N_A_34_481#_c_425_n 0.0153258f $X=0.68 $Y=0.84 $X2=0 $Y2=0
cc_306 N_SCE_c_295_n N_A_34_481#_c_425_n 0.00268217f $X=2.125 $Y=2.21 $X2=0
+ $Y2=0
cc_307 N_SCE_c_298_n N_A_34_481#_c_425_n 0.0107796f $X=0.94 $Y=2.08 $X2=0 $Y2=0
cc_308 N_SCE_c_299_n N_A_34_481#_c_425_n 0.00140678f $X=0.935 $Y=2.105 $X2=0
+ $Y2=0
cc_309 N_SCE_c_285_n N_A_34_481#_c_427_n 0.00791508f $X=0.29 $Y=1.915 $X2=0
+ $Y2=0
cc_310 N_SCE_c_286_n N_A_34_481#_c_427_n 0.0072063f $X=0.68 $Y=0.84 $X2=0 $Y2=0
cc_311 N_SCE_c_287_n N_A_34_481#_c_427_n 0.00711875f $X=0.365 $Y=0.84 $X2=0
+ $Y2=0
cc_312 N_SCE_c_288_n N_A_34_481#_c_427_n 0.00437996f $X=0.755 $Y=0.765 $X2=0
+ $Y2=0
cc_313 N_SCE_c_285_n N_A_34_481#_c_428_n 0.0190334f $X=0.29 $Y=1.915 $X2=0 $Y2=0
cc_314 N_SCE_M1022_g N_A_34_481#_c_428_n 0.00608969f $X=0.51 $Y=2.725 $X2=0
+ $Y2=0
cc_315 N_SCE_c_298_n N_A_34_481#_c_428_n 0.0201679f $X=0.94 $Y=2.08 $X2=0 $Y2=0
cc_316 N_SCE_c_299_n N_A_34_481#_c_428_n 0.0290517f $X=0.935 $Y=2.105 $X2=0
+ $Y2=0
cc_317 N_SCE_c_286_n N_A_34_481#_c_429_n 0.00631576f $X=0.68 $Y=0.84 $X2=0 $Y2=0
cc_318 N_SCE_c_298_n N_A_34_481#_c_429_n 0.00795051f $X=0.94 $Y=2.08 $X2=0 $Y2=0
cc_319 N_SCE_c_299_n N_A_34_481#_c_429_n 0.0128743f $X=0.935 $Y=2.105 $X2=0
+ $Y2=0
cc_320 N_SCE_c_286_n N_A_34_481#_c_430_n 0.00610353f $X=0.68 $Y=0.84 $X2=0 $Y2=0
cc_321 N_SCE_c_287_n N_A_34_481#_c_430_n 8.25904e-19 $X=0.365 $Y=0.84 $X2=0
+ $Y2=0
cc_322 N_SCE_c_285_n N_A_34_481#_c_431_n 0.0132635f $X=0.29 $Y=1.915 $X2=0 $Y2=0
cc_323 N_SCE_c_286_n N_A_34_481#_c_431_n 2.37e-19 $X=0.68 $Y=0.84 $X2=0 $Y2=0
cc_324 N_SCE_c_295_n N_SCD_M1011_g 0.00573978f $X=2.125 $Y=2.21 $X2=0 $Y2=0
cc_325 N_SCE_c_295_n N_SCD_c_492_n 0.00186378f $X=2.125 $Y=2.21 $X2=0 $Y2=0
cc_326 N_SCE_c_290_n N_SCD_c_492_n 0.00413658f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_327 N_SCE_c_291_n N_SCD_c_492_n 0.0106879f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_328 N_SCE_M1006_g N_SCD_M1036_g 0.0401713f $X=2.315 $Y=0.445 $X2=0 $Y2=0
cc_329 N_SCE_c_290_n N_SCD_M1036_g 0.00192393f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_330 N_SCE_c_291_n N_SCD_M1036_g 0.0412137f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_331 N_SCE_c_295_n SCD 0.00614105f $X=2.125 $Y=2.21 $X2=0 $Y2=0
cc_332 N_SCE_c_290_n SCD 0.0780921f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_333 N_SCE_c_291_n SCD 0.00366337f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_334 N_SCE_c_295_n N_SCD_c_495_n 0.00346186f $X=2.125 $Y=2.21 $X2=0 $Y2=0
cc_335 N_SCE_c_290_n N_SCD_c_495_n 0.00304767f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_336 N_SCE_c_290_n N_SCD_c_496_n 0.00198758f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_337 N_SCE_c_295_n N_CLK_M1009_g 4.73515e-19 $X=2.125 $Y=2.21 $X2=0 $Y2=0
cc_338 N_SCE_M1022_g N_VPWR_c_1609_n 0.0115345f $X=0.51 $Y=2.725 $X2=0 $Y2=0
cc_339 N_SCE_M1034_g N_VPWR_c_1609_n 0.015217f $X=0.94 $Y=2.725 $X2=0 $Y2=0
cc_340 N_SCE_c_298_n N_VPWR_c_1609_n 6.93842e-19 $X=0.94 $Y=2.08 $X2=0 $Y2=0
cc_341 N_SCE_c_299_n N_VPWR_c_1609_n 0.023196f $X=0.935 $Y=2.105 $X2=0 $Y2=0
cc_342 N_SCE_M1022_g N_VPWR_c_1622_n 0.00445056f $X=0.51 $Y=2.725 $X2=0 $Y2=0
cc_343 N_SCE_M1034_g N_VPWR_c_1623_n 0.00445056f $X=0.94 $Y=2.725 $X2=0 $Y2=0
cc_344 N_SCE_M1022_g N_VPWR_c_1608_n 0.00876571f $X=0.51 $Y=2.725 $X2=0 $Y2=0
cc_345 N_SCE_M1034_g N_VPWR_c_1608_n 0.0079903f $X=0.94 $Y=2.725 $X2=0 $Y2=0
cc_346 N_SCE_M1006_g N_A_275_481#_c_1770_n 0.0233343f $X=2.315 $Y=0.445 $X2=0
+ $Y2=0
cc_347 N_SCE_c_290_n N_A_275_481#_c_1770_n 0.00877309f $X=2.29 $Y=1.16 $X2=0
+ $Y2=0
cc_348 N_SCE_c_291_n N_A_275_481#_c_1770_n 0.00353247f $X=2.29 $Y=1.16 $X2=0
+ $Y2=0
cc_349 N_SCE_c_295_n N_A_275_481#_c_1785_n 0.0358543f $X=2.125 $Y=2.21 $X2=0
+ $Y2=0
cc_350 N_SCE_c_295_n N_A_275_481#_c_1772_n 0.0034472f $X=2.125 $Y=2.21 $X2=0
+ $Y2=0
cc_351 N_SCE_c_290_n N_A_275_481#_c_1772_n 0.00264304f $X=2.29 $Y=1.16 $X2=0
+ $Y2=0
cc_352 N_SCE_c_295_n N_A_275_481#_c_1788_n 0.023158f $X=2.125 $Y=2.21 $X2=0
+ $Y2=0
cc_353 N_SCE_c_288_n N_VGND_c_1931_n 0.0104856f $X=0.755 $Y=0.765 $X2=0 $Y2=0
cc_354 N_SCE_M1006_g N_VGND_c_1932_n 0.00143462f $X=2.315 $Y=0.445 $X2=0 $Y2=0
cc_355 N_SCE_c_286_n N_VGND_c_1939_n 8.2951e-19 $X=0.68 $Y=0.84 $X2=0 $Y2=0
cc_356 N_SCE_c_288_n N_VGND_c_1939_n 0.00486043f $X=0.755 $Y=0.765 $X2=0 $Y2=0
cc_357 N_SCE_M1006_g N_VGND_c_1941_n 0.00364515f $X=2.315 $Y=0.445 $X2=0 $Y2=0
cc_358 N_SCE_c_286_n N_VGND_c_1953_n 9.49268e-19 $X=0.68 $Y=0.84 $X2=0 $Y2=0
cc_359 N_SCE_c_288_n N_VGND_c_1953_n 0.0095519f $X=0.755 $Y=0.765 $X2=0 $Y2=0
cc_360 N_SCE_M1006_g N_VGND_c_1953_n 0.00612358f $X=2.315 $Y=0.445 $X2=0 $Y2=0
cc_361 N_D_c_378_n N_A_34_481#_M1032_g 0.0622134f $X=1.545 $Y=0.765 $X2=0 $Y2=0
cc_362 D N_A_34_481#_M1032_g 0.0156011f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_363 D N_A_34_481#_c_423_n 0.0253782f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_364 N_D_c_380_n N_A_34_481#_c_423_n 0.0288434f $X=1.75 $Y=0.93 $X2=0 $Y2=0
cc_365 N_D_M1039_g N_A_34_481#_M1008_g 0.0249992f $X=1.3 $Y=2.725 $X2=0 $Y2=0
cc_366 D N_A_34_481#_M1008_g 0.0149962f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_367 N_D_c_383_n N_A_34_481#_M1008_g 0.0206622f $X=1.39 $Y=1.86 $X2=0 $Y2=0
cc_368 D N_A_34_481#_c_425_n 0.00486457f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_369 D N_A_34_481#_c_426_n 0.0118508f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_370 N_D_c_383_n N_A_34_481#_c_426_n 0.0180994f $X=1.39 $Y=1.86 $X2=0 $Y2=0
cc_371 D N_A_34_481#_c_429_n 0.0277655f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_372 N_D_M1039_g N_VPWR_c_1609_n 0.00269808f $X=1.3 $Y=2.725 $X2=0 $Y2=0
cc_373 N_D_M1039_g N_VPWR_c_1623_n 0.0053602f $X=1.3 $Y=2.725 $X2=0 $Y2=0
cc_374 N_D_M1039_g N_VPWR_c_1608_n 0.0105051f $X=1.3 $Y=2.725 $X2=0 $Y2=0
cc_375 N_D_c_378_n N_A_275_481#_c_1770_n 0.00556873f $X=1.545 $Y=0.765 $X2=0
+ $Y2=0
cc_376 D N_A_275_481#_c_1770_n 0.0250734f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_377 N_D_c_380_n N_A_275_481#_c_1770_n 0.00203442f $X=1.75 $Y=0.93 $X2=0 $Y2=0
cc_378 N_D_M1039_g N_A_275_481#_c_1788_n 0.00790438f $X=1.3 $Y=2.725 $X2=0 $Y2=0
cc_379 N_D_c_378_n N_VGND_c_1931_n 0.0022187f $X=1.545 $Y=0.765 $X2=0 $Y2=0
cc_380 D N_VGND_c_1931_n 0.00214357f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_381 N_D_c_378_n N_VGND_c_1941_n 0.0054833f $X=1.545 $Y=0.765 $X2=0 $Y2=0
cc_382 N_D_c_378_n N_VGND_c_1953_n 0.00671354f $X=1.545 $Y=0.765 $X2=0 $Y2=0
cc_383 D N_VGND_c_1953_n 0.0181181f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_384 N_A_34_481#_M1008_g N_SCD_c_492_n 0.0711824f $X=1.84 $Y=2.725 $X2=0 $Y2=0
cc_385 N_A_34_481#_M1008_g N_SCD_c_496_n 0.00237696f $X=1.84 $Y=2.725 $X2=0
+ $Y2=0
cc_386 N_A_34_481#_c_428_n N_VPWR_c_1609_n 0.0232759f $X=0.295 $Y=2.55 $X2=0
+ $Y2=0
cc_387 N_A_34_481#_c_428_n N_VPWR_c_1622_n 0.0173955f $X=0.295 $Y=2.55 $X2=0
+ $Y2=0
cc_388 N_A_34_481#_M1008_g N_VPWR_c_1623_n 0.00383441f $X=1.84 $Y=2.725 $X2=0
+ $Y2=0
cc_389 N_A_34_481#_M1008_g N_VPWR_c_1608_n 0.0055441f $X=1.84 $Y=2.725 $X2=0
+ $Y2=0
cc_390 N_A_34_481#_c_428_n N_VPWR_c_1608_n 0.00998284f $X=0.295 $Y=2.55 $X2=0
+ $Y2=0
cc_391 N_A_34_481#_M1032_g N_A_275_481#_c_1770_n 8.48142e-19 $X=1.185 $Y=0.445
+ $X2=0 $Y2=0
cc_392 N_A_34_481#_M1008_g N_A_275_481#_c_1785_n 0.00817803f $X=1.84 $Y=2.725
+ $X2=0 $Y2=0
cc_393 N_A_34_481#_M1008_g N_A_275_481#_c_1788_n 0.00772288f $X=1.84 $Y=2.725
+ $X2=0 $Y2=0
cc_394 N_A_34_481#_M1032_g N_VGND_c_1931_n 0.0110793f $X=1.185 $Y=0.445 $X2=0
+ $Y2=0
cc_395 N_A_34_481#_c_425_n N_VGND_c_1931_n 0.00601606f $X=1.11 $Y=1.29 $X2=0
+ $Y2=0
cc_396 N_A_34_481#_c_429_n N_VGND_c_1931_n 0.00321439f $X=0.77 $Y=1.29 $X2=0
+ $Y2=0
cc_397 N_A_34_481#_c_430_n N_VGND_c_1939_n 0.0288984f $X=0.54 $Y=0.445 $X2=0
+ $Y2=0
cc_398 N_A_34_481#_M1032_g N_VGND_c_1941_n 0.00486043f $X=1.185 $Y=0.445 $X2=0
+ $Y2=0
cc_399 N_A_34_481#_M1013_s N_VGND_c_1953_n 0.00269609f $X=0.415 $Y=0.235 $X2=0
+ $Y2=0
cc_400 N_A_34_481#_M1032_g N_VGND_c_1953_n 0.0042918f $X=1.185 $Y=0.445 $X2=0
+ $Y2=0
cc_401 N_A_34_481#_c_430_n N_VGND_c_1953_n 0.0190046f $X=0.54 $Y=0.445 $X2=0
+ $Y2=0
cc_402 N_SCD_M1036_g N_CLK_c_534_n 0.0182245f $X=2.74 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_403 SCD N_CLK_c_534_n 6.04135e-19 $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_404 N_SCD_c_496_n N_CLK_M1009_g 0.0182245f $X=2.74 $Y=2.04 $X2=0 $Y2=0
cc_405 N_SCD_M1036_g N_CLK_M1023_g 0.0425805f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_406 N_SCD_M1011_g N_VPWR_c_1610_n 0.0105165f $X=2.2 $Y=2.725 $X2=0 $Y2=0
cc_407 N_SCD_M1011_g N_VPWR_c_1623_n 0.00391581f $X=2.2 $Y=2.725 $X2=0 $Y2=0
cc_408 N_SCD_M1011_g N_VPWR_c_1608_n 0.00638569f $X=2.2 $Y=2.725 $X2=0 $Y2=0
cc_409 N_SCD_M1036_g N_A_275_481#_c_1770_n 0.00536607f $X=2.74 $Y=0.445 $X2=0
+ $Y2=0
cc_410 N_SCD_M1011_g N_A_275_481#_c_1785_n 0.0136183f $X=2.2 $Y=2.725 $X2=0
+ $Y2=0
cc_411 SCD N_A_275_481#_c_1785_n 0.0103322f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_412 N_SCD_c_495_n N_A_275_481#_c_1785_n 0.00590663f $X=2.475 $Y=2.04 $X2=0
+ $Y2=0
cc_413 N_SCD_c_496_n N_A_275_481#_c_1785_n 0.00421804f $X=2.74 $Y=2.04 $X2=0
+ $Y2=0
cc_414 N_SCD_M1036_g N_A_275_481#_c_1771_n 0.0131345f $X=2.74 $Y=0.445 $X2=0
+ $Y2=0
cc_415 SCD N_A_275_481#_c_1771_n 0.0113634f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_416 N_SCD_M1011_g N_A_275_481#_c_1772_n 0.00422734f $X=2.2 $Y=2.725 $X2=0
+ $Y2=0
cc_417 N_SCD_M1036_g N_A_275_481#_c_1772_n 0.0120281f $X=2.74 $Y=0.445 $X2=0
+ $Y2=0
cc_418 SCD N_A_275_481#_c_1772_n 0.0810801f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_419 N_SCD_M1011_g N_A_275_481#_c_1806_n 0.00368091f $X=2.2 $Y=2.725 $X2=0
+ $Y2=0
cc_420 N_SCD_M1011_g N_A_275_481#_c_1788_n 0.00146911f $X=2.2 $Y=2.725 $X2=0
+ $Y2=0
cc_421 N_SCD_M1036_g N_VGND_c_1932_n 0.00835962f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_422 N_SCD_M1036_g N_VGND_c_1941_n 0.00355956f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_423 N_SCD_M1036_g N_VGND_c_1953_n 0.00424676f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_424 N_CLK_c_534_n N_A_640_481#_c_1125_n 0.0286511f $X=3.125 $Y=1.66 $X2=0
+ $Y2=0
cc_425 CLK N_A_640_481#_c_1125_n 0.00557347f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_426 N_CLK_c_534_n N_A_640_481#_c_1133_n 6.16535e-19 $X=3.125 $Y=1.66 $X2=0
+ $Y2=0
cc_427 N_CLK_c_534_n N_A_640_481#_c_1135_n 0.00224146f $X=3.125 $Y=1.66 $X2=0
+ $Y2=0
cc_428 CLK N_A_640_481#_c_1135_n 0.0399378f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_429 CLK N_A_640_481#_c_1145_n 0.0166676f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_430 N_CLK_M1009_g N_A_640_481#_c_1146_n 0.00407906f $X=3.125 $Y=2.725 $X2=0
+ $Y2=0
cc_431 CLK N_A_640_481#_c_1146_n 0.00888105f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_432 N_CLK_c_534_n N_A_640_481#_c_1136_n 8.27617e-19 $X=3.125 $Y=1.66 $X2=0
+ $Y2=0
cc_433 N_CLK_M1023_g N_A_640_481#_c_1136_n 0.00350824f $X=3.17 $Y=0.445 $X2=0
+ $Y2=0
cc_434 CLK N_A_640_481#_c_1136_n 0.0845367f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_435 N_CLK_M1009_g N_VPWR_c_1610_n 0.00393481f $X=3.125 $Y=2.725 $X2=0 $Y2=0
cc_436 N_CLK_M1009_g N_VPWR_c_1624_n 0.00327695f $X=3.125 $Y=2.725 $X2=0 $Y2=0
cc_437 N_CLK_M1009_g N_VPWR_c_1608_n 0.00667022f $X=3.125 $Y=2.725 $X2=0 $Y2=0
cc_438 N_CLK_M1023_g N_A_275_481#_c_1771_n 0.00530376f $X=3.17 $Y=0.445 $X2=0
+ $Y2=0
cc_439 N_CLK_c_534_n N_A_275_481#_c_1772_n 0.00342111f $X=3.125 $Y=1.66 $X2=0
+ $Y2=0
cc_440 N_CLK_M1009_g N_A_275_481#_c_1772_n 0.0270915f $X=3.125 $Y=2.725 $X2=0
+ $Y2=0
cc_441 N_CLK_M1023_g N_A_275_481#_c_1772_n 0.00651567f $X=3.17 $Y=0.445 $X2=0
+ $Y2=0
cc_442 CLK N_A_275_481#_c_1772_n 0.0724411f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_443 N_CLK_M1009_g N_A_275_481#_c_1806_n 0.00843126f $X=3.125 $Y=2.725 $X2=0
+ $Y2=0
cc_444 N_CLK_M1009_g N_A_275_481#_c_1776_n 0.0120447f $X=3.125 $Y=2.725 $X2=0
+ $Y2=0
cc_445 N_CLK_M1009_g N_A_275_481#_c_1777_n 0.00352175f $X=3.125 $Y=2.725 $X2=0
+ $Y2=0
cc_446 N_CLK_M1009_g N_A_275_481#_c_1816_n 0.00592956f $X=3.125 $Y=2.725 $X2=0
+ $Y2=0
cc_447 N_CLK_M1009_g N_A_275_481#_c_1779_n 0.00315613f $X=3.125 $Y=2.725 $X2=0
+ $Y2=0
cc_448 N_CLK_M1023_g N_VGND_c_1932_n 0.011491f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_449 N_CLK_M1023_g N_VGND_c_1943_n 0.00486043f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_450 N_CLK_c_534_n N_VGND_c_1953_n 7.83929e-19 $X=3.125 $Y=1.66 $X2=0 $Y2=0
cc_451 N_CLK_M1023_g N_VGND_c_1953_n 0.00975473f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_452 CLK N_VGND_c_1953_n 0.00142635f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_453 N_A_901_441#_M1018_g N_A_1274_401#_M1031_g 0.00102402f $X=5.655 $Y=2.525
+ $X2=0 $Y2=0
cc_454 N_A_901_441#_M1025_g N_A_1274_401#_M1015_g 0.0778942f $X=6.15 $Y=0.805
+ $X2=0 $Y2=0
cc_455 N_A_901_441#_c_577_n N_A_1274_401#_M1015_g 0.00353751f $X=5.655 $Y=1.71
+ $X2=0 $Y2=0
cc_456 N_A_901_441#_c_582_n N_A_1274_401#_M1015_g 0.0122324f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_457 N_A_901_441#_c_587_n N_A_1274_401#_M1015_g 0.00118604f $X=6.095 $Y=1.46
+ $X2=0 $Y2=0
cc_458 N_A_901_441#_c_582_n N_A_1274_401#_c_745_n 0.0237576f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_459 N_A_901_441#_c_597_n N_A_1274_401#_c_746_n 0.0247501f $X=8.955 $Y=1.865
+ $X2=0 $Y2=0
cc_460 N_A_901_441#_c_607_p N_A_1274_401#_c_746_n 0.00422847f $X=7.985 $Y=1.865
+ $X2=0 $Y2=0
cc_461 N_A_901_441#_c_582_n N_A_1274_401#_c_747_n 0.00724449f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_462 N_A_901_441#_c_575_n N_A_1274_401#_c_740_n 0.0148814f $X=9.525 $Y=1.35
+ $X2=0 $Y2=0
cc_463 N_A_901_441#_c_580_n N_A_1274_401#_c_740_n 0.00945986f $X=9.975 $Y=1.515
+ $X2=0 $Y2=0
cc_464 N_A_901_441#_c_597_n N_A_1274_401#_c_740_n 0.00603101f $X=8.955 $Y=1.865
+ $X2=0 $Y2=0
cc_465 N_A_901_441#_c_612_p N_A_1274_401#_c_740_n 0.0131874f $X=9.125 $Y=1.515
+ $X2=0 $Y2=0
cc_466 N_A_901_441#_c_585_n N_A_1274_401#_c_740_n 0.0476954f $X=9.625 $Y=1.515
+ $X2=0 $Y2=0
cc_467 N_A_901_441#_M1012_g N_A_1274_401#_c_766_n 0.00116943f $X=10.05 $Y=2.65
+ $X2=0 $Y2=0
cc_468 N_A_901_441#_M1012_g N_A_1274_401#_c_748_n 0.00814299f $X=10.05 $Y=2.65
+ $X2=0 $Y2=0
cc_469 N_A_901_441#_c_579_n N_A_1274_401#_c_748_n 0.010303f $X=9.6 $Y=1.515
+ $X2=0 $Y2=0
cc_470 N_A_901_441#_c_585_n N_A_1274_401#_c_748_n 0.0213831f $X=9.625 $Y=1.515
+ $X2=0 $Y2=0
cc_471 N_A_901_441#_c_597_n N_A_1274_401#_c_749_n 0.0126727f $X=8.955 $Y=1.865
+ $X2=0 $Y2=0
cc_472 N_A_901_441#_c_585_n N_A_1274_401#_c_749_n 0.0136506f $X=9.625 $Y=1.515
+ $X2=0 $Y2=0
cc_473 N_A_901_441#_c_575_n N_A_1274_401#_c_742_n 0.00276977f $X=9.525 $Y=1.35
+ $X2=0 $Y2=0
cc_474 N_A_901_441#_M1012_g N_A_1274_401#_c_742_n 0.00288395f $X=10.05 $Y=2.65
+ $X2=0 $Y2=0
cc_475 N_A_901_441#_c_580_n N_A_1274_401#_c_742_n 0.0157384f $X=9.975 $Y=1.515
+ $X2=0 $Y2=0
cc_476 N_A_901_441#_c_585_n N_A_1274_401#_c_742_n 0.014321f $X=9.625 $Y=1.515
+ $X2=0 $Y2=0
cc_477 N_A_901_441#_c_577_n N_A_1274_401#_c_751_n 0.00102402f $X=5.655 $Y=1.71
+ $X2=0 $Y2=0
cc_478 N_A_901_441#_c_582_n N_A_1274_401#_c_751_n 0.006283f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_479 N_A_901_441#_c_582_n N_A_1146_463#_M1004_g 0.0142932f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_480 N_A_901_441#_c_583_n N_A_1146_463#_M1004_g 0.00492812f $X=7.9 $Y=1.78
+ $X2=0 $Y2=0
cc_481 N_A_901_441#_c_607_p N_A_1146_463#_M1004_g 2.73505e-19 $X=7.985 $Y=1.865
+ $X2=0 $Y2=0
cc_482 N_A_901_441#_c_582_n N_A_1146_463#_c_868_n 7.52953e-19 $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_483 N_A_901_441#_c_579_n N_A_1146_463#_c_870_n 0.0389376f $X=9.6 $Y=1.515
+ $X2=0 $Y2=0
cc_484 N_A_901_441#_c_584_n N_A_1146_463#_c_870_n 0.00415539f $X=9.04 $Y=1.78
+ $X2=0 $Y2=0
cc_485 N_A_901_441#_c_612_p N_A_1146_463#_c_870_n 0.00928735f $X=9.125 $Y=1.515
+ $X2=0 $Y2=0
cc_486 N_A_901_441#_c_585_n N_A_1146_463#_c_870_n 0.00501671f $X=9.625 $Y=1.515
+ $X2=0 $Y2=0
cc_487 N_A_901_441#_c_597_n N_A_1146_463#_M1019_g 0.0109798f $X=8.955 $Y=1.865
+ $X2=0 $Y2=0
cc_488 N_A_901_441#_c_584_n N_A_1146_463#_M1019_g 0.00626049f $X=9.04 $Y=1.78
+ $X2=0 $Y2=0
cc_489 N_A_901_441#_c_575_n N_A_1146_463#_c_871_n 0.0329718f $X=9.525 $Y=1.35
+ $X2=0 $Y2=0
cc_490 N_A_901_441#_c_582_n N_A_1146_463#_c_872_n 0.0113882f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_491 N_A_901_441#_c_597_n N_A_1146_463#_c_873_n 0.0127332f $X=8.955 $Y=1.865
+ $X2=0 $Y2=0
cc_492 N_A_901_441#_M1018_g N_A_1146_463#_c_887_n 0.00324927f $X=5.655 $Y=2.525
+ $X2=0 $Y2=0
cc_493 N_A_901_441#_M1025_g N_A_1146_463#_c_904_n 0.0068621f $X=6.15 $Y=0.805
+ $X2=0 $Y2=0
cc_494 N_A_901_441#_M1025_g N_A_1146_463#_c_874_n 0.0106216f $X=6.15 $Y=0.805
+ $X2=0 $Y2=0
cc_495 N_A_901_441#_c_582_n N_A_1146_463#_c_874_n 0.0615864f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_496 N_A_901_441#_c_587_n N_A_1146_463#_c_874_n 0.0089045f $X=6.095 $Y=1.46
+ $X2=0 $Y2=0
cc_497 N_A_901_441#_M1025_g N_A_1146_463#_c_875_n 0.00346656f $X=6.15 $Y=0.805
+ $X2=0 $Y2=0
cc_498 N_A_901_441#_c_578_n N_A_1146_463#_c_875_n 0.00582336f $X=6.075 $Y=1.54
+ $X2=0 $Y2=0
cc_499 N_A_901_441#_c_587_n N_A_1146_463#_c_875_n 0.0110368f $X=6.095 $Y=1.46
+ $X2=0 $Y2=0
cc_500 N_A_901_441#_c_582_n N_A_1146_463#_c_878_n 0.0544245f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_501 N_A_901_441#_c_597_n N_A_1146_463#_c_878_n 0.00521101f $X=8.955 $Y=1.865
+ $X2=0 $Y2=0
cc_502 N_A_901_441#_c_582_n N_A_1146_463#_c_879_n 0.00344531f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_503 N_A_901_441#_c_582_n N_A_1146_463#_c_880_n 0.0105869f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_504 N_A_901_441#_c_583_n N_A_1146_463#_c_880_n 0.00489445f $X=7.9 $Y=1.78
+ $X2=0 $Y2=0
cc_505 N_A_901_441#_c_597_n N_A_1146_463#_c_880_n 0.012751f $X=8.955 $Y=1.865
+ $X2=0 $Y2=0
cc_506 N_A_901_441#_c_597_n N_A_1146_463#_c_881_n 0.0303035f $X=8.955 $Y=1.865
+ $X2=0 $Y2=0
cc_507 N_A_901_441#_c_612_p N_A_1146_463#_c_881_n 0.0150684f $X=9.125 $Y=1.515
+ $X2=0 $Y2=0
cc_508 N_A_901_441#_M1025_g N_A_1146_463#_c_882_n 0.00363706f $X=6.15 $Y=0.805
+ $X2=0 $Y2=0
cc_509 N_A_901_441#_c_577_n N_A_1146_463#_c_882_n 0.0158121f $X=5.655 $Y=1.71
+ $X2=0 $Y2=0
cc_510 N_A_901_441#_c_578_n N_A_1146_463#_c_882_n 0.00845696f $X=6.075 $Y=1.54
+ $X2=0 $Y2=0
cc_511 N_A_901_441#_c_587_n N_A_1146_463#_c_882_n 0.023122f $X=6.095 $Y=1.46
+ $X2=0 $Y2=0
cc_512 N_A_901_441#_M1018_g N_A_1146_463#_c_889_n 0.00569062f $X=5.655 $Y=2.525
+ $X2=0 $Y2=0
cc_513 N_A_901_441#_c_577_n N_A_1146_463#_c_889_n 0.00653804f $X=5.655 $Y=1.71
+ $X2=0 $Y2=0
cc_514 N_A_901_441#_c_578_n N_A_1146_463#_c_889_n 0.00556555f $X=6.075 $Y=1.54
+ $X2=0 $Y2=0
cc_515 N_A_901_441#_c_587_n N_A_1146_463#_c_889_n 0.0055184f $X=6.095 $Y=1.46
+ $X2=0 $Y2=0
cc_516 N_A_901_441#_c_582_n N_A_1146_463#_c_927_n 0.0147533f $X=7.815 $Y=1.46
+ $X2=0 $Y2=0
cc_517 N_A_901_441#_c_582_n N_SET_B_c_1012_n 0.00608034f $X=7.815 $Y=1.46
+ $X2=-0.19 $Y2=-0.245
cc_518 N_A_901_441#_c_597_n N_SET_B_c_1014_n 0.0116734f $X=8.955 $Y=1.865 $X2=0
+ $Y2=0
cc_519 N_A_901_441#_c_607_p N_SET_B_c_1014_n 0.0103383f $X=7.985 $Y=1.865 $X2=0
+ $Y2=0
cc_520 N_A_901_441#_c_582_n N_SET_B_M1041_g 0.00373004f $X=7.815 $Y=1.46 $X2=0
+ $Y2=0
cc_521 N_A_901_441#_c_583_n N_SET_B_M1041_g 0.00761636f $X=7.9 $Y=1.78 $X2=0
+ $Y2=0
cc_522 N_A_901_441#_c_597_n N_SET_B_M1041_g 0.00352644f $X=8.955 $Y=1.865 $X2=0
+ $Y2=0
cc_523 N_A_901_441#_M1012_g N_SET_B_c_1017_n 0.00506374f $X=10.05 $Y=2.65 $X2=0
+ $Y2=0
cc_524 N_A_901_441#_c_582_n N_SET_B_c_1017_n 0.0057605f $X=7.815 $Y=1.46 $X2=0
+ $Y2=0
cc_525 N_A_901_441#_c_597_n N_SET_B_c_1017_n 0.0367639f $X=8.955 $Y=1.865 $X2=0
+ $Y2=0
cc_526 N_A_901_441#_c_607_p N_SET_B_c_1017_n 0.00525051f $X=7.985 $Y=1.865 $X2=0
+ $Y2=0
cc_527 N_A_901_441#_c_585_n N_SET_B_c_1017_n 0.00830424f $X=9.625 $Y=1.515 $X2=0
+ $Y2=0
cc_528 N_A_901_441#_c_582_n N_SET_B_c_1018_n 0.00328768f $X=7.815 $Y=1.46 $X2=0
+ $Y2=0
cc_529 N_A_901_441#_c_607_p N_SET_B_c_1018_n 2.02271e-19 $X=7.985 $Y=1.865 $X2=0
+ $Y2=0
cc_530 N_A_901_441#_c_582_n N_SET_B_c_1019_n 0.0155058f $X=7.815 $Y=1.46 $X2=0
+ $Y2=0
cc_531 N_A_901_441#_c_607_p N_SET_B_c_1019_n 0.0124651f $X=7.985 $Y=1.865 $X2=0
+ $Y2=0
cc_532 N_A_901_441#_c_586_n N_A_640_481#_c_1124_n 0.00753443f $X=5.01 $Y=1.54
+ $X2=0 $Y2=0
cc_533 N_A_901_441#_c_595_n N_A_640_481#_M1017_g 0.0204638f $X=4.645 $Y=2.35
+ $X2=0 $Y2=0
cc_534 N_A_901_441#_c_586_n N_A_640_481#_M1017_g 0.00352508f $X=5.01 $Y=1.54
+ $X2=0 $Y2=0
cc_535 N_A_901_441#_M1018_g N_A_640_481#_c_1139_n 0.0104164f $X=5.655 $Y=2.525
+ $X2=0 $Y2=0
cc_536 N_A_901_441#_c_581_n N_A_640_481#_M1026_g 0.00963415f $X=4.84 $Y=0.565
+ $X2=0 $Y2=0
cc_537 N_A_901_441#_c_581_n N_A_640_481#_c_1128_n 0.00491654f $X=4.84 $Y=0.565
+ $X2=0 $Y2=0
cc_538 N_A_901_441#_M1025_g N_A_640_481#_M1024_g 0.0135865f $X=6.15 $Y=0.805
+ $X2=0 $Y2=0
cc_539 N_A_901_441#_c_577_n N_A_640_481#_M1024_g 0.00872692f $X=5.655 $Y=1.71
+ $X2=0 $Y2=0
cc_540 N_A_901_441#_c_581_n N_A_640_481#_M1024_g 0.00462114f $X=4.84 $Y=0.565
+ $X2=0 $Y2=0
cc_541 N_A_901_441#_M1025_g N_A_640_481#_c_1131_n 0.0103162f $X=6.15 $Y=0.805
+ $X2=0 $Y2=0
cc_542 N_A_901_441#_c_575_n N_A_640_481#_c_1131_n 0.0103123f $X=9.525 $Y=1.35
+ $X2=0 $Y2=0
cc_543 N_A_901_441#_M1018_g N_A_640_481#_M1000_g 0.0128352f $X=5.655 $Y=2.525
+ $X2=0 $Y2=0
cc_544 N_A_901_441#_c_578_n N_A_640_481#_M1000_g 0.00338827f $X=6.075 $Y=1.54
+ $X2=0 $Y2=0
cc_545 N_A_901_441#_c_587_n N_A_640_481#_M1000_g 8.69449e-19 $X=6.095 $Y=1.46
+ $X2=0 $Y2=0
cc_546 N_A_901_441#_M1012_g N_A_640_481#_M1040_g 0.0187007f $X=10.05 $Y=2.65
+ $X2=0 $Y2=0
cc_547 N_A_901_441#_c_579_n N_A_640_481#_M1040_g 0.00988962f $X=9.6 $Y=1.515
+ $X2=0 $Y2=0
cc_548 N_A_901_441#_c_575_n N_A_640_481#_M1030_g 0.0170607f $X=9.525 $Y=1.35
+ $X2=0 $Y2=0
cc_549 N_A_901_441#_c_580_n N_A_640_481#_M1030_g 0.00492181f $X=9.975 $Y=1.515
+ $X2=0 $Y2=0
cc_550 N_A_901_441#_c_576_n N_A_640_481#_c_1133_n 0.0222029f $X=5.58 $Y=1.71
+ $X2=0 $Y2=0
cc_551 N_A_901_441#_c_586_n N_A_640_481#_c_1133_n 0.00583185f $X=5.01 $Y=1.54
+ $X2=0 $Y2=0
cc_552 N_A_901_441#_c_595_n N_A_640_481#_c_1145_n 0.0100478f $X=4.645 $Y=2.35
+ $X2=0 $Y2=0
cc_553 N_A_901_441#_c_581_n N_A_640_481#_c_1136_n 0.0189731f $X=4.84 $Y=0.565
+ $X2=0 $Y2=0
cc_554 N_A_901_441#_c_586_n N_A_640_481#_c_1136_n 0.0387019f $X=5.01 $Y=1.54
+ $X2=0 $Y2=0
cc_555 N_A_901_441#_c_581_n N_A_640_481#_c_1137_n 0.00349615f $X=4.84 $Y=0.565
+ $X2=0 $Y2=0
cc_556 N_A_901_441#_c_580_n N_A_2067_92#_M1035_g 0.00618968f $X=9.975 $Y=1.515
+ $X2=0 $Y2=0
cc_557 N_A_901_441#_M1012_g N_A_2067_92#_M1001_g 0.0458806f $X=10.05 $Y=2.65
+ $X2=0 $Y2=0
cc_558 N_A_901_441#_c_580_n N_A_2067_92#_c_1261_n 0.0458806f $X=9.975 $Y=1.515
+ $X2=0 $Y2=0
cc_559 N_A_901_441#_c_575_n N_A_1920_119#_c_1376_n 0.00526473f $X=9.525 $Y=1.35
+ $X2=0 $Y2=0
cc_560 N_A_901_441#_c_580_n N_A_1920_119#_c_1376_n 4.78075e-19 $X=9.975 $Y=1.515
+ $X2=0 $Y2=0
cc_561 N_A_901_441#_M1012_g N_A_1920_119#_c_1347_n 0.00270572f $X=10.05 $Y=2.65
+ $X2=0 $Y2=0
cc_562 N_A_901_441#_c_580_n N_A_1920_119#_c_1347_n 0.00166958f $X=9.975 $Y=1.515
+ $X2=0 $Y2=0
cc_563 N_A_901_441#_M1012_g N_A_1920_119#_c_1366_n 0.0239397f $X=10.05 $Y=2.65
+ $X2=0 $Y2=0
cc_564 N_A_901_441#_c_580_n N_A_1920_119#_c_1366_n 6.32705e-19 $X=9.975 $Y=1.515
+ $X2=0 $Y2=0
cc_565 N_A_901_441#_c_597_n N_VPWR_M1010_d 0.00264755f $X=8.955 $Y=1.865 $X2=0
+ $Y2=0
cc_566 N_A_901_441#_M1012_g N_VPWR_c_1626_n 0.00372033f $X=10.05 $Y=2.65 $X2=0
+ $Y2=0
cc_567 N_A_901_441#_M1018_g N_VPWR_c_1608_n 9.39239e-19 $X=5.655 $Y=2.525 $X2=0
+ $Y2=0
cc_568 N_A_901_441#_M1012_g N_VPWR_c_1608_n 0.00514438f $X=10.05 $Y=2.65 $X2=0
+ $Y2=0
cc_569 N_A_901_441#_M1012_g N_VPWR_c_1633_n 7.86949e-19 $X=10.05 $Y=2.65 $X2=0
+ $Y2=0
cc_570 N_A_901_441#_M1017_d N_A_275_481#_c_1778_n 0.00567354f $X=4.505 $Y=2.205
+ $X2=0 $Y2=0
cc_571 N_A_901_441#_c_576_n N_A_275_481#_c_1778_n 0.00543855f $X=5.58 $Y=1.71
+ $X2=0 $Y2=0
cc_572 N_A_901_441#_c_595_n N_A_275_481#_c_1778_n 0.0450089f $X=4.645 $Y=2.35
+ $X2=0 $Y2=0
cc_573 N_A_901_441#_M1025_g N_A_275_481#_c_1773_n 2.02886e-19 $X=6.15 $Y=0.805
+ $X2=0 $Y2=0
cc_574 N_A_901_441#_c_576_n N_A_275_481#_c_1773_n 0.0054225f $X=5.58 $Y=1.71
+ $X2=0 $Y2=0
cc_575 N_A_901_441#_c_581_n N_A_275_481#_c_1773_n 0.0284489f $X=4.84 $Y=0.565
+ $X2=0 $Y2=0
cc_576 N_A_901_441#_M1018_g N_A_275_481#_c_1780_n 0.00247583f $X=5.655 $Y=2.525
+ $X2=0 $Y2=0
cc_577 N_A_901_441#_c_576_n N_A_275_481#_c_1780_n 0.00367562f $X=5.58 $Y=1.71
+ $X2=0 $Y2=0
cc_578 N_A_901_441#_c_595_n N_A_275_481#_c_1780_n 0.0417343f $X=4.645 $Y=2.35
+ $X2=0 $Y2=0
cc_579 N_A_901_441#_M1018_g N_A_275_481#_c_1774_n 0.00626074f $X=5.655 $Y=2.525
+ $X2=0 $Y2=0
cc_580 N_A_901_441#_M1025_g N_A_275_481#_c_1774_n 9.0111e-19 $X=6.15 $Y=0.805
+ $X2=0 $Y2=0
cc_581 N_A_901_441#_c_576_n N_A_275_481#_c_1774_n 0.0385495f $X=5.58 $Y=1.71
+ $X2=0 $Y2=0
cc_582 N_A_901_441#_c_581_n N_A_275_481#_c_1774_n 0.0194208f $X=4.84 $Y=0.565
+ $X2=0 $Y2=0
cc_583 N_A_901_441#_c_586_n N_A_275_481#_c_1774_n 0.0417343f $X=5.01 $Y=1.54
+ $X2=0 $Y2=0
cc_584 N_A_901_441#_c_586_n N_VGND_c_1933_n 0.00116267f $X=5.01 $Y=1.54 $X2=0
+ $Y2=0
cc_585 N_A_901_441#_M1025_g N_VGND_c_1934_n 0.00146293f $X=6.15 $Y=0.805 $X2=0
+ $Y2=0
cc_586 N_A_901_441#_c_581_n N_VGND_c_1945_n 0.00991649f $X=4.84 $Y=0.565 $X2=0
+ $Y2=0
cc_587 N_A_901_441#_M1025_g N_VGND_c_1953_n 9.39239e-19 $X=6.15 $Y=0.805 $X2=0
+ $Y2=0
cc_588 N_A_901_441#_c_575_n N_VGND_c_1953_n 9.39239e-19 $X=9.525 $Y=1.35 $X2=0
+ $Y2=0
cc_589 N_A_901_441#_c_581_n N_VGND_c_1953_n 0.00947276f $X=4.84 $Y=0.565 $X2=0
+ $Y2=0
cc_590 N_A_1274_401#_M1031_g N_A_1146_463#_M1004_g 0.00933972f $X=6.445 $Y=2.525
+ $X2=0 $Y2=0
cc_591 N_A_1274_401#_M1015_g N_A_1146_463#_M1004_g 0.0168497f $X=6.51 $Y=0.805
+ $X2=0 $Y2=0
cc_592 N_A_1274_401#_c_747_n N_A_1146_463#_M1004_g 0.024848f $X=7.48 $Y=2.385
+ $X2=0 $Y2=0
cc_593 N_A_1274_401#_c_751_n N_A_1146_463#_M1004_g 0.0184106f $X=6.51 $Y=1.99
+ $X2=0 $Y2=0
cc_594 N_A_1274_401#_c_738_n N_A_1146_463#_c_868_n 0.0012118f $X=8.515 $Y=0.745
+ $X2=0 $Y2=0
cc_595 N_A_1274_401#_c_738_n N_A_1146_463#_c_869_n 0.00940549f $X=8.515 $Y=0.745
+ $X2=0 $Y2=0
cc_596 N_A_1274_401#_c_746_n N_A_1146_463#_M1019_g 0.0132203f $X=9.305 $Y=2.385
+ $X2=0 $Y2=0
cc_597 N_A_1274_401#_c_766_n N_A_1146_463#_M1019_g 0.00641714f $X=9.39 $Y=2.3
+ $X2=0 $Y2=0
cc_598 N_A_1274_401#_c_749_n N_A_1146_463#_M1019_g 0.00103442f $X=9.475 $Y=1.865
+ $X2=0 $Y2=0
cc_599 N_A_1274_401#_c_739_n N_A_1146_463#_c_871_n 0.00420606f $X=8.6 $Y=1.08
+ $X2=0 $Y2=0
cc_600 N_A_1274_401#_c_740_n N_A_1146_463#_c_871_n 0.0161952f $X=9.96 $Y=1.165
+ $X2=0 $Y2=0
cc_601 N_A_1274_401#_c_738_n N_A_1146_463#_c_873_n 0.00126606f $X=8.515 $Y=0.745
+ $X2=0 $Y2=0
cc_602 N_A_1274_401#_c_740_n N_A_1146_463#_c_873_n 0.0112383f $X=9.96 $Y=1.165
+ $X2=0 $Y2=0
cc_603 N_A_1274_401#_c_741_n N_A_1146_463#_c_873_n 0.00429044f $X=8.685 $Y=1.165
+ $X2=0 $Y2=0
cc_604 N_A_1274_401#_M1031_g N_A_1146_463#_c_887_n 0.00269184f $X=6.445 $Y=2.525
+ $X2=0 $Y2=0
cc_605 N_A_1274_401#_M1015_g N_A_1146_463#_c_904_n 0.001439f $X=6.51 $Y=0.805
+ $X2=0 $Y2=0
cc_606 N_A_1274_401#_M1015_g N_A_1146_463#_c_874_n 0.0145926f $X=6.51 $Y=0.805
+ $X2=0 $Y2=0
cc_607 N_A_1274_401#_M1015_g N_A_1146_463#_c_876_n 7.64345e-19 $X=6.51 $Y=0.805
+ $X2=0 $Y2=0
cc_608 N_A_1274_401#_c_738_n N_A_1146_463#_c_876_n 0.0177154f $X=8.515 $Y=0.745
+ $X2=0 $Y2=0
cc_609 N_A_1274_401#_M1015_g N_A_1146_463#_c_877_n 0.017168f $X=6.51 $Y=0.805
+ $X2=0 $Y2=0
cc_610 N_A_1274_401#_c_738_n N_A_1146_463#_c_877_n 0.00214633f $X=8.515 $Y=0.745
+ $X2=0 $Y2=0
cc_611 N_A_1274_401#_c_738_n N_A_1146_463#_c_878_n 0.0600575f $X=8.515 $Y=0.745
+ $X2=0 $Y2=0
cc_612 N_A_1274_401#_c_739_n N_A_1146_463#_c_878_n 0.00442407f $X=8.6 $Y=1.08
+ $X2=0 $Y2=0
cc_613 N_A_1274_401#_c_741_n N_A_1146_463#_c_878_n 0.0112429f $X=8.685 $Y=1.165
+ $X2=0 $Y2=0
cc_614 N_A_1274_401#_c_741_n N_A_1146_463#_c_879_n 0.003613f $X=8.685 $Y=1.165
+ $X2=0 $Y2=0
cc_615 N_A_1274_401#_c_738_n N_A_1146_463#_c_881_n 0.00547362f $X=8.515 $Y=0.745
+ $X2=0 $Y2=0
cc_616 N_A_1274_401#_c_740_n N_A_1146_463#_c_881_n 0.00645161f $X=9.96 $Y=1.165
+ $X2=0 $Y2=0
cc_617 N_A_1274_401#_c_741_n N_A_1146_463#_c_881_n 0.0136959f $X=8.685 $Y=1.165
+ $X2=0 $Y2=0
cc_618 N_A_1274_401#_M1015_g N_A_1146_463#_c_882_n 0.00181757f $X=6.51 $Y=0.805
+ $X2=0 $Y2=0
cc_619 N_A_1274_401#_c_745_n N_A_1146_463#_c_889_n 0.0120811f $X=7.005 $Y=2.047
+ $X2=0 $Y2=0
cc_620 N_A_1274_401#_c_751_n N_A_1146_463#_c_889_n 0.0023594f $X=6.51 $Y=1.99
+ $X2=0 $Y2=0
cc_621 N_A_1274_401#_c_747_n N_SET_B_c_1012_n 7.55298e-19 $X=7.48 $Y=2.385
+ $X2=-0.19 $Y2=-0.245
cc_622 N_A_1274_401#_c_746_n N_SET_B_M1010_g 0.00893946f $X=9.305 $Y=2.385 $X2=0
+ $Y2=0
cc_623 N_A_1274_401#_c_747_n N_SET_B_M1010_g 0.0107839f $X=7.48 $Y=2.385 $X2=0
+ $Y2=0
cc_624 N_A_1274_401#_c_746_n N_SET_B_c_1014_n 0.0172817f $X=9.305 $Y=2.385 $X2=0
+ $Y2=0
cc_625 N_A_1274_401#_c_738_n N_SET_B_M1041_g 0.0142584f $X=8.515 $Y=0.745 $X2=0
+ $Y2=0
cc_626 N_A_1274_401#_c_739_n N_SET_B_M1041_g 0.00545837f $X=8.6 $Y=1.08 $X2=0
+ $Y2=0
cc_627 N_A_1274_401#_c_741_n N_SET_B_M1041_g 0.00106951f $X=8.685 $Y=1.165 $X2=0
+ $Y2=0
cc_628 N_A_1274_401#_c_746_n N_SET_B_c_1017_n 0.0485176f $X=9.305 $Y=2.385 $X2=0
+ $Y2=0
cc_629 N_A_1274_401#_c_766_n N_SET_B_c_1017_n 0.0210576f $X=9.39 $Y=2.3 $X2=0
+ $Y2=0
cc_630 N_A_1274_401#_c_748_n N_SET_B_c_1017_n 0.0222502f $X=9.96 $Y=1.865 $X2=0
+ $Y2=0
cc_631 N_A_1274_401#_c_746_n N_SET_B_c_1018_n 0.00249512f $X=9.305 $Y=2.385
+ $X2=0 $Y2=0
cc_632 N_A_1274_401#_c_747_n N_SET_B_c_1018_n 0.0146797f $X=7.48 $Y=2.385 $X2=0
+ $Y2=0
cc_633 N_A_1274_401#_c_746_n N_SET_B_c_1019_n 0.0104763f $X=9.305 $Y=2.385 $X2=0
+ $Y2=0
cc_634 N_A_1274_401#_c_747_n N_SET_B_c_1019_n 0.0253592f $X=7.48 $Y=2.385 $X2=0
+ $Y2=0
cc_635 N_A_1274_401#_M1015_g N_A_640_481#_c_1131_n 0.0103107f $X=6.51 $Y=0.805
+ $X2=0 $Y2=0
cc_636 N_A_1274_401#_c_738_n N_A_640_481#_c_1131_n 0.0173134f $X=8.515 $Y=0.745
+ $X2=0 $Y2=0
cc_637 N_A_1274_401#_M1031_g N_A_640_481#_M1000_g 0.0401842f $X=6.445 $Y=2.525
+ $X2=0 $Y2=0
cc_638 N_A_1274_401#_M1031_g N_A_640_481#_c_1142_n 0.0103562f $X=6.445 $Y=2.525
+ $X2=0 $Y2=0
cc_639 N_A_1274_401#_c_746_n N_A_640_481#_c_1142_n 0.00998269f $X=9.305 $Y=2.385
+ $X2=0 $Y2=0
cc_640 N_A_1274_401#_c_747_n N_A_640_481#_c_1142_n 0.00506137f $X=7.48 $Y=2.385
+ $X2=0 $Y2=0
cc_641 N_A_1274_401#_c_746_n N_A_640_481#_M1040_g 0.00489752f $X=9.305 $Y=2.385
+ $X2=0 $Y2=0
cc_642 N_A_1274_401#_c_766_n N_A_640_481#_M1040_g 0.00852829f $X=9.39 $Y=2.3
+ $X2=0 $Y2=0
cc_643 N_A_1274_401#_c_748_n N_A_640_481#_M1040_g 0.00389161f $X=9.96 $Y=1.865
+ $X2=0 $Y2=0
cc_644 N_A_1274_401#_c_749_n N_A_640_481#_M1040_g 7.98072e-19 $X=9.475 $Y=1.865
+ $X2=0 $Y2=0
cc_645 N_A_1274_401#_c_740_n N_A_640_481#_M1030_g 0.00619426f $X=9.96 $Y=1.165
+ $X2=0 $Y2=0
cc_646 N_A_1274_401#_c_740_n N_A_2067_92#_M1035_g 0.00103892f $X=9.96 $Y=1.165
+ $X2=0 $Y2=0
cc_647 N_A_1274_401#_c_742_n N_A_2067_92#_M1035_g 0.00192352f $X=10.045 $Y=1.78
+ $X2=0 $Y2=0
cc_648 N_A_1274_401#_c_748_n N_A_2067_92#_c_1261_n 6.19699e-19 $X=9.96 $Y=1.865
+ $X2=0 $Y2=0
cc_649 N_A_1274_401#_c_740_n N_A_1920_119#_M1038_d 0.00229396f $X=9.96 $Y=1.165
+ $X2=-0.19 $Y2=-0.245
cc_650 N_A_1274_401#_c_740_n N_A_1920_119#_c_1376_n 0.0357075f $X=9.96 $Y=1.165
+ $X2=0 $Y2=0
cc_651 N_A_1274_401#_c_740_n N_A_1920_119#_c_1347_n 0.013784f $X=9.96 $Y=1.165
+ $X2=0 $Y2=0
cc_652 N_A_1274_401#_c_748_n N_A_1920_119#_c_1347_n 0.0136857f $X=9.96 $Y=1.865
+ $X2=0 $Y2=0
cc_653 N_A_1274_401#_c_742_n N_A_1920_119#_c_1347_n 0.0382489f $X=10.045 $Y=1.78
+ $X2=0 $Y2=0
cc_654 N_A_1274_401#_c_748_n N_A_1920_119#_c_1366_n 0.0312059f $X=9.96 $Y=1.865
+ $X2=0 $Y2=0
cc_655 N_A_1274_401#_c_746_n N_VPWR_M1010_d 0.0224217f $X=9.305 $Y=2.385 $X2=0
+ $Y2=0
cc_656 N_A_1274_401#_M1031_g N_VPWR_c_1611_n 0.0104579f $X=6.445 $Y=2.525 $X2=0
+ $Y2=0
cc_657 N_A_1274_401#_c_745_n N_VPWR_c_1611_n 0.025438f $X=7.005 $Y=2.047 $X2=0
+ $Y2=0
cc_658 N_A_1274_401#_c_751_n N_VPWR_c_1611_n 0.00174265f $X=6.51 $Y=1.99 $X2=0
+ $Y2=0
cc_659 N_A_1274_401#_c_746_n N_VPWR_c_1616_n 0.0933781f $X=9.305 $Y=2.385 $X2=0
+ $Y2=0
cc_660 N_A_1274_401#_c_747_n N_VPWR_c_1617_n 0.00740629f $X=7.48 $Y=2.385 $X2=0
+ $Y2=0
cc_661 N_A_1274_401#_M1031_g N_VPWR_c_1608_n 8.51577e-19 $X=6.445 $Y=2.525 $X2=0
+ $Y2=0
cc_662 N_A_1274_401#_c_746_n N_VPWR_c_1608_n 0.0265544f $X=9.305 $Y=2.385 $X2=0
+ $Y2=0
cc_663 N_A_1274_401#_c_747_n N_VPWR_c_1608_n 0.0120286f $X=7.48 $Y=2.385 $X2=0
+ $Y2=0
cc_664 N_A_1274_401#_c_746_n A_1818_379# 0.00488734f $X=9.305 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_665 N_A_1274_401#_c_766_n A_1818_379# 0.00487705f $X=9.39 $Y=2.3 $X2=-0.19
+ $Y2=-0.245
cc_666 N_A_1274_401#_c_749_n A_1818_379# 4.96617e-19 $X=9.475 $Y=1.865 $X2=-0.19
+ $Y2=-0.245
cc_667 N_A_1274_401#_c_738_n N_VGND_M1041_d 0.0146293f $X=8.515 $Y=0.745 $X2=0
+ $Y2=0
cc_668 N_A_1274_401#_c_739_n N_VGND_M1041_d 0.00546782f $X=8.6 $Y=1.08 $X2=0
+ $Y2=0
cc_669 N_A_1274_401#_c_740_n N_VGND_M1041_d 0.00472249f $X=9.96 $Y=1.165 $X2=0
+ $Y2=0
cc_670 N_A_1274_401#_M1015_g N_VGND_c_1934_n 0.00912632f $X=6.51 $Y=0.805 $X2=0
+ $Y2=0
cc_671 N_A_1274_401#_c_738_n N_VGND_c_1935_n 0.0180968f $X=8.515 $Y=0.745 $X2=0
+ $Y2=0
cc_672 N_A_1274_401#_c_739_n N_VGND_c_1935_n 0.00400778f $X=8.6 $Y=1.08 $X2=0
+ $Y2=0
cc_673 N_A_1274_401#_c_740_n N_VGND_c_1935_n 0.0144005f $X=9.96 $Y=1.165 $X2=0
+ $Y2=0
cc_674 N_A_1274_401#_c_738_n N_VGND_c_1949_n 0.0205444f $X=8.515 $Y=0.745 $X2=0
+ $Y2=0
cc_675 N_A_1274_401#_M1015_g N_VGND_c_1953_n 7.88961e-19 $X=6.51 $Y=0.805 $X2=0
+ $Y2=0
cc_676 N_A_1274_401#_c_738_n N_VGND_c_1953_n 0.03142f $X=8.515 $Y=0.745 $X2=0
+ $Y2=0
cc_677 N_A_1274_401#_c_738_n A_1575_119# 0.00236933f $X=8.515 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_678 N_A_1274_401#_c_740_n A_1848_119# 0.00366293f $X=9.96 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_679 N_A_1146_463#_M1004_g N_SET_B_c_1012_n 0.0207932f $X=7.1 $Y=2.525
+ $X2=-0.19 $Y2=-0.245
cc_680 N_A_1146_463#_c_868_n N_SET_B_c_1012_n 0.0082113f $X=7.725 $Y=1.2
+ $X2=-0.19 $Y2=-0.245
cc_681 N_A_1146_463#_M1004_g N_SET_B_M1010_g 0.0151842f $X=7.1 $Y=2.525 $X2=0
+ $Y2=0
cc_682 N_A_1146_463#_c_878_n N_SET_B_c_1014_n 8.9408e-19 $X=8.165 $Y=1.115 $X2=0
+ $Y2=0
cc_683 N_A_1146_463#_c_869_n N_SET_B_M1041_g 0.0526152f $X=7.8 $Y=1.125 $X2=0
+ $Y2=0
cc_684 N_A_1146_463#_M1019_g N_SET_B_M1041_g 0.00663354f $X=9.015 $Y=2.315 $X2=0
+ $Y2=0
cc_685 N_A_1146_463#_c_873_n N_SET_B_M1041_g 0.0218021f $X=8.94 $Y=1.515 $X2=0
+ $Y2=0
cc_686 N_A_1146_463#_c_878_n N_SET_B_M1041_g 0.0112352f $X=8.165 $Y=1.115 $X2=0
+ $Y2=0
cc_687 N_A_1146_463#_c_879_n N_SET_B_M1041_g 0.00901501f $X=8.25 $Y=1.42 $X2=0
+ $Y2=0
cc_688 N_A_1146_463#_c_880_n N_SET_B_M1041_g 0.0053499f $X=8.335 $Y=1.515 $X2=0
+ $Y2=0
cc_689 N_A_1146_463#_M1019_g N_SET_B_c_1017_n 0.00627024f $X=9.015 $Y=2.315
+ $X2=0 $Y2=0
cc_690 N_A_1146_463#_M1004_g N_SET_B_c_1019_n 0.00314611f $X=7.1 $Y=2.525 $X2=0
+ $Y2=0
cc_691 N_A_1146_463#_c_887_n N_A_640_481#_c_1139_n 0.00312067f $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_692 N_A_1146_463#_c_875_n N_A_640_481#_M1024_g 0.0128835f $X=6.1 $Y=1.115
+ $X2=0 $Y2=0
cc_693 N_A_1146_463#_c_869_n N_A_640_481#_c_1131_n 0.00978449f $X=7.8 $Y=1.125
+ $X2=0 $Y2=0
cc_694 N_A_1146_463#_c_871_n N_A_640_481#_c_1131_n 0.0104164f $X=9.165 $Y=1.35
+ $X2=0 $Y2=0
cc_695 N_A_1146_463#_c_904_n N_A_640_481#_c_1131_n 0.00335508f $X=5.935 $Y=0.805
+ $X2=0 $Y2=0
cc_696 N_A_1146_463#_c_876_n N_A_640_481#_c_1131_n 6.85903e-19 $X=7.155 $Y=0.69
+ $X2=0 $Y2=0
cc_697 N_A_1146_463#_c_877_n N_A_640_481#_c_1131_n 0.015841f $X=7.155 $Y=0.69
+ $X2=0 $Y2=0
cc_698 N_A_1146_463#_c_887_n N_A_640_481#_M1000_g 0.0105414f $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_699 N_A_1146_463#_M1004_g N_A_640_481#_c_1142_n 0.00979048f $X=7.1 $Y=2.525
+ $X2=0 $Y2=0
cc_700 N_A_1146_463#_M1019_g N_A_640_481#_c_1142_n 0.0100709f $X=9.015 $Y=2.315
+ $X2=0 $Y2=0
cc_701 N_A_1146_463#_M1019_g N_A_640_481#_M1040_g 0.0315321f $X=9.015 $Y=2.315
+ $X2=0 $Y2=0
cc_702 N_A_1146_463#_c_871_n N_A_1920_119#_c_1376_n 7.50289e-19 $X=9.165 $Y=1.35
+ $X2=0 $Y2=0
cc_703 N_A_1146_463#_M1004_g N_VPWR_c_1611_n 0.00569408f $X=7.1 $Y=2.525 $X2=0
+ $Y2=0
cc_704 N_A_1146_463#_c_887_n N_VPWR_c_1611_n 0.0107323f $X=5.87 $Y=2.525 $X2=0
+ $Y2=0
cc_705 N_A_1146_463#_c_887_n N_VPWR_c_1614_n 0.00453007f $X=5.87 $Y=2.525 $X2=0
+ $Y2=0
cc_706 N_A_1146_463#_M1004_g N_VPWR_c_1608_n 9.39239e-19 $X=7.1 $Y=2.525 $X2=0
+ $Y2=0
cc_707 N_A_1146_463#_M1019_g N_VPWR_c_1608_n 9.39239e-19 $X=9.015 $Y=2.315 $X2=0
+ $Y2=0
cc_708 N_A_1146_463#_c_887_n N_VPWR_c_1608_n 0.00751411f $X=5.87 $Y=2.525 $X2=0
+ $Y2=0
cc_709 N_A_1146_463#_M1019_g N_VPWR_c_1632_n 0.00783343f $X=9.015 $Y=2.315 $X2=0
+ $Y2=0
cc_710 N_A_1146_463#_c_904_n N_A_275_481#_c_1773_n 0.00346795f $X=5.935 $Y=0.805
+ $X2=0 $Y2=0
cc_711 N_A_1146_463#_c_875_n N_A_275_481#_c_1773_n 0.00336607f $X=6.1 $Y=1.115
+ $X2=0 $Y2=0
cc_712 N_A_1146_463#_c_887_n N_A_275_481#_c_1774_n 0.0151431f $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_713 N_A_1146_463#_c_875_n N_A_275_481#_c_1774_n 0.0143747f $X=6.1 $Y=1.115
+ $X2=0 $Y2=0
cc_714 N_A_1146_463#_c_882_n N_A_275_481#_c_1774_n 0.0607369f $X=5.83 $Y=1.885
+ $X2=0 $Y2=0
cc_715 N_A_1146_463#_c_904_n N_VGND_c_1934_n 0.00706431f $X=5.935 $Y=0.805 $X2=0
+ $Y2=0
cc_716 N_A_1146_463#_c_874_n N_VGND_c_1934_n 0.0245421f $X=7.06 $Y=1.115 $X2=0
+ $Y2=0
cc_717 N_A_1146_463#_c_876_n N_VGND_c_1934_n 0.025108f $X=7.155 $Y=0.69 $X2=0
+ $Y2=0
cc_718 N_A_1146_463#_c_877_n N_VGND_c_1934_n 0.00305784f $X=7.155 $Y=0.69 $X2=0
+ $Y2=0
cc_719 N_A_1146_463#_c_871_n N_VGND_c_1935_n 0.00523689f $X=9.165 $Y=1.35 $X2=0
+ $Y2=0
cc_720 N_A_1146_463#_c_904_n N_VGND_c_1945_n 0.00419215f $X=5.935 $Y=0.805 $X2=0
+ $Y2=0
cc_721 N_A_1146_463#_c_876_n N_VGND_c_1949_n 0.00441547f $X=7.155 $Y=0.69 $X2=0
+ $Y2=0
cc_722 N_A_1146_463#_c_869_n N_VGND_c_1953_n 9.39239e-19 $X=7.8 $Y=1.125 $X2=0
+ $Y2=0
cc_723 N_A_1146_463#_c_871_n N_VGND_c_1953_n 9.39239e-19 $X=9.165 $Y=1.35 $X2=0
+ $Y2=0
cc_724 N_A_1146_463#_c_904_n N_VGND_c_1953_n 0.00667772f $X=5.935 $Y=0.805 $X2=0
+ $Y2=0
cc_725 N_A_1146_463#_c_876_n N_VGND_c_1953_n 0.00522436f $X=7.155 $Y=0.69 $X2=0
+ $Y2=0
cc_726 N_A_1146_463#_c_877_n N_VGND_c_1953_n 9.07343e-19 $X=7.155 $Y=0.69 $X2=0
+ $Y2=0
cc_727 N_SET_B_M1041_g N_A_640_481#_c_1131_n 0.00978449f $X=8.16 $Y=0.805 $X2=0
+ $Y2=0
cc_728 N_SET_B_M1010_g N_A_640_481#_c_1142_n 0.0100242f $X=7.53 $Y=2.525 $X2=0
+ $Y2=0
cc_729 N_SET_B_c_1017_n N_A_640_481#_M1040_g 0.00716819f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_730 N_SET_B_M1028_g N_A_2067_92#_M1035_g 0.0496019f $X=10.77 $Y=0.8 $X2=0
+ $Y2=0
cc_731 N_SET_B_c_1017_n N_A_2067_92#_M1001_g 0.00152374f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_732 SET_B N_A_2067_92#_M1001_g 3.7234e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_733 N_SET_B_c_1021_n N_A_2067_92#_M1001_g 0.0109645f $X=11.365 $Y=2.035 $X2=0
+ $Y2=0
cc_734 N_SET_B_c_1022_n N_A_2067_92#_M1001_g 0.00182333f $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_735 N_SET_B_c_1010_n N_A_2067_92#_c_1262_n 0.0102543f $X=10.845 $Y=1.215
+ $X2=0 $Y2=0
cc_736 SET_B N_A_2067_92#_c_1262_n 0.00776449f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_737 N_SET_B_c_1021_n N_A_2067_92#_c_1262_n 3.7153e-19 $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_738 N_SET_B_c_1022_n N_A_2067_92#_c_1262_n 0.062493f $X=11.365 $Y=2.035 $X2=0
+ $Y2=0
cc_739 N_SET_B_c_1011_n N_A_2067_92#_c_1262_n 0.0140888f $X=11.365 $Y=1.87 $X2=0
+ $Y2=0
cc_740 N_SET_B_c_1010_n N_A_2067_92#_c_1263_n 0.0185926f $X=10.845 $Y=1.215
+ $X2=0 $Y2=0
cc_741 N_SET_B_c_1017_n N_A_2067_92#_c_1263_n 0.00405182f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_742 SET_B N_A_2067_92#_c_1263_n 0.00786681f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_743 N_SET_B_c_1022_n N_A_2067_92#_c_1263_n 0.00843153f $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_744 N_SET_B_c_1011_n N_A_2067_92#_c_1263_n 0.019011f $X=11.365 $Y=1.87 $X2=0
+ $Y2=0
cc_745 N_SET_B_M1028_g N_A_2067_92#_c_1264_n 0.00426562f $X=10.77 $Y=0.8 $X2=0
+ $Y2=0
cc_746 N_SET_B_c_1009_n N_A_2067_92#_c_1264_n 0.00921093f $X=11.23 $Y=1.215
+ $X2=0 $Y2=0
cc_747 N_SET_B_c_1011_n N_A_2067_92#_c_1264_n 0.011227f $X=11.365 $Y=1.87 $X2=0
+ $Y2=0
cc_748 N_SET_B_M1003_g N_A_2067_92#_c_1270_n 0.00273354f $X=11.275 $Y=2.65 $X2=0
+ $Y2=0
cc_749 N_SET_B_c_1021_n N_A_2067_92#_c_1270_n 0.00462001f $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_750 N_SET_B_c_1022_n N_A_2067_92#_c_1270_n 0.00805685f $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_751 N_SET_B_c_1011_n N_A_2067_92#_c_1270_n 0.0026404f $X=11.365 $Y=1.87 $X2=0
+ $Y2=0
cc_752 N_SET_B_c_1021_n N_A_2067_92#_c_1265_n 0.00360281f $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_753 N_SET_B_c_1011_n N_A_2067_92#_c_1265_n 0.00380406f $X=11.365 $Y=1.87
+ $X2=0 $Y2=0
cc_754 N_SET_B_c_1017_n N_A_1920_119#_M1040_d 0.0032883f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_755 N_SET_B_c_1009_n N_A_1920_119#_M1033_g 0.00887762f $X=11.23 $Y=1.215
+ $X2=0 $Y2=0
cc_756 N_SET_B_c_1011_n N_A_1920_119#_c_1342_n 0.00887762f $X=11.365 $Y=1.87
+ $X2=0 $Y2=0
cc_757 N_SET_B_M1028_g N_A_1920_119#_c_1376_n 8.9164e-19 $X=10.77 $Y=0.8 $X2=0
+ $Y2=0
cc_758 N_SET_B_M1028_g N_A_1920_119#_c_1347_n 0.00250506f $X=10.77 $Y=0.8 $X2=0
+ $Y2=0
cc_759 N_SET_B_c_1017_n N_A_1920_119#_c_1347_n 0.025134f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_760 SET_B N_A_1920_119#_c_1347_n 4.10462e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_761 N_SET_B_c_1022_n N_A_1920_119#_c_1347_n 0.0141212f $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_762 N_SET_B_M1003_g N_A_1920_119#_c_1365_n 0.0143617f $X=11.275 $Y=2.65 $X2=0
+ $Y2=0
cc_763 N_SET_B_c_1017_n N_A_1920_119#_c_1365_n 0.00750503f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_764 SET_B N_A_1920_119#_c_1365_n 0.0081505f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_765 N_SET_B_c_1021_n N_A_1920_119#_c_1365_n 0.00464481f $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_766 N_SET_B_c_1022_n N_A_1920_119#_c_1365_n 0.0635431f $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_767 N_SET_B_c_1017_n N_A_1920_119#_c_1366_n 0.0250142f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_768 SET_B N_A_1920_119#_c_1366_n 0.00115698f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_769 N_SET_B_c_1022_n N_A_1920_119#_c_1366_n 7.32248e-19 $X=11.365 $Y=2.035
+ $X2=0 $Y2=0
cc_770 N_SET_B_M1003_g N_A_1920_119#_c_1367_n 0.00119979f $X=11.275 $Y=2.65
+ $X2=0 $Y2=0
cc_771 N_SET_B_M1003_g N_A_1920_119#_c_1369_n 0.00198317f $X=11.275 $Y=2.65
+ $X2=0 $Y2=0
cc_772 N_SET_B_c_1017_n N_VPWR_M1010_d 0.00414437f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_773 N_SET_B_M1010_g N_VPWR_c_1616_n 0.0079202f $X=7.53 $Y=2.525 $X2=0 $Y2=0
cc_774 N_SET_B_M1003_g N_VPWR_c_1618_n 0.00422592f $X=11.275 $Y=2.65 $X2=0 $Y2=0
cc_775 N_SET_B_M1010_g N_VPWR_c_1608_n 9.39239e-19 $X=7.53 $Y=2.525 $X2=0 $Y2=0
cc_776 N_SET_B_M1003_g N_VPWR_c_1608_n 0.00432128f $X=11.275 $Y=2.65 $X2=0 $Y2=0
cc_777 N_SET_B_M1003_g N_VPWR_c_1633_n 0.00728187f $X=11.275 $Y=2.65 $X2=0 $Y2=0
cc_778 N_SET_B_c_1017_n N_VPWR_c_1633_n 4.21254e-19 $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_779 N_SET_B_c_1017_n A_1818_379# 0.00378377f $X=10.655 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_780 N_SET_B_M1041_g N_VGND_c_1935_n 0.00443606f $X=8.16 $Y=0.805 $X2=0 $Y2=0
cc_781 N_SET_B_M1028_g N_VGND_c_1936_n 0.0112936f $X=10.77 $Y=0.8 $X2=0 $Y2=0
cc_782 N_SET_B_c_1009_n N_VGND_c_1936_n 0.00708939f $X=11.23 $Y=1.215 $X2=0
+ $Y2=0
cc_783 N_SET_B_M1028_g N_VGND_c_1947_n 0.00360926f $X=10.77 $Y=0.8 $X2=0 $Y2=0
cc_784 N_SET_B_M1041_g N_VGND_c_1953_n 9.39239e-19 $X=8.16 $Y=0.805 $X2=0 $Y2=0
cc_785 N_SET_B_M1028_g N_VGND_c_1953_n 0.00402538f $X=10.77 $Y=0.8 $X2=0 $Y2=0
cc_786 N_A_640_481#_M1030_g N_A_2067_92#_M1035_g 0.0428235f $X=10.05 $Y=0.8
+ $X2=0 $Y2=0
cc_787 N_A_640_481#_c_1131_n N_A_1920_119#_c_1376_n 0.00496121f $X=9.975 $Y=0.18
+ $X2=0 $Y2=0
cc_788 N_A_640_481#_M1030_g N_A_1920_119#_c_1376_n 0.015579f $X=10.05 $Y=0.8
+ $X2=0 $Y2=0
cc_789 N_A_640_481#_M1030_g N_A_1920_119#_c_1347_n 0.00177836f $X=10.05 $Y=0.8
+ $X2=0 $Y2=0
cc_790 N_A_640_481#_M1040_g N_A_1920_119#_c_1366_n 8.18186e-19 $X=9.525 $Y=2.44
+ $X2=0 $Y2=0
cc_791 N_A_640_481#_c_1145_n N_VPWR_M1017_s 0.00542835f $X=3.925 $Y=2.332 $X2=0
+ $Y2=0
cc_792 N_A_640_481#_c_1136_n N_VPWR_M1017_s 4.51595e-19 $X=4.04 $Y=1.06 $X2=0
+ $Y2=0
cc_793 N_A_640_481#_M1000_g N_VPWR_c_1611_n 0.00819663f $X=6.085 $Y=2.525 $X2=0
+ $Y2=0
cc_794 N_A_640_481#_c_1142_n N_VPWR_c_1611_n 0.0258744f $X=9.45 $Y=3.15 $X2=0
+ $Y2=0
cc_795 N_A_640_481#_c_1140_n N_VPWR_c_1614_n 0.0607245f $X=4.505 $Y=3.15 $X2=0
+ $Y2=0
cc_796 N_A_640_481#_c_1142_n N_VPWR_c_1616_n 0.0248186f $X=9.45 $Y=3.15 $X2=0
+ $Y2=0
cc_797 N_A_640_481#_c_1142_n N_VPWR_c_1617_n 0.0236757f $X=9.45 $Y=3.15 $X2=0
+ $Y2=0
cc_798 N_A_640_481#_c_1142_n N_VPWR_c_1625_n 0.0248635f $X=9.45 $Y=3.15 $X2=0
+ $Y2=0
cc_799 N_A_640_481#_c_1142_n N_VPWR_c_1626_n 0.026094f $X=9.45 $Y=3.15 $X2=0
+ $Y2=0
cc_800 N_A_640_481#_c_1139_n N_VPWR_c_1608_n 0.04073f $X=6.01 $Y=3.15 $X2=0
+ $Y2=0
cc_801 N_A_640_481#_c_1140_n N_VPWR_c_1608_n 0.00635961f $X=4.505 $Y=3.15 $X2=0
+ $Y2=0
cc_802 N_A_640_481#_c_1142_n N_VPWR_c_1608_n 0.0704171f $X=9.45 $Y=3.15 $X2=0
+ $Y2=0
cc_803 N_A_640_481#_c_1144_n N_VPWR_c_1608_n 0.00847591f $X=6.085 $Y=3.15 $X2=0
+ $Y2=0
cc_804 N_A_640_481#_M1017_g N_VPWR_c_1631_n 0.0106378f $X=4.43 $Y=2.525 $X2=0
+ $Y2=0
cc_805 N_A_640_481#_c_1142_n N_VPWR_c_1632_n 0.0248186f $X=9.45 $Y=3.15 $X2=0
+ $Y2=0
cc_806 N_A_640_481#_M1040_g N_VPWR_c_1632_n 0.00617305f $X=9.525 $Y=2.44 $X2=0
+ $Y2=0
cc_807 N_A_640_481#_c_1146_n N_A_275_481#_c_1772_n 0.0150923f $X=3.435 $Y=2.332
+ $X2=0 $Y2=0
cc_808 N_A_640_481#_M1009_d N_A_275_481#_c_1776_n 0.00310085f $X=3.2 $Y=2.405
+ $X2=0 $Y2=0
cc_809 N_A_640_481#_c_1231_p N_A_275_481#_c_1776_n 0.013177f $X=3.34 $Y=2.56
+ $X2=0 $Y2=0
cc_810 N_A_640_481#_c_1145_n N_A_275_481#_c_1776_n 0.00641687f $X=3.925 $Y=2.332
+ $X2=0 $Y2=0
cc_811 N_A_640_481#_M1017_g N_A_275_481#_c_1778_n 0.0192241f $X=4.43 $Y=2.525
+ $X2=0 $Y2=0
cc_812 N_A_640_481#_c_1139_n N_A_275_481#_c_1778_n 0.0129855f $X=6.01 $Y=3.15
+ $X2=0 $Y2=0
cc_813 N_A_640_481#_c_1145_n N_A_275_481#_c_1778_n 0.026692f $X=3.925 $Y=2.332
+ $X2=0 $Y2=0
cc_814 N_A_640_481#_c_1128_n N_A_275_481#_c_1773_n 0.00592128f $X=5.645 $Y=0.18
+ $X2=0 $Y2=0
cc_815 N_A_640_481#_M1024_g N_A_275_481#_c_1773_n 0.00662626f $X=5.72 $Y=0.805
+ $X2=0 $Y2=0
cc_816 N_A_640_481#_M1017_g N_A_275_481#_c_1779_n 0.00428509f $X=4.43 $Y=2.525
+ $X2=0 $Y2=0
cc_817 N_A_640_481#_c_1231_p N_A_275_481#_c_1779_n 0.00820338f $X=3.34 $Y=2.56
+ $X2=0 $Y2=0
cc_818 N_A_640_481#_c_1145_n N_A_275_481#_c_1779_n 0.0133487f $X=3.925 $Y=2.332
+ $X2=0 $Y2=0
cc_819 N_A_640_481#_c_1139_n N_A_275_481#_c_1780_n 0.00611256f $X=6.01 $Y=3.15
+ $X2=0 $Y2=0
cc_820 N_A_640_481#_M1024_g N_A_275_481#_c_1774_n 7.42931e-19 $X=5.72 $Y=0.805
+ $X2=0 $Y2=0
cc_821 N_A_640_481#_c_1124_n N_VGND_c_1933_n 0.00866424f $X=4.55 $Y=0.97 $X2=0
+ $Y2=0
cc_822 N_A_640_481#_c_1129_n N_VGND_c_1933_n 0.0108372f $X=4.7 $Y=0.18 $X2=0
+ $Y2=0
cc_823 N_A_640_481#_c_1135_n N_VGND_c_1933_n 0.0281203f $X=3.925 $Y=0.495 $X2=0
+ $Y2=0
cc_824 N_A_640_481#_c_1136_n N_VGND_c_1933_n 0.0053397f $X=4.04 $Y=1.06 $X2=0
+ $Y2=0
cc_825 N_A_640_481#_c_1131_n N_VGND_c_1934_n 0.0255466f $X=9.975 $Y=0.18 $X2=0
+ $Y2=0
cc_826 N_A_640_481#_c_1131_n N_VGND_c_1935_n 0.0186949f $X=9.975 $Y=0.18 $X2=0
+ $Y2=0
cc_827 N_A_640_481#_c_1131_n N_VGND_c_1936_n 0.0064106f $X=9.975 $Y=0.18 $X2=0
+ $Y2=0
cc_828 N_A_640_481#_c_1135_n N_VGND_c_1943_n 0.0383115f $X=3.925 $Y=0.495 $X2=0
+ $Y2=0
cc_829 N_A_640_481#_c_1129_n N_VGND_c_1945_n 0.0616402f $X=4.7 $Y=0.18 $X2=0
+ $Y2=0
cc_830 N_A_640_481#_c_1131_n N_VGND_c_1947_n 0.0327748f $X=9.975 $Y=0.18 $X2=0
+ $Y2=0
cc_831 N_A_640_481#_c_1131_n N_VGND_c_1949_n 0.0535816f $X=9.975 $Y=0.18 $X2=0
+ $Y2=0
cc_832 N_A_640_481#_M1023_d N_VGND_c_1953_n 0.0026808f $X=3.245 $Y=0.235 $X2=0
+ $Y2=0
cc_833 N_A_640_481#_c_1128_n N_VGND_c_1953_n 0.0315689f $X=5.645 $Y=0.18 $X2=0
+ $Y2=0
cc_834 N_A_640_481#_c_1129_n N_VGND_c_1953_n 0.0113744f $X=4.7 $Y=0.18 $X2=0
+ $Y2=0
cc_835 N_A_640_481#_c_1131_n N_VGND_c_1953_n 0.131777f $X=9.975 $Y=0.18 $X2=0
+ $Y2=0
cc_836 N_A_640_481#_c_1134_n N_VGND_c_1953_n 0.00842121f $X=5.72 $Y=0.18 $X2=0
+ $Y2=0
cc_837 N_A_640_481#_c_1135_n N_VGND_c_1953_n 0.0306558f $X=3.925 $Y=0.495 $X2=0
+ $Y2=0
cc_838 N_A_2067_92#_c_1264_n N_A_1920_119#_M1033_g 0.00987996f $X=11.6 $Y=0.96
+ $X2=0 $Y2=0
cc_839 N_A_2067_92#_c_1265_n N_A_1920_119#_M1033_g 0.0113999f $X=12.062 $Y=1.622
+ $X2=0 $Y2=0
cc_840 N_A_2067_92#_c_1270_n N_A_1920_119#_c_1341_n 0.00341502f $X=12.062
+ $Y=2.465 $X2=0 $Y2=0
cc_841 N_A_2067_92#_c_1265_n N_A_1920_119#_c_1341_n 0.01211f $X=12.062 $Y=1.622
+ $X2=0 $Y2=0
cc_842 N_A_2067_92#_c_1265_n N_A_1920_119#_c_1342_n 0.00639904f $X=12.062
+ $Y=1.622 $X2=0 $Y2=0
cc_843 N_A_2067_92#_c_1270_n N_A_1920_119#_M1016_g 0.00383727f $X=12.062
+ $Y=2.465 $X2=0 $Y2=0
cc_844 N_A_2067_92#_c_1272_n N_A_1920_119#_M1016_g 0.00356526f $X=12.18 $Y=2.63
+ $X2=0 $Y2=0
cc_845 N_A_2067_92#_c_1265_n N_A_1920_119#_M1002_g 5.12329e-19 $X=12.062
+ $Y=1.622 $X2=0 $Y2=0
cc_846 N_A_2067_92#_M1035_g N_A_1920_119#_c_1376_n 0.0109127f $X=10.41 $Y=0.8
+ $X2=0 $Y2=0
cc_847 N_A_2067_92#_M1035_g N_A_1920_119#_c_1347_n 0.0241091f $X=10.41 $Y=0.8
+ $X2=0 $Y2=0
cc_848 N_A_2067_92#_M1001_g N_A_1920_119#_c_1347_n 0.00810268f $X=10.41 $Y=2.65
+ $X2=0 $Y2=0
cc_849 N_A_2067_92#_c_1261_n N_A_1920_119#_c_1347_n 0.0120986f $X=10.41 $Y=1.665
+ $X2=0 $Y2=0
cc_850 N_A_2067_92#_c_1262_n N_A_1920_119#_c_1347_n 0.0183896f $X=11.375
+ $Y=1.622 $X2=0 $Y2=0
cc_851 N_A_2067_92#_M1001_g N_A_1920_119#_c_1365_n 0.00356302f $X=10.41 $Y=2.65
+ $X2=0 $Y2=0
cc_852 N_A_2067_92#_c_1263_n N_A_1920_119#_c_1365_n 0.00493371f $X=10.825
+ $Y=1.665 $X2=0 $Y2=0
cc_853 N_A_2067_92#_c_1270_n N_A_1920_119#_c_1365_n 0.00899269f $X=12.062
+ $Y=2.465 $X2=0 $Y2=0
cc_854 N_A_2067_92#_c_1265_n N_A_1920_119#_c_1365_n 0.00479695f $X=12.062
+ $Y=1.622 $X2=0 $Y2=0
cc_855 N_A_2067_92#_M1001_g N_A_1920_119#_c_1366_n 0.0195129f $X=10.41 $Y=2.65
+ $X2=0 $Y2=0
cc_856 N_A_2067_92#_c_1272_n N_A_1920_119#_c_1367_n 0.0140686f $X=12.18 $Y=2.63
+ $X2=0 $Y2=0
cc_857 N_A_2067_92#_c_1272_n N_A_1920_119#_c_1368_n 0.0245975f $X=12.18 $Y=2.63
+ $X2=0 $Y2=0
cc_858 N_A_2067_92#_c_1270_n N_A_1920_119#_c_1348_n 0.0392691f $X=12.062
+ $Y=2.465 $X2=0 $Y2=0
cc_859 N_A_2067_92#_c_1265_n N_A_1920_119#_c_1348_n 0.0131024f $X=12.062
+ $Y=1.622 $X2=0 $Y2=0
cc_860 N_A_2067_92#_c_1272_n N_A_1920_119#_c_1348_n 0.00165852f $X=12.18 $Y=2.63
+ $X2=0 $Y2=0
cc_861 N_A_2067_92#_c_1270_n N_A_1920_119#_c_1371_n 0.00798365f $X=12.062
+ $Y=2.465 $X2=0 $Y2=0
cc_862 N_A_2067_92#_c_1265_n N_A_1920_119#_c_1349_n 0.00387227f $X=12.062
+ $Y=1.622 $X2=0 $Y2=0
cc_863 N_A_2067_92#_c_1270_n N_A_1920_119#_c_1374_n 0.00356677f $X=12.062
+ $Y=2.465 $X2=0 $Y2=0
cc_864 N_A_2067_92#_M1001_g N_VPWR_c_1626_n 0.00422593f $X=10.41 $Y=2.65 $X2=0
+ $Y2=0
cc_865 N_A_2067_92#_M1001_g N_VPWR_c_1608_n 0.00432128f $X=10.41 $Y=2.65 $X2=0
+ $Y2=0
cc_866 N_A_2067_92#_M1001_g N_VPWR_c_1633_n 0.00865656f $X=10.41 $Y=2.65 $X2=0
+ $Y2=0
cc_867 N_A_2067_92#_M1035_g N_VGND_c_1936_n 0.0017112f $X=10.41 $Y=0.8 $X2=0
+ $Y2=0
cc_868 N_A_2067_92#_c_1262_n N_VGND_c_1936_n 0.0110421f $X=11.375 $Y=1.622 $X2=0
+ $Y2=0
cc_869 N_A_2067_92#_c_1264_n N_VGND_c_1936_n 0.0113573f $X=11.6 $Y=0.96 $X2=0
+ $Y2=0
cc_870 N_A_2067_92#_c_1265_n N_VGND_c_1937_n 0.0101004f $X=12.062 $Y=1.622 $X2=0
+ $Y2=0
cc_871 N_A_2067_92#_M1035_g N_VGND_c_1947_n 0.00338477f $X=10.41 $Y=0.8 $X2=0
+ $Y2=0
cc_872 N_A_2067_92#_M1035_g N_VGND_c_1953_n 0.00479212f $X=10.41 $Y=0.8 $X2=0
+ $Y2=0
cc_873 N_A_2067_92#_c_1264_n N_VGND_c_1953_n 0.0145247f $X=11.6 $Y=0.96 $X2=0
+ $Y2=0
cc_874 N_A_1920_119#_c_1352_n N_A_2582_150#_c_1545_n 0.00585139f $X=14.665
+ $Y=0.765 $X2=0 $Y2=0
cc_875 N_A_1920_119#_c_1355_n N_A_2582_150#_c_1545_n 3.65735e-19 $X=13.57
+ $Y=0.415 $X2=0 $Y2=0
cc_876 N_A_1920_119#_c_1352_n N_A_2582_150#_c_1546_n 0.0171697f $X=14.665
+ $Y=0.765 $X2=0 $Y2=0
cc_877 N_A_1920_119#_c_1353_n N_A_2582_150#_c_1546_n 0.00571257f $X=14.75
+ $Y=1.505 $X2=0 $Y2=0
cc_878 N_A_1920_119#_c_1441_p N_A_2582_150#_c_1546_n 0.00200094f $X=13.57
+ $Y=0.415 $X2=0 $Y2=0
cc_879 N_A_1920_119#_c_1355_n N_A_2582_150#_c_1546_n 0.0165059f $X=13.57
+ $Y=0.415 $X2=0 $Y2=0
cc_880 N_A_1920_119#_c_1356_n N_A_2582_150#_c_1546_n 0.0241269f $X=14.772
+ $Y=1.34 $X2=0 $Y2=0
cc_881 N_A_1920_119#_M1007_g N_A_2582_150#_M1027_g 0.0199652f $X=14.725 $Y=2.465
+ $X2=0 $Y2=0
cc_882 N_A_1920_119#_c_1353_n N_A_2582_150#_c_1548_n 0.00110581f $X=14.75
+ $Y=1.505 $X2=0 $Y2=0
cc_883 N_A_1920_119#_c_1354_n N_A_2582_150#_c_1548_n 0.020418f $X=14.75 $Y=1.505
+ $X2=0 $Y2=0
cc_884 N_A_1920_119#_c_1344_n N_A_2582_150#_c_1549_n 0.00488638f $X=13.405
+ $Y=0.6 $X2=0 $Y2=0
cc_885 N_A_1920_119#_c_1350_n N_A_2582_150#_c_1549_n 0.0195112f $X=13.405
+ $Y=0.535 $X2=0 $Y2=0
cc_886 N_A_1920_119#_c_1441_p N_A_2582_150#_c_1549_n 0.00467366f $X=13.57
+ $Y=0.415 $X2=0 $Y2=0
cc_887 N_A_1920_119#_c_1355_n N_A_2582_150#_c_1549_n 0.00234459f $X=13.57
+ $Y=0.415 $X2=0 $Y2=0
cc_888 N_A_1920_119#_c_1360_n N_A_2582_150#_c_1550_n 0.00642072f $X=13.09
+ $Y=2.05 $X2=0 $Y2=0
cc_889 N_A_1920_119#_M1002_g N_A_2582_150#_c_1550_n 0.00173232f $X=12.835
+ $Y=0.96 $X2=0 $Y2=0
cc_890 N_A_1920_119#_c_1344_n N_A_2582_150#_c_1550_n 0.00126559f $X=13.405
+ $Y=0.6 $X2=0 $Y2=0
cc_891 N_A_1920_119#_c_1349_n N_A_2582_150#_c_1550_n 0.0131188f $X=12.71 $Y=1.59
+ $X2=0 $Y2=0
cc_892 N_A_1920_119#_c_1350_n N_A_2582_150#_c_1550_n 0.00509733f $X=13.405
+ $Y=0.535 $X2=0 $Y2=0
cc_893 N_A_1920_119#_c_1441_p N_A_2582_150#_c_1550_n 0.0119044f $X=13.57
+ $Y=0.415 $X2=0 $Y2=0
cc_894 N_A_1920_119#_c_1355_n N_A_2582_150#_c_1550_n 0.00114489f $X=13.57
+ $Y=0.415 $X2=0 $Y2=0
cc_895 N_A_1920_119#_M1002_g N_A_2582_150#_c_1551_n 0.00182147f $X=12.835
+ $Y=0.96 $X2=0 $Y2=0
cc_896 N_A_1920_119#_c_1348_n N_A_2582_150#_c_1551_n 0.0164307f $X=12.6 $Y=2.26
+ $X2=0 $Y2=0
cc_897 N_A_1920_119#_c_1349_n N_A_2582_150#_c_1551_n 0.00901245f $X=12.71
+ $Y=1.59 $X2=0 $Y2=0
cc_898 N_A_1920_119#_c_1360_n N_A_2582_150#_c_1554_n 0.00791869f $X=13.09
+ $Y=2.05 $X2=0 $Y2=0
cc_899 N_A_1920_119#_c_1348_n N_A_2582_150#_c_1554_n 0.0053112f $X=12.6 $Y=2.26
+ $X2=0 $Y2=0
cc_900 N_A_1920_119#_c_1374_n N_A_2582_150#_c_1554_n 2.5501e-19 $X=12.5 $Y=1.755
+ $X2=0 $Y2=0
cc_901 N_A_1920_119#_M1002_g N_A_2582_150#_c_1552_n 0.0056542f $X=12.835 $Y=0.96
+ $X2=0 $Y2=0
cc_902 N_A_1920_119#_c_1346_n N_A_2582_150#_c_1552_n 0.0056542f $X=12.835
+ $Y=1.665 $X2=0 $Y2=0
cc_903 N_A_1920_119#_c_1348_n N_A_2582_150#_c_1552_n 6.14882e-19 $X=12.6 $Y=2.26
+ $X2=0 $Y2=0
cc_904 N_A_1920_119#_c_1349_n N_A_2582_150#_c_1552_n 3.43457e-19 $X=12.71
+ $Y=1.59 $X2=0 $Y2=0
cc_905 N_A_1920_119#_c_1441_p N_A_2582_150#_c_1552_n 0.00136298f $X=13.57
+ $Y=0.415 $X2=0 $Y2=0
cc_906 N_A_1920_119#_c_1355_n N_A_2582_150#_c_1552_n 0.0191884f $X=13.57
+ $Y=0.415 $X2=0 $Y2=0
cc_907 N_A_1920_119#_c_1346_n N_A_2582_150#_c_1556_n 0.00182147f $X=12.835
+ $Y=1.665 $X2=0 $Y2=0
cc_908 N_A_1920_119#_c_1365_n N_VPWR_M1001_d 0.00688095f $X=11.395 $Y=2.385
+ $X2=0 $Y2=0
cc_909 N_A_1920_119#_c_1371_n N_VPWR_M1016_d 0.00654931f $X=12.6 $Y=2.905 $X2=0
+ $Y2=0
cc_910 N_A_1920_119#_M1016_g N_VPWR_c_1612_n 0.00120832f $X=12.395 $Y=2.63 $X2=0
+ $Y2=0
cc_911 N_A_1920_119#_c_1360_n N_VPWR_c_1612_n 0.0108858f $X=13.09 $Y=2.05 $X2=0
+ $Y2=0
cc_912 N_A_1920_119#_c_1361_n N_VPWR_c_1612_n 0.0156877f $X=13.165 $Y=2.125
+ $X2=0 $Y2=0
cc_913 N_A_1920_119#_c_1368_n N_VPWR_c_1612_n 0.0147862f $X=12.515 $Y=2.99 $X2=0
+ $Y2=0
cc_914 N_A_1920_119#_c_1348_n N_VPWR_c_1612_n 0.00653726f $X=12.6 $Y=2.26 $X2=0
+ $Y2=0
cc_915 N_A_1920_119#_c_1371_n N_VPWR_c_1612_n 0.0487061f $X=12.6 $Y=2.905 $X2=0
+ $Y2=0
cc_916 N_A_1920_119#_c_1375_n N_VPWR_c_1612_n 2.86816e-19 $X=12.492 $Y=2.05
+ $X2=0 $Y2=0
cc_917 N_A_1920_119#_M1007_g N_VPWR_c_1613_n 0.00366932f $X=14.725 $Y=2.465
+ $X2=0 $Y2=0
cc_918 N_A_1920_119#_c_1354_n N_VPWR_c_1613_n 7.8075e-19 $X=14.75 $Y=1.505 $X2=0
+ $Y2=0
cc_919 N_A_1920_119#_M1016_g N_VPWR_c_1618_n 7.26245e-19 $X=12.395 $Y=2.63 $X2=0
+ $Y2=0
cc_920 N_A_1920_119#_c_1368_n N_VPWR_c_1618_n 0.0675282f $X=12.515 $Y=2.99 $X2=0
+ $Y2=0
cc_921 N_A_1920_119#_c_1369_n N_VPWR_c_1618_n 0.0186386f $X=11.655 $Y=2.99 $X2=0
+ $Y2=0
cc_922 N_A_1920_119#_c_1361_n N_VPWR_c_1620_n 0.00410575f $X=13.165 $Y=2.125
+ $X2=0 $Y2=0
cc_923 N_A_1920_119#_c_1366_n N_VPWR_c_1626_n 0.0156375f $X=10.48 $Y=2.385 $X2=0
+ $Y2=0
cc_924 N_A_1920_119#_M1007_g N_VPWR_c_1627_n 0.00585385f $X=14.725 $Y=2.465
+ $X2=0 $Y2=0
cc_925 N_A_1920_119#_c_1361_n N_VPWR_c_1608_n 0.00427039f $X=13.165 $Y=2.125
+ $X2=0 $Y2=0
cc_926 N_A_1920_119#_M1007_g N_VPWR_c_1608_n 0.0116689f $X=14.725 $Y=2.465 $X2=0
+ $Y2=0
cc_927 N_A_1920_119#_c_1365_n N_VPWR_c_1608_n 0.00764841f $X=11.395 $Y=2.385
+ $X2=0 $Y2=0
cc_928 N_A_1920_119#_c_1366_n N_VPWR_c_1608_n 0.0285712f $X=10.48 $Y=2.385 $X2=0
+ $Y2=0
cc_929 N_A_1920_119#_c_1368_n N_VPWR_c_1608_n 0.0389353f $X=12.515 $Y=2.99 $X2=0
+ $Y2=0
cc_930 N_A_1920_119#_c_1369_n N_VPWR_c_1608_n 0.0101082f $X=11.655 $Y=2.99 $X2=0
+ $Y2=0
cc_931 N_A_1920_119#_c_1365_n N_VPWR_c_1633_n 0.0486856f $X=11.395 $Y=2.385
+ $X2=0 $Y2=0
cc_932 N_A_1920_119#_c_1366_n N_VPWR_c_1633_n 0.00827853f $X=10.48 $Y=2.385
+ $X2=0 $Y2=0
cc_933 N_A_1920_119#_c_1367_n N_VPWR_c_1633_n 0.0128358f $X=11.49 $Y=2.655 $X2=0
+ $Y2=0
cc_934 N_A_1920_119#_c_1369_n N_VPWR_c_1633_n 0.0154742f $X=11.655 $Y=2.99 $X2=0
+ $Y2=0
cc_935 N_A_1920_119#_c_1366_n A_2025_488# 0.00214129f $X=10.48 $Y=2.385
+ $X2=-0.19 $Y2=-0.245
cc_936 N_A_1920_119#_c_1352_n N_Q_M1020_s 0.00729794f $X=14.665 $Y=0.765
+ $X2=-0.19 $Y2=-0.245
cc_937 N_A_1920_119#_c_1361_n N_Q_c_1898_n 0.00432728f $X=13.165 $Y=2.125 $X2=0
+ $Y2=0
cc_938 N_A_1920_119#_M1007_g N_Q_c_1898_n 0.00118725f $X=14.725 $Y=2.465 $X2=0
+ $Y2=0
cc_939 N_A_1920_119#_c_1352_n N_Q_c_1898_n 0.0223214f $X=14.665 $Y=0.765 $X2=0
+ $Y2=0
cc_940 N_A_1920_119#_c_1353_n N_Q_c_1898_n 0.0234802f $X=14.75 $Y=1.505 $X2=0
+ $Y2=0
cc_941 N_A_1920_119#_c_1354_n N_Q_c_1898_n 0.00103497f $X=14.75 $Y=1.505 $X2=0
+ $Y2=0
cc_942 N_A_1920_119#_c_1356_n N_Q_c_1898_n 2.87106e-19 $X=14.772 $Y=1.34 $X2=0
+ $Y2=0
cc_943 N_A_1920_119#_M1007_g Q_N 0.00580777f $X=14.725 $Y=2.465 $X2=0 $Y2=0
cc_944 N_A_1920_119#_c_1353_n Q_N 0.0454404f $X=14.75 $Y=1.505 $X2=0 $Y2=0
cc_945 N_A_1920_119#_c_1356_n Q_N 0.014513f $X=14.772 $Y=1.34 $X2=0 $Y2=0
cc_946 N_A_1920_119#_c_1354_n Q_N 0.00549175f $X=14.75 $Y=1.505 $X2=0 $Y2=0
cc_947 N_A_1920_119#_c_1349_n N_VGND_M1033_d 0.00695051f $X=12.71 $Y=1.59 $X2=0
+ $Y2=0
cc_948 N_A_1920_119#_c_1352_n N_VGND_M1020_d 0.0113627f $X=14.665 $Y=0.765 $X2=0
+ $Y2=0
cc_949 N_A_1920_119#_c_1353_n N_VGND_M1020_d 0.00485333f $X=14.75 $Y=1.505 $X2=0
+ $Y2=0
cc_950 N_A_1920_119#_M1033_g N_VGND_c_1936_n 0.00412438f $X=11.815 $Y=0.96 $X2=0
+ $Y2=0
cc_951 N_A_1920_119#_c_1376_n N_VGND_c_1936_n 0.0123356f $X=10.31 $Y=0.775 $X2=0
+ $Y2=0
cc_952 N_A_1920_119#_c_1347_n N_VGND_c_1936_n 0.00202899f $X=10.395 $Y=2.12
+ $X2=0 $Y2=0
cc_953 N_A_1920_119#_M1033_g N_VGND_c_1937_n 0.00611417f $X=11.815 $Y=0.96 $X2=0
+ $Y2=0
cc_954 N_A_1920_119#_c_1341_n N_VGND_c_1937_n 0.00589879f $X=12.32 $Y=1.665
+ $X2=0 $Y2=0
cc_955 N_A_1920_119#_c_1345_n N_VGND_c_1937_n 0.00312337f $X=12.91 $Y=0.6 $X2=0
+ $Y2=0
cc_956 N_A_1920_119#_c_1346_n N_VGND_c_1937_n 8.85401e-19 $X=12.835 $Y=1.665
+ $X2=0 $Y2=0
cc_957 N_A_1920_119#_c_1348_n N_VGND_c_1937_n 0.00495337f $X=12.6 $Y=2.26 $X2=0
+ $Y2=0
cc_958 N_A_1920_119#_c_1349_n N_VGND_c_1937_n 0.036996f $X=12.71 $Y=1.59 $X2=0
+ $Y2=0
cc_959 N_A_1920_119#_c_1351_n N_VGND_c_1937_n 0.0156186f $X=12.795 $Y=0.535
+ $X2=0 $Y2=0
cc_960 N_A_1920_119#_c_1352_n N_VGND_c_1938_n 0.0258699f $X=14.665 $Y=0.765
+ $X2=0 $Y2=0
cc_961 N_A_1920_119#_c_1355_n N_VGND_c_1938_n 8.98847e-19 $X=13.57 $Y=0.415
+ $X2=0 $Y2=0
cc_962 N_A_1920_119#_c_1356_n N_VGND_c_1938_n 0.00433503f $X=14.772 $Y=1.34
+ $X2=0 $Y2=0
cc_963 N_A_1920_119#_c_1376_n N_VGND_c_1947_n 0.0140327f $X=10.31 $Y=0.775 $X2=0
+ $Y2=0
cc_964 N_A_1920_119#_M1033_g N_VGND_c_1950_n 0.00355139f $X=11.815 $Y=0.96 $X2=0
+ $Y2=0
cc_965 N_A_1920_119#_c_1345_n N_VGND_c_1951_n 0.0027651f $X=12.91 $Y=0.6 $X2=0
+ $Y2=0
cc_966 N_A_1920_119#_c_1350_n N_VGND_c_1951_n 0.0175292f $X=13.405 $Y=0.535
+ $X2=0 $Y2=0
cc_967 N_A_1920_119#_c_1351_n N_VGND_c_1951_n 0.00539649f $X=12.795 $Y=0.535
+ $X2=0 $Y2=0
cc_968 N_A_1920_119#_c_1352_n N_VGND_c_1951_n 0.0101137f $X=14.665 $Y=0.765
+ $X2=0 $Y2=0
cc_969 N_A_1920_119#_c_1441_p N_VGND_c_1951_n 0.0146249f $X=13.57 $Y=0.415 $X2=0
+ $Y2=0
cc_970 N_A_1920_119#_c_1355_n N_VGND_c_1951_n 0.00871292f $X=13.57 $Y=0.415
+ $X2=0 $Y2=0
cc_971 N_A_1920_119#_c_1352_n N_VGND_c_1952_n 8.76405e-19 $X=14.665 $Y=0.765
+ $X2=0 $Y2=0
cc_972 N_A_1920_119#_c_1356_n N_VGND_c_1952_n 0.00542213f $X=14.772 $Y=1.34
+ $X2=0 $Y2=0
cc_973 N_A_1920_119#_M1033_g N_VGND_c_1953_n 0.0043622f $X=11.815 $Y=0.96 $X2=0
+ $Y2=0
cc_974 N_A_1920_119#_c_1376_n N_VGND_c_1953_n 0.0238805f $X=10.31 $Y=0.775 $X2=0
+ $Y2=0
cc_975 N_A_1920_119#_c_1350_n N_VGND_c_1953_n 0.0200699f $X=13.405 $Y=0.535
+ $X2=0 $Y2=0
cc_976 N_A_1920_119#_c_1351_n N_VGND_c_1953_n 0.00588742f $X=12.795 $Y=0.535
+ $X2=0 $Y2=0
cc_977 N_A_1920_119#_c_1352_n N_VGND_c_1953_n 0.0226804f $X=14.665 $Y=0.765
+ $X2=0 $Y2=0
cc_978 N_A_1920_119#_c_1441_p N_VGND_c_1953_n 0.0119019f $X=13.57 $Y=0.415 $X2=0
+ $Y2=0
cc_979 N_A_1920_119#_c_1355_n N_VGND_c_1953_n 0.0117998f $X=13.57 $Y=0.415 $X2=0
+ $Y2=0
cc_980 N_A_1920_119#_c_1356_n N_VGND_c_1953_n 0.00539454f $X=14.772 $Y=1.34
+ $X2=0 $Y2=0
cc_981 N_A_1920_119#_c_1376_n A_2025_118# 0.00558226f $X=10.31 $Y=0.775
+ $X2=-0.19 $Y2=-0.245
cc_982 N_A_2582_150#_c_1554_n N_VPWR_c_1612_n 0.0261249f $X=13.38 $Y=2.345 $X2=0
+ $Y2=0
cc_983 N_A_2582_150#_M1027_g N_VPWR_c_1613_n 0.00352797f $X=14.295 $Y=2.465
+ $X2=0 $Y2=0
cc_984 N_A_2582_150#_M1027_g N_VPWR_c_1620_n 0.00541359f $X=14.295 $Y=2.465
+ $X2=0 $Y2=0
cc_985 N_A_2582_150#_c_1554_n N_VPWR_c_1620_n 0.00773544f $X=13.38 $Y=2.345
+ $X2=0 $Y2=0
cc_986 N_A_2582_150#_M1027_g N_VPWR_c_1608_n 0.0109327f $X=14.295 $Y=2.465 $X2=0
+ $Y2=0
cc_987 N_A_2582_150#_c_1554_n N_VPWR_c_1608_n 0.00881366f $X=13.38 $Y=2.345
+ $X2=0 $Y2=0
cc_988 N_A_2582_150#_c_1545_n N_Q_c_1898_n 0.0182241f $X=14.22 $Y=1.415 $X2=0
+ $Y2=0
cc_989 N_A_2582_150#_c_1546_n N_Q_c_1898_n 0.0071643f $X=14.295 $Y=1.34 $X2=0
+ $Y2=0
cc_990 N_A_2582_150#_M1027_g N_Q_c_1898_n 0.0272235f $X=14.295 $Y=2.465 $X2=0
+ $Y2=0
cc_991 N_A_2582_150#_c_1548_n N_Q_c_1898_n 0.00233496f $X=14.295 $Y=1.415 $X2=0
+ $Y2=0
cc_992 N_A_2582_150#_c_1550_n N_Q_c_1898_n 0.0105836f $X=13.475 $Y=1.33 $X2=0
+ $Y2=0
cc_993 N_A_2582_150#_c_1551_n N_Q_c_1898_n 0.0293294f $X=13.475 $Y=1.64 $X2=0
+ $Y2=0
cc_994 N_A_2582_150#_c_1554_n N_Q_c_1898_n 0.0492516f $X=13.38 $Y=2.345 $X2=0
+ $Y2=0
cc_995 N_A_2582_150#_c_1552_n N_Q_c_1898_n 0.00511361f $X=13.56 $Y=1.325 $X2=0
+ $Y2=0
cc_996 N_A_2582_150#_c_1546_n N_VGND_c_1938_n 0.00449987f $X=14.295 $Y=1.34
+ $X2=0 $Y2=0
cc_997 N_A_2582_150#_c_1546_n N_VGND_c_1951_n 0.00436274f $X=14.295 $Y=1.34
+ $X2=0 $Y2=0
cc_998 N_A_2582_150#_c_1546_n N_VGND_c_1953_n 0.00539454f $X=14.295 $Y=1.34
+ $X2=0 $Y2=0
cc_999 N_VPWR_M1011_d N_A_275_481#_c_1785_n 0.0205958f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_1000 N_VPWR_c_1610_n N_A_275_481#_c_1785_n 0.0253821f $X=2.57 $Y=2.92 $X2=0
+ $Y2=0
cc_1001 N_VPWR_c_1623_n N_A_275_481#_c_1785_n 0.00811453f $X=2.405 $Y=3.33 $X2=0
+ $Y2=0
cc_1002 N_VPWR_c_1624_n N_A_275_481#_c_1785_n 0.00265072f $X=3.955 $Y=3.33 $X2=0
+ $Y2=0
cc_1003 N_VPWR_c_1608_n N_A_275_481#_c_1785_n 0.0216138f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1004 N_VPWR_M1011_d N_A_275_481#_c_1772_n 0.00118499f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_1005 N_VPWR_M1011_d N_A_275_481#_c_1806_n 0.00367779f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_1006 N_VPWR_c_1610_n N_A_275_481#_c_1806_n 0.0060774f $X=2.57 $Y=2.92 $X2=0
+ $Y2=0
cc_1007 N_VPWR_c_1624_n N_A_275_481#_c_1776_n 0.0317538f $X=3.955 $Y=3.33 $X2=0
+ $Y2=0
cc_1008 N_VPWR_c_1608_n N_A_275_481#_c_1776_n 0.0192319f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1009 N_VPWR_M1011_d N_A_275_481#_c_1777_n 0.00152369f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_1010 N_VPWR_c_1610_n N_A_275_481#_c_1777_n 0.0145763f $X=2.57 $Y=2.92 $X2=0
+ $Y2=0
cc_1011 N_VPWR_c_1624_n N_A_275_481#_c_1777_n 0.0113112f $X=3.955 $Y=3.33 $X2=0
+ $Y2=0
cc_1012 N_VPWR_c_1608_n N_A_275_481#_c_1777_n 0.0064524f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1013 N_VPWR_M1017_s N_A_275_481#_c_1778_n 0.0127752f $X=3.995 $Y=2.205 $X2=0
+ $Y2=0
cc_1014 N_VPWR_c_1614_n N_A_275_481#_c_1778_n 0.0205101f $X=6.505 $Y=3.33 $X2=0
+ $Y2=0
cc_1015 N_VPWR_c_1624_n N_A_275_481#_c_1778_n 0.00402338f $X=3.955 $Y=3.33 $X2=0
+ $Y2=0
cc_1016 N_VPWR_c_1608_n N_A_275_481#_c_1778_n 0.03385f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1017 N_VPWR_c_1631_n N_A_275_481#_c_1778_n 0.024406f $X=4.12 $Y=3.05 $X2=0
+ $Y2=0
cc_1018 N_VPWR_c_1609_n N_A_275_481#_c_1788_n 0.0168088f $X=0.725 $Y=2.55 $X2=0
+ $Y2=0
cc_1019 N_VPWR_c_1610_n N_A_275_481#_c_1788_n 0.00589986f $X=2.57 $Y=2.92 $X2=0
+ $Y2=0
cc_1020 N_VPWR_c_1623_n N_A_275_481#_c_1788_n 0.0156787f $X=2.405 $Y=3.33 $X2=0
+ $Y2=0
cc_1021 N_VPWR_c_1608_n N_A_275_481#_c_1788_n 0.0122278f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1022 N_VPWR_c_1624_n N_A_275_481#_c_1779_n 0.0109843f $X=3.955 $Y=3.33 $X2=0
+ $Y2=0
cc_1023 N_VPWR_c_1608_n N_A_275_481#_c_1779_n 0.00642982f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1024 N_VPWR_c_1631_n N_A_275_481#_c_1779_n 0.00837701f $X=4.12 $Y=3.05 $X2=0
+ $Y2=0
cc_1025 N_VPWR_c_1614_n N_A_275_481#_c_1780_n 0.00725716f $X=6.505 $Y=3.33 $X2=0
+ $Y2=0
cc_1026 N_VPWR_c_1608_n N_A_275_481#_c_1780_n 0.00839455f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1027 N_VPWR_c_1608_n N_Q_M1027_s 0.00215158f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1028 N_VPWR_c_1620_n N_Q_c_1898_n 0.0213875f $X=14.425 $Y=3.33 $X2=0 $Y2=0
cc_1029 N_VPWR_c_1608_n N_Q_c_1898_n 0.0127404f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1030 N_VPWR_c_1608_n N_Q_N_M1007_d 0.00336915f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1031 N_VPWR_c_1627_n Q_N 0.0303526f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1032 N_VPWR_c_1608_n Q_N 0.0170284f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1033 N_A_275_481#_c_1785_n A_383_481# 0.00281462f $X=2.905 $Y=2.56 $X2=-0.19
+ $Y2=-0.245
cc_1034 N_A_275_481#_c_1771_n N_VGND_M1036_d 0.00181469f $X=2.905 $Y=0.74 $X2=0
+ $Y2=0
cc_1035 N_A_275_481#_c_1770_n N_VGND_c_1931_n 0.0111072f $X=2.37 $Y=0.437 $X2=0
+ $Y2=0
cc_1036 N_A_275_481#_c_1770_n N_VGND_c_1932_n 0.0112538f $X=2.37 $Y=0.437 $X2=0
+ $Y2=0
cc_1037 N_A_275_481#_c_1771_n N_VGND_c_1932_n 0.0189468f $X=2.905 $Y=0.74 $X2=0
+ $Y2=0
cc_1038 N_A_275_481#_c_1770_n N_VGND_c_1941_n 0.0491986f $X=2.37 $Y=0.437 $X2=0
+ $Y2=0
cc_1039 N_A_275_481#_c_1771_n N_VGND_c_1941_n 0.00412567f $X=2.905 $Y=0.74 $X2=0
+ $Y2=0
cc_1040 N_A_275_481#_c_1773_n N_VGND_c_1945_n 0.008976f $X=5.365 $Y=1.035 $X2=0
+ $Y2=0
cc_1041 N_A_275_481#_M1014_d N_VGND_c_1953_n 0.00509637f $X=1.62 $Y=0.235 $X2=0
+ $Y2=0
cc_1042 N_A_275_481#_c_1770_n N_VGND_c_1953_n 0.0347174f $X=2.37 $Y=0.437 $X2=0
+ $Y2=0
cc_1043 N_A_275_481#_c_1771_n N_VGND_c_1953_n 0.00775634f $X=2.905 $Y=0.74 $X2=0
+ $Y2=0
cc_1044 N_A_275_481#_c_1773_n N_VGND_c_1953_n 0.0111108f $X=5.365 $Y=1.035 $X2=0
+ $Y2=0
cc_1045 N_A_275_481#_c_1770_n A_478_47# 0.0048345f $X=2.37 $Y=0.437 $X2=-0.19
+ $Y2=-0.245
cc_1046 Q_N N_VGND_c_1938_n 5.63305e-19 $X=15.035 $Y=0.47 $X2=0 $Y2=0
cc_1047 Q_N N_VGND_c_1952_n 0.0106706f $X=15.035 $Y=0.47 $X2=0 $Y2=0
cc_1048 Q_N N_VGND_c_1953_n 0.00971712f $X=15.035 $Y=0.47 $X2=0 $Y2=0
cc_1049 N_VGND_c_1953_n A_252_47# 0.00284246f $X=15.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1050 N_VGND_c_1953_n A_478_47# 0.00269325f $X=15.12 $Y=0 $X2=-0.19 $Y2=-0.245
