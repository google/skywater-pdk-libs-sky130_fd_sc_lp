* File: sky130_fd_sc_lp__clkbuflp_8.spice
* Created: Wed Sep  2 09:39:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkbuflp_8.pex.spice"
.subckt sky130_fd_sc_lp__clkbuflp_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_M1009_g A_110_47# VNB NSHORT L=0.15 W=0.64 AD=0.1696
+ AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75000.2 SB=75004.5
+ A=0.096 P=1.58 MULT=1
MM1001 A_110_47# N_A_M1001_g N_A_130_417#_M1001_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.5
+ SB=75004.2 A=0.096 P=1.58 MULT=1
MM1017 A_268_47# N_A_M1017_g N_A_130_417#_M1001_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75003.7 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g A_268_47# VNB NSHORT L=0.15 W=0.64 AD=0.255382
+ AS=0.0672 PD=1.57042 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75001.3
+ SB=75003.4 A=0.096 P=1.58 MULT=1
MM1005 A_534_47# N_A_130_417#_M1005_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.219468 PD=0.76 PS=1.34958 NRD=10.908 NRS=118.908 M=1 R=3.66667
+ SA=75002.3 SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1000 N_X_M1000_d N_A_130_417#_M1000_g A_534_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75002.7
+ SB=75002.6 A=0.0825 P=1.4 MULT=1
MM1002 N_X_M1000_d N_A_130_417#_M1002_g A_1008_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75003.1
+ SB=75002.1 A=0.0825 P=1.4 MULT=1
MM1016 A_1008_47# N_A_130_417#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75003.5
+ SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1010 A_692_47# N_A_130_417#_M1010_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75003.9
+ SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1006 N_X_M1006_d N_A_130_417#_M1006_g A_692_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75004.2
+ SB=75001 A=0.0825 P=1.4 MULT=1
MM1012 N_X_M1006_d N_A_130_417#_M1012_g A_850_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75004.7
+ SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1019 A_850_47# N_A_130_417#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75005
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_130_417#_M1007_s VPB PHIGHVT L=0.25 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125006
+ A=0.25 P=2.5 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_A_130_417#_M1007_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125005 A=0.25
+ P=2.5 MULT=1
MM1021 N_VPWR_M1015_d N_A_M1021_g N_A_130_417#_M1021_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125005 A=0.25
+ P=2.5 MULT=1
MM1022 N_VPWR_M1022_d N_A_M1022_g N_A_130_417#_M1021_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125004 A=0.25
+ P=2.5 MULT=1
MM1003 N_VPWR_M1022_d N_A_130_417#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125004 A=0.25
+ P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_130_417#_M1004_g N_X_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1008 N_VPWR_M1004_d N_A_130_417#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1013 N_VPWR_M1013_d N_A_130_417#_M1013_g N_X_M1008_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1014 N_VPWR_M1013_d N_A_130_417#_M1014_g N_X_M1014_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1018 N_VPWR_M1018_d N_A_130_417#_M1018_g N_X_M1014_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125005 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1020 N_VPWR_M1018_d N_A_130_417#_M1020_g N_X_M1020_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125005 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1023 N_VPWR_M1023_d N_A_130_417#_M1023_g N_X_M1020_s VPB PHIGHVT L=0.25 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125006 SB=125000
+ A=0.25 P=2.5 MULT=1
DX24_noxref VNB VPB NWDIODE A=14.1367 P=18.89
*
.include "sky130_fd_sc_lp__clkbuflp_8.pxi.spice"
*
.ends
*
*
