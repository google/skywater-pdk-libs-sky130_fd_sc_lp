* File: sky130_fd_sc_lp__o22ai_lp.pex.spice
* Created: Fri Aug 28 11:11:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22AI_LP%B1 3 9 10 11 12 15 17
r36 15 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.68 $Y=1.615
+ $X2=0.68 $Y2=1.78
r37 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.68 $Y=1.615
+ $X2=0.68 $Y2=1.45
r38 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.68
+ $Y=1.615 $X2=0.68 $Y2=1.615
r39 11 17 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=0.77 $Y=1.15 $X2=0.77
+ $Y2=1.45
r40 10 11 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=0.78 $Y=1 $X2=0.78
+ $Y2=1.15
r41 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.79 $Y=0.715 $X2=0.79
+ $Y2=1
r42 3 18 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=0.72 $Y=2.595
+ $X2=0.72 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_LP%B2 3 7 9 12
r37 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.615
+ $X2=1.25 $Y2=1.78
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.615
+ $X2=1.25 $Y2=1.45
r39 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.615 $X2=1.25 $Y2=1.615
r40 7 14 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.22 $Y=0.715
+ $X2=1.22 $Y2=1.45
r41 3 15 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=1.21 $Y=2.595
+ $X2=1.21 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_LP%A2 3 6 8 11 12 13
c36 11 0 1.64784e-19 $X=2.11 $Y=1.2
r37 11 14 63.2352 $w=6.2e-07 $l=5.05e-07 $layer=POLY_cond $X=1.965 $Y=1.2
+ $X2=1.965 $Y2=1.705
r38 11 13 50.0851 $w=6.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.965 $Y=1.2
+ $X2=1.965 $Y2=1.035
r39 11 12 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.11 $Y=1.2
+ $X2=2.11 $Y2=1.2
r40 8 12 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.11 $Y=1.295
+ $X2=2.11 $Y2=1.2
r41 6 14 221.124 $w=2.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.78 $Y=2.595
+ $X2=1.78 $Y2=1.705
r42 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.73 $Y=0.715
+ $X2=1.73 $Y2=1.035
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_LP%A1 3 6 9 10 11 12 15 16
r30 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.68 $Y=1.2
+ $X2=2.68 $Y2=1.2
r31 12 16 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.68 $Y=1.295
+ $X2=2.68 $Y2=1.2
r32 10 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.68 $Y=1.54
+ $X2=2.68 $Y2=1.2
r33 10 11 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.54
+ $X2=2.68 $Y2=1.705
r34 9 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.035
+ $X2=2.68 $Y2=1.2
r35 6 11 221.124 $w=2.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2.64 $Y=2.595
+ $X2=2.64 $Y2=1.705
r36 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.59 $Y=0.715 $X2=2.59
+ $Y2=1.035
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_LP%VPWR 1 2 9 13 16 17 18 19 20 21 34
r31 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r33 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 27 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 25 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 21 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 21 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 19 30 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.74 $Y=3.33 $X2=2.64
+ $Y2=3.33
r41 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.905 $Y2=3.33
r42 18 33 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=3.07 $Y=3.33 $X2=3.12
+ $Y2=3.33
r43 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=3.33
+ $X2=2.905 $Y2=3.33
r44 16 24 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=0.29 $Y=3.33 $X2=0.24
+ $Y2=3.33
r45 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.29 $Y=3.33
+ $X2=0.455 $Y2=3.33
r46 15 27 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.62 $Y=3.33 $X2=0.72
+ $Y2=3.33
r47 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.455 $Y2=3.33
r48 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=3.33
r49 11 13 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=2.4
r50 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.455 $Y=3.245
+ $X2=0.455 $Y2=3.33
r51 7 9 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.455 $Y=3.245
+ $X2=0.455 $Y2=2.475
r52 2 13 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=2.765
+ $Y=2.095 $X2=2.905 $Y2=2.4
r53 1 9 300 $w=1.7e-07 $l=4.46654e-07 $layer=licon1_PDIFF $count=2 $X=0.31
+ $Y=2.095 $X2=0.455 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_LP%Y 1 2 8 9 10 11 12 15 17 18
c45 9 0 1.64784e-19 $X=0.84 $Y=1.185
r46 17 18 9.52321 $w=4.74e-07 $l=3.7e-07 $layer=LI1_cond $X=1.362 $Y=2.405
+ $X2=1.362 $Y2=2.775
r47 17 23 0.128692 $w=4.74e-07 $l=5e-09 $layer=LI1_cond $X=1.362 $Y=2.405
+ $X2=1.362 $Y2=2.4
r48 13 15 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.005 $Y=1.1
+ $X2=1.005 $Y2=0.78
r49 11 23 9.13713 $w=4.74e-07 $l=4.73667e-07 $layer=LI1_cond $X=1.085 $Y=2.045
+ $X2=1.362 $Y2=2.4
r50 11 12 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.085 $Y=2.045
+ $X2=0.335 $Y2=2.045
r51 9 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.84 $Y=1.185
+ $X2=1.005 $Y2=1.1
r52 9 10 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.84 $Y=1.185
+ $X2=0.335 $Y2=1.185
r53 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.25 $Y=1.96
+ $X2=0.335 $Y2=2.045
r54 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.25 $Y=1.27
+ $X2=0.335 $Y2=1.185
r55 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.25 $Y=1.27 $X2=0.25
+ $Y2=1.96
r56 2 23 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=1.335
+ $Y=2.095 $X2=1.475 $Y2=2.4
r57 1 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.865
+ $Y=0.505 $X2=1.005 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_LP%A_70_101# 1 2 3 12 14 15 19 21 22 23 24 29
+ 30
r62 28 29 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.11 $Y=0.855
+ $X2=3.11 $Y2=1.885
r63 24 28 8.10976 $w=3.7e-07 $l=2.23495e-07 $layer=LI1_cond $X=3.025 $Y=0.67
+ $X2=3.11 $Y2=0.855
r64 24 26 6.85236 $w=3.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.025 $Y=0.67
+ $X2=2.805 $Y2=0.67
r65 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.025 $Y=1.97
+ $X2=3.11 $Y2=1.885
r66 22 23 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=3.025 $Y=1.97
+ $X2=1.765 $Y2=1.97
r67 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.68 $Y=1.885
+ $X2=1.765 $Y2=1.97
r68 21 30 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.68 $Y=1.885
+ $X2=1.68 $Y2=0.945
r69 17 30 9.87967 $w=4.13e-07 $l=2.07e-07 $layer=LI1_cond $X=1.557 $Y=0.738
+ $X2=1.557 $Y2=0.945
r70 17 19 0.638703 $w=4.13e-07 $l=2.3e-08 $layer=LI1_cond $X=1.557 $Y=0.738
+ $X2=1.557 $Y2=0.715
r71 16 19 7.77552 $w=4.13e-07 $l=2.8e-07 $layer=LI1_cond $X=1.557 $Y=0.435
+ $X2=1.557 $Y2=0.715
r72 14 16 8.50155 $w=1.7e-07 $l=2.45854e-07 $layer=LI1_cond $X=1.35 $Y=0.35
+ $X2=1.557 $Y2=0.435
r73 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.35 $Y=0.35 $X2=0.66
+ $Y2=0.35
r74 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.495 $Y=0.435
+ $X2=0.66 $Y2=0.35
r75 10 12 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.495 $Y=0.435
+ $X2=0.495 $Y2=0.7
r76 3 26 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.505 $X2=2.805 $Y2=0.67
r77 2 19 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=1.295
+ $Y=0.505 $X2=1.515 $Y2=0.715
r78 1 12 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.35
+ $Y=0.505 $X2=0.495 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_LP%VGND 1 6 8 10 20 21 24
r24 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r25 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r26 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r27 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.11
+ $Y2=0
r28 18 20 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=3.12
+ $Y2=0
r29 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r30 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r31 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.11
+ $Y2=0
r32 10 16 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.68
+ $Y2=0
r33 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r34 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r35 8 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r36 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0.085 $X2=2.11
+ $Y2=0
r37 4 6 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.67
r38 1 6 182 $w=1.7e-07 $l=3.78616e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.505 $X2=2.11 $Y2=0.67
.ends

