* File: sky130_fd_sc_lp__lsbufiso1p_lp.pxi.spice
* Created: Fri Aug 28 10:42:31 2020
* 
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%VGND N_VGND_M1014_s N_VGND_M1023_d
+ N_VGND_M1018_s N_VGND_M1012_s N_VGND_M1014_b N_VGND_c_12_p N_VGND_c_109_p
+ N_VGND_c_7_p N_VGND_c_76_p N_VGND_c_113_p VGND N_VGND_c_13_p N_VGND_c_95_p
+ N_VGND_c_77_p N_VGND_c_18_p N_VGND_c_8_p VGND
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%VGND
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%VPB N_VPB_M1011_b VPB VPB VPB VPB VPB VPB
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%VPB
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%DESTVPB N_DESTVPB_M1020_b DESTVPB DESTVPB
+ DESTVPB DESTVPB DESTVPB DESTVPB PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%DESTVPB
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_176_987# N_A_176_987#_M1022_d
+ N_A_176_987#_M1008_d N_A_176_987#_M1020_g N_A_176_987#_M1019_g
+ N_A_176_987#_c_260_n N_A_176_987#_c_253_n N_A_176_987#_c_262_n
+ N_A_176_987#_c_263_n N_A_176_987#_c_254_n N_A_176_987#_c_264_n
+ N_A_176_987#_c_257_n PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_176_987#
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A N_A_M1011_g N_A_c_331_n N_A_M1014_g
+ N_A_M1006_g N_A_c_340_n N_A_c_343_n N_A_M1004_g N_A_M1010_g N_A_c_349_n
+ N_A_M1000_g N_A_c_357_n N_A_c_359_n A N_A_c_363_n N_A_c_365_n
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_278_47# N_A_278_47#_M1010_d
+ N_A_278_47#_M1004_d N_A_278_47#_c_402_n N_A_278_47#_M1001_g
+ N_A_278_47#_c_404_n N_A_278_47#_c_407_n N_A_278_47#_c_410_n
+ N_A_278_47#_c_413_n N_A_278_47#_M1022_g N_A_278_47#_c_416_n
+ N_A_278_47#_c_429_n N_A_278_47#_c_419_n N_A_278_47#_c_422_n
+ N_A_278_47#_c_425_n N_A_278_47#_c_430_n N_A_278_47#_c_428_n
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_278_47#
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_123_718# N_A_123_718#_M1006_s
+ N_A_123_718#_M1020_s N_A_123_718#_c_492_n N_A_123_718#_M1007_g
+ N_A_123_718#_c_493_n N_A_123_718#_M1008_g N_A_123_718#_c_494_n
+ N_A_123_718#_c_473_n N_A_123_718#_M1017_g N_A_123_718#_M1009_g
+ N_A_123_718#_M1016_g N_A_123_718#_c_478_n N_A_123_718#_c_499_n
+ N_A_123_718#_c_481_n N_A_123_718#_c_482_n N_A_123_718#_c_501_n
+ N_A_123_718#_c_502_n N_A_123_718#_c_503_n N_A_123_718#_c_561_p
+ N_A_123_718#_c_504_n N_A_123_718#_c_483_n N_A_123_718#_c_484_n
+ N_A_123_718#_c_486_n N_A_123_718#_c_507_n N_A_123_718#_c_487_n
+ N_A_123_718#_c_510_n N_A_123_718#_c_488_n N_A_123_718#_c_489_n
+ N_A_123_718#_c_491_n PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_123_718#
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%SLEEP N_SLEEP_c_630_n N_SLEEP_M1018_g
+ N_SLEEP_M1015_g N_SLEEP_c_635_n N_SLEEP_M1013_g N_SLEEP_M1002_g
+ N_SLEEP_c_640_n N_SLEEP_c_641_n N_SLEEP_M1003_g SLEEP N_SLEEP_c_643_n
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%SLEEP
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_517_420# N_A_517_420#_M1013_d
+ N_A_517_420#_M1003_d N_A_517_420#_c_697_n N_A_517_420#_M1023_g
+ N_A_517_420#_c_700_n N_A_517_420#_c_705_n N_A_517_420#_c_709_n
+ N_A_517_420#_c_712_n N_A_517_420#_c_713_n N_A_517_420#_c_714_n
+ N_A_517_420#_M1021_g N_A_517_420#_c_716_n N_A_517_420#_M1005_g
+ N_A_517_420#_c_718_n N_A_517_420#_c_719_n N_A_517_420#_M1012_g
+ N_A_517_420#_c_723_n N_A_517_420#_c_724_n N_A_517_420#_c_726_n
+ N_A_517_420#_c_730_n N_A_517_420#_c_731_n N_A_517_420#_c_732_n
+ N_A_517_420#_c_733_n N_A_517_420#_c_736_n
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_517_420#
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%VPWR N_VPWR_M1011_s N_VPWR_c_797_n VPWR
+ N_VPWR_c_799_n N_VPWR_c_801_n N_VPWR_c_796_n N_VPWR_c_806_n VPWR
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%VPWR
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_278_1085# N_A_278_1085#_M1019_d
+ N_A_278_1085#_M1015_s N_A_278_1085#_c_827_n N_A_278_1085#_c_823_n
+ N_A_278_1085#_c_833_n N_A_278_1085#_c_824_n N_A_278_1085#_c_825_n
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_278_1085#
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%DESTPWR N_DESTPWR_M1015_d N_DESTPWR_M1005_d
+ N_DESTPWR_c_862_n N_DESTPWR_c_863_n N_DESTPWR_c_864_n N_DESTPWR_c_866_n
+ DESTPWR N_DESTPWR_c_867_n N_DESTPWR_c_868_n N_DESTPWR_c_861_n
+ N_DESTPWR_c_873_n DESTPWR PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%DESTPWR
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%X N_X_M1009_d N_X_M1021_s N_X_M1016_d
+ N_X_c_941_n N_X_c_942_n N_X_c_943_n X X X X X X X N_X_c_937_n X
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%X
x_PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_278_718# N_A_278_718#_M1000_d
+ N_A_278_718#_M1023_s N_A_278_718#_c_988_n N_A_278_718#_c_992_n
+ N_A_278_718#_c_993_n N_A_278_718#_c_999_n N_A_278_718#_c_1002_n
+ PM_SKY130_FD_SC_LP__LSBUFISO1P_LP%A_278_718#
cc_1 N_VGND_M1014_b VPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_2 N_VGND_M1014_b VPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=6.875 $Y2=0.47
cc_3 N_VGND_M1014_b DESTVPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_4 N_VGND_M1014_b DESTVPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=6.875 $Y2=0.47
cc_5 N_VGND_M1014_b N_A_176_987#_c_253_n 0.0155112f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_6 N_VGND_M1014_b N_A_176_987#_c_254_n 0.00431945f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_7 N_VGND_c_7_p N_A_176_987#_c_254_n 0.0120094f $X=2.865 $Y=4.155 $X2=0 $Y2=0
cc_8 N_VGND_c_8_p N_A_176_987#_c_254_n 0.00149965f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_9 N_VGND_M1014_b N_A_176_987#_c_257_n 0.0169579f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_10 N_VGND_M1014_b N_A_M1011_g 0.00622578f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_11 N_VGND_M1014_b N_A_c_331_n 0.0206818f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_12 N_VGND_c_12_p N_A_c_331_n 0.00818476f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_13 N_VGND_c_13_p N_A_c_331_n 9.22492e-19 $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_14 N_VGND_c_8_p N_A_c_331_n 7.18026e-19 $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_15 N_VGND_M1014_b N_A_M1006_g 0.0399099f $X=-0.025 $Y=-0.245 $X2=0.155
+ $Y2=0.84
cc_16 N_VGND_c_12_p N_A_M1006_g 0.00429861f $X=0.74 $Y=2.44 $X2=0.155 $Y2=0.84
cc_17 N_VGND_c_13_p N_A_M1006_g 0.00909137f $X=1.68 $Y=3.33 $X2=0.155 $Y2=0.84
cc_18 N_VGND_c_18_p N_A_M1006_g 0.00506743f $X=0.72 $Y=3.33 $X2=0.155 $Y2=0.84
cc_19 N_VGND_c_8_p N_A_M1006_g 0.0108583f $X=6.955 $Y=3.33 $X2=0.155 $Y2=0.84
cc_20 N_VGND_M1014_b N_A_c_340_n 0.0114117f $X=-0.025 $Y=-0.245 $X2=6.875
+ $Y2=0.47
cc_21 N_VGND_c_13_p N_A_c_340_n 5.14398e-19 $X=1.68 $Y=3.33 $X2=6.875 $Y2=0.47
cc_22 N_VGND_c_8_p N_A_c_340_n 0.00400159f $X=6.955 $Y=3.33 $X2=6.875 $Y2=0.47
cc_23 N_VGND_M1014_b N_A_c_343_n 0.00960464f $X=-0.025 $Y=-0.245 $X2=6.875
+ $Y2=0.84
cc_24 N_VGND_c_12_p N_A_c_343_n 0.00626201f $X=0.74 $Y=2.44 $X2=6.875 $Y2=0.84
cc_25 N_VGND_c_8_p N_A_c_343_n 0.00228999f $X=6.955 $Y=3.33 $X2=6.875 $Y2=0.84
cc_26 N_VGND_M1014_b N_A_M1004_g 0.00537455f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_27 N_VGND_M1014_b N_A_M1010_g 0.0097482f $X=-0.025 $Y=-0.245 $X2=0.24
+ $Y2=0.525
cc_28 N_VGND_c_12_p N_A_M1010_g 3.60856e-19 $X=0.74 $Y=2.44 $X2=0.24 $Y2=0.525
cc_29 N_VGND_M1014_b N_A_c_349_n 0.032122f $X=-0.025 $Y=-0.245 $X2=0.24
+ $Y2=0.525
cc_30 N_VGND_c_12_p N_A_c_349_n 5.98673e-19 $X=0.74 $Y=2.44 $X2=0.24 $Y2=0.525
cc_31 N_VGND_c_13_p N_A_c_349_n 0.0030635f $X=1.68 $Y=3.33 $X2=0.24 $Y2=0.525
cc_32 N_VGND_c_8_p N_A_c_349_n 0.00643718f $X=6.955 $Y=3.33 $X2=0.24 $Y2=0.525
cc_33 N_VGND_M1014_b N_A_M1000_g 0.029645f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_34 N_VGND_c_12_p N_A_M1000_g 8.81789e-19 $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_35 N_VGND_c_13_p N_A_M1000_g 0.0110813f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_36 N_VGND_c_8_p N_A_M1000_g 0.00964689f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_37 N_VGND_M1014_b N_A_c_357_n 0.00229529f $X=-0.025 $Y=-0.245 $X2=0.24
+ $Y2=1.295
cc_38 N_VGND_c_12_p N_A_c_357_n 0.0223008f $X=0.74 $Y=2.44 $X2=0.24 $Y2=1.295
cc_39 N_VGND_M1014_b N_A_c_359_n 0.00551809f $X=-0.025 $Y=-0.245 $X2=6.96
+ $Y2=0.525
cc_40 N_VGND_c_12_p N_A_c_359_n 0.0252639f $X=0.74 $Y=2.44 $X2=6.96 $Y2=0.525
cc_41 N_VGND_c_13_p N_A_c_359_n 0.0362016f $X=1.68 $Y=3.33 $X2=6.96 $Y2=0.525
cc_42 N_VGND_c_8_p N_A_c_359_n 0.0196655f $X=6.955 $Y=3.33 $X2=6.96 $Y2=0.525
cc_43 N_VGND_M1014_b N_A_c_363_n 0.0674831f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_44 N_VGND_c_12_p N_A_c_363_n 0.00213349f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_45 N_VGND_M1014_b N_A_c_365_n 0.0344278f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_46 N_VGND_c_12_p N_A_c_365_n 0.0262117f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_47 N_VGND_M1014_b N_A_278_47#_c_402_n 0.012966f $X=-0.025 $Y=-0.245
+ $X2=-0.025 $Y2=-0.19
cc_48 N_VGND_c_8_p N_A_278_47#_c_402_n 0.00222998f $X=6.955 $Y=3.33 $X2=-0.025
+ $Y2=-0.19
cc_49 N_VGND_M1014_b N_A_278_47#_c_404_n 0.00602992f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=0.84
cc_50 N_VGND_c_13_p N_A_278_47#_c_404_n 0.00312162f $X=1.68 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_51 N_VGND_c_8_p N_A_278_47#_c_404_n 2.63629e-19 $X=6.955 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_52 N_VGND_M1014_b N_A_278_47#_c_407_n 0.00857286f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=1.21
cc_53 N_VGND_c_13_p N_A_278_47#_c_407_n 0.00482701f $X=1.68 $Y=3.33 $X2=0.155
+ $Y2=1.21
cc_54 N_VGND_c_8_p N_A_278_47#_c_407_n 6.46318e-19 $X=6.955 $Y=3.33 $X2=0.155
+ $Y2=1.21
cc_55 N_VGND_M1014_b N_A_278_47#_c_410_n 0.0164815f $X=-0.025 $Y=-0.245
+ $X2=6.875 $Y2=0.84
cc_56 N_VGND_c_13_p N_A_278_47#_c_410_n 0.00507498f $X=1.68 $Y=3.33 $X2=6.875
+ $Y2=0.84
cc_57 N_VGND_c_8_p N_A_278_47#_c_410_n 0.00497945f $X=6.955 $Y=3.33 $X2=6.875
+ $Y2=0.84
cc_58 N_VGND_M1014_b N_A_278_47#_c_413_n 0.0162397f $X=-0.025 $Y=-0.245
+ $X2=6.875 $Y2=1.21
cc_59 N_VGND_c_7_p N_A_278_47#_c_413_n 0.00860948f $X=2.865 $Y=4.155 $X2=6.875
+ $Y2=1.21
cc_60 N_VGND_c_8_p N_A_278_47#_c_413_n 0.00271031f $X=6.955 $Y=3.33 $X2=6.875
+ $Y2=1.21
cc_61 N_VGND_M1014_b N_A_278_47#_c_416_n 0.00923091f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_62 N_VGND_c_13_p N_A_278_47#_c_416_n 0.00190461f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_63 N_VGND_c_8_p N_A_278_47#_c_416_n 0.00291644f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_64 N_VGND_M1014_b N_A_278_47#_c_419_n 0.0216596f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_65 N_VGND_c_13_p N_A_278_47#_c_419_n 0.00259986f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_66 N_VGND_c_8_p N_A_278_47#_c_419_n 0.00569686f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_67 N_VGND_M1014_b N_A_278_47#_c_422_n 0.00372993f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_68 N_VGND_c_13_p N_A_278_47#_c_422_n 0.0220216f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_69 N_VGND_c_8_p N_A_278_47#_c_422_n 0.012589f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_70 N_VGND_M1014_b N_A_278_47#_c_425_n 0.0371605f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_71 N_VGND_c_13_p N_A_278_47#_c_425_n 8.65569e-19 $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_72 N_VGND_c_8_p N_A_278_47#_c_425_n 0.00157003f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_73 N_VGND_M1014_b N_A_278_47#_c_428_n 0.0355797f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_74 N_VGND_M1014_b N_A_123_718#_c_473_n 0.0149084f $X=-0.025 $Y=-0.245
+ $X2=6.875 $Y2=1.21
cc_75 N_VGND_M1014_b N_A_123_718#_M1009_g 0.0472903f $X=-0.025 $Y=-0.245
+ $X2=0.24 $Y2=0.525
cc_76 N_VGND_c_76_p N_A_123_718#_M1009_g 0.00274215f $X=5.665 $Y=3.715 $X2=0.24
+ $Y2=0.525
cc_77 N_VGND_c_77_p N_A_123_718#_M1009_g 0.00525141f $X=6.81 $Y=3.33 $X2=0.24
+ $Y2=0.525
cc_78 N_VGND_c_8_p N_A_123_718#_M1009_g 0.0105621f $X=6.955 $Y=3.33 $X2=0.24
+ $Y2=0.525
cc_79 N_VGND_M1014_b N_A_123_718#_c_478_n 0.101989f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_80 N_VGND_c_18_p N_A_123_718#_c_478_n 0.0205041f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_81 N_VGND_c_8_p N_A_123_718#_c_478_n 0.0106717f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_82 N_VGND_M1014_b N_A_123_718#_c_481_n 0.0267048f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_83 N_VGND_M1014_b N_A_123_718#_c_482_n 0.00597888f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_84 N_VGND_M1014_b N_A_123_718#_c_483_n 0.00872825f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_85 N_VGND_M1014_b N_A_123_718#_c_484_n 0.0165559f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_86 N_VGND_c_76_p N_A_123_718#_c_484_n 0.0096556f $X=5.665 $Y=3.715 $X2=0
+ $Y2=0
cc_87 N_VGND_M1014_b N_A_123_718#_c_486_n 0.0152338f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_88 N_VGND_M1014_b N_A_123_718#_c_487_n 0.0119951f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_89 N_VGND_M1014_b N_A_123_718#_c_488_n 0.0063108f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_90 N_VGND_M1014_b N_A_123_718#_c_489_n 0.0150209f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_91 N_VGND_c_7_p N_A_123_718#_c_489_n 0.00116779f $X=2.865 $Y=4.155 $X2=0
+ $Y2=0
cc_92 N_VGND_M1014_b N_A_123_718#_c_491_n 0.0255523f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_93 N_VGND_M1014_b N_SLEEP_c_630_n 0.0164714f $X=-0.025 $Y=-0.245 $X2=0.155
+ $Y2=0.32
cc_94 N_VGND_c_7_p N_SLEEP_c_630_n 0.00923491f $X=2.865 $Y=4.155 $X2=0.155
+ $Y2=0.32
cc_95 N_VGND_c_95_p N_SLEEP_c_630_n 0.00153691f $X=5.5 $Y=3.33 $X2=0.155
+ $Y2=0.32
cc_96 N_VGND_c_8_p N_SLEEP_c_630_n 0.00245232f $X=6.955 $Y=3.33 $X2=0.155
+ $Y2=0.32
cc_97 N_VGND_M1014_b N_SLEEP_M1015_g 0.00647375f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_98 N_VGND_M1014_b N_SLEEP_c_635_n 0.0152475f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_99 N_VGND_c_7_p N_SLEEP_c_635_n 9.79299e-19 $X=2.865 $Y=4.155 $X2=0 $Y2=0
cc_100 N_VGND_c_95_p N_SLEEP_c_635_n 0.00171734f $X=5.5 $Y=3.33 $X2=0 $Y2=0
cc_101 N_VGND_c_8_p N_SLEEP_c_635_n 0.00243285f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_102 N_VGND_M1014_b N_SLEEP_M1002_g 0.00541457f $X=-0.025 $Y=-0.245 $X2=6.875
+ $Y2=0.84
cc_103 N_VGND_M1014_b N_SLEEP_c_640_n 0.0213497f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_104 N_VGND_M1014_b N_SLEEP_c_641_n 0.0425991f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_105 N_VGND_M1014_b N_SLEEP_M1003_g 0.0192696f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_106 N_VGND_M1014_b N_SLEEP_c_643_n 0.0119878f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_107 N_VGND_c_7_p N_SLEEP_c_643_n 0.0103371f $X=2.865 $Y=4.155 $X2=0 $Y2=0
cc_108 N_VGND_M1014_b N_A_517_420#_c_697_n 0.0273195f $X=-0.025 $Y=-0.245
+ $X2=-0.025 $Y2=-0.19
cc_109 N_VGND_c_109_p N_A_517_420#_c_697_n 0.0116122f $X=2.875 $Y=2.515
+ $X2=-0.025 $Y2=-0.19
cc_110 N_VGND_c_8_p N_A_517_420#_c_697_n 0.00596799f $X=6.955 $Y=3.33 $X2=-0.025
+ $Y2=-0.19
cc_111 N_VGND_M1014_b N_A_517_420#_c_700_n 0.0943772f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=0.84
cc_112 N_VGND_c_109_p N_A_517_420#_c_700_n 0.0124235f $X=2.875 $Y=2.515
+ $X2=0.155 $Y2=0.84
cc_113 N_VGND_c_113_p N_A_517_420#_c_700_n 0.00850832f $X=2.87 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_114 N_VGND_c_95_p N_A_517_420#_c_700_n 0.0351019f $X=5.5 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_115 N_VGND_c_8_p N_A_517_420#_c_700_n 0.0103238f $X=6.955 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_116 N_VGND_M1014_b N_A_517_420#_c_705_n 0.0101923f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=1.21
cc_117 N_VGND_c_109_p N_A_517_420#_c_705_n 8.23954e-19 $X=2.875 $Y=2.515
+ $X2=0.155 $Y2=1.21
cc_118 N_VGND_c_113_p N_A_517_420#_c_705_n 0.00129312f $X=2.87 $Y=3.33 $X2=0.155
+ $Y2=1.21
cc_119 N_VGND_c_8_p N_A_517_420#_c_705_n 0.00282686f $X=6.955 $Y=3.33 $X2=0.155
+ $Y2=1.21
cc_120 N_VGND_M1014_b N_A_517_420#_c_709_n 0.0467336f $X=-0.025 $Y=-0.245
+ $X2=6.875 $Y2=1.21
cc_121 N_VGND_c_95_p N_A_517_420#_c_709_n 0.0130561f $X=5.5 $Y=3.33 $X2=6.875
+ $Y2=1.21
cc_122 N_VGND_c_8_p N_A_517_420#_c_709_n 0.0140572f $X=6.955 $Y=3.33 $X2=6.875
+ $Y2=1.21
cc_123 N_VGND_M1014_b N_A_517_420#_c_712_n 0.0598505f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_124 N_VGND_M1014_b N_A_517_420#_c_713_n 0.0256106f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_125 N_VGND_M1014_b N_A_517_420#_c_714_n 0.0109051f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_126 N_VGND_M1014_b N_A_517_420#_M1021_g 0.0227467f $X=-0.025 $Y=-0.245
+ $X2=0.24 $Y2=0.525
cc_127 N_VGND_M1014_b N_A_517_420#_c_716_n 0.0152476f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_128 N_VGND_M1014_b N_A_517_420#_M1005_g 0.0173578f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_129 N_VGND_M1014_b N_A_517_420#_c_718_n 0.0231331f $X=-0.025 $Y=-0.245
+ $X2=6.96 $Y2=0.525
cc_130 N_VGND_M1014_b N_A_517_420#_c_719_n 0.0181137f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_131 N_VGND_c_76_p N_A_517_420#_c_719_n 0.017264f $X=5.665 $Y=3.715 $X2=0
+ $Y2=0
cc_132 N_VGND_c_77_p N_A_517_420#_c_719_n 0.00465098f $X=6.81 $Y=3.33 $X2=0
+ $Y2=0
cc_133 N_VGND_c_8_p N_A_517_420#_c_719_n 0.00803846f $X=6.955 $Y=3.33 $X2=0
+ $Y2=0
cc_134 N_VGND_M1014_b N_A_517_420#_c_723_n 0.0106787f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_135 N_VGND_M1014_b N_A_517_420#_c_724_n 0.0100249f $X=-0.025 $Y=-0.245
+ $X2=6.96 $Y2=1.295
cc_136 N_VGND_c_76_p N_A_517_420#_c_724_n 0.00506431f $X=5.665 $Y=3.715 $X2=6.96
+ $Y2=1.295
cc_137 N_VGND_M1014_b N_A_517_420#_c_726_n 0.019742f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_138 N_VGND_c_7_p N_A_517_420#_c_726_n 0.025063f $X=2.865 $Y=4.155 $X2=0 $Y2=0
cc_139 N_VGND_c_95_p N_A_517_420#_c_726_n 0.0400923f $X=5.5 $Y=3.33 $X2=0 $Y2=0
cc_140 N_VGND_c_8_p N_A_517_420#_c_726_n 0.0217427f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_141 N_VGND_M1014_b N_A_517_420#_c_730_n 0.0112138f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_142 N_VGND_M1014_b N_A_517_420#_c_731_n 0.0182874f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_143 N_VGND_M1014_b N_A_517_420#_c_732_n 0.00206795f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_144 N_VGND_M1014_b N_A_517_420#_c_733_n 0.0449483f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_145 N_VGND_c_95_p N_A_517_420#_c_733_n 0.00336816f $X=5.5 $Y=3.33 $X2=0 $Y2=0
cc_146 N_VGND_c_8_p N_A_517_420#_c_733_n 0.00254324f $X=6.955 $Y=3.33 $X2=0
+ $Y2=0
cc_147 N_VGND_M1014_b N_A_517_420#_c_736_n 0.0233371f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_148 N_VGND_c_95_p N_A_517_420#_c_736_n 0.00847838f $X=5.5 $Y=3.33 $X2=0 $Y2=0
cc_149 N_VGND_c_8_p N_A_517_420#_c_736_n 0.00641058f $X=6.955 $Y=3.33 $X2=0
+ $Y2=0
cc_150 N_VGND_M1014_b N_VPWR_c_796_n 0.302998f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_151 N_VGND_M1014_b N_DESTPWR_c_861_n 0.302998f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_152 N_VGND_M1014_b N_X_c_937_n 0.116044f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_153 N_VGND_c_76_p N_X_c_937_n 0.02158f $X=5.665 $Y=3.715 $X2=0 $Y2=0
cc_154 N_VGND_c_77_p N_X_c_937_n 0.0234355f $X=6.81 $Y=3.33 $X2=0 $Y2=0
cc_155 N_VGND_c_8_p N_X_c_937_n 0.0124904f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_156 N_VGND_M1014_b N_A_278_718#_c_988_n 0.00481358f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=0.47
cc_157 N_VGND_c_7_p N_A_278_718#_c_988_n 0.0127465f $X=2.865 $Y=4.155 $X2=0.155
+ $Y2=0.47
cc_158 N_VGND_c_13_p N_A_278_718#_c_988_n 0.03008f $X=1.68 $Y=3.33 $X2=0.155
+ $Y2=0.47
cc_159 N_VGND_c_8_p N_A_278_718#_c_988_n 0.0273016f $X=6.955 $Y=3.33 $X2=0.155
+ $Y2=0.47
cc_160 N_VGND_M1014_b N_A_278_718#_c_992_n 0.00602893f $X=-0.025 $Y=-0.245
+ $X2=6.875 $Y2=0.84
cc_161 N_VGND_M1014_b N_A_278_718#_c_993_n 0.00951612f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_162 N_VGND_c_109_p N_A_278_718#_c_993_n 0.00818712f $X=2.875 $Y=2.515 $X2=0
+ $Y2=0
cc_163 N_VGND_c_7_p N_A_278_718#_c_993_n 0.00977302f $X=2.865 $Y=4.155 $X2=0
+ $Y2=0
cc_164 N_VGND_c_113_p N_A_278_718#_c_993_n 0.009578f $X=2.87 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VGND_c_13_p N_A_278_718#_c_993_n 0.0115155f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_166 N_VGND_c_8_p N_A_278_718#_c_993_n 0.0299272f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_167 N_VGND_M1014_b N_A_278_718#_c_999_n 0.00440914f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_168 N_VGND_c_13_p N_A_278_718#_c_999_n 0.0199194f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_169 N_VGND_c_8_p N_A_278_718#_c_999_n 0.0106419f $X=6.955 $Y=3.33 $X2=0 $Y2=0
cc_170 N_VGND_M1014_b N_A_278_718#_c_1002_n 0.00150655f $X=-0.025 $Y=-0.245
+ $X2=0 $Y2=0
cc_171 N_VGND_c_109_p N_A_278_718#_c_1002_n 0.0254913f $X=2.875 $Y=2.515 $X2=0
+ $Y2=0
cc_172 N_VGND_c_8_p N_A_278_718#_c_1002_n 0.0150136f $X=6.955 $Y=3.33 $X2=0
+ $Y2=0
cc_173 N_VPB_M1011_b N_A_M1011_g 0.0389027f $X=-0.025 $Y=-0.19 $X2=2.74 $Y2=4.01
cc_174 VPB N_A_M1011_g 0.00621856f $X=0.155 $Y=0.47 $X2=2.74 $Y2=4.01
cc_175 N_VPB_M1011_b N_A_M1004_g 0.0358449f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_176 N_VPB_M1011_b N_A_c_365_n 0.0183257f $X=-0.025 $Y=-0.19 $X2=2.865
+ $Y2=3.415
cc_177 N_VPB_M1011_b N_A_278_47#_c_429_n 0.0369401f $X=-0.025 $Y=-0.19 $X2=0
+ $Y2=0
cc_178 N_VPB_M1011_b N_A_278_47#_c_430_n 0.00836222f $X=-0.025 $Y=-0.19 $X2=0.24
+ $Y2=3.245
cc_179 N_VPB_M1011_b N_A_278_47#_c_428_n 0.0164461f $X=-0.025 $Y=-0.19 $X2=0
+ $Y2=0
cc_180 N_VPB_M1011_b N_VPWR_c_797_n 0.0144492f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_797_n 0.0708842f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_182 N_VPB_M1011_b N_VPWR_c_799_n 0.0176917f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_799_n 0.0200925f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_184 N_VPB_M1011_b N_VPWR_c_801_n 0.195456f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_801_n 0.0200925f $X=6.875 $Y=0.47 $X2=0 $Y2=0
cc_186 N_VPB_M1011_b N_VPWR_c_796_n 0.269451f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_796_n 0.0115306f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_796_n 0.0115306f $X=6.875 $Y=0.47 $X2=0 $Y2=0
cc_189 N_VPB_M1011_b N_VPWR_c_806_n 0.00513431f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_190 N_DESTVPB_M1020_b N_A_176_987#_M1020_g 0.0210833f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_191 N_DESTVPB_M1020_b N_A_176_987#_M1019_g 0.0170453f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_192 N_DESTVPB_M1020_b N_A_176_987#_c_260_n 0.00720677f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_193 N_DESTVPB_M1020_b N_A_176_987#_c_253_n 0.00300753f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_194 N_DESTVPB_M1020_b N_A_176_987#_c_262_n 0.00470784f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_195 N_DESTVPB_M1020_b N_A_176_987#_c_263_n 0.00229064f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_196 N_DESTVPB_M1020_b N_A_176_987#_c_264_n 0.00192288f $X=-0.025 $Y=4.985
+ $X2=0.24 $Y2=3.245
cc_197 N_DESTVPB_M1020_b N_A_176_987#_c_257_n 0.0274464f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_198 N_DESTVPB_M1020_b N_A_123_718#_c_492_n 0.0130622f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_199 N_DESTVPB_M1020_b N_A_123_718#_c_493_n 0.0167244f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_200 N_DESTVPB_M1020_b N_A_123_718#_c_494_n 0.0141652f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_201 N_DESTVPB_M1020_b N_A_123_718#_c_473_n 0.0331088f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_202 N_DESTVPB_M1020_b N_A_123_718#_M1017_g 0.0212279f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_203 N_DESTVPB_M1020_b N_A_123_718#_M1016_g 0.0261663f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_204 DESTVPB N_A_123_718#_M1016_g 0.00227698f $X=6.875 $Y=5.28 $X2=0 $Y2=0
cc_205 N_DESTVPB_M1020_b N_A_123_718#_c_499_n 0.00931091f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_206 N_DESTVPB_M1020_b N_A_123_718#_c_482_n 3.94425e-19 $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_207 N_DESTVPB_M1020_b N_A_123_718#_c_501_n 0.0188543f $X=-0.025 $Y=4.985
+ $X2=0.575 $Y2=3.33
cc_208 N_DESTVPB_M1020_b N_A_123_718#_c_502_n 0.00125038f $X=-0.025 $Y=4.985
+ $X2=0.74 $Y2=2.44
cc_209 N_DESTVPB_M1020_b N_A_123_718#_c_503_n 0.00887275f $X=-0.025 $Y=4.985
+ $X2=0.74 $Y2=2.44
cc_210 N_DESTVPB_M1020_b N_A_123_718#_c_504_n 0.0230839f $X=-0.025 $Y=4.985
+ $X2=2.87 $Y2=2.515
cc_211 N_DESTVPB_M1020_b N_A_123_718#_c_483_n 0.00281474f $X=-0.025 $Y=4.985
+ $X2=2.875 $Y2=2.515
cc_212 N_DESTVPB_M1020_b N_A_123_718#_c_484_n 0.0178612f $X=-0.025 $Y=4.985
+ $X2=2.865 $Y2=3.415
cc_213 N_DESTVPB_M1020_b N_A_123_718#_c_507_n 0.00192794f $X=-0.025 $Y=4.985
+ $X2=5.665 $Y2=3.715
cc_214 N_DESTVPB_M1020_b N_A_123_718#_c_487_n 0.0165636f $X=-0.025 $Y=4.985
+ $X2=5.665 $Y2=3.715
cc_215 DESTVPB N_A_123_718#_c_487_n 0.0914628f $X=0.155 $Y=5.28 $X2=5.665
+ $Y2=3.715
cc_216 N_DESTVPB_M1020_b N_A_123_718#_c_510_n 0.00338836f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_217 N_DESTVPB_M1020_b N_A_123_718#_c_489_n 0.0375662f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_218 N_DESTVPB_M1020_b N_A_123_718#_c_491_n 0.0208973f $X=-0.025 $Y=4.985
+ $X2=3.12 $Y2=3.33
cc_219 N_DESTVPB_M1020_b N_SLEEP_M1015_g 0.035012f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_220 N_DESTVPB_M1020_b N_SLEEP_M1002_g 0.0295144f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_221 N_DESTVPB_M1020_b N_SLEEP_M1003_g 0.0340418f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_222 N_DESTVPB_M1020_b N_A_517_420#_M1021_g 0.0376072f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_223 N_DESTVPB_M1020_b N_A_517_420#_M1005_g 0.0295558f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_224 N_DESTVPB_M1020_b N_A_517_420#_c_732_n 0.00941765f $X=-0.025 $Y=4.985
+ $X2=0.575 $Y2=3.33
cc_225 N_DESTVPB_M1020_b N_A_278_1085#_c_823_n 0.0106837f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_226 N_DESTVPB_M1020_b N_A_278_1085#_c_824_n 4.74859e-19 $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_227 N_DESTVPB_M1020_b N_A_278_1085#_c_825_n 0.00837059f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_228 N_DESTVPB_M1020_b N_DESTPWR_c_862_n 0.0047158f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_229 N_DESTVPB_M1020_b N_DESTPWR_c_863_n 4.89148e-19 $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_230 N_DESTVPB_M1020_b N_DESTPWR_c_864_n 0.0819886f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_231 DESTVPB N_DESTPWR_c_864_n 0.0200925f $X=0.155 $Y=5.28 $X2=0 $Y2=0
cc_232 N_DESTVPB_M1020_b N_DESTPWR_c_866_n 0.00324402f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_233 N_DESTVPB_M1020_b N_DESTPWR_c_867_n 0.0546587f $X=-0.025 $Y=4.985
+ $X2=-0.025 $Y2=-0.245
cc_234 N_DESTVPB_M1020_b N_DESTPWR_c_868_n 0.0387302f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_235 DESTVPB N_DESTPWR_c_868_n 0.0200925f $X=6.875 $Y=5.28 $X2=0 $Y2=0
cc_236 N_DESTVPB_M1020_b N_DESTPWR_c_861_n 0.0793456f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_237 DESTVPB N_DESTPWR_c_861_n 0.0115306f $X=0.155 $Y=5.28 $X2=0 $Y2=0
cc_238 DESTVPB N_DESTPWR_c_861_n 0.0115306f $X=6.875 $Y=5.28 $X2=0 $Y2=0
cc_239 N_DESTVPB_M1020_b N_DESTPWR_c_873_n 0.00436868f $X=-0.025 $Y=4.985
+ $X2=0.39 $Y2=3.33
cc_240 N_DESTVPB_M1020_b N_X_c_941_n 0.00499003f $X=-0.025 $Y=4.985 $X2=0 $Y2=0
cc_241 N_DESTVPB_M1020_b N_X_c_942_n 0.00863934f $X=-0.025 $Y=4.985 $X2=0 $Y2=0
cc_242 N_DESTVPB_M1020_b N_X_c_943_n 0.00924941f $X=-0.025 $Y=4.985 $X2=0 $Y2=0
cc_243 N_DESTVPB_M1020_b X 0.00192634f $X=-0.025 $Y=4.985 $X2=0 $Y2=0
cc_244 DESTVPB X 0.0138061f $X=6.875 $Y=5.28 $X2=0 $Y2=0
cc_245 N_DESTVPB_M1020_b X 0.00959313f $X=-0.025 $Y=4.985 $X2=0 $Y2=0
cc_246 DESTVPB X 0.0615054f $X=6.875 $Y=5.28 $X2=0 $Y2=0
cc_247 N_DESTVPB_M1020_b N_X_c_937_n 0.0126699f $X=-0.025 $Y=4.985 $X2=0 $Y2=0
cc_248 DESTVPB N_X_c_937_n 0.0152519f $X=6.875 $Y=5.28 $X2=0 $Y2=0
cc_249 N_A_176_987#_c_257_n N_A_M1006_g 0.00436304f $X=1.315 $Y=5.1 $X2=0 $Y2=0
cc_250 N_A_176_987#_c_257_n N_A_M1000_g 0.00436304f $X=1.315 $Y=5.1 $X2=0 $Y2=0
cc_251 N_A_176_987#_c_254_n N_A_278_47#_c_402_n 0.00155306f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_252 N_A_176_987#_c_253_n N_A_278_47#_c_413_n 0.00534252f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_253 N_A_176_987#_c_254_n N_A_278_47#_c_413_n 0.00599326f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_254 N_A_176_987#_c_260_n N_A_123_718#_c_492_n 0.0137915f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_255 N_A_176_987#_c_262_n N_A_123_718#_c_492_n 0.00182938f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_256 N_A_176_987#_c_260_n N_A_123_718#_c_493_n 0.0137481f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_257 N_A_176_987#_c_262_n N_A_123_718#_c_493_n 0.00899114f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_258 N_A_176_987#_c_264_n N_A_123_718#_c_493_n 0.0015814f $X=2.155 $Y=5.355
+ $X2=0 $Y2=0
cc_259 N_A_176_987#_c_253_n N_A_123_718#_c_494_n 0.0113062f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_260 N_A_176_987#_c_264_n N_A_123_718#_c_494_n 0.00779865f $X=2.155 $Y=5.355
+ $X2=0 $Y2=0
cc_261 N_A_176_987#_M1019_g N_A_123_718#_c_473_n 0.0275551f $X=1.315 $Y=5.925
+ $X2=0 $Y2=0
cc_262 N_A_176_987#_c_260_n N_A_123_718#_c_473_n 0.00279508f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_263 N_A_176_987#_c_253_n N_A_123_718#_c_473_n 0.00893677f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_264 N_A_176_987#_c_263_n N_A_123_718#_c_473_n 0.00130944f $X=1.165 $Y=5.1
+ $X2=0 $Y2=0
cc_265 N_A_176_987#_c_257_n N_A_123_718#_c_473_n 0.0219836f $X=1.315 $Y=5.1
+ $X2=0 $Y2=0
cc_266 N_A_176_987#_M1020_g N_A_123_718#_c_499_n 0.0139667f $X=0.955 $Y=5.925
+ $X2=0 $Y2=0
cc_267 N_A_176_987#_c_260_n N_A_123_718#_c_481_n 0.00619807f $X=2.155 $Y=5.44
+ $X2=0.24 $Y2=3.855
cc_268 N_A_176_987#_c_253_n N_A_123_718#_c_481_n 0.00714341f $X=2.24 $Y=5.355
+ $X2=0.24 $Y2=3.855
cc_269 N_A_176_987#_c_263_n N_A_123_718#_c_481_n 0.0252464f $X=1.165 $Y=5.1
+ $X2=0.24 $Y2=3.855
cc_270 N_A_176_987#_c_257_n N_A_123_718#_c_481_n 0.0102483f $X=1.315 $Y=5.1
+ $X2=0.24 $Y2=3.855
cc_271 N_A_176_987#_c_253_n N_A_123_718#_c_482_n 0.00682589f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_272 N_A_176_987#_c_263_n N_A_123_718#_c_482_n 0.00138846f $X=1.165 $Y=5.1
+ $X2=0 $Y2=0
cc_273 N_A_176_987#_c_257_n N_A_123_718#_c_482_n 0.00132465f $X=1.315 $Y=5.1
+ $X2=0 $Y2=0
cc_274 N_A_176_987#_M1020_g N_A_123_718#_c_507_n 0.00381798f $X=0.955 $Y=5.925
+ $X2=5.665 $Y2=3.715
cc_275 N_A_176_987#_M1019_g N_A_123_718#_c_507_n 0.00296352f $X=1.315 $Y=5.925
+ $X2=5.665 $Y2=3.715
cc_276 N_A_176_987#_c_263_n N_A_123_718#_c_507_n 0.00581585f $X=1.165 $Y=5.1
+ $X2=5.665 $Y2=3.715
cc_277 N_A_176_987#_c_263_n N_A_123_718#_c_487_n 0.0299155f $X=1.165 $Y=5.1
+ $X2=5.665 $Y2=3.715
cc_278 N_A_176_987#_c_257_n N_A_123_718#_c_487_n 0.0143834f $X=1.315 $Y=5.1
+ $X2=5.665 $Y2=3.715
cc_279 N_A_176_987#_c_260_n N_A_123_718#_c_510_n 0.0290917f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_280 N_A_176_987#_c_253_n N_A_123_718#_c_510_n 0.0107546f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_281 N_A_176_987#_c_263_n N_A_123_718#_c_510_n 0.0129286f $X=1.165 $Y=5.1
+ $X2=0 $Y2=0
cc_282 N_A_176_987#_c_257_n N_A_123_718#_c_510_n 0.00119275f $X=1.315 $Y=5.1
+ $X2=0 $Y2=0
cc_283 N_A_176_987#_c_253_n N_A_123_718#_c_488_n 0.0247133f $X=2.24 $Y=5.355
+ $X2=6.96 $Y2=3.855
cc_284 N_A_176_987#_c_253_n N_A_123_718#_c_489_n 0.00266561f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_285 N_A_176_987#_c_254_n N_A_123_718#_c_489_n 0.00195932f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_286 N_A_176_987#_c_253_n N_SLEEP_c_630_n 0.00210636f $X=2.24 $Y=5.355
+ $X2=0.615 $Y2=2.23
cc_287 N_A_176_987#_c_254_n N_SLEEP_c_630_n 0.00282641f $X=2.32 $Y=4.235
+ $X2=0.615 $Y2=2.23
cc_288 N_A_176_987#_c_253_n N_SLEEP_M1015_g 8.14403e-19 $X=2.24 $Y=5.355 $X2=0
+ $Y2=0
cc_289 N_A_176_987#_c_264_n N_SLEEP_M1015_g 0.00227452f $X=2.155 $Y=5.355 $X2=0
+ $Y2=0
cc_290 N_A_176_987#_c_253_n N_SLEEP_c_641_n 0.00165252f $X=2.24 $Y=5.355 $X2=0
+ $Y2=0
cc_291 N_A_176_987#_c_253_n N_SLEEP_c_643_n 0.0156705f $X=2.24 $Y=5.355 $X2=0
+ $Y2=0
cc_292 N_A_176_987#_c_263_n A_206_1085# 0.00200208f $X=1.165 $Y=5.1 $X2=0.615
+ $Y2=2.23
cc_293 N_A_176_987#_c_260_n N_A_278_1085#_M1019_d 0.00176461f $X=2.155 $Y=5.44
+ $X2=0.615 $Y2=2.23
cc_294 N_A_176_987#_M1020_g N_A_278_1085#_c_827_n 0.00145208f $X=0.955 $Y=5.925
+ $X2=0 $Y2=0
cc_295 N_A_176_987#_M1019_g N_A_278_1085#_c_827_n 0.0102531f $X=1.315 $Y=5.925
+ $X2=0 $Y2=0
cc_296 N_A_176_987#_c_260_n N_A_278_1085#_c_827_n 0.0171383f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_297 N_A_176_987#_c_262_n N_A_278_1085#_c_827_n 0.0120446f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_298 N_A_176_987#_M1008_d N_A_278_1085#_c_823_n 0.00559995f $X=2.18 $Y=5.425
+ $X2=0 $Y2=0
cc_299 N_A_176_987#_c_262_n N_A_278_1085#_c_823_n 0.019416f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_300 N_A_176_987#_M1020_g N_A_278_1085#_c_833_n 4.5542e-19 $X=0.955 $Y=5.925
+ $X2=0 $Y2=0
cc_301 N_A_176_987#_M1019_g N_A_278_1085#_c_833_n 0.00285177f $X=1.315 $Y=5.925
+ $X2=0 $Y2=0
cc_302 N_A_176_987#_c_262_n N_A_278_1085#_c_825_n 0.0374058f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_303 N_A_176_987#_c_264_n N_A_278_1085#_c_825_n 0.00449869f $X=2.155 $Y=5.355
+ $X2=0 $Y2=0
cc_304 N_A_176_987#_c_260_n A_364_1085# 0.00366293f $X=2.155 $Y=5.44 $X2=0.615
+ $Y2=2.23
cc_305 N_A_176_987#_M1020_g N_DESTPWR_c_864_n 0.00518588f $X=0.955 $Y=5.925
+ $X2=0 $Y2=0
cc_306 N_A_176_987#_M1019_g N_DESTPWR_c_864_n 0.00547432f $X=1.315 $Y=5.925
+ $X2=0 $Y2=0
cc_307 N_A_176_987#_M1008_d N_DESTPWR_c_861_n 0.00232737f $X=2.18 $Y=5.425 $X2=0
+ $Y2=0
cc_308 N_A_176_987#_M1020_g N_DESTPWR_c_861_n 0.0103683f $X=0.955 $Y=5.925 $X2=0
+ $Y2=0
cc_309 N_A_176_987#_M1019_g N_DESTPWR_c_861_n 0.00979813f $X=1.315 $Y=5.925
+ $X2=0 $Y2=0
cc_310 N_A_176_987#_M1022_d N_A_278_718#_c_988_n 0.00426626f $X=2.18 $Y=3.59
+ $X2=0 $Y2=0
cc_311 N_A_176_987#_c_254_n N_A_278_718#_c_988_n 0.0126536f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_312 N_A_176_987#_c_254_n N_A_278_718#_c_999_n 0.00705761f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_313 N_A_M1000_g N_A_278_47#_c_407_n 0.0237825f $X=1.315 $Y=4.01 $X2=0 $Y2=0
cc_314 N_A_c_349_n N_A_278_47#_c_410_n 0.00454236f $X=1.315 $Y=3.14 $X2=0 $Y2=0
cc_315 N_A_M1011_g N_A_278_47#_c_429_n 0.00339963f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_316 N_A_M1004_g N_A_278_47#_c_429_n 0.0148505f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_317 N_A_c_349_n N_A_278_47#_c_419_n 0.00346449f $X=1.315 $Y=3.14 $X2=0 $Y2=0
cc_318 N_A_c_359_n N_A_278_47#_c_419_n 0.0154334f $X=1.405 $Y=2.925 $X2=0 $Y2=0
cc_319 N_A_M1010_g N_A_278_47#_c_422_n 0.00232378f $X=1.315 $Y=2.44 $X2=0 $Y2=0
cc_320 N_A_c_349_n N_A_278_47#_c_422_n 3.97765e-19 $X=1.315 $Y=3.14 $X2=0 $Y2=0
cc_321 N_A_c_357_n N_A_278_47#_c_422_n 0.00510196f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_322 N_A_c_359_n N_A_278_47#_c_422_n 0.0247675f $X=1.405 $Y=2.925 $X2=0 $Y2=0
cc_323 N_A_c_349_n N_A_278_47#_c_425_n 0.0171629f $X=1.315 $Y=3.14 $X2=-0.025
+ $Y2=-0.245
cc_324 N_A_c_359_n N_A_278_47#_c_425_n 0.00191938f $X=1.405 $Y=2.925 $X2=-0.025
+ $Y2=-0.245
cc_325 N_A_M1004_g N_A_278_47#_c_430_n 0.00684213f $X=1.315 $Y=0.735 $X2=0.24
+ $Y2=3.245
cc_326 N_A_M1004_g N_A_278_47#_c_428_n 0.0272488f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_327 N_A_c_357_n N_A_278_47#_c_428_n 0.0140219f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_328 N_A_c_365_n N_A_278_47#_c_428_n 0.0500336f $X=1.16 $Y=1.832 $X2=0 $Y2=0
cc_329 N_A_M1006_g N_A_123_718#_c_478_n 0.00781951f $X=0.955 $Y=4.01 $X2=-0.025
+ $Y2=-0.245
cc_330 N_A_M1006_g N_A_123_718#_c_481_n 0.00392017f $X=0.955 $Y=4.01 $X2=0.24
+ $Y2=3.855
cc_331 N_A_M1000_g N_A_123_718#_c_481_n 0.00352781f $X=1.315 $Y=4.01 $X2=0.24
+ $Y2=3.855
cc_332 N_A_M1011_g N_VPWR_c_797_n 0.0213886f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_333 N_A_M1004_g N_VPWR_c_797_n 0.00375886f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_334 N_A_c_363_n N_VPWR_c_797_n 0.00119966f $X=1.315 $Y=1.96 $X2=0 $Y2=0
cc_335 N_A_c_365_n N_VPWR_c_797_n 0.0154497f $X=1.16 $Y=1.832 $X2=0 $Y2=0
cc_336 N_A_M1011_g N_VPWR_c_801_n 0.00486043f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_337 N_A_M1004_g N_VPWR_c_801_n 0.00549284f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_338 N_A_M1011_g N_VPWR_c_796_n 0.00814425f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_339 N_A_M1004_g N_VPWR_c_796_n 0.0111098f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_340 N_A_M1006_g N_A_278_718#_c_999_n 0.00250397f $X=0.955 $Y=4.01 $X2=0 $Y2=0
cc_341 N_A_M1000_g N_A_278_718#_c_999_n 0.0175796f $X=1.315 $Y=4.01 $X2=0 $Y2=0
cc_342 N_A_278_47#_c_402_n N_A_123_718#_c_473_n 0.006115f $X=1.745 $Y=3.515
+ $X2=0 $Y2=0
cc_343 N_A_278_47#_c_413_n N_A_123_718#_c_473_n 0.00407187f $X=2.105 $Y=3.515
+ $X2=0 $Y2=0
cc_344 N_A_278_47#_c_402_n N_A_123_718#_c_481_n 5.99168e-19 $X=1.745 $Y=3.515
+ $X2=0.24 $Y2=3.855
cc_345 N_A_278_47#_c_402_n N_A_123_718#_c_510_n 8.15435e-19 $X=1.745 $Y=3.515
+ $X2=0 $Y2=0
cc_346 N_A_278_47#_c_413_n N_SLEEP_c_643_n 2.77866e-19 $X=2.105 $Y=3.515 $X2=0
+ $Y2=0
cc_347 N_A_278_47#_c_425_n N_A_517_420#_c_697_n 0.00490025f $X=1.98 $Y=2.925
+ $X2=0 $Y2=0
cc_348 N_A_278_47#_c_410_n N_A_517_420#_c_705_n 0.00490025f $X=2.07 $Y=3.365
+ $X2=0 $Y2=0
cc_349 N_A_278_47#_c_429_n N_VPWR_c_797_n 0.0305839f $X=1.53 $Y=0.38 $X2=0 $Y2=0
cc_350 N_A_278_47#_c_429_n N_VPWR_c_801_n 0.0211337f $X=1.53 $Y=0.38 $X2=0 $Y2=0
cc_351 N_A_278_47#_M1004_d N_VPWR_c_796_n 0.00215406f $X=1.39 $Y=0.235 $X2=0
+ $Y2=0
cc_352 N_A_278_47#_c_429_n N_VPWR_c_796_n 0.0132819f $X=1.53 $Y=0.38 $X2=0 $Y2=0
cc_353 N_A_278_47#_c_402_n N_A_278_718#_c_988_n 0.012303f $X=1.745 $Y=3.515
+ $X2=0 $Y2=0
cc_354 N_A_278_47#_c_404_n N_A_278_718#_c_988_n 5.62214e-19 $X=1.995 $Y=3.44
+ $X2=0 $Y2=0
cc_355 N_A_278_47#_c_413_n N_A_278_718#_c_988_n 0.0151615f $X=2.105 $Y=3.515
+ $X2=0 $Y2=0
cc_356 N_A_278_47#_c_419_n N_A_278_718#_c_992_n 0.0144198f $X=1.98 $Y=2.605
+ $X2=0 $Y2=0
cc_357 N_A_278_47#_c_422_n N_A_278_718#_c_992_n 0.036567f $X=1.98 $Y=2.925 $X2=0
+ $Y2=0
cc_358 N_A_278_47#_c_425_n N_A_278_718#_c_992_n 0.00279589f $X=1.98 $Y=2.925
+ $X2=0 $Y2=0
cc_359 N_A_278_47#_c_428_n N_A_278_718#_c_992_n 0.00349796f $X=1.53 $Y=2.44
+ $X2=0 $Y2=0
cc_360 N_A_278_47#_c_410_n N_A_278_718#_c_993_n 6.18037e-19 $X=2.07 $Y=3.365
+ $X2=0 $Y2=0
cc_361 N_A_278_47#_c_416_n N_A_278_718#_c_993_n 0.00617354f $X=2.087 $Y=3.44
+ $X2=0 $Y2=0
cc_362 N_A_278_47#_c_402_n N_A_278_718#_c_999_n 0.00138154f $X=1.745 $Y=3.515
+ $X2=0 $Y2=0
cc_363 N_A_278_47#_c_410_n N_A_278_718#_c_1002_n 0.00279589f $X=2.07 $Y=3.365
+ $X2=0 $Y2=0
cc_364 N_A_123_718#_c_501_n N_SLEEP_M1015_g 0.0156186f $X=3.63 $Y=5.182 $X2=0
+ $Y2=0
cc_365 N_A_123_718#_c_488_n N_SLEEP_M1015_g 8.95485e-19 $X=2.58 $Y=5.1 $X2=0
+ $Y2=0
cc_366 N_A_123_718#_c_489_n N_SLEEP_M1015_g 0.0216008f $X=2.58 $Y=5.1 $X2=0
+ $Y2=0
cc_367 N_A_123_718#_c_501_n N_SLEEP_M1002_g 0.0205619f $X=3.63 $Y=5.182 $X2=0
+ $Y2=0
cc_368 N_A_123_718#_c_502_n N_SLEEP_M1002_g 0.00589813f $X=3.715 $Y=6.235 $X2=0
+ $Y2=0
cc_369 N_A_123_718#_c_501_n N_SLEEP_c_641_n 6.5474e-19 $X=3.63 $Y=5.182 $X2=0
+ $Y2=0
cc_370 N_A_123_718#_c_501_n N_SLEEP_M1003_g 0.00387019f $X=3.63 $Y=5.182 $X2=0
+ $Y2=0
cc_371 N_A_123_718#_c_502_n N_SLEEP_M1003_g 0.0161684f $X=3.715 $Y=6.235 $X2=0
+ $Y2=0
cc_372 N_A_123_718#_c_503_n N_SLEEP_M1003_g 0.0137631f $X=4.34 $Y=6.32 $X2=0
+ $Y2=0
cc_373 N_A_123_718#_c_561_p N_SLEEP_M1003_g 0.00114517f $X=3.8 $Y=6.32 $X2=0
+ $Y2=0
cc_374 N_A_123_718#_c_504_n N_SLEEP_M1003_g 0.00396339f $X=4.427 $Y=6.235 $X2=0
+ $Y2=0
cc_375 N_A_123_718#_c_483_n N_SLEEP_M1003_g 8.11573e-19 $X=4.515 $Y=5.03 $X2=0
+ $Y2=0
cc_376 N_A_123_718#_c_501_n N_SLEEP_c_643_n 0.0465697f $X=3.63 $Y=5.182 $X2=0
+ $Y2=0
cc_377 N_A_123_718#_c_503_n N_A_517_420#_M1003_d 0.00726325f $X=4.34 $Y=6.32
+ $X2=2.735 $Y2=2.23
cc_378 N_A_123_718#_c_484_n N_A_517_420#_c_714_n 0.01922f $X=5.97 $Y=5.03 $X2=0
+ $Y2=0
cc_379 N_A_123_718#_c_504_n N_A_517_420#_M1021_g 0.00657811f $X=4.427 $Y=6.235
+ $X2=0 $Y2=0
cc_380 N_A_123_718#_c_484_n N_A_517_420#_M1021_g 0.024411f $X=5.97 $Y=5.03 $X2=0
+ $Y2=0
cc_381 N_A_123_718#_c_484_n N_A_517_420#_c_716_n 0.00106595f $X=5.97 $Y=5.03
+ $X2=0 $Y2=0
cc_382 N_A_123_718#_M1009_g N_A_517_420#_M1005_g 0.00495086f $X=6.24 $Y=4.01
+ $X2=0 $Y2=0
cc_383 N_A_123_718#_c_484_n N_A_517_420#_M1005_g 0.0199892f $X=5.97 $Y=5.03
+ $X2=0 $Y2=0
cc_384 N_A_123_718#_c_491_n N_A_517_420#_M1005_g 0.0470057f $X=6.24 $Y=5.03
+ $X2=0 $Y2=0
cc_385 N_A_123_718#_c_484_n N_A_517_420#_c_718_n 0.00827873f $X=5.97 $Y=5.03
+ $X2=0 $Y2=0
cc_386 N_A_123_718#_c_491_n N_A_517_420#_c_718_n 0.0113492f $X=6.24 $Y=5.03
+ $X2=0 $Y2=0
cc_387 N_A_123_718#_M1009_g N_A_517_420#_c_719_n 0.0721639f $X=6.24 $Y=4.01
+ $X2=0.24 $Y2=2.39
cc_388 N_A_123_718#_c_501_n N_A_517_420#_c_731_n 0.0173336f $X=3.63 $Y=5.182
+ $X2=0 $Y2=0
cc_389 N_A_123_718#_c_483_n N_A_517_420#_c_731_n 0.00407387f $X=4.515 $Y=5.03
+ $X2=0 $Y2=0
cc_390 N_A_123_718#_c_501_n N_A_517_420#_c_732_n 0.0165741f $X=3.63 $Y=5.182
+ $X2=0.575 $Y2=3.33
cc_391 N_A_123_718#_c_502_n N_A_517_420#_c_732_n 0.0314219f $X=3.715 $Y=6.235
+ $X2=0.575 $Y2=3.33
cc_392 N_A_123_718#_c_503_n N_A_517_420#_c_732_n 0.0121011f $X=4.34 $Y=6.32
+ $X2=0.575 $Y2=3.33
cc_393 N_A_123_718#_c_504_n N_A_517_420#_c_732_n 0.064803f $X=4.427 $Y=6.235
+ $X2=0.575 $Y2=3.33
cc_394 N_A_123_718#_c_483_n N_A_517_420#_c_732_n 0.02434f $X=4.515 $Y=5.03
+ $X2=0.575 $Y2=3.33
cc_395 N_A_123_718#_c_492_n N_A_278_1085#_c_827_n 0.0106887f $X=1.745 $Y=5.35
+ $X2=0 $Y2=0
cc_396 N_A_123_718#_c_493_n N_A_278_1085#_c_827_n 0.00187953f $X=2.105 $Y=5.35
+ $X2=0 $Y2=0
cc_397 N_A_123_718#_c_499_n N_A_278_1085#_c_827_n 0.0188335f $X=0.74 $Y=6.28
+ $X2=0 $Y2=0
cc_398 N_A_123_718#_c_492_n N_A_278_1085#_c_823_n 0.010046f $X=1.745 $Y=5.35
+ $X2=0 $Y2=0
cc_399 N_A_123_718#_c_493_n N_A_278_1085#_c_823_n 0.0151541f $X=2.105 $Y=5.35
+ $X2=0 $Y2=0
cc_400 N_A_123_718#_c_492_n N_A_278_1085#_c_833_n 5.81207e-19 $X=1.745 $Y=5.35
+ $X2=0 $Y2=0
cc_401 N_A_123_718#_c_499_n N_A_278_1085#_c_833_n 0.00629328f $X=0.74 $Y=6.28
+ $X2=0 $Y2=0
cc_402 N_A_123_718#_c_493_n N_A_278_1085#_c_825_n 0.00426399f $X=2.105 $Y=5.35
+ $X2=0 $Y2=0
cc_403 N_A_123_718#_c_501_n N_A_278_1085#_c_825_n 0.0235948f $X=3.63 $Y=5.182
+ $X2=0 $Y2=0
cc_404 N_A_123_718#_c_489_n N_A_278_1085#_c_825_n 0.00115449f $X=2.58 $Y=5.1
+ $X2=0 $Y2=0
cc_405 N_A_123_718#_c_501_n N_DESTPWR_c_862_n 0.0139854f $X=3.63 $Y=5.182 $X2=0
+ $Y2=0
cc_406 N_A_123_718#_M1017_g N_DESTPWR_c_863_n 0.0157312f $X=5.88 $Y=5.925 $X2=0
+ $Y2=0
cc_407 N_A_123_718#_M1016_g N_DESTPWR_c_863_n 0.00298741f $X=6.24 $Y=5.925 $X2=0
+ $Y2=0
cc_408 N_A_123_718#_c_492_n N_DESTPWR_c_864_n 0.00357842f $X=1.745 $Y=5.35 $X2=0
+ $Y2=0
cc_409 N_A_123_718#_c_493_n N_DESTPWR_c_864_n 0.00357877f $X=2.105 $Y=5.35 $X2=0
+ $Y2=0
cc_410 N_A_123_718#_c_499_n N_DESTPWR_c_864_n 0.0224101f $X=0.74 $Y=6.28 $X2=0
+ $Y2=0
cc_411 N_A_123_718#_c_503_n N_DESTPWR_c_867_n 0.0449568f $X=4.34 $Y=6.32
+ $X2=-0.025 $Y2=-0.245
cc_412 N_A_123_718#_c_561_p N_DESTPWR_c_867_n 0.00953907f $X=3.8 $Y=6.32
+ $X2=-0.025 $Y2=-0.245
cc_413 N_A_123_718#_M1017_g N_DESTPWR_c_868_n 0.00486043f $X=5.88 $Y=5.925 $X2=0
+ $Y2=0
cc_414 N_A_123_718#_M1016_g N_DESTPWR_c_868_n 0.0054895f $X=6.24 $Y=5.925 $X2=0
+ $Y2=0
cc_415 N_A_123_718#_M1020_s N_DESTPWR_c_861_n 0.00215158f $X=0.615 $Y=5.425
+ $X2=0 $Y2=0
cc_416 N_A_123_718#_c_492_n N_DESTPWR_c_861_n 0.00516571f $X=1.745 $Y=5.35 $X2=0
+ $Y2=0
cc_417 N_A_123_718#_c_493_n N_DESTPWR_c_861_n 0.0066108f $X=2.105 $Y=5.35 $X2=0
+ $Y2=0
cc_418 N_A_123_718#_M1017_g N_DESTPWR_c_861_n 0.00814425f $X=5.88 $Y=5.925 $X2=0
+ $Y2=0
cc_419 N_A_123_718#_M1016_g N_DESTPWR_c_861_n 0.0111095f $X=6.24 $Y=5.925 $X2=0
+ $Y2=0
cc_420 N_A_123_718#_c_499_n N_DESTPWR_c_861_n 0.0132444f $X=0.74 $Y=6.28 $X2=0
+ $Y2=0
cc_421 N_A_123_718#_c_503_n N_DESTPWR_c_861_n 0.0264391f $X=4.34 $Y=6.32 $X2=0
+ $Y2=0
cc_422 N_A_123_718#_c_561_p N_DESTPWR_c_861_n 0.00658105f $X=3.8 $Y=6.32 $X2=0
+ $Y2=0
cc_423 N_A_123_718#_c_561_p A_717_1085# 9.38685e-19 $X=3.8 $Y=6.32 $X2=0.615
+ $Y2=2.23
cc_424 N_A_123_718#_c_504_n N_X_c_941_n 0.0130569f $X=4.427 $Y=6.235 $X2=0 $Y2=0
cc_425 N_A_123_718#_c_484_n N_X_c_941_n 0.0237492f $X=5.97 $Y=5.03 $X2=0 $Y2=0
cc_426 N_A_123_718#_c_503_n N_X_c_942_n 0.0136484f $X=4.34 $Y=6.32 $X2=0 $Y2=0
cc_427 N_A_123_718#_c_504_n N_X_c_942_n 0.0464642f $X=4.427 $Y=6.235 $X2=0 $Y2=0
cc_428 N_A_123_718#_M1017_g N_X_c_943_n 0.0140575f $X=5.88 $Y=5.925 $X2=0 $Y2=0
cc_429 N_A_123_718#_M1016_g N_X_c_943_n 0.0144352f $X=6.24 $Y=5.925 $X2=0 $Y2=0
cc_430 N_A_123_718#_c_484_n N_X_c_943_n 0.0622623f $X=5.97 $Y=5.03 $X2=0 $Y2=0
cc_431 N_A_123_718#_c_491_n N_X_c_943_n 9.24294e-19 $X=6.24 $Y=5.03 $X2=0 $Y2=0
cc_432 N_A_123_718#_M1016_g X 3.84662e-19 $X=6.24 $Y=5.925 $X2=0 $Y2=0
cc_433 N_A_123_718#_M1017_g X 0.0026051f $X=5.88 $Y=5.925 $X2=0 $Y2=0
cc_434 N_A_123_718#_M1016_g X 0.0133868f $X=6.24 $Y=5.925 $X2=0 $Y2=0
cc_435 N_A_123_718#_M1017_g N_X_c_937_n 0.00112036f $X=5.88 $Y=5.925 $X2=0 $Y2=0
cc_436 N_A_123_718#_M1009_g N_X_c_937_n 0.0388936f $X=6.24 $Y=4.01 $X2=0 $Y2=0
cc_437 N_A_123_718#_M1016_g N_X_c_937_n 0.00837854f $X=6.24 $Y=5.925 $X2=0 $Y2=0
cc_438 N_A_123_718#_c_484_n N_X_c_937_n 0.0201866f $X=5.97 $Y=5.03 $X2=0 $Y2=0
cc_439 N_A_123_718#_c_491_n N_X_c_937_n 0.0128845f $X=6.24 $Y=5.03 $X2=0 $Y2=0
cc_440 N_A_123_718#_c_478_n N_A_278_718#_c_999_n 0.0147015f $X=0.74 $Y=3.75
+ $X2=0 $Y2=0
cc_441 N_A_123_718#_c_481_n N_A_278_718#_c_999_n 0.0239528f $X=1.52 $Y=4.735
+ $X2=0 $Y2=0
cc_442 N_SLEEP_c_630_n N_A_517_420#_c_700_n 0.0024026f $X=3.08 $Y=4.505 $X2=0
+ $Y2=0
cc_443 N_SLEEP_c_635_n N_A_517_420#_c_700_n 0.00239275f $X=3.44 $Y=4.505 $X2=0
+ $Y2=0
cc_444 N_SLEEP_c_640_n N_A_517_420#_c_714_n 0.00499312f $X=3.795 $Y=4.58 $X2=0
+ $Y2=0
cc_445 N_SLEEP_c_630_n N_A_517_420#_c_726_n 9.80946e-19 $X=3.08 $Y=4.505
+ $X2=0.24 $Y2=3.855
cc_446 N_SLEEP_c_635_n N_A_517_420#_c_726_n 0.00974027f $X=3.44 $Y=4.505
+ $X2=0.24 $Y2=3.855
cc_447 N_SLEEP_c_640_n N_A_517_420#_c_726_n 0.00115892f $X=3.795 $Y=4.58
+ $X2=0.24 $Y2=3.855
cc_448 N_SLEEP_c_641_n N_A_517_420#_c_726_n 0.00200184f $X=3.585 $Y=4.58
+ $X2=0.24 $Y2=3.855
cc_449 N_SLEEP_c_635_n N_A_517_420#_c_730_n 0.00830112f $X=3.44 $Y=4.505 $X2=0
+ $Y2=0
cc_450 N_SLEEP_c_640_n N_A_517_420#_c_730_n 0.0171351f $X=3.795 $Y=4.58 $X2=0
+ $Y2=0
cc_451 N_SLEEP_c_641_n N_A_517_420#_c_730_n 6.97724e-19 $X=3.585 $Y=4.58 $X2=0
+ $Y2=0
cc_452 N_SLEEP_M1003_g N_A_517_420#_c_730_n 0.00409965f $X=3.87 $Y=5.925 $X2=0
+ $Y2=0
cc_453 N_SLEEP_c_643_n N_A_517_420#_c_730_n 0.0182819f $X=3.255 $Y=4.705 $X2=0
+ $Y2=0
cc_454 N_SLEEP_c_640_n N_A_517_420#_c_731_n 2.17082e-19 $X=3.795 $Y=4.58 $X2=0
+ $Y2=0
cc_455 N_SLEEP_c_641_n N_A_517_420#_c_731_n 0.00145826f $X=3.585 $Y=4.58 $X2=0
+ $Y2=0
cc_456 N_SLEEP_M1003_g N_A_517_420#_c_731_n 0.0182564f $X=3.87 $Y=5.925 $X2=0
+ $Y2=0
cc_457 N_SLEEP_c_643_n N_A_517_420#_c_731_n 0.0148003f $X=3.255 $Y=4.705 $X2=0
+ $Y2=0
cc_458 N_SLEEP_M1003_g N_A_517_420#_c_732_n 0.0148374f $X=3.87 $Y=5.925
+ $X2=0.575 $Y2=3.33
cc_459 N_SLEEP_c_635_n N_A_517_420#_c_733_n 0.00136449f $X=3.44 $Y=4.505
+ $X2=0.74 $Y2=2.44
cc_460 N_SLEEP_c_640_n N_A_517_420#_c_733_n 0.00195107f $X=3.795 $Y=4.58
+ $X2=0.74 $Y2=2.44
cc_461 N_SLEEP_M1015_g N_A_278_1085#_c_824_n 0.00196162f $X=3.08 $Y=5.925 $X2=0
+ $Y2=0
cc_462 N_SLEEP_M1015_g N_A_278_1085#_c_825_n 0.00829071f $X=3.08 $Y=5.925 $X2=0
+ $Y2=0
cc_463 N_SLEEP_M1015_g N_DESTPWR_c_862_n 0.00271808f $X=3.08 $Y=5.925 $X2=0
+ $Y2=0
cc_464 N_SLEEP_M1002_g N_DESTPWR_c_862_n 0.00271808f $X=3.51 $Y=5.925 $X2=0
+ $Y2=0
cc_465 N_SLEEP_M1015_g N_DESTPWR_c_864_n 0.00547432f $X=3.08 $Y=5.925 $X2=0
+ $Y2=0
cc_466 N_SLEEP_M1002_g N_DESTPWR_c_867_n 0.00585385f $X=3.51 $Y=5.925 $X2=-0.025
+ $Y2=-0.245
cc_467 N_SLEEP_M1003_g N_DESTPWR_c_867_n 0.0035787f $X=3.87 $Y=5.925 $X2=-0.025
+ $Y2=-0.245
cc_468 N_SLEEP_M1015_g N_DESTPWR_c_861_n 0.0110556f $X=3.08 $Y=5.925 $X2=0 $Y2=0
cc_469 N_SLEEP_M1002_g N_DESTPWR_c_861_n 0.0105424f $X=3.51 $Y=5.925 $X2=0 $Y2=0
cc_470 N_SLEEP_M1003_g N_DESTPWR_c_861_n 0.00661079f $X=3.87 $Y=5.925 $X2=0
+ $Y2=0
cc_471 N_A_517_420#_M1021_g N_DESTPWR_c_863_n 0.00298741f $X=5.09 $Y=5.925 $X2=0
+ $Y2=0
cc_472 N_A_517_420#_M1005_g N_DESTPWR_c_863_n 0.0157312f $X=5.45 $Y=5.925 $X2=0
+ $Y2=0
cc_473 N_A_517_420#_M1021_g N_DESTPWR_c_867_n 0.0054895f $X=5.09 $Y=5.925
+ $X2=-0.025 $Y2=-0.245
cc_474 N_A_517_420#_M1005_g N_DESTPWR_c_867_n 0.00486043f $X=5.45 $Y=5.925
+ $X2=-0.025 $Y2=-0.245
cc_475 N_A_517_420#_M1003_d N_DESTPWR_c_861_n 0.00232737f $X=3.945 $Y=5.425
+ $X2=0 $Y2=0
cc_476 N_A_517_420#_M1021_g N_DESTPWR_c_861_n 0.0111095f $X=5.09 $Y=5.925 $X2=0
+ $Y2=0
cc_477 N_A_517_420#_M1005_g N_DESTPWR_c_861_n 0.00814425f $X=5.45 $Y=5.925 $X2=0
+ $Y2=0
cc_478 N_A_517_420#_M1021_g N_X_c_941_n 8.0539e-19 $X=5.09 $Y=5.925 $X2=0 $Y2=0
cc_479 N_A_517_420#_M1021_g N_X_c_942_n 0.0133868f $X=5.09 $Y=5.925 $X2=0 $Y2=0
cc_480 N_A_517_420#_M1005_g N_X_c_942_n 0.0026051f $X=5.45 $Y=5.925 $X2=0 $Y2=0
cc_481 N_A_517_420#_M1021_g N_X_c_943_n 0.0109191f $X=5.09 $Y=5.925 $X2=0 $Y2=0
cc_482 N_A_517_420#_M1005_g N_X_c_943_n 0.0140575f $X=5.45 $Y=5.925 $X2=0 $Y2=0
cc_483 N_A_517_420#_c_719_n N_X_c_937_n 0.00400661f $X=5.88 $Y=4.505 $X2=0 $Y2=0
cc_484 N_A_517_420#_c_697_n N_A_278_718#_c_993_n 0.00164072f $X=2.66 $Y=3.145
+ $X2=0 $Y2=0
cc_485 N_A_517_420#_c_697_n N_A_278_718#_c_1002_n 9.25134e-19 $X=2.66 $Y=3.145
+ $X2=0 $Y2=0
cc_486 N_VPWR_c_796_n A_206_47# 0.00899413f $X=6.96 $Y=0 $X2=0.615 $Y2=2.23
cc_487 A_206_1085# N_DESTPWR_c_861_n 0.00899413f $X=1.03 $Y=5.425 $X2=0 $Y2=0
cc_488 N_A_278_1085#_c_823_n A_364_1085# 0.00456442f $X=2.7 $Y=6.32 $X2=0.155
+ $Y2=5.495
cc_489 N_A_278_1085#_c_823_n N_DESTPWR_c_864_n 0.0585658f $X=2.7 $Y=6.32 $X2=0
+ $Y2=0
cc_490 N_A_278_1085#_c_833_n N_DESTPWR_c_864_n 0.019107f $X=1.695 $Y=6.32 $X2=0
+ $Y2=0
cc_491 N_A_278_1085#_c_824_n N_DESTPWR_c_864_n 0.021147f $X=2.865 $Y=6.235 $X2=0
+ $Y2=0
cc_492 N_A_278_1085#_M1019_d N_DESTPWR_c_861_n 0.00223559f $X=1.39 $Y=5.425
+ $X2=0 $Y2=0
cc_493 N_A_278_1085#_M1015_s N_DESTPWR_c_861_n 0.00219347f $X=2.735 $Y=5.425
+ $X2=0 $Y2=0
cc_494 N_A_278_1085#_c_823_n N_DESTPWR_c_861_n 0.0365269f $X=2.7 $Y=6.32 $X2=0
+ $Y2=0
cc_495 N_A_278_1085#_c_833_n N_DESTPWR_c_861_n 0.0124689f $X=1.695 $Y=6.32 $X2=0
+ $Y2=0
cc_496 N_A_278_1085#_c_824_n N_DESTPWR_c_861_n 0.0126374f $X=2.865 $Y=6.235
+ $X2=0 $Y2=0
cc_497 A_364_1085# N_DESTPWR_c_861_n 0.00168889f $X=1.82 $Y=5.425 $X2=0 $Y2=0
cc_498 N_DESTPWR_c_861_n A_717_1085# 0.00325419f $X=6.96 $Y=6.66 $X2=0.615
+ $Y2=2.23
cc_499 N_DESTPWR_c_861_n N_X_M1021_s 0.00231914f $X=6.96 $Y=6.66 $X2=2.735
+ $Y2=2.23
cc_500 N_DESTPWR_c_861_n N_X_M1016_d 0.00215158f $X=6.96 $Y=6.66 $X2=2.74
+ $Y2=4.01
cc_501 N_DESTPWR_c_863_n N_X_c_942_n 0.02158f $X=5.665 $Y=5.925 $X2=0 $Y2=0
cc_502 N_DESTPWR_c_867_n N_X_c_942_n 0.0210192f $X=5.5 $Y=6.66 $X2=0 $Y2=0
cc_503 N_DESTPWR_c_861_n N_X_c_942_n 0.0125689f $X=6.96 $Y=6.66 $X2=0 $Y2=0
cc_504 N_DESTPWR_M1005_d N_X_c_943_n 0.00176461f $X=5.525 $Y=5.425 $X2=0 $Y2=0
cc_505 N_DESTPWR_c_863_n N_X_c_943_n 0.0170777f $X=5.665 $Y=5.925 $X2=0 $Y2=0
cc_506 N_DESTPWR_c_863_n X 0.02158f $X=5.665 $Y=5.925 $X2=0 $Y2=0
cc_507 N_DESTPWR_c_868_n X 0.0210467f $X=6.96 $Y=6.66 $X2=0 $Y2=0
cc_508 N_DESTPWR_c_861_n X 0.0125689f $X=6.96 $Y=6.66 $X2=0 $Y2=0
cc_509 N_DESTPWR_c_861_n A_1033_1085# 0.00899413f $X=6.96 $Y=6.66 $X2=0.615
+ $Y2=2.23
cc_510 N_DESTPWR_c_861_n A_1191_1085# 0.00899413f $X=6.96 $Y=6.66 $X2=0.615
+ $Y2=2.23
cc_511 N_X_c_943_n A_1033_1085# 0.00366293f $X=6.29 $Y=5.505 $X2=0.615 $Y2=2.23
cc_512 N_X_c_943_n A_1191_1085# 0.00366293f $X=6.29 $Y=5.505 $X2=0.615 $Y2=2.23
cc_513 N_A_278_718#_c_988_n A_364_718# 0.00366293f $X=2.315 $Y=3.67 $X2=0.615
+ $Y2=2.23
