* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__lsbufiso0p_lp A DESTPWR DESTVPB SLEEP VGND VPB VPWR X
X0 a_206_1085# a_176_987# a_278_1085# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A a_206_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_123_718# a_176_987# a_206_1085# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_1096_1085# a_123_718# X DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_123_718# a_1096_718# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_278_718# a_517_420# VGND VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 DESTPWR SLEEP a_1096_1085# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_206_718# A a_278_718# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_364_718# a_278_47# a_176_987# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_278_1085# SLEEP DESTPWR DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_206_446# A a_278_47# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_123_718# A a_206_718# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_278_718# a_278_47# a_364_718# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_206_47# A a_278_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND A a_206_446# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 DESTPWR SLEEP a_789_1085# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND SLEEP a_631_802# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_364_1085# a_123_718# a_176_987# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_938_718# SLEEP VGND VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_278_1085# a_123_718# a_364_1085# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 X SLEEP a_938_718# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_1096_718# a_123_718# X VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_631_802# SLEEP a_517_420# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_789_1085# SLEEP a_517_420# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
