* File: sky130_fd_sc_lp__nand2_0.pxi.spice
* Created: Wed Sep  2 10:02:28 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2_0%B N_B_c_31_n N_B_M1000_g N_B_M1003_g N_B_c_34_n B
+ B B B N_B_c_36_n PM_SKY130_FD_SC_LP__NAND2_0%B
x_PM_SKY130_FD_SC_LP__NAND2_0%A N_A_M1001_g N_A_c_65_n N_A_M1002_g N_A_c_67_n A
+ A A A N_A_c_69_n PM_SKY130_FD_SC_LP__NAND2_0%A
x_PM_SKY130_FD_SC_LP__NAND2_0%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_c_92_n
+ N_VPWR_c_93_n N_VPWR_c_94_n N_VPWR_c_95_n VPWR N_VPWR_c_96_n N_VPWR_c_91_n
+ PM_SKY130_FD_SC_LP__NAND2_0%VPWR
x_PM_SKY130_FD_SC_LP__NAND2_0%Y N_Y_M1001_d N_Y_M1000_d N_Y_c_112_n Y Y Y Y Y Y
+ Y N_Y_c_121_n PM_SKY130_FD_SC_LP__NAND2_0%Y
x_PM_SKY130_FD_SC_LP__NAND2_0%VGND N_VGND_M1003_s N_VGND_c_137_n N_VGND_c_138_n
+ VGND N_VGND_c_139_n N_VGND_c_140_n PM_SKY130_FD_SC_LP__NAND2_0%VGND
cc_1 VNB N_B_c_31_n 0.0202004f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.293
cc_2 VNB N_B_M1000_g 0.0091255f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.63
cc_3 VNB N_B_M1003_g 0.0268657f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_4 VNB N_B_c_34_n 0.0275627f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.51
cc_5 VNB B 0.0348786f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_B_c_36_n 0.0272544f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.005
cc_7 VNB N_A_M1001_g 0.0279297f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.51
cc_8 VNB N_A_c_65_n 0.0253344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_M1002_g 0.00912628f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_10 VNB N_A_c_67_n 0.0225363f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.51
cc_11 VNB A 0.0346214f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_12 VNB N_A_c_69_n 0.0225363f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.005
cc_13 VNB N_VPWR_c_91_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.005
cc_14 VNB N_Y_c_112_n 0.0146291f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_15 VNB Y 0.00746953f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.51
cc_16 VNB N_VGND_c_137_n 0.0126323f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.63
cc_17 VNB N_VGND_c_138_n 0.0195287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_139_n 0.0277722f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_19 VNB N_VGND_c_140_n 0.108843f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VPB N_B_M1000_g 0.0566387f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.63
cc_21 VPB B 0.0245417f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_22 VPB N_A_M1002_g 0.0568021f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.445
cc_23 VPB A 0.0246608f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_24 VPB N_VPWR_c_92_n 0.0120225f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.84
cc_25 VPB N_VPWR_c_93_n 0.0380505f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.445
cc_26 VPB N_VPWR_c_94_n 0.0123961f $X=-0.19 $Y=1.655 $X2=0.402 $Y2=1.51
cc_27 VPB N_VPWR_c_95_n 0.0382776f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_28 VPB N_VPWR_c_96_n 0.0156608f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_91_n 0.0548521f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.005
cc_30 VPB Y 0.0153505f $X=-0.19 $Y=1.655 $X2=0.402 $Y2=1.51
cc_31 N_B_M1003_g N_A_M1001_g 0.018627f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_32 N_B_c_31_n N_A_c_65_n 0.018627f $X=0.402 $Y=1.293 $X2=0 $Y2=0
cc_33 N_B_M1000_g N_A_M1002_g 0.0330237f $X=0.505 $Y=2.63 $X2=0 $Y2=0
cc_34 N_B_c_34_n N_A_c_67_n 0.018627f $X=0.402 $Y=1.51 $X2=0 $Y2=0
cc_35 N_B_c_36_n A 4.96749e-19 $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_36 N_B_c_36_n N_A_c_69_n 0.018627f $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_37 N_B_M1000_g N_VPWR_c_93_n 0.0107396f $X=0.505 $Y=2.63 $X2=0 $Y2=0
cc_38 B N_VPWR_c_93_n 0.0288227f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_39 N_B_M1000_g N_VPWR_c_95_n 5.189e-19 $X=0.505 $Y=2.63 $X2=0 $Y2=0
cc_40 N_B_M1000_g N_VPWR_c_96_n 0.00550536f $X=0.505 $Y=2.63 $X2=0 $Y2=0
cc_41 N_B_M1000_g N_VPWR_c_91_n 0.005282f $X=0.505 $Y=2.63 $X2=0 $Y2=0
cc_42 N_B_c_31_n Y 0.00528529f $X=0.402 $Y=1.293 $X2=0 $Y2=0
cc_43 N_B_M1000_g Y 0.00931179f $X=0.505 $Y=2.63 $X2=0 $Y2=0
cc_44 N_B_M1003_g Y 0.0109331f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_45 N_B_c_34_n Y 0.00525324f $X=0.402 $Y=1.51 $X2=0 $Y2=0
cc_46 B Y 0.0954349f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_47 N_B_c_36_n Y 0.00490132f $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_48 N_B_M1003_g N_Y_c_121_n 0.00680023f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_49 N_B_M1003_g N_VGND_c_138_n 0.00495318f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_50 B N_VGND_c_138_n 0.0170081f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_51 N_B_c_36_n N_VGND_c_138_n 0.00179982f $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_52 N_B_M1003_g N_VGND_c_139_n 0.00563132f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_53 N_B_M1003_g N_VGND_c_140_n 0.0112381f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_54 B N_VGND_c_140_n 0.00417553f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_55 N_B_c_36_n N_VGND_c_140_n 8.97026e-19 $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_56 N_A_M1002_g N_VPWR_c_93_n 4.96635e-19 $X=0.935 $Y=2.63 $X2=0 $Y2=0
cc_57 N_A_M1002_g N_VPWR_c_95_n 0.0126707f $X=0.935 $Y=2.63 $X2=0 $Y2=0
cc_58 A N_VPWR_c_95_n 0.0305157f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_59 N_A_M1002_g N_VPWR_c_96_n 0.0047441f $X=0.935 $Y=2.63 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_VPWR_c_91_n 0.00455844f $X=0.935 $Y=2.63 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_Y_c_112_n 0.0157886f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_62 A N_Y_c_112_n 0.0187654f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_63 N_A_c_69_n N_Y_c_112_n 0.00139689f $X=1.07 $Y=1.005 $X2=0 $Y2=0
cc_64 N_A_M1001_g Y 0.0187766f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_65 A Y 0.0984922f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_66 N_A_M1001_g N_VGND_c_139_n 0.00363059f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_VGND_c_140_n 0.0063805f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_68 A N_VGND_c_140_n 0.00222705f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_69 N_VPWR_c_93_n Y 0.0267484f $X=0.29 $Y=2.455 $X2=0 $Y2=0
cc_70 N_VPWR_c_95_n Y 0.0269916f $X=1.15 $Y=2.455 $X2=0 $Y2=0
cc_71 N_VPWR_c_96_n Y 0.00892288f $X=0.985 $Y=3.33 $X2=0 $Y2=0
cc_72 N_VPWR_c_91_n Y 0.00763575f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_73 N_Y_c_112_n N_VGND_c_139_n 0.0256433f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_74 N_Y_c_121_n N_VGND_c_139_n 0.0106426f $X=0.71 $Y=0.61 $X2=0 $Y2=0
cc_75 N_Y_M1001_d N_VGND_c_140_n 0.0021695f $X=1.01 $Y=0.235 $X2=0 $Y2=0
cc_76 N_Y_c_112_n N_VGND_c_140_n 0.0181066f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_77 N_Y_c_121_n N_VGND_c_140_n 0.00799541f $X=0.71 $Y=0.61 $X2=0 $Y2=0
cc_78 N_Y_c_121_n A_124_47# 0.001301f $X=0.71 $Y=0.61 $X2=-0.19 $Y2=-0.245
cc_79 N_VGND_c_140_n A_124_47# 0.00193852f $X=1.2 $Y=0 $X2=-0.19 $Y2=-0.245
