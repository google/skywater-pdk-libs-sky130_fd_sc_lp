* NGSPICE file created from sky130_fd_sc_lp__a22o_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_94_249# A1 a_340_49# VNB nshort w=840000u l=150000u
+  ad=4.452e+11p pd=4.42e+06u as=1.764e+11p ps=2.1e+06u
M1001 X a_94_249# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=9.114e+11p ps=7.21e+06u
M1002 VGND a_94_249# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A1 a_326_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.2096e+12p pd=9.48e+06u as=7.056e+11p ps=6.16e+06u
M1004 a_94_249# B1 a_326_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=6.678e+11p pd=6.1e+06u as=0p ps=0u
M1005 a_340_49# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_610_49# B2 VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1007 a_94_249# B1 a_610_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_94_249# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1009 a_326_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_326_367# B2 a_94_249# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_94_249# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

