* File: sky130_fd_sc_lp__mux2i_0.pex.spice
* Created: Wed Sep  2 10:00:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2I_0%S 3 7 9 11 16 20 22 25 26 27 29 30 31 34 35
+ 37 38 43 48 50
c114 34 0 8.81432e-20 $X=2.975 $Y=1.79
r115 43 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.845
+ $X2=0.665 $Y2=2.01
r116 43 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.845
+ $X2=0.665 $Y2=1.68
r117 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.665
+ $Y=1.845 $X2=0.665 $Y2=1.845
r118 38 50 2.85154 $w=3.55e-07 $l=1.17e-07 $layer=LI1_cond $X=0.712 $Y=2.127
+ $X2=0.712 $Y2=2.01
r119 38 50 0.973895 $w=3.53e-07 $l=3e-08 $layer=LI1_cond $X=0.712 $Y=1.98
+ $X2=0.712 $Y2=2.01
r120 38 44 4.38253 $w=3.53e-07 $l=1.35e-07 $layer=LI1_cond $X=0.712 $Y=1.98
+ $X2=0.712 $Y2=1.845
r121 37 44 5.84337 $w=3.53e-07 $l=1.8e-07 $layer=LI1_cond $X=0.712 $Y=1.665
+ $X2=0.712 $Y2=1.845
r122 35 49 81.3905 $w=5.4e-07 $l=5.05e-07 $layer=POLY_cond $X=2.87 $Y=1.79
+ $X2=2.87 $Y2=2.295
r123 35 48 47.7034 $w=5.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.87 $Y=1.79
+ $X2=2.87 $Y2=1.625
r124 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.975
+ $Y=1.79 $X2=2.975 $Y2=1.79
r125 32 34 30.5184 $w=2.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.005 $Y=2.505
+ $X2=3.005 $Y2=1.79
r126 30 32 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.87 $Y=2.59
+ $X2=3.005 $Y2=2.505
r127 30 31 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.87 $Y=2.59
+ $X2=2.555 $Y2=2.59
r128 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.47 $Y=2.675
+ $X2=2.555 $Y2=2.59
r129 28 29 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.47 $Y=2.675
+ $X2=2.47 $Y2=2.905
r130 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.385 $Y=2.99
+ $X2=2.47 $Y2=2.905
r131 26 27 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.385 $Y=2.99
+ $X2=1.67 $Y2=2.99
r132 25 27 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.57 $Y=2.905
+ $X2=1.67 $Y2=2.99
r133 24 25 36.6 $w=1.98e-07 $l=6.6e-07 $layer=LI1_cond $X=1.57 $Y=2.245 $X2=1.57
+ $Y2=2.905
r134 23 38 4.33824 $w=2.35e-07 $l=1.78e-07 $layer=LI1_cond $X=0.89 $Y=2.127
+ $X2=0.712 $Y2=2.127
r135 22 24 6.87405 $w=2.35e-07 $l=1.60387e-07 $layer=LI1_cond $X=1.47 $Y=2.127
+ $X2=1.57 $Y2=2.245
r136 22 23 28.4433 $w=2.33e-07 $l=5.8e-07 $layer=LI1_cond $X=1.47 $Y=2.127
+ $X2=0.89 $Y2=2.127
r137 18 20 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.495 $Y=0.845
+ $X2=2.675 $Y2=0.845
r138 16 49 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.675 $Y=2.775
+ $X2=2.675 $Y2=2.295
r139 12 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.675 $Y=0.92
+ $X2=2.675 $Y2=0.845
r140 12 48 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.675 $Y=0.92
+ $X2=2.675 $Y2=1.625
r141 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.495 $Y=0.77
+ $X2=2.495 $Y2=0.845
r142 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.495 $Y=0.77
+ $X2=2.495 $Y2=0.45
r143 7 46 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.755 $Y=2.775
+ $X2=0.755 $Y2=2.01
r144 3 45 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=0.575 $Y=0.45
+ $X2=0.575 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_0%A_47_48# 1 2 9 11 14 17 18 19 22 26 32 33 35
+ 37 38
c71 32 0 1.75857e-20 $X=1.055 $Y=0.935
c72 19 0 1.56142e-19 $X=1.055 $Y=1.44
r73 37 38 7.20939 $w=6.18e-07 $l=1.85e-07 $layer=LI1_cond $X=0.395 $Y=2.6
+ $X2=0.395 $Y2=2.415
r74 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.055
+ $Y=0.935 $X2=1.055 $Y2=0.935
r75 30 35 0.275373 $w=5.75e-07 $l=2.2e-07 $layer=LI1_cond $X=0.525 $Y=1.072
+ $X2=0.305 $Y2=1.072
r76 30 32 11.0247 $w=5.73e-07 $l=5.3e-07 $layer=LI1_cond $X=0.525 $Y=1.072
+ $X2=1.055 $Y2=1.072
r77 28 35 7.47898 $w=3.6e-07 $l=3.25552e-07 $layer=LI1_cond $X=0.225 $Y=1.36
+ $X2=0.305 $Y2=1.072
r78 28 38 43.4224 $w=2.78e-07 $l=1.055e-06 $layer=LI1_cond $X=0.225 $Y=1.36
+ $X2=0.225 $Y2=2.415
r79 24 35 7.47898 $w=3.6e-07 $l=2.87e-07 $layer=LI1_cond $X=0.305 $Y=0.785
+ $X2=0.305 $Y2=1.072
r80 24 26 8.77428 $w=4.38e-07 $l=3.35e-07 $layer=LI1_cond $X=0.305 $Y=0.785
+ $X2=0.305 $Y2=0.45
r81 20 22 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.145 $Y=2.125
+ $X2=1.385 $Y2=2.125
r82 18 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.055 $Y=1.275
+ $X2=1.055 $Y2=0.935
r83 18 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.275
+ $X2=1.055 $Y2=1.44
r84 17 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=0.77
+ $X2=1.055 $Y2=0.935
r85 12 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.385 $Y=2.2
+ $X2=1.385 $Y2=2.125
r86 12 14 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.385 $Y=2.2
+ $X2=1.385 $Y2=2.775
r87 11 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.145 $Y=2.05
+ $X2=1.145 $Y2=2.125
r88 11 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.145 $Y=2.05
+ $X2=1.145 $Y2=1.44
r89 9 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.145 $Y=0.45
+ $X2=1.145 $Y2=0.77
r90 2 37 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.415
+ $Y=2.455 $X2=0.54 $Y2=2.6
r91 1 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.24 $X2=0.36 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_0%A0 3 6 8 10 18 20 23 24 38
c59 38 0 1.56142e-19 $X=2.195 $Y=1.095
c60 18 0 1.97676e-19 $X=1.625 $Y=0.935
c61 6 0 8.81432e-20 $X=2.25 $Y=2.775
r62 23 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.9
+ $X2=2.195 $Y2=2.065
r63 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.195
+ $Y=1.9 $X2=2.195 $Y2=1.9
r64 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=0.935
+ $X2=1.625 $Y2=0.77
r65 10 38 0.734434 $w=5.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.16 $Y=1.095
+ $X2=2.195 $Y2=1.095
r66 10 38 3.93508 $w=3.3e-07 $l=2.85e-07 $layer=LI1_cond $X=2.195 $Y=1.38
+ $X2=2.195 $Y2=1.095
r67 10 24 13.8229 $w=4.98e-07 $l=5.2e-07 $layer=LI1_cond $X=2.195 $Y=1.38
+ $X2=2.195 $Y2=1.9
r68 8 10 11.2263 $w=5.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.625 $Y=1.095
+ $X2=2.16 $Y2=1.095
r69 8 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=0.935 $X2=1.625 $Y2=0.935
r70 6 26 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.25 $Y=2.775
+ $X2=2.25 $Y2=2.065
r71 3 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.535 $Y=0.45
+ $X2=1.535 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_0%A1 3 5 9 11 12 15
c51 15 0 1.75857e-20 $X=1.64 $Y=1.42
c52 12 0 1.97676e-19 $X=1.68 $Y=1.665
c53 5 0 1.8102e-21 $X=2.03 $Y=1.42
r54 18 20 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.64 $Y=1.645
+ $X2=1.64 $Y2=1.81
r55 15 18 36.0651 $w=3.6e-07 $l=2.25e-07 $layer=POLY_cond $X=1.64 $Y=1.42
+ $X2=1.64 $Y2=1.645
r56 12 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.645 $X2=1.625 $Y2=1.645
r57 11 12 16.8893 $w=2.88e-07 $l=4.25e-07 $layer=LI1_cond $X=1.2 $Y=1.695
+ $X2=1.625 $Y2=1.695
r58 7 9 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=2.105 $Y=1.345
+ $X2=2.105 $Y2=0.45
r59 6 15 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.82 $Y=1.42 $X2=1.64
+ $Y2=1.42
r60 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.03 $Y=1.42
+ $X2=2.105 $Y2=1.345
r61 5 6 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.03 $Y=1.42 $X2=1.82
+ $Y2=1.42
r62 3 20 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=1.745 $Y=2.775
+ $X2=1.745 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_0%VPWR 1 2 9 13 15 16 17 18 20 31 33
r44 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 28 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 25 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=3.33
+ $X2=1.065 $Y2=3.33
r49 25 27 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=1.23 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=1.065 $Y2=3.33
r53 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=0.72
+ $Y2=3.33
r54 18 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 18 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 16 27 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.89 $Y2=3.33
r58 15 30 4.66471 $w=1.7e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=3.33
+ $X2=2.89 $Y2=3.33
r60 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=3.245
+ $X2=2.89 $Y2=3.33
r61 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.89 $Y=3.245
+ $X2=2.89 $Y2=2.97
r62 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=3.245
+ $X2=1.065 $Y2=3.33
r63 7 9 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=1.065 $Y=3.245
+ $X2=1.065 $Y2=2.6
r64 2 13 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=2.75
+ $Y=2.455 $X2=2.89 $Y2=2.97
r65 1 9 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=0.83
+ $Y=2.455 $X2=1.065 $Y2=2.6
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_0%Y 1 2 9 11 12 14 15 16
c49 11 0 1.8102e-21 $X=2.53 $Y=2.25
r50 16 19 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=2.16 $Y=0.462
+ $X2=1.825 $Y2=0.462
r51 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.53 $Y=0.462
+ $X2=2.16 $Y2=0.462
r52 13 15 7.97992 $w=3.55e-07 $l=2.16365e-07 $layer=LI1_cond $X=2.615 $Y=0.64
+ $X2=2.53 $Y2=0.462
r53 13 14 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=2.615 $Y=0.64
+ $X2=2.615 $Y2=2.165
r54 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.53 $Y=2.25
+ $X2=2.615 $Y2=2.165
r55 11 12 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.53 $Y=2.25
+ $X2=2.17 $Y2=2.25
r56 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.005 $Y=2.335
+ $X2=2.17 $Y2=2.25
r57 7 9 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.005 $Y=2.335
+ $X2=2.005 $Y2=2.62
r58 2 9 600 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=2.455 $X2=2.005 $Y2=2.62
r59 1 19 182 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_NDIFF $count=1 $X=1.61
+ $Y=0.24 $X2=1.825 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_0%VGND 1 2 11 13 15 17 19 28 32
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r43 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r45 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r46 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 20 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.87
+ $Y2=0
r48 20 22 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r49 19 31 4.00852 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=3.115
+ $Y2=0
r50 19 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.64
+ $Y2=0
r51 17 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r52 17 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r53 13 31 3.23954 $w=2.65e-07 $l=1.49579e-07 $layer=LI1_cond $X=3.002 $Y=0.085
+ $X2=3.115 $Y2=0
r54 13 15 15.8733 $w=2.63e-07 $l=3.65e-07 $layer=LI1_cond $X=3.002 $Y=0.085
+ $X2=3.002 $Y2=0.45
r55 9 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=0.085 $X2=0.87
+ $Y2=0
r56 9 11 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.87 $Y=0.085
+ $X2=0.87 $Y2=0.45
r57 2 15 182 $w=1.7e-07 $l=4.93964e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.24 $X2=2.97 $Y2=0.45
r58 1 11 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.24 $X2=0.87 $Y2=0.45
.ends

