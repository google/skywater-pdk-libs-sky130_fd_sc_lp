# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__fa_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__fa_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 0.440000 7.235000 0.670000 ;
        RECT 6.905000 0.265000 7.235000 0.440000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125000 1.235000 4.710000 1.405000 ;
        RECT 3.125000 1.405000 3.775000 1.565000 ;
        RECT 3.605000 1.565000 3.775000 2.100000 ;
        RECT 3.605000 2.100000 4.210000 2.165000 ;
        RECT 3.605000 2.165000 9.135000 2.270000 ;
        RECT 4.040000 2.270000 9.135000 2.335000 ;
        RECT 4.435000 1.180000 4.710000 1.235000 ;
        RECT 4.435000 1.405000 4.710000 1.565000 ;
        RECT 8.820000 1.605000 9.135000 2.165000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.939000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.955000 1.590000 4.225000 1.750000 ;
        RECT 3.955000 1.750000 4.560000 1.815000 ;
        RECT 3.955000 1.815000 8.610000 1.920000 ;
        RECT 4.390000 1.920000 8.610000 1.985000 ;
        RECT 6.800000 1.550000 7.080000 1.815000 ;
        RECT 8.280000 1.605000 8.610000 1.815000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.405000 0.545000 0.865000 ;
        RECT 0.115000 0.865000 0.445000 2.935000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.115000 0.310000 10.470000 1.040000 ;
        RECT 10.115000 2.075000 10.470000 3.065000 ;
        RECT 10.300000 1.040000 10.470000 2.075000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.245000 10.560000 3.415000 ;
      RECT 0.645000  1.895000  0.975000 3.245000 ;
      RECT 0.700000  1.045000  1.030000 1.545000 ;
      RECT 0.700000  1.545000  2.945000 1.715000 ;
      RECT 1.005000  0.085000  1.575000 0.865000 ;
      RECT 1.205000  1.895000  2.415000 2.065000 ;
      RECT 1.205000  2.065000  1.535000 3.065000 ;
      RECT 1.405000  0.865000  1.575000 1.195000 ;
      RECT 1.405000  1.195000  2.595000 1.365000 ;
      RECT 1.735000  2.245000  2.065000 3.245000 ;
      RECT 1.755000  0.320000  4.230000 0.490000 ;
      RECT 1.755000  0.490000  2.085000 1.015000 ;
      RECT 2.245000  2.065000  2.415000 2.095000 ;
      RECT 2.245000  2.095000  3.075000 2.265000 ;
      RECT 2.265000  0.685000  2.595000 1.195000 ;
      RECT 2.265000  2.445000  2.595000 2.895000 ;
      RECT 2.265000  2.895000  4.390000 3.065000 ;
      RECT 2.775000  0.830000  5.060000 1.000000 ;
      RECT 2.775000  1.000000  3.605000 1.055000 ;
      RECT 2.775000  1.055000  2.945000 1.545000 ;
      RECT 2.775000  1.715000  2.945000 1.745000 ;
      RECT 2.775000  1.745000  3.425000 1.915000 ;
      RECT 2.825000  2.265000  3.075000 2.715000 ;
      RECT 3.250000  0.685000  3.580000 0.830000 ;
      RECT 3.255000  1.915000  3.425000 2.450000 ;
      RECT 3.255000  2.450000  3.860000 2.715000 ;
      RECT 3.900000  0.490000  4.230000 0.650000 ;
      RECT 4.060000  2.515000  4.390000 2.895000 ;
      RECT 4.490000  0.085000  4.820000 0.650000 ;
      RECT 4.690000  2.515000  5.020000 3.245000 ;
      RECT 4.890000  1.000000  5.060000 1.465000 ;
      RECT 4.890000  1.465000  6.620000 1.635000 ;
      RECT 5.080000  0.320000  5.410000 0.650000 ;
      RECT 5.220000  2.515000  7.845000 2.685000 ;
      RECT 5.220000  2.685000  5.550000 3.065000 ;
      RECT 5.240000  0.650000  5.410000 1.115000 ;
      RECT 5.240000  1.115000  6.270000 1.285000 ;
      RECT 5.590000  0.085000  5.920000 0.935000 ;
      RECT 5.750000  2.865000  6.080000 3.245000 ;
      RECT 6.100000  0.850000  7.745000 1.020000 ;
      RECT 6.100000  1.020000  6.270000 1.115000 ;
      RECT 6.450000  1.200000  7.430000 1.305000 ;
      RECT 6.450000  1.305000  8.010000 1.370000 ;
      RECT 6.450000  1.370000  6.620000 1.465000 ;
      RECT 7.260000  1.370000  8.010000 1.635000 ;
      RECT 7.415000  0.685000  7.745000 0.850000 ;
      RECT 7.515000  2.685000  7.845000 3.065000 ;
      RECT 7.975000  0.685000  8.360000 1.125000 ;
      RECT 8.045000  2.515000  9.485000 2.685000 ;
      RECT 8.045000  2.685000  8.375000 3.065000 ;
      RECT 8.190000  1.125000  8.360000 1.220000 ;
      RECT 8.190000  1.220000 10.120000 1.390000 ;
      RECT 9.270000  0.085000  9.600000 0.770000 ;
      RECT 9.315000  1.390000  9.485000 2.515000 ;
      RECT 9.665000  2.075000  9.915000 3.245000 ;
      RECT 9.820000  1.390000 10.120000 1.890000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_lp__fa_lp
END LIBRARY
