* File: sky130_fd_sc_lp__clkinv_0.pxi.spice
* Created: Fri Aug 28 10:17:21 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINV_0%A N_A_M1000_g N_A_M1001_g A A A A N_A_c_22_n
+ PM_SKY130_FD_SC_LP__CLKINV_0%A
x_PM_SKY130_FD_SC_LP__CLKINV_0%VPWR N_VPWR_M1001_s N_VPWR_c_41_n N_VPWR_c_42_n
+ VPWR N_VPWR_c_43_n N_VPWR_c_40_n PM_SKY130_FD_SC_LP__CLKINV_0%VPWR
x_PM_SKY130_FD_SC_LP__CLKINV_0%Y N_Y_M1000_d N_Y_M1001_d N_Y_c_53_n Y Y Y Y Y Y
+ Y PM_SKY130_FD_SC_LP__CLKINV_0%Y
x_PM_SKY130_FD_SC_LP__CLKINV_0%VGND N_VGND_M1000_s N_VGND_c_66_n N_VGND_c_67_n
+ VGND N_VGND_c_68_n N_VGND_c_69_n PM_SKY130_FD_SC_LP__CLKINV_0%VGND
cc_1 VNB N_A_M1000_g 0.0290158f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.56
cc_2 VNB N_A_M1001_g 0.00168831f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.63
cc_3 VNB A 0.0340643f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_4 VNB N_A_c_22_n 0.0850037f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_5 VNB N_VPWR_c_40_n 0.0442671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_Y_c_53_n 0.0152597f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB Y 0.047681f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_VGND_c_66_n 0.0115566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_VGND_c_67_n 0.0215368f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.63
cc_10 VNB N_VGND_c_68_n 0.0166435f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_11 VNB N_VGND_c_69_n 0.0900768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VPB N_A_M1001_g 0.0571374f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.63
cc_13 VPB A 0.0276907f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_14 VPB N_VPWR_c_41_n 0.0111987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_15 VPB N_VPWR_c_42_n 0.0409159f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.63
cc_16 VPB N_VPWR_c_43_n 0.0176876f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_17 VPB N_VPWR_c_40_n 0.0493087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_18 VPB Y 0.0639382f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_19 N_A_M1001_g N_VPWR_c_42_n 0.00569522f $X=0.485 $Y=2.63 $X2=0 $Y2=0
cc_20 A N_VPWR_c_42_n 0.0274534f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_21 N_A_c_22_n N_VPWR_c_42_n 8.55346e-19 $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_22 N_A_M1001_g N_VPWR_c_43_n 0.00570944f $X=0.485 $Y=2.63 $X2=0 $Y2=0
cc_23 N_A_M1001_g N_VPWR_c_40_n 0.00542671f $X=0.485 $Y=2.63 $X2=0 $Y2=0
cc_24 N_A_M1000_g N_Y_c_53_n 6.61049e-19 $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_25 N_A_M1000_g Y 0.0224292f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_26 A Y 0.103567f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_27 N_A_c_22_n Y 0.0224292f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_28 N_A_M1000_g N_VGND_c_67_n 0.0142623f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_29 A N_VGND_c_67_n 0.0242687f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_30 N_A_c_22_n N_VGND_c_67_n 0.00161326f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_31 N_A_M1000_g N_VGND_c_68_n 0.00396895f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_32 N_A_M1000_g N_VGND_c_69_n 0.00789173f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_33 A N_VGND_c_69_n 0.00185499f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_34 N_VPWR_c_42_n Y 0.00147627f $X=0.27 $Y=2.465 $X2=0 $Y2=0
cc_35 N_VPWR_c_43_n Y 0.0125142f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_36 N_VPWR_c_40_n Y 0.011055f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_37 N_Y_c_53_n N_VGND_c_68_n 0.00968744f $X=0.7 $Y=0.56 $X2=0 $Y2=0
cc_38 N_Y_c_53_n N_VGND_c_69_n 0.00962496f $X=0.7 $Y=0.56 $X2=0 $Y2=0
cc_39 Y N_VGND_c_69_n 0.0014137f $X=0.635 $Y=0.84 $X2=0 $Y2=0
