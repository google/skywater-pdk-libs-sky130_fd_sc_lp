* File: sky130_fd_sc_lp__dfsbp_2.pxi.spice
* Created: Fri Aug 28 10:22:46 2020
* 
x_PM_SKY130_FD_SC_LP__DFSBP_2%CLK N_CLK_M1002_g N_CLK_M1000_g CLK CLK
+ N_CLK_c_264_n N_CLK_c_265_n PM_SKY130_FD_SC_LP__DFSBP_2%CLK
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_129_179# N_A_129_179#_M1002_d
+ N_A_129_179#_M1000_d N_A_129_179#_c_318_n N_A_129_179#_M1036_g
+ N_A_129_179#_c_319_n N_A_129_179#_M1006_g N_A_129_179#_M1033_g
+ N_A_129_179#_c_290_n N_A_129_179#_c_291_n N_A_129_179#_M1028_g
+ N_A_129_179#_M1009_g N_A_129_179#_M1020_g N_A_129_179#_c_323_n
+ N_A_129_179#_c_293_n N_A_129_179#_c_325_n N_A_129_179#_c_294_n
+ N_A_129_179#_c_326_n N_A_129_179#_c_295_n N_A_129_179#_c_296_n
+ N_A_129_179#_c_297_n N_A_129_179#_c_298_n N_A_129_179#_c_299_n
+ N_A_129_179#_c_300_n N_A_129_179#_c_301_n N_A_129_179#_c_328_n
+ N_A_129_179#_c_302_n N_A_129_179#_c_303_n N_A_129_179#_c_304_n
+ N_A_129_179#_c_305_n N_A_129_179#_c_306_n N_A_129_179#_c_307_n
+ N_A_129_179#_c_308_n N_A_129_179#_c_309_n N_A_129_179#_c_329_n
+ N_A_129_179#_c_310_n N_A_129_179#_c_331_n N_A_129_179#_c_332_n
+ N_A_129_179#_c_311_n N_A_129_179#_c_312_n N_A_129_179#_c_313_n
+ N_A_129_179#_c_314_n N_A_129_179#_c_315_n N_A_129_179#_c_316_n
+ N_A_129_179#_c_317_n PM_SKY130_FD_SC_LP__DFSBP_2%A_129_179#
x_PM_SKY130_FD_SC_LP__DFSBP_2%D N_D_M1032_g N_D_M1008_g D D D N_D_c_556_n
+ N_D_c_559_n PM_SKY130_FD_SC_LP__DFSBP_2%D
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_721_99# N_A_721_99#_M1023_s N_A_721_99#_M1019_d
+ N_A_721_99#_c_600_n N_A_721_99#_M1025_g N_A_721_99#_M1031_g
+ N_A_721_99#_c_601_n N_A_721_99#_c_602_n N_A_721_99#_c_608_n
+ N_A_721_99#_c_609_n N_A_721_99#_c_603_n N_A_721_99#_c_604_n
+ N_A_721_99#_c_610_n N_A_721_99#_c_611_n N_A_721_99#_c_612_n
+ N_A_721_99#_c_613_n N_A_721_99#_c_605_n N_A_721_99#_c_678_p
+ N_A_721_99#_c_614_n N_A_721_99#_c_606_n N_A_721_99#_c_616_n
+ PM_SKY130_FD_SC_LP__DFSBP_2%A_721_99#
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_593_125# N_A_593_125#_M1033_d
+ N_A_593_125#_M1037_d N_A_593_125#_M1019_g N_A_593_125#_M1023_g
+ N_A_593_125#_c_703_n N_A_593_125#_M1003_g N_A_593_125#_c_704_n
+ N_A_593_125#_c_705_n N_A_593_125#_c_706_n N_A_593_125#_M1010_g
+ N_A_593_125#_c_707_n N_A_593_125#_c_716_n N_A_593_125#_c_708_n
+ N_A_593_125#_c_718_n N_A_593_125#_c_719_n N_A_593_125#_c_720_n
+ N_A_593_125#_c_721_n N_A_593_125#_c_722_n N_A_593_125#_c_709_n
+ N_A_593_125#_c_710_n N_A_593_125#_c_724_n N_A_593_125#_c_767_n
+ N_A_593_125#_c_725_n N_A_593_125#_c_726_n N_A_593_125#_c_727_n
+ N_A_593_125#_c_711_n N_A_593_125#_c_729_n
+ PM_SKY130_FD_SC_LP__DFSBP_2%A_593_125#
x_PM_SKY130_FD_SC_LP__DFSBP_2%SET_B N_SET_B_M1022_g N_SET_B_c_877_n
+ N_SET_B_M1017_g N_SET_B_M1005_g N_SET_B_c_880_n N_SET_B_M1014_g
+ N_SET_B_c_882_n N_SET_B_c_883_n N_SET_B_c_884_n N_SET_B_c_885_n
+ N_SET_B_c_928_n N_SET_B_c_886_n N_SET_B_c_929_n N_SET_B_c_887_n
+ N_SET_B_c_888_n N_SET_B_c_889_n N_SET_B_c_890_n SET_B N_SET_B_c_891_n SET_B
+ PM_SKY130_FD_SC_LP__DFSBP_2%SET_B
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_191_21# N_A_191_21#_M1036_s N_A_191_21#_M1006_s
+ N_A_191_21#_c_994_n N_A_191_21#_c_995_n N_A_191_21#_c_1003_n
+ N_A_191_21#_c_1004_n N_A_191_21#_M1037_g N_A_191_21#_M1021_g
+ N_A_191_21#_c_997_n N_A_191_21#_M1026_g N_A_191_21#_M1029_g
+ N_A_191_21#_c_999_n N_A_191_21#_c_1000_n N_A_191_21#_c_1007_n
+ N_A_191_21#_c_1008_n N_A_191_21#_c_1001_n
+ PM_SKY130_FD_SC_LP__DFSBP_2%A_191_21#
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_1533_258# N_A_1533_258#_M1007_s
+ N_A_1533_258#_M1024_s N_A_1533_258#_M1013_g N_A_1533_258#_c_1126_n
+ N_A_1533_258#_c_1127_n N_A_1533_258#_M1011_g N_A_1533_258#_c_1128_n
+ N_A_1533_258#_c_1129_n N_A_1533_258#_c_1135_n N_A_1533_258#_c_1130_n
+ N_A_1533_258#_c_1131_n N_A_1533_258#_c_1137_n N_A_1533_258#_c_1132_n
+ N_A_1533_258#_c_1133_n PM_SKY130_FD_SC_LP__DFSBP_2%A_1533_258#
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_1360_451# N_A_1360_451#_M1020_d
+ N_A_1360_451#_M1009_d N_A_1360_451#_M1005_d N_A_1360_451#_c_1210_n
+ N_A_1360_451#_M1024_g N_A_1360_451#_M1007_g N_A_1360_451#_c_1212_n
+ N_A_1360_451#_M1004_g N_A_1360_451#_M1015_g N_A_1360_451#_c_1215_n
+ N_A_1360_451#_M1035_g N_A_1360_451#_M1030_g N_A_1360_451#_c_1218_n
+ N_A_1360_451#_M1034_g N_A_1360_451#_M1018_g N_A_1360_451#_c_1221_n
+ N_A_1360_451#_c_1222_n N_A_1360_451#_c_1223_n N_A_1360_451#_c_1224_n
+ N_A_1360_451#_c_1225_n N_A_1360_451#_c_1226_n N_A_1360_451#_c_1227_n
+ N_A_1360_451#_c_1228_n N_A_1360_451#_c_1238_n N_A_1360_451#_c_1249_n
+ N_A_1360_451#_c_1229_n N_A_1360_451#_c_1239_n N_A_1360_451#_c_1230_n
+ PM_SKY130_FD_SC_LP__DFSBP_2%A_1360_451#
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_2227_367# N_A_2227_367#_M1018_d
+ N_A_2227_367#_M1034_d N_A_2227_367#_M1012_g N_A_2227_367#_M1001_g
+ N_A_2227_367#_c_1366_n N_A_2227_367#_c_1367_n N_A_2227_367#_M1027_g
+ N_A_2227_367#_M1016_g N_A_2227_367#_c_1369_n N_A_2227_367#_c_1370_n
+ N_A_2227_367#_c_1377_n N_A_2227_367#_c_1371_n N_A_2227_367#_c_1372_n
+ N_A_2227_367#_c_1373_n N_A_2227_367#_c_1374_n
+ PM_SKY130_FD_SC_LP__DFSBP_2%A_2227_367#
x_PM_SKY130_FD_SC_LP__DFSBP_2%VPWR N_VPWR_M1000_s N_VPWR_M1006_d N_VPWR_M1031_d
+ N_VPWR_M1017_d N_VPWR_M1013_d N_VPWR_M1024_d N_VPWR_M1035_d N_VPWR_M1001_d
+ N_VPWR_M1016_d N_VPWR_c_1420_n N_VPWR_c_1421_n N_VPWR_c_1422_n N_VPWR_c_1423_n
+ N_VPWR_c_1424_n N_VPWR_c_1425_n N_VPWR_c_1426_n N_VPWR_c_1427_n
+ N_VPWR_c_1428_n N_VPWR_c_1429_n VPWR N_VPWR_c_1430_n N_VPWR_c_1431_n
+ N_VPWR_c_1432_n N_VPWR_c_1433_n N_VPWR_c_1434_n N_VPWR_c_1435_n
+ N_VPWR_c_1436_n N_VPWR_c_1437_n N_VPWR_c_1438_n N_VPWR_c_1439_n
+ N_VPWR_c_1440_n N_VPWR_c_1441_n N_VPWR_c_1442_n N_VPWR_c_1443_n
+ N_VPWR_c_1444_n N_VPWR_c_1419_n PM_SKY130_FD_SC_LP__DFSBP_2%VPWR
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_507_125# N_A_507_125#_M1032_d
+ N_A_507_125#_M1008_d N_A_507_125#_c_1573_n N_A_507_125#_c_1574_n
+ N_A_507_125#_c_1575_n N_A_507_125#_c_1592_n
+ PM_SKY130_FD_SC_LP__DFSBP_2%A_507_125#
x_PM_SKY130_FD_SC_LP__DFSBP_2%Q_N N_Q_N_M1015_d N_Q_N_M1004_s Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1611_n PM_SKY130_FD_SC_LP__DFSBP_2%Q_N
x_PM_SKY130_FD_SC_LP__DFSBP_2%Q N_Q_M1012_d N_Q_M1001_s Q N_Q_c_1631_n
+ PM_SKY130_FD_SC_LP__DFSBP_2%Q
x_PM_SKY130_FD_SC_LP__DFSBP_2%VGND N_VGND_M1002_s N_VGND_M1036_d N_VGND_M1025_d
+ N_VGND_M1022_d N_VGND_M1014_d N_VGND_M1007_d N_VGND_M1030_s N_VGND_M1012_s
+ N_VGND_M1027_s N_VGND_c_1648_n N_VGND_c_1649_n N_VGND_c_1650_n N_VGND_c_1651_n
+ N_VGND_c_1652_n N_VGND_c_1653_n N_VGND_c_1654_n N_VGND_c_1655_n
+ N_VGND_c_1656_n N_VGND_c_1657_n N_VGND_c_1658_n N_VGND_c_1659_n
+ N_VGND_c_1660_n N_VGND_c_1661_n N_VGND_c_1662_n N_VGND_c_1663_n VGND
+ N_VGND_c_1664_n N_VGND_c_1665_n N_VGND_c_1666_n N_VGND_c_1667_n
+ N_VGND_c_1668_n N_VGND_c_1669_n N_VGND_c_1670_n N_VGND_c_1671_n
+ N_VGND_c_1672_n N_VGND_c_1673_n N_VGND_c_1674_n
+ PM_SKY130_FD_SC_LP__DFSBP_2%VGND
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_1173_125# N_A_1173_125#_M1003_d
+ N_A_1173_125#_M1026_d N_A_1173_125#_c_1795_n N_A_1173_125#_c_1796_n
+ N_A_1173_125#_c_1797_n PM_SKY130_FD_SC_LP__DFSBP_2%A_1173_125#
x_PM_SKY130_FD_SC_LP__DFSBP_2%A_1280_159# N_A_1280_159#_M1020_s
+ N_A_1280_159#_M1011_s N_A_1280_159#_c_1822_n N_A_1280_159#_c_1823_n
+ N_A_1280_159#_c_1824_n N_A_1280_159#_c_1825_n
+ PM_SKY130_FD_SC_LP__DFSBP_2%A_1280_159#
cc_1 VNB N_CLK_M1002_g 0.027345f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.105
cc_2 VNB N_CLK_c_264_n 0.0207654f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.65
cc_3 VNB N_CLK_c_265_n 0.0153157f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.65
cc_4 VNB N_A_129_179#_M1033_g 0.0303014f $X=-0.19 $Y=-0.245 $X2=0.467 $Y2=1.815
cc_5 VNB N_A_129_179#_c_290_n 0.0498267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_129_179#_c_291_n 0.00746415f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.665
cc_7 VNB N_A_129_179#_M1020_g 0.0197192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_129_179#_c_293_n 0.0101122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_129_179#_c_294_n 0.00346977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_129_179#_c_295_n 0.00443533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_129_179#_c_296_n 0.0083242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_129_179#_c_297_n 0.00399416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_129_179#_c_298_n 0.0218403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_129_179#_c_299_n 0.00200511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_129_179#_c_300_n 0.00292147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_129_179#_c_301_n 0.00357568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_129_179#_c_302_n 0.0130502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_129_179#_c_303_n 0.00820925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_129_179#_c_304_n 0.0180314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_129_179#_c_305_n 0.00405453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_129_179#_c_306_n 8.21017e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_129_179#_c_307_n 0.00450953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_129_179#_c_308_n 0.00154637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_129_179#_c_309_n 0.0175327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_129_179#_c_310_n 0.00311569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_129_179#_c_311_n 0.031916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_129_179#_c_312_n 0.00546989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_129_179#_c_313_n 0.00116809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_129_179#_c_314_n 0.00473844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_129_179#_c_315_n 0.00114695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_129_179#_c_316_n 0.0166216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_129_179#_c_317_n 0.0167784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_D_M1032_g 0.024863f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.105
cc_34 VNB D 0.0148843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_D_c_556_n 0.0506414f $X=-0.19 $Y=-0.245 $X2=0.467 $Y2=1.485
cc_36 VNB N_A_721_99#_c_600_n 0.0145198f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.295
cc_37 VNB N_A_721_99#_c_601_n 0.0343226f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.65
cc_38 VNB N_A_721_99#_c_602_n 0.00890883f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.65
cc_39 VNB N_A_721_99#_c_603_n 0.012542f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=2.035
cc_40 VNB N_A_721_99#_c_604_n 0.0204147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_721_99#_c_605_n 0.00479249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_721_99#_c_606_n 0.00699236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_593_125#_M1023_g 0.0282805f $X=-0.19 $Y=-0.245 $X2=0.467 $Y2=1.65
cc_44 VNB N_A_593_125#_c_703_n 0.0176926f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.65
cc_45 VNB N_A_593_125#_c_704_n 0.0227287f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.65
cc_46 VNB N_A_593_125#_c_705_n 0.00819466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_593_125#_c_706_n 0.00812845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_593_125#_c_707_n 0.00917315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_593_125#_c_708_n 0.00498914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_593_125#_c_709_n 0.00388207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_593_125#_c_710_n 0.00154637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_593_125#_c_711_n 0.001989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_SET_B_M1022_g 0.031275f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.105
cc_54 VNB N_SET_B_M1014_g 0.0605817f $X=-0.19 $Y=-0.245 $X2=0.467 $Y2=1.815
cc_55 VNB N_A_191_21#_c_994_n 0.0644258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_191_21#_c_995_n 0.142083f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_57 VNB N_A_191_21#_M1021_g 0.0332428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_191_21#_c_997_n 0.292083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_191_21#_M1026_g 0.047845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_191_21#_c_999_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_191_21#_c_1000_n 0.00827035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_191_21#_c_1001_n 0.0508588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1533_258#_M1013_g 0.0144565f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_64 VNB N_A_1533_258#_c_1126_n 0.0150791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1533_258#_c_1127_n 0.0103137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1533_258#_c_1128_n 0.0311361f $X=-0.19 $Y=-0.245 $X2=0.467
+ $Y2=1.485
cc_67 VNB N_A_1533_258#_c_1129_n 0.042453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1533_258#_c_1130_n 0.00304327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1533_258#_c_1131_n 0.00369788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1533_258#_c_1132_n 0.00767571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1533_258#_c_1133_n 0.0205998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1360_451#_c_1210_n 0.0275866f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_73 VNB N_A_1360_451#_M1007_g 0.0311595f $X=-0.19 $Y=-0.245 $X2=0.467
+ $Y2=1.485
cc_74 VNB N_A_1360_451#_c_1212_n 0.0158915f $X=-0.19 $Y=-0.245 $X2=0.312
+ $Y2=1.65
cc_75 VNB N_A_1360_451#_M1004_g 0.00906478f $X=-0.19 $Y=-0.245 $X2=0.312
+ $Y2=2.035
cc_76 VNB N_A_1360_451#_M1015_g 0.0272052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1360_451#_c_1215_n 0.00950863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1360_451#_M1035_g 0.00850052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1360_451#_M1030_g 0.0264171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1360_451#_c_1218_n 0.01503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1360_451#_M1034_g 0.0108726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1360_451#_M1018_g 0.0301274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1360_451#_c_1221_n 0.00302468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1360_451#_c_1222_n 0.00302468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1360_451#_c_1223_n 0.00779661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1360_451#_c_1224_n 0.00173353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1360_451#_c_1225_n 4.03688e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1360_451#_c_1226_n 0.0176629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1360_451#_c_1227_n 3.09182e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1360_451#_c_1228_n 0.0258826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1360_451#_c_1229_n 0.00107514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1360_451#_c_1230_n 0.00310098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2227_367#_c_1366_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.65
cc_94 VNB N_A_2227_367#_c_1367_n 0.019242f $X=-0.19 $Y=-0.245 $X2=0.467
+ $Y2=1.485
cc_95 VNB N_A_2227_367#_M1016_g 0.0127436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2227_367#_c_1369_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2227_367#_c_1370_n 0.00795178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2227_367#_c_1371_n 0.00831328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2227_367#_c_1372_n 0.00325142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2227_367#_c_1373_n 0.0286122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2227_367#_c_1374_n 0.0176741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VPWR_c_1419_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_507_125#_c_1573_n 0.00424025f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_104 VNB N_A_507_125#_c_1574_n 0.00302783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_507_125#_c_1575_n 0.00464982f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.65
cc_106 VNB N_Q_N_c_1611_n 0.00574359f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=2.035
cc_107 VNB N_Q_c_1631_n 0.00700489f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_108 VNB N_VGND_c_1648_n 0.0131994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1649_n 0.042409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1650_n 0.00842751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1651_n 0.0150969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1652_n 0.0169475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1653_n 0.0238188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1654_n 0.0214063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1655_n 0.0170443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1656_n 0.0237637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1657_n 0.0259125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1658_n 0.0111613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1659_n 0.0515345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1660_n 0.0338008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1661_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1662_n 0.0403309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1663_n 0.0034624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1664_n 0.0353057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1665_n 0.0741046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1666_n 0.0151073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1667_n 0.0206107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1668_n 0.0166935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1669_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1670_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1671_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1672_n 0.00548201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1673_n 0.0058666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1674_n 0.669354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_1173_125#_c_1795_n 0.0121706f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_136 VNB N_A_1173_125#_c_1796_n 0.00494035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_1173_125#_c_1797_n 0.0322206f $X=-0.19 $Y=-0.245 $X2=0.467
+ $Y2=1.65
cc_138 VNB N_A_1280_159#_c_1822_n 0.00448357f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_139 VNB N_A_1280_159#_c_1823_n 0.0038588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_1280_159#_c_1824_n 0.00336181f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.65
cc_141 VNB N_A_1280_159#_c_1825_n 0.00836698f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.65
cc_142 VPB N_CLK_M1000_g 0.0243486f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.295
cc_143 VPB N_CLK_c_264_n 0.0198887f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.65
cc_144 VPB N_CLK_c_265_n 0.0235981f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.65
cc_145 VPB N_A_129_179#_c_318_n 0.048967f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.295
cc_146 VPB N_A_129_179#_c_319_n 0.0173493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_129_179#_c_290_n 0.00440239f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_129_179#_M1028_g 0.0359776f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_129_179#_M1009_g 0.0255636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_129_179#_c_323_n 0.0212718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_129_179#_c_293_n 0.0142931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_129_179#_c_325_n 0.0164999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_129_179#_c_326_n 0.00357419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_129_179#_c_301_n 0.00142676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_129_179#_c_328_n 0.0277169f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_129_179#_c_329_n 0.00526208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_129_179#_c_310_n 0.0107537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_129_179#_c_331_n 0.00787763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_129_179#_c_332_n 0.0628535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_129_179#_c_315_n 0.00142111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_D_M1008_g 0.0215991f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.295
cc_162 VPB D 0.013361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_D_c_559_n 0.032237f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.665
cc_164 VPB N_A_721_99#_M1031_g 0.0196795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_721_99#_c_608_n 0.0156066f $X=-0.19 $Y=1.655 $X2=0.467 $Y2=1.485
cc_166 VPB N_A_721_99#_c_609_n 0.00803772f $X=-0.19 $Y=1.655 $X2=0.467 $Y2=1.815
cc_167 VPB N_A_721_99#_c_610_n 8.61815e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_721_99#_c_611_n 0.0382403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_721_99#_c_612_n 0.00716669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_721_99#_c_613_n 0.0029358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_721_99#_c_614_n 0.00651506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_721_99#_c_606_n 0.00938535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_721_99#_c_616_n 0.0268406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_593_125#_M1019_g 0.0324763f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_175 VPB N_A_593_125#_c_706_n 0.00308755f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_593_125#_M1010_g 0.0226933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_593_125#_c_707_n 0.00784992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_593_125#_c_716_n 0.0177599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_593_125#_c_708_n 0.0114586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_593_125#_c_718_n 0.00107182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_593_125#_c_719_n 0.00865829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_593_125#_c_720_n 0.00632449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_593_125#_c_721_n 0.0150433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_593_125#_c_722_n 0.00325835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_593_125#_c_709_n 0.00407459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_593_125#_c_724_n 0.0040683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_593_125#_c_725_n 0.00240893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_593_125#_c_726_n 0.00104991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_593_125#_c_727_n 0.0326005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_593_125#_c_711_n 0.00231519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_593_125#_c_729_n 0.0349705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_SET_B_M1022_g 0.0107258f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.105
cc_193 VPB N_SET_B_c_877_n 0.0334051f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.815
cc_194 VPB N_SET_B_M1017_g 0.0305799f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.295
cc_195 VPB N_SET_B_M1005_g 0.0247822f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_SET_B_c_880_n 0.0252791f $X=-0.19 $Y=1.655 $X2=0.467 $Y2=1.65
cc_197 VPB N_SET_B_M1014_g 0.00980511f $X=-0.19 $Y=1.655 $X2=0.467 $Y2=1.815
cc_198 VPB N_SET_B_c_882_n 0.0158038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_SET_B_c_883_n 0.0306698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_SET_B_c_884_n 0.0059433f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=2.035
cc_201 VPB N_SET_B_c_885_n 0.002006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_SET_B_c_886_n 0.0140524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_SET_B_c_887_n 0.00834845f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_SET_B_c_888_n 0.00449279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_SET_B_c_889_n 0.00688987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_SET_B_c_890_n 0.0163745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_SET_B_c_891_n 0.031901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_191_21#_c_994_n 0.00578679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_191_21#_c_1003_n 0.0886979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_191_21#_c_1004_n 0.0589354f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_191_21#_M1037_g 0.0477022f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.65
cc_212 VPB N_A_191_21#_M1026_g 0.0407153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_191_21#_c_1007_n 0.00664975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_191_21#_c_1008_n 0.0178943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_1533_258#_M1013_g 0.043806f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_216 VPB N_A_1533_258#_c_1135_n 0.00229952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_1533_258#_c_1131_n 0.00345607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_1533_258#_c_1137_n 0.00973131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1360_451#_c_1210_n 0.00515011f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_220 VPB N_A_1360_451#_M1024_g 0.032783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_1360_451#_M1004_g 0.0220982f $X=-0.19 $Y=1.655 $X2=0.312
+ $Y2=2.035
cc_222 VPB N_A_1360_451#_M1035_g 0.0223393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_1360_451#_M1034_g 0.0244548f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_1360_451#_c_1225_n 0.00450494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1360_451#_c_1227_n 0.0148557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_1360_451#_c_1238_n 9.43289e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_1360_451#_c_1239_n 0.0181494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_2227_367#_M1001_g 0.0230537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_2227_367#_M1016_g 0.0272176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_2227_367#_c_1377_n 0.0187079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_2227_367#_c_1371_n 0.00762681f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_2227_367#_c_1372_n 9.93106e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_2227_367#_c_1373_n 0.00762447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1420_n 0.0145833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1421_n 0.0423907f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1422_n 0.00768148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1423_n 0.0058114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1424_n 0.0223217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1425_n 0.0314809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1426_n 0.0353172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1427_n 0.0315732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1428_n 0.0111354f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1429_n 0.0585971f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1430_n 0.0409844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1431_n 0.0315251f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1432_n 0.0371076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1433_n 0.0504907f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1434_n 0.0152911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1435_n 0.0218423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1436_n 0.016215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1437_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1438_n 0.0410899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1439_n 0.0164657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1440_n 0.00535614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1441_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1442_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1443_n 0.00641775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1444_n 0.00584071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1419_n 0.133645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_507_125#_c_1574_n 0.0081072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_Q_N_c_1611_n 0.0014608f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=2.035
cc_262 VPB N_Q_c_1631_n 0.00462283f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_263 N_CLK_M1002_g N_A_129_179#_c_294_n 0.0121541f $X=0.57 $Y=1.105 $X2=0
+ $Y2=0
cc_264 N_CLK_M1000_g N_A_129_179#_c_326_n 0.00253252f $X=0.57 $Y=2.295 $X2=0
+ $Y2=0
cc_265 N_CLK_M1000_g N_A_129_179#_c_329_n 3.34329e-19 $X=0.57 $Y=2.295 $X2=0
+ $Y2=0
cc_266 N_CLK_c_264_n N_A_129_179#_c_310_n 0.0127526f $X=0.455 $Y=1.65 $X2=0
+ $Y2=0
cc_267 N_CLK_c_265_n N_A_129_179#_c_310_n 0.047649f $X=0.455 $Y=1.65 $X2=0 $Y2=0
cc_268 N_CLK_M1002_g N_A_191_21#_c_994_n 0.0146384f $X=0.57 $Y=1.105 $X2=0 $Y2=0
cc_269 N_CLK_M1000_g N_A_191_21#_c_1004_n 0.00244164f $X=0.57 $Y=2.295 $X2=0
+ $Y2=0
cc_270 N_CLK_c_264_n N_A_191_21#_c_1004_n 0.0146384f $X=0.455 $Y=1.65 $X2=0
+ $Y2=0
cc_271 N_CLK_M1002_g N_A_191_21#_c_1000_n 7.15243e-19 $X=0.57 $Y=1.105 $X2=0
+ $Y2=0
cc_272 N_CLK_c_265_n N_VPWR_M1000_s 0.00288507f $X=0.455 $Y=1.65 $X2=-0.19
+ $Y2=-0.245
cc_273 N_CLK_M1000_g N_VPWR_c_1421_n 0.00867625f $X=0.57 $Y=2.295 $X2=0 $Y2=0
cc_274 N_CLK_c_264_n N_VPWR_c_1421_n 7.43702e-19 $X=0.455 $Y=1.65 $X2=0 $Y2=0
cc_275 N_CLK_c_265_n N_VPWR_c_1421_n 0.0242732f $X=0.455 $Y=1.65 $X2=0 $Y2=0
cc_276 N_CLK_M1000_g N_VPWR_c_1430_n 0.00308317f $X=0.57 $Y=2.295 $X2=0 $Y2=0
cc_277 N_CLK_M1000_g N_VPWR_c_1419_n 0.00374015f $X=0.57 $Y=2.295 $X2=0 $Y2=0
cc_278 N_CLK_M1002_g N_VGND_c_1649_n 0.00452984f $X=0.57 $Y=1.105 $X2=0 $Y2=0
cc_279 N_CLK_c_264_n N_VGND_c_1649_n 0.00118434f $X=0.455 $Y=1.65 $X2=0 $Y2=0
cc_280 N_CLK_c_265_n N_VGND_c_1649_n 0.0191222f $X=0.455 $Y=1.65 $X2=0 $Y2=0
cc_281 N_CLK_M1002_g N_VGND_c_1660_n 0.00297774f $X=0.57 $Y=1.105 $X2=0 $Y2=0
cc_282 N_CLK_M1002_g N_VGND_c_1674_n 0.00400849f $X=0.57 $Y=1.105 $X2=0 $Y2=0
cc_283 N_A_129_179#_M1033_g N_D_M1032_g 0.0111052f $X=2.89 $Y=0.835 $X2=0 $Y2=0
cc_284 N_A_129_179#_c_296_n N_D_M1032_g 0.00597132f $X=2.24 $Y=1.105 $X2=0 $Y2=0
cc_285 N_A_129_179#_c_297_n N_D_M1032_g 0.0140154f $X=2.325 $Y=1.015 $X2=0 $Y2=0
cc_286 N_A_129_179#_c_298_n N_D_M1032_g 0.00303342f $X=3.465 $Y=0.34 $X2=0 $Y2=0
cc_287 N_A_129_179#_c_317_n N_D_M1032_g 0.00782226f $X=1.51 $Y=1.155 $X2=0 $Y2=0
cc_288 N_A_129_179#_c_319_n N_D_M1008_g 0.0137622f $X=1.86 $Y=3.075 $X2=0 $Y2=0
cc_289 N_A_129_179#_c_319_n D 0.00960782f $X=1.86 $Y=3.075 $X2=0 $Y2=0
cc_290 N_A_129_179#_c_296_n D 0.0346831f $X=2.24 $Y=1.105 $X2=0 $Y2=0
cc_291 N_A_129_179#_c_312_n D 0.00722848f $X=1.675 $Y=1.25 $X2=0 $Y2=0
cc_292 N_A_129_179#_c_291_n N_D_c_556_n 0.0130822f $X=2.965 $Y=1.49 $X2=0 $Y2=0
cc_293 N_A_129_179#_c_296_n N_D_c_556_n 0.0118177f $X=2.24 $Y=1.105 $X2=0 $Y2=0
cc_294 N_A_129_179#_c_311_n N_D_c_556_n 0.0110954f $X=1.51 $Y=1.32 $X2=0 $Y2=0
cc_295 N_A_129_179#_c_312_n N_D_c_556_n 7.41463e-19 $X=1.675 $Y=1.25 $X2=0 $Y2=0
cc_296 N_A_129_179#_c_319_n N_D_c_559_n 0.00855983f $X=1.86 $Y=3.075 $X2=0 $Y2=0
cc_297 N_A_129_179#_c_300_n N_A_721_99#_c_600_n 0.0129718f $X=3.555 $Y=1.125
+ $X2=0 $Y2=0
cc_298 N_A_129_179#_c_302_n N_A_721_99#_c_600_n 0.005146f $X=4.255 $Y=1.21 $X2=0
+ $Y2=0
cc_299 N_A_129_179#_c_303_n N_A_721_99#_c_600_n 0.00260063f $X=4.34 $Y=1.125
+ $X2=0 $Y2=0
cc_300 N_A_129_179#_c_313_n N_A_721_99#_c_600_n 7.90794e-19 $X=3.56 $Y=1.21
+ $X2=0 $Y2=0
cc_301 N_A_129_179#_c_302_n N_A_721_99#_c_601_n 0.0257801f $X=4.255 $Y=1.21
+ $X2=0 $Y2=0
cc_302 N_A_129_179#_M1033_g N_A_721_99#_c_602_n 0.00141955f $X=2.89 $Y=0.835
+ $X2=0 $Y2=0
cc_303 N_A_129_179#_c_290_n N_A_721_99#_c_602_n 0.00859568f $X=3.245 $Y=1.49
+ $X2=0 $Y2=0
cc_304 N_A_129_179#_c_301_n N_A_721_99#_c_602_n 9.98501e-19 $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_305 N_A_129_179#_c_302_n N_A_721_99#_c_602_n 0.00323441f $X=4.255 $Y=1.21
+ $X2=0 $Y2=0
cc_306 N_A_129_179#_c_313_n N_A_721_99#_c_602_n 0.00234479f $X=3.56 $Y=1.21
+ $X2=0 $Y2=0
cc_307 N_A_129_179#_M1028_g N_A_721_99#_c_609_n 0.051335f $X=3.43 $Y=2.885 $X2=0
+ $Y2=0
cc_308 N_A_129_179#_c_323_n N_A_721_99#_c_609_n 6.628e-19 $X=3.54 $Y=2.185 $X2=0
+ $Y2=0
cc_309 N_A_129_179#_c_290_n N_A_721_99#_c_603_n 5.45373e-19 $X=3.245 $Y=1.49
+ $X2=0 $Y2=0
cc_310 N_A_129_179#_c_301_n N_A_721_99#_c_603_n 0.008597f $X=3.56 $Y=1.68 $X2=0
+ $Y2=0
cc_311 N_A_129_179#_c_302_n N_A_721_99#_c_603_n 0.0337911f $X=4.255 $Y=1.21
+ $X2=0 $Y2=0
cc_312 N_A_129_179#_c_290_n N_A_721_99#_c_604_n 0.00716668f $X=3.245 $Y=1.49
+ $X2=0 $Y2=0
cc_313 N_A_129_179#_c_301_n N_A_721_99#_c_604_n 0.00500197f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_314 N_A_129_179#_M1028_g N_A_721_99#_c_611_n 0.00265253f $X=3.43 $Y=2.885
+ $X2=0 $Y2=0
cc_315 N_A_129_179#_c_302_n N_A_721_99#_c_605_n 0.0143256f $X=4.255 $Y=1.21
+ $X2=0 $Y2=0
cc_316 N_A_129_179#_c_303_n N_A_721_99#_c_605_n 0.0175547f $X=4.34 $Y=1.125
+ $X2=0 $Y2=0
cc_317 N_A_129_179#_c_304_n N_A_721_99#_c_605_n 0.0156461f $X=4.975 $Y=0.617
+ $X2=0 $Y2=0
cc_318 N_A_129_179#_c_308_n N_A_721_99#_c_605_n 0.00940407f $X=5.145 $Y=1.25
+ $X2=0 $Y2=0
cc_319 N_A_129_179#_c_301_n N_A_721_99#_c_606_n 4.24593e-19 $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_320 N_A_129_179#_c_328_n N_A_721_99#_c_606_n 0.00570195f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_321 N_A_129_179#_c_301_n N_A_721_99#_c_616_n 7.07317e-19 $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_322 N_A_129_179#_c_328_n N_A_721_99#_c_616_n 0.0135668f $X=3.56 $Y=1.68 $X2=0
+ $Y2=0
cc_323 N_A_129_179#_c_303_n N_A_593_125#_M1023_g 0.00285417f $X=4.34 $Y=1.125
+ $X2=0 $Y2=0
cc_324 N_A_129_179#_c_304_n N_A_593_125#_M1023_g 0.00838885f $X=4.975 $Y=0.617
+ $X2=0 $Y2=0
cc_325 N_A_129_179#_c_306_n N_A_593_125#_M1023_g 0.00843012f $X=5.06 $Y=1.165
+ $X2=0 $Y2=0
cc_326 N_A_129_179#_c_308_n N_A_593_125#_M1023_g 0.00319947f $X=5.145 $Y=1.25
+ $X2=0 $Y2=0
cc_327 N_A_129_179#_c_304_n N_A_593_125#_c_703_n 7.76621e-19 $X=4.975 $Y=0.617
+ $X2=0 $Y2=0
cc_328 N_A_129_179#_c_307_n N_A_593_125#_c_703_n 0.0154992f $X=6.025 $Y=1.25
+ $X2=0 $Y2=0
cc_329 N_A_129_179#_c_314_n N_A_593_125#_c_703_n 0.00226804f $X=6.11 $Y=1.25
+ $X2=0 $Y2=0
cc_330 N_A_129_179#_c_307_n N_A_593_125#_c_704_n 0.00400694f $X=6.025 $Y=1.25
+ $X2=0 $Y2=0
cc_331 N_A_129_179#_c_309_n N_A_593_125#_c_704_n 0.00474552f $X=6.65 $Y=1.44
+ $X2=0 $Y2=0
cc_332 N_A_129_179#_c_314_n N_A_593_125#_c_704_n 0.0104093f $X=6.11 $Y=1.25
+ $X2=0 $Y2=0
cc_333 N_A_129_179#_c_316_n N_A_593_125#_c_704_n 0.00475896f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_334 N_A_129_179#_c_293_n N_A_593_125#_c_706_n 0.00475896f $X=6.815 $Y=1.86
+ $X2=0 $Y2=0
cc_335 N_A_129_179#_c_315_n N_A_593_125#_c_706_n 0.0010135f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_336 N_A_129_179#_c_325_n N_A_593_125#_M1010_g 0.0465421f $X=6.815 $Y=2.025
+ $X2=0 $Y2=0
cc_337 N_A_129_179#_M1033_g N_A_593_125#_c_708_n 0.00467152f $X=2.89 $Y=0.835
+ $X2=0 $Y2=0
cc_338 N_A_129_179#_c_290_n N_A_593_125#_c_708_n 0.0170136f $X=3.245 $Y=1.49
+ $X2=0 $Y2=0
cc_339 N_A_129_179#_c_300_n N_A_593_125#_c_708_n 0.00892024f $X=3.555 $Y=1.125
+ $X2=0 $Y2=0
cc_340 N_A_129_179#_c_301_n N_A_593_125#_c_708_n 0.0642533f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_341 N_A_129_179#_c_328_n N_A_593_125#_c_708_n 0.00939992f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_342 N_A_129_179#_c_313_n N_A_593_125#_c_708_n 0.0142228f $X=3.56 $Y=1.21
+ $X2=0 $Y2=0
cc_343 N_A_129_179#_M1028_g N_A_593_125#_c_718_n 0.00993759f $X=3.43 $Y=2.885
+ $X2=0 $Y2=0
cc_344 N_A_129_179#_M1028_g N_A_593_125#_c_719_n 0.0113241f $X=3.43 $Y=2.885
+ $X2=0 $Y2=0
cc_345 N_A_129_179#_c_323_n N_A_593_125#_c_719_n 0.00371302f $X=3.54 $Y=2.185
+ $X2=0 $Y2=0
cc_346 N_A_129_179#_c_301_n N_A_593_125#_c_719_n 0.0142377f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_347 N_A_129_179#_M1028_g N_A_593_125#_c_720_n 0.0016665f $X=3.43 $Y=2.885
+ $X2=0 $Y2=0
cc_348 N_A_129_179#_c_301_n N_A_593_125#_c_720_n 0.0143484f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_349 N_A_129_179#_c_328_n N_A_593_125#_c_720_n 0.00169928f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_350 N_A_129_179#_c_301_n N_A_593_125#_c_722_n 0.0138148f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_351 N_A_129_179#_c_328_n N_A_593_125#_c_722_n 0.00162093f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_352 N_A_129_179#_c_302_n N_A_593_125#_c_722_n 0.00491785f $X=4.255 $Y=1.21
+ $X2=0 $Y2=0
cc_353 N_A_129_179#_c_307_n N_A_593_125#_c_709_n 0.0387059f $X=6.025 $Y=1.25
+ $X2=0 $Y2=0
cc_354 N_A_129_179#_c_308_n N_A_593_125#_c_710_n 0.0158834f $X=5.145 $Y=1.25
+ $X2=0 $Y2=0
cc_355 N_A_129_179#_c_293_n N_A_593_125#_c_724_n 0.0010902f $X=6.815 $Y=1.86
+ $X2=0 $Y2=0
cc_356 N_A_129_179#_c_307_n N_A_593_125#_c_724_n 0.00822994f $X=6.025 $Y=1.25
+ $X2=0 $Y2=0
cc_357 N_A_129_179#_c_309_n N_A_593_125#_c_724_n 0.0153454f $X=6.65 $Y=1.44
+ $X2=0 $Y2=0
cc_358 N_A_129_179#_c_314_n N_A_593_125#_c_724_n 0.0123692f $X=6.11 $Y=1.25
+ $X2=0 $Y2=0
cc_359 N_A_129_179#_c_315_n N_A_593_125#_c_724_n 0.0186662f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_360 N_A_129_179#_c_290_n N_A_593_125#_c_767_n 0.00354088f $X=3.245 $Y=1.49
+ $X2=0 $Y2=0
cc_361 N_A_129_179#_c_298_n N_A_593_125#_c_767_n 0.0140831f $X=3.465 $Y=0.34
+ $X2=0 $Y2=0
cc_362 N_A_129_179#_c_300_n N_A_593_125#_c_767_n 0.0243265f $X=3.555 $Y=1.125
+ $X2=0 $Y2=0
cc_363 N_A_129_179#_c_290_n N_A_593_125#_c_725_n 0.00149275f $X=3.245 $Y=1.49
+ $X2=0 $Y2=0
cc_364 N_A_129_179#_M1028_g N_A_593_125#_c_725_n 0.00305188f $X=3.43 $Y=2.885
+ $X2=0 $Y2=0
cc_365 N_A_129_179#_c_307_n N_A_593_125#_c_711_n 0.0128514f $X=6.025 $Y=1.25
+ $X2=0 $Y2=0
cc_366 N_A_129_179#_c_314_n N_A_593_125#_c_711_n 0.00129487f $X=6.11 $Y=1.25
+ $X2=0 $Y2=0
cc_367 N_A_129_179#_c_293_n N_A_593_125#_c_729_n 0.0465421f $X=6.815 $Y=1.86
+ $X2=0 $Y2=0
cc_368 N_A_129_179#_c_309_n N_A_593_125#_c_729_n 0.00570931f $X=6.65 $Y=1.44
+ $X2=0 $Y2=0
cc_369 N_A_129_179#_c_315_n N_A_593_125#_c_729_n 0.00116243f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_370 N_A_129_179#_c_306_n N_SET_B_M1022_g 0.00199816f $X=5.06 $Y=1.165 $X2=0
+ $Y2=0
cc_371 N_A_129_179#_c_307_n N_SET_B_M1022_g 0.0145974f $X=6.025 $Y=1.25 $X2=0
+ $Y2=0
cc_372 N_A_129_179#_c_314_n N_SET_B_M1022_g 4.55586e-19 $X=6.11 $Y=1.25 $X2=0
+ $Y2=0
cc_373 N_A_129_179#_c_307_n N_SET_B_c_883_n 3.56767e-19 $X=6.025 $Y=1.25 $X2=0
+ $Y2=0
cc_374 N_A_129_179#_M1009_g N_SET_B_c_886_n 0.015393f $X=6.725 $Y=2.675 $X2=0
+ $Y2=0
cc_375 N_A_129_179#_M1009_g N_SET_B_c_887_n 0.002224f $X=6.725 $Y=2.675 $X2=0
+ $Y2=0
cc_376 N_A_129_179#_M1009_g N_SET_B_c_890_n 0.0014208f $X=6.725 $Y=2.675 $X2=0
+ $Y2=0
cc_377 N_A_129_179#_c_295_n N_A_191_21#_M1036_s 0.00212773f $X=1.44 $Y=1.25
+ $X2=-0.19 $Y2=-0.245
cc_378 N_A_129_179#_c_312_n N_A_191_21#_M1036_s 3.07096e-19 $X=1.675 $Y=1.25
+ $X2=-0.19 $Y2=-0.245
cc_379 N_A_129_179#_c_295_n N_A_191_21#_c_994_n 0.0266023f $X=1.44 $Y=1.25 $X2=0
+ $Y2=0
cc_380 N_A_129_179#_c_310_n N_A_191_21#_c_994_n 0.00950992f $X=0.82 $Y=2.29
+ $X2=0 $Y2=0
cc_381 N_A_129_179#_c_311_n N_A_191_21#_c_994_n 0.0213315f $X=1.51 $Y=1.32 $X2=0
+ $Y2=0
cc_382 N_A_129_179#_c_317_n N_A_191_21#_c_994_n 0.0148371f $X=1.51 $Y=1.155
+ $X2=0 $Y2=0
cc_383 N_A_129_179#_M1033_g N_A_191_21#_c_995_n 0.00737859f $X=2.89 $Y=0.835
+ $X2=0 $Y2=0
cc_384 N_A_129_179#_c_298_n N_A_191_21#_c_995_n 0.0130282f $X=3.465 $Y=0.34
+ $X2=0 $Y2=0
cc_385 N_A_129_179#_c_299_n N_A_191_21#_c_995_n 0.0037969f $X=2.41 $Y=0.34 $X2=0
+ $Y2=0
cc_386 N_A_129_179#_c_317_n N_A_191_21#_c_995_n 0.00894172f $X=1.51 $Y=1.155
+ $X2=0 $Y2=0
cc_387 N_A_129_179#_c_319_n N_A_191_21#_c_1003_n 0.010543f $X=1.86 $Y=3.075
+ $X2=0 $Y2=0
cc_388 N_A_129_179#_c_291_n N_A_191_21#_c_1003_n 0.0121548f $X=2.965 $Y=1.49
+ $X2=0 $Y2=0
cc_389 N_A_129_179#_c_296_n N_A_191_21#_c_1003_n 0.00514576f $X=2.24 $Y=1.105
+ $X2=0 $Y2=0
cc_390 N_A_129_179#_c_328_n N_A_191_21#_c_1003_n 0.0170459f $X=3.56 $Y=1.68
+ $X2=0 $Y2=0
cc_391 N_A_129_179#_c_311_n N_A_191_21#_c_1003_n 0.00544528f $X=1.51 $Y=1.32
+ $X2=0 $Y2=0
cc_392 N_A_129_179#_c_312_n N_A_191_21#_c_1003_n 7.72495e-19 $X=1.675 $Y=1.25
+ $X2=0 $Y2=0
cc_393 N_A_129_179#_c_295_n N_A_191_21#_c_1004_n 0.00666461f $X=1.44 $Y=1.25
+ $X2=0 $Y2=0
cc_394 N_A_129_179#_c_310_n N_A_191_21#_c_1004_n 0.0017546f $X=0.82 $Y=2.29
+ $X2=0 $Y2=0
cc_395 N_A_129_179#_c_311_n N_A_191_21#_c_1004_n 0.0106046f $X=1.51 $Y=1.32
+ $X2=0 $Y2=0
cc_396 N_A_129_179#_c_323_n N_A_191_21#_M1037_g 0.0170459f $X=3.54 $Y=2.185
+ $X2=0 $Y2=0
cc_397 N_A_129_179#_M1033_g N_A_191_21#_M1021_g 0.0126054f $X=2.89 $Y=0.835
+ $X2=0 $Y2=0
cc_398 N_A_129_179#_c_290_n N_A_191_21#_M1021_g 0.00984703f $X=3.245 $Y=1.49
+ $X2=0 $Y2=0
cc_399 N_A_129_179#_c_298_n N_A_191_21#_M1021_g 0.0161928f $X=3.465 $Y=0.34
+ $X2=0 $Y2=0
cc_400 N_A_129_179#_c_300_n N_A_191_21#_M1021_g 0.00933004f $X=3.555 $Y=1.125
+ $X2=0 $Y2=0
cc_401 N_A_129_179#_c_313_n N_A_191_21#_M1021_g 3.44891e-19 $X=3.56 $Y=1.21
+ $X2=0 $Y2=0
cc_402 N_A_129_179#_M1020_g N_A_191_21#_c_997_n 0.00350215f $X=6.74 $Y=1.005
+ $X2=0 $Y2=0
cc_403 N_A_129_179#_c_298_n N_A_191_21#_c_997_n 0.00483986f $X=3.465 $Y=0.34
+ $X2=0 $Y2=0
cc_404 N_A_129_179#_c_304_n N_A_191_21#_c_997_n 0.012816f $X=4.975 $Y=0.617
+ $X2=0 $Y2=0
cc_405 N_A_129_179#_c_305_n N_A_191_21#_c_997_n 0.00361151f $X=4.425 $Y=0.617
+ $X2=0 $Y2=0
cc_406 N_A_129_179#_M1009_g N_A_191_21#_M1026_g 0.0159033f $X=6.725 $Y=2.675
+ $X2=0 $Y2=0
cc_407 N_A_129_179#_M1020_g N_A_191_21#_M1026_g 0.0105048f $X=6.74 $Y=1.005
+ $X2=0 $Y2=0
cc_408 N_A_129_179#_c_315_n N_A_191_21#_M1026_g 4.57845e-19 $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_409 N_A_129_179#_c_316_n N_A_191_21#_M1026_g 0.0412676f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_410 N_A_129_179#_c_295_n N_A_191_21#_c_1000_n 0.0457443f $X=1.44 $Y=1.25
+ $X2=0 $Y2=0
cc_411 N_A_129_179#_c_311_n N_A_191_21#_c_1000_n 8.85732e-19 $X=1.51 $Y=1.32
+ $X2=0 $Y2=0
cc_412 N_A_129_179#_c_317_n N_A_191_21#_c_1000_n 0.00625578f $X=1.51 $Y=1.155
+ $X2=0 $Y2=0
cc_413 N_A_129_179#_c_319_n N_A_191_21#_c_1007_n 0.00221658f $X=1.86 $Y=3.075
+ $X2=0 $Y2=0
cc_414 N_A_129_179#_c_295_n N_A_191_21#_c_1007_n 0.0163261f $X=1.44 $Y=1.25
+ $X2=0 $Y2=0
cc_415 N_A_129_179#_c_310_n N_A_191_21#_c_1007_n 0.0286688f $X=0.82 $Y=2.29
+ $X2=0 $Y2=0
cc_416 N_A_129_179#_c_311_n N_A_191_21#_c_1007_n 6.5784e-19 $X=1.51 $Y=1.32
+ $X2=0 $Y2=0
cc_417 N_A_129_179#_c_318_n N_A_191_21#_c_1008_n 0.00881577f $X=1.785 $Y=3.15
+ $X2=0 $Y2=0
cc_418 N_A_129_179#_c_319_n N_A_191_21#_c_1008_n 4.3695e-19 $X=1.86 $Y=3.075
+ $X2=0 $Y2=0
cc_419 N_A_129_179#_c_329_n N_A_191_21#_c_1008_n 0.0214136f $X=0.785 $Y=2.455
+ $X2=0 $Y2=0
cc_420 N_A_129_179#_c_331_n N_A_191_21#_c_1008_n 0.0114897f $X=1.05 $Y=2.94
+ $X2=0 $Y2=0
cc_421 N_A_129_179#_c_332_n N_A_191_21#_c_1008_n 8.487e-19 $X=1.05 $Y=2.94 $X2=0
+ $Y2=0
cc_422 N_A_129_179#_c_295_n N_A_191_21#_c_1001_n 6.73946e-19 $X=1.44 $Y=1.25
+ $X2=0 $Y2=0
cc_423 N_A_129_179#_c_317_n N_A_191_21#_c_1001_n 0.00109563f $X=1.51 $Y=1.155
+ $X2=0 $Y2=0
cc_424 N_A_129_179#_M1020_g N_A_1360_451#_c_1224_n 0.00332074f $X=6.74 $Y=1.005
+ $X2=0 $Y2=0
cc_425 N_A_129_179#_c_315_n N_A_1360_451#_c_1224_n 0.00397349f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_426 N_A_129_179#_c_316_n N_A_1360_451#_c_1224_n 3.00531e-19 $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_427 N_A_129_179#_M1009_g N_A_1360_451#_c_1225_n 0.00484065f $X=6.725 $Y=2.675
+ $X2=0 $Y2=0
cc_428 N_A_129_179#_c_293_n N_A_1360_451#_c_1225_n 0.00266675f $X=6.815 $Y=1.86
+ $X2=0 $Y2=0
cc_429 N_A_129_179#_c_315_n N_A_1360_451#_c_1225_n 0.0323999f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_430 N_A_129_179#_M1009_g N_A_1360_451#_c_1238_n 0.00363344f $X=6.725 $Y=2.675
+ $X2=0 $Y2=0
cc_431 N_A_129_179#_c_325_n N_A_1360_451#_c_1238_n 0.00298915f $X=6.815 $Y=2.025
+ $X2=0 $Y2=0
cc_432 N_A_129_179#_c_315_n N_A_1360_451#_c_1238_n 0.00415428f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_433 N_A_129_179#_c_315_n N_A_1360_451#_c_1249_n 0.00437103f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_434 N_A_129_179#_c_316_n N_A_1360_451#_c_1249_n 0.00332863f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_435 N_A_129_179#_c_315_n N_A_1360_451#_c_1229_n 0.0156355f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_436 N_A_129_179#_c_316_n N_A_1360_451#_c_1229_n 0.00126599f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_437 N_A_129_179#_c_326_n N_VPWR_c_1421_n 0.00996365f $X=0.835 $Y=2.775 $X2=0
+ $Y2=0
cc_438 N_A_129_179#_c_329_n N_VPWR_c_1421_n 0.0133194f $X=0.785 $Y=2.455 $X2=0
+ $Y2=0
cc_439 N_A_129_179#_c_331_n N_VPWR_c_1421_n 0.0229244f $X=1.05 $Y=2.94 $X2=0
+ $Y2=0
cc_440 N_A_129_179#_c_332_n N_VPWR_c_1421_n 0.00496991f $X=1.05 $Y=2.94 $X2=0
+ $Y2=0
cc_441 N_A_129_179#_c_319_n N_VPWR_c_1422_n 0.00971978f $X=1.86 $Y=3.075 $X2=0
+ $Y2=0
cc_442 N_A_129_179#_c_329_n N_VPWR_c_1430_n 4.8884e-19 $X=0.785 $Y=2.455 $X2=0
+ $Y2=0
cc_443 N_A_129_179#_c_331_n N_VPWR_c_1430_n 0.0321165f $X=1.05 $Y=2.94 $X2=0
+ $Y2=0
cc_444 N_A_129_179#_c_332_n N_VPWR_c_1430_n 0.0304409f $X=1.05 $Y=2.94 $X2=0
+ $Y2=0
cc_445 N_A_129_179#_M1009_g N_VPWR_c_1432_n 0.00357877f $X=6.725 $Y=2.675 $X2=0
+ $Y2=0
cc_446 N_A_129_179#_M1028_g N_VPWR_c_1438_n 0.00557327f $X=3.43 $Y=2.885 $X2=0
+ $Y2=0
cc_447 N_A_129_179#_M1028_g N_VPWR_c_1439_n 0.00202503f $X=3.43 $Y=2.885 $X2=0
+ $Y2=0
cc_448 N_A_129_179#_c_318_n N_VPWR_c_1419_n 0.0269116f $X=1.785 $Y=3.15 $X2=0
+ $Y2=0
cc_449 N_A_129_179#_M1028_g N_VPWR_c_1419_n 0.00624007f $X=3.43 $Y=2.885 $X2=0
+ $Y2=0
cc_450 N_A_129_179#_M1009_g N_VPWR_c_1419_n 0.00665366f $X=6.725 $Y=2.675 $X2=0
+ $Y2=0
cc_451 N_A_129_179#_c_329_n N_VPWR_c_1419_n 8.12108e-19 $X=0.785 $Y=2.455 $X2=0
+ $Y2=0
cc_452 N_A_129_179#_c_331_n N_VPWR_c_1419_n 0.0173353f $X=1.05 $Y=2.94 $X2=0
+ $Y2=0
cc_453 N_A_129_179#_c_332_n N_VPWR_c_1419_n 0.0101219f $X=1.05 $Y=2.94 $X2=0
+ $Y2=0
cc_454 N_A_129_179#_M1033_g N_A_507_125#_c_1573_n 0.00233192f $X=2.89 $Y=0.835
+ $X2=0 $Y2=0
cc_455 N_A_129_179#_c_296_n N_A_507_125#_c_1573_n 0.0134955f $X=2.24 $Y=1.105
+ $X2=0 $Y2=0
cc_456 N_A_129_179#_c_298_n N_A_507_125#_c_1573_n 0.0113353f $X=3.465 $Y=0.34
+ $X2=0 $Y2=0
cc_457 N_A_129_179#_c_290_n N_A_507_125#_c_1574_n 5.09075e-19 $X=3.245 $Y=1.49
+ $X2=0 $Y2=0
cc_458 N_A_129_179#_c_291_n N_A_507_125#_c_1574_n 0.00647846f $X=2.965 $Y=1.49
+ $X2=0 $Y2=0
cc_459 N_A_129_179#_M1028_g N_A_507_125#_c_1574_n 2.57031e-19 $X=3.43 $Y=2.885
+ $X2=0 $Y2=0
cc_460 N_A_129_179#_M1033_g N_A_507_125#_c_1575_n 0.009724f $X=2.89 $Y=0.835
+ $X2=0 $Y2=0
cc_461 N_A_129_179#_c_291_n N_A_507_125#_c_1575_n 0.00106526f $X=2.965 $Y=1.49
+ $X2=0 $Y2=0
cc_462 N_A_129_179#_c_296_n N_VGND_M1036_d 0.0109597f $X=2.24 $Y=1.105 $X2=0
+ $Y2=0
cc_463 N_A_129_179#_c_297_n N_VGND_M1036_d 0.00492505f $X=2.325 $Y=1.015 $X2=0
+ $Y2=0
cc_464 N_A_129_179#_c_307_n N_VGND_M1022_d 0.00324203f $X=6.025 $Y=1.25 $X2=0
+ $Y2=0
cc_465 N_A_129_179#_c_296_n N_VGND_c_1650_n 0.026707f $X=2.24 $Y=1.105 $X2=0
+ $Y2=0
cc_466 N_A_129_179#_c_297_n N_VGND_c_1650_n 0.0313073f $X=2.325 $Y=1.015 $X2=0
+ $Y2=0
cc_467 N_A_129_179#_c_299_n N_VGND_c_1650_n 0.0144411f $X=2.41 $Y=0.34 $X2=0
+ $Y2=0
cc_468 N_A_129_179#_c_317_n N_VGND_c_1650_n 0.00357032f $X=1.51 $Y=1.155 $X2=0
+ $Y2=0
cc_469 N_A_129_179#_c_298_n N_VGND_c_1651_n 0.0147862f $X=3.465 $Y=0.34 $X2=0
+ $Y2=0
cc_470 N_A_129_179#_c_300_n N_VGND_c_1651_n 0.0391467f $X=3.555 $Y=1.125 $X2=0
+ $Y2=0
cc_471 N_A_129_179#_c_302_n N_VGND_c_1651_n 0.0213336f $X=4.255 $Y=1.21 $X2=0
+ $Y2=0
cc_472 N_A_129_179#_c_303_n N_VGND_c_1651_n 0.0171789f $X=4.34 $Y=1.125 $X2=0
+ $Y2=0
cc_473 N_A_129_179#_c_305_n N_VGND_c_1651_n 0.0169818f $X=4.425 $Y=0.617 $X2=0
+ $Y2=0
cc_474 N_A_129_179#_c_304_n N_VGND_c_1652_n 0.0132958f $X=4.975 $Y=0.617 $X2=0
+ $Y2=0
cc_475 N_A_129_179#_c_306_n N_VGND_c_1652_n 0.0115452f $X=5.06 $Y=1.165 $X2=0
+ $Y2=0
cc_476 N_A_129_179#_c_307_n N_VGND_c_1652_n 0.0218816f $X=6.025 $Y=1.25 $X2=0
+ $Y2=0
cc_477 N_A_129_179#_c_298_n N_VGND_c_1662_n 0.0797213f $X=3.465 $Y=0.34 $X2=0
+ $Y2=0
cc_478 N_A_129_179#_c_299_n N_VGND_c_1662_n 0.0115893f $X=2.41 $Y=0.34 $X2=0
+ $Y2=0
cc_479 N_A_129_179#_c_304_n N_VGND_c_1664_n 0.0178889f $X=4.975 $Y=0.617 $X2=0
+ $Y2=0
cc_480 N_A_129_179#_c_305_n N_VGND_c_1664_n 0.00451713f $X=4.425 $Y=0.617 $X2=0
+ $Y2=0
cc_481 N_A_129_179#_c_298_n N_VGND_c_1674_n 0.041484f $X=3.465 $Y=0.34 $X2=0
+ $Y2=0
cc_482 N_A_129_179#_c_299_n N_VGND_c_1674_n 0.00583135f $X=2.41 $Y=0.34 $X2=0
+ $Y2=0
cc_483 N_A_129_179#_c_304_n N_VGND_c_1674_n 0.0200966f $X=4.975 $Y=0.617 $X2=0
+ $Y2=0
cc_484 N_A_129_179#_c_305_n N_VGND_c_1674_n 0.00494968f $X=4.425 $Y=0.617 $X2=0
+ $Y2=0
cc_485 N_A_129_179#_c_317_n N_VGND_c_1674_n 7.97988e-19 $X=1.51 $Y=1.155 $X2=0
+ $Y2=0
cc_486 N_A_129_179#_c_300_n A_679_125# 0.00354114f $X=3.555 $Y=1.125 $X2=-0.19
+ $Y2=-0.245
cc_487 N_A_129_179#_c_307_n N_A_1173_125#_M1003_d 0.00137045f $X=6.025 $Y=1.25
+ $X2=-0.19 $Y2=-0.245
cc_488 N_A_129_179#_c_314_n N_A_1173_125#_M1003_d 0.00150852f $X=6.11 $Y=1.25
+ $X2=-0.19 $Y2=-0.245
cc_489 N_A_129_179#_M1020_g N_A_1173_125#_c_1795_n 5.34611e-19 $X=6.74 $Y=1.005
+ $X2=0 $Y2=0
cc_490 N_A_129_179#_c_307_n N_A_1173_125#_c_1795_n 0.00837991f $X=6.025 $Y=1.25
+ $X2=0 $Y2=0
cc_491 N_A_129_179#_c_314_n N_A_1173_125#_c_1795_n 0.0124422f $X=6.11 $Y=1.25
+ $X2=0 $Y2=0
cc_492 N_A_129_179#_M1020_g N_A_1173_125#_c_1797_n 5.0188e-19 $X=6.74 $Y=1.005
+ $X2=0 $Y2=0
cc_493 N_A_129_179#_c_309_n N_A_1280_159#_c_1822_n 0.0199761f $X=6.65 $Y=1.44
+ $X2=0 $Y2=0
cc_494 N_A_129_179#_c_314_n N_A_1280_159#_c_1822_n 3.93442e-19 $X=6.11 $Y=1.25
+ $X2=0 $Y2=0
cc_495 N_A_129_179#_M1020_g N_A_1280_159#_c_1823_n 0.00279758f $X=6.74 $Y=1.005
+ $X2=0 $Y2=0
cc_496 N_A_129_179#_M1020_g N_A_1280_159#_c_1825_n 0.00883891f $X=6.74 $Y=1.005
+ $X2=0 $Y2=0
cc_497 N_A_129_179#_c_315_n N_A_1280_159#_c_1825_n 0.00464538f $X=6.815 $Y=1.52
+ $X2=0 $Y2=0
cc_498 N_D_M1032_g N_A_191_21#_c_995_n 0.00752747f $X=2.46 $Y=0.835 $X2=0 $Y2=0
cc_499 D N_A_191_21#_c_1003_n 0.0342476f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_500 N_D_c_556_n N_A_191_21#_c_1003_n 0.029157f $X=2.08 $Y=1.45 $X2=0 $Y2=0
cc_501 N_D_c_559_n N_A_191_21#_c_1003_n 0.0218496f $X=2.51 $Y=2.35 $X2=0 $Y2=0
cc_502 D N_A_191_21#_c_1004_n 0.00512068f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_503 N_D_M1008_g N_A_191_21#_M1037_g 0.0149098f $X=2.53 $Y=2.885 $X2=0 $Y2=0
cc_504 D N_A_191_21#_M1037_g 0.00153212f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_505 N_D_c_559_n N_A_191_21#_M1037_g 0.0203401f $X=2.51 $Y=2.35 $X2=0 $Y2=0
cc_506 D N_A_191_21#_c_1007_n 0.0234922f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_507 D N_A_191_21#_c_1008_n 0.00792237f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_508 D N_VPWR_M1006_d 0.0031099f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_509 N_D_M1008_g N_VPWR_c_1422_n 0.00869842f $X=2.53 $Y=2.885 $X2=0 $Y2=0
cc_510 D N_VPWR_c_1422_n 0.0290203f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_511 N_D_M1008_g N_VPWR_c_1438_n 0.00585385f $X=2.53 $Y=2.885 $X2=0 $Y2=0
cc_512 N_D_M1008_g N_VPWR_c_1419_n 0.00732179f $X=2.53 $Y=2.885 $X2=0 $Y2=0
cc_513 D N_VPWR_c_1419_n 0.0138055f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_514 N_D_c_559_n N_VPWR_c_1419_n 8.0553e-19 $X=2.51 $Y=2.35 $X2=0 $Y2=0
cc_515 N_D_M1032_g N_A_507_125#_c_1573_n 0.00296197f $X=2.46 $Y=0.835 $X2=0
+ $Y2=0
cc_516 N_D_M1008_g N_A_507_125#_c_1574_n 0.00360993f $X=2.53 $Y=2.885 $X2=0
+ $Y2=0
cc_517 D N_A_507_125#_c_1574_n 0.0799506f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_518 N_D_c_556_n N_A_507_125#_c_1574_n 7.47818e-19 $X=2.08 $Y=1.45 $X2=0 $Y2=0
cc_519 N_D_c_559_n N_A_507_125#_c_1574_n 0.00205307f $X=2.51 $Y=2.35 $X2=0 $Y2=0
cc_520 N_D_M1032_g N_A_507_125#_c_1575_n 0.00374076f $X=2.46 $Y=0.835 $X2=0
+ $Y2=0
cc_521 D N_A_507_125#_c_1575_n 0.0046057f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_522 N_D_c_559_n N_A_507_125#_c_1592_n 9.60095e-19 $X=2.51 $Y=2.35 $X2=0 $Y2=0
cc_523 N_D_M1032_g N_VGND_c_1650_n 0.00114026f $X=2.46 $Y=0.835 $X2=0 $Y2=0
cc_524 N_A_721_99#_c_612_n N_A_593_125#_M1019_g 0.0133357f $X=4.845 $Y=2.58
+ $X2=0 $Y2=0
cc_525 N_A_721_99#_c_614_n N_A_593_125#_M1019_g 0.00238401f $X=4.995 $Y=2.58
+ $X2=0 $Y2=0
cc_526 N_A_721_99#_c_601_n N_A_593_125#_M1023_g 0.00607474f $X=3.965 $Y=1.23
+ $X2=0 $Y2=0
cc_527 N_A_721_99#_c_603_n N_A_593_125#_M1023_g 0.00259146f $X=4.595 $Y=1.555
+ $X2=0 $Y2=0
cc_528 N_A_721_99#_c_605_n N_A_593_125#_M1023_g 0.00452617f $X=4.69 $Y=1.055
+ $X2=0 $Y2=0
cc_529 N_A_721_99#_c_603_n N_A_593_125#_c_707_n 0.00718775f $X=4.595 $Y=1.555
+ $X2=0 $Y2=0
cc_530 N_A_721_99#_c_606_n N_A_593_125#_c_707_n 0.00426753f $X=4.13 $Y=1.715
+ $X2=0 $Y2=0
cc_531 N_A_721_99#_c_616_n N_A_593_125#_c_707_n 0.0140327f $X=4.26 $Y=2.185
+ $X2=0 $Y2=0
cc_532 N_A_721_99#_c_612_n N_A_593_125#_c_716_n 0.00131741f $X=4.845 $Y=2.58
+ $X2=0 $Y2=0
cc_533 N_A_721_99#_c_614_n N_A_593_125#_c_716_n 0.00404009f $X=4.995 $Y=2.58
+ $X2=0 $Y2=0
cc_534 N_A_721_99#_c_602_n N_A_593_125#_c_708_n 3.77146e-19 $X=3.755 $Y=1.23
+ $X2=0 $Y2=0
cc_535 N_A_721_99#_c_609_n N_A_593_125#_c_718_n 0.00206805f $X=3.865 $Y=2.47
+ $X2=0 $Y2=0
cc_536 N_A_721_99#_c_608_n N_A_593_125#_c_719_n 0.00768345f $X=4.095 $Y=2.47
+ $X2=0 $Y2=0
cc_537 N_A_721_99#_c_609_n N_A_593_125#_c_719_n 0.00903489f $X=3.865 $Y=2.47
+ $X2=0 $Y2=0
cc_538 N_A_721_99#_c_610_n N_A_593_125#_c_719_n 0.00956029f $X=4.26 $Y=2.35
+ $X2=0 $Y2=0
cc_539 N_A_721_99#_c_611_n N_A_593_125#_c_719_n 3.68444e-19 $X=4.26 $Y=2.35
+ $X2=0 $Y2=0
cc_540 N_A_721_99#_c_613_n N_A_593_125#_c_719_n 0.003229f $X=4.345 $Y=2.58 $X2=0
+ $Y2=0
cc_541 N_A_721_99#_c_610_n N_A_593_125#_c_720_n 0.0122958f $X=4.26 $Y=2.35 $X2=0
+ $Y2=0
cc_542 N_A_721_99#_c_616_n N_A_593_125#_c_720_n 0.00457678f $X=4.26 $Y=2.185
+ $X2=0 $Y2=0
cc_543 N_A_721_99#_c_608_n N_A_593_125#_c_721_n 0.00178804f $X=4.095 $Y=2.47
+ $X2=0 $Y2=0
cc_544 N_A_721_99#_c_603_n N_A_593_125#_c_721_n 0.0601718f $X=4.595 $Y=1.555
+ $X2=0 $Y2=0
cc_545 N_A_721_99#_c_610_n N_A_593_125#_c_721_n 0.0177346f $X=4.26 $Y=2.35 $X2=0
+ $Y2=0
cc_546 N_A_721_99#_c_611_n N_A_593_125#_c_721_n 0.00311711f $X=4.26 $Y=2.35
+ $X2=0 $Y2=0
cc_547 N_A_721_99#_c_612_n N_A_593_125#_c_721_n 0.0250067f $X=4.845 $Y=2.58
+ $X2=0 $Y2=0
cc_548 N_A_721_99#_c_614_n N_A_593_125#_c_721_n 0.026748f $X=4.995 $Y=2.58 $X2=0
+ $Y2=0
cc_549 N_A_721_99#_c_606_n N_A_593_125#_c_721_n 0.00185554f $X=4.13 $Y=1.715
+ $X2=0 $Y2=0
cc_550 N_A_721_99#_c_616_n N_A_593_125#_c_721_n 0.014303f $X=4.26 $Y=2.185 $X2=0
+ $Y2=0
cc_551 N_A_721_99#_c_601_n N_A_593_125#_c_722_n 0.00227501f $X=3.965 $Y=1.23
+ $X2=0 $Y2=0
cc_552 N_A_721_99#_c_603_n N_A_593_125#_c_722_n 0.00244137f $X=4.595 $Y=1.555
+ $X2=0 $Y2=0
cc_553 N_A_721_99#_c_606_n N_A_593_125#_c_722_n 4.28635e-19 $X=4.13 $Y=1.715
+ $X2=0 $Y2=0
cc_554 N_A_721_99#_c_603_n N_A_593_125#_c_710_n 0.0117515f $X=4.595 $Y=1.555
+ $X2=0 $Y2=0
cc_555 N_A_721_99#_c_600_n N_A_593_125#_c_767_n 2.7236e-19 $X=3.68 $Y=1.155
+ $X2=0 $Y2=0
cc_556 N_A_721_99#_c_610_n N_A_593_125#_c_727_n 0.0014158f $X=4.26 $Y=2.35 $X2=0
+ $Y2=0
cc_557 N_A_721_99#_c_611_n N_A_593_125#_c_727_n 0.0219164f $X=4.26 $Y=2.35 $X2=0
+ $Y2=0
cc_558 N_A_721_99#_c_614_n N_SET_B_M1017_g 0.00488417f $X=4.995 $Y=2.58 $X2=0
+ $Y2=0
cc_559 N_A_721_99#_c_678_p N_SET_B_c_882_n 0.00451478f $X=5.625 $Y=2.885 $X2=0
+ $Y2=0
cc_560 N_A_721_99#_c_678_p N_SET_B_c_883_n 3.45206e-19 $X=5.625 $Y=2.885 $X2=0
+ $Y2=0
cc_561 N_A_721_99#_c_678_p N_SET_B_c_884_n 0.0125312f $X=5.625 $Y=2.885 $X2=0
+ $Y2=0
cc_562 N_A_721_99#_c_678_p N_SET_B_c_890_n 0.013142f $X=5.625 $Y=2.885 $X2=0
+ $Y2=0
cc_563 N_A_721_99#_c_600_n N_A_191_21#_M1021_g 0.0395734f $X=3.68 $Y=1.155 $X2=0
+ $Y2=0
cc_564 N_A_721_99#_c_600_n N_A_191_21#_c_997_n 0.00885751f $X=3.68 $Y=1.155
+ $X2=0 $Y2=0
cc_565 N_A_721_99#_c_612_n N_VPWR_c_1431_n 0.00266742f $X=4.845 $Y=2.58 $X2=0
+ $Y2=0
cc_566 N_A_721_99#_c_678_p N_VPWR_c_1431_n 0.0383048f $X=5.625 $Y=2.885 $X2=0
+ $Y2=0
cc_567 N_A_721_99#_c_614_n N_VPWR_c_1431_n 0.0203369f $X=4.995 $Y=2.58 $X2=0
+ $Y2=0
cc_568 N_A_721_99#_M1031_g N_VPWR_c_1438_n 0.00486043f $X=3.79 $Y=2.885 $X2=0
+ $Y2=0
cc_569 N_A_721_99#_M1031_g N_VPWR_c_1439_n 0.0111655f $X=3.79 $Y=2.885 $X2=0
+ $Y2=0
cc_570 N_A_721_99#_c_608_n N_VPWR_c_1439_n 0.00900995f $X=4.095 $Y=2.47 $X2=0
+ $Y2=0
cc_571 N_A_721_99#_c_611_n N_VPWR_c_1439_n 0.00145126f $X=4.26 $Y=2.35 $X2=0
+ $Y2=0
cc_572 N_A_721_99#_c_612_n N_VPWR_c_1439_n 0.0229397f $X=4.845 $Y=2.58 $X2=0
+ $Y2=0
cc_573 N_A_721_99#_c_613_n N_VPWR_c_1439_n 0.0142803f $X=4.345 $Y=2.58 $X2=0
+ $Y2=0
cc_574 N_A_721_99#_M1019_d N_VPWR_c_1419_n 0.00836111f $X=4.8 $Y=2.675 $X2=0
+ $Y2=0
cc_575 N_A_721_99#_M1031_g N_VPWR_c_1419_n 0.00433829f $X=3.79 $Y=2.885 $X2=0
+ $Y2=0
cc_576 N_A_721_99#_c_612_n N_VPWR_c_1419_n 0.0055126f $X=4.845 $Y=2.58 $X2=0
+ $Y2=0
cc_577 N_A_721_99#_c_613_n N_VPWR_c_1419_n 7.94568e-19 $X=4.345 $Y=2.58 $X2=0
+ $Y2=0
cc_578 N_A_721_99#_c_678_p N_VPWR_c_1419_n 0.0223617f $X=5.625 $Y=2.885 $X2=0
+ $Y2=0
cc_579 N_A_721_99#_c_614_n N_VPWR_c_1419_n 0.0115376f $X=4.995 $Y=2.58 $X2=0
+ $Y2=0
cc_580 N_A_721_99#_c_600_n N_VGND_c_1651_n 0.00387122f $X=3.68 $Y=1.155 $X2=0
+ $Y2=0
cc_581 N_A_721_99#_c_601_n N_VGND_c_1651_n 0.00188648f $X=3.965 $Y=1.23 $X2=0
+ $Y2=0
cc_582 N_A_721_99#_c_600_n N_VGND_c_1674_n 6.99321e-19 $X=3.68 $Y=1.155 $X2=0
+ $Y2=0
cc_583 N_A_593_125#_M1023_g N_SET_B_M1022_g 0.0449202f $X=4.905 $Y=1.055 $X2=0
+ $Y2=0
cc_584 N_A_593_125#_c_703_n N_SET_B_M1022_g 0.0202577f $X=5.79 $Y=1.375 $X2=0
+ $Y2=0
cc_585 N_A_593_125#_c_709_n N_SET_B_M1022_g 0.0148444f $X=5.675 $Y=1.59 $X2=0
+ $Y2=0
cc_586 N_A_593_125#_c_726_n N_SET_B_M1022_g 0.00231085f $X=4.897 $Y=1.815 $X2=0
+ $Y2=0
cc_587 N_A_593_125#_c_711_n N_SET_B_M1022_g 0.00366407f $X=5.76 $Y=1.59 $X2=0
+ $Y2=0
cc_588 N_A_593_125#_c_705_n N_SET_B_c_877_n 0.00502007f $X=5.865 $Y=1.45 $X2=0
+ $Y2=0
cc_589 N_A_593_125#_M1010_g N_SET_B_c_877_n 0.0302471f $X=6.365 $Y=2.675 $X2=0
+ $Y2=0
cc_590 N_A_593_125#_c_721_n N_SET_B_c_877_n 2.98074e-19 $X=4.65 $Y=1.9 $X2=0
+ $Y2=0
cc_591 N_A_593_125#_c_724_n N_SET_B_c_877_n 0.00150423f $X=6.245 $Y=1.87 $X2=0
+ $Y2=0
cc_592 N_A_593_125#_c_727_n N_SET_B_c_877_n 0.00224731f $X=4.815 $Y=1.9 $X2=0
+ $Y2=0
cc_593 N_A_593_125#_c_711_n N_SET_B_c_877_n 0.00795516f $X=5.76 $Y=1.59 $X2=0
+ $Y2=0
cc_594 N_A_593_125#_c_729_n N_SET_B_c_877_n 0.0107833f $X=6.365 $Y=1.87 $X2=0
+ $Y2=0
cc_595 N_A_593_125#_c_707_n N_SET_B_c_882_n 0.0449202f $X=4.815 $Y=1.77 $X2=0
+ $Y2=0
cc_596 N_A_593_125#_c_721_n N_SET_B_c_882_n 0.00231085f $X=4.65 $Y=1.9 $X2=0
+ $Y2=0
cc_597 N_A_593_125#_c_709_n N_SET_B_c_883_n 0.00563519f $X=5.675 $Y=1.59 $X2=0
+ $Y2=0
cc_598 N_A_593_125#_c_711_n N_SET_B_c_883_n 0.0033956f $X=5.76 $Y=1.59 $X2=0
+ $Y2=0
cc_599 N_A_593_125#_M1019_g N_SET_B_c_884_n 0.00213647f $X=4.725 $Y=2.885 $X2=0
+ $Y2=0
cc_600 N_A_593_125#_c_716_n N_SET_B_c_884_n 0.00241352f $X=4.815 $Y=2.415 $X2=0
+ $Y2=0
cc_601 N_A_593_125#_c_721_n N_SET_B_c_884_n 0.0109318f $X=4.65 $Y=1.9 $X2=0
+ $Y2=0
cc_602 N_A_593_125#_c_727_n N_SET_B_c_884_n 4.10171e-19 $X=4.815 $Y=1.9 $X2=0
+ $Y2=0
cc_603 N_A_593_125#_c_721_n N_SET_B_c_885_n 0.0284124f $X=4.65 $Y=1.9 $X2=0
+ $Y2=0
cc_604 N_A_593_125#_c_709_n N_SET_B_c_885_n 0.0148292f $X=5.675 $Y=1.59 $X2=0
+ $Y2=0
cc_605 N_A_593_125#_c_727_n N_SET_B_c_885_n 3.36314e-19 $X=4.815 $Y=1.9 $X2=0
+ $Y2=0
cc_606 N_A_593_125#_c_711_n N_SET_B_c_885_n 0.0129894f $X=5.76 $Y=1.59 $X2=0
+ $Y2=0
cc_607 N_A_593_125#_M1010_g N_SET_B_c_928_n 0.00752983f $X=6.365 $Y=2.675 $X2=0
+ $Y2=0
cc_608 N_A_593_125#_M1010_g N_SET_B_c_929_n 0.00309817f $X=6.365 $Y=2.675 $X2=0
+ $Y2=0
cc_609 N_A_593_125#_M1010_g N_SET_B_c_890_n 0.0166066f $X=6.365 $Y=2.675 $X2=0
+ $Y2=0
cc_610 N_A_593_125#_c_709_n N_SET_B_c_890_n 0.00597811f $X=5.675 $Y=1.59 $X2=0
+ $Y2=0
cc_611 N_A_593_125#_c_724_n N_SET_B_c_890_n 0.0446859f $X=6.245 $Y=1.87 $X2=0
+ $Y2=0
cc_612 N_A_593_125#_c_711_n N_SET_B_c_890_n 0.013042f $X=5.76 $Y=1.59 $X2=0
+ $Y2=0
cc_613 N_A_593_125#_c_729_n N_SET_B_c_890_n 0.00528626f $X=6.365 $Y=1.87 $X2=0
+ $Y2=0
cc_614 N_A_593_125#_c_708_n N_A_191_21#_c_1003_n 0.00415203f $X=3.205 $Y=2.365
+ $X2=0 $Y2=0
cc_615 N_A_593_125#_c_718_n N_A_191_21#_M1037_g 0.00254874f $X=3.21 $Y=2.88
+ $X2=0 $Y2=0
cc_616 N_A_593_125#_c_725_n N_A_191_21#_M1037_g 0.00138805f $X=3.245 $Y=2.45
+ $X2=0 $Y2=0
cc_617 N_A_593_125#_c_708_n N_A_191_21#_M1021_g 0.00371794f $X=3.205 $Y=2.365
+ $X2=0 $Y2=0
cc_618 N_A_593_125#_c_767_n N_A_191_21#_M1021_g 0.00481844f $X=3.205 $Y=0.835
+ $X2=0 $Y2=0
cc_619 N_A_593_125#_M1023_g N_A_191_21#_c_997_n 0.00305421f $X=4.905 $Y=1.055
+ $X2=0 $Y2=0
cc_620 N_A_593_125#_c_703_n N_A_191_21#_c_997_n 0.00894529f $X=5.79 $Y=1.375
+ $X2=0 $Y2=0
cc_621 N_A_593_125#_c_724_n N_A_1360_451#_c_1225_n 2.45002e-19 $X=6.245 $Y=1.87
+ $X2=0 $Y2=0
cc_622 N_A_593_125#_M1010_g N_A_1360_451#_c_1238_n 2.51316e-19 $X=6.365 $Y=2.675
+ $X2=0 $Y2=0
cc_623 N_A_593_125#_M1010_g N_VPWR_c_1423_n 0.00360226f $X=6.365 $Y=2.675 $X2=0
+ $Y2=0
cc_624 N_A_593_125#_M1019_g N_VPWR_c_1431_n 0.0035715f $X=4.725 $Y=2.885 $X2=0
+ $Y2=0
cc_625 N_A_593_125#_M1010_g N_VPWR_c_1432_n 0.00577794f $X=6.365 $Y=2.675 $X2=0
+ $Y2=0
cc_626 N_A_593_125#_c_718_n N_VPWR_c_1438_n 0.0134961f $X=3.21 $Y=2.88 $X2=0
+ $Y2=0
cc_627 N_A_593_125#_M1019_g N_VPWR_c_1439_n 0.00995557f $X=4.725 $Y=2.885 $X2=0
+ $Y2=0
cc_628 N_A_593_125#_c_718_n N_VPWR_c_1439_n 0.00722348f $X=3.21 $Y=2.88 $X2=0
+ $Y2=0
cc_629 N_A_593_125#_c_719_n N_VPWR_c_1439_n 0.00604969f $X=3.825 $Y=2.45 $X2=0
+ $Y2=0
cc_630 N_A_593_125#_M1037_d N_VPWR_c_1419_n 0.00540229f $X=3.035 $Y=2.675 $X2=0
+ $Y2=0
cc_631 N_A_593_125#_M1019_g N_VPWR_c_1419_n 0.00563653f $X=4.725 $Y=2.885 $X2=0
+ $Y2=0
cc_632 N_A_593_125#_M1010_g N_VPWR_c_1419_n 0.00638175f $X=6.365 $Y=2.675 $X2=0
+ $Y2=0
cc_633 N_A_593_125#_c_718_n N_VPWR_c_1419_n 0.00978375f $X=3.21 $Y=2.88 $X2=0
+ $Y2=0
cc_634 N_A_593_125#_c_719_n N_VPWR_c_1419_n 0.0156424f $X=3.825 $Y=2.45 $X2=0
+ $Y2=0
cc_635 N_A_593_125#_c_708_n N_A_507_125#_c_1573_n 0.0133322f $X=3.205 $Y=2.365
+ $X2=0 $Y2=0
cc_636 N_A_593_125#_c_708_n N_A_507_125#_c_1574_n 0.0675233f $X=3.205 $Y=2.365
+ $X2=0 $Y2=0
cc_637 N_A_593_125#_c_718_n N_A_507_125#_c_1574_n 0.0118228f $X=3.21 $Y=2.88
+ $X2=0 $Y2=0
cc_638 N_A_593_125#_c_725_n N_A_507_125#_c_1574_n 0.0137656f $X=3.245 $Y=2.45
+ $X2=0 $Y2=0
cc_639 N_A_593_125#_c_708_n N_A_507_125#_c_1575_n 0.0127318f $X=3.205 $Y=2.365
+ $X2=0 $Y2=0
cc_640 N_A_593_125#_c_718_n N_A_507_125#_c_1592_n 0.0249791f $X=3.21 $Y=2.88
+ $X2=0 $Y2=0
cc_641 N_A_593_125#_c_703_n N_VGND_c_1652_n 0.00956091f $X=5.79 $Y=1.375 $X2=0
+ $Y2=0
cc_642 N_A_593_125#_c_703_n N_VGND_c_1674_n 7.97988e-19 $X=5.79 $Y=1.375 $X2=0
+ $Y2=0
cc_643 N_A_593_125#_c_703_n N_A_1173_125#_c_1795_n 0.00311519f $X=5.79 $Y=1.375
+ $X2=0 $Y2=0
cc_644 N_A_593_125#_c_704_n N_A_1173_125#_c_1795_n 9.39241e-19 $X=6.08 $Y=1.45
+ $X2=0 $Y2=0
cc_645 N_A_593_125#_c_703_n N_A_1280_159#_c_1822_n 0.0043559f $X=5.79 $Y=1.375
+ $X2=0 $Y2=0
cc_646 N_SET_B_M1022_g N_A_191_21#_c_997_n 0.00462072f $X=5.265 $Y=1.055 $X2=0
+ $Y2=0
cc_647 N_SET_B_c_886_n N_A_191_21#_M1026_g 0.00574715f $X=7.43 $Y=2.99 $X2=0
+ $Y2=0
cc_648 N_SET_B_c_887_n N_A_191_21#_M1026_g 0.00633999f $X=7.525 $Y=2.905 $X2=0
+ $Y2=0
cc_649 N_SET_B_c_888_n N_A_191_21#_M1026_g 0.0027235f $X=7.62 $Y=1.93 $X2=0
+ $Y2=0
cc_650 N_SET_B_c_887_n N_A_1533_258#_M1013_g 0.00707104f $X=7.525 $Y=2.905 $X2=0
+ $Y2=0
cc_651 N_SET_B_c_889_n N_A_1533_258#_M1013_g 0.0203719f $X=8.26 $Y=1.93 $X2=0
+ $Y2=0
cc_652 N_SET_B_c_891_n N_A_1533_258#_M1013_g 0.0291276f $X=8.26 $Y=1.84 $X2=0
+ $Y2=0
cc_653 N_SET_B_c_889_n N_A_1533_258#_c_1126_n 0.00146309f $X=8.26 $Y=1.93 $X2=0
+ $Y2=0
cc_654 N_SET_B_c_880_n N_A_1533_258#_c_1128_n 4.21308e-19 $X=8.595 $Y=1.84 $X2=0
+ $Y2=0
cc_655 N_SET_B_M1014_g N_A_1533_258#_c_1128_n 0.0193453f $X=8.67 $Y=0.665 $X2=0
+ $Y2=0
cc_656 N_SET_B_c_889_n N_A_1533_258#_c_1129_n 2.5116e-19 $X=8.26 $Y=1.93 $X2=0
+ $Y2=0
cc_657 N_SET_B_c_891_n N_A_1533_258#_c_1129_n 0.0105541f $X=8.26 $Y=1.84 $X2=0
+ $Y2=0
cc_658 N_SET_B_c_880_n N_A_1533_258#_c_1137_n 0.00214962f $X=8.595 $Y=1.84 $X2=0
+ $Y2=0
cc_659 N_SET_B_M1014_g N_A_1533_258#_c_1132_n 0.0045537f $X=8.67 $Y=0.665 $X2=0
+ $Y2=0
cc_660 N_SET_B_M1014_g N_A_1533_258#_c_1133_n 0.0707301f $X=8.67 $Y=0.665 $X2=0
+ $Y2=0
cc_661 N_SET_B_c_886_n N_A_1360_451#_M1009_d 0.00522477f $X=7.43 $Y=2.99 $X2=0
+ $Y2=0
cc_662 N_SET_B_M1014_g N_A_1360_451#_c_1210_n 0.0060441f $X=8.67 $Y=0.665 $X2=0
+ $Y2=0
cc_663 N_SET_B_c_887_n N_A_1360_451#_c_1225_n 0.0211874f $X=7.525 $Y=2.905 $X2=0
+ $Y2=0
cc_664 N_SET_B_c_888_n N_A_1360_451#_c_1225_n 0.0255037f $X=7.62 $Y=1.93 $X2=0
+ $Y2=0
cc_665 N_SET_B_c_890_n N_A_1360_451#_c_1225_n 0.0045826f $X=6.435 $Y=2.347 $X2=0
+ $Y2=0
cc_666 N_SET_B_c_888_n N_A_1360_451#_c_1226_n 0.0154702f $X=7.62 $Y=1.93 $X2=0
+ $Y2=0
cc_667 N_SET_B_c_889_n N_A_1360_451#_c_1226_n 0.0531623f $X=8.26 $Y=1.93 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_891_n N_A_1360_451#_c_1226_n 0.00756919f $X=8.26 $Y=1.84 $X2=0
+ $Y2=0
cc_669 N_SET_B_M1005_g N_A_1360_451#_c_1227_n 0.0051627f $X=8.17 $Y=2.465 $X2=0
+ $Y2=0
cc_670 N_SET_B_c_880_n N_A_1360_451#_c_1227_n 0.012719f $X=8.595 $Y=1.84 $X2=0
+ $Y2=0
cc_671 N_SET_B_M1014_g N_A_1360_451#_c_1227_n 0.00693867f $X=8.67 $Y=0.665 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_889_n N_A_1360_451#_c_1227_n 0.0245334f $X=8.26 $Y=1.93 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_891_n N_A_1360_451#_c_1227_n 0.00442186f $X=8.26 $Y=1.84 $X2=0
+ $Y2=0
cc_674 N_SET_B_M1014_g N_A_1360_451#_c_1228_n 0.00832756f $X=8.67 $Y=0.665 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_886_n N_A_1360_451#_c_1238_n 0.0293966f $X=7.43 $Y=2.99 $X2=0
+ $Y2=0
cc_676 N_SET_B_c_887_n N_A_1360_451#_c_1238_n 0.0241886f $X=7.525 $Y=2.905 $X2=0
+ $Y2=0
cc_677 N_SET_B_c_880_n N_A_1360_451#_c_1239_n 0.00354461f $X=8.595 $Y=1.84 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_889_n N_A_1360_451#_c_1239_n 0.00487842f $X=8.26 $Y=1.93 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_891_n N_A_1360_451#_c_1239_n 0.00511371f $X=8.26 $Y=1.84 $X2=0
+ $Y2=0
cc_680 N_SET_B_M1014_g N_A_1360_451#_c_1230_n 0.00844761f $X=8.67 $Y=0.665 $X2=0
+ $Y2=0
cc_681 N_SET_B_c_890_n N_VPWR_M1017_d 0.00241037f $X=6.435 $Y=2.347 $X2=0 $Y2=0
cc_682 N_SET_B_M1017_g N_VPWR_c_1423_n 0.00837592f $X=5.84 $Y=2.885 $X2=0 $Y2=0
cc_683 N_SET_B_c_890_n N_VPWR_c_1423_n 0.0204684f $X=6.435 $Y=2.347 $X2=0 $Y2=0
cc_684 N_SET_B_M1005_g N_VPWR_c_1424_n 0.00381165f $X=8.17 $Y=2.465 $X2=0 $Y2=0
cc_685 N_SET_B_c_886_n N_VPWR_c_1424_n 0.0149189f $X=7.43 $Y=2.99 $X2=0 $Y2=0
cc_686 N_SET_B_c_887_n N_VPWR_c_1424_n 0.0323689f $X=7.525 $Y=2.905 $X2=0 $Y2=0
cc_687 N_SET_B_c_889_n N_VPWR_c_1424_n 0.0197276f $X=8.26 $Y=1.93 $X2=0 $Y2=0
cc_688 N_SET_B_M1017_g N_VPWR_c_1431_n 0.00585385f $X=5.84 $Y=2.885 $X2=0 $Y2=0
cc_689 N_SET_B_c_886_n N_VPWR_c_1432_n 0.0631017f $X=7.43 $Y=2.99 $X2=0 $Y2=0
cc_690 N_SET_B_c_929_n N_VPWR_c_1432_n 0.00953907f $X=6.605 $Y=2.99 $X2=0 $Y2=0
cc_691 N_SET_B_M1005_g N_VPWR_c_1433_n 0.00399858f $X=8.17 $Y=2.465 $X2=0 $Y2=0
cc_692 N_SET_B_M1017_g N_VPWR_c_1419_n 0.00810941f $X=5.84 $Y=2.885 $X2=0 $Y2=0
cc_693 N_SET_B_M1005_g N_VPWR_c_1419_n 0.0046122f $X=8.17 $Y=2.465 $X2=0 $Y2=0
cc_694 N_SET_B_c_886_n N_VPWR_c_1419_n 0.0377143f $X=7.43 $Y=2.99 $X2=0 $Y2=0
cc_695 N_SET_B_c_929_n N_VPWR_c_1419_n 0.00658633f $X=6.605 $Y=2.99 $X2=0 $Y2=0
cc_696 N_SET_B_c_890_n N_VPWR_c_1419_n 0.0146323f $X=6.435 $Y=2.347 $X2=0 $Y2=0
cc_697 N_SET_B_c_929_n A_1288_451# 9.38685e-19 $X=6.605 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_698 N_SET_B_c_887_n A_1468_451# 0.00749677f $X=7.525 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_699 N_SET_B_M1022_g N_VGND_c_1652_n 0.00278037f $X=5.265 $Y=1.055 $X2=0 $Y2=0
cc_700 N_SET_B_M1014_g N_VGND_c_1653_n 0.0118443f $X=8.67 $Y=0.665 $X2=0 $Y2=0
cc_701 N_SET_B_M1014_g N_VGND_c_1665_n 0.00429764f $X=8.67 $Y=0.665 $X2=0 $Y2=0
cc_702 N_SET_B_M1022_g N_VGND_c_1674_n 9.7053e-19 $X=5.265 $Y=1.055 $X2=0 $Y2=0
cc_703 N_SET_B_M1014_g N_VGND_c_1674_n 0.00435987f $X=8.67 $Y=0.665 $X2=0 $Y2=0
cc_704 N_SET_B_M1014_g N_A_1280_159#_c_1824_n 8.23231e-19 $X=8.67 $Y=0.665 $X2=0
+ $Y2=0
cc_705 N_A_191_21#_M1026_g N_A_1533_258#_c_1127_n 0.0494849f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_706 N_A_191_21#_M1026_g N_A_1533_258#_c_1128_n 0.00115549f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_707 N_A_191_21#_M1026_g N_A_1533_258#_c_1129_n 0.00423865f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_708 N_A_191_21#_M1026_g N_A_1360_451#_c_1224_n 0.00886484f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_709 N_A_191_21#_M1026_g N_A_1360_451#_c_1225_n 0.0175386f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_710 N_A_191_21#_M1026_g N_A_1360_451#_c_1226_n 0.0102332f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_711 N_A_191_21#_M1026_g N_A_1360_451#_c_1238_n 0.00976692f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_712 N_A_191_21#_M1026_g N_A_1360_451#_c_1249_n 0.0103784f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_713 N_A_191_21#_M1026_g N_A_1360_451#_c_1229_n 0.00184921f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_714 N_A_191_21#_c_1008_n N_VPWR_c_1422_n 0.00821782f $X=1.612 $Y=2.475 $X2=0
+ $Y2=0
cc_715 N_A_191_21#_c_1008_n N_VPWR_c_1430_n 0.0112439f $X=1.612 $Y=2.475 $X2=0
+ $Y2=0
cc_716 N_A_191_21#_M1037_g N_VPWR_c_1438_n 0.0049848f $X=2.96 $Y=2.885 $X2=0
+ $Y2=0
cc_717 N_A_191_21#_M1037_g N_VPWR_c_1419_n 0.00891106f $X=2.96 $Y=2.885 $X2=0
+ $Y2=0
cc_718 N_A_191_21#_c_1008_n N_VPWR_c_1419_n 0.0166153f $X=1.612 $Y=2.475 $X2=0
+ $Y2=0
cc_719 N_A_191_21#_c_1003_n N_A_507_125#_c_1574_n 0.0108985f $X=2.885 $Y=1.9
+ $X2=0 $Y2=0
cc_720 N_A_191_21#_M1037_g N_A_507_125#_c_1574_n 0.0155774f $X=2.96 $Y=2.885
+ $X2=0 $Y2=0
cc_721 N_A_191_21#_c_1003_n N_A_507_125#_c_1575_n 0.00489743f $X=2.885 $Y=1.9
+ $X2=0 $Y2=0
cc_722 N_A_191_21#_M1037_g N_A_507_125#_c_1592_n 0.00493751f $X=2.96 $Y=2.885
+ $X2=0 $Y2=0
cc_723 N_A_191_21#_c_994_n N_VGND_c_1649_n 0.00141128f $X=1.06 $Y=1.725 $X2=0
+ $Y2=0
cc_724 N_A_191_21#_c_1000_n N_VGND_c_1649_n 0.0226174f $X=1.12 $Y=0.35 $X2=0
+ $Y2=0
cc_725 N_A_191_21#_c_1001_n N_VGND_c_1649_n 0.00730385f $X=1.12 $Y=0.18 $X2=0
+ $Y2=0
cc_726 N_A_191_21#_c_995_n N_VGND_c_1650_n 0.0258691f $X=3.245 $Y=0.18 $X2=0
+ $Y2=0
cc_727 N_A_191_21#_c_1000_n N_VGND_c_1650_n 0.0389712f $X=1.12 $Y=0.35 $X2=0
+ $Y2=0
cc_728 N_A_191_21#_c_1001_n N_VGND_c_1650_n 9.97882e-19 $X=1.12 $Y=0.18 $X2=0
+ $Y2=0
cc_729 N_A_191_21#_M1021_g N_VGND_c_1651_n 8.25021e-19 $X=3.32 $Y=0.835 $X2=0
+ $Y2=0
cc_730 N_A_191_21#_c_997_n N_VGND_c_1651_n 0.0221195f $X=7.19 $Y=0.18 $X2=0
+ $Y2=0
cc_731 N_A_191_21#_c_997_n N_VGND_c_1652_n 0.0258253f $X=7.19 $Y=0.18 $X2=0
+ $Y2=0
cc_732 N_A_191_21#_c_1000_n N_VGND_c_1660_n 0.0399799f $X=1.12 $Y=0.35 $X2=0
+ $Y2=0
cc_733 N_A_191_21#_c_1001_n N_VGND_c_1660_n 0.0196246f $X=1.12 $Y=0.18 $X2=0
+ $Y2=0
cc_734 N_A_191_21#_c_995_n N_VGND_c_1662_n 0.0417864f $X=3.245 $Y=0.18 $X2=0
+ $Y2=0
cc_735 N_A_191_21#_c_997_n N_VGND_c_1664_n 0.0364619f $X=7.19 $Y=0.18 $X2=0
+ $Y2=0
cc_736 N_A_191_21#_c_997_n N_VGND_c_1665_n 0.0358398f $X=7.19 $Y=0.18 $X2=0
+ $Y2=0
cc_737 N_A_191_21#_c_995_n N_VGND_c_1674_n 0.046268f $X=3.245 $Y=0.18 $X2=0
+ $Y2=0
cc_738 N_A_191_21#_c_997_n N_VGND_c_1674_n 0.097996f $X=7.19 $Y=0.18 $X2=0 $Y2=0
cc_739 N_A_191_21#_c_999_n N_VGND_c_1674_n 0.00370846f $X=3.32 $Y=0.18 $X2=0
+ $Y2=0
cc_740 N_A_191_21#_c_1000_n N_VGND_c_1674_n 0.0202224f $X=1.12 $Y=0.35 $X2=0
+ $Y2=0
cc_741 N_A_191_21#_c_1001_n N_VGND_c_1674_n 0.0102769f $X=1.12 $Y=0.18 $X2=0
+ $Y2=0
cc_742 N_A_191_21#_c_997_n N_A_1173_125#_c_1796_n 0.00640469f $X=7.19 $Y=0.18
+ $X2=0 $Y2=0
cc_743 N_A_191_21#_c_997_n N_A_1173_125#_c_1797_n 0.0197706f $X=7.19 $Y=0.18
+ $X2=0 $Y2=0
cc_744 N_A_191_21#_M1026_g N_A_1173_125#_c_1797_n 0.0152496f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_745 N_A_191_21#_M1026_g N_A_1280_159#_c_1824_n 0.00321849f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_746 N_A_191_21#_M1026_g N_A_1280_159#_c_1825_n 0.0144458f $X=7.265 $Y=0.895
+ $X2=0 $Y2=0
cc_747 N_A_1533_258#_c_1131_n N_A_1360_451#_c_1210_n 0.00420153f $X=9.92
+ $Y=1.815 $X2=0 $Y2=0
cc_748 N_A_1533_258#_c_1137_n N_A_1360_451#_c_1210_n 0.00422235f $X=9.365 $Y=1.9
+ $X2=0 $Y2=0
cc_749 N_A_1533_258#_c_1132_n N_A_1360_451#_c_1210_n 0.00569925f $X=9.405
+ $Y=0.865 $X2=0 $Y2=0
cc_750 N_A_1533_258#_c_1135_n N_A_1360_451#_M1024_g 0.0115399f $X=9.835 $Y=1.9
+ $X2=0 $Y2=0
cc_751 N_A_1533_258#_c_1137_n N_A_1360_451#_M1024_g 0.00733576f $X=9.365 $Y=1.9
+ $X2=0 $Y2=0
cc_752 N_A_1533_258#_c_1128_n N_A_1360_451#_M1007_g 6.00194e-19 $X=9.24 $Y=1.11
+ $X2=0 $Y2=0
cc_753 N_A_1533_258#_c_1130_n N_A_1360_451#_M1007_g 0.0120911f $X=9.835 $Y=1.15
+ $X2=0 $Y2=0
cc_754 N_A_1533_258#_c_1131_n N_A_1360_451#_M1007_g 0.00222611f $X=9.92 $Y=1.815
+ $X2=0 $Y2=0
cc_755 N_A_1533_258#_c_1132_n N_A_1360_451#_M1007_g 0.0111805f $X=9.405 $Y=0.865
+ $X2=0 $Y2=0
cc_756 N_A_1533_258#_c_1135_n N_A_1360_451#_c_1212_n 0.00195296f $X=9.835 $Y=1.9
+ $X2=0 $Y2=0
cc_757 N_A_1533_258#_c_1130_n N_A_1360_451#_c_1212_n 0.00126753f $X=9.835
+ $Y=1.15 $X2=0 $Y2=0
cc_758 N_A_1533_258#_c_1131_n N_A_1360_451#_c_1212_n 0.0139777f $X=9.92 $Y=1.815
+ $X2=0 $Y2=0
cc_759 N_A_1533_258#_c_1135_n N_A_1360_451#_M1004_g 0.0010712f $X=9.835 $Y=1.9
+ $X2=0 $Y2=0
cc_760 N_A_1533_258#_c_1131_n N_A_1360_451#_M1004_g 0.00312471f $X=9.92 $Y=1.815
+ $X2=0 $Y2=0
cc_761 N_A_1533_258#_c_1137_n N_A_1360_451#_M1004_g 5.35638e-19 $X=9.365 $Y=1.9
+ $X2=0 $Y2=0
cc_762 N_A_1533_258#_c_1130_n N_A_1360_451#_M1015_g 0.00162955f $X=9.835 $Y=1.15
+ $X2=0 $Y2=0
cc_763 N_A_1533_258#_c_1131_n N_A_1360_451#_M1015_g 8.65672e-19 $X=9.92 $Y=1.815
+ $X2=0 $Y2=0
cc_764 N_A_1533_258#_c_1132_n N_A_1360_451#_M1015_g 5.10709e-19 $X=9.405
+ $Y=0.865 $X2=0 $Y2=0
cc_765 N_A_1533_258#_c_1127_n N_A_1360_451#_c_1224_n 7.08497e-19 $X=7.815
+ $Y=1.365 $X2=0 $Y2=0
cc_766 N_A_1533_258#_M1013_g N_A_1360_451#_c_1225_n 0.00128172f $X=7.74 $Y=2.465
+ $X2=0 $Y2=0
cc_767 N_A_1533_258#_M1013_g N_A_1360_451#_c_1226_n 0.00946709f $X=7.74 $Y=2.465
+ $X2=0 $Y2=0
cc_768 N_A_1533_258#_c_1126_n N_A_1360_451#_c_1226_n 0.00810888f $X=8.025
+ $Y=1.365 $X2=0 $Y2=0
cc_769 N_A_1533_258#_c_1127_n N_A_1360_451#_c_1226_n 0.00372155f $X=7.815
+ $Y=1.365 $X2=0 $Y2=0
cc_770 N_A_1533_258#_c_1128_n N_A_1360_451#_c_1226_n 0.0361217f $X=9.24 $Y=1.11
+ $X2=0 $Y2=0
cc_771 N_A_1533_258#_c_1129_n N_A_1360_451#_c_1226_n 0.0100114f $X=8.19 $Y=1.15
+ $X2=0 $Y2=0
cc_772 N_A_1533_258#_c_1137_n N_A_1360_451#_c_1227_n 0.0143623f $X=9.365 $Y=1.9
+ $X2=0 $Y2=0
cc_773 N_A_1533_258#_c_1128_n N_A_1360_451#_c_1228_n 0.0429489f $X=9.24 $Y=1.11
+ $X2=0 $Y2=0
cc_774 N_A_1533_258#_c_1135_n N_A_1360_451#_c_1228_n 0.00870314f $X=9.835 $Y=1.9
+ $X2=0 $Y2=0
cc_775 N_A_1533_258#_c_1130_n N_A_1360_451#_c_1228_n 0.00591813f $X=9.835
+ $Y=1.15 $X2=0 $Y2=0
cc_776 N_A_1533_258#_c_1131_n N_A_1360_451#_c_1228_n 0.0179126f $X=9.92 $Y=1.815
+ $X2=0 $Y2=0
cc_777 N_A_1533_258#_c_1137_n N_A_1360_451#_c_1228_n 0.0262619f $X=9.365 $Y=1.9
+ $X2=0 $Y2=0
cc_778 N_A_1533_258#_c_1132_n N_A_1360_451#_c_1228_n 0.0267562f $X=9.405
+ $Y=0.865 $X2=0 $Y2=0
cc_779 N_A_1533_258#_c_1128_n N_A_1360_451#_c_1230_n 0.0138972f $X=9.24 $Y=1.11
+ $X2=0 $Y2=0
cc_780 N_A_1533_258#_c_1135_n N_VPWR_M1024_d 0.0042876f $X=9.835 $Y=1.9 $X2=0
+ $Y2=0
cc_781 N_A_1533_258#_M1013_g N_VPWR_c_1424_n 0.0079873f $X=7.74 $Y=2.465 $X2=0
+ $Y2=0
cc_782 N_A_1533_258#_c_1135_n N_VPWR_c_1425_n 0.0212739f $X=9.835 $Y=1.9 $X2=0
+ $Y2=0
cc_783 N_A_1533_258#_c_1137_n N_VPWR_c_1425_n 0.00384115f $X=9.365 $Y=1.9 $X2=0
+ $Y2=0
cc_784 N_A_1533_258#_M1013_g N_VPWR_c_1432_n 0.00332367f $X=7.74 $Y=2.465 $X2=0
+ $Y2=0
cc_785 N_A_1533_258#_M1013_g N_VPWR_c_1419_n 0.00387424f $X=7.74 $Y=2.465 $X2=0
+ $Y2=0
cc_786 N_A_1533_258#_c_1135_n N_Q_N_c_1611_n 0.00133226f $X=9.835 $Y=1.9 $X2=0
+ $Y2=0
cc_787 N_A_1533_258#_c_1130_n N_Q_N_c_1611_n 0.0114431f $X=9.835 $Y=1.15 $X2=0
+ $Y2=0
cc_788 N_A_1533_258#_c_1131_n N_Q_N_c_1611_n 0.0361618f $X=9.92 $Y=1.815 $X2=0
+ $Y2=0
cc_789 N_A_1533_258#_c_1130_n N_VGND_M1007_d 0.00329355f $X=9.835 $Y=1.15 $X2=0
+ $Y2=0
cc_790 N_A_1533_258#_c_1128_n N_VGND_c_1653_n 0.0251776f $X=9.24 $Y=1.11 $X2=0
+ $Y2=0
cc_791 N_A_1533_258#_c_1132_n N_VGND_c_1653_n 0.00885527f $X=9.405 $Y=0.865
+ $X2=0 $Y2=0
cc_792 N_A_1533_258#_c_1133_n N_VGND_c_1653_n 0.00176217f $X=8.205 $Y=0.985
+ $X2=0 $Y2=0
cc_793 N_A_1533_258#_c_1132_n N_VGND_c_1654_n 0.00495237f $X=9.405 $Y=0.865
+ $X2=0 $Y2=0
cc_794 N_A_1533_258#_c_1130_n N_VGND_c_1655_n 0.0209047f $X=9.835 $Y=1.15 $X2=0
+ $Y2=0
cc_795 N_A_1533_258#_c_1132_n N_VGND_c_1655_n 0.0134837f $X=9.405 $Y=0.865 $X2=0
+ $Y2=0
cc_796 N_A_1533_258#_c_1133_n N_VGND_c_1665_n 0.00494981f $X=8.205 $Y=0.985
+ $X2=0 $Y2=0
cc_797 N_A_1533_258#_c_1132_n N_VGND_c_1674_n 0.00933518f $X=9.405 $Y=0.865
+ $X2=0 $Y2=0
cc_798 N_A_1533_258#_c_1133_n N_VGND_c_1674_n 0.00519032f $X=8.205 $Y=0.985
+ $X2=0 $Y2=0
cc_799 N_A_1533_258#_c_1133_n N_A_1173_125#_c_1797_n 0.00406297f $X=8.205
+ $Y=0.985 $X2=0 $Y2=0
cc_800 N_A_1533_258#_c_1126_n N_A_1280_159#_c_1824_n 0.0032694f $X=8.025
+ $Y=1.365 $X2=0 $Y2=0
cc_801 N_A_1533_258#_c_1128_n N_A_1280_159#_c_1824_n 0.0147335f $X=9.24 $Y=1.11
+ $X2=0 $Y2=0
cc_802 N_A_1533_258#_c_1129_n N_A_1280_159#_c_1824_n 0.00491826f $X=8.19 $Y=1.15
+ $X2=0 $Y2=0
cc_803 N_A_1533_258#_c_1133_n N_A_1280_159#_c_1824_n 0.00554515f $X=8.205
+ $Y=0.985 $X2=0 $Y2=0
cc_804 N_A_1533_258#_c_1127_n N_A_1280_159#_c_1825_n 0.0032694f $X=7.815
+ $Y=1.365 $X2=0 $Y2=0
cc_805 N_A_1360_451#_M1030_g N_A_2227_367#_c_1370_n 0.00138693f $X=10.575
+ $Y=0.655 $X2=0 $Y2=0
cc_806 N_A_1360_451#_M1018_g N_A_2227_367#_c_1370_n 0.0147566f $X=11.1 $Y=0.865
+ $X2=0 $Y2=0
cc_807 N_A_1360_451#_c_1223_n N_A_2227_367#_c_1370_n 6.11479e-19 $X=11.08
+ $Y=1.41 $X2=0 $Y2=0
cc_808 N_A_1360_451#_M1034_g N_A_2227_367#_c_1377_n 0.00679221f $X=11.06
+ $Y=2.155 $X2=0 $Y2=0
cc_809 N_A_1360_451#_M1034_g N_A_2227_367#_c_1372_n 0.00704323f $X=11.06
+ $Y=2.155 $X2=0 $Y2=0
cc_810 N_A_1360_451#_c_1223_n N_A_2227_367#_c_1372_n 0.0108835f $X=11.08 $Y=1.41
+ $X2=0 $Y2=0
cc_811 N_A_1360_451#_M1034_g N_A_2227_367#_c_1373_n 0.00237661f $X=11.06
+ $Y=2.155 $X2=0 $Y2=0
cc_812 N_A_1360_451#_c_1223_n N_A_2227_367#_c_1373_n 0.00230239f $X=11.08
+ $Y=1.41 $X2=0 $Y2=0
cc_813 N_A_1360_451#_M1024_g N_VPWR_c_1425_n 0.00534536f $X=9.58 $Y=2.045 $X2=0
+ $Y2=0
cc_814 N_A_1360_451#_c_1212_n N_VPWR_c_1425_n 4.36491e-19 $X=10.03 $Y=1.41 $X2=0
+ $Y2=0
cc_815 N_A_1360_451#_M1004_g N_VPWR_c_1425_n 0.0156731f $X=10.105 $Y=2.465 $X2=0
+ $Y2=0
cc_816 N_A_1360_451#_M1035_g N_VPWR_c_1425_n 7.86599e-19 $X=10.535 $Y=2.465
+ $X2=0 $Y2=0
cc_817 N_A_1360_451#_M1035_g N_VPWR_c_1426_n 0.00783454f $X=10.535 $Y=2.465
+ $X2=0 $Y2=0
cc_818 N_A_1360_451#_c_1218_n N_VPWR_c_1426_n 0.00700485f $X=10.985 $Y=1.41
+ $X2=0 $Y2=0
cc_819 N_A_1360_451#_M1034_g N_VPWR_c_1426_n 0.00571559f $X=11.06 $Y=2.155 $X2=0
+ $Y2=0
cc_820 N_A_1360_451#_M1034_g N_VPWR_c_1427_n 0.00399067f $X=11.06 $Y=2.155 $X2=0
+ $Y2=0
cc_821 N_A_1360_451#_c_1239_n N_VPWR_c_1433_n 0.00647361f $X=8.61 $Y=2.44 $X2=0
+ $Y2=0
cc_822 N_A_1360_451#_M1004_g N_VPWR_c_1434_n 0.00486043f $X=10.105 $Y=2.465
+ $X2=0 $Y2=0
cc_823 N_A_1360_451#_M1035_g N_VPWR_c_1434_n 0.00579312f $X=10.535 $Y=2.465
+ $X2=0 $Y2=0
cc_824 N_A_1360_451#_M1034_g N_VPWR_c_1435_n 0.00312414f $X=11.06 $Y=2.155 $X2=0
+ $Y2=0
cc_825 N_A_1360_451#_M1009_d N_VPWR_c_1419_n 0.00224358f $X=6.8 $Y=2.255 $X2=0
+ $Y2=0
cc_826 N_A_1360_451#_M1004_g N_VPWR_c_1419_n 0.00824727f $X=10.105 $Y=2.465
+ $X2=0 $Y2=0
cc_827 N_A_1360_451#_M1035_g N_VPWR_c_1419_n 0.011752f $X=10.535 $Y=2.465 $X2=0
+ $Y2=0
cc_828 N_A_1360_451#_M1034_g N_VPWR_c_1419_n 0.00410284f $X=11.06 $Y=2.155 $X2=0
+ $Y2=0
cc_829 N_A_1360_451#_c_1239_n N_VPWR_c_1419_n 0.0120614f $X=8.61 $Y=2.44 $X2=0
+ $Y2=0
cc_830 N_A_1360_451#_M1004_g N_Q_N_c_1611_n 0.00334796f $X=10.105 $Y=2.465 $X2=0
+ $Y2=0
cc_831 N_A_1360_451#_M1015_g N_Q_N_c_1611_n 0.002957f $X=10.145 $Y=0.655 $X2=0
+ $Y2=0
cc_832 N_A_1360_451#_c_1215_n N_Q_N_c_1611_n 0.010581f $X=10.46 $Y=1.41 $X2=0
+ $Y2=0
cc_833 N_A_1360_451#_M1035_g N_Q_N_c_1611_n 0.0217774f $X=10.535 $Y=2.465 $X2=0
+ $Y2=0
cc_834 N_A_1360_451#_M1030_g N_Q_N_c_1611_n 0.00703187f $X=10.575 $Y=0.655 $X2=0
+ $Y2=0
cc_835 N_A_1360_451#_M1034_g N_Q_N_c_1611_n 0.00166796f $X=11.06 $Y=2.155 $X2=0
+ $Y2=0
cc_836 N_A_1360_451#_c_1222_n N_Q_N_c_1611_n 0.00696109f $X=10.555 $Y=1.41 $X2=0
+ $Y2=0
cc_837 N_A_1360_451#_M1007_g N_VGND_c_1653_n 0.00425581f $X=9.62 $Y=0.865 $X2=0
+ $Y2=0
cc_838 N_A_1360_451#_M1007_g N_VGND_c_1654_n 0.00385987f $X=9.62 $Y=0.865 $X2=0
+ $Y2=0
cc_839 N_A_1360_451#_M1007_g N_VGND_c_1655_n 0.0064429f $X=9.62 $Y=0.865 $X2=0
+ $Y2=0
cc_840 N_A_1360_451#_c_1212_n N_VGND_c_1655_n 7.3941e-19 $X=10.03 $Y=1.41 $X2=0
+ $Y2=0
cc_841 N_A_1360_451#_M1015_g N_VGND_c_1655_n 0.00337289f $X=10.145 $Y=0.655
+ $X2=0 $Y2=0
cc_842 N_A_1360_451#_M1015_g N_VGND_c_1656_n 6.90821e-19 $X=10.145 $Y=0.655
+ $X2=0 $Y2=0
cc_843 N_A_1360_451#_M1030_g N_VGND_c_1656_n 0.020303f $X=10.575 $Y=0.655 $X2=0
+ $Y2=0
cc_844 N_A_1360_451#_c_1218_n N_VGND_c_1656_n 0.00770539f $X=10.985 $Y=1.41
+ $X2=0 $Y2=0
cc_845 N_A_1360_451#_M1018_g N_VGND_c_1656_n 0.00435171f $X=11.1 $Y=0.865 $X2=0
+ $Y2=0
cc_846 N_A_1360_451#_M1018_g N_VGND_c_1657_n 0.00520592f $X=11.1 $Y=0.865 $X2=0
+ $Y2=0
cc_847 N_A_1360_451#_M1015_g N_VGND_c_1666_n 0.00585385f $X=10.145 $Y=0.655
+ $X2=0 $Y2=0
cc_848 N_A_1360_451#_M1030_g N_VGND_c_1666_n 0.00525069f $X=10.575 $Y=0.655
+ $X2=0 $Y2=0
cc_849 N_A_1360_451#_M1018_g N_VGND_c_1667_n 0.00385987f $X=11.1 $Y=0.865 $X2=0
+ $Y2=0
cc_850 N_A_1360_451#_M1007_g N_VGND_c_1674_n 0.0046122f $X=9.62 $Y=0.865 $X2=0
+ $Y2=0
cc_851 N_A_1360_451#_M1015_g N_VGND_c_1674_n 0.0118358f $X=10.145 $Y=0.655 $X2=0
+ $Y2=0
cc_852 N_A_1360_451#_M1030_g N_VGND_c_1674_n 0.00886509f $X=10.575 $Y=0.655
+ $X2=0 $Y2=0
cc_853 N_A_1360_451#_M1018_g N_VGND_c_1674_n 0.0046122f $X=11.1 $Y=0.865 $X2=0
+ $Y2=0
cc_854 N_A_1360_451#_M1020_d N_A_1280_159#_c_1825_n 0.00467306f $X=6.815
+ $Y=0.795 $X2=0 $Y2=0
cc_855 N_A_1360_451#_c_1226_n N_A_1280_159#_c_1825_n 0.0209952f $X=8.525
+ $Y=1.495 $X2=0 $Y2=0
cc_856 N_A_1360_451#_c_1249_n N_A_1280_159#_c_1825_n 0.0232747f $X=7.165
+ $Y=1.075 $X2=0 $Y2=0
cc_857 N_A_2227_367#_c_1377_n N_VPWR_c_1426_n 0.00232431f $X=11.275 $Y=1.98
+ $X2=0 $Y2=0
cc_858 N_A_2227_367#_M1001_g N_VPWR_c_1427_n 0.00671101f $X=12.05 $Y=2.465 $X2=0
+ $Y2=0
cc_859 N_A_2227_367#_c_1377_n N_VPWR_c_1427_n 0.0462938f $X=11.275 $Y=1.98 $X2=0
+ $Y2=0
cc_860 N_A_2227_367#_c_1371_n N_VPWR_c_1427_n 0.0227997f $X=11.89 $Y=1.51 $X2=0
+ $Y2=0
cc_861 N_A_2227_367#_c_1373_n N_VPWR_c_1427_n 0.00562998f $X=11.925 $Y=1.42
+ $X2=0 $Y2=0
cc_862 N_A_2227_367#_M1016_g N_VPWR_c_1429_n 0.00777219f $X=12.48 $Y=2.465 $X2=0
+ $Y2=0
cc_863 N_A_2227_367#_M1001_g N_VPWR_c_1436_n 0.00583607f $X=12.05 $Y=2.465 $X2=0
+ $Y2=0
cc_864 N_A_2227_367#_M1016_g N_VPWR_c_1436_n 0.00585385f $X=12.48 $Y=2.465 $X2=0
+ $Y2=0
cc_865 N_A_2227_367#_M1001_g N_VPWR_c_1419_n 0.0117786f $X=12.05 $Y=2.465 $X2=0
+ $Y2=0
cc_866 N_A_2227_367#_M1016_g N_VPWR_c_1419_n 0.011446f $X=12.48 $Y=2.465 $X2=0
+ $Y2=0
cc_867 N_A_2227_367#_c_1377_n N_VPWR_c_1419_n 0.0122878f $X=11.275 $Y=1.98 $X2=0
+ $Y2=0
cc_868 N_A_2227_367#_c_1366_n N_Q_c_1631_n 0.0163556f $X=12.405 $Y=1.42 $X2=0
+ $Y2=0
cc_869 N_A_2227_367#_c_1367_n N_Q_c_1631_n 0.00345904f $X=12.48 $Y=1.345 $X2=0
+ $Y2=0
cc_870 N_A_2227_367#_M1016_g N_Q_c_1631_n 0.00954344f $X=12.48 $Y=2.465 $X2=0
+ $Y2=0
cc_871 N_A_2227_367#_c_1370_n N_Q_c_1631_n 0.00434396f $X=11.315 $Y=0.865 $X2=0
+ $Y2=0
cc_872 N_A_2227_367#_c_1371_n N_Q_c_1631_n 0.026332f $X=11.89 $Y=1.51 $X2=0
+ $Y2=0
cc_873 N_A_2227_367#_c_1373_n N_Q_c_1631_n 0.00664526f $X=11.925 $Y=1.42 $X2=0
+ $Y2=0
cc_874 N_A_2227_367#_c_1374_n N_Q_c_1631_n 0.00248293f $X=11.925 $Y=1.345 $X2=0
+ $Y2=0
cc_875 N_A_2227_367#_c_1370_n N_VGND_c_1656_n 0.0156172f $X=11.315 $Y=0.865
+ $X2=0 $Y2=0
cc_876 N_A_2227_367#_c_1370_n N_VGND_c_1657_n 0.0363594f $X=11.315 $Y=0.865
+ $X2=0 $Y2=0
cc_877 N_A_2227_367#_c_1371_n N_VGND_c_1657_n 0.0227997f $X=11.89 $Y=1.51 $X2=0
+ $Y2=0
cc_878 N_A_2227_367#_c_1373_n N_VGND_c_1657_n 0.00562998f $X=11.925 $Y=1.42
+ $X2=0 $Y2=0
cc_879 N_A_2227_367#_c_1374_n N_VGND_c_1657_n 0.00543982f $X=11.925 $Y=1.345
+ $X2=0 $Y2=0
cc_880 N_A_2227_367#_c_1367_n N_VGND_c_1659_n 0.00751159f $X=12.48 $Y=1.345
+ $X2=0 $Y2=0
cc_881 N_A_2227_367#_c_1370_n N_VGND_c_1667_n 0.0050336f $X=11.315 $Y=0.865
+ $X2=0 $Y2=0
cc_882 N_A_2227_367#_c_1367_n N_VGND_c_1668_n 0.00559701f $X=12.48 $Y=1.345
+ $X2=0 $Y2=0
cc_883 N_A_2227_367#_c_1374_n N_VGND_c_1668_n 0.00558361f $X=11.925 $Y=1.345
+ $X2=0 $Y2=0
cc_884 N_A_2227_367#_c_1367_n N_VGND_c_1674_n 0.00537853f $X=12.48 $Y=1.345
+ $X2=0 $Y2=0
cc_885 N_A_2227_367#_c_1370_n N_VGND_c_1674_n 0.00944273f $X=11.315 $Y=0.865
+ $X2=0 $Y2=0
cc_886 N_A_2227_367#_c_1374_n N_VGND_c_1674_n 0.00537853f $X=11.925 $Y=1.345
+ $X2=0 $Y2=0
cc_887 N_VPWR_c_1419_n N_A_507_125#_M1008_d 0.002703f $X=12.72 $Y=3.33 $X2=0
+ $Y2=0
cc_888 N_VPWR_c_1422_n N_A_507_125#_c_1574_n 4.04269e-19 $X=2.195 $Y=2.82 $X2=0
+ $Y2=0
cc_889 N_VPWR_c_1438_n N_A_507_125#_c_1592_n 0.0133682f $X=3.84 $Y=3.125 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_1419_n N_A_507_125#_c_1592_n 0.0110139f $X=12.72 $Y=3.33 $X2=0
+ $Y2=0
cc_891 N_VPWR_c_1419_n A_701_535# 0.0029401f $X=12.72 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_892 N_VPWR_c_1419_n A_1288_451# 0.00168878f $X=12.72 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_893 N_VPWR_c_1419_n N_Q_N_M1004_s 0.00380103f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_894 N_VPWR_c_1426_n N_Q_N_c_1611_n 0.0437697f $X=10.845 $Y=1.98 $X2=0 $Y2=0
cc_895 N_VPWR_c_1434_n N_Q_N_c_1611_n 0.0143246f $X=10.645 $Y=3.33 $X2=0 $Y2=0
cc_896 N_VPWR_c_1419_n N_Q_N_c_1611_n 0.00916141f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_897 N_VPWR_c_1419_n N_Q_M1001_s 0.00345315f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_898 N_VPWR_c_1429_n N_Q_c_1631_n 0.00153478f $X=12.695 $Y=1.98 $X2=0 $Y2=0
cc_899 N_VPWR_c_1436_n N_Q_c_1631_n 0.0144039f $X=12.56 $Y=3.33 $X2=0 $Y2=0
cc_900 N_VPWR_c_1419_n N_Q_c_1631_n 0.00944728f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_901 N_VPWR_c_1429_n N_VGND_c_1659_n 0.0121422f $X=12.695 $Y=1.98 $X2=0 $Y2=0
cc_902 N_Q_N_c_1611_n N_VGND_c_1656_n 0.0324873f $X=10.36 $Y=0.42 $X2=0 $Y2=0
cc_903 N_Q_N_c_1611_n N_VGND_c_1666_n 0.0142265f $X=10.36 $Y=0.42 $X2=0 $Y2=0
cc_904 N_Q_N_M1015_d N_VGND_c_1674_n 0.00362709f $X=10.22 $Y=0.235 $X2=0 $Y2=0
cc_905 N_Q_N_c_1611_n N_VGND_c_1674_n 0.00925289f $X=10.36 $Y=0.42 $X2=0 $Y2=0
cc_906 N_Q_c_1631_n N_VGND_c_1657_n 0.0303144f $X=12.265 $Y=0.54 $X2=0 $Y2=0
cc_907 N_Q_c_1631_n N_VGND_c_1659_n 0.00306956f $X=12.265 $Y=0.54 $X2=0 $Y2=0
cc_908 N_Q_c_1631_n N_VGND_c_1668_n 0.00985247f $X=12.265 $Y=0.54 $X2=0 $Y2=0
cc_909 N_Q_c_1631_n N_VGND_c_1674_n 0.00883833f $X=12.265 $Y=0.54 $X2=0 $Y2=0
cc_910 N_VGND_c_1674_n N_A_1173_125#_M1026_d 0.00213412f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_911 N_VGND_c_1652_n N_A_1173_125#_c_1795_n 0.0263517f $X=5.575 $Y=0.87 $X2=0
+ $Y2=0
cc_912 N_VGND_c_1652_n N_A_1173_125#_c_1796_n 0.0176923f $X=5.575 $Y=0.87 $X2=0
+ $Y2=0
cc_913 N_VGND_c_1665_n N_A_1173_125#_c_1796_n 0.017523f $X=8.72 $Y=0 $X2=0 $Y2=0
cc_914 N_VGND_c_1674_n N_A_1173_125#_c_1796_n 0.00902319f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_915 N_VGND_c_1665_n N_A_1173_125#_c_1797_n 0.0955147f $X=8.72 $Y=0 $X2=0
+ $Y2=0
cc_916 N_VGND_c_1674_n N_A_1173_125#_c_1797_n 0.0540983f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_917 N_VGND_c_1653_n N_A_1280_159#_c_1824_n 0.0104909f $X=8.885 $Y=0.665 $X2=0
+ $Y2=0
cc_918 N_VGND_c_1665_n N_A_1280_159#_c_1824_n 0.007665f $X=8.72 $Y=0 $X2=0 $Y2=0
cc_919 N_VGND_c_1674_n N_A_1280_159#_c_1824_n 0.0106464f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_920 N_VGND_c_1665_n N_A_1280_159#_c_1825_n 0.00345594f $X=8.72 $Y=0 $X2=0
+ $Y2=0
cc_921 N_VGND_c_1674_n N_A_1280_159#_c_1825_n 0.00747751f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_922 N_A_1173_125#_c_1795_n N_A_1280_159#_c_1822_n 0.0139722f $X=6.005 $Y=0.83
+ $X2=0 $Y2=0
cc_923 N_A_1173_125#_c_1795_n N_A_1280_159#_c_1823_n 0.0134196f $X=6.005 $Y=0.83
+ $X2=0 $Y2=0
cc_924 N_A_1173_125#_c_1797_n N_A_1280_159#_c_1823_n 0.0237422f $X=7.575 $Y=0.37
+ $X2=0 $Y2=0
cc_925 N_A_1173_125#_M1026_d N_A_1280_159#_c_1825_n 0.0106867f $X=7.34 $Y=0.575
+ $X2=0 $Y2=0
cc_926 N_A_1173_125#_c_1797_n N_A_1280_159#_c_1825_n 0.0718422f $X=7.575 $Y=0.37
+ $X2=0 $Y2=0
