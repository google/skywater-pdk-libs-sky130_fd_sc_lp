# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xor3_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__xor3_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.605000 1.315000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.002000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.775000 1.550000 3.235000 1.565000 ;
        RECT 2.775000 1.565000 4.425000 1.895000 ;
        RECT 3.615000 1.155000 3.945000 1.565000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.245000 1.180000 9.955000 1.565000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.125000 2.095000 10.925000 2.265000 ;
        RECT 10.125000 2.265000 10.455000 3.065000 ;
        RECT 10.675000 0.685000 10.925000 2.095000 ;
        RECT 10.675000 2.265000 10.925000 2.890000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.265000  0.545000  0.595000 1.095000 ;
      RECT  0.265000  1.095000  1.735000 1.425000 ;
      RECT  0.265000  1.425000  0.655000 2.330000 ;
      RECT  0.265000  2.330000  1.535000 2.500000 ;
      RECT  0.265000  2.500000  0.655000 3.065000 ;
      RECT  0.855000  2.680000  1.185000 3.245000 ;
      RECT  1.055000  0.085000  1.385000 0.915000 ;
      RECT  1.365000  2.500000  1.535000 2.895000 ;
      RECT  1.365000  2.895000  3.840000 3.065000 ;
      RECT  1.565000  0.265000  4.150000 0.435000 ;
      RECT  1.565000  0.435000  1.735000 1.095000 ;
      RECT  1.915000  0.810000  2.845000 1.005000 ;
      RECT  1.915000  1.005000  2.245000 2.715000 ;
      RECT  2.425000  1.185000  3.435000 1.355000 ;
      RECT  2.425000  1.355000  2.595000 2.075000 ;
      RECT  2.425000  2.075000  4.190000 2.245000 ;
      RECT  2.425000  2.245000  2.775000 2.715000 ;
      RECT  2.515000  0.625000  2.845000 0.810000 ;
      RECT  3.105000  0.615000  3.435000 1.185000 ;
      RECT  3.510000  2.425000  3.840000 2.895000 ;
      RECT  3.820000  0.435000  4.150000 0.685000 ;
      RECT  4.020000  2.245000  4.190000 2.895000 ;
      RECT  4.020000  2.895000  6.080000 3.065000 ;
      RECT  4.330000  0.310000  4.660000 1.035000 ;
      RECT  4.330000  1.035000  4.500000 1.215000 ;
      RECT  4.330000  1.215000  4.775000 1.385000 ;
      RECT  4.390000  2.310000  4.775000 2.715000 ;
      RECT  4.605000  1.385000  4.775000 2.310000 ;
      RECT  4.840000  0.575000  5.170000 1.035000 ;
      RECT  4.955000  1.035000  5.170000 1.040000 ;
      RECT  4.955000  1.040000  5.125000 1.960000 ;
      RECT  4.955000  1.960000  5.250000 2.715000 ;
      RECT  5.305000  1.450000  5.730000 1.780000 ;
      RECT  5.350000  0.265000  5.730000 0.425000 ;
      RECT  5.350000  0.425000  6.100000 0.595000 ;
      RECT  5.480000  1.780000  5.730000 2.715000 ;
      RECT  5.560000  0.595000  6.100000 0.885000 ;
      RECT  5.560000  0.885000  5.730000 1.450000 ;
      RECT  5.910000  1.150000  7.290000 1.320000 ;
      RECT  5.910000  1.320000  6.080000 2.895000 ;
      RECT  6.260000  1.960000  6.430000 3.245000 ;
      RECT  6.560000  0.085000  6.890000 0.885000 ;
      RECT  6.615000  1.320000  6.785000 2.010000 ;
      RECT  6.615000  2.010000  7.070000 3.050000 ;
      RECT  6.965000  1.500000  8.135000 1.565000 ;
      RECT  6.965000  1.565000  7.640000 1.830000 ;
      RECT  7.120000  0.595000  7.450000 1.055000 ;
      RECT  7.120000  1.055000  7.290000 1.150000 ;
      RECT  7.270000  2.010000  7.600000 2.895000 ;
      RECT  7.270000  2.895000  9.415000 3.065000 ;
      RECT  7.470000  1.235000  8.135000 1.500000 ;
      RECT  7.630000  0.265000 10.145000 0.435000 ;
      RECT  7.630000  0.435000  7.960000 1.055000 ;
      RECT  7.800000  2.010000  8.485000 2.715000 ;
      RECT  8.140000  0.615000  8.485000 1.055000 ;
      RECT  8.315000  1.055000  8.485000 2.010000 ;
      RECT  8.665000  0.685000  9.065000 2.715000 ;
      RECT  9.245000  1.745000 10.465000 1.915000 ;
      RECT  9.245000  1.915000  9.415000 2.895000 ;
      RECT  9.595000  2.095000  9.925000 3.245000 ;
      RECT  9.775000  0.775000 10.495000 1.000000 ;
      RECT  9.870000  0.435000 10.145000 0.595000 ;
      RECT 10.135000  1.235000 10.465000 1.745000 ;
      RECT 10.325000  0.085000 10.495000 0.775000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  0.840000  2.245000 1.010000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  2.320000  4.645000 2.490000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  0.840000  5.125000 1.010000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  2.320000  8.005000 2.490000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
    LAYER met1 ;
      RECT 2.015000 0.810000 2.305000 0.855000 ;
      RECT 2.015000 0.855000 5.185000 0.995000 ;
      RECT 2.015000 0.995000 2.305000 1.040000 ;
      RECT 4.415000 2.290000 4.705000 2.335000 ;
      RECT 4.415000 2.335000 8.065000 2.475000 ;
      RECT 4.415000 2.475000 4.705000 2.520000 ;
      RECT 4.895000 0.810000 5.185000 0.855000 ;
      RECT 4.895000 0.995000 5.185000 1.040000 ;
      RECT 7.775000 2.290000 8.065000 2.335000 ;
      RECT 7.775000 2.475000 8.065000 2.520000 ;
  END
END sky130_fd_sc_lp__xor3_lp
END LIBRARY
