* File: sky130_fd_sc_lp__a2111o_0.pex.spice
* Created: Fri Aug 28 09:45:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111O_0%A_80_159# 1 2 3 11 14 18 20 21 22 23 25 26
+ 29 33 35 39 43 44
c86 29 0 2.86757e-20 $X=1.27 $Y=2.525
c87 25 0 1.24001e-19 $X=1.105 $Y=2.14
r88 43 46 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=0.96
+ $X2=0.605 $Y2=0.795
r89 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.645
+ $Y=0.96 $X2=0.645 $Y2=0.96
r90 37 39 15.8178 $w=2.53e-07 $l=3.5e-07 $layer=LI1_cond $X=2.617 $Y=0.795
+ $X2=2.617 $Y2=0.445
r91 36 44 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.51 $Y=0.88
+ $X2=1.377 $Y2=0.88
r92 35 37 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=2.49 $Y=0.88
+ $X2=2.617 $Y2=0.795
r93 35 36 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=2.49 $Y=0.88
+ $X2=1.51 $Y2=0.88
r94 31 44 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.377 $Y=0.795
+ $X2=1.377 $Y2=0.88
r95 31 33 15.2209 $w=2.63e-07 $l=3.5e-07 $layer=LI1_cond $X=1.377 $Y=0.795
+ $X2=1.377 $Y2=0.445
r96 27 29 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=1.24 $Y=2.225 $X2=1.24
+ $Y2=2.525
r97 25 27 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.105 $Y=2.14
+ $X2=1.24 $Y2=2.225
r98 25 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.105 $Y=2.14
+ $X2=0.81 $Y2=2.14
r99 24 42 4.53113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.81 $Y=0.88
+ $X2=0.672 $Y2=0.88
r100 23 44 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.245 $Y=0.88
+ $X2=1.377 $Y2=0.88
r101 23 24 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.245 $Y=0.88
+ $X2=0.81 $Y2=0.88
r102 22 26 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=0.672 $Y=2.055
+ $X2=0.81 $Y2=2.14
r103 21 42 2.79091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.672 $Y=0.965
+ $X2=0.672 $Y2=0.88
r104 21 22 45.6786 $w=2.73e-07 $l=1.09e-06 $layer=LI1_cond $X=0.672 $Y=0.965
+ $X2=0.672 $Y2=2.055
r105 18 46 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.735 $Y=0.445
+ $X2=0.735 $Y2=0.795
r106 14 20 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=0.475 $Y=2.735
+ $X2=0.475 $Y2=1.465
r107 11 20 51.3336 $w=4.1e-07 $l=2.05e-07 $layer=POLY_cond $X=0.605 $Y=1.26
+ $X2=0.605 $Y2=1.465
r108 10 43 5.42589 $w=4.1e-07 $l=4e-08 $layer=POLY_cond $X=0.605 $Y=1 $X2=0.605
+ $Y2=0.96
r109 10 11 35.2683 $w=4.1e-07 $l=2.6e-07 $layer=POLY_cond $X=0.605 $Y=1
+ $X2=0.605 $Y2=1.26
r110 3 29 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=2.38 $X2=1.27 $Y2=2.525
r111 2 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.62 $Y2=0.445
r112 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.24
+ $Y=0.235 $X2=1.38 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_0%D1 3 6 7 9 12 13 16 18 19 23
c54 3 0 1.94051e-19 $X=1.165 $Y=0.445
r55 18 19 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.177 $Y=1.295
+ $X2=1.177 $Y2=1.665
r56 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.215
+ $Y=1.37 $X2=1.215 $Y2=1.37
r57 14 16 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.305 $Y=2.195
+ $X2=1.485 $Y2=2.195
r58 12 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.215 $Y=1.71
+ $X2=1.215 $Y2=1.37
r59 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=1.71
+ $X2=1.215 $Y2=1.875
r60 11 23 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=1.205
+ $X2=1.215 $Y2=1.37
r61 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.485 $Y=2.27
+ $X2=1.485 $Y2=2.195
r62 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.485 $Y=2.27
+ $X2=1.485 $Y2=2.7
r63 6 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.305 $Y=2.12
+ $X2=1.305 $Y2=2.195
r64 6 13 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.305 $Y=2.12
+ $X2=1.305 $Y2=1.875
r65 3 11 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.165 $Y=0.445
+ $X2=1.165 $Y2=1.205
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_0%C1 3 6 11 15 17 18 19 20 21 22 29 31
c55 18 0 3.57794e-19 $X=1.68 $Y=1.295
c56 11 0 1.52676e-19 $X=1.875 $Y=2.7
r57 29 31 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.375
+ $X2=1.77 $Y2=1.21
r58 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.785
+ $Y=1.375 $X2=1.785 $Y2=1.375
r59 21 22 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.707 $Y=2.405
+ $X2=1.707 $Y2=2.775
r60 20 21 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.707 $Y=2.035
+ $X2=1.707 $Y2=2.405
r61 19 20 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.707 $Y=1.665
+ $X2=1.707 $Y2=2.035
r62 19 30 10.2833 $w=3.23e-07 $l=2.9e-07 $layer=LI1_cond $X=1.707 $Y=1.665
+ $X2=1.707 $Y2=1.375
r63 18 30 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=1.707 $Y=1.295
+ $X2=1.707 $Y2=1.375
r64 13 15 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.595 $Y=0.92
+ $X2=1.71 $Y2=0.92
r65 11 17 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.875 $Y=2.7
+ $X2=1.875 $Y2=1.88
r66 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.71 $Y=0.995
+ $X2=1.71 $Y2=0.92
r67 7 31 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.71 $Y=0.995
+ $X2=1.71 $Y2=1.21
r68 6 17 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.77 $Y=1.7 $X2=1.77
+ $Y2=1.88
r69 5 29 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.77 $Y=1.39 $X2=1.77
+ $Y2=1.375
r70 5 6 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.77 $Y=1.39 $X2=1.77
+ $Y2=1.7
r71 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.595 $Y=0.845
+ $X2=1.595 $Y2=0.92
r72 1 3 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.595 $Y=0.845 $X2=1.595
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_0%B1 3 7 11 12 13 14 15 16 23 34
c52 13 0 9.52314e-20 $X=2.16 $Y=1.295
c53 7 0 2.63615e-19 $X=2.405 $Y=0.445
r54 25 34 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=2.225 $Y=2.085
+ $X2=2.225 $Y2=2.035
r55 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.325
+ $Y=1.375 $X2=2.325 $Y2=1.375
r56 15 16 13.5904 $w=2.72e-07 $l=3.03e-07 $layer=LI1_cond $X=2.225 $Y=2.102
+ $X2=2.225 $Y2=2.405
r57 15 25 1.44022 $w=3.7e-07 $l=1.7e-08 $layer=LI1_cond $X=2.225 $Y=2.102
+ $X2=2.225 $Y2=2.085
r58 15 34 0.560648 $w=3.68e-07 $l=1.8e-08 $layer=LI1_cond $X=2.225 $Y=2.017
+ $X2=2.225 $Y2=2.035
r59 14 15 10.9638 $w=3.68e-07 $l=3.52e-07 $layer=LI1_cond $X=2.225 $Y=1.665
+ $X2=2.225 $Y2=2.017
r60 14 24 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.225 $Y=1.665
+ $X2=2.225 $Y2=1.375
r61 13 24 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=2.225 $Y=1.295
+ $X2=2.225 $Y2=1.375
r62 11 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.325 $Y=1.715
+ $X2=2.325 $Y2=1.375
r63 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.715
+ $X2=2.325 $Y2=1.88
r64 10 23 44.4756 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.21
+ $X2=2.325 $Y2=1.375
r65 7 10 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.405 $Y=0.445
+ $X2=2.405 $Y2=1.21
r66 3 12 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.265 $Y=2.7
+ $X2=2.265 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_0%A1 1 2 5 9 11 12 13 14
c51 12 0 9.98724e-20 $X=3.12 $Y=0.925
c52 9 0 1.37156e-19 $X=2.91 $Y=2.7
c53 5 0 9.52314e-20 $X=2.835 $Y=0.445
r54 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3 $Y=1.335
+ $X2=3 $Y2=1.335
r55 14 20 11.3524 $w=3.33e-07 $l=3.3e-07 $layer=LI1_cond $X=3.082 $Y=1.665
+ $X2=3.082 $Y2=1.335
r56 13 20 1.37605 $w=3.33e-07 $l=4e-08 $layer=LI1_cond $X=3.082 $Y=1.295
+ $X2=3.082 $Y2=1.335
r57 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.082 $Y=0.925
+ $X2=3.082 $Y2=1.295
r58 9 11 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.91 $Y=2.7 $X2=2.91
+ $Y2=1.84
r59 3 19 40.7576 $w=4.29e-07 $l=2.18952e-07 $layer=POLY_cond $X=2.835 $Y=1.165
+ $X2=2.947 $Y2=1.335
r60 3 5 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.835 $Y=1.165
+ $X2=2.835 $Y2=0.445
r61 2 11 42.3913 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=2.947 $Y=1.623
+ $X2=2.947 $Y2=1.84
r62 1 19 5.76184 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=2.947 $Y=1.387
+ $X2=2.947 $Y2=1.335
r63 1 2 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=2.947 $Y=1.387
+ $X2=2.947 $Y2=1.623
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_0%A2 1 3 6 9 13 17 20 21 22 23 28
c38 21 0 2.46084e-20 $X=3.6 $Y=0.925
r39 22 23 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=1.295
+ $X2=3.587 $Y2=1.665
r40 21 22 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=0.925
+ $X2=3.587 $Y2=1.295
r41 21 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.005 $X2=3.57 $Y2=1.005
r42 19 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.57 $Y=1.345
+ $X2=3.57 $Y2=1.005
r43 19 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.345
+ $X2=3.57 $Y2=1.51
r44 15 17 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=3.34 $Y=2.155
+ $X2=3.48 $Y2=2.155
r45 13 28 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.57 $Y=0.93
+ $X2=3.57 $Y2=1.005
r46 10 13 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=3.195 $Y=0.855
+ $X2=3.57 $Y2=0.855
r47 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.48 $Y=2.08 $X2=3.48
+ $Y2=2.155
r48 9 20 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.48 $Y=2.08 $X2=3.48
+ $Y2=1.51
r49 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.34 $Y=2.23 $X2=3.34
+ $Y2=2.155
r50 4 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.34 $Y=2.23 $X2=3.34
+ $Y2=2.7
r51 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.195 $Y=0.78
+ $X2=3.195 $Y2=0.855
r52 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.195 $Y=0.78
+ $X2=3.195 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_0%X 1 2 7 8 9 10 11 12 13 44
r16 22 39 1.70047 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.225 $Y=0.61
+ $X2=0.225 $Y2=0.445
r17 13 35 8.84912 $w=2.78e-07 $l=2.15e-07 $layer=LI1_cond $X=0.225 $Y=2.775
+ $X2=0.225 $Y2=2.56
r18 12 35 6.3796 $w=2.78e-07 $l=1.55e-07 $layer=LI1_cond $X=0.225 $Y=2.405
+ $X2=0.225 $Y2=2.56
r19 11 12 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=2.035
+ $X2=0.225 $Y2=2.405
r20 10 11 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=2.035
r21 9 10 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r22 8 9 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r23 7 44 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=0.445 $X2=0.52
+ $Y2=0.445
r24 7 39 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.24 $Y=0.445
+ $X2=0.225 $Y2=0.445
r25 7 8 12.3476 $w=2.78e-07 $l=3e-07 $layer=LI1_cond $X=0.225 $Y=0.625 $X2=0.225
+ $Y2=0.925
r26 7 22 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=0.225 $Y=0.625
+ $X2=0.225 $Y2=0.61
r27 2 35 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.415 $X2=0.26 $Y2=2.56
r28 1 44 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.395
+ $Y=0.235 $X2=0.52 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_0%VPWR 1 2 9 13 15 17 22 32 33 36 39
r44 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r48 30 39 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.255 $Y=3.33
+ $X2=3.122 $Y2=3.33
r49 30 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.255 $Y=3.33
+ $X2=3.6 $Y2=3.33
r50 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 23 36 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.695 $Y2=3.33
r56 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 22 39 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.99 $Y=3.33
+ $X2=3.122 $Y2=3.33
r58 22 28 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.99 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 17 36 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.695 $Y2=3.33
r62 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 11 39 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.122 $Y=3.245
+ $X2=3.122 $Y2=3.33
r66 11 13 30.8768 $w=2.63e-07 $l=7.1e-07 $layer=LI1_cond $X=3.122 $Y=3.245
+ $X2=3.122 $Y2=2.535
r67 7 36 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=3.33
r68 7 9 24.3093 $w=3.18e-07 $l=6.75e-07 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=2.57
r69 2 13 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=2.38 $X2=3.125 $Y2=2.535
r70 1 9 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.415 $X2=0.69 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_0%A_468_476# 1 2 10 11 12 15 20
c34 15 0 1.12547e-19 $X=3.555 $Y=2.525
r35 18 20 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.48 $Y=2.875
+ $X2=2.7 $Y2=2.875
r36 13 15 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=3.572 $Y=2.19
+ $X2=3.572 $Y2=2.525
r37 11 13 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=3.425 $Y=2.105
+ $X2=3.572 $Y2=2.19
r38 11 12 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.425 $Y=2.105
+ $X2=2.82 $Y2=2.105
r39 8 20 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=2.71 $X2=2.7
+ $Y2=2.875
r40 8 10 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=2.7 $Y=2.71 $X2=2.7
+ $Y2=2.525
r41 7 12 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.7 $Y=2.19
+ $X2=2.82 $Y2=2.105
r42 7 10 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=2.7 $Y=2.19 $X2=2.7
+ $Y2=2.525
r43 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.415
+ $Y=2.38 $X2=3.555 $Y2=2.525
r44 1 18 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=2.38 $X2=2.48 $Y2=2.875
r45 1 10 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=2.38 $X2=2.695 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_0%VGND 1 2 3 12 16 18 20 21 22 28 36 42 45
r49 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 41 42 10.1707 $w=6.93e-07 $l=1.3e-07 $layer=LI1_cond $X=2.19 $Y=0.262
+ $X2=2.32 $Y2=0.262
r51 38 41 0.516293 $w=6.93e-07 $l=3e-08 $layer=LI1_cond $X=2.16 $Y=0.262
+ $X2=2.19 $Y2=0.262
r52 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r53 34 38 8.26068 $w=6.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.262
+ $X2=2.16 $Y2=0.262
r54 34 36 7.9334 $w=6.93e-07 $l=4.17027e-08 $layer=LI1_cond $X=1.68 $Y=0.262
+ $X2=1.68 $Y2=0.262
r55 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 32 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r57 32 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r58 31 42 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=2.32
+ $Y2=0
r59 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r60 28 44 4.92749 $w=1.7e-07 $l=3.12e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.527
+ $Y2=0
r61 28 31 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.12
+ $Y2=0
r62 26 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r63 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r64 22 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r65 22 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r66 20 25 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.72
+ $Y2=0
r67 20 21 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.945
+ $Y2=0
r68 16 44 3.2692 $w=3.8e-07 $l=1.58915e-07 $layer=LI1_cond $X=3.405 $Y=0.085
+ $X2=3.527 $Y2=0
r69 16 18 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.405 $Y=0.085
+ $X2=3.405 $Y2=0.445
r70 15 21 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=0.945
+ $Y2=0
r71 15 36 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=1.68
+ $Y2=0
r72 10 21 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.945 $Y=0.085
+ $X2=0.945 $Y2=0
r73 10 12 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.945 $Y=0.085
+ $X2=0.945 $Y2=0.445
r74 3 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.27
+ $Y=0.235 $X2=3.41 $Y2=0.445
r75 2 41 91 $w=1.7e-07 $l=6.16117e-07 $layer=licon1_NDIFF $count=2 $X=1.67
+ $Y=0.235 $X2=2.19 $Y2=0.445
r76 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.81
+ $Y=0.235 $X2=0.95 $Y2=0.445
.ends

