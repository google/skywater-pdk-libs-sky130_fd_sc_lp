* File: sky130_fd_sc_lp__o22ai_lp.pxi.spice
* Created: Wed Sep  2 10:20:57 2020
* 
x_PM_SKY130_FD_SC_LP__O22AI_LP%B1 N_B1_M1005_g N_B1_M1007_g N_B1_c_61_n
+ N_B1_c_62_n B1 N_B1_c_64_n N_B1_c_65_n PM_SKY130_FD_SC_LP__O22AI_LP%B1
x_PM_SKY130_FD_SC_LP__O22AI_LP%B2 N_B2_M1000_g N_B2_M1004_g B2 N_B2_c_99_n
+ PM_SKY130_FD_SC_LP__O22AI_LP%B2
x_PM_SKY130_FD_SC_LP__O22AI_LP%A2 N_A2_M1003_g N_A2_M1006_g A2 N_A2_c_134_n
+ N_A2_c_135_n N_A2_c_136_n PM_SKY130_FD_SC_LP__O22AI_LP%A2
x_PM_SKY130_FD_SC_LP__O22AI_LP%A1 N_A1_M1002_g N_A1_M1001_g N_A1_c_170_n
+ N_A1_c_171_n N_A1_c_172_n A1 N_A1_c_173_n N_A1_c_174_n
+ PM_SKY130_FD_SC_LP__O22AI_LP%A1
x_PM_SKY130_FD_SC_LP__O22AI_LP%VPWR N_VPWR_M1005_s N_VPWR_M1001_d N_VPWR_c_201_n
+ N_VPWR_c_202_n N_VPWR_c_203_n N_VPWR_c_204_n N_VPWR_c_205_n N_VPWR_c_206_n
+ N_VPWR_c_207_n VPWR N_VPWR_c_200_n PM_SKY130_FD_SC_LP__O22AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O22AI_LP%Y N_Y_M1007_d N_Y_M1000_d N_Y_c_233_n N_Y_c_234_n
+ N_Y_c_235_n N_Y_c_237_n N_Y_c_238_n N_Y_c_250_n Y Y
+ PM_SKY130_FD_SC_LP__O22AI_LP%Y
x_PM_SKY130_FD_SC_LP__O22AI_LP%A_70_101# N_A_70_101#_M1007_s N_A_70_101#_M1004_d
+ N_A_70_101#_M1002_d N_A_70_101#_c_279_n N_A_70_101#_c_280_n
+ N_A_70_101#_c_281_n N_A_70_101#_c_282_n N_A_70_101#_c_283_n
+ N_A_70_101#_c_288_n N_A_70_101#_c_289_n N_A_70_101#_c_284_n
+ N_A_70_101#_c_285_n N_A_70_101#_c_286_n PM_SKY130_FD_SC_LP__O22AI_LP%A_70_101#
x_PM_SKY130_FD_SC_LP__O22AI_LP%VGND N_VGND_M1003_d N_VGND_c_341_n VGND
+ N_VGND_c_342_n N_VGND_c_343_n N_VGND_c_344_n N_VGND_c_345_n
+ PM_SKY130_FD_SC_LP__O22AI_LP%VGND
cc_1 VNB N_B1_c_61_n 0.017291f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1
cc_2 VNB N_B1_c_62_n 0.0121797f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.15
cc_3 VNB B1 0.0016928f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_B1_c_64_n 0.0209338f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.615
cc_5 VNB N_B1_c_65_n 0.0179336f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.45
cc_6 VNB N_B2_M1004_g 0.0389534f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1
cc_7 VNB B2 0.00357468f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.715
cc_8 VNB N_B2_c_99_n 0.019572f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_9 VNB N_A2_c_134_n 0.0783242f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.15
cc_10 VNB N_A2_c_135_n 0.00313393f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_11 VNB N_A2_c_136_n 0.0192201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_c_170_n 0.0239601f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.715
cc_13 VNB N_A1_c_171_n 0.026086f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1
cc_14 VNB N_A1_c_172_n 0.00887541f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.15
cc_15 VNB N_A1_c_173_n 0.0178431f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.615
cc_16 VNB N_A1_c_174_n 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.615
cc_17 VNB N_VPWR_c_200_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_233_n 0.0188537f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.715
cc_19 VNB N_Y_c_234_n 0.022138f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.715
cc_20 VNB N_Y_c_235_n 0.0149163f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1
cc_21 VNB N_A_70_101#_c_279_n 0.0196638f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_22 VNB N_A_70_101#_c_280_n 0.0143962f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.615
cc_23 VNB N_A_70_101#_c_281_n 0.0106412f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.615
cc_24 VNB N_A_70_101#_c_282_n 6.89024e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_70_101#_c_283_n 0.00606562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_70_101#_c_284_n 0.0264477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_70_101#_c_285_n 0.0382371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_70_101#_c_286_n 0.00827576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_341_n 0.0179687f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.45
cc_30 VNB N_VGND_c_342_n 0.0508107f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1
cc_31 VNB N_VGND_c_343_n 0.0333497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_344_n 0.236451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_345_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_B1_M1005_g 0.0383824f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.595
cc_35 VPB B1 7.47102e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_36 VPB N_B1_c_64_n 0.0119057f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.615
cc_37 VPB N_B2_M1000_g 0.0351053f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.595
cc_38 VPB B2 0.00110633f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.715
cc_39 VPB N_B2_c_99_n 0.0110927f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_40 VPB N_A2_M1006_g 0.0434758f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.45
cc_41 VPB N_A2_c_134_n 0.015211f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.15
cc_42 VPB N_A2_c_135_n 0.00313998f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_43 VPB N_A1_M1001_g 0.0505261f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.45
cc_44 VPB N_A1_c_172_n 0.00611381f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.15
cc_45 VPB N_A1_c_174_n 7.56276e-19 $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.615
cc_46 VPB N_VPWR_c_201_n 0.032591f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.715
cc_47 VPB N_VPWR_c_202_n 0.0354389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_203_n 0.0113717f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.615
cc_49 VPB N_VPWR_c_204_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.45
cc_50 VPB N_VPWR_c_205_n 0.0113717f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.78
cc_51 VPB N_VPWR_c_206_n 0.0601852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_207_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_200_n 0.0600214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_Y_c_233_n 0.0149425f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.715
cc_55 VPB N_Y_c_237_n 0.0152699f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.15
cc_56 VPB N_Y_c_238_n 0.0132327f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_57 VPB N_A_70_101#_c_283_n 0.00183801f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_70_101#_c_288_n 0.0562692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_70_101#_c_289_n 0.00266732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_70_101#_c_285_n 0.0114395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 N_B1_M1005_g N_B2_M1000_g 0.0481014f $X=0.72 $Y=2.595 $X2=0 $Y2=0
cc_62 N_B1_c_61_n N_B2_M1004_g 0.0191111f $X=0.78 $Y=1 $X2=0 $Y2=0
cc_63 N_B1_c_65_n N_B2_M1004_g 0.0134693f $X=0.68 $Y=1.45 $X2=0 $Y2=0
cc_64 B1 B2 0.0188003f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_65 N_B1_c_64_n B2 0.00121489f $X=0.68 $Y=1.615 $X2=0 $Y2=0
cc_66 B1 N_B2_c_99_n 0.00121489f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_67 N_B1_c_64_n N_B2_c_99_n 0.0481014f $X=0.68 $Y=1.615 $X2=0 $Y2=0
cc_68 N_B1_M1005_g N_VPWR_c_201_n 0.0227289f $X=0.72 $Y=2.595 $X2=0 $Y2=0
cc_69 N_B1_M1005_g N_VPWR_c_206_n 0.008763f $X=0.72 $Y=2.595 $X2=0 $Y2=0
cc_70 N_B1_M1005_g N_VPWR_c_200_n 0.0144563f $X=0.72 $Y=2.595 $X2=0 $Y2=0
cc_71 N_B1_M1005_g N_Y_c_233_n 0.00590404f $X=0.72 $Y=2.595 $X2=0 $Y2=0
cc_72 B1 N_Y_c_233_n 0.0237562f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_73 N_B1_c_64_n N_Y_c_233_n 0.00735127f $X=0.68 $Y=1.615 $X2=0 $Y2=0
cc_74 N_B1_c_65_n N_Y_c_233_n 0.00500796f $X=0.68 $Y=1.45 $X2=0 $Y2=0
cc_75 N_B1_c_62_n N_Y_c_234_n 0.00677362f $X=0.78 $Y=1.15 $X2=0 $Y2=0
cc_76 B1 N_Y_c_234_n 0.0228535f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_77 N_B1_c_64_n N_Y_c_234_n 0.00123714f $X=0.68 $Y=1.615 $X2=0 $Y2=0
cc_78 N_B1_c_65_n N_Y_c_234_n 0.00783751f $X=0.68 $Y=1.45 $X2=0 $Y2=0
cc_79 N_B1_M1005_g N_Y_c_237_n 0.02318f $X=0.72 $Y=2.595 $X2=0 $Y2=0
cc_80 B1 N_Y_c_237_n 0.022783f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_81 N_B1_c_64_n N_Y_c_237_n 5.5002e-19 $X=0.68 $Y=1.615 $X2=0 $Y2=0
cc_82 N_B1_c_61_n N_Y_c_250_n 0.00794847f $X=0.78 $Y=1 $X2=0 $Y2=0
cc_83 N_B1_c_62_n N_Y_c_250_n 0.00548272f $X=0.78 $Y=1.15 $X2=0 $Y2=0
cc_84 N_B1_M1005_g Y 0.00423856f $X=0.72 $Y=2.595 $X2=0 $Y2=0
cc_85 N_B1_c_61_n N_A_70_101#_c_279_n 0.0108472f $X=0.78 $Y=1 $X2=0 $Y2=0
cc_86 N_B1_c_61_n N_A_70_101#_c_280_n 0.00918035f $X=0.78 $Y=1 $X2=0 $Y2=0
cc_87 N_B1_c_62_n N_A_70_101#_c_280_n 3.92696e-19 $X=0.78 $Y=1.15 $X2=0 $Y2=0
cc_88 N_B1_c_61_n N_VGND_c_342_n 7.10185e-19 $X=0.78 $Y=1 $X2=0 $Y2=0
cc_89 N_B2_M1000_g N_A2_M1006_g 0.0256771f $X=1.21 $Y=2.595 $X2=0 $Y2=0
cc_90 B2 N_A2_c_134_n 3.70835e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_91 N_B2_c_99_n N_A2_c_134_n 0.0174296f $X=1.25 $Y=1.615 $X2=0 $Y2=0
cc_92 N_B2_M1004_g N_A2_c_136_n 0.0250388f $X=1.22 $Y=0.715 $X2=0 $Y2=0
cc_93 N_B2_M1000_g N_VPWR_c_201_n 0.00174029f $X=1.21 $Y=2.595 $X2=0 $Y2=0
cc_94 N_B2_M1000_g N_VPWR_c_206_n 0.00599594f $X=1.21 $Y=2.595 $X2=0 $Y2=0
cc_95 N_B2_M1000_g N_VPWR_c_200_n 0.0078732f $X=1.21 $Y=2.595 $X2=0 $Y2=0
cc_96 N_B2_M1004_g N_Y_c_234_n 0.00514826f $X=1.22 $Y=0.715 $X2=0 $Y2=0
cc_97 B2 N_Y_c_234_n 0.00668272f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_98 N_B2_c_99_n N_Y_c_234_n 4.5416e-19 $X=1.25 $Y=1.615 $X2=0 $Y2=0
cc_99 N_B2_M1004_g N_Y_c_250_n 0.00827463f $X=1.22 $Y=0.715 $X2=0 $Y2=0
cc_100 N_B2_M1000_g Y 0.0424805f $X=1.21 $Y=2.595 $X2=0 $Y2=0
cc_101 B2 Y 0.0200591f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_102 N_B2_c_99_n Y 2.91808e-19 $X=1.25 $Y=1.615 $X2=0 $Y2=0
cc_103 N_B2_M1004_g N_A_70_101#_c_280_n 0.0107384f $X=1.22 $Y=0.715 $X2=0 $Y2=0
cc_104 N_B2_M1004_g N_A_70_101#_c_282_n 0.00437741f $X=1.22 $Y=0.715 $X2=0 $Y2=0
cc_105 N_B2_M1000_g N_A_70_101#_c_283_n 0.00200769f $X=1.21 $Y=2.595 $X2=0 $Y2=0
cc_106 N_B2_M1004_g N_A_70_101#_c_283_n 0.00562145f $X=1.22 $Y=0.715 $X2=0 $Y2=0
cc_107 B2 N_A_70_101#_c_283_n 0.0237562f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_B2_c_99_n N_A_70_101#_c_283_n 0.00187395f $X=1.25 $Y=1.615 $X2=0 $Y2=0
cc_109 N_B2_M1000_g N_A_70_101#_c_289_n 0.00263659f $X=1.21 $Y=2.595 $X2=0 $Y2=0
cc_110 B2 N_A_70_101#_c_286_n 0.00235712f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_B2_c_99_n N_A_70_101#_c_286_n 4.16578e-19 $X=1.25 $Y=1.615 $X2=0 $Y2=0
cc_112 N_B2_M1004_g N_VGND_c_342_n 7.10185e-19 $X=1.22 $Y=0.715 $X2=0 $Y2=0
cc_113 N_A2_M1006_g N_A1_M1001_g 0.0373426f $X=1.78 $Y=2.595 $X2=0 $Y2=0
cc_114 N_A2_c_136_n N_A1_c_170_n 0.007872f $X=1.965 $Y=1.035 $X2=0 $Y2=0
cc_115 N_A2_c_134_n N_A1_c_173_n 0.0363669f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_116 N_A2_c_135_n N_A1_c_173_n 0.00246051f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_117 N_A2_c_134_n N_A1_c_174_n 0.00278026f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_118 N_A2_c_135_n N_A1_c_174_n 0.0381134f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_119 N_A2_M1006_g N_VPWR_c_206_n 0.00975641f $X=1.78 $Y=2.595 $X2=0 $Y2=0
cc_120 N_A2_M1006_g N_VPWR_c_200_n 0.0178616f $X=1.78 $Y=2.595 $X2=0 $Y2=0
cc_121 N_A2_c_136_n N_Y_c_250_n 2.50334e-19 $X=1.965 $Y=1.035 $X2=0 $Y2=0
cc_122 N_A2_M1006_g Y 0.00112784f $X=1.78 $Y=2.595 $X2=0 $Y2=0
cc_123 N_A2_c_136_n N_A_70_101#_c_280_n 0.00366333f $X=1.965 $Y=1.035 $X2=0
+ $Y2=0
cc_124 N_A2_c_136_n N_A_70_101#_c_282_n 0.00600164f $X=1.965 $Y=1.035 $X2=0
+ $Y2=0
cc_125 N_A2_M1006_g N_A_70_101#_c_283_n 0.00952929f $X=1.78 $Y=2.595 $X2=0 $Y2=0
cc_126 N_A2_c_134_n N_A_70_101#_c_283_n 0.0200488f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_127 N_A2_c_135_n N_A_70_101#_c_283_n 0.0457028f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_128 N_A2_c_136_n N_A_70_101#_c_283_n 0.00473841f $X=1.965 $Y=1.035 $X2=0
+ $Y2=0
cc_129 N_A2_M1006_g N_A_70_101#_c_288_n 0.0177928f $X=1.78 $Y=2.595 $X2=0 $Y2=0
cc_130 N_A2_c_134_n N_A_70_101#_c_288_n 0.00392401f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_131 N_A2_c_135_n N_A_70_101#_c_288_n 0.0250673f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_132 N_A2_M1006_g N_A_70_101#_c_289_n 0.00840428f $X=1.78 $Y=2.595 $X2=0 $Y2=0
cc_133 N_A2_c_136_n N_A_70_101#_c_286_n 0.00697638f $X=1.965 $Y=1.035 $X2=0
+ $Y2=0
cc_134 N_A2_c_134_n N_VGND_c_341_n 0.0025495f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_135 N_A2_c_135_n N_VGND_c_341_n 0.0273869f $X=2.11 $Y=1.2 $X2=0 $Y2=0
cc_136 N_A2_c_136_n N_VGND_c_341_n 0.00503743f $X=1.965 $Y=1.035 $X2=0 $Y2=0
cc_137 N_A2_c_136_n N_VGND_c_342_n 0.00181207f $X=1.965 $Y=1.035 $X2=0 $Y2=0
cc_138 N_A2_c_136_n N_VGND_c_344_n 0.00134369f $X=1.965 $Y=1.035 $X2=0 $Y2=0
cc_139 N_A1_M1001_g N_VPWR_c_202_n 0.0477254f $X=2.64 $Y=2.595 $X2=0 $Y2=0
cc_140 N_A1_M1001_g N_VPWR_c_206_n 0.008763f $X=2.64 $Y=2.595 $X2=0 $Y2=0
cc_141 N_A1_M1001_g N_VPWR_c_200_n 0.0152194f $X=2.64 $Y=2.595 $X2=0 $Y2=0
cc_142 N_A1_M1001_g N_A_70_101#_c_288_n 0.0247542f $X=2.64 $Y=2.595 $X2=0 $Y2=0
cc_143 N_A1_c_172_n N_A_70_101#_c_288_n 5.43485e-19 $X=2.68 $Y=1.705 $X2=0 $Y2=0
cc_144 N_A1_c_174_n N_A_70_101#_c_288_n 0.0241279f $X=2.68 $Y=1.2 $X2=0 $Y2=0
cc_145 N_A1_c_170_n N_A_70_101#_c_284_n 0.00686846f $X=2.68 $Y=1.035 $X2=0 $Y2=0
cc_146 N_A1_c_173_n N_A_70_101#_c_284_n 0.00115594f $X=2.68 $Y=1.2 $X2=0 $Y2=0
cc_147 N_A1_c_174_n N_A_70_101#_c_284_n 0.0138564f $X=2.68 $Y=1.2 $X2=0 $Y2=0
cc_148 N_A1_M1001_g N_A_70_101#_c_285_n 0.00590404f $X=2.64 $Y=2.595 $X2=0 $Y2=0
cc_149 N_A1_c_170_n N_A_70_101#_c_285_n 0.00486989f $X=2.68 $Y=1.035 $X2=0 $Y2=0
cc_150 N_A1_c_173_n N_A_70_101#_c_285_n 0.0148853f $X=2.68 $Y=1.2 $X2=0 $Y2=0
cc_151 N_A1_c_174_n N_A_70_101#_c_285_n 0.0481606f $X=2.68 $Y=1.2 $X2=0 $Y2=0
cc_152 N_A1_c_170_n N_VGND_c_341_n 0.00678909f $X=2.68 $Y=1.035 $X2=0 $Y2=0
cc_153 N_A1_c_170_n N_VGND_c_343_n 0.00463701f $X=2.68 $Y=1.035 $X2=0 $Y2=0
cc_154 N_A1_c_170_n N_VGND_c_344_n 0.00503886f $X=2.68 $Y=1.035 $X2=0 $Y2=0
cc_155 N_VPWR_c_200_n A_169_419# 0.010279f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_156 N_VPWR_c_200_n N_Y_M1000_d 0.00304713f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_157 N_VPWR_M1005_s N_Y_c_237_n 0.00234811f $X=0.31 $Y=2.095 $X2=0 $Y2=0
cc_158 N_VPWR_c_201_n N_Y_c_237_n 0.0174952f $X=0.455 $Y=2.475 $X2=0 $Y2=0
cc_159 N_VPWR_M1005_s N_Y_c_238_n 3.31869e-19 $X=0.31 $Y=2.095 $X2=0 $Y2=0
cc_160 N_VPWR_c_201_n N_Y_c_238_n 0.00386824f $X=0.455 $Y=2.475 $X2=0 $Y2=0
cc_161 N_VPWR_c_201_n Y 0.0261152f $X=0.455 $Y=2.475 $X2=0 $Y2=0
cc_162 N_VPWR_c_206_n Y 0.0328859f $X=2.74 $Y=3.33 $X2=0 $Y2=0
cc_163 N_VPWR_c_200_n Y 0.0202504f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VPWR_c_200_n A_381_419# 0.0262099f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_165 N_VPWR_c_202_n N_A_70_101#_c_288_n 0.0237066f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_166 A_169_419# N_Y_c_237_n 0.0048076f $X=0.845 $Y=2.095 $X2=2.905 $Y2=3.245
cc_167 N_Y_c_234_n N_A_70_101#_c_279_n 0.0255667f $X=0.84 $Y=1.185 $X2=0 $Y2=0
cc_168 N_Y_c_234_n N_A_70_101#_c_280_n 0.00420989f $X=0.84 $Y=1.185 $X2=0 $Y2=0
cc_169 N_Y_c_250_n N_A_70_101#_c_280_n 0.019558f $X=1.005 $Y=0.78 $X2=0 $Y2=0
cc_170 N_Y_c_234_n N_A_70_101#_c_283_n 0.00680274f $X=0.84 $Y=1.185 $X2=0 $Y2=0
cc_171 N_Y_c_250_n N_A_70_101#_c_283_n 0.00582789f $X=1.005 $Y=0.78 $X2=0 $Y2=0
cc_172 Y N_A_70_101#_c_289_n 0.00793068f $X=1.115 $Y=2.69 $X2=0 $Y2=0
cc_173 N_Y_c_250_n N_A_70_101#_c_286_n 0.0126136f $X=1.005 $Y=0.78 $X2=0 $Y2=0
cc_174 N_A_70_101#_c_280_n N_VGND_c_341_n 0.0141653f $X=1.35 $Y=0.35 $X2=0 $Y2=0
cc_175 N_A_70_101#_c_282_n N_VGND_c_341_n 0.031766f $X=1.515 $Y=0.715 $X2=0
+ $Y2=0
cc_176 N_A_70_101#_c_284_n N_VGND_c_341_n 0.0165754f $X=3.025 $Y=0.67 $X2=0
+ $Y2=0
cc_177 N_A_70_101#_c_280_n N_VGND_c_342_n 0.0697644f $X=1.35 $Y=0.35 $X2=0 $Y2=0
cc_178 N_A_70_101#_c_281_n N_VGND_c_342_n 0.0221876f $X=0.66 $Y=0.35 $X2=0 $Y2=0
cc_179 N_A_70_101#_c_284_n N_VGND_c_343_n 0.0153972f $X=3.025 $Y=0.67 $X2=0
+ $Y2=0
cc_180 N_A_70_101#_c_280_n N_VGND_c_344_n 0.0418368f $X=1.35 $Y=0.35 $X2=0 $Y2=0
cc_181 N_A_70_101#_c_281_n N_VGND_c_344_n 0.0127558f $X=0.66 $Y=0.35 $X2=0 $Y2=0
cc_182 N_A_70_101#_c_284_n N_VGND_c_344_n 0.0184091f $X=3.025 $Y=0.67 $X2=0
+ $Y2=0
