* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__buflp_4 A VGND VNB VPB VPWR X
X0 X a_84_21# a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VPWR A a_886_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_114_47# a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND a_84_21# a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 X a_84_21# a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 X a_84_21# a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_886_47# A a_84_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_114_367# a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_114_47# a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR a_84_21# a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 X a_84_21# a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_886_367# A a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_114_367# a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VPWR a_84_21# a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VGND a_84_21# a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_114_47# a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VGND A a_886_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_114_47# a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_114_367# a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_114_367# a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
