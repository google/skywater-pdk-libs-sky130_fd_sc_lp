* File: sky130_fd_sc_lp__nand3_4.pxi.spice
* Created: Wed Sep  2 10:04:24 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3_4%A N_A_M1006_g N_A_M1000_g N_A_M1014_g N_A_M1009_g
+ N_A_M1018_g N_A_M1016_g N_A_M1019_g N_A_M1023_g A A A N_A_c_97_n
+ PM_SKY130_FD_SC_LP__NAND3_4%A
x_PM_SKY130_FD_SC_LP__NAND3_4%B N_B_M1002_g N_B_M1004_g N_B_M1010_g N_B_M1011_g
+ N_B_M1013_g N_B_M1012_g N_B_M1020_g N_B_M1022_g N_B_c_240_p N_B_c_173_n
+ N_B_c_181_n N_B_c_182_n N_B_c_211_p N_B_c_174_n N_B_c_175_n N_B_c_191_p B B B
+ B N_B_c_176_n PM_SKY130_FD_SC_LP__NAND3_4%B
x_PM_SKY130_FD_SC_LP__NAND3_4%C N_C_M1003_g N_C_M1001_g N_C_M1005_g N_C_M1008_g
+ N_C_M1007_g N_C_M1017_g N_C_M1015_g N_C_M1021_g C C C N_C_c_299_n N_C_c_300_n
+ PM_SKY130_FD_SC_LP__NAND3_4%C
x_PM_SKY130_FD_SC_LP__NAND3_4%VPWR N_VPWR_M1000_s N_VPWR_M1009_s N_VPWR_M1023_s
+ N_VPWR_M1011_s N_VPWR_M1003_s N_VPWR_M1017_s N_VPWR_M1022_s N_VPWR_c_379_n
+ N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n
+ N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n N_VPWR_c_389_n
+ N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n VPWR N_VPWR_c_393_n
+ N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_398_n
+ N_VPWR_c_378_n PM_SKY130_FD_SC_LP__NAND3_4%VPWR
x_PM_SKY130_FD_SC_LP__NAND3_4%Y N_Y_M1006_d N_Y_M1018_d N_Y_M1000_d N_Y_M1016_d
+ N_Y_M1004_d N_Y_M1012_d N_Y_M1008_d N_Y_M1021_d N_Y_c_577_p N_Y_c_494_n
+ N_Y_c_550_n N_Y_c_487_n N_Y_c_488_n N_Y_c_503_n N_Y_c_582_p N_Y_c_489_n
+ N_Y_c_490_n N_Y_c_556_n N_Y_c_493_n N_Y_c_528_n N_Y_c_530_n N_Y_c_534_n
+ N_Y_c_535_n N_Y_c_491_n N_Y_c_536_n N_Y_c_537_n N_Y_c_538_n N_Y_c_539_n Y
+ PM_SKY130_FD_SC_LP__NAND3_4%Y
x_PM_SKY130_FD_SC_LP__NAND3_4%A_33_57# N_A_33_57#_M1006_s N_A_33_57#_M1014_s
+ N_A_33_57#_M1019_s N_A_33_57#_M1010_s N_A_33_57#_M1020_s N_A_33_57#_c_588_n
+ N_A_33_57#_c_589_n N_A_33_57#_c_590_n N_A_33_57#_c_603_n N_A_33_57#_c_591_n
+ N_A_33_57#_c_592_n N_A_33_57#_c_593_n N_A_33_57#_c_654_p N_A_33_57#_c_594_n
+ N_A_33_57#_c_595_n N_A_33_57#_c_596_n N_A_33_57#_c_597_n
+ PM_SKY130_FD_SC_LP__NAND3_4%A_33_57#
x_PM_SKY130_FD_SC_LP__NAND3_4%A_460_57# N_A_460_57#_M1002_d N_A_460_57#_M1013_d
+ N_A_460_57#_M1005_s N_A_460_57#_M1015_s N_A_460_57#_c_675_n
+ N_A_460_57#_c_672_n N_A_460_57#_c_673_n N_A_460_57#_c_674_n
+ N_A_460_57#_c_683_n N_A_460_57#_c_685_n N_A_460_57#_c_691_n
+ N_A_460_57#_c_693_n N_A_460_57#_c_686_n N_A_460_57#_c_695_n
+ PM_SKY130_FD_SC_LP__NAND3_4%A_460_57#
x_PM_SKY130_FD_SC_LP__NAND3_4%VGND N_VGND_M1001_d N_VGND_M1007_d N_VGND_c_730_n
+ N_VGND_c_731_n N_VGND_c_732_n N_VGND_c_733_n VGND N_VGND_c_734_n
+ N_VGND_c_735_n N_VGND_c_736_n N_VGND_c_737_n PM_SKY130_FD_SC_LP__NAND3_4%VGND
cc_1 VNB N_A_M1006_g 0.0303619f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.705
cc_2 VNB N_A_M1014_g 0.0209412f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.705
cc_3 VNB N_A_M1018_g 0.0209088f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.705
cc_4 VNB N_A_M1019_g 0.0221501f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.705
cc_5 VNB A 0.0142891f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_6 VNB N_A_c_97_n 0.0782539f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.51
cc_7 VNB N_B_M1002_g 0.0211114f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.705
cc_8 VNB N_B_M1010_g 0.0209962f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.705
cc_9 VNB N_B_M1013_g 0.0216173f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.705
cc_10 VNB N_B_M1020_g 0.0283972f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.705
cc_11 VNB N_B_c_173_n 0.00119566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_c_174_n 0.00179127f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.51
cc_13 VNB N_B_c_175_n 0.0354903f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.51
cc_14 VNB N_B_c_176_n 0.049162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C_M1001_g 0.0214704f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_16 VNB N_C_M1005_g 0.0206383f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.705
cc_17 VNB N_C_M1007_g 0.0206383f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.705
cc_18 VNB N_C_M1015_g 0.0209072f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.705
cc_19 VNB N_C_c_299_n 0.00326791f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=1.51
cc_20 VNB N_C_c_300_n 0.0684191f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.572
cc_21 VNB N_VPWR_c_378_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_487_n 0.0041582f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_23 VNB N_Y_c_488_n 0.00295979f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_24 VNB N_Y_c_489_n 0.00210962f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.51
cc_25 VNB N_Y_c_490_n 0.00314197f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_26 VNB N_Y_c_491_n 0.00107665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_33_57#_c_588_n 0.0305845f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.705
cc_28 VNB N_A_33_57#_c_589_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_33_57#_c_590_n 0.0094534f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=1.675
cc_30 VNB N_A_33_57#_c_591_n 0.00391652f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.705
cc_31 VNB N_A_33_57#_c_592_n 0.00329143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_33_57#_c_593_n 0.00381743f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_33 VNB N_A_33_57#_c_594_n 0.0293107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_33_57#_c_595_n 0.033073f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.51
cc_35 VNB N_A_33_57#_c_596_n 0.00203565f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.51
cc_36 VNB N_A_33_57#_c_597_n 0.00172363f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.51
cc_37 VNB N_A_460_57#_c_672_n 0.00213603f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.345
cc_38 VNB N_A_460_57#_c_673_n 0.00203727f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.705
cc_39 VNB N_A_460_57#_c_674_n 0.00225555f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.705
cc_40 VNB N_VGND_c_730_n 0.00327323f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.345
cc_41 VNB N_VGND_c_731_n 0.00144947f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.675
cc_42 VNB N_VGND_c_732_n 0.0872428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_733_n 0.00432892f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.345
cc_44 VNB N_VGND_c_734_n 0.0133858f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.705
cc_45 VNB N_VGND_c_735_n 0.0278026f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_46 VNB N_VGND_c_736_n 0.316954f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_47 VNB N_VGND_c_737_n 0.00497796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_A_M1000_g 0.0235869f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_49 VPB N_A_M1009_g 0.0179345f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_50 VPB N_A_M1016_g 0.0181927f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=2.465
cc_51 VPB N_A_M1023_g 0.0171979f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=2.465
cc_52 VPB A 0.015547f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_53 VPB N_A_c_97_n 0.0170558f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=1.51
cc_54 VPB N_B_M1004_g 0.0181468f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_55 VPB N_B_M1011_g 0.0182296f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_56 VPB N_B_M1012_g 0.0181427f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=2.465
cc_57 VPB N_B_M1022_g 0.0216056f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=2.465
cc_58 VPB N_B_c_181_n 0.00134103f $X=-0.19 $Y=1.655 $X2=0.465 $Y2=1.51
cc_59 VPB N_B_c_182_n 0.00583361f $X=-0.19 $Y=1.655 $X2=0.465 $Y2=1.51
cc_60 VPB N_B_c_174_n 0.00322055f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.51
cc_61 VPB N_B_c_175_n 0.0071052f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.51
cc_62 VPB N_B_c_176_n 0.00864527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_C_M1003_g 0.0184778f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.705
cc_64 VPB N_C_M1008_g 0.0184882f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_65 VPB N_C_M1017_g 0.0179387f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=2.465
cc_66 VPB N_C_M1021_g 0.0181284f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=2.465
cc_67 VPB N_C_c_299_n 0.0100671f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=1.51
cc_68 VPB N_C_c_300_n 0.0151719f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.572
cc_69 VPB N_VPWR_c_379_n 0.0119347f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=2.465
cc_70 VPB N_VPWR_c_380_n 0.0483636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_381_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.815 $Y2=2.465
cc_72 VPB N_VPWR_c_382_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_73 VPB N_VPWR_c_383_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.465 $Y2=1.51
cc_74 VPB N_VPWR_c_384_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.51
cc_75 VPB N_VPWR_c_385_n 0.00208088f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.51
cc_76 VPB N_VPWR_c_386_n 3.14366e-19 $X=-0.19 $Y=1.655 $X2=1.385 $Y2=1.51
cc_77 VPB N_VPWR_c_387_n 0.0103398f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=1.51
cc_78 VPB N_VPWR_c_388_n 0.0352627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_389_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.572
cc_80 VPB N_VPWR_c_390_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_391_n 0.0130339f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.572
cc_82 VPB N_VPWR_c_392_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.572
cc_83 VPB N_VPWR_c_393_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_394_n 0.014796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_395_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_396_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_397_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_398_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_378_n 0.0458496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_Y_c_490_n 0.0026594f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.51
cc_91 VPB N_Y_c_493_n 0.00464507f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.51
cc_92 N_A_M1019_g N_B_M1002_g 0.0151551f $X=1.795 $Y=0.705 $X2=0 $Y2=0
cc_93 N_A_M1023_g N_B_M1004_g 0.0200315f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_c_97_n N_B_c_176_n 0.0227024f $X=1.795 $Y=1.51 $X2=0 $Y2=0
cc_95 N_A_M1000_g N_VPWR_c_380_n 0.0203774f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A_M1009_g N_VPWR_c_380_n 7.26038e-19 $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_97 A N_VPWR_c_380_n 0.0258897f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A_c_97_n N_VPWR_c_380_n 8.28013e-19 $X=1.795 $Y=1.51 $X2=0 $Y2=0
cc_99 N_A_M1000_g N_VPWR_c_381_n 6.77662e-19 $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_M1009_g N_VPWR_c_381_n 0.0149184f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A_M1016_g N_VPWR_c_381_n 0.0149184f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_M1023_g N_VPWR_c_381_n 6.77662e-19 $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_M1016_g N_VPWR_c_382_n 7.21513e-19 $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A_M1023_g N_VPWR_c_382_n 0.0139801f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A_M1016_g N_VPWR_c_389_n 0.00486043f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_M1023_g N_VPWR_c_389_n 0.00486043f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_M1000_g N_VPWR_c_393_n 0.00486043f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_M1009_g N_VPWR_c_393_n 0.00486043f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_M1000_g N_VPWR_c_378_n 0.00824727f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A_M1009_g N_VPWR_c_378_n 0.00824727f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_M1016_g N_VPWR_c_378_n 0.00824727f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_M1023_g N_VPWR_c_378_n 0.00824727f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_113 A N_Y_c_494_n 0.0154822f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A_c_97_n N_Y_c_494_n 6.51484e-19 $X=1.795 $Y=1.51 $X2=0 $Y2=0
cc_115 N_A_M1014_g N_Y_c_487_n 0.0118617f $X=0.935 $Y=0.705 $X2=0 $Y2=0
cc_116 N_A_M1018_g N_Y_c_487_n 0.0158466f $X=1.365 $Y=0.705 $X2=0 $Y2=0
cc_117 A N_Y_c_487_n 0.0367403f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_118 N_A_c_97_n N_Y_c_487_n 0.00246131f $X=1.795 $Y=1.51 $X2=0 $Y2=0
cc_119 N_A_M1006_g N_Y_c_488_n 0.00315266f $X=0.505 $Y=0.705 $X2=0 $Y2=0
cc_120 A N_Y_c_488_n 0.0185322f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A_c_97_n N_Y_c_488_n 0.00254802f $X=1.795 $Y=1.51 $X2=0 $Y2=0
cc_122 N_A_M1009_g N_Y_c_503_n 0.0125192f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_M1016_g N_Y_c_503_n 0.0171019f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_124 A N_Y_c_503_n 0.0305479f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A_c_97_n N_Y_c_503_n 5.79315e-19 $X=1.795 $Y=1.51 $X2=0 $Y2=0
cc_126 N_A_M1018_g N_Y_c_489_n 0.00297011f $X=1.365 $Y=0.705 $X2=0 $Y2=0
cc_127 N_A_M1019_g N_Y_c_489_n 0.00260622f $X=1.795 $Y=0.705 $X2=0 $Y2=0
cc_128 A N_Y_c_489_n 0.00206445f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A_c_97_n N_Y_c_489_n 0.0080396f $X=1.795 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A_M1016_g N_Y_c_490_n 0.00356303f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A_M1023_g N_Y_c_490_n 0.0150689f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_132 A N_Y_c_490_n 0.0253263f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A_c_97_n N_Y_c_490_n 0.0252603f $X=1.795 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A_M1019_g N_Y_c_491_n 0.00120657f $X=1.795 $Y=0.705 $X2=0 $Y2=0
cc_135 N_A_M1006_g N_A_33_57#_c_588_n 0.00371035f $X=0.505 $Y=0.705 $X2=0 $Y2=0
cc_136 A N_A_33_57#_c_588_n 0.0196911f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A_c_97_n N_A_33_57#_c_588_n 0.00293822f $X=1.795 $Y=1.51 $X2=0 $Y2=0
cc_138 N_A_M1006_g N_A_33_57#_c_589_n 0.0126328f $X=0.505 $Y=0.705 $X2=0 $Y2=0
cc_139 N_A_M1014_g N_A_33_57#_c_589_n 0.00835698f $X=0.935 $Y=0.705 $X2=0 $Y2=0
cc_140 N_A_M1006_g N_A_33_57#_c_603_n 5.231e-19 $X=0.505 $Y=0.705 $X2=0 $Y2=0
cc_141 N_A_M1014_g N_A_33_57#_c_603_n 0.00629337f $X=0.935 $Y=0.705 $X2=0 $Y2=0
cc_142 N_A_M1018_g N_A_33_57#_c_603_n 0.00624891f $X=1.365 $Y=0.705 $X2=0 $Y2=0
cc_143 N_A_M1019_g N_A_33_57#_c_603_n 5.24123e-19 $X=1.795 $Y=0.705 $X2=0 $Y2=0
cc_144 N_A_M1018_g N_A_33_57#_c_591_n 0.00831042f $X=1.365 $Y=0.705 $X2=0 $Y2=0
cc_145 N_A_M1019_g N_A_33_57#_c_591_n 0.0123266f $X=1.795 $Y=0.705 $X2=0 $Y2=0
cc_146 N_A_M1019_g N_A_33_57#_c_593_n 0.00114873f $X=1.795 $Y=0.705 $X2=0 $Y2=0
cc_147 N_A_M1014_g N_A_33_57#_c_596_n 9.09899e-19 $X=0.935 $Y=0.705 $X2=0 $Y2=0
cc_148 N_A_M1018_g N_A_33_57#_c_596_n 9.09899e-19 $X=1.365 $Y=0.705 $X2=0 $Y2=0
cc_149 N_A_M1006_g N_VGND_c_732_n 0.00325902f $X=0.505 $Y=0.705 $X2=0 $Y2=0
cc_150 N_A_M1014_g N_VGND_c_732_n 0.00325872f $X=0.935 $Y=0.705 $X2=0 $Y2=0
cc_151 N_A_M1018_g N_VGND_c_732_n 0.00325872f $X=1.365 $Y=0.705 $X2=0 $Y2=0
cc_152 N_A_M1019_g N_VGND_c_732_n 0.00325902f $X=1.795 $Y=0.705 $X2=0 $Y2=0
cc_153 N_A_M1006_g N_VGND_c_736_n 0.00553347f $X=0.505 $Y=0.705 $X2=0 $Y2=0
cc_154 N_A_M1014_g N_VGND_c_736_n 0.00486898f $X=0.935 $Y=0.705 $X2=0 $Y2=0
cc_155 N_A_M1018_g N_VGND_c_736_n 0.00486898f $X=1.365 $Y=0.705 $X2=0 $Y2=0
cc_156 N_A_M1019_g N_VGND_c_736_n 0.00488654f $X=1.795 $Y=0.705 $X2=0 $Y2=0
cc_157 N_B_M1012_g N_C_M1003_g 0.035511f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B_c_181_n N_C_M1003_g 0.00114957f $X=2.987 $Y=1.92 $X2=0 $Y2=0
cc_159 N_B_c_191_p N_C_M1003_g 0.0118166f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_160 N_B_M1013_g N_C_M1001_g 0.0197813f $X=3.105 $Y=0.705 $X2=0 $Y2=0
cc_161 N_B_c_191_p N_C_M1008_g 0.0118715f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_162 N_B_c_191_p N_C_M1017_g 0.0116622f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_163 N_B_M1020_g N_C_M1015_g 0.029161f $X=5.285 $Y=0.705 $X2=0 $Y2=0
cc_164 N_B_M1022_g N_C_M1021_g 0.029161f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_165 N_B_c_182_n N_C_M1021_g 0.00251031f $X=5.315 $Y=1.92 $X2=0 $Y2=0
cc_166 N_B_c_191_p N_C_M1021_g 0.0116073f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_167 N_B_M1012_g N_C_c_299_n 4.79398e-19 $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_168 N_B_c_173_n N_C_c_299_n 0.012772f $X=2.987 $Y=1.605 $X2=0 $Y2=0
cc_169 N_B_c_181_n N_C_c_299_n 0.0100853f $X=2.987 $Y=1.92 $X2=0 $Y2=0
cc_170 N_B_c_174_n N_C_c_299_n 0.0190624f $X=5.375 $Y=1.51 $X2=0 $Y2=0
cc_171 N_B_c_175_n N_C_c_299_n 4.07599e-19 $X=5.375 $Y=1.51 $X2=0 $Y2=0
cc_172 N_B_c_191_p N_C_c_299_n 0.102488f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_173 N_B_c_176_n N_C_c_299_n 5.0426e-19 $X=3.105 $Y=1.51 $X2=0 $Y2=0
cc_174 N_B_c_173_n N_C_c_300_n 2.22064e-19 $X=2.987 $Y=1.605 $X2=0 $Y2=0
cc_175 N_B_c_174_n N_C_c_300_n 6.18792e-19 $X=5.375 $Y=1.51 $X2=0 $Y2=0
cc_176 N_B_c_175_n N_C_c_300_n 0.029161f $X=5.375 $Y=1.51 $X2=0 $Y2=0
cc_177 N_B_c_191_p N_C_c_300_n 0.00222779f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_178 N_B_c_176_n N_C_c_300_n 0.02316f $X=3.105 $Y=1.51 $X2=0 $Y2=0
cc_179 N_B_c_211_p N_VPWR_M1011_s 0.00229733f $X=3.18 $Y=2.02 $X2=0 $Y2=0
cc_180 N_B_c_191_p N_VPWR_M1003_s 0.00393014f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_181 N_B_c_191_p N_VPWR_M1017_s 0.00334942f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_182 N_B_c_182_n N_VPWR_M1022_s 0.00332446f $X=5.315 $Y=1.92 $X2=0 $Y2=0
cc_183 N_B_c_191_p N_VPWR_M1022_s 0.00915499f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_184 N_B_M1004_g N_VPWR_c_382_n 0.0139613f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_185 N_B_M1011_g N_VPWR_c_382_n 7.59846e-19 $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B_M1004_g N_VPWR_c_383_n 5.82718e-19 $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_187 N_B_M1011_g N_VPWR_c_383_n 0.0106726f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_188 N_B_M1012_g N_VPWR_c_383_n 0.0105703f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_189 N_B_M1012_g N_VPWR_c_384_n 0.00486043f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_190 N_B_M1012_g N_VPWR_c_385_n 5.75816e-19 $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B_M1022_g N_VPWR_c_386_n 5.75816e-19 $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_192 N_B_M1022_g N_VPWR_c_388_n 0.0170434f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_193 N_B_c_174_n N_VPWR_c_388_n 0.00382425f $X=5.375 $Y=1.51 $X2=0 $Y2=0
cc_194 N_B_c_175_n N_VPWR_c_388_n 8.11454e-19 $X=5.375 $Y=1.51 $X2=0 $Y2=0
cc_195 N_B_c_191_p N_VPWR_c_388_n 0.00312145f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_196 N_B_M1004_g N_VPWR_c_391_n 0.00486043f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_197 N_B_M1011_g N_VPWR_c_391_n 0.00486043f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_198 N_B_M1022_g N_VPWR_c_395_n 0.00486043f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_199 N_B_M1004_g N_VPWR_c_378_n 0.00824727f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_200 N_B_M1011_g N_VPWR_c_378_n 0.00824727f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_201 N_B_M1012_g N_VPWR_c_378_n 0.0082726f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B_M1022_g N_VPWR_c_378_n 0.0082726f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B_c_191_p N_Y_M1012_d 0.0051211f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_204 N_B_c_191_p N_Y_M1008_d 0.00334509f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_205 N_B_c_191_p N_Y_M1021_d 0.00528357f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_206 N_B_c_176_n N_Y_c_489_n 4.35391e-19 $X=3.105 $Y=1.51 $X2=0 $Y2=0
cc_207 N_B_M1004_g N_Y_c_490_n 0.00256252f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B_c_240_p N_Y_c_490_n 0.0155044f $X=2.795 $Y=1.515 $X2=0 $Y2=0
cc_209 N_B_c_176_n N_Y_c_490_n 0.00335598f $X=3.105 $Y=1.51 $X2=0 $Y2=0
cc_210 N_B_M1004_g N_Y_c_493_n 0.0129249f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_211 N_B_M1011_g N_Y_c_493_n 0.00279785f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_212 N_B_c_240_p N_Y_c_493_n 0.0343563f $X=2.795 $Y=1.515 $X2=0 $Y2=0
cc_213 N_B_c_181_n N_Y_c_493_n 0.00863112f $X=2.987 $Y=1.92 $X2=0 $Y2=0
cc_214 N_B_c_176_n N_Y_c_493_n 0.00327622f $X=3.105 $Y=1.51 $X2=0 $Y2=0
cc_215 N_B_M1011_g N_Y_c_528_n 0.00556109f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_216 N_B_M1012_g N_Y_c_528_n 9.57732e-19 $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_217 N_B_M1011_g N_Y_c_530_n 0.0142032f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B_M1012_g N_Y_c_530_n 0.0122068f $X=3.105 $Y=2.465 $X2=0 $Y2=0
cc_219 N_B_c_211_p N_Y_c_530_n 0.0249007f $X=3.18 $Y=2.02 $X2=0 $Y2=0
cc_220 N_B_c_176_n N_Y_c_530_n 2.86047e-19 $X=3.105 $Y=1.51 $X2=0 $Y2=0
cc_221 N_B_c_191_p N_Y_c_534_n 0.0349355f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_222 N_B_c_191_p N_Y_c_535_n 0.0327296f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_223 N_B_M1011_g N_Y_c_536_n 0.0016312f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_224 N_B_c_191_p N_Y_c_537_n 0.0136549f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_225 N_B_c_191_p N_Y_c_538_n 0.0136549f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_226 N_B_c_191_p N_Y_c_539_n 0.0136549f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_227 N_B_M1002_g N_A_33_57#_c_591_n 2.42902e-19 $X=2.225 $Y=0.705 $X2=0 $Y2=0
cc_228 N_B_M1002_g N_A_33_57#_c_592_n 0.0137234f $X=2.225 $Y=0.705 $X2=0 $Y2=0
cc_229 N_B_M1010_g N_A_33_57#_c_592_n 0.0124229f $X=2.655 $Y=0.705 $X2=0 $Y2=0
cc_230 N_B_c_240_p N_A_33_57#_c_592_n 0.0423704f $X=2.795 $Y=1.515 $X2=0 $Y2=0
cc_231 N_B_c_176_n N_A_33_57#_c_592_n 0.00255068f $X=3.105 $Y=1.51 $X2=0 $Y2=0
cc_232 N_B_M1013_g N_A_33_57#_c_594_n 0.0129017f $X=3.105 $Y=0.705 $X2=0 $Y2=0
cc_233 N_B_M1020_g N_A_33_57#_c_594_n 0.014789f $X=5.285 $Y=0.705 $X2=0 $Y2=0
cc_234 N_B_c_173_n N_A_33_57#_c_594_n 0.0134113f $X=2.987 $Y=1.605 $X2=0 $Y2=0
cc_235 N_B_c_174_n N_A_33_57#_c_594_n 0.0271395f $X=5.375 $Y=1.51 $X2=0 $Y2=0
cc_236 N_B_c_175_n N_A_33_57#_c_594_n 0.00459237f $X=5.375 $Y=1.51 $X2=0 $Y2=0
cc_237 N_B_c_191_p N_A_33_57#_c_594_n 0.0112237f $X=5.2 $Y=2.02 $X2=0 $Y2=0
cc_238 N_B_M1020_g N_A_33_57#_c_595_n 0.00365969f $X=5.285 $Y=0.705 $X2=0 $Y2=0
cc_239 N_B_c_240_p N_A_33_57#_c_597_n 0.00157138f $X=2.795 $Y=1.515 $X2=0 $Y2=0
cc_240 N_B_c_173_n N_A_33_57#_c_597_n 0.0185941f $X=2.987 $Y=1.605 $X2=0 $Y2=0
cc_241 N_B_c_176_n N_A_33_57#_c_597_n 0.00314894f $X=3.105 $Y=1.51 $X2=0 $Y2=0
cc_242 N_B_M1002_g N_A_460_57#_c_675_n 0.0053946f $X=2.225 $Y=0.705 $X2=0 $Y2=0
cc_243 N_B_M1010_g N_A_460_57#_c_675_n 0.00717622f $X=2.655 $Y=0.705 $X2=0 $Y2=0
cc_244 N_B_M1013_g N_A_460_57#_c_675_n 6.67552e-19 $X=3.105 $Y=0.705 $X2=0 $Y2=0
cc_245 N_B_M1010_g N_A_460_57#_c_672_n 0.00856015f $X=2.655 $Y=0.705 $X2=0 $Y2=0
cc_246 N_B_M1013_g N_A_460_57#_c_672_n 0.00959783f $X=3.105 $Y=0.705 $X2=0 $Y2=0
cc_247 N_B_M1002_g N_A_460_57#_c_673_n 0.00223164f $X=2.225 $Y=0.705 $X2=0 $Y2=0
cc_248 N_B_M1010_g N_A_460_57#_c_673_n 9.09899e-19 $X=2.655 $Y=0.705 $X2=0 $Y2=0
cc_249 N_B_M1013_g N_A_460_57#_c_674_n 4.71487e-19 $X=3.105 $Y=0.705 $X2=0 $Y2=0
cc_250 N_B_M1010_g N_A_460_57#_c_683_n 5.97429e-19 $X=2.655 $Y=0.705 $X2=0 $Y2=0
cc_251 N_B_M1013_g N_A_460_57#_c_683_n 0.00480975f $X=3.105 $Y=0.705 $X2=0 $Y2=0
cc_252 N_B_M1013_g N_A_460_57#_c_685_n 0.00149689f $X=3.105 $Y=0.705 $X2=0 $Y2=0
cc_253 N_B_M1020_g N_A_460_57#_c_686_n 0.00319371f $X=5.285 $Y=0.705 $X2=0 $Y2=0
cc_254 N_B_M1020_g N_VGND_c_731_n 0.00173041f $X=5.285 $Y=0.705 $X2=0 $Y2=0
cc_255 N_B_M1002_g N_VGND_c_732_n 0.0050097f $X=2.225 $Y=0.705 $X2=0 $Y2=0
cc_256 N_B_M1010_g N_VGND_c_732_n 0.00325872f $X=2.655 $Y=0.705 $X2=0 $Y2=0
cc_257 N_B_M1013_g N_VGND_c_732_n 0.00325896f $X=3.105 $Y=0.705 $X2=0 $Y2=0
cc_258 N_B_M1020_g N_VGND_c_735_n 0.00512259f $X=5.285 $Y=0.705 $X2=0 $Y2=0
cc_259 N_B_M1002_g N_VGND_c_736_n 0.00951894f $X=2.225 $Y=0.705 $X2=0 $Y2=0
cc_260 N_B_M1010_g N_VGND_c_736_n 0.00490447f $X=2.655 $Y=0.705 $X2=0 $Y2=0
cc_261 N_B_M1013_g N_VGND_c_736_n 0.00497112f $X=3.105 $Y=0.705 $X2=0 $Y2=0
cc_262 N_B_M1020_g N_VGND_c_736_n 0.0102916f $X=5.285 $Y=0.705 $X2=0 $Y2=0
cc_263 N_C_M1003_g N_VPWR_c_383_n 5.75816e-19 $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_264 N_C_M1003_g N_VPWR_c_384_n 0.00486043f $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_265 N_C_M1003_g N_VPWR_c_385_n 0.0103526f $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_266 N_C_M1008_g N_VPWR_c_385_n 0.00241634f $X=3.995 $Y=2.465 $X2=0 $Y2=0
cc_267 N_C_M1008_g N_VPWR_c_386_n 5.88023e-19 $X=3.995 $Y=2.465 $X2=0 $Y2=0
cc_268 N_C_M1017_g N_VPWR_c_386_n 0.0106396f $X=4.425 $Y=2.465 $X2=0 $Y2=0
cc_269 N_C_M1021_g N_VPWR_c_386_n 0.0105703f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_270 N_C_M1021_g N_VPWR_c_388_n 6.24191e-19 $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_271 N_C_M1008_g N_VPWR_c_394_n 0.00585385f $X=3.995 $Y=2.465 $X2=0 $Y2=0
cc_272 N_C_M1017_g N_VPWR_c_394_n 0.00486043f $X=4.425 $Y=2.465 $X2=0 $Y2=0
cc_273 N_C_M1021_g N_VPWR_c_395_n 0.00486043f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_274 N_C_M1003_g N_VPWR_c_378_n 0.0082726f $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_275 N_C_M1008_g N_VPWR_c_378_n 0.0106981f $X=3.995 $Y=2.465 $X2=0 $Y2=0
cc_276 N_C_M1017_g N_VPWR_c_378_n 0.00824727f $X=4.425 $Y=2.465 $X2=0 $Y2=0
cc_277 N_C_M1021_g N_VPWR_c_378_n 0.0082726f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_278 N_C_M1003_g N_Y_c_534_n 0.0124371f $X=3.535 $Y=2.465 $X2=0 $Y2=0
cc_279 N_C_M1008_g N_Y_c_534_n 0.0131711f $X=3.995 $Y=2.465 $X2=0 $Y2=0
cc_280 N_C_M1017_g N_Y_c_535_n 0.0122129f $X=4.425 $Y=2.465 $X2=0 $Y2=0
cc_281 N_C_M1021_g N_Y_c_535_n 0.0122595f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_282 N_C_M1001_g N_A_33_57#_c_594_n 0.0106164f $X=3.565 $Y=0.705 $X2=0 $Y2=0
cc_283 N_C_M1005_g N_A_33_57#_c_594_n 0.0104926f $X=3.995 $Y=0.705 $X2=0 $Y2=0
cc_284 N_C_M1007_g N_A_33_57#_c_594_n 0.0104926f $X=4.425 $Y=0.705 $X2=0 $Y2=0
cc_285 N_C_M1015_g N_A_33_57#_c_594_n 0.010446f $X=4.855 $Y=0.705 $X2=0 $Y2=0
cc_286 N_C_c_299_n N_A_33_57#_c_594_n 0.113366f $X=4.575 $Y=1.51 $X2=0 $Y2=0
cc_287 N_C_c_300_n N_A_33_57#_c_594_n 0.00998783f $X=4.855 $Y=1.51 $X2=0 $Y2=0
cc_288 N_C_M1001_g N_A_460_57#_c_674_n 0.00208971f $X=3.565 $Y=0.705 $X2=0 $Y2=0
cc_289 N_C_M1001_g N_A_460_57#_c_683_n 0.00460791f $X=3.565 $Y=0.705 $X2=0 $Y2=0
cc_290 N_C_M1005_g N_A_460_57#_c_683_n 6.67119e-19 $X=3.995 $Y=0.705 $X2=0 $Y2=0
cc_291 N_C_M1001_g N_A_460_57#_c_685_n 4.26794e-19 $X=3.565 $Y=0.705 $X2=0 $Y2=0
cc_292 N_C_M1001_g N_A_460_57#_c_691_n 0.00938051f $X=3.565 $Y=0.705 $X2=0 $Y2=0
cc_293 N_C_M1005_g N_A_460_57#_c_691_n 0.00961846f $X=3.995 $Y=0.705 $X2=0 $Y2=0
cc_294 N_C_M1005_g N_A_460_57#_c_693_n 7.95083e-19 $X=3.995 $Y=0.705 $X2=0 $Y2=0
cc_295 N_C_M1007_g N_A_460_57#_c_693_n 8.04766e-19 $X=4.425 $Y=0.705 $X2=0 $Y2=0
cc_296 N_C_M1007_g N_A_460_57#_c_695_n 0.00961846f $X=4.425 $Y=0.705 $X2=0 $Y2=0
cc_297 N_C_M1015_g N_A_460_57#_c_695_n 0.00989361f $X=4.855 $Y=0.705 $X2=0 $Y2=0
cc_298 N_C_M1001_g N_VGND_c_730_n 0.00248612f $X=3.565 $Y=0.705 $X2=0 $Y2=0
cc_299 N_C_M1005_g N_VGND_c_730_n 0.00894883f $X=3.995 $Y=0.705 $X2=0 $Y2=0
cc_300 N_C_M1007_g N_VGND_c_730_n 0.00126341f $X=4.425 $Y=0.705 $X2=0 $Y2=0
cc_301 N_C_M1005_g N_VGND_c_731_n 0.00126504f $X=3.995 $Y=0.705 $X2=0 $Y2=0
cc_302 N_C_M1007_g N_VGND_c_731_n 0.00927215f $X=4.425 $Y=0.705 $X2=0 $Y2=0
cc_303 N_C_M1015_g N_VGND_c_731_n 0.0103911f $X=4.855 $Y=0.705 $X2=0 $Y2=0
cc_304 N_C_M1001_g N_VGND_c_732_n 0.00391619f $X=3.565 $Y=0.705 $X2=0 $Y2=0
cc_305 N_C_M1005_g N_VGND_c_734_n 0.00331555f $X=3.995 $Y=0.705 $X2=0 $Y2=0
cc_306 N_C_M1007_g N_VGND_c_734_n 0.00331555f $X=4.425 $Y=0.705 $X2=0 $Y2=0
cc_307 N_C_M1015_g N_VGND_c_735_n 0.00331737f $X=4.855 $Y=0.705 $X2=0 $Y2=0
cc_308 N_C_M1001_g N_VGND_c_736_n 0.00554734f $X=3.565 $Y=0.705 $X2=0 $Y2=0
cc_309 N_C_M1005_g N_VGND_c_736_n 0.00415929f $X=3.995 $Y=0.705 $X2=0 $Y2=0
cc_310 N_C_M1007_g N_VGND_c_736_n 0.00415929f $X=4.425 $Y=0.705 $X2=0 $Y2=0
cc_311 N_C_M1015_g N_VGND_c_736_n 0.00418057f $X=4.855 $Y=0.705 $X2=0 $Y2=0
cc_312 N_VPWR_c_378_n N_Y_M1000_d 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_313 N_VPWR_c_378_n N_Y_M1016_d 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_314 N_VPWR_c_378_n N_Y_M1004_d 0.00571434f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_315 N_VPWR_c_378_n N_Y_M1012_d 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_316 N_VPWR_c_378_n N_Y_M1008_d 0.00501859f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_317 N_VPWR_c_378_n N_Y_M1021_d 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_318 N_VPWR_c_393_n N_Y_c_550_n 0.0124525f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_319 N_VPWR_c_378_n N_Y_c_550_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_M1009_s N_Y_c_503_n 0.00333424f $X=1.03 $Y=1.835 $X2=0 $Y2=0
cc_321 N_VPWR_c_381_n N_Y_c_503_n 0.0171443f $X=1.17 $Y=2.355 $X2=0 $Y2=0
cc_322 N_VPWR_M1023_s N_Y_c_490_n 5.81731e-19 $X=1.89 $Y=1.835 $X2=0 $Y2=0
cc_323 N_VPWR_c_382_n N_Y_c_490_n 0.00663404f $X=2.03 $Y=2.2 $X2=0 $Y2=0
cc_324 N_VPWR_c_389_n N_Y_c_556_n 0.0124525f $X=1.865 $Y=3.33 $X2=0 $Y2=0
cc_325 N_VPWR_c_378_n N_Y_c_556_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_326 N_VPWR_M1023_s N_Y_c_493_n 0.00119058f $X=1.89 $Y=1.835 $X2=0 $Y2=0
cc_327 N_VPWR_c_382_n N_Y_c_493_n 0.0109431f $X=2.03 $Y=2.2 $X2=0 $Y2=0
cc_328 N_VPWR_M1011_s N_Y_c_530_n 0.00344196f $X=2.75 $Y=1.835 $X2=0 $Y2=0
cc_329 N_VPWR_c_383_n N_Y_c_530_n 0.0170777f $X=2.89 $Y=2.755 $X2=0 $Y2=0
cc_330 N_VPWR_M1003_s N_Y_c_534_n 0.00405824f $X=3.61 $Y=1.835 $X2=0 $Y2=0
cc_331 N_VPWR_c_385_n N_Y_c_534_n 0.0177324f $X=3.75 $Y=2.755 $X2=0 $Y2=0
cc_332 N_VPWR_M1017_s N_Y_c_535_n 0.00344593f $X=4.5 $Y=1.835 $X2=0 $Y2=0
cc_333 N_VPWR_c_386_n N_Y_c_535_n 0.0170777f $X=4.64 $Y=2.755 $X2=0 $Y2=0
cc_334 N_VPWR_c_391_n N_Y_c_536_n 0.0120977f $X=2.725 $Y=3.33 $X2=0 $Y2=0
cc_335 N_VPWR_c_378_n N_Y_c_536_n 0.00691495f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_336 N_VPWR_c_384_n N_Y_c_537_n 0.0124525f $X=3.585 $Y=3.33 $X2=0 $Y2=0
cc_337 N_VPWR_c_378_n N_Y_c_537_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_338 N_VPWR_c_394_n N_Y_c_538_n 0.0128073f $X=4.475 $Y=3.33 $X2=0 $Y2=0
cc_339 N_VPWR_c_378_n N_Y_c_538_n 0.00769778f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_340 N_VPWR_c_395_n N_Y_c_539_n 0.0124525f $X=5.335 $Y=3.33 $X2=0 $Y2=0
cc_341 N_VPWR_c_378_n N_Y_c_539_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_342 N_Y_c_487_n N_A_33_57#_M1014_s 0.00176461f $X=1.485 $Y=1.14 $X2=0 $Y2=0
cc_343 N_Y_c_488_n N_A_33_57#_c_588_n 0.00166817f $X=0.815 $Y=1.14 $X2=0 $Y2=0
cc_344 N_Y_M1006_d N_A_33_57#_c_589_n 0.00176461f $X=0.58 $Y=0.285 $X2=0 $Y2=0
cc_345 N_Y_c_577_p N_A_33_57#_c_589_n 0.0125606f $X=0.72 $Y=0.76 $X2=0 $Y2=0
cc_346 N_Y_c_487_n N_A_33_57#_c_589_n 0.00284209f $X=1.485 $Y=1.14 $X2=0 $Y2=0
cc_347 N_Y_c_487_n N_A_33_57#_c_603_n 0.0169714f $X=1.485 $Y=1.14 $X2=0 $Y2=0
cc_348 N_Y_M1018_d N_A_33_57#_c_591_n 0.00176461f $X=1.44 $Y=0.285 $X2=0 $Y2=0
cc_349 N_Y_c_487_n N_A_33_57#_c_591_n 0.00284209f $X=1.485 $Y=1.14 $X2=0 $Y2=0
cc_350 N_Y_c_582_p N_A_33_57#_c_591_n 0.0126348f $X=1.58 $Y=0.76 $X2=0 $Y2=0
cc_351 N_Y_c_493_n N_A_33_57#_c_592_n 0.00216048f $X=2.365 $Y=1.86 $X2=0 $Y2=0
cc_352 N_Y_c_489_n N_A_33_57#_c_593_n 0.00253398f $X=1.602 $Y=1.425 $X2=0 $Y2=0
cc_353 N_Y_c_490_n N_A_33_57#_c_593_n 0.0110214f $X=1.6 $Y=2.1 $X2=0 $Y2=0
cc_354 N_Y_c_493_n N_A_33_57#_c_593_n 0.00406057f $X=2.365 $Y=1.86 $X2=0 $Y2=0
cc_355 N_Y_c_491_n N_A_33_57#_c_593_n 0.00926935f $X=1.597 $Y=1.14 $X2=0 $Y2=0
cc_356 N_A_33_57#_c_592_n N_A_460_57#_M1002_d 0.00176461f $X=2.775 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_357 N_A_33_57#_c_594_n N_A_460_57#_M1013_d 0.00208352f $X=5.405 $Y=1.17 $X2=0
+ $Y2=0
cc_358 N_A_33_57#_c_594_n N_A_460_57#_M1005_s 0.00176891f $X=5.405 $Y=1.17 $X2=0
+ $Y2=0
cc_359 N_A_33_57#_c_594_n N_A_460_57#_M1015_s 0.00176891f $X=5.405 $Y=1.17 $X2=0
+ $Y2=0
cc_360 N_A_33_57#_c_592_n N_A_460_57#_c_675_n 0.017036f $X=2.775 $Y=1.17 $X2=0
+ $Y2=0
cc_361 N_A_33_57#_M1010_s N_A_460_57#_c_672_n 0.00221305f $X=2.73 $Y=0.285 $X2=0
+ $Y2=0
cc_362 N_A_33_57#_c_592_n N_A_460_57#_c_672_n 0.00272017f $X=2.775 $Y=1.17 $X2=0
+ $Y2=0
cc_363 N_A_33_57#_c_654_p N_A_460_57#_c_672_n 0.011248f $X=2.89 $Y=0.81 $X2=0
+ $Y2=0
cc_364 N_A_33_57#_c_594_n N_A_460_57#_c_672_n 0.00315715f $X=5.405 $Y=1.17 $X2=0
+ $Y2=0
cc_365 N_A_33_57#_c_591_n N_A_460_57#_c_673_n 0.00855299f $X=1.88 $Y=0.34 $X2=0
+ $Y2=0
cc_366 N_A_33_57#_c_594_n N_A_460_57#_c_685_n 0.0173432f $X=5.405 $Y=1.17 $X2=0
+ $Y2=0
cc_367 N_A_33_57#_c_594_n N_A_460_57#_c_691_n 0.0898091f $X=5.405 $Y=1.17 $X2=0
+ $Y2=0
cc_368 N_A_33_57#_c_594_n N_VGND_M1001_d 0.00176891f $X=5.405 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_369 N_A_33_57#_c_594_n N_VGND_M1007_d 0.00176891f $X=5.405 $Y=1.17 $X2=0
+ $Y2=0
cc_370 N_A_33_57#_c_595_n N_VGND_c_731_n 0.00440788f $X=5.5 $Y=0.43 $X2=0 $Y2=0
cc_371 N_A_33_57#_c_589_n N_VGND_c_732_n 0.0352183f $X=0.985 $Y=0.34 $X2=0 $Y2=0
cc_372 N_A_33_57#_c_590_n N_VGND_c_732_n 0.021506f $X=0.425 $Y=0.34 $X2=0 $Y2=0
cc_373 N_A_33_57#_c_591_n N_VGND_c_732_n 0.05167f $X=1.88 $Y=0.34 $X2=0 $Y2=0
cc_374 N_A_33_57#_c_596_n N_VGND_c_732_n 0.023347f $X=1.15 $Y=0.34 $X2=0 $Y2=0
cc_375 N_A_33_57#_c_595_n N_VGND_c_735_n 0.0173955f $X=5.5 $Y=0.43 $X2=0 $Y2=0
cc_376 N_A_33_57#_c_589_n N_VGND_c_736_n 0.0197959f $X=0.985 $Y=0.34 $X2=0 $Y2=0
cc_377 N_A_33_57#_c_590_n N_VGND_c_736_n 0.0116633f $X=0.425 $Y=0.34 $X2=0 $Y2=0
cc_378 N_A_33_57#_c_591_n N_VGND_c_736_n 0.0287313f $X=1.88 $Y=0.34 $X2=0 $Y2=0
cc_379 N_A_33_57#_c_595_n N_VGND_c_736_n 0.00998284f $X=5.5 $Y=0.43 $X2=0 $Y2=0
cc_380 N_A_33_57#_c_596_n N_VGND_c_736_n 0.0125753f $X=1.15 $Y=0.34 $X2=0 $Y2=0
cc_381 N_A_460_57#_c_691_n N_VGND_M1001_d 0.00335318f $X=4.065 $Y=0.807
+ $X2=-0.19 $Y2=-0.245
cc_382 N_A_460_57#_c_695_n N_VGND_M1007_d 0.00335318f $X=4.93 $Y=0.807 $X2=0
+ $Y2=0
cc_383 N_A_460_57#_c_674_n N_VGND_c_730_n 0.00833645f $X=3.34 $Y=0.425 $X2=0
+ $Y2=0
cc_384 N_A_460_57#_c_691_n N_VGND_c_730_n 0.0147753f $X=4.065 $Y=0.807 $X2=0
+ $Y2=0
cc_385 N_A_460_57#_c_695_n N_VGND_c_731_n 0.0165001f $X=4.93 $Y=0.807 $X2=0
+ $Y2=0
cc_386 N_A_460_57#_c_672_n N_VGND_c_732_n 0.03588f $X=3.175 $Y=0.34 $X2=0 $Y2=0
cc_387 N_A_460_57#_c_673_n N_VGND_c_732_n 0.0234284f $X=2.605 $Y=0.34 $X2=0
+ $Y2=0
cc_388 N_A_460_57#_c_674_n N_VGND_c_732_n 0.0235331f $X=3.34 $Y=0.425 $X2=0
+ $Y2=0
cc_389 N_A_460_57#_c_691_n N_VGND_c_732_n 0.00197392f $X=4.065 $Y=0.807 $X2=0
+ $Y2=0
cc_390 N_A_460_57#_c_691_n N_VGND_c_734_n 0.00152385f $X=4.065 $Y=0.807 $X2=0
+ $Y2=0
cc_391 N_A_460_57#_c_693_n N_VGND_c_734_n 0.00363847f $X=4.355 $Y=0.807 $X2=0
+ $Y2=0
cc_392 N_A_460_57#_c_695_n N_VGND_c_734_n 0.00152385f $X=4.93 $Y=0.807 $X2=0
+ $Y2=0
cc_393 N_A_460_57#_c_686_n N_VGND_c_735_n 0.00385932f $X=5.07 $Y=0.83 $X2=0
+ $Y2=0
cc_394 N_A_460_57#_c_695_n N_VGND_c_735_n 0.00158787f $X=4.93 $Y=0.807 $X2=0
+ $Y2=0
cc_395 N_A_460_57#_c_672_n N_VGND_c_736_n 0.0201952f $X=3.175 $Y=0.34 $X2=0
+ $Y2=0
cc_396 N_A_460_57#_c_673_n N_VGND_c_736_n 0.0125908f $X=2.605 $Y=0.34 $X2=0
+ $Y2=0
cc_397 N_A_460_57#_c_674_n N_VGND_c_736_n 0.012728f $X=3.34 $Y=0.425 $X2=0 $Y2=0
cc_398 N_A_460_57#_c_691_n N_VGND_c_736_n 0.00738139f $X=4.065 $Y=0.807 $X2=0
+ $Y2=0
cc_399 N_A_460_57#_c_693_n N_VGND_c_736_n 0.00788332f $X=4.355 $Y=0.807 $X2=0
+ $Y2=0
cc_400 N_A_460_57#_c_686_n N_VGND_c_736_n 0.00822401f $X=5.07 $Y=0.83 $X2=0
+ $Y2=0
cc_401 N_A_460_57#_c_695_n N_VGND_c_736_n 0.00645782f $X=4.93 $Y=0.807 $X2=0
+ $Y2=0
