* File: sky130_fd_sc_lp__buflp_1.pxi.spice
* Created: Wed Sep  2 09:36:27 2020
* 
x_PM_SKY130_FD_SC_LP__BUFLP_1%A_86_21# N_A_86_21#_M1004_d N_A_86_21#_M1001_d
+ N_A_86_21#_M1003_g N_A_86_21#_M1002_g N_A_86_21#_c_38_n N_A_86_21#_M1000_g
+ N_A_86_21#_M1005_g N_A_86_21#_c_40_n N_A_86_21#_c_41_n N_A_86_21#_c_42_n
+ N_A_86_21#_c_50_p N_A_86_21#_c_70_p N_A_86_21#_c_43_n N_A_86_21#_c_44_n
+ N_A_86_21#_c_45_n PM_SKY130_FD_SC_LP__BUFLP_1%A_86_21#
x_PM_SKY130_FD_SC_LP__BUFLP_1%A N_A_c_100_n N_A_M1006_g N_A_M1007_g N_A_c_102_n
+ N_A_M1004_g N_A_M1001_g A A A A N_A_c_104_n N_A_c_105_n
+ PM_SKY130_FD_SC_LP__BUFLP_1%A
x_PM_SKY130_FD_SC_LP__BUFLP_1%X N_X_M1003_s N_X_M1002_s X X X X X X X
+ N_X_c_138_n PM_SKY130_FD_SC_LP__BUFLP_1%X
x_PM_SKY130_FD_SC_LP__BUFLP_1%VPWR N_VPWR_M1005_d N_VPWR_c_157_n VPWR
+ N_VPWR_c_158_n N_VPWR_c_159_n N_VPWR_c_156_n N_VPWR_c_161_n
+ PM_SKY130_FD_SC_LP__BUFLP_1%VPWR
x_PM_SKY130_FD_SC_LP__BUFLP_1%VGND N_VGND_M1000_d N_VGND_c_186_n VGND
+ N_VGND_c_187_n N_VGND_c_188_n N_VGND_c_189_n N_VGND_c_190_n
+ PM_SKY130_FD_SC_LP__BUFLP_1%VGND
cc_1 VNB N_A_86_21#_M1003_g 0.0304496f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_2 VNB N_A_86_21#_M1002_g 0.00838554f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_3 VNB N_A_86_21#_c_38_n 0.00943917f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.44
cc_4 VNB N_A_86_21#_M1005_g 0.00771979f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.465
cc_5 VNB N_A_86_21#_c_40_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.44
cc_6 VNB N_A_86_21#_c_41_n 0.00329981f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.35
cc_7 VNB N_A_86_21#_c_42_n 0.0305808f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.35
cc_8 VNB N_A_86_21#_c_43_n 0.0317039f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=2.16
cc_9 VNB N_A_86_21#_c_44_n 0.018522f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=0.825
cc_10 VNB N_A_86_21#_c_45_n 0.0175959f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.185
cc_11 VNB N_A_c_100_n 0.0179359f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.655
cc_12 VNB N_A_M1007_g 0.00715834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_c_102_n 0.0203703f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_14 VNB N_A_M1001_g 0.00677055f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_15 VNB N_A_c_104_n 5.6343e-19 $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.35
cc_16 VNB N_A_c_105_n 0.0363177f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.35
cc_17 VNB N_X_c_138_n 0.0555506f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.465
cc_18 VNB N_VPWR_c_156_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.465
cc_19 VNB N_VGND_c_186_n 0.0150056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_187_n 0.0279551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_188_n 0.0364828f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.185
cc_22 VNB N_VGND_c_189_n 0.164917f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.655
cc_23 VNB N_VGND_c_190_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.465
cc_24 VPB N_A_86_21#_M1002_g 0.0239104f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_25 VPB N_A_86_21#_M1005_g 0.0220789f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=2.465
cc_26 VPB N_A_86_21#_c_43_n 0.0463216f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=2.16
cc_27 VPB N_A_M1007_g 0.0294441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_A_M1001_g 0.0314603f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_29 VPB N_A_c_104_n 0.00816223f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.35
cc_30 VPB N_X_c_138_n 0.0547566f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=2.465
cc_31 VPB N_VPWR_c_157_n 0.0200748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_158_n 0.0279551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_159_n 0.0346039f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=2.465
cc_34 VPB N_VPWR_c_156_n 0.0648065f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=2.465
cc_35 VPB N_VPWR_c_161_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.015
cc_36 N_A_86_21#_c_41_n N_A_c_100_n 0.00387076f $X=0.985 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_37 N_A_86_21#_c_50_p N_A_c_100_n 0.0138311f $X=1.905 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_38 N_A_86_21#_c_44_n N_A_c_100_n 0.00104262f $X=2.07 $Y=0.825 $X2=-0.19
+ $Y2=-0.245
cc_39 N_A_86_21#_c_45_n N_A_c_100_n 0.0161693f $X=0.985 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_40 N_A_86_21#_M1005_g N_A_M1007_g 0.0209225f $X=0.895 $Y=2.465 $X2=0 $Y2=0
cc_41 N_A_86_21#_c_50_p N_A_c_102_n 0.0121016f $X=1.905 $Y=0.93 $X2=0 $Y2=0
cc_42 N_A_86_21#_c_43_n N_A_c_102_n 0.0267409f $X=2.07 $Y=2.16 $X2=0 $Y2=0
cc_43 N_A_86_21#_c_44_n N_A_c_102_n 0.00654625f $X=2.07 $Y=0.825 $X2=0 $Y2=0
cc_44 N_A_86_21#_M1005_g N_A_c_104_n 0.00187809f $X=0.895 $Y=2.465 $X2=0 $Y2=0
cc_45 N_A_86_21#_c_41_n N_A_c_104_n 0.0160099f $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_46 N_A_86_21#_c_42_n N_A_c_104_n 0.00119681f $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_47 N_A_86_21#_c_50_p N_A_c_104_n 0.0229327f $X=1.905 $Y=0.93 $X2=0 $Y2=0
cc_48 N_A_86_21#_c_43_n N_A_c_104_n 0.0828479f $X=2.07 $Y=2.16 $X2=0 $Y2=0
cc_49 N_A_86_21#_c_41_n N_A_c_105_n 0.00137729f $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_50 N_A_86_21#_c_42_n N_A_c_105_n 0.0184429f $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_51 N_A_86_21#_c_50_p N_A_c_105_n 4.22969e-19 $X=1.905 $Y=0.93 $X2=0 $Y2=0
cc_52 N_A_86_21#_M1003_g N_X_c_138_n 0.0258467f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_53 N_A_86_21#_M1002_g N_X_c_138_n 0.0358711f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_54 N_A_86_21#_M1005_g N_X_c_138_n 0.00504859f $X=0.895 $Y=2.465 $X2=0 $Y2=0
cc_55 N_A_86_21#_c_40_n N_X_c_138_n 0.00657988f $X=0.505 $Y=1.44 $X2=0 $Y2=0
cc_56 N_A_86_21#_c_41_n N_X_c_138_n 0.0202513f $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_57 N_A_86_21#_c_70_p N_X_c_138_n 0.00732751f $X=1.15 $Y=0.93 $X2=0 $Y2=0
cc_58 N_A_86_21#_c_45_n N_X_c_138_n 0.00320916f $X=0.985 $Y=1.185 $X2=0 $Y2=0
cc_59 N_A_86_21#_M1002_g N_VPWR_c_157_n 0.00475339f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_60 N_A_86_21#_M1005_g N_VPWR_c_157_n 0.0303995f $X=0.895 $Y=2.465 $X2=0 $Y2=0
cc_61 N_A_86_21#_c_41_n N_VPWR_c_157_n 0.0116937f $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_62 N_A_86_21#_c_42_n N_VPWR_c_157_n 0.00132119f $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_63 N_A_86_21#_M1002_g N_VPWR_c_158_n 0.0054895f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A_86_21#_M1005_g N_VPWR_c_158_n 0.00486043f $X=0.895 $Y=2.465 $X2=0
+ $Y2=0
cc_65 N_A_86_21#_c_43_n N_VPWR_c_159_n 0.0048213f $X=2.07 $Y=2.16 $X2=0 $Y2=0
cc_66 N_A_86_21#_M1002_g N_VPWR_c_156_n 0.0108635f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_67 N_A_86_21#_M1005_g N_VPWR_c_156_n 0.00823808f $X=0.895 $Y=2.465 $X2=0
+ $Y2=0
cc_68 N_A_86_21#_c_43_n N_VPWR_c_156_n 0.00741569f $X=2.07 $Y=2.16 $X2=0 $Y2=0
cc_69 N_A_86_21#_c_41_n N_VGND_M1000_d 7.81051e-19 $X=0.985 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_70 N_A_86_21#_c_50_p N_VGND_M1000_d 0.00994505f $X=1.905 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A_86_21#_c_70_p N_VGND_M1000_d 0.00133164f $X=1.15 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_86_21#_M1003_g N_VGND_c_186_n 0.00237575f $X=0.505 $Y=0.655 $X2=0
+ $Y2=0
cc_73 N_A_86_21#_c_42_n N_VGND_c_186_n 5.99084e-19 $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_74 N_A_86_21#_c_50_p N_VGND_c_186_n 0.00983688f $X=1.905 $Y=0.93 $X2=0 $Y2=0
cc_75 N_A_86_21#_c_70_p N_VGND_c_186_n 0.0127977f $X=1.15 $Y=0.93 $X2=0 $Y2=0
cc_76 N_A_86_21#_c_44_n N_VGND_c_186_n 0.00113117f $X=2.07 $Y=0.825 $X2=0 $Y2=0
cc_77 N_A_86_21#_c_45_n N_VGND_c_186_n 0.0143371f $X=0.985 $Y=1.185 $X2=0 $Y2=0
cc_78 N_A_86_21#_M1003_g N_VGND_c_187_n 0.0054895f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_79 N_A_86_21#_c_45_n N_VGND_c_187_n 0.00486043f $X=0.985 $Y=1.185 $X2=0 $Y2=0
cc_80 N_A_86_21#_c_44_n N_VGND_c_188_n 0.00652217f $X=2.07 $Y=0.825 $X2=0 $Y2=0
cc_81 N_A_86_21#_M1003_g N_VGND_c_189_n 0.0108635f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_82 N_A_86_21#_c_50_p N_VGND_c_189_n 0.0211757f $X=1.905 $Y=0.93 $X2=0 $Y2=0
cc_83 N_A_86_21#_c_70_p N_VGND_c_189_n 0.00469772f $X=1.15 $Y=0.93 $X2=0 $Y2=0
cc_84 N_A_86_21#_c_44_n N_VGND_c_189_n 0.00986372f $X=2.07 $Y=0.825 $X2=0 $Y2=0
cc_85 N_A_86_21#_c_45_n N_VGND_c_189_n 0.00451072f $X=0.985 $Y=1.185 $X2=0 $Y2=0
cc_86 N_A_86_21#_c_50_p A_308_131# 0.00374661f $X=1.905 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A_M1007_g N_VPWR_c_157_n 0.0078972f $X=1.465 $Y=2.335 $X2=0 $Y2=0
cc_88 N_A_c_104_n N_VPWR_c_157_n 0.0849057f $X=1.61 $Y=1.35 $X2=0 $Y2=0
cc_89 N_A_M1007_g N_VPWR_c_159_n 0.00183215f $X=1.465 $Y=2.335 $X2=0 $Y2=0
cc_90 N_A_M1001_g N_VPWR_c_159_n 0.00359134f $X=1.855 $Y=2.335 $X2=0 $Y2=0
cc_91 N_A_c_104_n N_VPWR_c_159_n 0.0113794f $X=1.61 $Y=1.35 $X2=0 $Y2=0
cc_92 N_A_M1007_g N_VPWR_c_156_n 0.00170177f $X=1.465 $Y=2.335 $X2=0 $Y2=0
cc_93 N_A_M1001_g N_VPWR_c_156_n 0.00413287f $X=1.855 $Y=2.335 $X2=0 $Y2=0
cc_94 N_A_c_104_n N_VPWR_c_156_n 0.0121336f $X=1.61 $Y=1.35 $X2=0 $Y2=0
cc_95 N_A_c_100_n N_VGND_c_186_n 0.00350177f $X=1.465 $Y=1.185 $X2=0 $Y2=0
cc_96 N_A_c_100_n N_VGND_c_188_n 0.00399858f $X=1.465 $Y=1.185 $X2=0 $Y2=0
cc_97 N_A_c_102_n N_VGND_c_188_n 0.00385415f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_98 N_A_c_100_n N_VGND_c_189_n 0.0046122f $X=1.465 $Y=1.185 $X2=0 $Y2=0
cc_99 N_A_c_102_n N_VGND_c_189_n 0.0046122f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_100 N_X_c_138_n N_VPWR_c_157_n 0.0399176f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_101 N_X_c_138_n N_VPWR_c_158_n 0.0210192f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_102 N_X_M1002_s N_VPWR_c_156_n 0.00231914f $X=0.145 $Y=1.835 $X2=0 $Y2=0
cc_103 N_X_c_138_n N_VPWR_c_156_n 0.0125689f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_104 N_X_c_138_n N_VGND_c_186_n 0.0133059f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_105 N_X_c_138_n N_VGND_c_187_n 0.0210192f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_106 N_X_M1003_s N_VGND_c_189_n 0.00231914f $X=0.145 $Y=0.235 $X2=0 $Y2=0
cc_107 N_X_c_138_n N_VGND_c_189_n 0.0125689f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_108 A_116_367# N_VPWR_c_156_n 0.010279f $X=0.58 $Y=1.835 $X2=2.16 $Y2=3.33
cc_109 A_116_47# N_VGND_c_189_n 0.010279f $X=0.58 $Y=0.235 $X2=2.16 $Y2=0
