* File: sky130_fd_sc_lp__nand4_lp.pxi.spice
* Created: Wed Sep  2 10:05:48 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4_LP%D N_D_M1005_g N_D_M1002_g D N_D_c_51_n N_D_c_52_n
+ PM_SKY130_FD_SC_LP__NAND4_LP%D
x_PM_SKY130_FD_SC_LP__NAND4_LP%C N_C_M1006_g N_C_M1000_g N_C_c_78_n N_C_c_79_n
+ N_C_c_80_n C C C N_C_c_82_n PM_SKY130_FD_SC_LP__NAND4_LP%C
x_PM_SKY130_FD_SC_LP__NAND4_LP%B N_B_M1003_g N_B_c_120_n N_B_M1007_g N_B_c_122_n
+ N_B_c_123_n B B B N_B_c_125_n PM_SKY130_FD_SC_LP__NAND4_LP%B
x_PM_SKY130_FD_SC_LP__NAND4_LP%A N_A_M1001_g N_A_M1004_g A A N_A_c_165_n
+ N_A_c_166_n PM_SKY130_FD_SC_LP__NAND4_LP%A
x_PM_SKY130_FD_SC_LP__NAND4_LP%VPWR N_VPWR_M1005_s N_VPWR_M1000_d N_VPWR_M1004_d
+ N_VPWR_c_195_n N_VPWR_c_196_n N_VPWR_c_197_n N_VPWR_c_198_n N_VPWR_c_199_n
+ N_VPWR_c_200_n VPWR N_VPWR_c_201_n N_VPWR_c_202_n N_VPWR_c_194_n
+ PM_SKY130_FD_SC_LP__NAND4_LP%VPWR
x_PM_SKY130_FD_SC_LP__NAND4_LP%Y N_Y_M1001_d N_Y_M1005_d N_Y_M1007_d N_Y_c_234_n
+ N_Y_c_235_n N_Y_c_236_n N_Y_c_237_n N_Y_c_253_n N_Y_c_232_n N_Y_c_238_n Y Y Y
+ PM_SKY130_FD_SC_LP__NAND4_LP%Y
x_PM_SKY130_FD_SC_LP__NAND4_LP%VGND N_VGND_M1002_s N_VGND_c_288_n N_VGND_c_289_n
+ VGND N_VGND_c_290_n N_VGND_c_291_n PM_SKY130_FD_SC_LP__NAND4_LP%VGND
cc_1 VNB N_D_M1005_g 0.0151994f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.545
cc_2 VNB N_D_M1002_g 0.025878f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_3 VNB N_D_c_51_n 0.0801597f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.99
cc_4 VNB N_D_c_52_n 0.0291871f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.99
cc_5 VNB N_C_M1000_g 0.0144108f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_6 VNB N_C_c_78_n 0.0167706f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_C_c_79_n 0.0213929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_C_c_80_n 0.0126979f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.99
cc_9 VNB C 0.00632868f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.99
cc_10 VNB N_C_c_82_n 0.0156432f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.16
cc_11 VNB N_B_c_120_n 0.0138802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_M1007_g 0.0143666f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_13 VNB N_B_c_122_n 0.0182558f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_B_c_123_n 0.0238729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB B 0.00153492f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.99
cc_16 VNB N_B_c_125_n 0.0167626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_M1001_g 0.0481698f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.545
cc_18 VNB N_A_c_165_n 0.0719506f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.825
cc_19 VNB N_A_c_166_n 0.0268366f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.495
cc_20 VNB N_VPWR_c_194_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_232_n 0.00690682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Y 0.0294351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_288_n 0.0138745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_289_n 0.0183356f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_25 VNB N_VGND_c_290_n 0.0638673f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.495
cc_26 VNB N_VGND_c_291_n 0.173695f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.16
cc_27 VPB N_D_M1005_g 0.0518981f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.545
cc_28 VPB N_C_M1000_g 0.0376326f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.445
cc_29 VPB N_B_M1007_g 0.0376854f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.445
cc_30 VPB N_A_M1004_g 0.0408091f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.445
cc_31 VPB N_A_c_165_n 0.0250555f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=0.825
cc_32 VPB N_A_c_166_n 0.0121459f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.495
cc_33 VPB N_VPWR_c_195_n 0.0119948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_196_n 0.0479643f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.99
cc_35 VPB N_VPWR_c_197_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.16
cc_36 VPB N_VPWR_c_198_n 0.00446486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_199_n 0.0155402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_200_n 0.0497319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_201_n 0.0210253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_202_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_194_n 0.0557981f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_Y_c_234_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.99
cc_43 VPB N_Y_c_235_n 0.00991661f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.16
cc_44 VPB N_Y_c_236_n 0.00908361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_Y_c_237_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_Y_c_238_n 0.00764869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 N_D_c_51_n N_C_M1000_g 0.0361379f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_48 N_D_c_52_n N_C_M1000_g 2.92318e-19 $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_49 N_D_M1002_g N_C_c_78_n 0.0380062f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_50 N_D_M1002_g C 0.0018677f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_51 N_D_c_51_n C 0.00249171f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_52 N_D_c_52_n C 0.0264703f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_53 N_D_c_51_n N_C_c_82_n 0.0391014f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_54 N_D_c_52_n N_C_c_82_n 0.00171651f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_55 N_D_M1005_g N_VPWR_c_196_n 0.0239979f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_56 N_D_c_51_n N_VPWR_c_196_n 0.00456474f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_57 N_D_c_52_n N_VPWR_c_196_n 0.012628f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_58 N_D_M1005_g N_VPWR_c_197_n 0.00769046f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_59 N_D_M1005_g N_VPWR_c_198_n 9.45383e-19 $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_60 N_D_M1005_g N_VPWR_c_194_n 0.0134474f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_61 N_D_M1005_g N_Y_c_234_n 0.0289408f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_62 N_D_M1005_g N_Y_c_236_n 0.0115348f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_63 N_D_M1002_g N_VGND_c_289_n 0.0131971f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_64 N_D_c_51_n N_VGND_c_289_n 0.00758869f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_65 N_D_c_52_n N_VGND_c_289_n 0.0240373f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_66 N_D_M1002_g N_VGND_c_290_n 0.00486043f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_67 N_D_M1002_g N_VGND_c_291_n 0.00779546f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_68 N_D_c_51_n N_VGND_c_291_n 7.74273e-19 $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_69 N_D_c_52_n N_VGND_c_291_n 0.0048771f $X=0.385 $Y=0.99 $X2=0 $Y2=0
cc_70 N_C_c_80_n N_B_c_120_n 0.0117523f $X=1.065 $Y=1.435 $X2=0 $Y2=0
cc_71 N_C_M1000_g N_B_M1007_g 0.0344708f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_72 N_C_c_78_n N_B_c_122_n 0.0186614f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_73 C N_B_c_122_n 0.00652031f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_74 N_C_c_79_n N_B_c_123_n 0.0117523f $X=1.065 $Y=1.27 $X2=0 $Y2=0
cc_75 N_C_c_78_n B 2.96101e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_76 C B 0.0760026f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_77 N_C_c_82_n B 7.56445e-19 $X=1.065 $Y=0.93 $X2=0 $Y2=0
cc_78 N_C_c_82_n N_B_c_125_n 0.0117523f $X=1.065 $Y=0.93 $X2=0 $Y2=0
cc_79 N_C_M1000_g N_VPWR_c_196_n 9.45383e-19 $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_80 N_C_M1000_g N_VPWR_c_197_n 0.00769046f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_81 N_C_M1000_g N_VPWR_c_198_n 0.022508f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_82 N_C_M1000_g N_VPWR_c_194_n 0.0134474f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_83 N_C_M1000_g N_Y_c_234_n 0.0238595f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_84 N_C_M1000_g N_Y_c_235_n 0.0184366f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_85 C N_Y_c_235_n 0.0174964f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_86 N_C_M1000_g N_Y_c_236_n 0.0028345f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_87 N_C_c_80_n N_Y_c_236_n 5.18336e-19 $X=1.065 $Y=1.435 $X2=0 $Y2=0
cc_88 C N_Y_c_236_n 0.00634621f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_89 N_C_M1000_g N_Y_c_237_n 0.00105185f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_90 N_C_c_78_n N_VGND_c_289_n 0.00264669f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_91 C N_VGND_c_289_n 0.00843548f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_92 N_C_c_78_n N_VGND_c_290_n 0.00394642f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_93 C N_VGND_c_290_n 0.0111981f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_94 N_C_c_82_n N_VGND_c_290_n 4.70837e-19 $X=1.065 $Y=0.93 $X2=0 $Y2=0
cc_95 N_C_c_78_n N_VGND_c_291_n 0.00586352f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_96 C N_VGND_c_291_n 0.0127858f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_97 C A_210_47# 0.00489415f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_98 N_B_c_122_n N_A_M1001_g 0.0176431f $X=1.635 $Y=0.765 $X2=0 $Y2=0
cc_99 B N_A_M1001_g 0.00186938f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_100 N_B_c_125_n N_A_M1001_g 0.017633f $X=1.635 $Y=0.93 $X2=0 $Y2=0
cc_101 N_B_M1007_g N_A_c_165_n 0.033445f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_102 N_B_c_123_n N_A_c_165_n 0.017633f $X=1.635 $Y=1.27 $X2=0 $Y2=0
cc_103 N_B_M1007_g N_VPWR_c_198_n 0.0215101f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_104 N_B_M1007_g N_VPWR_c_201_n 0.00804781f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_105 N_B_M1007_g N_VPWR_c_194_n 0.0140691f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_106 N_B_M1007_g N_Y_c_234_n 0.00104367f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_107 N_B_c_120_n N_Y_c_235_n 2.52689e-19 $X=1.635 $Y=1.435 $X2=0 $Y2=0
cc_108 N_B_M1007_g N_Y_c_235_n 0.0187384f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_109 B N_Y_c_235_n 0.0153701f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_110 N_B_M1007_g N_Y_c_237_n 0.0244878f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_111 N_B_c_122_n N_Y_c_253_n 0.00474793f $X=1.635 $Y=0.765 $X2=0 $Y2=0
cc_112 B N_Y_c_253_n 0.0192422f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_113 N_B_M1007_g N_Y_c_232_n 0.00474141f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_114 N_B_c_122_n N_Y_c_232_n 2.0904e-19 $X=1.635 $Y=0.765 $X2=0 $Y2=0
cc_115 B N_Y_c_232_n 0.0549769f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_116 N_B_c_125_n N_Y_c_232_n 0.00379786f $X=1.635 $Y=0.93 $X2=0 $Y2=0
cc_117 N_B_c_120_n N_Y_c_238_n 2.93245e-19 $X=1.635 $Y=1.435 $X2=0 $Y2=0
cc_118 N_B_M1007_g N_Y_c_238_n 0.0028345f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_119 B N_Y_c_238_n 0.00428354f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_120 N_B_c_122_n N_VGND_c_290_n 0.00394642f $X=1.635 $Y=0.765 $X2=0 $Y2=0
cc_121 B N_VGND_c_290_n 0.00930091f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_122 N_B_c_125_n N_VGND_c_290_n 4.68308e-19 $X=1.635 $Y=0.93 $X2=0 $Y2=0
cc_123 N_B_c_122_n N_VGND_c_291_n 0.00629536f $X=1.635 $Y=0.765 $X2=0 $Y2=0
cc_124 B N_VGND_c_291_n 0.0106938f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_125 B A_324_47# 0.00361625f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_126 N_A_M1004_g N_VPWR_c_198_n 9.38445e-19 $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_127 N_A_M1004_g N_VPWR_c_200_n 0.0270912f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_128 N_A_c_165_n N_VPWR_c_200_n 0.00246051f $X=2.495 $Y=1.275 $X2=0 $Y2=0
cc_129 N_A_c_166_n N_VPWR_c_200_n 0.022184f $X=2.495 $Y=1.275 $X2=0 $Y2=0
cc_130 N_A_M1004_g N_VPWR_c_201_n 0.00741874f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_131 N_A_M1004_g N_VPWR_c_194_n 0.0132069f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_132 N_A_M1004_g N_Y_c_237_n 0.0329166f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_133 N_A_M1001_g N_Y_c_253_n 0.00841515f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A_M1001_g N_Y_c_232_n 0.0224889f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_135 N_A_c_165_n N_Y_c_232_n 0.0161678f $X=2.495 $Y=1.275 $X2=0 $Y2=0
cc_136 N_A_c_166_n N_Y_c_232_n 0.0393073f $X=2.495 $Y=1.275 $X2=0 $Y2=0
cc_137 N_A_M1004_g N_Y_c_238_n 0.0042969f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_138 N_A_c_165_n N_Y_c_238_n 0.00390814f $X=2.495 $Y=1.275 $X2=0 $Y2=0
cc_139 N_A_c_166_n N_Y_c_238_n 0.00815308f $X=2.495 $Y=1.275 $X2=0 $Y2=0
cc_140 N_A_M1001_g Y 0.00434769f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A_c_165_n Y 0.00691503f $X=2.495 $Y=1.275 $X2=0 $Y2=0
cc_142 N_A_c_166_n Y 0.018248f $X=2.495 $Y=1.275 $X2=0 $Y2=0
cc_143 N_A_M1001_g N_VGND_c_290_n 0.00359812f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A_M1001_g N_VGND_c_291_n 0.00697519f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_145 N_VPWR_c_196_n N_Y_c_234_n 0.0685263f $X=0.3 $Y=2.19 $X2=0 $Y2=0
cc_146 N_VPWR_c_197_n N_Y_c_234_n 0.021949f $X=1.195 $Y=3.33 $X2=0 $Y2=0
cc_147 N_VPWR_c_198_n N_Y_c_234_n 0.0685263f $X=1.36 $Y=2.19 $X2=0 $Y2=0
cc_148 N_VPWR_c_194_n N_Y_c_234_n 0.0124703f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_149 N_VPWR_c_198_n N_Y_c_235_n 0.0262847f $X=1.36 $Y=2.19 $X2=0 $Y2=0
cc_150 N_VPWR_c_198_n N_Y_c_237_n 0.0670852f $X=1.36 $Y=2.19 $X2=0 $Y2=0
cc_151 N_VPWR_c_200_n N_Y_c_237_n 0.0401237f $X=2.495 $Y=2.19 $X2=0 $Y2=0
cc_152 N_VPWR_c_201_n N_Y_c_237_n 0.0273857f $X=2.33 $Y=3.33 $X2=0 $Y2=0
cc_153 N_VPWR_c_194_n N_Y_c_237_n 0.0153677f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_154 N_Y_c_253_n N_VGND_c_290_n 0.00914355f $X=2.065 $Y=0.675 $X2=0 $Y2=0
cc_155 Y N_VGND_c_290_n 0.0368266f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_156 N_Y_M1001_d N_VGND_c_291_n 0.00233022f $X=2.19 $Y=0.235 $X2=0 $Y2=0
cc_157 N_Y_c_253_n N_VGND_c_291_n 0.00607116f $X=2.065 $Y=0.675 $X2=0 $Y2=0
cc_158 Y N_VGND_c_291_n 0.0228969f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_159 N_Y_c_253_n A_324_47# 0.00486731f $X=2.065 $Y=0.675 $X2=-0.19 $Y2=-0.245
cc_160 N_VGND_c_291_n A_132_47# 0.00960097f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_161 N_VGND_c_291_n A_210_47# 0.00995342f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_162 N_VGND_c_291_n A_324_47# 0.00984608f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
