* File: sky130_fd_sc_lp__nand3b_lp.pex.spice
* Created: Fri Aug 28 10:50:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3B_LP%A_90_247# 1 2 9 13 15 16 17 20 21 23 24 29
+ 34 35 36
c67 23 0 1.41654e-19 $X=2.435 $Y=1.285
c68 9 0 9.90479e-20 $X=0.625 $Y=2.58
r69 34 35 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=2.225
+ $X2=2.56 $Y2=2.06
r70 31 36 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.68 $Y=1.37
+ $X2=2.6 $Y2=1.285
r71 31 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.68 $Y=1.37 $X2=2.68
+ $Y2=2.06
r72 27 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=1.2 $X2=2.6
+ $Y2=1.285
r73 27 29 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.6 $Y=1.2 $X2=2.6
+ $Y2=0.955
r74 23 36 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.435 $Y=1.285
+ $X2=2.6 $Y2=1.285
r75 23 24 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=2.435 $Y=1.285
+ $X2=0.78 $Y2=1.285
r76 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.615
+ $Y=1.4 $X2=0.615 $Y2=1.4
r77 18 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.615 $Y=1.37
+ $X2=0.78 $Y2=1.285
r78 18 20 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.615 $Y=1.37
+ $X2=0.615 $Y2=1.4
r79 16 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.615 $Y=1.74
+ $X2=0.615 $Y2=1.4
r80 16 17 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=1.74
+ $X2=0.615 $Y2=1.905
r81 15 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=1.235
+ $X2=0.615 $Y2=1.4
r82 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.705 $Y=0.915
+ $X2=0.705 $Y2=1.235
r83 9 17 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.625 $Y=2.58
+ $X2=0.625 $Y2=1.905
r84 2 34 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.38
+ $Y=2.08 $X2=2.52 $Y2=2.225
r85 1 29 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.705 $X2=2.6 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_LP%B 3 7 9 12
c36 9 0 9.90479e-20 $X=1.2 $Y=1.665
c37 7 0 6.44281e-20 $X=1.155 $Y=2.58
c38 3 0 3.97458e-20 $X=1.095 $Y=0.915
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.755
+ $X2=1.155 $Y2=1.59
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.755 $X2=1.155 $Y2=1.755
r41 9 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.155 $Y=1.665
+ $X2=1.155 $Y2=1.755
r42 5 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.92
+ $X2=1.155 $Y2=1.755
r43 5 7 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.155 $Y=1.92
+ $X2=1.155 $Y2=2.58
r44 3 14 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.095 $Y=0.915
+ $X2=1.095 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_LP%C 1 3 8 12 14 15 19 21
c43 15 0 3.97458e-20 $X=2.16 $Y=1.665
c44 1 0 6.90867e-20 $X=1.485 $Y=1.2
r45 19 22 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.715
+ $X2=1.725 $Y2=1.88
r46 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.715
+ $X2=1.725 $Y2=1.55
r47 14 15 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.715
+ $X2=2.16 $Y2=1.715
r48 14 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.715 $X2=1.725 $Y2=1.715
r49 10 12 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.485 $Y=1.275
+ $X2=1.635 $Y2=1.275
r50 8 22 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.685 $Y=2.58 $X2=1.685
+ $Y2=1.88
r51 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.635 $Y=1.35
+ $X2=1.635 $Y2=1.275
r52 4 21 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.635 $Y=1.35 $X2=1.635
+ $Y2=1.55
r53 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.485 $Y=1.2
+ $X2=1.485 $Y2=1.275
r54 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.485 $Y=1.2 $X2=1.485
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_LP%A_N 1 3 6 11 13 14 15 23
c37 23 0 1.41654e-19 $X=2.385 $Y=0.43
c38 15 0 6.90867e-20 $X=2.64 $Y=0.555
r39 21 23 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.21 $Y=0.43
+ $X2=2.385 $Y2=0.43
r40 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=0.43 $X2=2.21 $Y2=0.43
r41 18 21 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.025 $Y=0.43
+ $X2=2.21 $Y2=0.43
r42 15 22 12.2358 $w=4.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.64 $Y=0.467
+ $X2=2.21 $Y2=0.467
r43 14 22 1.42277 $w=4.03e-07 $l=5e-08 $layer=LI1_cond $X=2.16 $Y=0.467 $X2=2.21
+ $Y2=0.467
r44 12 13 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.295 $Y=1.495
+ $X2=2.295 $Y2=1.645
r45 11 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.385 $Y=0.915
+ $X2=2.385 $Y2=1.495
r46 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=0.595
+ $X2=2.385 $Y2=0.43
r47 8 11 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.385 $Y=0.595
+ $X2=2.385 $Y2=0.915
r48 6 13 232.304 $w=2.5e-07 $l=9.35e-07 $layer=POLY_cond $X=2.255 $Y=2.58
+ $X2=2.255 $Y2=1.645
r49 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.025 $Y=0.595
+ $X2=2.025 $Y2=0.43
r50 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.025 $Y=0.595
+ $X2=2.025 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_LP%Y 1 2 3 10 11 14 19 21 22 23 24
c44 19 0 6.44281e-20 $X=0.36 $Y=2.25
r45 23 24 9.89858 $w=5.78e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=0.73 $X2=1.2
+ $Y2=0.73
r46 23 32 4.74307 $w=5.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.72 $Y=0.73
+ $X2=0.49 $Y2=0.73
r47 22 29 2.24098 $w=5.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.185 $Y=0.73
+ $X2=0.27 $Y2=0.73
r48 22 32 3.98005 $w=5.78e-07 $l=1.93e-07 $layer=LI1_cond $X=0.297 $Y=0.73
+ $X2=0.49 $Y2=0.73
r49 22 29 0.556795 $w=5.78e-07 $l=2.7e-08 $layer=LI1_cond $X=0.297 $Y=0.73
+ $X2=0.27 $Y2=0.73
r50 15 19 3.41642 $w=1.7e-07 $l=2.16963e-07 $layer=LI1_cond $X=0.525 $Y=2.185
+ $X2=0.312 $Y2=2.177
r51 14 21 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=2.185
+ $X2=1.42 $Y2=2.185
r52 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.255 $Y=2.185
+ $X2=0.525 $Y2=2.185
r53 11 19 3.17288 $w=2.97e-07 $l=1.66772e-07 $layer=LI1_cond $X=0.185 $Y=2.085
+ $X2=0.312 $Y2=2.177
r54 10 22 7.64568 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=0.185 $Y=1.02
+ $X2=0.185 $Y2=0.73
r55 10 11 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=0.185 $Y=1.02
+ $X2=0.185 $Y2=2.085
r56 3 21 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=1.28
+ $Y=2.08 $X2=1.42 $Y2=2.265
r57 2 19 300 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=2 $X=0.215
+ $Y=2.08 $X2=0.36 $Y2=2.25
r58 1 32 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.345
+ $Y=0.705 $X2=0.49 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_LP%VPWR 1 2 9 13 18 19 21 22 23 33 34
r37 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r40 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 23 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 23 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 21 30 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.95 $Y2=3.33
r45 20 33 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.95 $Y2=3.33
r47 18 26 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.89 $Y2=3.33
r49 17 30 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.89 $Y2=3.33
r51 13 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.95 $Y=2.225
+ $X2=1.95 $Y2=2.935
r52 11 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=3.33
r53 11 16 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=2.935
r54 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245 $X2=0.89
+ $Y2=3.33
r55 7 9 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.89 $Y=3.245 $X2=0.89
+ $Y2=2.775
r56 2 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.81
+ $Y=2.08 $X2=1.95 $Y2=2.935
r57 2 13 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.81
+ $Y=2.08 $X2=1.95 $Y2=2.225
r58 1 9 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=0.75
+ $Y=2.08 $X2=0.89 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_LP%VGND 1 6 8 10 20 21 24
r26 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r27 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r28 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r29 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.7
+ $Y2=0
r30 18 20 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.64
+ $Y2=0
r31 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r32 13 17 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r33 12 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r34 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.7
+ $Y2=0
r36 10 16 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.2
+ $Y2=0
r37 8 25 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r38 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r39 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r40 4 6 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0.85
r41 1 6 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.705 $X2=1.7 $Y2=0.85
.ends

