* File: sky130_fd_sc_lp__and2_lp2.pxi.spice
* Created: Wed Sep  2 09:30:34 2020
* 
x_PM_SKY130_FD_SC_LP__AND2_LP2%A_99_21# N_A_99_21#_M1002_d N_A_99_21#_M1004_d
+ N_A_99_21#_c_43_n N_A_99_21#_M1001_g N_A_99_21#_M1000_g N_A_99_21#_M1006_g
+ N_A_99_21#_c_45_n N_A_99_21#_c_46_n N_A_99_21#_c_83_p N_A_99_21#_c_47_n
+ N_A_99_21#_c_48_n N_A_99_21#_c_53_n N_A_99_21#_c_54_n N_A_99_21#_c_55_n
+ N_A_99_21#_c_49_n N_A_99_21#_c_50_n PM_SKY130_FD_SC_LP__AND2_LP2%A_99_21#
x_PM_SKY130_FD_SC_LP__AND2_LP2%B N_B_M1004_g N_B_M1003_g B N_B_c_115_n
+ PM_SKY130_FD_SC_LP__AND2_LP2%B
x_PM_SKY130_FD_SC_LP__AND2_LP2%A N_A_M1002_g N_A_M1005_g A A N_A_c_152_n
+ PM_SKY130_FD_SC_LP__AND2_LP2%A
x_PM_SKY130_FD_SC_LP__AND2_LP2%X N_X_M1001_s N_X_M1000_s X X X X X X X
+ N_X_c_180_n X PM_SKY130_FD_SC_LP__AND2_LP2%X
x_PM_SKY130_FD_SC_LP__AND2_LP2%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_c_203_n
+ N_VPWR_c_204_n N_VPWR_c_205_n N_VPWR_c_206_n N_VPWR_c_207_n VPWR
+ N_VPWR_c_208_n N_VPWR_c_202_n PM_SKY130_FD_SC_LP__AND2_LP2%VPWR
x_PM_SKY130_FD_SC_LP__AND2_LP2%VGND N_VGND_M1006_d N_VGND_c_233_n VGND
+ N_VGND_c_234_n N_VGND_c_235_n N_VGND_c_236_n N_VGND_c_237_n
+ PM_SKY130_FD_SC_LP__AND2_LP2%VGND
cc_1 VNB N_A_99_21#_c_43_n 0.0350817f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.775
cc_2 VNB N_A_99_21#_M1000_g 0.0115564f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.545
cc_3 VNB N_A_99_21#_c_45_n 0.0192025f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.925
cc_4 VNB N_A_99_21#_c_46_n 0.0186478f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.485
cc_5 VNB N_A_99_21#_c_47_n 0.00344355f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_6 VNB N_A_99_21#_c_48_n 0.0333322f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.9
cc_7 VNB N_A_99_21#_c_49_n 0.0216047f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=0.47
cc_8 VNB N_A_99_21#_c_50_n 0.0315214f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.98
cc_9 VNB N_B_M1004_g 0.0105455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_M1003_g 0.0362229f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.775
cc_11 VNB B 0.00542876f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.445
cc_12 VNB N_B_c_115_n 0.025981f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.545
cc_13 VNB N_A_M1002_g 0.0470233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A 0.0273558f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.445
cc_15 VNB N_A_c_152_n 0.0596194f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.775
cc_16 VNB X 0.0515624f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.775
cc_17 VNB N_X_c_180_n 0.0160497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_202_n 0.103974f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=0.815
cc_19 VNB N_VGND_c_233_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_234_n 0.0286414f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.485
cc_21 VNB N_VGND_c_235_n 0.0327565f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.925
cc_22 VNB N_VGND_c_236_n 0.157267f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.775
cc_23 VNB N_VGND_c_237_n 0.00437061f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.485
cc_24 VPB N_A_99_21#_M1000_g 0.0450391f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.545
cc_25 VPB N_A_99_21#_c_47_n 3.90385e-19 $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_26 VPB N_A_99_21#_c_53_n 0.0219615f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=1.76
cc_27 VPB N_A_99_21#_c_54_n 0.0023733f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=1.76
cc_28 VPB N_A_99_21#_c_55_n 0.00524774f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=2.19
cc_29 VPB N_B_M1004_g 0.0380384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_A_M1005_g 0.0373128f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.775
cc_31 VPB A 0.0117093f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.445
cc_32 VPB N_A_c_152_n 0.0257782f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.775
cc_33 VPB X 0.0193338f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.775
cc_34 VPB X 0.0397435f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.545
cc_35 VPB X 0.0177926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_203_n 0.00437013f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.445
cc_37 VPB N_VPWR_c_204_n 0.0131113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_205_n 0.0462566f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.445
cc_39 VPB N_VPWR_c_206_n 0.0227455f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.3
cc_40 VPB N_VPWR_c_207_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.485
cc_41 VPB N_VPWR_c_208_n 0.0196598f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=1.845
cc_42 VPB N_VPWR_c_202_n 0.0538616f $X=-0.19 $Y=1.655 $X2=1.965 $Y2=0.815
cc_43 N_A_99_21#_M1000_g N_B_M1004_g 0.0312405f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_44 N_A_99_21#_c_47_n N_B_M1004_g 0.00389427f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_45 N_A_99_21#_c_53_n N_B_M1004_g 0.0205325f $X=1.34 $Y=1.76 $X2=0 $Y2=0
cc_46 N_A_99_21#_c_55_n N_B_M1004_g 0.0236728f $X=1.505 $Y=2.19 $X2=0 $Y2=0
cc_47 N_A_99_21#_c_43_n N_B_M1003_g 0.0208471f $X=0.57 $Y=0.775 $X2=0 $Y2=0
cc_48 N_A_99_21#_c_47_n N_B_M1003_g 0.00101368f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_49 N_A_99_21#_c_48_n N_B_M1003_g 0.0117058f $X=1.8 $Y=0.9 $X2=0 $Y2=0
cc_50 N_A_99_21#_c_49_n N_B_M1003_g 0.0019366f $X=1.965 $Y=0.47 $X2=0 $Y2=0
cc_51 N_A_99_21#_c_50_n N_B_M1003_g 0.00724505f $X=0.7 $Y=0.98 $X2=0 $Y2=0
cc_52 N_A_99_21#_c_47_n B 0.0216025f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_53 N_A_99_21#_c_48_n B 0.024713f $X=1.8 $Y=0.9 $X2=0 $Y2=0
cc_54 N_A_99_21#_c_53_n B 0.0251189f $X=1.34 $Y=1.76 $X2=0 $Y2=0
cc_55 N_A_99_21#_c_50_n B 0.00198057f $X=0.7 $Y=0.98 $X2=0 $Y2=0
cc_56 N_A_99_21#_M1000_g N_B_c_115_n 4.56578e-19 $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_57 N_A_99_21#_c_47_n N_B_c_115_n 4.23476e-19 $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_58 N_A_99_21#_c_48_n N_B_c_115_n 0.00467238f $X=1.8 $Y=0.9 $X2=0 $Y2=0
cc_59 N_A_99_21#_c_53_n N_B_c_115_n 0.00211855f $X=1.34 $Y=1.76 $X2=0 $Y2=0
cc_60 N_A_99_21#_c_50_n N_B_c_115_n 0.0171423f $X=0.7 $Y=0.98 $X2=0 $Y2=0
cc_61 N_A_99_21#_c_48_n N_A_M1002_g 0.017166f $X=1.8 $Y=0.9 $X2=0 $Y2=0
cc_62 N_A_99_21#_c_49_n N_A_M1002_g 0.0129267f $X=1.965 $Y=0.47 $X2=0 $Y2=0
cc_63 N_A_99_21#_c_55_n N_A_M1005_g 0.00577342f $X=1.505 $Y=2.19 $X2=0 $Y2=0
cc_64 N_A_99_21#_c_48_n A 0.0238987f $X=1.8 $Y=0.9 $X2=0 $Y2=0
cc_65 N_A_99_21#_c_53_n A 0.0131495f $X=1.34 $Y=1.76 $X2=0 $Y2=0
cc_66 N_A_99_21#_c_48_n N_A_c_152_n 0.00341253f $X=1.8 $Y=0.9 $X2=0 $Y2=0
cc_67 N_A_99_21#_c_53_n N_A_c_152_n 0.00214617f $X=1.34 $Y=1.76 $X2=0 $Y2=0
cc_68 N_A_99_21#_c_43_n X 0.0228994f $X=0.57 $Y=0.775 $X2=0 $Y2=0
cc_69 N_A_99_21#_M1000_g X 0.00859311f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_70 N_A_99_21#_c_83_p X 0.0132565f $X=0.7 $Y=0.985 $X2=0 $Y2=0
cc_71 N_A_99_21#_c_47_n X 0.0515194f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_72 N_A_99_21#_c_54_n X 0.0140758f $X=0.865 $Y=1.76 $X2=0 $Y2=0
cc_73 N_A_99_21#_M1000_g X 0.0141535f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_74 N_A_99_21#_c_43_n N_X_c_180_n 0.00825755f $X=0.57 $Y=0.775 $X2=0 $Y2=0
cc_75 N_A_99_21#_M1000_g X 0.00489193f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_76 N_A_99_21#_c_46_n X 0.00151505f $X=0.68 $Y=1.485 $X2=0 $Y2=0
cc_77 N_A_99_21#_c_54_n X 0.00639216f $X=0.865 $Y=1.76 $X2=0 $Y2=0
cc_78 N_A_99_21#_M1000_g N_VPWR_c_203_n 0.0237294f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_79 N_A_99_21#_c_53_n N_VPWR_c_203_n 0.0219858f $X=1.34 $Y=1.76 $X2=0 $Y2=0
cc_80 N_A_99_21#_c_54_n N_VPWR_c_203_n 0.00459312f $X=0.865 $Y=1.76 $X2=0 $Y2=0
cc_81 N_A_99_21#_c_55_n N_VPWR_c_203_n 0.0685263f $X=1.505 $Y=2.19 $X2=0 $Y2=0
cc_82 N_A_99_21#_c_55_n N_VPWR_c_205_n 0.0319273f $X=1.505 $Y=2.19 $X2=0 $Y2=0
cc_83 N_A_99_21#_M1000_g N_VPWR_c_206_n 0.00769046f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_84 N_A_99_21#_c_55_n N_VPWR_c_208_n 0.0220321f $X=1.505 $Y=2.19 $X2=0 $Y2=0
cc_85 N_A_99_21#_M1000_g N_VPWR_c_202_n 0.0141652f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_86 N_A_99_21#_c_55_n N_VPWR_c_202_n 0.0125808f $X=1.505 $Y=2.19 $X2=0 $Y2=0
cc_87 N_A_99_21#_c_43_n N_VGND_c_233_n 0.0140029f $X=0.57 $Y=0.775 $X2=0 $Y2=0
cc_88 N_A_99_21#_c_48_n N_VGND_c_233_n 0.0201328f $X=1.8 $Y=0.9 $X2=0 $Y2=0
cc_89 N_A_99_21#_c_49_n N_VGND_c_233_n 0.0117218f $X=1.965 $Y=0.47 $X2=0 $Y2=0
cc_90 N_A_99_21#_c_43_n N_VGND_c_234_n 0.0103386f $X=0.57 $Y=0.775 $X2=0 $Y2=0
cc_91 N_A_99_21#_c_45_n N_VGND_c_234_n 5.88488e-19 $X=0.75 $Y=0.925 $X2=0 $Y2=0
cc_92 N_A_99_21#_c_49_n N_VGND_c_235_n 0.0198636f $X=1.965 $Y=0.47 $X2=0 $Y2=0
cc_93 N_A_99_21#_M1002_d N_VGND_c_236_n 0.00232985f $X=1.825 $Y=0.235 $X2=0
+ $Y2=0
cc_94 N_A_99_21#_c_43_n N_VGND_c_236_n 0.0119795f $X=0.57 $Y=0.775 $X2=0 $Y2=0
cc_95 N_A_99_21#_c_45_n N_VGND_c_236_n 7.97054e-19 $X=0.75 $Y=0.925 $X2=0 $Y2=0
cc_96 N_A_99_21#_c_83_p N_VGND_c_236_n 0.0115459f $X=0.7 $Y=0.985 $X2=0 $Y2=0
cc_97 N_A_99_21#_c_48_n N_VGND_c_236_n 0.0198725f $X=1.8 $Y=0.9 $X2=0 $Y2=0
cc_98 N_A_99_21#_c_49_n N_VGND_c_236_n 0.0126008f $X=1.965 $Y=0.47 $X2=0 $Y2=0
cc_99 N_B_M1003_g N_A_M1002_g 0.0374546f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_100 N_B_M1004_g A 9.36281e-19 $X=1.24 $Y=2.545 $X2=0 $Y2=0
cc_101 B A 0.0122965f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B_c_115_n A 3.24794e-19 $X=1.27 $Y=1.33 $X2=0 $Y2=0
cc_103 N_B_M1004_g N_A_c_152_n 0.0278304f $X=1.24 $Y=2.545 $X2=0 $Y2=0
cc_104 B N_A_c_152_n 0.00144188f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B_c_115_n N_A_c_152_n 0.0374546f $X=1.27 $Y=1.33 $X2=0 $Y2=0
cc_106 N_B_M1004_g X 2.76166e-19 $X=1.24 $Y=2.545 $X2=0 $Y2=0
cc_107 N_B_M1004_g N_VPWR_c_203_n 0.0225438f $X=1.24 $Y=2.545 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_VPWR_c_205_n 9.39135e-19 $X=1.24 $Y=2.545 $X2=0 $Y2=0
cc_109 N_B_M1004_g N_VPWR_c_208_n 0.00769046f $X=1.24 $Y=2.545 $X2=0 $Y2=0
cc_110 N_B_M1004_g N_VPWR_c_202_n 0.0134968f $X=1.24 $Y=2.545 $X2=0 $Y2=0
cc_111 N_B_M1003_g N_VGND_c_233_n 0.0119809f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_112 N_B_M1003_g N_VGND_c_235_n 0.00486043f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_113 N_B_M1003_g N_VGND_c_236_n 0.0044857f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A_M1005_g N_VPWR_c_203_n 8.90692e-19 $X=1.8 $Y=2.545 $X2=0 $Y2=0
cc_115 N_A_M1005_g N_VPWR_c_205_n 0.0207571f $X=1.8 $Y=2.545 $X2=0 $Y2=0
cc_116 A N_VPWR_c_205_n 0.0269634f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_117 N_A_c_152_n N_VPWR_c_205_n 0.00196918f $X=2.015 $Y=1.33 $X2=0 $Y2=0
cc_118 N_A_M1005_g N_VPWR_c_208_n 0.00802402f $X=1.8 $Y=2.545 $X2=0 $Y2=0
cc_119 N_A_M1005_g N_VPWR_c_202_n 0.014386f $X=1.8 $Y=2.545 $X2=0 $Y2=0
cc_120 N_A_M1002_g N_VGND_c_233_n 0.00228379f $X=1.75 $Y=0.445 $X2=0 $Y2=0
cc_121 N_A_M1002_g N_VGND_c_235_n 0.00549284f $X=1.75 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_M1002_g N_VGND_c_236_n 0.00734919f $X=1.75 $Y=0.445 $X2=0 $Y2=0
cc_123 X N_VPWR_c_203_n 0.0705698f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_124 X N_VPWR_c_206_n 0.0324829f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_125 X N_VPWR_c_202_n 0.0185782f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_126 N_X_c_180_n N_VGND_c_233_n 0.0125123f $X=0.355 $Y=0.45 $X2=0 $Y2=0
cc_127 N_X_c_180_n N_VGND_c_234_n 0.0231678f $X=0.355 $Y=0.45 $X2=0 $Y2=0
cc_128 N_X_M1001_s N_VGND_c_236_n 0.00233022f $X=0.21 $Y=0.235 $X2=0 $Y2=0
cc_129 N_X_c_180_n N_VGND_c_236_n 0.0149093f $X=0.355 $Y=0.45 $X2=0 $Y2=0
cc_130 A_129_47# N_VGND_c_236_n 0.00299993f $X=0.645 $Y=0.235 $X2=2.16 $Y2=0
cc_131 N_VGND_c_236_n A_287_47# 0.00343208f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
