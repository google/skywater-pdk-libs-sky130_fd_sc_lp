* File: sky130_fd_sc_lp__a211oi_0.pxi.spice
* Created: Wed Sep  2 09:17:57 2020
* 
x_PM_SKY130_FD_SC_LP__A211OI_0%A2 N_A2_c_65_n N_A2_c_66_n N_A2_c_67_n
+ N_A2_M1003_g N_A2_M1000_g N_A2_c_69_n N_A2_c_74_n A2 A2 A2 N_A2_c_71_n
+ PM_SKY130_FD_SC_LP__A211OI_0%A2
x_PM_SKY130_FD_SC_LP__A211OI_0%A1 N_A1_M1007_g N_A1_M1005_g A1 A1 A1
+ N_A1_c_106_n PM_SKY130_FD_SC_LP__A211OI_0%A1
x_PM_SKY130_FD_SC_LP__A211OI_0%B1 N_B1_M1001_g N_B1_c_145_n N_B1_M1002_g
+ N_B1_c_146_n B1 B1 N_B1_c_148_n PM_SKY130_FD_SC_LP__A211OI_0%B1
x_PM_SKY130_FD_SC_LP__A211OI_0%C1 N_C1_M1006_g N_C1_c_182_n N_C1_M1004_g
+ N_C1_c_190_n N_C1_c_191_n N_C1_c_183_n N_C1_c_184_n N_C1_c_192_n N_C1_c_185_n
+ N_C1_c_186_n N_C1_c_194_n C1 C1 C1 C1 C1 N_C1_c_188_n
+ PM_SKY130_FD_SC_LP__A211OI_0%C1
x_PM_SKY130_FD_SC_LP__A211OI_0%A_57_483# N_A_57_483#_M1003_s N_A_57_483#_M1005_d
+ N_A_57_483#_c_228_n N_A_57_483#_c_229_n N_A_57_483#_c_230_n
+ N_A_57_483#_c_231_n PM_SKY130_FD_SC_LP__A211OI_0%A_57_483#
x_PM_SKY130_FD_SC_LP__A211OI_0%VPWR N_VPWR_M1003_d N_VPWR_c_257_n VPWR
+ N_VPWR_c_258_n N_VPWR_c_256_n N_VPWR_c_260_n PM_SKY130_FD_SC_LP__A211OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A211OI_0%Y N_Y_M1007_d N_Y_M1004_d N_Y_M1006_d N_Y_c_282_n
+ N_Y_c_283_n N_Y_c_284_n N_Y_c_287_n N_Y_c_288_n N_Y_c_285_n Y Y
+ PM_SKY130_FD_SC_LP__A211OI_0%Y
x_PM_SKY130_FD_SC_LP__A211OI_0%VGND N_VGND_M1000_s N_VGND_M1001_d N_VGND_c_330_n
+ N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n VGND N_VGND_c_334_n
+ N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n PM_SKY130_FD_SC_LP__A211OI_0%VGND
cc_1 VNB N_A2_c_65_n 0.0089214f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.115
cc_2 VNB N_A2_c_66_n 0.020585f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.89
cc_3 VNB N_A2_c_67_n 0.0189051f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.89
cc_4 VNB N_A2_M1000_g 0.0240417f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.445
cc_5 VNB N_A2_c_69_n 0.0185685f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_6 VNB A2 0.0380206f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB N_A2_c_71_n 0.0306068f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_8 VNB N_A1_M1007_g 0.0409318f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.89
cc_9 VNB A1 0.0129374f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.815
cc_10 VNB N_A1_c_106_n 0.0433685f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.19
cc_11 VNB N_B1_M1001_g 0.0376952f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.89
cc_12 VNB N_B1_c_145_n 0.0214883f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.735
cc_13 VNB N_B1_c_146_n 0.00431603f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.445
cc_14 VNB B1 0.00238458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_c_148_n 0.0279435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C1_c_182_n 0.0194856f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.265
cc_17 VNB N_C1_c_183_n 0.0357189f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.445
cc_18 VNB N_C1_c_184_n 0.00863714f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.445
cc_19 VNB N_C1_c_185_n 0.0210164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C1_c_186_n 0.0249189f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.19
cc_21 VNB C1 0.0199738f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_22 VNB N_C1_c_188_n 0.0198748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_256_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.19
cc_24 VNB N_Y_c_282_n 0.00251955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_283_n 0.00977993f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_26 VNB N_Y_c_284_n 0.0119595f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_27 VNB N_Y_c_285_n 0.0127901f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB Y 0.0456563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_330_n 0.0173617f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.815
cc_30 VNB N_VGND_c_331_n 0.00522139f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.965
cc_31 VNB N_VGND_c_332_n 0.0112126f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.19
cc_32 VNB N_VGND_c_333_n 0.00510915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_334_n 0.0270577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_335_n 0.0284339f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_35 VNB N_VGND_c_336_n 0.171553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_337_n 0.00497572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A2_c_65_n 0.0317333f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.115
cc_38 VPB N_A2_M1003_g 0.0217563f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.735
cc_39 VPB N_A2_c_74_n 0.0280019f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.19
cc_40 VPB A2 0.0152097f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_41 VPB N_A1_M1005_g 0.0410404f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.735
cc_42 VPB A1 0.00461564f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.815
cc_43 VPB N_A1_c_106_n 0.0257586f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.19
cc_44 VPB N_B1_M1002_g 0.0417591f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.815
cc_45 VPB N_B1_c_146_n 0.0231929f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.445
cc_46 VPB B1 0.00992453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_C1_M1006_g 0.0242983f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.89
cc_48 VPB N_C1_c_190_n 0.0447641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_C1_c_191_n 0.0117613f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.815
cc_50 VPB N_C1_c_192_n 0.0101843f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.51
cc_51 VPB N_C1_c_186_n 0.00526959f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.19
cc_52 VPB N_C1_c_194_n 0.0197542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB C1 0.0681815f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_54 VPB N_A_57_483#_c_228_n 0.0357102f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.815
cc_55 VPB N_A_57_483#_c_229_n 0.0192009f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.445
cc_56 VPB N_A_57_483#_c_230_n 0.0119046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_57_483#_c_231_n 0.00364545f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.51
cc_58 VPB N_VPWR_c_257_n 0.00852303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_258_n 0.054226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_256_n 0.0778876f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.19
cc_61 VPB N_VPWR_c_260_n 0.0269556f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_62 VPB N_Y_c_287_n 6.48292e-19 $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.19
cc_63 VPB N_Y_c_288_n 0.00271036f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.19
cc_64 VPB N_Y_c_285_n 0.0117254f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_65 N_A2_M1000_g N_A1_M1007_g 0.044597f $X=0.665 $Y=0.445 $X2=0 $Y2=0
cc_66 N_A2_c_71_n N_A1_M1007_g 0.00201677f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_67 N_A2_c_65_n N_A1_M1005_g 0.00413016f $X=0.36 $Y=2.115 $X2=0 $Y2=0
cc_68 N_A2_c_74_n N_A1_M1005_g 0.0188617f $X=0.625 $Y=2.19 $X2=0 $Y2=0
cc_69 N_A2_c_66_n A1 0.00807882f $X=0.59 $Y=0.89 $X2=0 $Y2=0
cc_70 N_A2_M1000_g A1 0.00442283f $X=0.665 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A2_c_74_n A1 5.43156e-19 $X=0.625 $Y=2.19 $X2=0 $Y2=0
cc_72 A2 A1 0.0871402f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_73 N_A2_c_71_n A1 0.00545023f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_74 N_A2_c_66_n N_A1_c_106_n 0.00360272f $X=0.59 $Y=0.89 $X2=0 $Y2=0
cc_75 N_A2_c_74_n N_A1_c_106_n 0.00138566f $X=0.625 $Y=2.19 $X2=0 $Y2=0
cc_76 A2 N_A1_c_106_n 7.11739e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_77 N_A2_c_71_n N_A1_c_106_n 0.0342266f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_78 N_A2_M1003_g N_A_57_483#_c_228_n 0.0048436f $X=0.625 $Y=2.735 $X2=0 $Y2=0
cc_79 N_A2_c_74_n N_A_57_483#_c_228_n 0.00845809f $X=0.625 $Y=2.19 $X2=0 $Y2=0
cc_80 N_A2_c_74_n N_A_57_483#_c_229_n 0.0121202f $X=0.625 $Y=2.19 $X2=0 $Y2=0
cc_81 N_A2_c_65_n N_A_57_483#_c_230_n 0.00457385f $X=0.36 $Y=2.115 $X2=0 $Y2=0
cc_82 N_A2_c_74_n N_A_57_483#_c_230_n 0.00589646f $X=0.625 $Y=2.19 $X2=0 $Y2=0
cc_83 A2 N_A_57_483#_c_230_n 0.0155144f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A2_M1003_g N_VPWR_c_257_n 0.00290389f $X=0.625 $Y=2.735 $X2=0 $Y2=0
cc_85 N_A2_M1003_g N_VPWR_c_256_n 0.0111207f $X=0.625 $Y=2.735 $X2=0 $Y2=0
cc_86 N_A2_M1003_g N_VPWR_c_260_n 0.00545548f $X=0.625 $Y=2.735 $X2=0 $Y2=0
cc_87 N_A2_c_67_n N_VGND_c_330_n 0.00624537f $X=0.435 $Y=0.89 $X2=0 $Y2=0
cc_88 N_A2_M1000_g N_VGND_c_330_n 0.0132149f $X=0.665 $Y=0.445 $X2=0 $Y2=0
cc_89 A2 N_VGND_c_330_n 0.0123838f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_90 N_A2_M1000_g N_VGND_c_334_n 0.00486043f $X=0.665 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A2_M1000_g N_VGND_c_336_n 0.00441005f $X=0.665 $Y=0.445 $X2=0 $Y2=0
cc_92 A2 N_VGND_c_336_n 0.00886598f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_93 N_A1_M1007_g N_B1_M1001_g 0.0308587f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A1_M1005_g N_B1_c_146_n 0.0308587f $X=1.055 $Y=2.735 $X2=0 $Y2=0
cc_95 N_A1_M1007_g B1 0.00264116f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_96 A1 B1 0.021724f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_97 A1 N_B1_c_148_n 0.00228403f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_98 N_A1_c_106_n N_B1_c_148_n 0.0308587f $X=0.84 $Y=1.37 $X2=0 $Y2=0
cc_99 N_A1_M1005_g N_A_57_483#_c_229_n 0.0208818f $X=1.055 $Y=2.735 $X2=0 $Y2=0
cc_100 A1 N_A_57_483#_c_229_n 0.0310922f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_101 N_A1_c_106_n N_A_57_483#_c_229_n 0.00202686f $X=0.84 $Y=1.37 $X2=0 $Y2=0
cc_102 N_A1_M1005_g N_A_57_483#_c_231_n 0.00280552f $X=1.055 $Y=2.735 $X2=0
+ $Y2=0
cc_103 N_A1_M1005_g N_VPWR_c_257_n 0.00290389f $X=1.055 $Y=2.735 $X2=0 $Y2=0
cc_104 N_A1_M1005_g N_VPWR_c_258_n 0.00545548f $X=1.055 $Y=2.735 $X2=0 $Y2=0
cc_105 N_A1_M1005_g N_VPWR_c_256_n 0.0103349f $X=1.055 $Y=2.735 $X2=0 $Y2=0
cc_106 N_A1_M1007_g N_Y_c_282_n 0.00338039f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A1_M1007_g N_Y_c_284_n 0.00178313f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_108 A1 N_Y_c_284_n 0.0183233f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_109 N_A1_M1007_g N_VGND_c_330_n 0.00226547f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_110 A1 N_VGND_c_330_n 0.00148016f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_111 N_A1_M1007_g N_VGND_c_334_n 0.00585385f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_112 N_A1_M1007_g N_VGND_c_336_n 0.0109269f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_113 A1 N_VGND_c_336_n 0.0142595f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_114 N_B1_M1001_g N_C1_c_182_n 0.0191602f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_115 N_B1_M1002_g N_C1_c_191_n 0.0565932f $X=1.485 $Y=2.735 $X2=0 $Y2=0
cc_116 N_B1_c_146_n N_C1_c_191_n 0.00307841f $X=1.627 $Y=1.825 $X2=0 $Y2=0
cc_117 N_B1_c_148_n N_C1_c_184_n 2.78785e-19 $X=1.68 $Y=1.32 $X2=0 $Y2=0
cc_118 N_B1_c_148_n N_C1_c_185_n 0.00393922f $X=1.68 $Y=1.32 $X2=0 $Y2=0
cc_119 N_B1_c_146_n N_C1_c_186_n 0.00393922f $X=1.627 $Y=1.825 $X2=0 $Y2=0
cc_120 N_B1_c_145_n N_C1_c_188_n 0.00393922f $X=1.627 $Y=1.608 $X2=0 $Y2=0
cc_121 N_B1_M1002_g N_A_57_483#_c_229_n 0.00663186f $X=1.485 $Y=2.735 $X2=0
+ $Y2=0
cc_122 N_B1_M1002_g N_A_57_483#_c_231_n 0.0164898f $X=1.485 $Y=2.735 $X2=0 $Y2=0
cc_123 N_B1_M1002_g N_VPWR_c_258_n 0.00511358f $X=1.485 $Y=2.735 $X2=0 $Y2=0
cc_124 N_B1_M1002_g N_VPWR_c_256_n 0.00961121f $X=1.485 $Y=2.735 $X2=0 $Y2=0
cc_125 N_B1_M1001_g N_Y_c_282_n 0.00183869f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_126 N_B1_M1001_g N_Y_c_283_n 0.0154422f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_127 B1 N_Y_c_283_n 0.0274113f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_128 N_B1_c_148_n N_Y_c_283_n 0.00299308f $X=1.68 $Y=1.32 $X2=0 $Y2=0
cc_129 N_B1_M1002_g N_Y_c_287_n 0.00192575f $X=1.485 $Y=2.735 $X2=0 $Y2=0
cc_130 N_B1_M1001_g N_Y_c_285_n 0.00309041f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_131 N_B1_M1002_g N_Y_c_285_n 0.0066799f $X=1.485 $Y=2.735 $X2=0 $Y2=0
cc_132 B1 N_Y_c_285_n 0.0516337f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_133 N_B1_c_148_n N_Y_c_285_n 0.00650433f $X=1.68 $Y=1.32 $X2=0 $Y2=0
cc_134 N_B1_M1001_g Y 0.00176926f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_135 N_B1_M1001_g N_VGND_c_331_n 0.00316145f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_136 N_B1_M1001_g N_VGND_c_334_n 0.00585385f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_137 N_B1_M1001_g N_VGND_c_336_n 0.00619488f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_138 N_C1_c_191_n N_A_57_483#_c_229_n 5.86632e-19 $X=1.95 $Y=2.14 $X2=0 $Y2=0
cc_139 N_C1_M1006_g N_A_57_483#_c_231_n 0.0024211f $X=1.875 $Y=2.735 $X2=0 $Y2=0
cc_140 N_C1_M1006_g N_VPWR_c_258_n 0.00511358f $X=1.875 $Y=2.735 $X2=0 $Y2=0
cc_141 C1 N_VPWR_c_258_n 0.0159574f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_142 N_C1_M1006_g N_VPWR_c_256_n 0.0105915f $X=1.875 $Y=2.735 $X2=0 $Y2=0
cc_143 C1 N_VPWR_c_256_n 0.0147466f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_144 N_C1_c_184_n N_Y_c_283_n 0.00884902f $X=1.99 $Y=0.84 $X2=0 $Y2=0
cc_145 N_C1_M1006_g N_Y_c_287_n 0.00391162f $X=1.875 $Y=2.735 $X2=0 $Y2=0
cc_146 N_C1_c_190_n N_Y_c_287_n 0.00139575f $X=2.33 $Y=2.14 $X2=0 $Y2=0
cc_147 N_C1_M1006_g N_Y_c_288_n 0.00940891f $X=1.875 $Y=2.735 $X2=0 $Y2=0
cc_148 N_C1_M1006_g N_Y_c_285_n 0.00502273f $X=1.875 $Y=2.735 $X2=0 $Y2=0
cc_149 N_C1_c_190_n N_Y_c_285_n 0.0188194f $X=2.33 $Y=2.14 $X2=0 $Y2=0
cc_150 N_C1_c_185_n N_Y_c_285_n 0.0149636f $X=2.495 $Y=1.21 $X2=0 $Y2=0
cc_151 C1 N_Y_c_285_n 0.137929f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_152 N_C1_c_182_n Y 0.00384783f $X=1.915 $Y=0.765 $X2=0 $Y2=0
cc_153 N_C1_c_183_n Y 0.0284285f $X=2.33 $Y=0.84 $X2=0 $Y2=0
cc_154 N_C1_c_184_n Y 3.18249e-19 $X=1.99 $Y=0.84 $X2=0 $Y2=0
cc_155 N_C1_c_185_n Y 0.00926866f $X=2.495 $Y=1.21 $X2=0 $Y2=0
cc_156 C1 Y 0.0365605f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_157 N_C1_c_188_n Y 0.0014092f $X=2.495 $Y=1.375 $X2=0 $Y2=0
cc_158 N_C1_c_182_n N_VGND_c_331_n 0.00316145f $X=1.915 $Y=0.765 $X2=0 $Y2=0
cc_159 N_C1_c_182_n N_VGND_c_335_n 0.00585385f $X=1.915 $Y=0.765 $X2=0 $Y2=0
cc_160 N_C1_c_183_n N_VGND_c_335_n 0.00122753f $X=2.33 $Y=0.84 $X2=0 $Y2=0
cc_161 N_C1_c_182_n N_VGND_c_336_n 0.00756718f $X=1.915 $Y=0.765 $X2=0 $Y2=0
cc_162 N_C1_c_183_n N_VGND_c_336_n 2.04166e-19 $X=2.33 $Y=0.84 $X2=0 $Y2=0
cc_163 N_A_57_483#_c_228_n N_VPWR_c_257_n 0.00307927f $X=0.41 $Y=2.56 $X2=0
+ $Y2=0
cc_164 N_A_57_483#_c_229_n N_VPWR_c_257_n 0.0218758f $X=1.14 $Y=2.135 $X2=0
+ $Y2=0
cc_165 N_A_57_483#_c_231_n N_VPWR_c_257_n 0.00307927f $X=1.27 $Y=2.56 $X2=0
+ $Y2=0
cc_166 N_A_57_483#_c_231_n N_VPWR_c_258_n 0.0209199f $X=1.27 $Y=2.56 $X2=0 $Y2=0
cc_167 N_A_57_483#_c_228_n N_VPWR_c_256_n 0.0113912f $X=0.41 $Y=2.56 $X2=0 $Y2=0
cc_168 N_A_57_483#_c_231_n N_VPWR_c_256_n 0.0112813f $X=1.27 $Y=2.56 $X2=0 $Y2=0
cc_169 N_A_57_483#_c_228_n N_VPWR_c_260_n 0.0210042f $X=0.41 $Y=2.56 $X2=0 $Y2=0
cc_170 N_A_57_483#_c_231_n N_Y_c_287_n 0.0211329f $X=1.27 $Y=2.56 $X2=0 $Y2=0
cc_171 N_A_57_483#_c_229_n N_Y_c_285_n 0.00543582f $X=1.14 $Y=2.135 $X2=0 $Y2=0
cc_172 N_A_57_483#_c_231_n N_Y_c_285_n 0.00528749f $X=1.27 $Y=2.56 $X2=0 $Y2=0
cc_173 N_VPWR_c_258_n N_Y_c_288_n 0.0205614f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_174 N_VPWR_c_256_n N_Y_c_288_n 0.011087f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_175 N_Y_c_283_n N_VGND_c_331_n 0.0168955f $X=1.985 $Y=0.882 $X2=0 $Y2=0
cc_176 N_Y_c_282_n N_VGND_c_334_n 0.0126158f $X=1.27 $Y=0.445 $X2=0 $Y2=0
cc_177 Y N_VGND_c_335_n 0.0470144f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_178 N_Y_M1007_d N_VGND_c_336_n 0.0030402f $X=1.13 $Y=0.235 $X2=0 $Y2=0
cc_179 N_Y_M1004_d N_VGND_c_336_n 0.00508616f $X=1.99 $Y=0.235 $X2=0 $Y2=0
cc_180 N_Y_c_282_n N_VGND_c_336_n 0.0095345f $X=1.27 $Y=0.445 $X2=0 $Y2=0
cc_181 N_Y_c_283_n N_VGND_c_336_n 0.0107597f $X=1.985 $Y=0.882 $X2=0 $Y2=0
cc_182 Y N_VGND_c_336_n 0.03106f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_183 N_VGND_c_336_n A_148_47# 0.00328875f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
