* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 a_357_365# a_250_70# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR GATE_N a_250_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VPWR a_789_99# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_567_125# a_250_70# a_639_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_789_99# a_639_125# a_1009_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_1009_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND a_789_99# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 Q a_789_99# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND a_27_468# a_567_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_27_468# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 VPWR a_789_99# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND a_789_99# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_748_447# a_789_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 Q a_789_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 Q a_789_99# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_639_125# a_250_70# a_748_447# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 Q a_789_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_725_125# a_789_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_27_468# a_567_447# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_567_447# a_357_365# a_639_125# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_357_365# a_250_70# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 a_27_468# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VGND GATE_N a_250_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_789_99# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_639_125# a_357_365# a_725_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VPWR a_639_125# a_789_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
