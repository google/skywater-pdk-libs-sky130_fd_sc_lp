* File: sky130_fd_sc_lp__o21bai_1.pxi.spice
* Created: Wed Sep  2 10:17:28 2020
* 
x_PM_SKY130_FD_SC_LP__O21BAI_1%B1_N N_B1_N_M1005_g N_B1_N_c_62_n N_B1_N_c_63_n
+ N_B1_N_c_64_n N_B1_N_M1000_g N_B1_N_c_59_n B1_N B1_N N_B1_N_c_61_n
+ PM_SKY130_FD_SC_LP__O21BAI_1%B1_N
x_PM_SKY130_FD_SC_LP__O21BAI_1%A_27_69# N_A_27_69#_M1005_s N_A_27_69#_M1000_s
+ N_A_27_69#_c_96_n N_A_27_69#_M1006_g N_A_27_69#_M1003_g N_A_27_69#_c_98_n
+ N_A_27_69#_c_99_n N_A_27_69#_c_100_n N_A_27_69#_c_101_n N_A_27_69#_c_102_n
+ N_A_27_69#_c_103_n N_A_27_69#_c_107_n N_A_27_69#_c_104_n N_A_27_69#_c_105_n
+ PM_SKY130_FD_SC_LP__O21BAI_1%A_27_69#
x_PM_SKY130_FD_SC_LP__O21BAI_1%A2 N_A2_M1002_g N_A2_M1007_g A2 A2 N_A2_c_162_n
+ PM_SKY130_FD_SC_LP__O21BAI_1%A2
x_PM_SKY130_FD_SC_LP__O21BAI_1%A1 N_A1_M1004_g N_A1_M1001_g A1 N_A1_c_196_n
+ N_A1_c_197_n PM_SKY130_FD_SC_LP__O21BAI_1%A1
x_PM_SKY130_FD_SC_LP__O21BAI_1%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_c_218_n
+ N_VPWR_c_219_n N_VPWR_c_220_n VPWR N_VPWR_c_221_n N_VPWR_c_222_n
+ N_VPWR_c_223_n N_VPWR_c_217_n PM_SKY130_FD_SC_LP__O21BAI_1%VPWR
x_PM_SKY130_FD_SC_LP__O21BAI_1%Y N_Y_M1006_s N_Y_M1003_d N_Y_c_248_n N_Y_c_249_n
+ N_Y_c_250_n N_Y_c_254_n Y Y Y N_Y_c_273_n PM_SKY130_FD_SC_LP__O21BAI_1%Y
x_PM_SKY130_FD_SC_LP__O21BAI_1%VGND N_VGND_M1005_d N_VGND_M1002_d N_VGND_c_288_n
+ N_VGND_c_289_n VGND N_VGND_c_290_n N_VGND_c_291_n N_VGND_c_292_n
+ N_VGND_c_293_n N_VGND_c_294_n N_VGND_c_295_n PM_SKY130_FD_SC_LP__O21BAI_1%VGND
x_PM_SKY130_FD_SC_LP__O21BAI_1%A_310_47# N_A_310_47#_M1006_d N_A_310_47#_M1004_d
+ N_A_310_47#_c_341_n N_A_310_47#_c_326_n N_A_310_47#_c_327_n
+ N_A_310_47#_c_328_n PM_SKY130_FD_SC_LP__O21BAI_1%A_310_47#
cc_1 VNB N_B1_N_M1005_g 0.0484513f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.555
cc_2 VNB N_B1_N_c_59_n 0.0255561f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.755
cc_3 VNB B1_N 0.0213221f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_N_c_61_n 0.0185474f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_5 VNB N_A_27_69#_c_96_n 0.0202858f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.905
cc_6 VNB N_A_27_69#_M1003_g 0.00843927f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.755
cc_7 VNB N_A_27_69#_c_98_n 0.0647351f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A_27_69#_c_99_n 0.0113633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_69#_c_100_n 0.0186231f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_10 VNB N_A_27_69#_c_101_n 0.0116258f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.295
cc_11 VNB N_A_27_69#_c_102_n 0.00964421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_69#_c_103_n 0.00341776f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.35
cc_13 VNB N_A_27_69#_c_104_n 0.00241694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_69#_c_105_n 0.00247096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_M1002_g 0.0246102f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.555
cc_16 VNB A2 0.00623266f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_17 VNB N_A2_c_162_n 0.0238184f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_A1_M1004_g 0.0289707f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.555
cc_19 VNB N_A1_M1001_g 0.00176104f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.905
cc_20 VNB N_A1_c_196_n 0.0462599f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_A1_c_197_n 0.0112016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_217_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_248_n 0.00695726f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.225
cc_24 VNB N_Y_c_249_n 0.0024809f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.755
cc_25 VNB N_Y_c_250_n 0.00187087f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_26 VNB N_VGND_c_288_n 0.00921285f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.225
cc_27 VNB N_VGND_c_289_n 0.00294193f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_28 VNB N_VGND_c_290_n 0.0166455f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_29 VNB N_VGND_c_291_n 0.0293362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_292_n 0.0174185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_293_n 0.178975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_294_n 0.00596836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_295_n 0.00525267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_310_47#_c_326_n 0.0142202f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.185
cc_35 VNB N_A_310_47#_c_327_n 0.00304301f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.755
cc_36 VNB N_A_310_47#_c_328_n 0.030161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_B1_N_c_62_n 0.0327469f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.83
cc_38 VPB N_B1_N_c_63_n 0.0281749f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.83
cc_39 VPB N_B1_N_c_64_n 0.023865f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=1.905
cc_40 VPB N_B1_N_c_59_n 0.0086463f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.755
cc_41 VPB B1_N 0.014528f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_42 VPB N_A_27_69#_M1003_g 0.0243035f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.755
cc_43 VPB N_A_27_69#_c_107_n 0.0145953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_27_69#_c_104_n 0.00540395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A2_M1007_g 0.0190863f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=1.905
cc_46 VPB A2 0.0111966f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.35
cc_47 VPB N_A2_c_162_n 0.00716793f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_48 VPB N_A1_M1001_g 0.0246229f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=1.905
cc_49 VPB N_A1_c_197_n 0.0067895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_218_n 0.0254691f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.225
cc_51 VPB N_VPWR_c_219_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.185
cc_52 VPB N_VPWR_c_220_n 0.0484246f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_53 VPB N_VPWR_c_221_n 0.0361928f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.35
cc_54 VPB N_VPWR_c_222_n 0.0275337f $X=-0.19 $Y=1.655 $X2=0.3 $Y2=1.665
cc_55 VPB N_VPWR_c_223_n 0.00558929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_217_n 0.0806604f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_249_n 0.00162046f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.755
cc_58 N_B1_N_c_62_n N_A_27_69#_M1003_g 0.0169613f $X=0.875 $Y=1.83 $X2=0 $Y2=0
cc_59 N_B1_N_c_62_n N_A_27_69#_c_98_n 0.01377f $X=0.875 $Y=1.83 $X2=0 $Y2=0
cc_60 B1_N N_A_27_69#_c_98_n 3.16664e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_B1_N_c_61_n N_A_27_69#_c_98_n 0.0173668f $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_62 N_B1_N_M1005_g N_A_27_69#_c_100_n 0.0036463f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_63 N_B1_N_M1005_g N_A_27_69#_c_101_n 0.0157034f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_64 B1_N N_A_27_69#_c_101_n 0.0122793f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_B1_N_c_61_n N_A_27_69#_c_101_n 3.10808e-19 $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_66 B1_N N_A_27_69#_c_102_n 0.0236734f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B1_N_c_61_n N_A_27_69#_c_102_n 0.00104355f $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_68 N_B1_N_M1005_g N_A_27_69#_c_103_n 0.00621279f $X=0.475 $Y=0.555 $X2=0
+ $Y2=0
cc_69 N_B1_N_c_62_n N_A_27_69#_c_107_n 0.00430601f $X=0.875 $Y=1.83 $X2=0 $Y2=0
cc_70 N_B1_N_c_64_n N_A_27_69#_c_107_n 0.00618781f $X=0.95 $Y=1.905 $X2=0 $Y2=0
cc_71 N_B1_N_c_62_n N_A_27_69#_c_104_n 0.0146055f $X=0.875 $Y=1.83 $X2=0 $Y2=0
cc_72 N_B1_N_c_64_n N_A_27_69#_c_104_n 0.00443069f $X=0.95 $Y=1.905 $X2=0 $Y2=0
cc_73 N_B1_N_c_59_n N_A_27_69#_c_104_n 0.0056174f $X=0.385 $Y=1.755 $X2=0 $Y2=0
cc_74 B1_N N_A_27_69#_c_104_n 0.0287162f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_B1_N_c_62_n N_A_27_69#_c_105_n 0.00144349f $X=0.875 $Y=1.83 $X2=0 $Y2=0
cc_76 B1_N N_A_27_69#_c_105_n 0.0268779f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_B1_N_c_61_n N_A_27_69#_c_105_n 0.0021517f $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_78 N_B1_N_c_64_n N_VPWR_c_218_n 0.00466732f $X=0.95 $Y=1.905 $X2=0 $Y2=0
cc_79 N_B1_N_c_64_n N_VPWR_c_221_n 0.00297774f $X=0.95 $Y=1.905 $X2=0 $Y2=0
cc_80 N_B1_N_c_64_n N_VPWR_c_217_n 0.00400849f $X=0.95 $Y=1.905 $X2=0 $Y2=0
cc_81 N_B1_N_M1005_g N_Y_c_248_n 0.00506059f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_82 N_B1_N_c_62_n N_Y_c_249_n 0.00159791f $X=0.875 $Y=1.83 $X2=0 $Y2=0
cc_83 N_B1_N_c_64_n N_Y_c_254_n 0.00155315f $X=0.95 $Y=1.905 $X2=0 $Y2=0
cc_84 N_B1_N_M1005_g N_VGND_c_288_n 0.0134564f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_85 N_B1_N_M1005_g N_VGND_c_290_n 0.00400407f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_86 N_B1_N_M1005_g N_VGND_c_293_n 0.00423498f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_87 N_A_27_69#_c_96_n N_A2_M1002_g 0.0228398f $X=1.475 $Y=1.185 $X2=0 $Y2=0
cc_88 N_A_27_69#_M1003_g N_A2_M1007_g 0.0341139f $X=1.475 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_27_69#_c_99_n A2 0.00319033f $X=1.475 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A_27_69#_c_99_n N_A2_c_162_n 0.0207057f $X=1.475 $Y=1.35 $X2=0 $Y2=0
cc_91 N_A_27_69#_M1003_g N_VPWR_c_218_n 0.0186484f $X=1.475 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A_27_69#_M1003_g N_VPWR_c_222_n 0.00486043f $X=1.475 $Y=2.465 $X2=0
+ $Y2=0
cc_93 N_A_27_69#_M1003_g N_VPWR_c_217_n 0.00870566f $X=1.475 $Y=2.465 $X2=0
+ $Y2=0
cc_94 N_A_27_69#_c_96_n N_Y_c_248_n 0.00874334f $X=1.475 $Y=1.185 $X2=0 $Y2=0
cc_95 N_A_27_69#_c_101_n N_Y_c_248_n 0.0149964f $X=0.685 $Y=0.93 $X2=0 $Y2=0
cc_96 N_A_27_69#_c_96_n N_Y_c_249_n 0.00341979f $X=1.475 $Y=1.185 $X2=0 $Y2=0
cc_97 N_A_27_69#_M1003_g N_Y_c_249_n 0.0112355f $X=1.475 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_27_69#_c_98_n N_Y_c_249_n 0.0168331f $X=1.4 $Y=1.35 $X2=0 $Y2=0
cc_99 N_A_27_69#_c_99_n N_Y_c_249_n 0.00414826f $X=1.475 $Y=1.35 $X2=0 $Y2=0
cc_100 N_A_27_69#_c_103_n N_Y_c_249_n 0.00812764f $X=0.797 $Y=1.185 $X2=0 $Y2=0
cc_101 N_A_27_69#_c_104_n N_Y_c_249_n 0.0188091f $X=0.735 $Y=2.06 $X2=0 $Y2=0
cc_102 N_A_27_69#_c_105_n N_Y_c_249_n 0.0238398f $X=0.955 $Y=1.35 $X2=0 $Y2=0
cc_103 N_A_27_69#_c_96_n N_Y_c_250_n 0.0014982f $X=1.475 $Y=1.185 $X2=0 $Y2=0
cc_104 N_A_27_69#_c_98_n N_Y_c_250_n 0.00706616f $X=1.4 $Y=1.35 $X2=0 $Y2=0
cc_105 N_A_27_69#_M1003_g N_Y_c_254_n 0.00193556f $X=1.475 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_27_69#_c_104_n N_Y_c_254_n 0.00804668f $X=0.735 $Y=2.06 $X2=0 $Y2=0
cc_107 N_A_27_69#_M1003_g Y 0.0165063f $X=1.475 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_27_69#_c_96_n N_VGND_c_288_n 0.00302881f $X=1.475 $Y=1.185 $X2=0
+ $Y2=0
cc_109 N_A_27_69#_c_98_n N_VGND_c_288_n 2.47191e-19 $X=1.4 $Y=1.35 $X2=0 $Y2=0
cc_110 N_A_27_69#_c_101_n N_VGND_c_288_n 0.0245596f $X=0.685 $Y=0.93 $X2=0 $Y2=0
cc_111 N_A_27_69#_c_96_n N_VGND_c_289_n 0.00120547f $X=1.475 $Y=1.185 $X2=0
+ $Y2=0
cc_112 N_A_27_69#_c_100_n N_VGND_c_290_n 0.00959495f $X=0.26 $Y=0.55 $X2=0 $Y2=0
cc_113 N_A_27_69#_c_96_n N_VGND_c_291_n 0.00571722f $X=1.475 $Y=1.185 $X2=0
+ $Y2=0
cc_114 N_A_27_69#_c_96_n N_VGND_c_293_n 0.0118059f $X=1.475 $Y=1.185 $X2=0 $Y2=0
cc_115 N_A_27_69#_c_100_n N_VGND_c_293_n 0.00929928f $X=0.26 $Y=0.55 $X2=0 $Y2=0
cc_116 N_A_27_69#_c_101_n N_VGND_c_293_n 0.00809342f $X=0.685 $Y=0.93 $X2=0
+ $Y2=0
cc_117 N_A_27_69#_c_96_n N_A_310_47#_c_327_n 0.0011462f $X=1.475 $Y=1.185 $X2=0
+ $Y2=0
cc_118 N_A2_M1002_g N_A1_M1004_g 0.0189043f $X=1.91 $Y=0.655 $X2=0 $Y2=0
cc_119 N_A2_M1007_g N_A1_M1001_g 0.0565254f $X=2.045 $Y=2.465 $X2=0 $Y2=0
cc_120 A2 N_A1_c_196_n 0.00273151f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A2_c_162_n N_A1_c_196_n 0.0565254f $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_122 A2 N_A1_c_197_n 0.031643f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A2_c_162_n N_A1_c_197_n 3.09141e-19 $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_124 N_A2_M1007_g N_VPWR_c_218_n 0.00110221f $X=2.045 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A2_M1007_g N_VPWR_c_220_n 0.00451984f $X=2.045 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A2_M1007_g N_VPWR_c_222_n 0.00585385f $X=2.045 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A2_M1007_g N_VPWR_c_217_n 0.0111635f $X=2.045 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A2_M1002_g N_Y_c_249_n 7.70841e-19 $X=1.91 $Y=0.655 $X2=0 $Y2=0
cc_129 N_A2_M1007_g N_Y_c_249_n 8.56942e-19 $X=2.045 $Y=2.465 $X2=0 $Y2=0
cc_130 A2 N_Y_c_249_n 0.0300366f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A2_c_162_n N_Y_c_249_n 3.83119e-19 $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_132 A2 N_Y_c_273_n 0.0266664f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A2_c_162_n N_Y_c_273_n 0.00103656f $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A2_M1002_g N_VGND_c_289_n 0.00999251f $X=1.91 $Y=0.655 $X2=0 $Y2=0
cc_135 N_A2_M1002_g N_VGND_c_291_n 0.00564095f $X=1.91 $Y=0.655 $X2=0 $Y2=0
cc_136 N_A2_M1002_g N_VGND_c_293_n 0.00952034f $X=1.91 $Y=0.655 $X2=0 $Y2=0
cc_137 N_A2_M1002_g N_A_310_47#_c_326_n 0.0143442f $X=1.91 $Y=0.655 $X2=0 $Y2=0
cc_138 A2 N_A_310_47#_c_326_n 0.0337419f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A2_c_162_n N_A_310_47#_c_326_n 0.00426311f $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_140 A2 N_A_310_47#_c_327_n 0.0203237f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_141 N_A2_c_162_n N_A_310_47#_c_327_n 0.0012077f $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_142 N_A1_M1001_g N_VPWR_c_220_n 0.0296373f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A1_c_196_n N_VPWR_c_220_n 0.00146498f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_144 N_A1_c_197_n N_VPWR_c_220_n 0.026128f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_145 N_A1_M1001_g N_VPWR_c_222_n 0.00486043f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A1_M1001_g N_VPWR_c_217_n 0.00818711f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A1_M1004_g N_VGND_c_289_n 0.00327002f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_VGND_c_292_n 0.00585385f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_149 N_A1_M1004_g N_VGND_c_293_n 0.0116566f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_150 N_A1_M1004_g N_A_310_47#_c_326_n 0.018817f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_151 N_A1_c_196_n N_A_310_47#_c_326_n 0.00705552f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_152 N_A1_c_197_n N_A_310_47#_c_326_n 0.0300801f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_153 N_VPWR_c_217_n N_Y_M1003_d 0.00659813f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_154 N_VPWR_M1000_d N_Y_c_249_n 0.00106458f $X=1.025 $Y=2.015 $X2=0 $Y2=0
cc_155 N_VPWR_M1000_d N_Y_c_254_n 0.00314001f $X=1.025 $Y=2.015 $X2=0 $Y2=0
cc_156 N_VPWR_c_218_n N_Y_c_254_n 0.0100034f $X=1.26 $Y=2.38 $X2=0 $Y2=0
cc_157 N_VPWR_c_218_n Y 0.0010324f $X=1.26 $Y=2.38 $X2=0 $Y2=0
cc_158 N_VPWR_c_222_n Y 0.0222962f $X=2.455 $Y=3.33 $X2=0 $Y2=0
cc_159 N_VPWR_c_217_n Y 0.0127519f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_c_217_n A_424_367# 0.00899413f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_161 N_Y_c_248_n N_VGND_c_288_n 0.0287497f $X=1.245 $Y=0.38 $X2=0 $Y2=0
cc_162 N_Y_c_248_n N_VGND_c_291_n 0.0210788f $X=1.245 $Y=0.38 $X2=0 $Y2=0
cc_163 N_Y_M1006_s N_VGND_c_293_n 0.00227725f $X=1.12 $Y=0.235 $X2=0 $Y2=0
cc_164 N_Y_c_248_n N_VGND_c_293_n 0.0126375f $X=1.245 $Y=0.38 $X2=0 $Y2=0
cc_165 N_Y_c_249_n N_A_310_47#_c_327_n 0.0117685f $X=1.325 $Y=1.93 $X2=0 $Y2=0
cc_166 N_VGND_c_293_n N_A_310_47#_M1006_d 0.00418911f $X=2.64 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_167 N_VGND_c_293_n N_A_310_47#_M1004_d 0.00215158f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_168 N_VGND_c_291_n N_A_310_47#_c_341_n 0.0140459f $X=1.98 $Y=0 $X2=0 $Y2=0
cc_169 N_VGND_c_293_n N_A_310_47#_c_341_n 0.00886411f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_170 N_VGND_M1002_d N_A_310_47#_c_326_n 0.00245557f $X=1.985 $Y=0.235 $X2=0
+ $Y2=0
cc_171 N_VGND_c_289_n N_A_310_47#_c_326_n 0.0190564f $X=2.145 $Y=0.38 $X2=0
+ $Y2=0
cc_172 N_VGND_c_292_n N_A_310_47#_c_328_n 0.0194077f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_173 N_VGND_c_293_n N_A_310_47#_c_328_n 0.0117799f $X=2.64 $Y=0 $X2=0 $Y2=0
