* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 a_215_367# a_27_49# a_300_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_49# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_27_49# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR C a_215_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_215_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND a_215_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_372_47# C a_444_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_444_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_215_367# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR a_27_49# a_215_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_300_47# B a_372_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_215_367# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
