* File: sky130_fd_sc_lp__a311oi_lp.pex.spice
* Created: Wed Sep  2 09:25:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311OI_LP%A1 3 5 8 10 11 14 15
c34 14 0 2.52663e-20 $X=0.415 $Y=0.975
r35 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=0.975
+ $X2=0.415 $Y2=1.14
r36 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=0.975
+ $X2=0.415 $Y2=0.81
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=0.975 $X2=0.415 $Y2=0.975
r38 11 15 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.24 $Y=0.975
+ $X2=0.415 $Y2=0.975
r39 10 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.495 $Y=1.9
+ $X2=0.495 $Y2=1.14
r40 8 16 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.505 $Y=0.445
+ $X2=0.505 $Y2=0.81
r41 3 10 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.545 $Y=2.025
+ $X2=0.545 $Y2=1.9
r42 3 5 100.256 $w=2.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.545 $Y=2.025
+ $X2=0.545 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_LP%A2 3 7 9 10 15 16
r48 15 17 4.78808 $w=3.02e-07 $l=3e-08 $layer=POLY_cond $X=1.045 $Y=1.675
+ $X2=1.075 $Y2=1.675
r49 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.045
+ $Y=1.675 $X2=1.045 $Y2=1.675
r50 13 15 23.9404 $w=3.02e-07 $l=1.5e-07 $layer=POLY_cond $X=0.895 $Y=1.675
+ $X2=1.045 $Y2=1.675
r51 10 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.72 $Y=1.675
+ $X2=1.045 $Y2=1.675
r52 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.675
+ $X2=0.72 $Y2=1.675
r53 5 17 7.29241 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.84
+ $X2=1.075 $Y2=1.675
r54 5 7 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.075 $Y=1.84
+ $X2=1.075 $Y2=2.545
r55 1 13 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.51
+ $X2=0.895 $Y2=1.675
r56 1 3 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=0.895 $Y=1.51
+ $X2=0.895 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_LP%A3 3 7 12 15 16 17 21
r44 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.585
+ $Y=1.335 $X2=1.585 $Y2=1.335
r45 17 22 10.1415 $w=3.73e-07 $l=3.3e-07 $layer=LI1_cond $X=1.607 $Y=1.665
+ $X2=1.607 $Y2=1.335
r46 16 22 1.22927 $w=3.73e-07 $l=4e-08 $layer=LI1_cond $X=1.607 $Y=1.295
+ $X2=1.607 $Y2=1.335
r47 14 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.585 $Y=1.675
+ $X2=1.585 $Y2=1.335
r48 14 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.675
+ $X2=1.585 $Y2=1.84
r49 12 21 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=1.585 $Y=1.27
+ $X2=1.585 $Y2=1.335
r50 9 12 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.285 $Y=1.195 $X2=1.585
+ $Y2=1.195
r51 7 15 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.625 $Y=2.545
+ $X2=1.625 $Y2=1.84
r52 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.285 $Y=1.12
+ $X2=1.285 $Y2=1.195
r53 1 3 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.285 $Y=1.12
+ $X2=1.285 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_LP%B1 1 3 4 5 6 8 11 13 16 17 18 19 20 24
c65 24 0 2.87134e-20 $X=2.155 $Y=1.335
r66 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.155 $Y=1.295
+ $X2=2.155 $Y2=1.665
r67 19 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.155
+ $Y=1.335 $X2=2.155 $Y2=1.335
r68 17 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.155 $Y=1.675
+ $X2=2.155 $Y2=1.335
r69 16 24 44.4756 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.17
+ $X2=2.155 $Y2=1.335
r70 11 17 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.84
+ $X2=2.155 $Y2=1.675
r71 11 13 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.155 $Y=1.84
+ $X2=2.155 $Y2=2.545
r72 9 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.075 $Y=0.88
+ $X2=2.075 $Y2=0.805
r73 9 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.075 $Y=0.88
+ $X2=2.075 $Y2=1.17
r74 6 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.075 $Y=0.73
+ $X2=2.075 $Y2=0.805
r75 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.075 $Y=0.73 $X2=2.075
+ $Y2=0.445
r76 4 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2 $Y=0.805 $X2=2.075
+ $Y2=0.805
r77 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2 $Y=0.805 $X2=1.79
+ $Y2=0.805
r78 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.715 $Y=0.73
+ $X2=1.79 $Y2=0.805
r79 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.715 $Y=0.73 $X2=1.715
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_LP%C1 1 3 8 10 11 13 17 19 20 23 24 25
r53 23 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.51
+ $X2=2.725 $Y2=1.675
r54 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.51
+ $X2=2.725 $Y2=1.345
r55 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.725
+ $Y=1.51 $X2=2.725 $Y2=1.51
r56 20 24 4.89394 $w=3.63e-07 $l=1.55e-07 $layer=LI1_cond $X=2.707 $Y=1.665
+ $X2=2.707 $Y2=1.51
r57 19 26 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.635 $Y=1.915
+ $X2=2.635 $Y2=1.675
r58 16 17 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.635 $Y=0.855
+ $X2=2.865 $Y2=0.855
r59 14 16 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=2.505 $Y=0.855
+ $X2=2.635 $Y2=0.855
r60 11 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=0.78
+ $X2=2.865 $Y2=0.855
r61 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.865 $Y=0.78
+ $X2=2.865 $Y2=0.445
r62 8 19 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.685 $Y=2.04
+ $X2=2.685 $Y2=1.915
r63 8 10 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.685 $Y=2.04
+ $X2=2.685 $Y2=2.545
r64 4 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.635 $Y=0.93
+ $X2=2.635 $Y2=0.855
r65 4 25 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=2.635 $Y=0.93
+ $X2=2.635 $Y2=1.345
r66 1 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=0.78
+ $X2=2.505 $Y2=0.855
r67 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.505 $Y=0.78
+ $X2=2.505 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_LP%VPWR 1 2 7 9 13 17 19 26 27 33
r37 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r39 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 23 26 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 21 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.34 $Y2=3.33
r43 21 23 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 19 27 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 19 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 19 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 15 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.34 $Y=3.245
+ $X2=1.34 $Y2=3.33
r48 15 17 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.34 $Y=3.245
+ $X2=1.34 $Y2=2.535
r49 14 30 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r50 13 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=3.33
+ $X2=1.34 $Y2=3.33
r51 13 14 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.175 $Y=3.33
+ $X2=0.445 $Y2=3.33
r52 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.19 $X2=0.28
+ $Y2=2.9
r53 7 30 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r54 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.9
r55 2 17 300 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=2 $X=1.2
+ $Y=2.045 $X2=1.34 $Y2=2.535
r56 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r57 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_LP%A_134_409# 1 2 11 13 14 19
r35 17 19 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.89 $Y=2.19 $X2=1.89
+ $Y2=2.9
r36 13 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.725 $Y=2.105
+ $X2=1.89 $Y2=2.19
r37 13 14 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.725 $Y=2.105
+ $X2=0.975 $Y2=2.105
r38 9 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.81 $Y=2.19
+ $X2=0.975 $Y2=2.105
r39 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.19 $X2=0.81
+ $Y2=2.9
r40 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=2.045 $X2=1.89 $Y2=2.9
r41 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=2.045 $X2=1.89 $Y2=2.19
r42 1 11 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.9
r43 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_LP%Y 1 2 3 10 13 14 15 18 24 29 33 35 36 37
+ 40 42
c87 14 0 2.87134e-20 $X=2.125 $Y=0.905
c88 13 0 2.52663e-20 $X=0.845 $Y=0.82
r89 37 42 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=3.12 $Y=0.925
+ $X2=3.155 $Y2=0.925
r90 37 40 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=0.925
+ $X2=3.005 $Y2=0.925
r91 35 36 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.012 $Y=2.19
+ $X2=3.012 $Y2=2.025
r92 29 31 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.29 $Y=0.445 $X2=0.29
+ $Y2=0.545
r93 26 42 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.155 $Y=1.04
+ $X2=3.155 $Y2=0.925
r94 26 36 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=3.155 $Y=1.04
+ $X2=3.155 $Y2=2.025
r95 22 35 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=3.012 $Y=2.252
+ $X2=3.012 $Y2=2.19
r96 22 24 17.0343 $w=4.53e-07 $l=6.48e-07 $layer=LI1_cond $X=3.012 $Y=2.252
+ $X2=3.012 $Y2=2.9
r97 21 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0.905
+ $X2=2.29 $Y2=0.905
r98 21 40 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.455 $Y=0.905
+ $X2=3.005 $Y2=0.905
r99 16 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.82 $X2=2.29
+ $Y2=0.905
r100 16 18 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.29 $Y=0.82
+ $X2=2.29 $Y2=0.47
r101 14 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0.905
+ $X2=2.29 $Y2=0.905
r102 14 15 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=2.125 $Y=0.905
+ $X2=0.93 $Y2=0.905
r103 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.845 $Y=0.82
+ $X2=0.93 $Y2=0.905
r104 12 13 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.845 $Y=0.63
+ $X2=0.845 $Y2=0.82
r105 11 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=0.545
+ $X2=0.29 $Y2=0.545
r106 10 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.76 $Y=0.545
+ $X2=0.845 $Y2=0.63
r107 10 11 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.76 $Y=0.545
+ $X2=0.455 $Y2=0.545
r108 3 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.045 $X2=2.95 $Y2=2.19
r109 3 24 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.045 $X2=2.95 $Y2=2.9
r110 2 18 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.15
+ $Y=0.235 $X2=2.29 $Y2=0.47
r111 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.235 $X2=0.29 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_LP%VGND 1 2 9 11 13 16 17 18 27 36
r54 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r55 33 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r56 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r57 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r58 27 35 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r59 27 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r60 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r61 22 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r62 21 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r63 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r64 18 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r65 18 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r66 18 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r67 16 25 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.2
+ $Y2=0
r68 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.5
+ $Y2=0
r69 15 29 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.665 $Y=0 $X2=1.68
+ $Y2=0
r70 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=0 $X2=1.5
+ $Y2=0
r71 11 35 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r72 11 13 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.42
r73 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=0.085 $X2=1.5
+ $Y2=0
r74 7 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.5 $Y=0.085 $X2=1.5
+ $Y2=0.425
r75 2 13 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.42
r76 1 9 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.36
+ $Y=0.235 $X2=1.5 $Y2=0.425
.ends

