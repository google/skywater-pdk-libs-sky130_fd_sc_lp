* File: sky130_fd_sc_lp__o31a_1.pex.spice
* Created: Wed Sep  2 10:24:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31A_1%A_86_23# 1 2 9 12 16 17 19 20 23 25 29 32 34
+ 35 37
c69 16 0 8.21982e-20 $X=0.64 $Y=1.36
r70 32 35 50.8333 $w=1.78e-07 $l=8.25e-07 $layer=LI1_cond $X=3.185 $Y=1.93
+ $X2=3.185 $Y2=1.105
r71 27 35 10.429 $w=4.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.05 $Y=0.88
+ $X2=3.05 $Y2=1.105
r72 27 29 12.2266 $w=4.48e-07 $l=4.6e-07 $layer=LI1_cond $X=3.05 $Y=0.88
+ $X2=3.05 $Y2=0.42
r73 26 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=2.015
+ $X2=2.455 $Y2=2.015
r74 25 32 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.095 $Y=2.015
+ $X2=3.185 $Y2=1.93
r75 25 26 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.095 $Y=2.015
+ $X2=2.62 $Y2=2.015
r76 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=2.1
+ $X2=2.455 $Y2=2.015
r77 21 23 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.455 $Y=2.1
+ $X2=2.455 $Y2=2.485
r78 19 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=2.015
+ $X2=2.455 $Y2=2.015
r79 19 20 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=2.29 $Y=2.015
+ $X2=0.805 $Y2=2.015
r80 17 38 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.617 $Y=1.36
+ $X2=0.617 $Y2=1.525
r81 17 37 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.617 $Y=1.36
+ $X2=0.617 $Y2=1.195
r82 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.36 $X2=0.64 $Y2=1.36
r83 14 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.68 $Y=1.93
+ $X2=0.805 $Y2=2.015
r84 14 16 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=0.68 $Y=1.93
+ $X2=0.68 $Y2=1.36
r85 12 38 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=0.505 $Y=2.465 $X2=0.505
+ $Y2=1.525
r86 9 37 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.505 $Y=0.665
+ $X2=0.505 $Y2=1.195
r87 2 34 600 $w=1.7e-07 $l=2.54558e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.835 $X2=2.455 $Y2=2.015
r88 2 23 300 $w=1.7e-07 $l=7.34507e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=1.835 $X2=2.455 $Y2=2.485
r89 1 29 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.815
+ $Y=0.245 $X2=2.955 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_1%A1 3 6 8 9 13 15
c36 15 0 8.21982e-20 $X=1.205 $Y=1.21
c37 8 0 6.86178e-20 $X=1.2 $Y=1.295
r38 13 16 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.205 $Y=1.375
+ $X2=1.205 $Y2=1.54
r39 13 15 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.205 $Y=1.375
+ $X2=1.205 $Y2=1.21
r40 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.16 $Y=1.295 $X2=1.16
+ $Y2=1.665
r41 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.375 $X2=1.2 $Y2=1.375
r42 6 16 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.3 $Y=2.465 $X2=1.3
+ $Y2=1.54
r43 3 15 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.3 $Y=0.665 $X2=1.3
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_1%A2 3 7 9 12 13
c38 7 0 6.86178e-20 $X=1.76 $Y=2.465
r39 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.51
+ $X2=1.75 $Y2=1.675
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.51
+ $X2=1.75 $Y2=1.345
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.51 $X2=1.75 $Y2=1.51
r42 9 13 5.3322 $w=3.33e-07 $l=1.55e-07 $layer=LI1_cond $X=1.667 $Y=1.665
+ $X2=1.667 $Y2=1.51
r43 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.76 $Y=2.465
+ $X2=1.76 $Y2=1.675
r44 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.755 $Y=0.665
+ $X2=1.755 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_1%A3 3 7 9 12 13
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.51
+ $X2=2.29 $Y2=1.675
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.51
+ $X2=2.29 $Y2=1.345
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.51 $X2=2.29 $Y2=1.51
r39 9 13 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.19 $Y=1.665
+ $X2=2.19 $Y2=1.51
r40 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.31 $Y=0.665
+ $X2=2.31 $Y2=1.345
r41 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.2 $Y=2.465 $X2=2.2
+ $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_1%B1 3 7 9 12 13
r32 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.51
+ $X2=2.83 $Y2=1.675
r33 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.51
+ $X2=2.83 $Y2=1.345
r34 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.83
+ $Y=1.51 $X2=2.83 $Y2=1.51
r35 9 13 5.27625 $w=4.13e-07 $l=1.9e-07 $layer=LI1_cond $X=2.64 $Y=1.552
+ $X2=2.83 $Y2=1.552
r36 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.74 $Y=2.465
+ $X2=2.74 $Y2=1.675
r37 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.74 $Y=0.665
+ $X2=2.74 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_1%X 1 2 7 8 9 10 11 12 13 22
r10 13 40 5.18599 $w=2.98e-07 $l=1.35e-07 $layer=LI1_cond $X=0.235 $Y=2.775
+ $X2=0.235 $Y2=2.91
r11 12 13 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=2.405
+ $X2=0.235 $Y2=2.775
r12 11 12 16.3263 $w=2.98e-07 $l=4.25e-07 $layer=LI1_cond $X=0.235 $Y=1.98
+ $X2=0.235 $Y2=2.405
r13 10 11 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=0.235 $Y=1.665
+ $X2=0.235 $Y2=1.98
r14 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.665
r15 8 9 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=0.925
+ $X2=0.235 $Y2=1.295
r16 7 8 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=0.555
+ $X2=0.235 $Y2=0.925
r17 7 22 5.18599 $w=2.98e-07 $l=1.35e-07 $layer=LI1_cond $X=0.235 $Y=0.555
+ $X2=0.235 $Y2=0.42
r18 2 40 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.91
r19 2 11 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=1.98
r20 1 22 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.245 $X2=0.29 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_1%VPWR 1 2 9 11 13 15 17 22 28 34
r38 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 29 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 28 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 23 28 13.6095 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=0.902 $Y2=3.33
r45 23 25 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 22 33 4.51706 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.79 $Y=3.33
+ $X2=3.075 $Y2=3.33
r47 22 25 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=3.33 $X2=2.64
+ $Y2=3.33
r48 20 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 17 28 13.6095 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.902 $Y2=3.33
r51 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 15 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 11 33 3.24911 $w=3.3e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=3.075 $Y2=3.33
r55 11 13 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=2.955 $Y2=2.385
r56 7 28 2.84707 $w=6.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.902 $Y=3.245
+ $X2=0.902 $Y2=3.33
r57 7 9 15.3167 $w=6.93e-07 $l=8.9e-07 $layer=LI1_cond $X=0.902 $Y=3.245
+ $X2=0.902 $Y2=2.355
r58 2 13 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=2.815
+ $Y=1.835 $X2=2.955 $Y2=2.385
r59 1 9 150 $w=1.7e-07 $l=7.30068e-07 $layer=licon1_PDIFF $count=4 $X=0.58
+ $Y=1.835 $X2=1.085 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r43 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r46 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.2 $Y=0 $X2=2.035
+ $Y2=0
r48 27 29 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.2 $Y=0 $X2=3.12
+ $Y2=0
r49 23 33 13.6095 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=0.902
+ $Y2=0
r50 23 25 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.68
+ $Y2=0
r51 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=2.035
+ $Y2=0
r52 22 25 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.68
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 13.6095 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.902
+ $Y2=0
r56 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.24
+ $Y2=0
r57 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r58 15 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r59 15 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=0.085
+ $X2=2.035 $Y2=0
r61 11 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.035 $Y=0.085
+ $X2=2.035 $Y2=0.37
r62 7 33 2.84707 $w=6.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.902 $Y=0.085
+ $X2=0.902 $Y2=0
r63 7 9 5.24898 $w=6.93e-07 $l=3.05e-07 $layer=LI1_cond $X=0.902 $Y=0.085
+ $X2=0.902 $Y2=0.39
r64 2 13 91 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=2 $X=1.83
+ $Y=0.245 $X2=2.035 $Y2=0.37
r65 1 9 45.5 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_NDIFF $count=4 $X=0.58
+ $Y=0.245 $X2=1.085 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_1%A_275_49# 1 2 9 11 12 15
r31 13 15 23.6554 $w=2.83e-07 $l=5.85e-07 $layer=LI1_cond $X=2.512 $Y=1.005
+ $X2=2.512 $Y2=0.42
r32 11 13 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=2.37 $Y=1.09
+ $X2=2.512 $Y2=1.005
r33 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.37 $Y=1.09 $X2=1.7
+ $Y2=1.09
r34 7 12 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=1.577 $Y=1.005
+ $X2=1.7 $Y2=1.09
r35 7 9 27.5175 $w=2.43e-07 $l=5.85e-07 $layer=LI1_cond $X=1.577 $Y=1.005
+ $X2=1.577 $Y2=0.42
r36 2 15 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.385
+ $Y=0.245 $X2=2.525 $Y2=0.42
r37 1 9 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=1.375
+ $Y=0.245 $X2=1.54 $Y2=0.42
.ends

