* File: sky130_fd_sc_lp__nand2b_lp.pex.spice
* Created: Wed Sep  2 10:03:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2B_LP%A_N 1 3 7 10 12 14 16 17 18 19 22 23 24
c49 10 0 2.56727e-20 $X=0.69 $Y=2.595
r50 22 24 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.39
+ $X2=0.63 $Y2=1.225
r51 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.65
+ $Y=1.39 $X2=0.65 $Y2=1.39
r52 19 23 9.05491 $w=3.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.66 $Y=1.665
+ $X2=0.66 $Y2=1.39
r53 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.88 $Y=0.75 $X2=0.88
+ $Y2=0.465
r54 13 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.595 $Y=0.825
+ $X2=0.52 $Y2=0.825
r55 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.805 $Y=0.825
+ $X2=0.88 $Y2=0.75
r56 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.805 $Y=0.825
+ $X2=0.595 $Y2=0.825
r57 10 18 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.69 $Y=2.595 $X2=0.69
+ $Y2=1.895
r58 7 18 34.9505 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=0.63 $Y=1.71
+ $X2=0.63 $Y2=1.895
r59 6 22 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=0.63 $Y=1.41 $X2=0.63
+ $Y2=1.39
r60 6 7 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=0.63 $Y=1.41 $X2=0.63
+ $Y2=1.71
r61 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.9 $X2=0.52
+ $Y2=0.825
r62 4 24 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.52 $Y=0.9 $X2=0.52
+ $Y2=1.225
r63 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.75 $X2=0.52
+ $Y2=0.825
r64 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.75 $X2=0.52
+ $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_LP%B 1 3 7 11 12 15 16
r42 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.22
+ $Y=1.39 $X2=1.22 $Y2=1.39
r43 12 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.39
r44 11 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.22 $Y=1.73
+ $X2=1.22 $Y2=1.39
r45 10 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.225
+ $X2=1.22 $Y2=1.39
r46 7 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.31 $Y=0.465
+ $X2=1.31 $Y2=1.225
r47 1 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.895
+ $X2=1.22 $Y2=1.73
r48 1 3 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.22 $Y=1.895 $X2=1.22
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_LP%A_32_51# 1 2 9 13 17 18 21 27 31 33 34 36
+ 37
r70 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.79
+ $Y=1.04 $X2=1.79 $Y2=1.04
r71 33 34 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.362 $Y=2.24
+ $X2=0.362 $Y2=2.075
r72 28 31 2.79892 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.47 $Y=0.96
+ $X2=0.302 $Y2=0.96
r73 27 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=0.96
+ $X2=1.79 $Y2=0.96
r74 27 28 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.625 $Y=0.96
+ $X2=0.47 $Y2=0.96
r75 23 31 3.67481 $w=2.52e-07 $l=1.19143e-07 $layer=LI1_cond $X=0.22 $Y=1.045
+ $X2=0.302 $Y2=0.96
r76 23 34 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.22 $Y=1.045
+ $X2=0.22 $Y2=2.075
r77 19 31 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=0.302 $Y=0.875
+ $X2=0.302 $Y2=0.96
r78 19 21 13.5885 $w=3.33e-07 $l=3.95e-07 $layer=LI1_cond $X=0.302 $Y=0.875
+ $X2=0.302 $Y2=0.48
r79 17 37 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.79 $Y=1.38
+ $X2=1.79 $Y2=1.04
r80 17 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.38
+ $X2=1.79 $Y2=1.545
r81 16 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=0.875
+ $X2=1.79 $Y2=1.04
r82 13 18 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.75 $Y=2.595
+ $X2=1.75 $Y2=1.545
r83 9 16 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.7 $Y=0.465 $X2=1.7
+ $Y2=0.875
r84 2 33 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=2.095 $X2=0.425 $Y2=2.24
r85 1 21 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.255 $X2=0.305 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_LP%VPWR 1 2 9 13 15 18 19 20 26 32
r34 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 29 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 26 31 4.65202 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=2.157 $Y2=3.33
r38 26 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 20 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 18 23 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.79 $Y=3.33 $X2=0.72
+ $Y2=3.33
r43 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=3.33
+ $X2=0.955 $Y2=3.33
r44 17 28 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.12 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=3.33
+ $X2=0.955 $Y2=3.33
r46 13 31 3.11416 $w=3.3e-07 $l=1.17346e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.157 $Y2=3.33
r47 13 15 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=2.495
r48 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.955 $Y=2.24
+ $X2=0.955 $Y2=2.95
r49 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=3.245
+ $X2=0.955 $Y2=3.33
r50 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.955 $Y=3.245
+ $X2=0.955 $Y2=2.95
r51 2 15 300 $w=1.7e-07 $l=4.91935e-07 $layer=licon1_PDIFF $count=2 $X=1.875
+ $Y=2.095 $X2=2.08 $Y2=2.495
r52 1 12 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.815
+ $Y=2.095 $X2=0.955 $Y2=2.95
r53 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.815
+ $Y=2.095 $X2=0.955 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_LP%Y 1 2 7 9 12 16 18 19 24
c36 7 0 2.56727e-20 $X=1.527 $Y=2.15
r37 19 24 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=2.035
+ $X2=2.135 $Y2=2.035
r38 19 24 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=2.135 $Y2=2.035
r39 18 25 4.87637 $w=2.3e-07 $l=2.08e-07 $layer=LI1_cond $X=1.527 $Y=2.035
+ $X2=1.735 $Y2=2.035
r40 18 19 17.7877 $w=2.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.75 $Y=2.035
+ $X2=2.105 $Y2=2.035
r41 18 25 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.75 $Y=2.035
+ $X2=1.735 $Y2=2.035
r42 14 16 8.1743 $w=4.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.915 $Y=0.48
+ $X2=2.22 $Y2=0.48
r43 12 19 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.22 $Y=1.92
+ $X2=2.22 $Y2=2.035
r44 11 16 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.22 $Y=0.695
+ $X2=2.22 $Y2=0.48
r45 11 12 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=2.22 $Y=0.695
+ $X2=2.22 $Y2=1.92
r46 7 18 2.69607 $w=4.15e-07 $l=1.15e-07 $layer=LI1_cond $X=1.527 $Y=2.15
+ $X2=1.527 $Y2=2.035
r47 7 9 2.49927 $w=4.13e-07 $l=9e-08 $layer=LI1_cond $X=1.527 $Y=2.15 $X2=1.527
+ $Y2=2.24
r48 2 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.345
+ $Y=2.095 $X2=1.485 $Y2=2.24
r49 1 14 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.255 $X2=1.915 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_LP%VGND 1 6 8 10 17 18 21
r26 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.095
+ $Y2=0
r28 15 17 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=2.16
+ $Y2=0
r29 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=1.095
+ $Y2=0
r31 10 12 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=0.72
+ $Y2=0
r32 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r33 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r34 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=0.085
+ $X2=1.095 $Y2=0
r36 4 6 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.095 $Y=0.085
+ $X2=1.095 $Y2=0.465
r37 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.955
+ $Y=0.255 $X2=1.095 $Y2=0.465
.ends

