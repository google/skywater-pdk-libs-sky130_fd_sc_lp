* File: sky130_fd_sc_lp__dfrbp_lp.pxi.spice
* Created: Fri Aug 28 10:21:56 2020
* 
x_PM_SKY130_FD_SC_LP__DFRBP_LP%D N_D_M1043_g N_D_c_335_n N_D_c_336_n N_D_M1012_g
+ N_D_M1023_g N_D_c_329_n N_D_c_330_n N_D_c_331_n D D D N_D_c_333_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%D
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_662_90# N_A_662_90#_M1041_d N_A_662_90#_M1047_d
+ N_A_662_90#_c_392_n N_A_662_90#_M1045_g N_A_662_90#_M1010_g
+ N_A_662_90#_c_394_n N_A_662_90#_M1019_g N_A_662_90#_c_396_n
+ N_A_662_90#_c_397_n N_A_662_90#_M1021_g N_A_662_90#_c_398_n
+ N_A_662_90#_c_399_n N_A_662_90#_c_400_n N_A_662_90#_c_447_p
+ N_A_662_90#_c_401_n N_A_662_90#_c_402_n N_A_662_90#_c_403_n
+ N_A_662_90#_c_404_n N_A_662_90#_c_405_n N_A_662_90#_c_406_n
+ N_A_662_90#_c_407_n N_A_662_90#_c_408_n N_A_662_90#_c_409_n
+ N_A_662_90#_c_410_n N_A_662_90#_c_411_n PM_SKY130_FD_SC_LP__DFRBP_LP%A_662_90#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_817_90# N_A_817_90#_M1004_s N_A_817_90#_M1021_s
+ N_A_817_90#_M1000_s N_A_817_90#_M1044_d N_A_817_90#_M1003_g
+ N_A_817_90#_c_566_n N_A_817_90#_M1002_g N_A_817_90#_c_559_n
+ N_A_817_90#_c_560_n N_A_817_90#_c_561_n N_A_817_90#_c_569_n
+ N_A_817_90#_c_570_n N_A_817_90#_c_562_n N_A_817_90#_c_572_n
+ N_A_817_90#_c_573_n N_A_817_90#_c_563_n N_A_817_90#_c_575_n
+ N_A_817_90#_c_564_n N_A_817_90#_c_576_n N_A_817_90#_c_577_n
+ N_A_817_90#_c_578_n N_A_817_90#_c_579_n N_A_817_90#_c_565_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%A_817_90#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%RESET_B N_RESET_B_c_722_n N_RESET_B_M1014_g
+ N_RESET_B_M1022_g N_RESET_B_c_723_n N_RESET_B_c_724_n N_RESET_B_M1033_g
+ N_RESET_B_c_726_n N_RESET_B_c_727_n N_RESET_B_M1040_g N_RESET_B_c_729_n
+ N_RESET_B_c_730_n N_RESET_B_c_750_n N_RESET_B_M1009_g N_RESET_B_c_751_n
+ N_RESET_B_M1038_g N_RESET_B_c_731_n N_RESET_B_M1017_g N_RESET_B_M1029_g
+ N_RESET_B_M1001_g N_RESET_B_c_733_n N_RESET_B_c_734_n N_RESET_B_c_735_n
+ N_RESET_B_c_736_n N_RESET_B_c_737_n N_RESET_B_c_738_n N_RESET_B_c_739_n
+ N_RESET_B_c_740_n RESET_B N_RESET_B_c_742_n N_RESET_B_c_743_n
+ N_RESET_B_c_744_n N_RESET_B_c_745_n N_RESET_B_c_746_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%RESET_B
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_590_116# N_A_590_116#_M1016_d
+ N_A_590_116#_M1024_d N_A_590_116#_M1038_d N_A_590_116#_c_971_n
+ N_A_590_116#_c_972_n N_A_590_116#_c_973_n N_A_590_116#_M1004_g
+ N_A_590_116#_M1000_g N_A_590_116#_c_975_n N_A_590_116#_c_976_n
+ N_A_590_116#_M1005_g N_A_590_116#_M1007_g N_A_590_116#_c_978_n
+ N_A_590_116#_c_979_n N_A_590_116#_c_980_n N_A_590_116#_c_990_n
+ N_A_590_116#_c_991_n N_A_590_116#_c_981_n N_A_590_116#_c_993_n
+ N_A_590_116#_c_982_n N_A_590_116#_c_983_n N_A_590_116#_c_1056_n
+ N_A_590_116#_c_994_n N_A_590_116#_c_984_n N_A_590_116#_c_995_n
+ N_A_590_116#_c_996_n N_A_590_116#_c_997_n N_A_590_116#_c_985_n
+ N_A_590_116#_c_986_n PM_SKY130_FD_SC_LP__DFRBP_LP%A_590_116#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_560_90# N_A_560_90#_M1026_s N_A_560_90#_M1049_s
+ N_A_560_90#_M1016_g N_A_560_90#_M1024_g N_A_560_90#_c_1168_n
+ N_A_560_90#_c_1169_n N_A_560_90#_M1039_g N_A_560_90#_M1006_g
+ N_A_560_90#_c_1171_n N_A_560_90#_M1047_g N_A_560_90#_M1041_g
+ N_A_560_90#_c_1173_n N_A_560_90#_M1044_g N_A_560_90#_c_1153_n
+ N_A_560_90#_c_1154_n N_A_560_90#_M1036_g N_A_560_90#_c_1175_n
+ N_A_560_90#_c_1156_n N_A_560_90#_c_1177_n N_A_560_90#_c_1178_n
+ N_A_560_90#_c_1157_n N_A_560_90#_c_1158_n N_A_560_90#_c_1159_n
+ N_A_560_90#_c_1160_n N_A_560_90#_c_1246_p N_A_560_90#_c_1161_n
+ N_A_560_90#_c_1356_p N_A_560_90#_c_1162_n N_A_560_90#_c_1179_n
+ N_A_560_90#_c_1163_n N_A_560_90#_c_1164_n N_A_560_90#_c_1266_p
+ N_A_560_90#_c_1180_n N_A_560_90#_c_1165_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%A_560_90#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_2102_25# N_A_2102_25#_M1030_d
+ N_A_2102_25#_M1008_d N_A_2102_25#_M1032_g N_A_2102_25#_M1013_g
+ N_A_2102_25#_c_1392_n N_A_2102_25#_c_1393_n N_A_2102_25#_c_1394_n
+ N_A_2102_25#_c_1395_n N_A_2102_25#_c_1396_n N_A_2102_25#_c_1397_n
+ N_A_2102_25#_c_1398_n N_A_2102_25#_c_1399_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%A_2102_25#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_1799_379# N_A_1799_379#_M1021_d
+ N_A_1799_379#_M1019_d N_A_1799_379#_M1008_g N_A_1799_379#_M1030_g
+ N_A_1799_379#_c_1467_n N_A_1799_379#_c_1468_n N_A_1799_379#_M1020_g
+ N_A_1799_379#_M1050_g N_A_1799_379#_M1031_g N_A_1799_379#_c_1470_n
+ N_A_1799_379#_M1035_g N_A_1799_379#_M1011_g N_A_1799_379#_c_1473_n
+ N_A_1799_379#_M1042_g N_A_1799_379#_M1028_g N_A_1799_379#_c_1476_n
+ N_A_1799_379#_M1048_g N_A_1799_379#_M1025_g N_A_1799_379#_c_1479_n
+ N_A_1799_379#_c_1480_n N_A_1799_379#_c_1481_n N_A_1799_379#_c_1500_n
+ N_A_1799_379#_c_1482_n N_A_1799_379#_c_1483_n N_A_1799_379#_c_1502_n
+ N_A_1799_379#_c_1503_n N_A_1799_379#_c_1504_n N_A_1799_379#_c_1505_n
+ N_A_1799_379#_c_1506_n N_A_1799_379#_c_1507_n N_A_1799_379#_c_1508_n
+ N_A_1799_379#_c_1509_n N_A_1799_379#_c_1484_n N_A_1799_379#_c_1511_n
+ N_A_1799_379#_c_1485_n N_A_1799_379#_c_1486_n N_A_1799_379#_c_1487_n
+ N_A_1799_379#_c_1488_n N_A_1799_379#_c_1489_n N_A_1799_379#_c_1490_n
+ N_A_1799_379#_c_1491_n N_A_1799_379#_c_1492_n N_A_1799_379#_c_1493_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%A_1799_379#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%CLK N_CLK_M1026_g N_CLK_M1049_g N_CLK_c_1717_n
+ N_CLK_M1027_g N_CLK_M1034_g N_CLK_c_1720_n CLK CLK N_CLK_c_1722_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%CLK
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_3222_137# N_A_3222_137#_M1042_s
+ N_A_3222_137#_M1028_s N_A_3222_137#_M1015_g N_A_3222_137#_M1037_g
+ N_A_3222_137#_M1018_g N_A_3222_137#_M1046_g N_A_3222_137#_c_1776_n
+ N_A_3222_137#_c_1782_n N_A_3222_137#_c_1777_n N_A_3222_137#_c_1778_n
+ N_A_3222_137#_c_1779_n PM_SKY130_FD_SC_LP__DFRBP_LP%A_3222_137#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_27_457# N_A_27_457#_M1043_s N_A_27_457#_M1012_d
+ N_A_27_457#_c_1834_n N_A_27_457#_c_1835_n N_A_27_457#_c_1836_n
+ N_A_27_457#_c_1837_n N_A_27_457#_c_1838_n N_A_27_457#_c_1853_n
+ N_A_27_457#_c_1839_n PM_SKY130_FD_SC_LP__DFRBP_LP%A_27_457#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_111_457# N_A_111_457#_M1023_d
+ N_A_111_457#_M1043_d N_A_111_457#_M1010_d N_A_111_457#_c_1876_n
+ N_A_111_457#_c_1877_n N_A_111_457#_c_1878_n N_A_111_457#_c_1875_n
+ N_A_111_457#_c_1880_n N_A_111_457#_c_1881_n N_A_111_457#_c_1882_n
+ N_A_111_457#_c_1883_n N_A_111_457#_c_1884_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%A_111_457#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%VPWR N_VPWR_M1022_d N_VPWR_M1002_d N_VPWR_M1007_d
+ N_VPWR_M1013_d N_VPWR_M1001_d N_VPWR_M1034_d N_VPWR_M1025_d N_VPWR_c_1951_n
+ N_VPWR_c_1952_n N_VPWR_c_1953_n N_VPWR_c_1954_n N_VPWR_c_1955_n
+ N_VPWR_c_1956_n N_VPWR_c_1957_n N_VPWR_c_1958_n N_VPWR_c_1959_n
+ N_VPWR_c_1960_n N_VPWR_c_1961_n N_VPWR_c_1962_n N_VPWR_c_1963_n VPWR
+ N_VPWR_c_1964_n N_VPWR_c_1965_n N_VPWR_c_1966_n N_VPWR_c_1967_n
+ N_VPWR_c_1968_n N_VPWR_c_1950_n N_VPWR_c_1970_n N_VPWR_c_1971_n
+ N_VPWR_c_1972_n N_VPWR_c_1973_n PM_SKY130_FD_SC_LP__DFRBP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_484_411# N_A_484_411#_M1024_s
+ N_A_484_411#_M1002_s N_A_484_411#_c_2103_n N_A_484_411#_c_2104_n
+ N_A_484_411#_c_2105_n N_A_484_411#_c_2106_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%A_484_411#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_1712_379# N_A_1712_379#_M1019_s
+ N_A_1712_379#_M1013_s N_A_1712_379#_c_2146_n N_A_1712_379#_c_2147_n
+ N_A_1712_379#_c_2148_n N_A_1712_379#_c_2149_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%A_1712_379#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%A_2185_397# N_A_2185_397#_M1008_s
+ N_A_2185_397#_M1020_d N_A_2185_397#_c_2173_n N_A_2185_397#_c_2174_n
+ N_A_2185_397#_c_2175_n N_A_2185_397#_c_2176_n N_A_2185_397#_c_2177_n
+ N_A_2185_397#_c_2178_n N_A_2185_397#_c_2179_n N_A_2185_397#_c_2180_n
+ PM_SKY130_FD_SC_LP__DFRBP_LP%A_2185_397#
x_PM_SKY130_FD_SC_LP__DFRBP_LP%Q_N N_Q_N_M1035_d N_Q_N_M1011_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_2228_n PM_SKY130_FD_SC_LP__DFRBP_LP%Q_N
x_PM_SKY130_FD_SC_LP__DFRBP_LP%Q N_Q_M1018_d N_Q_M1046_d Q Q Q Q Q Q Q
+ N_Q_c_2251_n PM_SKY130_FD_SC_LP__DFRBP_LP%Q
x_PM_SKY130_FD_SC_LP__DFRBP_LP%VGND N_VGND_M1033_s N_VGND_M1040_d N_VGND_M1005_d
+ N_VGND_M1032_d N_VGND_M1027_d N_VGND_M1048_d N_VGND_c_2266_n N_VGND_c_2267_n
+ N_VGND_c_2268_n N_VGND_c_2269_n N_VGND_c_2270_n N_VGND_c_2271_n
+ N_VGND_c_2272_n VGND N_VGND_c_2273_n N_VGND_c_2274_n N_VGND_c_2275_n
+ N_VGND_c_2276_n N_VGND_c_2277_n N_VGND_c_2278_n N_VGND_c_2279_n
+ N_VGND_c_2280_n N_VGND_c_2281_n N_VGND_c_2282_n N_VGND_c_2283_n
+ N_VGND_c_2284_n N_VGND_c_2285_n PM_SKY130_FD_SC_LP__DFRBP_LP%VGND
cc_1 VNB N_D_M1012_g 0.00228913f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.68
cc_2 VNB N_D_c_329_n 0.0371067f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.47
cc_3 VNB N_D_c_330_n 0.0170688f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.24
cc_4 VNB N_D_c_331_n 0.0117934f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.075
cc_5 VNB D 0.0179831f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_6 VNB N_D_c_333_n 0.0189516f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.295
cc_7 VNB N_A_662_90#_c_392_n 0.0157877f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.62
cc_8 VNB N_A_662_90#_M1010_g 0.0130302f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.79
cc_9 VNB N_A_662_90#_c_394_n 0.093829f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.545
cc_10 VNB N_A_662_90#_M1019_g 0.0226994f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.545
cc_11 VNB N_A_662_90#_c_396_n 0.0299766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_662_90#_c_397_n 0.0206542f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.075
cc_13 VNB N_A_662_90#_c_398_n 0.00375964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_662_90#_c_399_n 0.0584096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_662_90#_c_400_n 0.0083081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_662_90#_c_401_n 0.0138475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_662_90#_c_402_n 0.0224935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_662_90#_c_403_n 0.00365429f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.295
cc_19 VNB N_A_662_90#_c_404_n 7.30072e-19 $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.295
cc_20 VNB N_A_662_90#_c_405_n 0.019756f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.555
cc_21 VNB N_A_662_90#_c_406_n 0.00277163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_662_90#_c_407_n 0.0128663f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.925
cc_23 VNB N_A_662_90#_c_408_n 0.00113092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_662_90#_c_409_n 0.0147784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_662_90#_c_410_n 0.00455983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_662_90#_c_411_n 0.00156651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_817_90#_M1003_g 0.0348439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_817_90#_c_559_n 0.0334112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_817_90#_c_560_n 0.00244282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_817_90#_c_561_n 0.00397298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_817_90#_c_562_n 0.0156172f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.555
cc_32 VNB N_A_817_90#_c_563_n 0.00354554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_817_90#_c_564_n 0.0217067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_817_90#_c_565_n 0.00100498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_RESET_B_c_722_n 0.0164148f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=3.075
cc_36 VNB N_RESET_B_c_723_n 0.0307487f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.68
cc_37 VNB N_RESET_B_c_724_n 0.0350471f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.68
cc_38 VNB N_RESET_B_M1033_g 0.0308527f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.545
cc_39 VNB N_RESET_B_c_726_n 0.220628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_RESET_B_c_727_n 0.0125935f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.545
cc_41 VNB N_RESET_B_M1040_g 0.0305854f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.075
cc_42 VNB N_RESET_B_c_729_n 0.0297827f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_43 VNB N_RESET_B_c_730_n 0.00596627f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.84
cc_44 VNB N_RESET_B_c_731_n 0.0107969f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.295
cc_45 VNB N_RESET_B_M1029_g 0.0388421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_RESET_B_c_733_n 0.0155168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_734_n 0.00231363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_RESET_B_c_735_n 0.0311795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_RESET_B_c_736_n 0.0255134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_c_737_n 7.11823e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_RESET_B_c_738_n 0.022755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_RESET_B_c_739_n 5.84685e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_RESET_B_c_740_n 0.00257692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB RESET_B 6.99951e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_RESET_B_c_742_n 0.0358283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_RESET_B_c_743_n 0.00523184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_c_744_n 0.0144561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_c_745_n 0.0225137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_RESET_B_c_746_n 0.00203128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_590_116#_c_971_n 0.0317387f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.68
cc_61 VNB N_A_590_116#_c_972_n 0.0174916f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.075
cc_62 VNB N_A_590_116#_c_973_n 0.0201031f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.79
cc_63 VNB N_A_590_116#_M1000_g 0.0200276f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.47
cc_64 VNB N_A_590_116#_c_975_n 0.00502958f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.24
cc_65 VNB N_A_590_116#_c_976_n 0.0181733f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_66 VNB N_A_590_116#_M1007_g 0.0201694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_590_116#_c_978_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_590_116#_c_979_n 0.00584545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_590_116#_c_980_n 0.00700779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_590_116#_c_981_n 0.00381702f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.925
cc_71 VNB N_A_590_116#_c_982_n 0.0177086f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.295
cc_72 VNB N_A_590_116#_c_983_n 0.00164143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_590_116#_c_984_n 0.00506651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_590_116#_c_985_n 0.00580661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_590_116#_c_986_n 0.032032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_560_90#_M1016_g 0.0497683f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.68
cc_77 VNB N_A_560_90#_M1039_g 0.00749286f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.075
cc_78 VNB N_A_560_90#_M1006_g 0.0296223f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_79 VNB N_A_560_90#_M1041_g 0.0317881f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.295
cc_80 VNB N_A_560_90#_M1044_g 0.00834745f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.925
cc_81 VNB N_A_560_90#_c_1153_n 0.0241269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_560_90#_c_1154_n 0.00925636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_560_90#_M1036_g 0.0323156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_560_90#_c_1156_n 0.0132692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_560_90#_c_1157_n 0.00196545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_560_90#_c_1158_n 0.059073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_560_90#_c_1159_n 0.0189801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_560_90#_c_1160_n 5.32607e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_560_90#_c_1161_n 0.0177089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_560_90#_c_1162_n 0.00866153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_560_90#_c_1163_n 0.0183484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_560_90#_c_1164_n 0.00645281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_560_90#_c_1165_n 0.00249638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2102_25#_M1032_g 0.0397833f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.68
cc_95 VNB N_A_2102_25#_M1013_g 0.0198389f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.79
cc_96 VNB N_A_2102_25#_c_1392_n 0.0245854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2102_25#_c_1393_n 0.00770327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2102_25#_c_1394_n 0.0133888f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_99 VNB N_A_2102_25#_c_1395_n 0.00467874f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=1.21
cc_100 VNB N_A_2102_25#_c_1396_n 0.0271511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2102_25#_c_1397_n 0.00311713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2102_25#_c_1398_n 0.0407017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2102_25#_c_1399_n 0.00283737f $X=-0.19 $Y=-0.245 $X2=2.15
+ $Y2=1.295
cc_104 VNB N_A_1799_379#_M1030_g 0.02833f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.79
cc_105 VNB N_A_1799_379#_c_1467_n 0.0295198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1799_379#_c_1468_n 0.0134078f $X=-0.19 $Y=-0.245 $X2=2.15
+ $Y2=1.545
cc_107 VNB N_A_1799_379#_M1050_g 0.0252356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1799_379#_c_1470_n 0.00502958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1799_379#_M1035_g 0.0283974f $X=-0.19 $Y=-0.245 $X2=2.15
+ $Y2=1.295
cc_110 VNB N_A_1799_379#_M1011_g 0.00935108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1799_379#_c_1473_n 0.0612896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1799_379#_M1042_g 0.0264366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1799_379#_M1028_g 0.00874667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1799_379#_c_1476_n 0.00502958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1799_379#_M1048_g 0.024082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_1799_379#_M1025_g 0.00696952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_1799_379#_c_1479_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_1799_379#_c_1480_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_1799_379#_c_1481_n 0.00487614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_1799_379#_c_1482_n 0.00764021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_1799_379#_c_1483_n 0.0015599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_1799_379#_c_1484_n 0.00790057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_1799_379#_c_1485_n 0.0222077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_1799_379#_c_1486_n 7.98171e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_1799_379#_c_1487_n 0.0168082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_1799_379#_c_1488_n 0.00235566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_1799_379#_c_1489_n 0.0102318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_1799_379#_c_1490_n 0.00359482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_1799_379#_c_1491_n 0.0347943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_1799_379#_c_1492_n 0.0413941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_1799_379#_c_1493_n 0.0301423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_CLK_M1026_g 0.0408888f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.495
cc_133 VNB N_CLK_M1049_g 0.0170139f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.62
cc_134 VNB N_CLK_c_1717_n 0.00563292f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.68
cc_135 VNB N_CLK_M1027_g 0.0338835f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.79
cc_136 VNB N_CLK_M1034_g 0.0202628f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.47
cc_137 VNB N_CLK_c_1720_n 0.00660243f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.24
cc_138 VNB CLK 0.0140569f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_139 VNB N_CLK_c_1722_n 0.0289116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_3222_137#_M1015_g 0.0226389f $X=-0.19 $Y=-0.245 $X2=1.805
+ $Y2=2.68
cc_141 VNB N_A_3222_137#_M1037_g 0.00101744f $X=-0.19 $Y=-0.245 $X2=2.06
+ $Y2=0.79
cc_142 VNB N_A_3222_137#_M1018_g 0.0249073f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.47
cc_143 VNB N_A_3222_137#_M1046_g 0.00112085f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=0.47
cc_144 VNB N_A_3222_137#_c_1776_n 0.0102002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_A_3222_137#_c_1777_n 0.0278334f $X=-0.19 $Y=-0.245 $X2=2.15
+ $Y2=1.295
cc_146 VNB N_A_3222_137#_c_1778_n 0.00152723f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=0.555
cc_147 VNB N_A_3222_137#_c_1779_n 0.0378831f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=0.925
cc_148 VNB N_A_111_457#_c_1875_n 0.0101429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VPWR_c_1950_n 0.760753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_Q_N_c_2228_n 0.0205568f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.84
cc_151 VNB N_Q_c_2251_n 0.0567461f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.84
cc_152 VNB N_VGND_c_2266_n 0.0389871f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.075
cc_153 VNB N_VGND_c_2267_n 0.00686134f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_154 VNB N_VGND_c_2268_n 0.0447885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2269_n 0.0193816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2270_n 0.0036965f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.295
cc_157 VNB N_VGND_c_2271_n 0.00299757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2272_n 0.0197306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2273_n 0.0357155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2274_n 0.0935127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2275_n 0.0949687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2276_n 0.0822514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2277_n 0.0628569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2278_n 0.0273851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2279_n 1.02519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2280_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2281_n 0.00632031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2282_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2283_n 0.00525412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2284_n 0.00514402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2285_n 0.00536178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VPB N_D_M1043_g 0.0416136f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.495
cc_173 VPB N_D_c_335_n 0.0916243f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=3.15
cc_174 VPB N_D_c_336_n 0.012806f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=3.15
cc_175 VPB N_D_M1012_g 0.0700537f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.68
cc_176 VPB N_A_662_90#_M1010_g 0.0355747f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.79
cc_177 VPB N_A_662_90#_M1019_g 0.0276482f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.545
cc_178 VPB N_A_662_90#_c_408_n 0.0112955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_817_90#_c_566_n 0.0179679f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.47
cc_180 VPB N_A_817_90#_M1002_g 0.0205836f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.24
cc_181 VPB N_A_817_90#_c_561_n 0.0237807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_817_90#_c_569_n 0.0243988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_817_90#_c_570_n 0.00333208f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.295
cc_184 VPB N_A_817_90#_c_562_n 0.00863103f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=0.555
cc_185 VPB N_A_817_90#_c_572_n 0.013701f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=0.925
cc_186 VPB N_A_817_90#_c_573_n 0.00851135f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=1.295
cc_187 VPB N_A_817_90#_c_563_n 0.00380005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_817_90#_c_575_n 0.0034822f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_817_90#_c_576_n 0.00349632f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_817_90#_c_577_n 2.09657e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_817_90#_c_578_n 0.00293488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_817_90#_c_579_n 0.00942575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_817_90#_c_565_n 0.00135473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_RESET_B_c_722_n 0.0164914f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=3.075
cc_195 VPB N_RESET_B_M1014_g 0.0393212f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.495
cc_196 VPB N_RESET_B_M1022_g 0.0340384f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.62
cc_197 VPB N_RESET_B_c_750_n 0.0164705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_RESET_B_c_751_n 0.0196896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_RESET_B_c_731_n 0.0133658f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.295
cc_200 VPB N_RESET_B_M1017_g 0.0223489f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.295
cc_201 VPB N_RESET_B_M1001_g 0.0209597f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=1.295
cc_202 VPB N_RESET_B_c_734_n 0.0558337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_RESET_B_c_736_n 0.0149375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_RESET_B_c_737_n 9.30065e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_RESET_B_c_738_n 0.0771286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_RESET_B_c_739_n 7.02262e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_740_n 0.00160081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB RESET_B 9.18192e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_590_116#_M1000_g 0.0234286f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.47
cc_210 VPB N_A_590_116#_M1007_g 0.0191472f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_590_116#_c_980_n 5.94689e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_590_116#_c_990_n 0.00347175f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.295
cc_213 VPB N_A_590_116#_c_991_n 0.0166539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_590_116#_c_981_n 4.75617e-19 $X=-0.19 $Y=1.655 $X2=1.94 $Y2=0.925
cc_215 VPB N_A_590_116#_c_993_n 0.0102584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_590_116#_c_994_n 0.00213814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_590_116#_c_995_n 0.00151808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_590_116#_c_996_n 0.00137324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_590_116#_c_997_n 0.00658792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_590_116#_c_985_n 0.00320028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_590_116#_c_986_n 0.0174682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_560_90#_M1016_g 0.00916085f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.68
cc_223 VPB N_A_560_90#_M1024_g 0.0519765f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.545
cc_224 VPB N_A_560_90#_c_1168_n 0.304904f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_560_90#_c_1169_n 0.012806f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.545
cc_226 VPB N_A_560_90#_M1039_g 0.0269633f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.075
cc_227 VPB N_A_560_90#_c_1171_n 0.00984309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_560_90#_M1047_g 0.0415956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_560_90#_c_1173_n 0.125212f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.295
cc_230 VPB N_A_560_90#_M1044_g 0.0253463f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=0.925
cc_231 VPB N_A_560_90#_c_1175_n 0.0222535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_560_90#_c_1156_n 0.0105623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_560_90#_c_1177_n 0.0257182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_560_90#_c_1178_n 0.00652136f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_560_90#_c_1179_n 0.0106415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_560_90#_c_1180_n 0.00204926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_560_90#_c_1165_n 0.00105389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_2102_25#_M1013_g 0.0888344f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.79
cc_239 VPB N_A_2102_25#_c_1394_n 0.00626278f $X=-0.19 $Y=1.655 $X2=1.595
+ $Y2=0.47
cc_240 VPB N_A_1799_379#_M1008_g 0.033539f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.68
cc_241 VPB N_A_1799_379#_M1020_g 0.0567833f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.47
cc_242 VPB N_A_1799_379#_M1031_g 0.0203634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1799_379#_M1011_g 0.023443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_1799_379#_M1028_g 0.0237323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_1799_379#_M1025_g 0.0219563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_1799_379#_c_1500_n 0.0186056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_1799_379#_c_1483_n 0.00221511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_1799_379#_c_1502_n 8.74713e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_1799_379#_c_1503_n 0.0189463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_1799_379#_c_1504_n 0.0100016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_1799_379#_c_1505_n 0.0220184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_1799_379#_c_1506_n 0.00307397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_1799_379#_c_1507_n 9.93275e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_1799_379#_c_1508_n 0.0212494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_1799_379#_c_1509_n 2.33253e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_A_1799_379#_c_1484_n 0.00118438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_1799_379#_c_1511_n 4.9792e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_1799_379#_c_1485_n 0.0169418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_1799_379#_c_1486_n 2.45591e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_1799_379#_c_1487_n 0.0104881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_1799_379#_c_1489_n 0.0276057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_1799_379#_c_1490_n 0.00311875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_1799_379#_c_1491_n 0.0109386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_1799_379#_c_1493_n 0.00992908f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_CLK_M1049_g 0.0225668f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.62
cc_266 VPB N_CLK_M1034_g 0.0217542f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.47
cc_267 VPB N_A_3222_137#_M1037_g 0.0215386f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.79
cc_268 VPB N_A_3222_137#_M1046_g 0.0234886f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.47
cc_269 VPB N_A_3222_137#_c_1782_n 0.0145016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_27_457#_c_1834_n 0.0362573f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.68
cc_271 VPB N_A_27_457#_c_1835_n 0.0146873f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=1.075
cc_272 VPB N_A_27_457#_c_1836_n 0.00956189f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.79
cc_273 VPB N_A_27_457#_c_1837_n 0.00235003f $X=-0.19 $Y=1.655 $X2=1.805
+ $Y2=1.545
cc_274 VPB N_A_27_457#_c_1838_n 0.00593433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_27_457#_c_1839_n 0.0073948f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.24
cc_276 VPB N_A_111_457#_c_1876_n 0.00282771f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.79
cc_277 VPB N_A_111_457#_c_1877_n 0.0311034f $X=-0.19 $Y=1.655 $X2=1.805
+ $Y2=1.545
cc_278 VPB N_A_111_457#_c_1878_n 0.0194149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_111_457#_c_1875_n 0.00597442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_A_111_457#_c_1880_n 6.46213e-19 $X=-0.19 $Y=1.655 $X2=1.595
+ $Y2=0.47
cc_281 VPB N_A_111_457#_c_1881_n 0.0132515f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.84
cc_282 VPB N_A_111_457#_c_1882_n 0.0028613f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_283 VPB N_A_111_457#_c_1883_n 0.00728957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_111_457#_c_1884_n 9.28569e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1951_n 0.00422685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_1952_n 0.0148966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_1953_n 0.0139786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_1954_n 0.0117443f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=0.555
cc_289 VPB N_VPWR_c_1955_n 0.00832397f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=0.925
cc_290 VPB N_VPWR_c_1956_n 0.0227373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1957_n 0.0256831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_1958_n 0.0701769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_1959_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_1960_n 0.0468907f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_1961_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_1962_n 0.0523754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_1963_n 0.00516759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_1964_n 0.0362112f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_1965_n 0.0536138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_1966_n 0.0912081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_1967_n 0.0579165f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_1968_n 0.0271876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_1950_n 0.192798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_1970_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_1971_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_1972_n 0.00356964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_1973_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_308 VPB N_A_484_411#_c_2103_n 0.0103219f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.68
cc_309 VPB N_A_484_411#_c_2104_n 0.0335241f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=1.075
cc_310 VPB N_A_484_411#_c_2105_n 0.00542972f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.79
cc_311 VPB N_A_484_411#_c_2106_n 0.0147855f $X=-0.19 $Y=1.655 $X2=1.805
+ $Y2=1.545
cc_312 VPB N_A_1712_379#_c_2146_n 0.0253826f $X=-0.19 $Y=1.655 $X2=1.805
+ $Y2=2.68
cc_313 VPB N_A_1712_379#_c_2147_n 0.0225146f $X=-0.19 $Y=1.655 $X2=2.06
+ $Y2=1.075
cc_314 VPB N_A_1712_379#_c_2148_n 0.00470318f $X=-0.19 $Y=1.655 $X2=2.06
+ $Y2=0.79
cc_315 VPB N_A_1712_379#_c_2149_n 0.00685658f $X=-0.19 $Y=1.655 $X2=1.805
+ $Y2=1.545
cc_316 VPB N_A_2185_397#_c_2173_n 0.0157695f $X=-0.19 $Y=1.655 $X2=1.805
+ $Y2=3.075
cc_317 VPB N_A_2185_397#_c_2174_n 0.0397115f $X=-0.19 $Y=1.655 $X2=1.805
+ $Y2=2.68
cc_318 VPB N_A_2185_397#_c_2175_n 0.00353434f $X=-0.19 $Y=1.655 $X2=1.805
+ $Y2=2.68
cc_319 VPB N_A_2185_397#_c_2176_n 0.0121987f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.79
cc_320 VPB N_A_2185_397#_c_2177_n 0.00870642f $X=-0.19 $Y=1.655 $X2=2.06
+ $Y2=0.79
cc_321 VPB N_A_2185_397#_c_2178_n 4.71231e-19 $X=-0.19 $Y=1.655 $X2=1.805
+ $Y2=1.545
cc_322 VPB N_A_2185_397#_c_2179_n 0.0195016f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.47
cc_323 VPB N_A_2185_397#_c_2180_n 0.0152146f $X=-0.19 $Y=1.655 $X2=2.15
+ $Y2=1.075
cc_324 VPB N_Q_N_c_2228_n 0.0275303f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.84
cc_325 VPB N_Q_c_2251_n 0.0543794f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.84
cc_326 N_D_M1012_g N_RESET_B_c_722_n 0.0201172f $X=1.805 $Y=2.68 $X2=-0.19
+ $Y2=-0.245
cc_327 N_D_M1043_g N_RESET_B_M1014_g 0.0126828f $X=0.48 $Y=2.495 $X2=0 $Y2=0
cc_328 N_D_c_335_n N_RESET_B_M1014_g 0.00737233f $X=1.73 $Y=3.15 $X2=0 $Y2=0
cc_329 N_D_c_335_n N_RESET_B_M1022_g 0.0085158f $X=1.73 $Y=3.15 $X2=0 $Y2=0
cc_330 N_D_c_329_n N_RESET_B_c_723_n 9.83269e-19 $X=2.15 $Y=1.47 $X2=0 $Y2=0
cc_331 N_D_c_330_n N_RESET_B_c_723_n 0.0221094f $X=2.15 $Y=1.24 $X2=0 $Y2=0
cc_332 D N_RESET_B_c_723_n 0.0105213f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_333 N_D_c_331_n N_RESET_B_M1033_g 0.0221094f $X=2.15 $Y=1.075 $X2=0 $Y2=0
cc_334 D N_RESET_B_M1033_g 0.0285538f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_335 N_D_c_331_n N_RESET_B_c_726_n 0.010097f $X=2.15 $Y=1.075 $X2=0 $Y2=0
cc_336 D N_RESET_B_c_726_n 0.00716522f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_337 N_D_M1012_g N_RESET_B_c_736_n 0.00495351f $X=1.805 $Y=2.68 $X2=0 $Y2=0
cc_338 N_D_c_329_n N_RESET_B_c_736_n 0.0100773f $X=2.15 $Y=1.47 $X2=0 $Y2=0
cc_339 D N_RESET_B_c_736_n 0.0225757f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_340 N_D_M1012_g N_RESET_B_c_737_n 2.32452e-19 $X=1.805 $Y=2.68 $X2=0 $Y2=0
cc_341 N_D_c_329_n N_RESET_B_c_737_n 2.81584e-19 $X=2.15 $Y=1.47 $X2=0 $Y2=0
cc_342 N_D_c_329_n N_RESET_B_c_742_n 0.0201172f $X=2.15 $Y=1.47 $X2=0 $Y2=0
cc_343 D N_RESET_B_c_742_n 0.00239423f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_344 N_D_c_333_n N_RESET_B_c_742_n 0.00263598f $X=2.15 $Y=1.295 $X2=0 $Y2=0
cc_345 N_D_c_329_n N_RESET_B_c_743_n 0.00250416f $X=2.15 $Y=1.47 $X2=0 $Y2=0
cc_346 N_D_c_330_n N_RESET_B_c_743_n 2.04979e-19 $X=2.15 $Y=1.24 $X2=0 $Y2=0
cc_347 D N_RESET_B_c_743_n 0.0213407f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_348 N_D_c_330_n N_A_560_90#_M1016_g 0.0105961f $X=2.15 $Y=1.24 $X2=0 $Y2=0
cc_349 N_D_c_331_n N_A_560_90#_M1016_g 0.00472602f $X=2.15 $Y=1.075 $X2=0 $Y2=0
cc_350 D N_A_560_90#_M1016_g 0.00407427f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_351 N_D_M1043_g N_A_27_457#_c_1834_n 0.00853225f $X=0.48 $Y=2.495 $X2=0 $Y2=0
cc_352 N_D_M1043_g N_A_27_457#_c_1835_n 0.0169992f $X=0.48 $Y=2.495 $X2=0 $Y2=0
cc_353 N_D_c_335_n N_A_27_457#_c_1835_n 0.0107537f $X=1.73 $Y=3.15 $X2=0 $Y2=0
cc_354 N_D_M1012_g N_A_27_457#_c_1835_n 7.2158e-19 $X=1.805 $Y=2.68 $X2=0 $Y2=0
cc_355 N_D_M1043_g N_A_27_457#_c_1837_n 0.00168893f $X=0.48 $Y=2.495 $X2=0 $Y2=0
cc_356 N_D_M1012_g N_A_27_457#_c_1837_n 6.62309e-19 $X=1.805 $Y=2.68 $X2=0 $Y2=0
cc_357 N_D_c_335_n N_A_27_457#_c_1838_n 0.00224846f $X=1.73 $Y=3.15 $X2=0 $Y2=0
cc_358 N_D_M1012_g N_A_27_457#_c_1838_n 0.0137717f $X=1.805 $Y=2.68 $X2=0 $Y2=0
cc_359 N_D_M1012_g N_A_27_457#_c_1839_n 8.26992e-19 $X=1.805 $Y=2.68 $X2=0 $Y2=0
cc_360 D N_A_111_457#_M1023_d 0.00422502f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_361 N_D_M1043_g N_A_111_457#_c_1876_n 0.012469f $X=0.48 $Y=2.495 $X2=0 $Y2=0
cc_362 N_D_M1012_g N_A_111_457#_c_1877_n 0.0141546f $X=1.805 $Y=2.68 $X2=0 $Y2=0
cc_363 N_D_c_329_n N_A_111_457#_c_1877_n 0.00677985f $X=2.15 $Y=1.47 $X2=0 $Y2=0
cc_364 D N_A_111_457#_c_1877_n 0.01216f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_365 N_D_M1012_g N_A_111_457#_c_1875_n 0.00672804f $X=1.805 $Y=2.68 $X2=0
+ $Y2=0
cc_366 N_D_c_330_n N_A_111_457#_c_1875_n 0.00757164f $X=2.15 $Y=1.24 $X2=0 $Y2=0
cc_367 N_D_c_331_n N_A_111_457#_c_1875_n 0.00146349f $X=2.15 $Y=1.075 $X2=0
+ $Y2=0
cc_368 D N_A_111_457#_c_1875_n 0.0712434f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_369 N_D_c_335_n N_VPWR_c_1951_n 0.022144f $X=1.73 $Y=3.15 $X2=0 $Y2=0
cc_370 N_D_M1012_g N_VPWR_c_1951_n 0.0104314f $X=1.805 $Y=2.68 $X2=0 $Y2=0
cc_371 N_D_c_335_n N_VPWR_c_1958_n 0.00486043f $X=1.73 $Y=3.15 $X2=0 $Y2=0
cc_372 N_D_c_336_n N_VPWR_c_1964_n 0.0247602f $X=0.555 $Y=3.15 $X2=0 $Y2=0
cc_373 N_D_c_335_n N_VPWR_c_1950_n 0.0276202f $X=1.73 $Y=3.15 $X2=0 $Y2=0
cc_374 N_D_c_336_n N_VPWR_c_1950_n 0.00557629f $X=0.555 $Y=3.15 $X2=0 $Y2=0
cc_375 N_D_M1012_g N_A_484_411#_c_2103_n 0.00127507f $X=1.805 $Y=2.68 $X2=0
+ $Y2=0
cc_376 N_D_M1012_g N_A_484_411#_c_2105_n 0.002698f $X=1.805 $Y=2.68 $X2=0 $Y2=0
cc_377 D N_VGND_c_2266_n 0.0164114f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_378 D N_VGND_c_2274_n 0.0240428f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_379 D N_VGND_c_2279_n 0.0253328f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_380 N_A_662_90#_c_402_n N_A_817_90#_M1004_s 0.0028778f $X=6.56 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_381 N_A_662_90#_c_392_n N_A_817_90#_M1003_g 0.0107777f $X=3.385 $Y=1.075
+ $X2=0 $Y2=0
cc_382 N_A_662_90#_c_398_n N_A_817_90#_M1003_g 0.00435608f $X=3.68 $Y=1.295
+ $X2=0 $Y2=0
cc_383 N_A_662_90#_c_399_n N_A_817_90#_M1003_g 0.0210385f $X=3.68 $Y=1.295 $X2=0
+ $Y2=0
cc_384 N_A_662_90#_c_400_n N_A_817_90#_M1003_g 0.0124348f $X=5.225 $Y=0.835
+ $X2=0 $Y2=0
cc_385 N_A_662_90#_M1010_g N_A_817_90#_c_559_n 0.002413f $X=3.465 $Y=2.265 $X2=0
+ $Y2=0
cc_386 N_A_662_90#_c_400_n N_A_817_90#_c_562_n 0.00584974f $X=5.225 $Y=0.835
+ $X2=0 $Y2=0
cc_387 N_A_662_90#_c_401_n N_A_817_90#_c_562_n 0.00416148f $X=5.31 $Y=0.75 $X2=0
+ $Y2=0
cc_388 N_A_662_90#_c_402_n N_A_817_90#_c_562_n 0.0195854f $X=6.56 $Y=0.35 $X2=0
+ $Y2=0
cc_389 N_A_662_90#_c_404_n N_A_817_90#_c_562_n 0.0269116f $X=6.645 $Y=1.175
+ $X2=0 $Y2=0
cc_390 N_A_662_90#_c_406_n N_A_817_90#_c_562_n 0.0133538f $X=6.73 $Y=1.26 $X2=0
+ $Y2=0
cc_391 N_A_662_90#_M1047_d N_A_817_90#_c_572_n 0.0115322f $X=7.76 $Y=2.065 $X2=0
+ $Y2=0
cc_392 N_A_662_90#_c_408_n N_A_817_90#_c_572_n 0.020035f $X=8.005 $Y=1.7 $X2=0
+ $Y2=0
cc_393 N_A_662_90#_M1019_g N_A_817_90#_c_573_n 0.00330453f $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_394 N_A_662_90#_c_408_n N_A_817_90#_c_573_n 0.0121726f $X=8.005 $Y=1.7 $X2=0
+ $Y2=0
cc_395 N_A_662_90#_c_394_n N_A_817_90#_c_563_n 0.00632052f $X=8.92 $Y=1.345
+ $X2=0 $Y2=0
cc_396 N_A_662_90#_M1019_g N_A_817_90#_c_563_n 0.00955883f $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_397 N_A_662_90#_c_409_n N_A_817_90#_c_563_n 0.0208072f $X=8.41 $Y=1.26 $X2=0
+ $Y2=0
cc_398 N_A_662_90#_c_394_n N_A_817_90#_c_575_n 2.32278e-19 $X=8.92 $Y=1.345
+ $X2=0 $Y2=0
cc_399 N_A_662_90#_c_408_n N_A_817_90#_c_575_n 0.0126021f $X=8.005 $Y=1.7 $X2=0
+ $Y2=0
cc_400 N_A_662_90#_c_409_n N_A_817_90#_c_575_n 0.0128148f $X=8.41 $Y=1.26 $X2=0
+ $Y2=0
cc_401 N_A_662_90#_c_394_n N_A_817_90#_c_564_n 0.0166808f $X=8.92 $Y=1.345 $X2=0
+ $Y2=0
cc_402 N_A_662_90#_M1019_g N_A_817_90#_c_564_n 0.0107753f $X=8.92 $Y=2.105 $X2=0
+ $Y2=0
cc_403 N_A_662_90#_c_396_n N_A_817_90#_c_564_n 0.016992f $X=9.305 $Y=1.06 $X2=0
+ $Y2=0
cc_404 N_A_662_90#_c_397_n N_A_817_90#_c_564_n 0.0105564f $X=9.38 $Y=0.985 $X2=0
+ $Y2=0
cc_405 N_A_662_90#_c_409_n N_A_817_90#_c_564_n 0.0129587f $X=8.41 $Y=1.26 $X2=0
+ $Y2=0
cc_406 N_A_662_90#_c_410_n N_A_817_90#_c_564_n 0.0370861f $X=8.575 $Y=0.84 $X2=0
+ $Y2=0
cc_407 N_A_662_90#_M1019_g N_A_817_90#_c_576_n 0.00228675f $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_408 N_A_662_90#_M1019_g N_A_817_90#_c_577_n 0.00315366f $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_409 N_A_662_90#_M1019_g N_A_817_90#_c_565_n 0.00497929f $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_410 N_A_662_90#_c_392_n N_RESET_B_c_726_n 0.0106323f $X=3.385 $Y=1.075 $X2=0
+ $Y2=0
cc_411 N_A_662_90#_c_400_n N_RESET_B_c_726_n 0.00421019f $X=5.225 $Y=0.835 $X2=0
+ $Y2=0
cc_412 N_A_662_90#_c_447_p N_RESET_B_c_726_n 0.00424542f $X=3.845 $Y=0.835 $X2=0
+ $Y2=0
cc_413 N_A_662_90#_c_400_n N_RESET_B_M1040_g 0.0140596f $X=5.225 $Y=0.835 $X2=0
+ $Y2=0
cc_414 N_A_662_90#_c_401_n N_RESET_B_M1040_g 0.00407526f $X=5.31 $Y=0.75 $X2=0
+ $Y2=0
cc_415 N_A_662_90#_c_400_n N_RESET_B_c_729_n 0.0101296f $X=5.225 $Y=0.835 $X2=0
+ $Y2=0
cc_416 N_A_662_90#_M1010_g N_RESET_B_c_736_n 0.00735173f $X=3.465 $Y=2.265 $X2=0
+ $Y2=0
cc_417 N_A_662_90#_c_398_n N_RESET_B_c_736_n 0.00902387f $X=3.68 $Y=1.295 $X2=0
+ $Y2=0
cc_418 N_A_662_90#_c_399_n N_RESET_B_c_736_n 0.00161792f $X=3.68 $Y=1.295 $X2=0
+ $Y2=0
cc_419 N_A_662_90#_M1047_d N_RESET_B_c_738_n 0.00108866f $X=7.76 $Y=2.065 $X2=0
+ $Y2=0
cc_420 N_A_662_90#_M1019_g N_RESET_B_c_738_n 0.00635394f $X=8.92 $Y=2.105 $X2=0
+ $Y2=0
cc_421 N_A_662_90#_c_396_n N_RESET_B_c_738_n 0.00329371f $X=9.305 $Y=1.06 $X2=0
+ $Y2=0
cc_422 N_A_662_90#_c_405_n N_RESET_B_c_738_n 0.0413111f $X=7.815 $Y=1.26 $X2=0
+ $Y2=0
cc_423 N_A_662_90#_c_406_n N_RESET_B_c_738_n 0.00815548f $X=6.73 $Y=1.26 $X2=0
+ $Y2=0
cc_424 N_A_662_90#_c_408_n N_RESET_B_c_738_n 0.0280152f $X=8.005 $Y=1.7 $X2=0
+ $Y2=0
cc_425 N_A_662_90#_c_409_n N_RESET_B_c_738_n 0.0083474f $X=8.41 $Y=1.26 $X2=0
+ $Y2=0
cc_426 N_A_662_90#_c_411_n N_RESET_B_c_738_n 0.00267592f $X=7.98 $Y=1.26 $X2=0
+ $Y2=0
cc_427 N_A_662_90#_c_402_n N_A_590_116#_c_971_n 0.00486531f $X=6.56 $Y=0.35
+ $X2=0 $Y2=0
cc_428 N_A_662_90#_c_402_n N_A_590_116#_c_972_n 0.00158614f $X=6.56 $Y=0.35
+ $X2=0 $Y2=0
cc_429 N_A_662_90#_c_402_n N_A_590_116#_c_973_n 0.0148463f $X=6.56 $Y=0.35 $X2=0
+ $Y2=0
cc_430 N_A_662_90#_c_404_n N_A_590_116#_c_973_n 0.0025225f $X=6.645 $Y=1.175
+ $X2=0 $Y2=0
cc_431 N_A_662_90#_c_406_n N_A_590_116#_M1000_g 6.92819e-19 $X=6.73 $Y=1.26
+ $X2=0 $Y2=0
cc_432 N_A_662_90#_c_404_n N_A_590_116#_c_975_n 0.00283201f $X=6.645 $Y=1.175
+ $X2=0 $Y2=0
cc_433 N_A_662_90#_c_406_n N_A_590_116#_c_975_n 0.00269129f $X=6.73 $Y=1.26
+ $X2=0 $Y2=0
cc_434 N_A_662_90#_c_402_n N_A_590_116#_c_976_n 0.00340599f $X=6.56 $Y=0.35
+ $X2=0 $Y2=0
cc_435 N_A_662_90#_c_404_n N_A_590_116#_c_976_n 0.0113871f $X=6.645 $Y=1.175
+ $X2=0 $Y2=0
cc_436 N_A_662_90#_c_405_n N_A_590_116#_M1007_g 0.00498529f $X=7.815 $Y=1.26
+ $X2=0 $Y2=0
cc_437 N_A_662_90#_c_406_n N_A_590_116#_M1007_g 9.74143e-19 $X=6.73 $Y=1.26
+ $X2=0 $Y2=0
cc_438 N_A_662_90#_c_404_n N_A_590_116#_c_979_n 0.00140451f $X=6.645 $Y=1.175
+ $X2=0 $Y2=0
cc_439 N_A_662_90#_c_405_n N_A_590_116#_c_979_n 0.0081388f $X=7.815 $Y=1.26
+ $X2=0 $Y2=0
cc_440 N_A_662_90#_c_392_n N_A_590_116#_c_980_n 0.00146007f $X=3.385 $Y=1.075
+ $X2=0 $Y2=0
cc_441 N_A_662_90#_M1010_g N_A_590_116#_c_980_n 0.00544828f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_442 N_A_662_90#_c_399_n N_A_590_116#_c_980_n 0.0103641f $X=3.68 $Y=1.295
+ $X2=0 $Y2=0
cc_443 N_A_662_90#_M1010_g N_A_590_116#_c_990_n 0.0044159f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_444 N_A_662_90#_M1010_g N_A_590_116#_c_991_n 0.0173458f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_445 N_A_662_90#_c_398_n N_A_590_116#_c_991_n 0.0165698f $X=3.68 $Y=1.295
+ $X2=0 $Y2=0
cc_446 N_A_662_90#_c_399_n N_A_590_116#_c_991_n 0.00374957f $X=3.68 $Y=1.295
+ $X2=0 $Y2=0
cc_447 N_A_662_90#_M1010_g N_A_590_116#_c_981_n 0.00347279f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_448 N_A_662_90#_c_398_n N_A_590_116#_c_981_n 0.0136416f $X=3.68 $Y=1.295
+ $X2=0 $Y2=0
cc_449 N_A_662_90#_c_399_n N_A_590_116#_c_981_n 0.0011522f $X=3.68 $Y=1.295
+ $X2=0 $Y2=0
cc_450 N_A_662_90#_M1010_g N_A_590_116#_c_993_n 0.0048519f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_451 N_A_662_90#_c_400_n N_A_590_116#_c_982_n 0.0779285f $X=5.225 $Y=0.835
+ $X2=0 $Y2=0
cc_452 N_A_662_90#_c_402_n N_A_590_116#_c_982_n 0.00418334f $X=6.56 $Y=0.35
+ $X2=0 $Y2=0
cc_453 N_A_662_90#_c_398_n N_A_590_116#_c_983_n 0.0137327f $X=3.68 $Y=1.295
+ $X2=0 $Y2=0
cc_454 N_A_662_90#_c_399_n N_A_590_116#_c_983_n 0.00118427f $X=3.68 $Y=1.295
+ $X2=0 $Y2=0
cc_455 N_A_662_90#_c_400_n N_A_590_116#_c_983_n 0.0107945f $X=5.225 $Y=0.835
+ $X2=0 $Y2=0
cc_456 N_A_662_90#_M1010_g N_A_590_116#_c_994_n 3.52713e-19 $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_457 N_A_662_90#_c_392_n N_A_590_116#_c_984_n 0.0107895f $X=3.385 $Y=1.075
+ $X2=0 $Y2=0
cc_458 N_A_662_90#_c_398_n N_A_590_116#_c_984_n 0.0344495f $X=3.68 $Y=1.295
+ $X2=0 $Y2=0
cc_459 N_A_662_90#_c_402_n N_A_590_116#_c_985_n 0.00921894f $X=6.56 $Y=0.35
+ $X2=0 $Y2=0
cc_460 N_A_662_90#_c_392_n N_A_560_90#_M1016_g 0.0241934f $X=3.385 $Y=1.075
+ $X2=0 $Y2=0
cc_461 N_A_662_90#_M1010_g N_A_560_90#_M1016_g 0.00775143f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_462 N_A_662_90#_M1010_g N_A_560_90#_c_1168_n 0.00281468f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_463 N_A_662_90#_c_404_n N_A_560_90#_M1006_g 8.95979e-19 $X=6.645 $Y=1.175
+ $X2=0 $Y2=0
cc_464 N_A_662_90#_c_405_n N_A_560_90#_M1006_g 0.0127676f $X=7.815 $Y=1.26 $X2=0
+ $Y2=0
cc_465 N_A_662_90#_c_407_n N_A_560_90#_M1006_g 0.00223078f $X=7.98 $Y=0.765
+ $X2=0 $Y2=0
cc_466 N_A_662_90#_c_408_n N_A_560_90#_M1047_g 0.0153929f $X=8.005 $Y=1.7 $X2=0
+ $Y2=0
cc_467 N_A_662_90#_c_394_n N_A_560_90#_M1041_g 0.00797815f $X=8.92 $Y=1.345
+ $X2=0 $Y2=0
cc_468 N_A_662_90#_c_405_n N_A_560_90#_M1041_g 0.00866618f $X=7.815 $Y=1.26
+ $X2=0 $Y2=0
cc_469 N_A_662_90#_c_407_n N_A_560_90#_M1041_g 0.0156674f $X=7.98 $Y=0.765 $X2=0
+ $Y2=0
cc_470 N_A_662_90#_c_410_n N_A_560_90#_M1041_g 2.66352e-19 $X=8.575 $Y=0.84
+ $X2=0 $Y2=0
cc_471 N_A_662_90#_c_411_n N_A_560_90#_M1041_g 0.00326373f $X=7.98 $Y=1.26 $X2=0
+ $Y2=0
cc_472 N_A_662_90#_M1019_g N_A_560_90#_c_1173_n 0.00501791f $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_473 N_A_662_90#_M1019_g N_A_560_90#_c_1154_n 0.0284357f $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_474 N_A_662_90#_c_396_n N_A_560_90#_c_1154_n 0.00502068f $X=9.305 $Y=1.06
+ $X2=0 $Y2=0
cc_475 N_A_662_90#_c_397_n N_A_560_90#_M1036_g 0.0104933f $X=9.38 $Y=0.985 $X2=0
+ $Y2=0
cc_476 N_A_662_90#_M1010_g N_A_560_90#_c_1175_n 0.0184464f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_477 N_A_662_90#_c_405_n N_A_560_90#_c_1156_n 0.0122481f $X=7.815 $Y=1.26
+ $X2=0 $Y2=0
cc_478 N_A_662_90#_c_408_n N_A_560_90#_c_1156_n 0.00936775f $X=8.005 $Y=1.7
+ $X2=0 $Y2=0
cc_479 N_A_662_90#_c_411_n N_A_560_90#_c_1156_n 3.2432e-19 $X=7.98 $Y=1.26 $X2=0
+ $Y2=0
cc_480 N_A_662_90#_c_397_n N_A_560_90#_c_1157_n 2.20265e-19 $X=9.38 $Y=0.985
+ $X2=0 $Y2=0
cc_481 N_A_662_90#_c_396_n N_A_560_90#_c_1158_n 0.0104933f $X=9.305 $Y=1.06
+ $X2=0 $Y2=0
cc_482 N_A_662_90#_M1019_g N_A_1799_379#_c_1500_n 5.67725e-19 $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_483 N_A_662_90#_c_394_n N_A_1799_379#_c_1482_n 0.00100043f $X=8.92 $Y=1.345
+ $X2=0 $Y2=0
cc_484 N_A_662_90#_c_396_n N_A_1799_379#_c_1482_n 0.00469698f $X=9.305 $Y=1.06
+ $X2=0 $Y2=0
cc_485 N_A_662_90#_c_397_n N_A_1799_379#_c_1482_n 0.0122639f $X=9.38 $Y=0.985
+ $X2=0 $Y2=0
cc_486 N_A_662_90#_c_392_n N_A_111_457#_c_1875_n 5.25498e-19 $X=3.385 $Y=1.075
+ $X2=0 $Y2=0
cc_487 N_A_662_90#_M1010_g N_A_111_457#_c_1875_n 3.11337e-19 $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_488 N_A_662_90#_M1010_g N_A_111_457#_c_1880_n 5.37666e-19 $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_489 N_A_662_90#_M1010_g N_A_111_457#_c_1881_n 0.00971106f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_490 N_A_662_90#_M1010_g N_A_111_457#_c_1883_n 0.00921713f $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_491 N_A_662_90#_M1010_g N_A_484_411#_c_2104_n 4.23818e-19 $X=3.465 $Y=2.265
+ $X2=0 $Y2=0
cc_492 N_A_662_90#_M1019_g N_A_1712_379#_c_2146_n 0.0119435f $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_493 N_A_662_90#_M1019_g N_A_1712_379#_c_2147_n 8.06636e-19 $X=8.92 $Y=2.105
+ $X2=0 $Y2=0
cc_494 N_A_662_90#_c_400_n N_VGND_M1040_d 0.0124933f $X=5.225 $Y=0.835 $X2=0
+ $Y2=0
cc_495 N_A_662_90#_c_400_n N_VGND_c_2267_n 0.0245808f $X=5.225 $Y=0.835 $X2=0
+ $Y2=0
cc_496 N_A_662_90#_c_401_n N_VGND_c_2267_n 0.0100349f $X=5.31 $Y=0.75 $X2=0
+ $Y2=0
cc_497 N_A_662_90#_c_403_n N_VGND_c_2267_n 0.0141772f $X=5.395 $Y=0.35 $X2=0
+ $Y2=0
cc_498 N_A_662_90#_c_400_n N_VGND_c_2268_n 0.00253519f $X=5.225 $Y=0.835 $X2=0
+ $Y2=0
cc_499 N_A_662_90#_c_402_n N_VGND_c_2268_n 0.0815652f $X=6.56 $Y=0.35 $X2=0
+ $Y2=0
cc_500 N_A_662_90#_c_403_n N_VGND_c_2268_n 0.0114298f $X=5.395 $Y=0.35 $X2=0
+ $Y2=0
cc_501 N_A_662_90#_c_402_n N_VGND_c_2269_n 0.0096064f $X=6.56 $Y=0.35 $X2=0
+ $Y2=0
cc_502 N_A_662_90#_c_404_n N_VGND_c_2269_n 0.0188551f $X=6.645 $Y=1.175 $X2=0
+ $Y2=0
cc_503 N_A_662_90#_c_405_n N_VGND_c_2269_n 0.0257663f $X=7.815 $Y=1.26 $X2=0
+ $Y2=0
cc_504 N_A_662_90#_c_407_n N_VGND_c_2269_n 0.0137622f $X=7.98 $Y=0.765 $X2=0
+ $Y2=0
cc_505 N_A_662_90#_c_400_n N_VGND_c_2274_n 0.0101455f $X=5.225 $Y=0.835 $X2=0
+ $Y2=0
cc_506 N_A_662_90#_c_447_p N_VGND_c_2274_n 0.00503514f $X=3.845 $Y=0.835 $X2=0
+ $Y2=0
cc_507 N_A_662_90#_c_394_n N_VGND_c_2275_n 0.0012308f $X=8.92 $Y=1.345 $X2=0
+ $Y2=0
cc_508 N_A_662_90#_c_397_n N_VGND_c_2275_n 0.00549284f $X=9.38 $Y=0.985 $X2=0
+ $Y2=0
cc_509 N_A_662_90#_c_407_n N_VGND_c_2275_n 0.00824843f $X=7.98 $Y=0.765 $X2=0
+ $Y2=0
cc_510 N_A_662_90#_c_410_n N_VGND_c_2275_n 0.00536945f $X=8.575 $Y=0.84 $X2=0
+ $Y2=0
cc_511 N_A_662_90#_c_392_n N_VGND_c_2279_n 0.00264436f $X=3.385 $Y=1.075 $X2=0
+ $Y2=0
cc_512 N_A_662_90#_c_397_n N_VGND_c_2279_n 0.0119473f $X=9.38 $Y=0.985 $X2=0
+ $Y2=0
cc_513 N_A_662_90#_c_400_n N_VGND_c_2279_n 0.0278247f $X=5.225 $Y=0.835 $X2=0
+ $Y2=0
cc_514 N_A_662_90#_c_447_p N_VGND_c_2279_n 0.00920177f $X=3.845 $Y=0.835 $X2=0
+ $Y2=0
cc_515 N_A_662_90#_c_402_n N_VGND_c_2279_n 0.0493534f $X=6.56 $Y=0.35 $X2=0
+ $Y2=0
cc_516 N_A_662_90#_c_403_n N_VGND_c_2279_n 0.00657111f $X=5.395 $Y=0.35 $X2=0
+ $Y2=0
cc_517 N_A_662_90#_c_407_n N_VGND_c_2279_n 0.0106779f $X=7.98 $Y=0.765 $X2=0
+ $Y2=0
cc_518 N_A_662_90#_c_410_n N_VGND_c_2279_n 0.00924883f $X=8.575 $Y=0.84 $X2=0
+ $Y2=0
cc_519 N_A_662_90#_c_398_n A_692_116# 0.00104581f $X=3.68 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_520 N_A_662_90#_c_400_n A_692_116# 0.0102478f $X=5.225 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_521 N_A_662_90#_c_447_p A_692_116# 0.00820126f $X=3.845 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_522 N_A_662_90#_c_400_n A_847_116# 0.00338781f $X=5.225 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_523 N_A_817_90#_M1003_g N_RESET_B_c_726_n 0.0106323f $X=4.16 $Y=0.79 $X2=0
+ $Y2=0
cc_524 N_A_817_90#_M1003_g N_RESET_B_M1040_g 0.0433853f $X=4.16 $Y=0.79 $X2=0
+ $Y2=0
cc_525 N_A_817_90#_c_559_n N_RESET_B_c_730_n 0.0133818f $X=4.54 $Y=1.605 $X2=0
+ $Y2=0
cc_526 N_A_817_90#_c_560_n N_RESET_B_c_730_n 2.62692e-19 $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_527 N_A_817_90#_c_579_n N_RESET_B_c_751_n 0.00320118f $X=6.215 $Y=2.01 $X2=0
+ $Y2=0
cc_528 N_A_817_90#_M1003_g N_RESET_B_c_733_n 0.00433964f $X=4.16 $Y=0.79 $X2=0
+ $Y2=0
cc_529 N_A_817_90#_c_566_n N_RESET_B_c_734_n 0.0147404f $X=4.54 $Y=2.125 $X2=0
+ $Y2=0
cc_530 N_A_817_90#_M1002_g N_RESET_B_c_734_n 0.0205792f $X=4.54 $Y=2.495 $X2=0
+ $Y2=0
cc_531 N_A_817_90#_c_560_n N_RESET_B_c_734_n 0.00125636f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_532 N_A_817_90#_c_561_n N_RESET_B_c_734_n 0.010517f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_533 N_A_817_90#_c_569_n N_RESET_B_c_734_n 0.0303828f $X=6.05 $Y=2.045 $X2=0
+ $Y2=0
cc_534 N_A_817_90#_c_579_n N_RESET_B_c_734_n 0.00256258f $X=6.215 $Y=2.01 $X2=0
+ $Y2=0
cc_535 N_A_817_90#_c_559_n N_RESET_B_c_736_n 0.00366889f $X=4.54 $Y=1.605 $X2=0
+ $Y2=0
cc_536 N_A_817_90#_c_560_n N_RESET_B_c_736_n 0.018793f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_537 N_A_817_90#_c_561_n N_RESET_B_c_736_n 0.00283661f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_538 N_A_817_90#_c_569_n N_RESET_B_c_736_n 0.00812408f $X=6.05 $Y=2.045 $X2=0
+ $Y2=0
cc_539 N_A_817_90#_c_569_n N_RESET_B_c_738_n 0.0220131f $X=6.05 $Y=2.045 $X2=0
+ $Y2=0
cc_540 N_A_817_90#_c_562_n N_RESET_B_c_738_n 0.0398741f $X=6.215 $Y=0.765 $X2=0
+ $Y2=0
cc_541 N_A_817_90#_c_572_n N_RESET_B_c_738_n 0.0613164f $X=8.27 $Y=2.13 $X2=0
+ $Y2=0
cc_542 N_A_817_90#_c_573_n N_RESET_B_c_738_n 0.0103583f $X=8.355 $Y=2.045 $X2=0
+ $Y2=0
cc_543 N_A_817_90#_c_563_n N_RESET_B_c_738_n 0.019369f $X=8.92 $Y=1.61 $X2=0
+ $Y2=0
cc_544 N_A_817_90#_c_575_n N_RESET_B_c_738_n 0.00499957f $X=8.44 $Y=1.61 $X2=0
+ $Y2=0
cc_545 N_A_817_90#_c_576_n N_RESET_B_c_738_n 0.0112562f $X=9.165 $Y=1.875 $X2=0
+ $Y2=0
cc_546 N_A_817_90#_c_578_n N_RESET_B_c_738_n 0.0168642f $X=9.67 $Y=2.04 $X2=0
+ $Y2=0
cc_547 N_A_817_90#_c_565_n N_RESET_B_c_738_n 0.0187168f $X=9.085 $Y=1.61 $X2=0
+ $Y2=0
cc_548 N_A_817_90#_c_559_n N_RESET_B_c_739_n 7.08405e-19 $X=4.54 $Y=1.605 $X2=0
+ $Y2=0
cc_549 N_A_817_90#_c_560_n N_RESET_B_c_739_n 0.00259401f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_550 N_A_817_90#_c_561_n N_RESET_B_c_739_n 6.86316e-19 $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_551 N_A_817_90#_c_569_n N_RESET_B_c_739_n 0.00748991f $X=6.05 $Y=2.045 $X2=0
+ $Y2=0
cc_552 N_A_817_90#_c_559_n N_RESET_B_c_740_n 0.00172568f $X=4.54 $Y=1.605 $X2=0
+ $Y2=0
cc_553 N_A_817_90#_c_560_n N_RESET_B_c_740_n 0.0181532f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_554 N_A_817_90#_c_569_n N_RESET_B_c_740_n 0.0203928f $X=6.05 $Y=2.045 $X2=0
+ $Y2=0
cc_555 N_A_817_90#_c_559_n N_RESET_B_c_744_n 0.010517f $X=4.54 $Y=1.605 $X2=0
+ $Y2=0
cc_556 N_A_817_90#_c_560_n N_RESET_B_c_744_n 4.9476e-19 $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_557 N_A_817_90#_c_562_n N_A_590_116#_c_971_n 0.0183884f $X=6.215 $Y=0.765
+ $X2=0 $Y2=0
cc_558 N_A_817_90#_c_562_n N_A_590_116#_c_973_n 0.00809451f $X=6.215 $Y=0.765
+ $X2=0 $Y2=0
cc_559 N_A_817_90#_c_562_n N_A_590_116#_M1000_g 0.0215608f $X=6.215 $Y=0.765
+ $X2=0 $Y2=0
cc_560 N_A_817_90#_c_572_n N_A_590_116#_M1000_g 0.0110224f $X=8.27 $Y=2.13 $X2=0
+ $Y2=0
cc_561 N_A_817_90#_c_579_n N_A_590_116#_M1000_g 0.0142638f $X=6.215 $Y=2.01
+ $X2=0 $Y2=0
cc_562 N_A_817_90#_c_562_n N_A_590_116#_c_976_n 3.81289e-19 $X=6.215 $Y=0.765
+ $X2=0 $Y2=0
cc_563 N_A_817_90#_c_562_n N_A_590_116#_M1007_g 0.00363484f $X=6.215 $Y=0.765
+ $X2=0 $Y2=0
cc_564 N_A_817_90#_c_572_n N_A_590_116#_M1007_g 0.0148182f $X=8.27 $Y=2.13 $X2=0
+ $Y2=0
cc_565 N_A_817_90#_c_579_n N_A_590_116#_M1007_g 0.00221988f $X=6.215 $Y=2.01
+ $X2=0 $Y2=0
cc_566 N_A_817_90#_c_562_n N_A_590_116#_c_978_n 0.002498f $X=6.215 $Y=0.765
+ $X2=0 $Y2=0
cc_567 N_A_817_90#_M1003_g N_A_590_116#_c_981_n 0.00936084f $X=4.16 $Y=0.79
+ $X2=0 $Y2=0
cc_568 N_A_817_90#_c_559_n N_A_590_116#_c_981_n 0.00775721f $X=4.54 $Y=1.605
+ $X2=0 $Y2=0
cc_569 N_A_817_90#_c_560_n N_A_590_116#_c_981_n 0.0152452f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_570 N_A_817_90#_c_561_n N_A_590_116#_c_981_n 0.00129071f $X=4.54 $Y=1.62
+ $X2=0 $Y2=0
cc_571 N_A_817_90#_c_566_n N_A_590_116#_c_993_n 0.00114878f $X=4.54 $Y=2.125
+ $X2=0 $Y2=0
cc_572 N_A_817_90#_M1002_g N_A_590_116#_c_993_n 0.00554532f $X=4.54 $Y=2.495
+ $X2=0 $Y2=0
cc_573 N_A_817_90#_c_560_n N_A_590_116#_c_993_n 0.0074868f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_574 N_A_817_90#_c_561_n N_A_590_116#_c_993_n 0.00231676f $X=4.54 $Y=1.62
+ $X2=0 $Y2=0
cc_575 N_A_817_90#_c_570_n N_A_590_116#_c_993_n 0.0130305f $X=4.705 $Y=2.045
+ $X2=0 $Y2=0
cc_576 N_A_817_90#_M1003_g N_A_590_116#_c_982_n 0.00399937f $X=4.16 $Y=0.79
+ $X2=0 $Y2=0
cc_577 N_A_817_90#_c_559_n N_A_590_116#_c_982_n 0.00612819f $X=4.54 $Y=1.605
+ $X2=0 $Y2=0
cc_578 N_A_817_90#_c_560_n N_A_590_116#_c_982_n 0.0228289f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_579 N_A_817_90#_M1003_g N_A_590_116#_c_983_n 0.00407089f $X=4.16 $Y=0.79
+ $X2=0 $Y2=0
cc_580 N_A_817_90#_c_566_n N_A_590_116#_c_1056_n 9.66291e-19 $X=4.54 $Y=2.125
+ $X2=0 $Y2=0
cc_581 N_A_817_90#_M1002_g N_A_590_116#_c_1056_n 0.0123512f $X=4.54 $Y=2.495
+ $X2=0 $Y2=0
cc_582 N_A_817_90#_c_569_n N_A_590_116#_c_1056_n 0.0478901f $X=6.05 $Y=2.045
+ $X2=0 $Y2=0
cc_583 N_A_817_90#_c_570_n N_A_590_116#_c_1056_n 0.0208205f $X=4.705 $Y=2.045
+ $X2=0 $Y2=0
cc_584 N_A_817_90#_c_560_n N_A_590_116#_c_996_n 0.0129838f $X=4.54 $Y=1.62 $X2=0
+ $Y2=0
cc_585 N_A_817_90#_c_561_n N_A_590_116#_c_996_n 0.00361698f $X=4.54 $Y=1.62
+ $X2=0 $Y2=0
cc_586 N_A_817_90#_c_569_n N_A_590_116#_c_997_n 0.0219661f $X=6.05 $Y=2.045
+ $X2=0 $Y2=0
cc_587 N_A_817_90#_c_579_n N_A_590_116#_c_997_n 0.0308305f $X=6.215 $Y=2.01
+ $X2=0 $Y2=0
cc_588 N_A_817_90#_c_569_n N_A_590_116#_c_985_n 0.021766f $X=6.05 $Y=2.045 $X2=0
+ $Y2=0
cc_589 N_A_817_90#_c_562_n N_A_590_116#_c_985_n 0.0493072f $X=6.215 $Y=0.765
+ $X2=0 $Y2=0
cc_590 N_A_817_90#_c_569_n N_A_590_116#_c_986_n 0.00221622f $X=6.05 $Y=2.045
+ $X2=0 $Y2=0
cc_591 N_A_817_90#_c_562_n N_A_590_116#_c_986_n 0.00420846f $X=6.215 $Y=0.765
+ $X2=0 $Y2=0
cc_592 N_A_817_90#_M1002_g N_A_560_90#_c_1168_n 0.00863568f $X=4.54 $Y=2.495
+ $X2=0 $Y2=0
cc_593 N_A_817_90#_c_579_n N_A_560_90#_c_1168_n 0.00610504f $X=6.215 $Y=2.01
+ $X2=0 $Y2=0
cc_594 N_A_817_90#_c_572_n N_A_560_90#_M1039_g 0.0157625f $X=8.27 $Y=2.13 $X2=0
+ $Y2=0
cc_595 N_A_817_90#_c_572_n N_A_560_90#_c_1171_n 6.38093e-19 $X=8.27 $Y=2.13
+ $X2=0 $Y2=0
cc_596 N_A_817_90#_c_572_n N_A_560_90#_M1047_g 0.0172406f $X=8.27 $Y=2.13 $X2=0
+ $Y2=0
cc_597 N_A_817_90#_c_573_n N_A_560_90#_M1047_g 0.00449453f $X=8.355 $Y=2.045
+ $X2=0 $Y2=0
cc_598 N_A_817_90#_c_572_n N_A_560_90#_c_1173_n 0.013239f $X=8.27 $Y=2.13 $X2=0
+ $Y2=0
cc_599 N_A_817_90#_c_576_n N_A_560_90#_M1044_g 0.00391186f $X=9.165 $Y=1.875
+ $X2=0 $Y2=0
cc_600 N_A_817_90#_c_578_n N_A_560_90#_M1044_g 0.0133883f $X=9.67 $Y=2.04 $X2=0
+ $Y2=0
cc_601 N_A_817_90#_c_565_n N_A_560_90#_M1044_g 0.00120402f $X=9.085 $Y=1.61
+ $X2=0 $Y2=0
cc_602 N_A_817_90#_c_578_n N_A_560_90#_c_1153_n 0.00112164f $X=9.67 $Y=2.04
+ $X2=0 $Y2=0
cc_603 N_A_817_90#_c_564_n N_A_560_90#_c_1154_n 0.00145821f $X=9.085 $Y=0.58
+ $X2=0 $Y2=0
cc_604 N_A_817_90#_c_572_n N_A_560_90#_c_1156_n 0.00244034f $X=8.27 $Y=2.13
+ $X2=0 $Y2=0
cc_605 N_A_817_90#_c_577_n N_A_1799_379#_M1019_d 0.00669584f $X=9.25 $Y=2.04
+ $X2=0 $Y2=0
cc_606 N_A_817_90#_c_578_n N_A_1799_379#_M1019_d 7.68253e-19 $X=9.67 $Y=2.04
+ $X2=0 $Y2=0
cc_607 N_A_817_90#_M1044_d N_A_1799_379#_c_1500_n 0.00868656f $X=9.53 $Y=1.895
+ $X2=0 $Y2=0
cc_608 N_A_817_90#_c_577_n N_A_1799_379#_c_1500_n 0.0139107f $X=9.25 $Y=2.04
+ $X2=0 $Y2=0
cc_609 N_A_817_90#_c_578_n N_A_1799_379#_c_1500_n 0.0291688f $X=9.67 $Y=2.04
+ $X2=0 $Y2=0
cc_610 N_A_817_90#_c_564_n N_A_1799_379#_c_1482_n 0.0713685f $X=9.085 $Y=0.58
+ $X2=0 $Y2=0
cc_611 N_A_817_90#_c_578_n N_A_1799_379#_c_1502_n 0.0208699f $X=9.67 $Y=2.04
+ $X2=0 $Y2=0
cc_612 N_A_817_90#_c_565_n N_A_1799_379#_c_1502_n 0.0125721f $X=9.085 $Y=1.61
+ $X2=0 $Y2=0
cc_613 N_A_817_90#_c_578_n N_A_1799_379#_c_1503_n 0.0260314f $X=9.67 $Y=2.04
+ $X2=0 $Y2=0
cc_614 N_A_817_90#_M1002_g N_A_111_457#_c_1881_n 0.00305671f $X=4.54 $Y=2.495
+ $X2=0 $Y2=0
cc_615 N_A_817_90#_M1002_g N_A_111_457#_c_1883_n 0.00226005f $X=4.54 $Y=2.495
+ $X2=0 $Y2=0
cc_616 N_A_817_90#_c_572_n N_VPWR_M1007_d 0.00712376f $X=8.27 $Y=2.13 $X2=0
+ $Y2=0
cc_617 N_A_817_90#_M1002_g N_VPWR_c_1952_n 0.0017192f $X=4.54 $Y=2.495 $X2=0
+ $Y2=0
cc_618 N_A_817_90#_c_572_n N_VPWR_c_1953_n 0.0209601f $X=8.27 $Y=2.13 $X2=0
+ $Y2=0
cc_619 N_A_817_90#_c_579_n N_VPWR_c_1953_n 0.0110409f $X=6.215 $Y=2.01 $X2=0
+ $Y2=0
cc_620 N_A_817_90#_c_579_n N_VPWR_c_1965_n 0.00701036f $X=6.215 $Y=2.01 $X2=0
+ $Y2=0
cc_621 N_A_817_90#_M1002_g N_VPWR_c_1950_n 9.49986e-19 $X=4.54 $Y=2.495 $X2=0
+ $Y2=0
cc_622 N_A_817_90#_c_579_n N_VPWR_c_1950_n 0.00885159f $X=6.215 $Y=2.01 $X2=0
+ $Y2=0
cc_623 N_A_817_90#_M1002_g N_A_484_411#_c_2106_n 0.00408969f $X=4.54 $Y=2.495
+ $X2=0 $Y2=0
cc_624 N_A_817_90#_c_572_n A_1301_373# 0.00511004f $X=8.27 $Y=2.13 $X2=-0.19
+ $Y2=-0.245
cc_625 N_A_817_90#_c_572_n A_1480_413# 0.00303348f $X=8.27 $Y=2.13 $X2=-0.19
+ $Y2=-0.245
cc_626 N_A_817_90#_c_572_n N_A_1712_379#_c_2146_n 0.0139102f $X=8.27 $Y=2.13
+ $X2=0 $Y2=0
cc_627 N_A_817_90#_c_573_n N_A_1712_379#_c_2146_n 0.0124095f $X=8.355 $Y=2.045
+ $X2=0 $Y2=0
cc_628 N_A_817_90#_c_563_n N_A_1712_379#_c_2146_n 0.0168539f $X=8.92 $Y=1.61
+ $X2=0 $Y2=0
cc_629 N_A_817_90#_c_577_n N_A_1712_379#_c_2146_n 0.0227357f $X=9.25 $Y=2.04
+ $X2=0 $Y2=0
cc_630 N_A_817_90#_c_564_n N_VGND_c_2275_n 0.0216625f $X=9.085 $Y=0.58 $X2=0
+ $Y2=0
cc_631 N_A_817_90#_M1021_s N_VGND_c_2279_n 0.00494841f $X=8.94 $Y=0.235 $X2=0
+ $Y2=0
cc_632 N_A_817_90#_M1003_g N_VGND_c_2279_n 0.00264436f $X=4.16 $Y=0.79 $X2=0
+ $Y2=0
cc_633 N_A_817_90#_c_564_n N_VGND_c_2279_n 0.0126859f $X=9.085 $Y=0.58 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_738_n N_A_590_116#_c_971_n 0.00173918f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_635 N_RESET_B_c_729_n N_A_590_116#_c_972_n 0.0046719f $X=4.945 $Y=1.15 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_738_n N_A_590_116#_M1000_g 0.00730632f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_637 N_RESET_B_c_738_n N_A_590_116#_M1007_g 0.00577517f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_638 N_RESET_B_c_736_n N_A_590_116#_c_980_n 0.0145579f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_639 N_RESET_B_c_736_n N_A_590_116#_c_991_n 0.0331767f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_736_n N_A_590_116#_c_981_n 0.0138866f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_729_n N_A_590_116#_c_982_n 0.0140877f $X=4.945 $Y=1.15 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_730_n N_A_590_116#_c_982_n 0.00562898f $X=4.625 $Y=1.15 $X2=0
+ $Y2=0
cc_643 N_RESET_B_c_733_n N_A_590_116#_c_982_n 0.00426976f $X=5.11 $Y=1.45 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_736_n N_A_590_116#_c_982_n 0.0154706f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_645 N_RESET_B_c_738_n N_A_590_116#_c_982_n 0.0108017f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_646 N_RESET_B_c_739_n N_A_590_116#_c_982_n 0.00275012f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_647 N_RESET_B_c_740_n N_A_590_116#_c_982_n 0.022822f $X=5.04 $Y=1.665 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_744_n N_A_590_116#_c_982_n 0.00471135f $X=5.11 $Y=1.615 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_750_n N_A_590_116#_c_1056_n 0.0102004f $X=5.11 $Y=2.16 $X2=0
+ $Y2=0
cc_650 N_RESET_B_c_751_n N_A_590_116#_c_1056_n 0.00707517f $X=5.47 $Y=2.16 $X2=0
+ $Y2=0
cc_651 N_RESET_B_c_734_n N_A_590_116#_c_1056_n 9.49066e-19 $X=5.11 $Y=1.845
+ $X2=0 $Y2=0
cc_652 N_RESET_B_c_736_n N_A_590_116#_c_1056_n 0.00667708f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_653 N_RESET_B_c_726_n N_A_590_116#_c_984_n 0.00439759f $X=4.475 $Y=0.165
+ $X2=0 $Y2=0
cc_654 N_RESET_B_c_736_n N_A_590_116#_c_984_n 0.00530525f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_655 N_RESET_B_c_736_n N_A_590_116#_c_995_n 0.0109164f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_656 N_RESET_B_c_736_n N_A_590_116#_c_996_n 0.0105791f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_750_n N_A_590_116#_c_997_n 0.00116325f $X=5.11 $Y=2.16 $X2=0
+ $Y2=0
cc_658 N_RESET_B_c_751_n N_A_590_116#_c_997_n 0.00631723f $X=5.47 $Y=2.16 $X2=0
+ $Y2=0
cc_659 N_RESET_B_c_733_n N_A_590_116#_c_985_n 9.9612e-19 $X=5.11 $Y=1.45 $X2=0
+ $Y2=0
cc_660 N_RESET_B_c_738_n N_A_590_116#_c_985_n 0.0282209f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_661 N_RESET_B_c_739_n N_A_590_116#_c_985_n 4.60294e-19 $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_662 N_RESET_B_c_740_n N_A_590_116#_c_985_n 0.0145351f $X=5.04 $Y=1.665 $X2=0
+ $Y2=0
cc_663 N_RESET_B_c_744_n N_A_590_116#_c_985_n 5.16937e-19 $X=5.11 $Y=1.615 $X2=0
+ $Y2=0
cc_664 N_RESET_B_c_733_n N_A_590_116#_c_986_n 0.0046719f $X=5.11 $Y=1.45 $X2=0
+ $Y2=0
cc_665 N_RESET_B_c_734_n N_A_590_116#_c_986_n 2.86051e-19 $X=5.11 $Y=1.845 $X2=0
+ $Y2=0
cc_666 N_RESET_B_c_738_n N_A_590_116#_c_986_n 0.002185f $X=12.095 $Y=1.665 $X2=0
+ $Y2=0
cc_667 N_RESET_B_c_740_n N_A_590_116#_c_986_n 0.00119018f $X=5.04 $Y=1.665 $X2=0
+ $Y2=0
cc_668 N_RESET_B_c_744_n N_A_590_116#_c_986_n 0.015728f $X=5.11 $Y=1.615 $X2=0
+ $Y2=0
cc_669 N_RESET_B_c_726_n N_A_560_90#_M1016_g 0.0106323f $X=4.475 $Y=0.165 $X2=0
+ $Y2=0
cc_670 N_RESET_B_c_736_n N_A_560_90#_M1016_g 0.0076323f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_671 N_RESET_B_c_750_n N_A_560_90#_c_1168_n 0.00863568f $X=5.11 $Y=2.16 $X2=0
+ $Y2=0
cc_672 N_RESET_B_c_751_n N_A_560_90#_c_1168_n 0.00858532f $X=5.47 $Y=2.16 $X2=0
+ $Y2=0
cc_673 N_RESET_B_c_738_n N_A_560_90#_M1039_g 0.00568563f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_674 N_RESET_B_c_738_n N_A_560_90#_M1047_g 0.00662169f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_675 N_RESET_B_c_738_n N_A_560_90#_M1044_g 0.00393136f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_676 N_RESET_B_c_736_n N_A_560_90#_c_1175_n 0.00468585f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_677 N_RESET_B_c_738_n N_A_560_90#_c_1156_n 0.0024749f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_678 N_RESET_B_c_738_n N_A_560_90#_c_1157_n 0.0022156f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_679 N_RESET_B_M1029_g N_A_560_90#_c_1161_n 0.0115366f $X=12.39 $Y=0.465 $X2=0
+ $Y2=0
cc_680 N_RESET_B_c_738_n N_A_2102_25#_M1013_g 0.00745256f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_681 N_RESET_B_c_738_n N_A_2102_25#_c_1392_n 0.0104823f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_682 N_RESET_B_M1029_g N_A_2102_25#_c_1393_n 0.00408231f $X=12.39 $Y=0.465
+ $X2=0 $Y2=0
cc_683 N_RESET_B_c_738_n N_A_2102_25#_c_1394_n 0.0236054f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_684 RESET_B N_A_2102_25#_c_1394_n 0.00263338f $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_685 N_RESET_B_c_745_n N_A_2102_25#_c_1394_n 0.014808f $X=12.29 $Y=1.275 $X2=0
+ $Y2=0
cc_686 N_RESET_B_c_746_n N_A_2102_25#_c_1394_n 0.0386327f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_687 N_RESET_B_M1029_g N_A_2102_25#_c_1396_n 0.0166883f $X=12.39 $Y=0.465
+ $X2=0 $Y2=0
cc_688 N_RESET_B_c_745_n N_A_2102_25#_c_1396_n 0.00210122f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_689 N_RESET_B_c_746_n N_A_2102_25#_c_1396_n 0.0198855f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_690 N_RESET_B_c_738_n N_A_2102_25#_c_1397_n 0.00208039f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_691 N_RESET_B_M1029_g N_A_2102_25#_c_1399_n 0.00311182f $X=12.39 $Y=0.465
+ $X2=0 $Y2=0
cc_692 N_RESET_B_c_745_n N_A_2102_25#_c_1399_n 0.00180239f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_693 N_RESET_B_c_746_n N_A_2102_25#_c_1399_n 0.00581749f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_694 N_RESET_B_c_731_n N_A_1799_379#_M1008_g 0.0100364f $X=12.18 $Y=1.78 $X2=0
+ $Y2=0
cc_695 N_RESET_B_c_738_n N_A_1799_379#_M1008_g 8.35195e-19 $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_696 N_RESET_B_M1029_g N_A_1799_379#_M1030_g 0.0545632f $X=12.39 $Y=0.465
+ $X2=0 $Y2=0
cc_697 N_RESET_B_M1001_g N_A_1799_379#_M1020_g 0.0128166f $X=12.54 $Y=2.195
+ $X2=0 $Y2=0
cc_698 N_RESET_B_c_738_n N_A_1799_379#_c_1483_n 0.00903322f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_699 N_RESET_B_c_738_n N_A_1799_379#_c_1502_n 0.0163825f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_700 N_RESET_B_c_738_n N_A_1799_379#_c_1503_n 0.0123672f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_701 N_RESET_B_M1017_g N_A_1799_379#_c_1504_n 7.78845e-19 $X=12.18 $Y=2.195
+ $X2=0 $Y2=0
cc_702 N_RESET_B_c_738_n N_A_1799_379#_c_1504_n 0.0114715f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_703 N_RESET_B_M1017_g N_A_1799_379#_c_1505_n 4.73841e-19 $X=12.18 $Y=2.195
+ $X2=0 $Y2=0
cc_704 N_RESET_B_M1017_g N_A_1799_379#_c_1507_n 0.012033f $X=12.18 $Y=2.195
+ $X2=0 $Y2=0
cc_705 N_RESET_B_M1001_g N_A_1799_379#_c_1507_n 5.53453e-19 $X=12.54 $Y=2.195
+ $X2=0 $Y2=0
cc_706 N_RESET_B_c_731_n N_A_1799_379#_c_1508_n 2.06137e-19 $X=12.18 $Y=1.78
+ $X2=0 $Y2=0
cc_707 N_RESET_B_M1001_g N_A_1799_379#_c_1508_n 0.0147393f $X=12.54 $Y=2.195
+ $X2=0 $Y2=0
cc_708 RESET_B N_A_1799_379#_c_1508_n 7.55376e-19 $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_709 N_RESET_B_c_746_n N_A_1799_379#_c_1508_n 0.011242f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_710 N_RESET_B_M1017_g N_A_1799_379#_c_1509_n 0.00670355f $X=12.18 $Y=2.195
+ $X2=0 $Y2=0
cc_711 RESET_B N_A_1799_379#_c_1509_n 0.00179858f $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_712 N_RESET_B_c_746_n N_A_1799_379#_c_1509_n 0.0102051f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_713 N_RESET_B_c_731_n N_A_1799_379#_c_1484_n 6.24711e-19 $X=12.18 $Y=1.78
+ $X2=0 $Y2=0
cc_714 N_RESET_B_c_746_n N_A_1799_379#_c_1484_n 0.00486366f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_715 N_RESET_B_c_731_n N_A_1799_379#_c_1511_n 0.00110299f $X=12.18 $Y=1.78
+ $X2=0 $Y2=0
cc_716 N_RESET_B_c_746_n N_A_1799_379#_c_1511_n 5.27597e-19 $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_738_n N_A_1799_379#_c_1486_n 0.0039996f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_718 N_RESET_B_c_738_n N_A_1799_379#_c_1487_n 0.0508357f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_719 N_RESET_B_c_738_n N_A_1799_379#_c_1488_n 0.0134061f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_720 N_RESET_B_c_731_n N_A_1799_379#_c_1489_n 0.0128166f $X=12.18 $Y=1.78
+ $X2=0 $Y2=0
cc_721 N_RESET_B_c_745_n N_A_1799_379#_c_1489_n 0.00635794f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_722 N_RESET_B_c_746_n N_A_1799_379#_c_1489_n 2.36087e-19 $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_723 N_RESET_B_c_735_n N_A_1799_379#_c_1491_n 0.0100364f $X=12.36 $Y=1.63
+ $X2=0 $Y2=0
cc_724 N_RESET_B_c_738_n N_A_1799_379#_c_1491_n 0.00282327f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_725 N_RESET_B_M1029_g N_A_1799_379#_c_1492_n 0.00635794f $X=12.39 $Y=0.465
+ $X2=0 $Y2=0
cc_726 N_RESET_B_c_746_n N_A_1799_379#_c_1492_n 0.00239262f $X=12.29 $Y=1.275
+ $X2=0 $Y2=0
cc_727 N_RESET_B_M1014_g N_A_27_457#_c_1835_n 0.00331137f $X=0.91 $Y=2.495 $X2=0
+ $Y2=0
cc_728 N_RESET_B_M1014_g N_A_27_457#_c_1837_n 0.0035397f $X=0.91 $Y=2.495 $X2=0
+ $Y2=0
cc_729 N_RESET_B_M1022_g N_A_27_457#_c_1837_n 0.00722825f $X=1.27 $Y=2.495 $X2=0
+ $Y2=0
cc_730 N_RESET_B_M1022_g N_A_27_457#_c_1838_n 0.00787625f $X=1.27 $Y=2.495 $X2=0
+ $Y2=0
cc_731 N_RESET_B_M1022_g N_A_27_457#_c_1853_n 0.00144522f $X=1.27 $Y=2.495 $X2=0
+ $Y2=0
cc_732 N_RESET_B_M1014_g N_A_111_457#_c_1876_n 0.00987937f $X=0.91 $Y=2.495
+ $X2=0 $Y2=0
cc_733 N_RESET_B_M1022_g N_A_111_457#_c_1876_n 0.00121987f $X=1.27 $Y=2.495
+ $X2=0 $Y2=0
cc_734 N_RESET_B_c_722_n N_A_111_457#_c_1877_n 2.06387e-19 $X=0.91 $Y=1.78 $X2=0
+ $Y2=0
cc_735 N_RESET_B_M1014_g N_A_111_457#_c_1877_n 0.0144626f $X=0.91 $Y=2.495 $X2=0
+ $Y2=0
cc_736 N_RESET_B_M1022_g N_A_111_457#_c_1877_n 0.0105936f $X=1.27 $Y=2.495 $X2=0
+ $Y2=0
cc_737 N_RESET_B_c_736_n N_A_111_457#_c_1877_n 0.0374123f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_738 N_RESET_B_c_737_n N_A_111_457#_c_1877_n 0.00313483f $X=1.345 $Y=1.665
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_743_n N_A_111_457#_c_1877_n 0.0204463f $X=1.15 $Y=1.275 $X2=0
+ $Y2=0
cc_740 N_RESET_B_M1014_g N_A_111_457#_c_1878_n 0.00513266f $X=0.91 $Y=2.495
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_726_n N_A_111_457#_c_1875_n 0.00450832f $X=4.475 $Y=0.165
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_736_n N_A_111_457#_c_1875_n 0.0416127f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_736_n N_A_111_457#_c_1883_n 0.00212706f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_736_n N_A_111_457#_c_1884_n 0.00742132f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_745 N_RESET_B_M1022_g N_VPWR_c_1951_n 0.00158668f $X=1.27 $Y=2.495 $X2=0
+ $Y2=0
cc_746 N_RESET_B_c_750_n N_VPWR_c_1952_n 0.00377627f $X=5.11 $Y=2.16 $X2=0 $Y2=0
cc_747 N_RESET_B_M1022_g N_VPWR_c_1950_n 8.57651e-19 $X=1.27 $Y=2.495 $X2=0
+ $Y2=0
cc_748 N_RESET_B_c_750_n N_VPWR_c_1950_n 9.49986e-19 $X=5.11 $Y=2.16 $X2=0 $Y2=0
cc_749 N_RESET_B_c_751_n N_VPWR_c_1950_n 9.49986e-19 $X=5.47 $Y=2.16 $X2=0 $Y2=0
cc_750 N_RESET_B_c_736_n N_A_484_411#_c_2103_n 7.91953e-19 $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_751 N_RESET_B_c_738_n N_A_1712_379#_c_2146_n 0.00666504f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_752 N_RESET_B_M1017_g N_A_2185_397#_c_2174_n 6.65587e-19 $X=12.18 $Y=2.195
+ $X2=0 $Y2=0
cc_753 N_RESET_B_M1001_g N_A_2185_397#_c_2176_n 0.00474054f $X=12.54 $Y=2.195
+ $X2=0 $Y2=0
cc_754 N_RESET_B_M1017_g N_A_2185_397#_c_2178_n 2.01539e-19 $X=12.18 $Y=2.195
+ $X2=0 $Y2=0
cc_755 N_RESET_B_M1001_g N_A_2185_397#_c_2178_n 0.00736212f $X=12.54 $Y=2.195
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_738_n N_A_2185_397#_c_2180_n 0.00854816f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_724_n N_VGND_c_2266_n 0.0044143f $X=1.345 $Y=1.185 $X2=0
+ $Y2=0
cc_758 N_RESET_B_M1033_g N_VGND_c_2266_n 0.00332485f $X=1.67 $Y=0.79 $X2=0 $Y2=0
cc_759 N_RESET_B_c_727_n N_VGND_c_2266_n 0.0113998f $X=1.745 $Y=0.165 $X2=0
+ $Y2=0
cc_760 N_RESET_B_c_737_n N_VGND_c_2266_n 9.47191e-19 $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_761 N_RESET_B_c_743_n N_VGND_c_2266_n 0.0221154f $X=1.15 $Y=1.275 $X2=0 $Y2=0
cc_762 N_RESET_B_c_726_n N_VGND_c_2267_n 0.0186759f $X=4.475 $Y=0.165 $X2=0
+ $Y2=0
cc_763 N_RESET_B_c_727_n N_VGND_c_2274_n 0.0838569f $X=1.745 $Y=0.165 $X2=0
+ $Y2=0
cc_764 N_RESET_B_M1029_g N_VGND_c_2276_n 0.00346682f $X=12.39 $Y=0.465 $X2=0
+ $Y2=0
cc_765 N_RESET_B_M1033_g N_VGND_c_2279_n 0.00157289f $X=1.67 $Y=0.79 $X2=0 $Y2=0
cc_766 N_RESET_B_c_726_n N_VGND_c_2279_n 0.0616494f $X=4.475 $Y=0.165 $X2=0
+ $Y2=0
cc_767 N_RESET_B_c_727_n N_VGND_c_2279_n 0.00479547f $X=1.745 $Y=0.165 $X2=0
+ $Y2=0
cc_768 N_RESET_B_M1040_g N_VGND_c_2279_n 0.00227535f $X=4.55 $Y=0.79 $X2=0 $Y2=0
cc_769 N_RESET_B_M1029_g N_VGND_c_2279_n 0.0063336f $X=12.39 $Y=0.465 $X2=0
+ $Y2=0
cc_770 N_A_590_116#_c_980_n N_A_560_90#_M1016_g 0.00517136f $X=3.25 $Y=1.685
+ $X2=0 $Y2=0
cc_771 N_A_590_116#_c_995_n N_A_560_90#_M1016_g 9.29005e-19 $X=3.25 $Y=1.77
+ $X2=0 $Y2=0
cc_772 N_A_590_116#_M1000_g N_A_560_90#_c_1168_n 0.00895007f $X=6.43 $Y=2.285
+ $X2=0 $Y2=0
cc_773 N_A_590_116#_M1007_g N_A_560_90#_c_1168_n 0.00894529f $X=6.79 $Y=2.285
+ $X2=0 $Y2=0
cc_774 N_A_590_116#_c_1056_n N_A_560_90#_c_1168_n 0.00709457f $X=5.52 $Y=2.395
+ $X2=0 $Y2=0
cc_775 N_A_590_116#_c_994_n N_A_560_90#_c_1168_n 3.24108e-19 $X=4.195 $Y=2.395
+ $X2=0 $Y2=0
cc_776 N_A_590_116#_c_997_n N_A_560_90#_c_1168_n 0.00589415f $X=5.685 $Y=2.395
+ $X2=0 $Y2=0
cc_777 N_A_590_116#_c_976_n N_A_560_90#_M1006_g 0.017821f $X=6.79 $Y=1.1 $X2=0
+ $Y2=0
cc_778 N_A_590_116#_c_990_n N_A_560_90#_c_1175_n 0.00171395f $X=3.25 $Y=2.2
+ $X2=0 $Y2=0
cc_779 N_A_590_116#_c_995_n N_A_560_90#_c_1175_n 7.28133e-19 $X=3.25 $Y=1.77
+ $X2=0 $Y2=0
cc_780 N_A_590_116#_M1007_g N_A_560_90#_c_1156_n 0.0457799f $X=6.79 $Y=2.285
+ $X2=0 $Y2=0
cc_781 N_A_590_116#_c_980_n N_A_111_457#_c_1875_n 0.0294957f $X=3.25 $Y=1.685
+ $X2=0 $Y2=0
cc_782 N_A_590_116#_c_990_n N_A_111_457#_c_1875_n 0.00471231f $X=3.25 $Y=2.2
+ $X2=0 $Y2=0
cc_783 N_A_590_116#_c_995_n N_A_111_457#_c_1875_n 0.00766544f $X=3.25 $Y=1.77
+ $X2=0 $Y2=0
cc_784 N_A_590_116#_c_990_n N_A_111_457#_c_1881_n 0.013238f $X=3.25 $Y=2.2 $X2=0
+ $Y2=0
cc_785 N_A_590_116#_c_990_n N_A_111_457#_c_1883_n 0.0125142f $X=3.25 $Y=2.2
+ $X2=0 $Y2=0
cc_786 N_A_590_116#_c_991_n N_A_111_457#_c_1883_n 0.0241864f $X=4.025 $Y=1.77
+ $X2=0 $Y2=0
cc_787 N_A_590_116#_c_993_n N_A_111_457#_c_1883_n 0.0209061f $X=4.11 $Y=2.31
+ $X2=0 $Y2=0
cc_788 N_A_590_116#_c_994_n N_A_111_457#_c_1883_n 0.0144409f $X=4.195 $Y=2.395
+ $X2=0 $Y2=0
cc_789 N_A_590_116#_c_990_n N_A_111_457#_c_1884_n 0.0102485f $X=3.25 $Y=2.2
+ $X2=0 $Y2=0
cc_790 N_A_590_116#_c_1056_n N_VPWR_M1002_d 0.00669362f $X=5.52 $Y=2.395 $X2=0
+ $Y2=0
cc_791 N_A_590_116#_c_1056_n N_VPWR_c_1952_n 0.0232582f $X=5.52 $Y=2.395 $X2=0
+ $Y2=0
cc_792 N_A_590_116#_c_997_n N_VPWR_c_1952_n 0.0013162f $X=5.685 $Y=2.395 $X2=0
+ $Y2=0
cc_793 N_A_590_116#_M1000_g N_VPWR_c_1953_n 0.00144992f $X=6.43 $Y=2.285 $X2=0
+ $Y2=0
cc_794 N_A_590_116#_M1007_g N_VPWR_c_1953_n 0.00939796f $X=6.79 $Y=2.285 $X2=0
+ $Y2=0
cc_795 N_A_590_116#_c_997_n N_VPWR_c_1965_n 0.00675783f $X=5.685 $Y=2.395 $X2=0
+ $Y2=0
cc_796 N_A_590_116#_M1000_g N_VPWR_c_1950_n 9.49986e-19 $X=6.43 $Y=2.285 $X2=0
+ $Y2=0
cc_797 N_A_590_116#_M1007_g N_VPWR_c_1950_n 7.97988e-19 $X=6.79 $Y=2.285 $X2=0
+ $Y2=0
cc_798 N_A_590_116#_c_1056_n N_VPWR_c_1950_n 0.0245291f $X=5.52 $Y=2.395 $X2=0
+ $Y2=0
cc_799 N_A_590_116#_c_994_n N_VPWR_c_1950_n 4.1868e-19 $X=4.195 $Y=2.395 $X2=0
+ $Y2=0
cc_800 N_A_590_116#_c_997_n N_VPWR_c_1950_n 0.00863128f $X=5.685 $Y=2.395 $X2=0
+ $Y2=0
cc_801 N_A_590_116#_c_993_n N_A_484_411#_M1002_s 4.45484e-19 $X=4.11 $Y=2.31
+ $X2=0 $Y2=0
cc_802 N_A_590_116#_c_1056_n N_A_484_411#_M1002_s 0.00669033f $X=5.52 $Y=2.395
+ $X2=0 $Y2=0
cc_803 N_A_590_116#_c_994_n N_A_484_411#_M1002_s 0.00214712f $X=4.195 $Y=2.395
+ $X2=0 $Y2=0
cc_804 N_A_590_116#_c_994_n N_A_484_411#_c_2104_n 0.00113153f $X=4.195 $Y=2.395
+ $X2=0 $Y2=0
cc_805 N_A_590_116#_c_1056_n N_A_484_411#_c_2106_n 0.0137311f $X=5.52 $Y=2.395
+ $X2=0 $Y2=0
cc_806 N_A_590_116#_c_994_n N_A_484_411#_c_2106_n 0.0112858f $X=4.195 $Y=2.395
+ $X2=0 $Y2=0
cc_807 N_A_590_116#_c_1056_n A_1037_457# 0.00181171f $X=5.52 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_808 N_A_590_116#_c_973_n N_VGND_c_2268_n 0.00298528f $X=6.43 $Y=1.1 $X2=0
+ $Y2=0
cc_809 N_A_590_116#_c_976_n N_VGND_c_2268_n 0.00471573f $X=6.79 $Y=1.1 $X2=0
+ $Y2=0
cc_810 N_A_590_116#_c_976_n N_VGND_c_2269_n 0.00942511f $X=6.79 $Y=1.1 $X2=0
+ $Y2=0
cc_811 N_A_590_116#_c_984_n N_VGND_c_2274_n 0.00639703f $X=3.17 $Y=0.79 $X2=0
+ $Y2=0
cc_812 N_A_590_116#_c_973_n N_VGND_c_2279_n 0.00450802f $X=6.43 $Y=1.1 $X2=0
+ $Y2=0
cc_813 N_A_590_116#_c_976_n N_VGND_c_2279_n 0.00941271f $X=6.79 $Y=1.1 $X2=0
+ $Y2=0
cc_814 N_A_590_116#_c_984_n N_VGND_c_2279_n 0.0102233f $X=3.17 $Y=0.79 $X2=0
+ $Y2=0
cc_815 N_A_560_90#_c_1161_n N_A_2102_25#_M1030_d 0.008727f $X=13.67 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_816 N_A_560_90#_M1036_g N_A_2102_25#_M1032_g 0.0203357f $X=9.925 $Y=0.465
+ $X2=0 $Y2=0
cc_817 N_A_560_90#_c_1157_n N_A_2102_25#_M1032_g 0.00423181f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_818 N_A_560_90#_c_1159_n N_A_2102_25#_M1032_g 0.0146937f $X=11.145 $Y=0.75
+ $X2=0 $Y2=0
cc_819 N_A_560_90#_c_1246_p N_A_2102_25#_M1032_g 0.00307933f $X=11.23 $Y=0.665
+ $X2=0 $Y2=0
cc_820 N_A_560_90#_c_1159_n N_A_2102_25#_c_1392_n 0.0356122f $X=11.145 $Y=0.75
+ $X2=0 $Y2=0
cc_821 N_A_560_90#_c_1161_n N_A_2102_25#_c_1392_n 0.0137373f $X=13.67 $Y=0.35
+ $X2=0 $Y2=0
cc_822 N_A_560_90#_c_1159_n N_A_2102_25#_c_1395_n 0.00804833f $X=11.145 $Y=0.75
+ $X2=0 $Y2=0
cc_823 N_A_560_90#_c_1246_p N_A_2102_25#_c_1395_n 0.00196023f $X=11.23 $Y=0.665
+ $X2=0 $Y2=0
cc_824 N_A_560_90#_c_1161_n N_A_2102_25#_c_1395_n 0.0123465f $X=13.67 $Y=0.35
+ $X2=0 $Y2=0
cc_825 N_A_560_90#_c_1161_n N_A_2102_25#_c_1396_n 0.073214f $X=13.67 $Y=0.35
+ $X2=0 $Y2=0
cc_826 N_A_560_90#_c_1162_n N_A_2102_25#_c_1396_n 0.00559569f $X=13.835 $Y=0.47
+ $X2=0 $Y2=0
cc_827 N_A_560_90#_c_1164_n N_A_2102_25#_c_1396_n 0.00697863f $X=14 $Y=0.815
+ $X2=0 $Y2=0
cc_828 N_A_560_90#_c_1157_n N_A_2102_25#_c_1397_n 0.0188003f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_829 N_A_560_90#_c_1158_n N_A_2102_25#_c_1397_n 0.00127159f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_830 N_A_560_90#_c_1159_n N_A_2102_25#_c_1397_n 0.0231602f $X=11.145 $Y=0.75
+ $X2=0 $Y2=0
cc_831 N_A_560_90#_c_1157_n N_A_2102_25#_c_1398_n 0.00121489f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_832 N_A_560_90#_c_1158_n N_A_2102_25#_c_1398_n 0.0292051f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_833 N_A_560_90#_c_1159_n N_A_2102_25#_c_1398_n 0.00124625f $X=11.145 $Y=0.75
+ $X2=0 $Y2=0
cc_834 N_A_560_90#_c_1161_n N_A_1799_379#_M1030_g 0.0115366f $X=13.67 $Y=0.35
+ $X2=0 $Y2=0
cc_835 N_A_560_90#_c_1179_n N_A_1799_379#_M1020_g 0.0055018f $X=13.865 $Y=2.11
+ $X2=0 $Y2=0
cc_836 N_A_560_90#_c_1180_n N_A_1799_379#_M1020_g 9.08881e-19 $X=14.03 $Y=2.025
+ $X2=0 $Y2=0
cc_837 N_A_560_90#_c_1163_n N_A_1799_379#_M1050_g 0.0160571f $X=15.165 $Y=0.815
+ $X2=0 $Y2=0
cc_838 N_A_560_90#_c_1165_n N_A_1799_379#_M1050_g 0.0112665f $X=15.25 $Y=1.94
+ $X2=0 $Y2=0
cc_839 N_A_560_90#_c_1266_p N_A_1799_379#_M1031_g 0.0185008f $X=15.165 $Y=2.025
+ $X2=0 $Y2=0
cc_840 N_A_560_90#_c_1165_n N_A_1799_379#_M1031_g 0.00587259f $X=15.25 $Y=1.94
+ $X2=0 $Y2=0
cc_841 N_A_560_90#_c_1165_n N_A_1799_379#_c_1470_n 0.00567731f $X=15.25 $Y=1.94
+ $X2=0 $Y2=0
cc_842 N_A_560_90#_c_1165_n N_A_1799_379#_M1035_g 0.00221686f $X=15.25 $Y=1.94
+ $X2=0 $Y2=0
cc_843 N_A_560_90#_c_1165_n N_A_1799_379#_M1011_g 0.00243642f $X=15.25 $Y=1.94
+ $X2=0 $Y2=0
cc_844 N_A_560_90#_c_1173_n N_A_1799_379#_c_1500_n 0.00442153f $X=9.38 $Y=2.92
+ $X2=0 $Y2=0
cc_845 N_A_560_90#_M1044_g N_A_1799_379#_c_1500_n 0.0164744f $X=9.455 $Y=2.315
+ $X2=0 $Y2=0
cc_846 N_A_560_90#_c_1153_n N_A_1799_379#_c_1482_n 0.0154056f $X=9.85 $Y=1.45
+ $X2=0 $Y2=0
cc_847 N_A_560_90#_c_1154_n N_A_1799_379#_c_1482_n 0.00445569f $X=9.53 $Y=1.45
+ $X2=0 $Y2=0
cc_848 N_A_560_90#_M1036_g N_A_1799_379#_c_1482_n 0.0219728f $X=9.925 $Y=0.465
+ $X2=0 $Y2=0
cc_849 N_A_560_90#_c_1157_n N_A_1799_379#_c_1482_n 0.0385881f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_850 N_A_560_90#_c_1160_n N_A_1799_379#_c_1482_n 0.0136434f $X=10.27 $Y=0.75
+ $X2=0 $Y2=0
cc_851 N_A_560_90#_c_1153_n N_A_1799_379#_c_1483_n 0.00789993f $X=9.85 $Y=1.45
+ $X2=0 $Y2=0
cc_852 N_A_560_90#_M1044_g N_A_1799_379#_c_1502_n 0.00710949f $X=9.455 $Y=2.315
+ $X2=0 $Y2=0
cc_853 N_A_560_90#_c_1153_n N_A_1799_379#_c_1502_n 0.0039834f $X=9.85 $Y=1.45
+ $X2=0 $Y2=0
cc_854 N_A_560_90#_M1044_g N_A_1799_379#_c_1503_n 0.00942f $X=9.455 $Y=2.315
+ $X2=0 $Y2=0
cc_855 N_A_560_90#_c_1179_n N_A_1799_379#_c_1508_n 0.00108915f $X=13.865 $Y=2.11
+ $X2=0 $Y2=0
cc_856 N_A_560_90#_c_1180_n N_A_1799_379#_c_1508_n 0.00884281f $X=14.03 $Y=2.025
+ $X2=0 $Y2=0
cc_857 N_A_560_90#_c_1180_n N_A_1799_379#_c_1511_n 0.00108914f $X=14.03 $Y=2.025
+ $X2=0 $Y2=0
cc_858 N_A_560_90#_c_1266_p N_A_1799_379#_c_1485_n 0.0416276f $X=15.165 $Y=2.025
+ $X2=0 $Y2=0
cc_859 N_A_560_90#_c_1180_n N_A_1799_379#_c_1485_n 0.0232639f $X=14.03 $Y=2.025
+ $X2=0 $Y2=0
cc_860 N_A_560_90#_c_1157_n N_A_1799_379#_c_1486_n 0.0121176f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_861 N_A_560_90#_c_1158_n N_A_1799_379#_c_1486_n 0.00564516f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_862 N_A_560_90#_c_1157_n N_A_1799_379#_c_1487_n 0.0113682f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_863 N_A_560_90#_c_1158_n N_A_1799_379#_c_1487_n 0.00499545f $X=10.105 $Y=1.18
+ $X2=0 $Y2=0
cc_864 N_A_560_90#_c_1163_n N_A_1799_379#_c_1490_n 0.00910984f $X=15.165
+ $Y=0.815 $X2=0 $Y2=0
cc_865 N_A_560_90#_c_1266_p N_A_1799_379#_c_1490_n 0.0193636f $X=15.165 $Y=2.025
+ $X2=0 $Y2=0
cc_866 N_A_560_90#_c_1165_n N_A_1799_379#_c_1490_n 0.0280814f $X=15.25 $Y=1.94
+ $X2=0 $Y2=0
cc_867 N_A_560_90#_c_1163_n N_A_1799_379#_c_1493_n 0.00142334f $X=15.165
+ $Y=0.815 $X2=0 $Y2=0
cc_868 N_A_560_90#_c_1266_p N_A_1799_379#_c_1493_n 0.00142518f $X=15.165
+ $Y=2.025 $X2=0 $Y2=0
cc_869 N_A_560_90#_c_1165_n N_A_1799_379#_c_1493_n 0.00599399f $X=15.25 $Y=1.94
+ $X2=0 $Y2=0
cc_870 N_A_560_90#_c_1161_n N_CLK_M1026_g 0.00329161f $X=13.67 $Y=0.35 $X2=0
+ $Y2=0
cc_871 N_A_560_90#_c_1162_n N_CLK_M1026_g 0.00643775f $X=13.835 $Y=0.47 $X2=0
+ $Y2=0
cc_872 N_A_560_90#_c_1163_n N_CLK_M1026_g 0.00855199f $X=15.165 $Y=0.815 $X2=0
+ $Y2=0
cc_873 N_A_560_90#_c_1164_n N_CLK_M1026_g 0.00420699f $X=14 $Y=0.815 $X2=0 $Y2=0
cc_874 N_A_560_90#_c_1179_n N_CLK_M1049_g 0.00884829f $X=13.865 $Y=2.11 $X2=0
+ $Y2=0
cc_875 N_A_560_90#_c_1266_p N_CLK_M1049_g 0.0104168f $X=15.165 $Y=2.025 $X2=0
+ $Y2=0
cc_876 N_A_560_90#_c_1180_n N_CLK_M1049_g 0.00236324f $X=14.03 $Y=2.025 $X2=0
+ $Y2=0
cc_877 N_A_560_90#_c_1163_n N_CLK_c_1717_n 0.00135471f $X=15.165 $Y=0.815 $X2=0
+ $Y2=0
cc_878 N_A_560_90#_c_1161_n N_CLK_M1027_g 4.79243e-19 $X=13.67 $Y=0.35 $X2=0
+ $Y2=0
cc_879 N_A_560_90#_c_1162_n N_CLK_M1027_g 0.001214f $X=13.835 $Y=0.47 $X2=0
+ $Y2=0
cc_880 N_A_560_90#_c_1163_n N_CLK_M1027_g 0.0172311f $X=15.165 $Y=0.815 $X2=0
+ $Y2=0
cc_881 N_A_560_90#_c_1165_n N_CLK_M1027_g 0.00209787f $X=15.25 $Y=1.94 $X2=0
+ $Y2=0
cc_882 N_A_560_90#_c_1179_n N_CLK_M1034_g 0.00192788f $X=13.865 $Y=2.11 $X2=0
+ $Y2=0
cc_883 N_A_560_90#_c_1266_p N_CLK_M1034_g 0.0152533f $X=15.165 $Y=2.025 $X2=0
+ $Y2=0
cc_884 N_A_560_90#_c_1165_n N_CLK_M1034_g 7.73481e-19 $X=15.25 $Y=1.94 $X2=0
+ $Y2=0
cc_885 N_A_560_90#_c_1161_n CLK 0.00327049f $X=13.67 $Y=0.35 $X2=0 $Y2=0
cc_886 N_A_560_90#_c_1163_n CLK 0.0192582f $X=15.165 $Y=0.815 $X2=0 $Y2=0
cc_887 N_A_560_90#_c_1164_n CLK 0.0270393f $X=14 $Y=0.815 $X2=0 $Y2=0
cc_888 N_A_560_90#_c_1164_n N_CLK_c_1722_n 0.00346378f $X=14 $Y=0.815 $X2=0
+ $Y2=0
cc_889 N_A_560_90#_M1016_g N_A_111_457#_c_1875_n 0.0285394f $X=2.875 $Y=0.79
+ $X2=0 $Y2=0
cc_890 N_A_560_90#_M1024_g N_A_111_457#_c_1875_n 3.171e-19 $X=3.035 $Y=2.265
+ $X2=0 $Y2=0
cc_891 N_A_560_90#_c_1175_n N_A_111_457#_c_1875_n 0.00614852f $X=3.035 $Y=1.87
+ $X2=0 $Y2=0
cc_892 N_A_560_90#_M1024_g N_A_111_457#_c_1880_n 0.0126979f $X=3.035 $Y=2.265
+ $X2=0 $Y2=0
cc_893 N_A_560_90#_M1024_g N_A_111_457#_c_1881_n 0.0124836f $X=3.035 $Y=2.265
+ $X2=0 $Y2=0
cc_894 N_A_560_90#_M1024_g N_A_111_457#_c_1882_n 0.00370163f $X=3.035 $Y=2.265
+ $X2=0 $Y2=0
cc_895 N_A_560_90#_M1024_g N_A_111_457#_c_1883_n 5.62766e-19 $X=3.035 $Y=2.265
+ $X2=0 $Y2=0
cc_896 N_A_560_90#_M1024_g N_A_111_457#_c_1884_n 0.00629865f $X=3.035 $Y=2.265
+ $X2=0 $Y2=0
cc_897 N_A_560_90#_c_1175_n N_A_111_457#_c_1884_n 0.00765319f $X=3.035 $Y=1.87
+ $X2=0 $Y2=0
cc_898 N_A_560_90#_c_1266_p N_VPWR_M1034_d 0.0135886f $X=15.165 $Y=2.025 $X2=0
+ $Y2=0
cc_899 N_A_560_90#_c_1168_n N_VPWR_c_1952_n 0.0253641f $X=7.25 $Y=3.15 $X2=0
+ $Y2=0
cc_900 N_A_560_90#_c_1168_n N_VPWR_c_1953_n 0.0250044f $X=7.25 $Y=3.15 $X2=0
+ $Y2=0
cc_901 N_A_560_90#_M1039_g N_VPWR_c_1953_n 0.0233116f $X=7.325 $Y=2.385 $X2=0
+ $Y2=0
cc_902 N_A_560_90#_c_1266_p N_VPWR_c_1956_n 0.0210122f $X=15.165 $Y=2.025 $X2=0
+ $Y2=0
cc_903 N_A_560_90#_c_1169_n N_VPWR_c_1958_n 0.0394739f $X=3.11 $Y=3.15 $X2=0
+ $Y2=0
cc_904 N_A_560_90#_c_1168_n N_VPWR_c_1965_n 0.0580539f $X=7.25 $Y=3.15 $X2=0
+ $Y2=0
cc_905 N_A_560_90#_c_1168_n N_VPWR_c_1966_n 0.00893687f $X=7.25 $Y=3.15 $X2=0
+ $Y2=0
cc_906 N_A_560_90#_c_1171_n N_VPWR_c_1966_n 0.0361119f $X=7.61 $Y=2.92 $X2=0
+ $Y2=0
cc_907 N_A_560_90#_c_1173_n N_VPWR_c_1966_n 0.00487243f $X=9.38 $Y=2.92 $X2=0
+ $Y2=0
cc_908 N_A_560_90#_c_1168_n N_VPWR_c_1950_n 0.105653f $X=7.25 $Y=3.15 $X2=0
+ $Y2=0
cc_909 N_A_560_90#_c_1169_n N_VPWR_c_1950_n 0.00604685f $X=3.11 $Y=3.15 $X2=0
+ $Y2=0
cc_910 N_A_560_90#_c_1171_n N_VPWR_c_1950_n 0.0363254f $X=7.61 $Y=2.92 $X2=0
+ $Y2=0
cc_911 N_A_560_90#_c_1177_n N_VPWR_c_1950_n 0.0115521f $X=7.325 $Y=2.92 $X2=0
+ $Y2=0
cc_912 N_A_560_90#_c_1179_n N_VPWR_c_1950_n 0.012638f $X=13.865 $Y=2.11 $X2=0
+ $Y2=0
cc_913 N_A_560_90#_M1024_g N_A_484_411#_c_2103_n 0.00754787f $X=3.035 $Y=2.265
+ $X2=0 $Y2=0
cc_914 N_A_560_90#_M1024_g N_A_484_411#_c_2104_n 0.0137753f $X=3.035 $Y=2.265
+ $X2=0 $Y2=0
cc_915 N_A_560_90#_c_1168_n N_A_484_411#_c_2104_n 0.01802f $X=7.25 $Y=3.15 $X2=0
+ $Y2=0
cc_916 N_A_560_90#_c_1168_n N_A_484_411#_c_2106_n 0.00789901f $X=7.25 $Y=3.15
+ $X2=0 $Y2=0
cc_917 N_A_560_90#_c_1173_n N_A_1712_379#_c_2146_n 0.0113632f $X=9.38 $Y=2.92
+ $X2=0 $Y2=0
cc_918 N_A_560_90#_M1044_g N_A_1712_379#_c_2146_n 0.00403939f $X=9.455 $Y=2.315
+ $X2=0 $Y2=0
cc_919 N_A_560_90#_c_1173_n N_A_1712_379#_c_2147_n 0.0284648f $X=9.38 $Y=2.92
+ $X2=0 $Y2=0
cc_920 N_A_560_90#_c_1173_n N_A_1712_379#_c_2148_n 0.0114268f $X=9.38 $Y=2.92
+ $X2=0 $Y2=0
cc_921 N_A_560_90#_c_1179_n N_A_2185_397#_c_2177_n 0.0131777f $X=13.865 $Y=2.11
+ $X2=0 $Y2=0
cc_922 N_A_560_90#_c_1179_n N_A_2185_397#_c_2179_n 0.00105883f $X=13.865 $Y=2.11
+ $X2=0 $Y2=0
cc_923 N_A_560_90#_c_1266_p A_2831_367# 0.00471068f $X=15.165 $Y=2.025 $X2=-0.19
+ $Y2=-0.245
cc_924 N_A_560_90#_c_1266_p A_3036_367# 0.00433061f $X=15.165 $Y=2.025 $X2=-0.19
+ $Y2=-0.245
cc_925 N_A_560_90#_c_1165_n N_Q_N_c_2228_n 0.0638485f $X=15.25 $Y=1.94 $X2=0
+ $Y2=0
cc_926 N_A_560_90#_c_1159_n N_VGND_M1032_d 0.00624466f $X=11.145 $Y=0.75 $X2=0
+ $Y2=0
cc_927 N_A_560_90#_c_1246_p N_VGND_M1032_d 0.0129791f $X=11.23 $Y=0.665 $X2=0
+ $Y2=0
cc_928 N_A_560_90#_c_1161_n N_VGND_M1032_d 0.0306952f $X=13.67 $Y=0.35 $X2=0
+ $Y2=0
cc_929 N_A_560_90#_c_1356_p N_VGND_M1032_d 0.00499578f $X=11.315 $Y=0.35 $X2=0
+ $Y2=0
cc_930 N_A_560_90#_c_1163_n N_VGND_M1027_d 0.00673723f $X=15.165 $Y=0.815 $X2=0
+ $Y2=0
cc_931 N_A_560_90#_M1006_g N_VGND_c_2269_n 0.00980526f $X=7.405 $Y=0.765 $X2=0
+ $Y2=0
cc_932 N_A_560_90#_M1036_g N_VGND_c_2270_n 0.00171477f $X=9.925 $Y=0.465 $X2=0
+ $Y2=0
cc_933 N_A_560_90#_c_1159_n N_VGND_c_2270_n 0.0196682f $X=11.145 $Y=0.75 $X2=0
+ $Y2=0
cc_934 N_A_560_90#_c_1246_p N_VGND_c_2270_n 0.00362732f $X=11.23 $Y=0.665 $X2=0
+ $Y2=0
cc_935 N_A_560_90#_c_1356_p N_VGND_c_2270_n 0.0138719f $X=11.315 $Y=0.35 $X2=0
+ $Y2=0
cc_936 N_A_560_90#_c_1161_n N_VGND_c_2271_n 0.00571183f $X=13.67 $Y=0.35 $X2=0
+ $Y2=0
cc_937 N_A_560_90#_c_1162_n N_VGND_c_2271_n 0.00362744f $X=13.835 $Y=0.47 $X2=0
+ $Y2=0
cc_938 N_A_560_90#_c_1163_n N_VGND_c_2271_n 0.0221947f $X=15.165 $Y=0.815 $X2=0
+ $Y2=0
cc_939 N_A_560_90#_M1006_g N_VGND_c_2275_n 0.00454183f $X=7.405 $Y=0.765 $X2=0
+ $Y2=0
cc_940 N_A_560_90#_M1041_g N_VGND_c_2275_n 0.00436277f $X=7.765 $Y=0.765 $X2=0
+ $Y2=0
cc_941 N_A_560_90#_M1036_g N_VGND_c_2275_n 0.00504125f $X=9.925 $Y=0.465 $X2=0
+ $Y2=0
cc_942 N_A_560_90#_c_1159_n N_VGND_c_2275_n 0.00539949f $X=11.145 $Y=0.75 $X2=0
+ $Y2=0
cc_943 N_A_560_90#_c_1160_n N_VGND_c_2275_n 0.00537453f $X=10.27 $Y=0.75 $X2=0
+ $Y2=0
cc_944 N_A_560_90#_c_1159_n N_VGND_c_2276_n 0.00292892f $X=11.145 $Y=0.75 $X2=0
+ $Y2=0
cc_945 N_A_560_90#_c_1161_n N_VGND_c_2276_n 0.154035f $X=13.67 $Y=0.35 $X2=0
+ $Y2=0
cc_946 N_A_560_90#_c_1356_p N_VGND_c_2276_n 0.011088f $X=11.315 $Y=0.35 $X2=0
+ $Y2=0
cc_947 N_A_560_90#_c_1163_n N_VGND_c_2276_n 0.00690612f $X=15.165 $Y=0.815 $X2=0
+ $Y2=0
cc_948 N_A_560_90#_c_1163_n N_VGND_c_2277_n 0.0065908f $X=15.165 $Y=0.815 $X2=0
+ $Y2=0
cc_949 N_A_560_90#_M1026_s N_VGND_c_2279_n 0.0023122f $X=13.69 $Y=0.24 $X2=0
+ $Y2=0
cc_950 N_A_560_90#_M1016_g N_VGND_c_2279_n 0.00264436f $X=2.875 $Y=0.79 $X2=0
+ $Y2=0
cc_951 N_A_560_90#_M1006_g N_VGND_c_2279_n 0.00489211f $X=7.405 $Y=0.765 $X2=0
+ $Y2=0
cc_952 N_A_560_90#_M1041_g N_VGND_c_2279_n 0.00489211f $X=7.765 $Y=0.765 $X2=0
+ $Y2=0
cc_953 N_A_560_90#_M1036_g N_VGND_c_2279_n 0.00950734f $X=9.925 $Y=0.465 $X2=0
+ $Y2=0
cc_954 N_A_560_90#_c_1159_n N_VGND_c_2279_n 0.0160668f $X=11.145 $Y=0.75 $X2=0
+ $Y2=0
cc_955 N_A_560_90#_c_1160_n N_VGND_c_2279_n 0.00948579f $X=10.27 $Y=0.75 $X2=0
+ $Y2=0
cc_956 N_A_560_90#_c_1161_n N_VGND_c_2279_n 0.0992618f $X=13.67 $Y=0.35 $X2=0
+ $Y2=0
cc_957 N_A_560_90#_c_1356_p N_VGND_c_2279_n 0.00654658f $X=11.315 $Y=0.35 $X2=0
+ $Y2=0
cc_958 N_A_560_90#_c_1163_n N_VGND_c_2279_n 0.0262856f $X=15.165 $Y=0.815 $X2=0
+ $Y2=0
cc_959 N_A_560_90#_c_1159_n A_2000_51# 0.00330762f $X=11.145 $Y=0.75 $X2=-0.19
+ $Y2=-0.245
cc_960 N_A_560_90#_c_1160_n A_2000_51# 0.00405433f $X=10.27 $Y=0.75 $X2=-0.19
+ $Y2=-0.245
cc_961 N_A_560_90#_c_1161_n A_2493_51# 0.00258465f $X=13.67 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_962 N_A_560_90#_c_1163_n A_3036_48# 0.00194172f $X=15.165 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_963 N_A_2102_25#_c_1396_n N_A_1799_379#_M1030_g 0.0196589f $X=13.11 $Y=0.7
+ $X2=0 $Y2=0
cc_964 N_A_2102_25#_c_1396_n N_A_1799_379#_c_1467_n 0.0148116f $X=13.11 $Y=0.7
+ $X2=0 $Y2=0
cc_965 N_A_2102_25#_M1013_g N_A_1799_379#_c_1500_n 0.00877897f $X=10.585
+ $Y=2.885 $X2=0 $Y2=0
cc_966 N_A_2102_25#_M1013_g N_A_1799_379#_c_1503_n 0.0180483f $X=10.585 $Y=2.885
+ $X2=0 $Y2=0
cc_967 N_A_2102_25#_c_1394_n N_A_1799_379#_c_1504_n 0.0450945f $X=11.85 $Y=2.165
+ $X2=0 $Y2=0
cc_968 N_A_2102_25#_c_1394_n N_A_1799_379#_c_1505_n 0.013324f $X=11.85 $Y=2.165
+ $X2=0 $Y2=0
cc_969 N_A_2102_25#_c_1394_n N_A_1799_379#_c_1507_n 0.0157539f $X=11.85 $Y=2.165
+ $X2=0 $Y2=0
cc_970 N_A_2102_25#_c_1394_n N_A_1799_379#_c_1509_n 0.0128131f $X=11.85 $Y=2.165
+ $X2=0 $Y2=0
cc_971 N_A_2102_25#_M1013_g N_A_1799_379#_c_1487_n 0.0152443f $X=10.585 $Y=2.885
+ $X2=0 $Y2=0
cc_972 N_A_2102_25#_c_1392_n N_A_1799_379#_c_1487_n 0.0147548f $X=11.765 $Y=1.1
+ $X2=0 $Y2=0
cc_973 N_A_2102_25#_c_1397_n N_A_1799_379#_c_1487_n 0.0211145f $X=10.675 $Y=1.1
+ $X2=0 $Y2=0
cc_974 N_A_2102_25#_c_1398_n N_A_1799_379#_c_1487_n 0.00124625f $X=10.675
+ $Y=1.18 $X2=0 $Y2=0
cc_975 N_A_2102_25#_M1013_g N_A_1799_379#_c_1488_n 8.19046e-19 $X=10.585
+ $Y=2.885 $X2=0 $Y2=0
cc_976 N_A_2102_25#_c_1392_n N_A_1799_379#_c_1488_n 0.0251609f $X=11.765 $Y=1.1
+ $X2=0 $Y2=0
cc_977 N_A_2102_25#_c_1394_n N_A_1799_379#_c_1488_n 0.0231991f $X=11.85 $Y=2.165
+ $X2=0 $Y2=0
cc_978 N_A_2102_25#_M1013_g N_A_1799_379#_c_1491_n 0.00534764f $X=10.585
+ $Y=2.885 $X2=0 $Y2=0
cc_979 N_A_2102_25#_c_1392_n N_A_1799_379#_c_1491_n 0.0091986f $X=11.765 $Y=1.1
+ $X2=0 $Y2=0
cc_980 N_A_2102_25#_c_1394_n N_A_1799_379#_c_1491_n 0.00804337f $X=11.85
+ $Y=2.165 $X2=0 $Y2=0
cc_981 N_A_2102_25#_c_1396_n N_CLK_M1026_g 9.97406e-19 $X=13.11 $Y=0.7 $X2=0
+ $Y2=0
cc_982 N_A_2102_25#_M1013_g N_VPWR_c_1954_n 0.0133978f $X=10.585 $Y=2.885 $X2=0
+ $Y2=0
cc_983 N_A_2102_25#_M1013_g N_VPWR_c_1966_n 0.00486043f $X=10.585 $Y=2.885 $X2=0
+ $Y2=0
cc_984 N_A_2102_25#_M1013_g N_VPWR_c_1950_n 0.00975473f $X=10.585 $Y=2.885 $X2=0
+ $Y2=0
cc_985 N_A_2102_25#_M1013_g N_A_1712_379#_c_2149_n 6.30273e-19 $X=10.585
+ $Y=2.885 $X2=0 $Y2=0
cc_986 N_A_2102_25#_M1013_g N_A_2185_397#_c_2173_n 0.0065793f $X=10.585 $Y=2.885
+ $X2=0 $Y2=0
cc_987 N_A_2102_25#_M1013_g N_A_2185_397#_c_2180_n 0.0157439f $X=10.585 $Y=2.885
+ $X2=0 $Y2=0
cc_988 N_A_2102_25#_c_1395_n N_VGND_M1032_d 0.00348367f $X=11.935 $Y=0.74 $X2=0
+ $Y2=0
cc_989 N_A_2102_25#_c_1396_n N_VGND_M1032_d 0.0040503f $X=13.11 $Y=0.7 $X2=0
+ $Y2=0
cc_990 N_A_2102_25#_M1032_g N_VGND_c_2270_n 0.0111895f $X=10.585 $Y=0.465 $X2=0
+ $Y2=0
cc_991 N_A_2102_25#_M1032_g N_VGND_c_2275_n 0.0034328f $X=10.585 $Y=0.465 $X2=0
+ $Y2=0
cc_992 N_A_2102_25#_M1032_g N_VGND_c_2279_n 0.00459614f $X=10.585 $Y=0.465 $X2=0
+ $Y2=0
cc_993 N_A_2102_25#_c_1396_n A_2493_51# 0.0013306f $X=13.11 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_994 N_A_1799_379#_c_1508_n N_CLK_M1049_g 5.27675e-19 $X=13.04 $Y=2.045 $X2=0
+ $Y2=0
cc_995 N_A_1799_379#_c_1511_n N_CLK_M1049_g 0.00131053f $X=13.205 $Y=1.96 $X2=0
+ $Y2=0
cc_996 N_A_1799_379#_c_1485_n N_CLK_M1049_g 0.0114367f $X=14.725 $Y=1.675 $X2=0
+ $Y2=0
cc_997 N_A_1799_379#_c_1489_n N_CLK_M1049_g 0.00535522f $X=13.205 $Y=1.755 $X2=0
+ $Y2=0
cc_998 N_A_1799_379#_M1050_g N_CLK_M1027_g 0.0242185f $X=15.105 $Y=0.66 $X2=0
+ $Y2=0
cc_999 N_A_1799_379#_M1031_g N_CLK_M1034_g 0.0159756f $X=15.105 $Y=2.465 $X2=0
+ $Y2=0
cc_1000 N_A_1799_379#_c_1485_n N_CLK_M1034_g 0.0145081f $X=14.725 $Y=1.675 $X2=0
+ $Y2=0
cc_1001 N_A_1799_379#_c_1490_n N_CLK_M1034_g 0.00162414f $X=14.89 $Y=1.51 $X2=0
+ $Y2=0
cc_1002 N_A_1799_379#_c_1493_n N_CLK_M1034_g 0.0218178f $X=15.18 $Y=1.51 $X2=0
+ $Y2=0
cc_1003 N_A_1799_379#_c_1485_n CLK 0.0521286f $X=14.725 $Y=1.675 $X2=0 $Y2=0
cc_1004 N_A_1799_379#_c_1490_n CLK 0.00257185f $X=14.89 $Y=1.51 $X2=0 $Y2=0
cc_1005 N_A_1799_379#_c_1492_n CLK 0.00788344f $X=13.205 $Y=1.59 $X2=0 $Y2=0
cc_1006 N_A_1799_379#_c_1485_n N_CLK_c_1722_n 0.00412671f $X=14.725 $Y=1.675
+ $X2=0 $Y2=0
cc_1007 N_A_1799_379#_c_1492_n N_CLK_c_1722_n 0.00396949f $X=13.205 $Y=1.59
+ $X2=0 $Y2=0
cc_1008 N_A_1799_379#_M1048_g N_A_3222_137#_M1015_g 0.0152262f $X=16.83 $Y=0.895
+ $X2=0 $Y2=0
cc_1009 N_A_1799_379#_M1025_g N_A_3222_137#_M1037_g 0.0166304f $X=16.83 $Y=2.155
+ $X2=0 $Y2=0
cc_1010 N_A_1799_379#_M1035_g N_A_3222_137#_c_1776_n 0.00178697f $X=15.465
+ $Y=0.66 $X2=0 $Y2=0
cc_1011 N_A_1799_379#_M1042_g N_A_3222_137#_c_1776_n 0.016733f $X=16.47 $Y=0.895
+ $X2=0 $Y2=0
cc_1012 N_A_1799_379#_M1048_g N_A_3222_137#_c_1776_n 0.00223078f $X=16.83
+ $Y=0.895 $X2=0 $Y2=0
cc_1013 N_A_1799_379#_M1011_g N_A_3222_137#_c_1782_n 0.00211777f $X=15.465
+ $Y=2.465 $X2=0 $Y2=0
cc_1014 N_A_1799_379#_M1028_g N_A_3222_137#_c_1782_n 0.0201599f $X=16.47
+ $Y=2.155 $X2=0 $Y2=0
cc_1015 N_A_1799_379#_M1025_g N_A_3222_137#_c_1782_n 0.0028674f $X=16.83
+ $Y=2.155 $X2=0 $Y2=0
cc_1016 N_A_1799_379#_M1042_g N_A_3222_137#_c_1777_n 0.00671173f $X=16.47
+ $Y=0.895 $X2=0 $Y2=0
cc_1017 N_A_1799_379#_M1028_g N_A_3222_137#_c_1777_n 0.00879129f $X=16.47
+ $Y=2.155 $X2=0 $Y2=0
cc_1018 N_A_1799_379#_c_1476_n N_A_3222_137#_c_1777_n 0.0038941f $X=16.755
+ $Y=1.42 $X2=0 $Y2=0
cc_1019 N_A_1799_379#_M1048_g N_A_3222_137#_c_1777_n 0.00859107f $X=16.83
+ $Y=0.895 $X2=0 $Y2=0
cc_1020 N_A_1799_379#_M1025_g N_A_3222_137#_c_1777_n 0.0123489f $X=16.83
+ $Y=2.155 $X2=0 $Y2=0
cc_1021 N_A_1799_379#_c_1480_n N_A_3222_137#_c_1777_n 0.00175146f $X=16.47
+ $Y=1.42 $X2=0 $Y2=0
cc_1022 N_A_1799_379#_c_1481_n N_A_3222_137#_c_1777_n 0.00434817f $X=16.83
+ $Y=1.42 $X2=0 $Y2=0
cc_1023 N_A_1799_379#_M1011_g N_A_3222_137#_c_1778_n 5.97095e-19 $X=15.465
+ $Y=2.465 $X2=0 $Y2=0
cc_1024 N_A_1799_379#_c_1473_n N_A_3222_137#_c_1778_n 0.0171919f $X=16.395
+ $Y=1.42 $X2=0 $Y2=0
cc_1025 N_A_1799_379#_M1042_g N_A_3222_137#_c_1778_n 8.79744e-19 $X=16.47
+ $Y=0.895 $X2=0 $Y2=0
cc_1026 N_A_1799_379#_M1028_g N_A_3222_137#_c_1778_n 0.0031355f $X=16.47
+ $Y=2.155 $X2=0 $Y2=0
cc_1027 N_A_1799_379#_c_1480_n N_A_3222_137#_c_1778_n 3.53117e-19 $X=16.47
+ $Y=1.42 $X2=0 $Y2=0
cc_1028 N_A_1799_379#_M1048_g N_A_3222_137#_c_1779_n 0.0103327f $X=16.83
+ $Y=0.895 $X2=0 $Y2=0
cc_1029 N_A_1799_379#_c_1508_n N_VPWR_M1001_d 0.00273362f $X=13.04 $Y=2.045
+ $X2=0 $Y2=0
cc_1030 N_A_1799_379#_M1020_g N_VPWR_c_1955_n 0.00462365f $X=13.115 $Y=2.76
+ $X2=0 $Y2=0
cc_1031 N_A_1799_379#_M1031_g N_VPWR_c_1956_n 0.0203993f $X=15.105 $Y=2.465
+ $X2=0 $Y2=0
cc_1032 N_A_1799_379#_M1011_g N_VPWR_c_1956_n 0.00333327f $X=15.465 $Y=2.465
+ $X2=0 $Y2=0
cc_1033 N_A_1799_379#_M1025_g N_VPWR_c_1957_n 0.0124152f $X=16.83 $Y=2.155 $X2=0
+ $Y2=0
cc_1034 N_A_1799_379#_M1020_g N_VPWR_c_1962_n 0.00441827f $X=13.115 $Y=2.76
+ $X2=0 $Y2=0
cc_1035 N_A_1799_379#_M1031_g N_VPWR_c_1967_n 0.00525069f $X=15.105 $Y=2.465
+ $X2=0 $Y2=0
cc_1036 N_A_1799_379#_M1011_g N_VPWR_c_1967_n 0.00549284f $X=15.465 $Y=2.465
+ $X2=0 $Y2=0
cc_1037 N_A_1799_379#_M1028_g N_VPWR_c_1967_n 0.00312414f $X=16.47 $Y=2.155
+ $X2=0 $Y2=0
cc_1038 N_A_1799_379#_M1025_g N_VPWR_c_1967_n 0.00312414f $X=16.83 $Y=2.155
+ $X2=0 $Y2=0
cc_1039 N_A_1799_379#_M1020_g N_VPWR_c_1950_n 0.00493098f $X=13.115 $Y=2.76
+ $X2=0 $Y2=0
cc_1040 N_A_1799_379#_M1031_g N_VPWR_c_1950_n 0.00876208f $X=15.105 $Y=2.465
+ $X2=0 $Y2=0
cc_1041 N_A_1799_379#_M1011_g N_VPWR_c_1950_n 0.0111098f $X=15.465 $Y=2.465
+ $X2=0 $Y2=0
cc_1042 N_A_1799_379#_M1028_g N_VPWR_c_1950_n 0.00410284f $X=16.47 $Y=2.155
+ $X2=0 $Y2=0
cc_1043 N_A_1799_379#_M1025_g N_VPWR_c_1950_n 0.00410284f $X=16.83 $Y=2.155
+ $X2=0 $Y2=0
cc_1044 N_A_1799_379#_c_1500_n N_A_1712_379#_c_2146_n 0.0246896f $X=9.935
+ $Y=2.55 $X2=0 $Y2=0
cc_1045 N_A_1799_379#_c_1500_n N_A_1712_379#_c_2147_n 0.0670753f $X=9.935
+ $Y=2.55 $X2=0 $Y2=0
cc_1046 N_A_1799_379#_c_1500_n N_A_1712_379#_c_2149_n 0.00481192f $X=9.935
+ $Y=2.55 $X2=0 $Y2=0
cc_1047 N_A_1799_379#_c_1506_n N_A_2185_397#_c_2173_n 0.0137879f $X=11.585
+ $Y=2.63 $X2=0 $Y2=0
cc_1048 N_A_1799_379#_M1008_g N_A_2185_397#_c_2174_n 6.65587e-19 $X=11.52
+ $Y=2.195 $X2=0 $Y2=0
cc_1049 N_A_1799_379#_c_1505_n N_A_2185_397#_c_2174_n 0.0487199f $X=12.115
+ $Y=2.63 $X2=0 $Y2=0
cc_1050 N_A_1799_379#_c_1506_n N_A_2185_397#_c_2174_n 0.012844f $X=11.585
+ $Y=2.63 $X2=0 $Y2=0
cc_1051 N_A_1799_379#_M1020_g N_A_2185_397#_c_2176_n 0.0024701f $X=13.115
+ $Y=2.76 $X2=0 $Y2=0
cc_1052 N_A_1799_379#_c_1505_n N_A_2185_397#_c_2176_n 0.0137879f $X=12.115
+ $Y=2.63 $X2=0 $Y2=0
cc_1053 N_A_1799_379#_c_1507_n N_A_2185_397#_c_2176_n 0.00442328f $X=12.2
+ $Y=2.545 $X2=0 $Y2=0
cc_1054 N_A_1799_379#_M1020_g N_A_2185_397#_c_2177_n 0.0134314f $X=13.115
+ $Y=2.76 $X2=0 $Y2=0
cc_1055 N_A_1799_379#_c_1508_n N_A_2185_397#_c_2177_n 0.0526231f $X=13.04
+ $Y=2.045 $X2=0 $Y2=0
cc_1056 N_A_1799_379#_c_1485_n N_A_2185_397#_c_2177_n 0.00464767f $X=14.725
+ $Y=1.675 $X2=0 $Y2=0
cc_1057 N_A_1799_379#_c_1489_n N_A_2185_397#_c_2177_n 8.74261e-19 $X=13.205
+ $Y=1.755 $X2=0 $Y2=0
cc_1058 N_A_1799_379#_c_1507_n N_A_2185_397#_c_2178_n 0.00952378f $X=12.2
+ $Y=2.545 $X2=0 $Y2=0
cc_1059 N_A_1799_379#_c_1508_n N_A_2185_397#_c_2178_n 0.0109114f $X=13.04
+ $Y=2.045 $X2=0 $Y2=0
cc_1060 N_A_1799_379#_M1020_g N_A_2185_397#_c_2179_n 0.00965784f $X=13.115
+ $Y=2.76 $X2=0 $Y2=0
cc_1061 N_A_1799_379#_M1008_g N_A_2185_397#_c_2180_n 0.00387094f $X=11.52
+ $Y=2.195 $X2=0 $Y2=0
cc_1062 N_A_1799_379#_c_1504_n N_A_2185_397#_c_2180_n 0.0277216f $X=11.5
+ $Y=2.545 $X2=0 $Y2=0
cc_1063 N_A_1799_379#_c_1487_n N_A_2185_397#_c_2180_n 0.0146211f $X=11.215
+ $Y=1.53 $X2=0 $Y2=0
cc_1064 N_A_1799_379#_c_1491_n N_A_2185_397#_c_2180_n 3.09527e-19 $X=11.52
+ $Y=1.53 $X2=0 $Y2=0
cc_1065 N_A_1799_379#_c_1508_n A_2451_397# 0.00366293f $X=13.04 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_1066 N_A_1799_379#_M1050_g N_Q_N_c_2228_n 0.0028171f $X=15.105 $Y=0.66 $X2=0
+ $Y2=0
cc_1067 N_A_1799_379#_M1031_g N_Q_N_c_2228_n 0.00302423f $X=15.105 $Y=2.465
+ $X2=0 $Y2=0
cc_1068 N_A_1799_379#_M1035_g N_Q_N_c_2228_n 0.0221542f $X=15.465 $Y=0.66 $X2=0
+ $Y2=0
cc_1069 N_A_1799_379#_M1011_g N_Q_N_c_2228_n 0.031729f $X=15.465 $Y=2.465 $X2=0
+ $Y2=0
cc_1070 N_A_1799_379#_c_1473_n N_Q_N_c_2228_n 0.0171532f $X=16.395 $Y=1.42 $X2=0
+ $Y2=0
cc_1071 N_A_1799_379#_M1042_g N_Q_N_c_2228_n 0.00459098f $X=16.47 $Y=0.895 $X2=0
+ $Y2=0
cc_1072 N_A_1799_379#_M1028_g N_Q_N_c_2228_n 0.00531397f $X=16.47 $Y=2.155 $X2=0
+ $Y2=0
cc_1073 N_A_1799_379#_c_1479_n N_Q_N_c_2228_n 0.00251562f $X=15.465 $Y=1.42
+ $X2=0 $Y2=0
cc_1074 N_A_1799_379#_c_1493_n N_Q_N_c_2228_n 4.82746e-19 $X=15.18 $Y=1.51 $X2=0
+ $Y2=0
cc_1075 N_A_1799_379#_M1050_g N_VGND_c_2271_n 0.00990464f $X=15.105 $Y=0.66
+ $X2=0 $Y2=0
cc_1076 N_A_1799_379#_M1048_g N_VGND_c_2272_n 0.0093704f $X=16.83 $Y=0.895 $X2=0
+ $Y2=0
cc_1077 N_A_1799_379#_c_1482_n N_VGND_c_2275_n 0.0197626f $X=9.595 $Y=0.58 $X2=0
+ $Y2=0
cc_1078 N_A_1799_379#_M1030_g N_VGND_c_2276_n 0.00346682f $X=12.78 $Y=0.465
+ $X2=0 $Y2=0
cc_1079 N_A_1799_379#_M1050_g N_VGND_c_2277_n 0.00434176f $X=15.105 $Y=0.66
+ $X2=0 $Y2=0
cc_1080 N_A_1799_379#_M1035_g N_VGND_c_2277_n 0.00544432f $X=15.465 $Y=0.66
+ $X2=0 $Y2=0
cc_1081 N_A_1799_379#_M1042_g N_VGND_c_2277_n 0.00371502f $X=16.47 $Y=0.895
+ $X2=0 $Y2=0
cc_1082 N_A_1799_379#_M1048_g N_VGND_c_2277_n 0.00385058f $X=16.83 $Y=0.895
+ $X2=0 $Y2=0
cc_1083 N_A_1799_379#_M1021_d N_VGND_c_2279_n 0.00230632f $X=9.455 $Y=0.235
+ $X2=0 $Y2=0
cc_1084 N_A_1799_379#_M1030_g N_VGND_c_2279_n 0.0063336f $X=12.78 $Y=0.465 $X2=0
+ $Y2=0
cc_1085 N_A_1799_379#_M1050_g N_VGND_c_2279_n 0.00650883f $X=15.105 $Y=0.66
+ $X2=0 $Y2=0
cc_1086 N_A_1799_379#_M1035_g N_VGND_c_2279_n 0.0110933f $X=15.465 $Y=0.66 $X2=0
+ $Y2=0
cc_1087 N_A_1799_379#_M1042_g N_VGND_c_2279_n 0.00453162f $X=16.47 $Y=0.895
+ $X2=0 $Y2=0
cc_1088 N_A_1799_379#_M1048_g N_VGND_c_2279_n 0.00453162f $X=16.83 $Y=0.895
+ $X2=0 $Y2=0
cc_1089 N_A_1799_379#_c_1482_n N_VGND_c_2279_n 0.0125808f $X=9.595 $Y=0.58 $X2=0
+ $Y2=0
cc_1090 N_CLK_M1034_g N_VPWR_c_1956_n 0.00783653f $X=14.44 $Y=2.155 $X2=0 $Y2=0
cc_1091 N_CLK_M1049_g N_VPWR_c_1962_n 0.00312414f $X=14.08 $Y=2.155 $X2=0 $Y2=0
cc_1092 N_CLK_M1034_g N_VPWR_c_1962_n 0.00312414f $X=14.44 $Y=2.155 $X2=0 $Y2=0
cc_1093 N_CLK_M1049_g N_VPWR_c_1950_n 0.00410284f $X=14.08 $Y=2.155 $X2=0 $Y2=0
cc_1094 N_CLK_M1034_g N_VPWR_c_1950_n 0.00410284f $X=14.44 $Y=2.155 $X2=0 $Y2=0
cc_1095 N_CLK_M1049_g N_A_2185_397#_c_2177_n 4.90203e-19 $X=14.08 $Y=2.155 $X2=0
+ $Y2=0
cc_1096 N_CLK_M1049_g N_A_2185_397#_c_2179_n 0.0029149f $X=14.08 $Y=2.155 $X2=0
+ $Y2=0
cc_1097 N_CLK_M1026_g N_VGND_c_2271_n 0.00200234f $X=14.05 $Y=0.45 $X2=0 $Y2=0
cc_1098 N_CLK_M1027_g N_VGND_c_2271_n 0.0106757f $X=14.44 $Y=0.45 $X2=0 $Y2=0
cc_1099 N_CLK_M1026_g N_VGND_c_2276_n 0.00421223f $X=14.05 $Y=0.45 $X2=0 $Y2=0
cc_1100 N_CLK_M1027_g N_VGND_c_2276_n 0.00361037f $X=14.44 $Y=0.45 $X2=0 $Y2=0
cc_1101 N_CLK_M1026_g N_VGND_c_2279_n 0.00730136f $X=14.05 $Y=0.45 $X2=0 $Y2=0
cc_1102 N_CLK_M1027_g N_VGND_c_2279_n 0.00425021f $X=14.44 $Y=0.45 $X2=0 $Y2=0
cc_1103 N_A_3222_137#_M1037_g N_VPWR_c_1957_n 0.0300646f $X=17.375 $Y=2.465
+ $X2=0 $Y2=0
cc_1104 N_A_3222_137#_M1046_g N_VPWR_c_1957_n 0.00468428f $X=17.735 $Y=2.465
+ $X2=0 $Y2=0
cc_1105 N_A_3222_137#_c_1782_n N_VPWR_c_1957_n 0.0203141f $X=16.255 $Y=1.98
+ $X2=0 $Y2=0
cc_1106 N_A_3222_137#_c_1777_n N_VPWR_c_1957_n 0.0275493f $X=17.44 $Y=1.47 $X2=0
+ $Y2=0
cc_1107 N_A_3222_137#_c_1779_n N_VPWR_c_1957_n 5.79521e-19 $X=17.735 $Y=1.47
+ $X2=0 $Y2=0
cc_1108 N_A_3222_137#_M1037_g N_VPWR_c_1968_n 0.00486043f $X=17.375 $Y=2.465
+ $X2=0 $Y2=0
cc_1109 N_A_3222_137#_M1046_g N_VPWR_c_1968_n 0.00549284f $X=17.735 $Y=2.465
+ $X2=0 $Y2=0
cc_1110 N_A_3222_137#_M1037_g N_VPWR_c_1950_n 0.00814425f $X=17.375 $Y=2.465
+ $X2=0 $Y2=0
cc_1111 N_A_3222_137#_M1046_g N_VPWR_c_1950_n 0.0107699f $X=17.735 $Y=2.465
+ $X2=0 $Y2=0
cc_1112 N_A_3222_137#_c_1782_n N_VPWR_c_1950_n 0.0128958f $X=16.255 $Y=1.98
+ $X2=0 $Y2=0
cc_1113 N_A_3222_137#_c_1776_n N_Q_N_c_2228_n 0.0412742f $X=16.255 $Y=0.895
+ $X2=0 $Y2=0
cc_1114 N_A_3222_137#_c_1782_n N_Q_N_c_2228_n 0.0554733f $X=16.255 $Y=1.98 $X2=0
+ $Y2=0
cc_1115 N_A_3222_137#_c_1778_n N_Q_N_c_2228_n 0.0212537f $X=16.255 $Y=1.47 $X2=0
+ $Y2=0
cc_1116 N_A_3222_137#_M1015_g N_Q_c_2251_n 0.00323857f $X=17.375 $Y=0.685 $X2=0
+ $Y2=0
cc_1117 N_A_3222_137#_M1037_g N_Q_c_2251_n 0.00430008f $X=17.375 $Y=2.465 $X2=0
+ $Y2=0
cc_1118 N_A_3222_137#_M1018_g N_Q_c_2251_n 0.0238324f $X=17.735 $Y=0.685 $X2=0
+ $Y2=0
cc_1119 N_A_3222_137#_M1046_g N_Q_c_2251_n 0.0300568f $X=17.735 $Y=2.465 $X2=0
+ $Y2=0
cc_1120 N_A_3222_137#_c_1777_n N_Q_c_2251_n 0.0250026f $X=17.44 $Y=1.47 $X2=0
+ $Y2=0
cc_1121 N_A_3222_137#_c_1779_n N_Q_c_2251_n 0.0121537f $X=17.735 $Y=1.47 $X2=0
+ $Y2=0
cc_1122 N_A_3222_137#_M1015_g N_VGND_c_2272_n 0.0221425f $X=17.375 $Y=0.685
+ $X2=0 $Y2=0
cc_1123 N_A_3222_137#_M1018_g N_VGND_c_2272_n 0.00336955f $X=17.735 $Y=0.685
+ $X2=0 $Y2=0
cc_1124 N_A_3222_137#_c_1776_n N_VGND_c_2272_n 0.0137622f $X=16.255 $Y=0.895
+ $X2=0 $Y2=0
cc_1125 N_A_3222_137#_c_1777_n N_VGND_c_2272_n 0.0275493f $X=17.44 $Y=1.47 $X2=0
+ $Y2=0
cc_1126 N_A_3222_137#_c_1779_n N_VGND_c_2272_n 5.79521e-19 $X=17.735 $Y=1.47
+ $X2=0 $Y2=0
cc_1127 N_A_3222_137#_c_1776_n N_VGND_c_2277_n 0.00619475f $X=16.255 $Y=0.895
+ $X2=0 $Y2=0
cc_1128 N_A_3222_137#_M1015_g N_VGND_c_2278_n 0.00461019f $X=17.375 $Y=0.685
+ $X2=0 $Y2=0
cc_1129 N_A_3222_137#_M1018_g N_VGND_c_2278_n 0.00520813f $X=17.735 $Y=0.685
+ $X2=0 $Y2=0
cc_1130 N_A_3222_137#_M1015_g N_VGND_c_2279_n 0.00803623f $X=17.375 $Y=0.685
+ $X2=0 $Y2=0
cc_1131 N_A_3222_137#_M1018_g N_VGND_c_2279_n 0.0104074f $X=17.735 $Y=0.685
+ $X2=0 $Y2=0
cc_1132 N_A_3222_137#_c_1776_n N_VGND_c_2279_n 0.00970591f $X=16.255 $Y=0.895
+ $X2=0 $Y2=0
cc_1133 N_A_27_457#_c_1834_n N_A_111_457#_c_1876_n 0.0172014f $X=0.265 $Y=2.495
+ $X2=0 $Y2=0
cc_1134 N_A_27_457#_c_1835_n N_A_111_457#_c_1876_n 0.0244976f $X=1.04 $Y=2.98
+ $X2=0 $Y2=0
cc_1135 N_A_27_457#_c_1837_n N_A_111_457#_c_1876_n 0.00874792f $X=1.125 $Y=2.895
+ $X2=0 $Y2=0
cc_1136 N_A_27_457#_c_1838_n N_A_111_457#_c_1877_n 0.065789f $X=1.935 $Y=2.395
+ $X2=0 $Y2=0
cc_1137 N_A_27_457#_c_1853_n N_A_111_457#_c_1877_n 0.0105422f $X=1.21 $Y=2.395
+ $X2=0 $Y2=0
cc_1138 N_A_27_457#_c_1853_n A_197_457# 0.00103727f $X=1.21 $Y=2.395 $X2=-0.19
+ $Y2=1.655
cc_1139 N_A_27_457#_c_1838_n N_VPWR_M1022_d 0.00497047f $X=1.935 $Y=2.395
+ $X2=-0.19 $Y2=1.655
cc_1140 N_A_27_457#_c_1835_n N_VPWR_c_1951_n 0.0127464f $X=1.04 $Y=2.98 $X2=0
+ $Y2=0
cc_1141 N_A_27_457#_c_1837_n N_VPWR_c_1951_n 0.0150227f $X=1.125 $Y=2.895 $X2=0
+ $Y2=0
cc_1142 N_A_27_457#_c_1838_n N_VPWR_c_1951_n 0.0204359f $X=1.935 $Y=2.395 $X2=0
+ $Y2=0
cc_1143 N_A_27_457#_c_1839_n N_VPWR_c_1951_n 0.0096883f $X=2.02 $Y=2.68 $X2=0
+ $Y2=0
cc_1144 N_A_27_457#_c_1839_n N_VPWR_c_1958_n 0.00854876f $X=2.02 $Y=2.68 $X2=0
+ $Y2=0
cc_1145 N_A_27_457#_c_1835_n N_VPWR_c_1964_n 0.0528019f $X=1.04 $Y=2.98 $X2=0
+ $Y2=0
cc_1146 N_A_27_457#_c_1836_n N_VPWR_c_1964_n 0.0168561f $X=0.35 $Y=2.98 $X2=0
+ $Y2=0
cc_1147 N_A_27_457#_c_1835_n N_VPWR_c_1950_n 0.0290283f $X=1.04 $Y=2.98 $X2=0
+ $Y2=0
cc_1148 N_A_27_457#_c_1836_n N_VPWR_c_1950_n 0.00967329f $X=0.35 $Y=2.98 $X2=0
+ $Y2=0
cc_1149 N_A_27_457#_c_1838_n N_VPWR_c_1950_n 0.0124543f $X=1.935 $Y=2.395 $X2=0
+ $Y2=0
cc_1150 N_A_27_457#_c_1839_n N_VPWR_c_1950_n 0.00872122f $X=2.02 $Y=2.68 $X2=0
+ $Y2=0
cc_1151 N_A_27_457#_c_1838_n N_A_484_411#_c_2103_n 0.0131471f $X=1.935 $Y=2.395
+ $X2=0 $Y2=0
cc_1152 N_A_27_457#_c_1839_n N_A_484_411#_c_2103_n 0.0294905f $X=2.02 $Y=2.68
+ $X2=0 $Y2=0
cc_1153 N_A_27_457#_c_1839_n N_A_484_411#_c_2105_n 0.00116004f $X=2.02 $Y=2.68
+ $X2=0 $Y2=0
cc_1154 N_A_111_457#_c_1877_n N_A_484_411#_M1024_s 0.00110883f $X=2.495 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_1155 N_A_111_457#_c_1880_n N_A_484_411#_M1024_s 0.00863065f $X=2.9 $Y=2.545
+ $X2=-0.19 $Y2=-0.245
cc_1156 N_A_111_457#_c_1884_n N_A_484_411#_M1024_s 0.0103041f $X=2.74 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_1157 N_A_111_457#_c_1877_n N_A_484_411#_c_2103_n 0.00827348f $X=2.495
+ $Y=2.045 $X2=0 $Y2=0
cc_1158 N_A_111_457#_c_1880_n N_A_484_411#_c_2103_n 0.0169039f $X=2.9 $Y=2.545
+ $X2=0 $Y2=0
cc_1159 N_A_111_457#_c_1882_n N_A_484_411#_c_2103_n 0.0140495f $X=2.985 $Y=2.63
+ $X2=0 $Y2=0
cc_1160 N_A_111_457#_c_1884_n N_A_484_411#_c_2103_n 0.0116368f $X=2.74 $Y=2.045
+ $X2=0 $Y2=0
cc_1161 N_A_111_457#_c_1881_n N_A_484_411#_c_2104_n 0.0599206f $X=3.515 $Y=2.63
+ $X2=0 $Y2=0
cc_1162 N_A_111_457#_c_1882_n N_A_484_411#_c_2104_n 0.0126496f $X=2.985 $Y=2.63
+ $X2=0 $Y2=0
cc_1163 N_A_111_457#_c_1881_n N_A_484_411#_c_2106_n 0.00419222f $X=3.515 $Y=2.63
+ $X2=0 $Y2=0
cc_1164 N_A_111_457#_c_1875_n N_VGND_c_2274_n 0.00652123f $X=2.66 $Y=0.79 $X2=0
+ $Y2=0
cc_1165 N_A_111_457#_c_1875_n N_VGND_c_2279_n 0.0103348f $X=2.66 $Y=0.79 $X2=0
+ $Y2=0
cc_1166 N_VPWR_c_1958_n N_A_484_411#_c_2104_n 0.0856245f $X=4.66 $Y=3.33 $X2=0
+ $Y2=0
cc_1167 N_VPWR_c_1950_n N_A_484_411#_c_2104_n 0.0485802f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1168 N_VPWR_c_1951_n N_A_484_411#_c_2105_n 0.00485018f $X=1.59 $Y=2.745 $X2=0
+ $Y2=0
cc_1169 N_VPWR_c_1958_n N_A_484_411#_c_2105_n 0.0168561f $X=4.66 $Y=3.33 $X2=0
+ $Y2=0
cc_1170 N_VPWR_c_1950_n N_A_484_411#_c_2105_n 0.00967329f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1171 N_VPWR_c_1952_n N_A_484_411#_c_2106_n 0.0226815f $X=4.825 $Y=2.825 $X2=0
+ $Y2=0
cc_1172 N_VPWR_c_1958_n N_A_484_411#_c_2106_n 0.0212726f $X=4.66 $Y=3.33 $X2=0
+ $Y2=0
cc_1173 N_VPWR_c_1950_n N_A_484_411#_c_2106_n 0.0112117f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1174 N_VPWR_c_1950_n N_A_1712_379#_M1013_s 0.00426945f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1175 N_VPWR_c_1966_n N_A_1712_379#_c_2147_n 0.0857091f $X=10.635 $Y=3.33
+ $X2=0 $Y2=0
cc_1176 N_VPWR_c_1950_n N_A_1712_379#_c_2147_n 0.0528788f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1177 N_VPWR_c_1966_n N_A_1712_379#_c_2148_n 0.0168561f $X=10.635 $Y=3.33
+ $X2=0 $Y2=0
cc_1178 N_VPWR_c_1950_n N_A_1712_379#_c_2148_n 0.00967329f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1179 N_VPWR_c_1954_n N_A_1712_379#_c_2149_n 0.0147694f $X=10.8 $Y=2.885 $X2=0
+ $Y2=0
cc_1180 N_VPWR_c_1966_n N_A_1712_379#_c_2149_n 0.0106732f $X=10.635 $Y=3.33
+ $X2=0 $Y2=0
cc_1181 N_VPWR_c_1950_n N_A_1712_379#_c_2149_n 0.00640972f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1182 N_VPWR_c_1954_n N_A_2185_397#_c_2173_n 0.0175221f $X=10.8 $Y=2.885 $X2=0
+ $Y2=0
cc_1183 N_VPWR_c_1955_n N_A_2185_397#_c_2174_n 0.0136857f $X=12.9 $Y=2.825 $X2=0
+ $Y2=0
cc_1184 N_VPWR_c_1960_n N_A_2185_397#_c_2174_n 0.0859881f $X=12.815 $Y=3.33
+ $X2=0 $Y2=0
cc_1185 N_VPWR_c_1950_n N_A_2185_397#_c_2174_n 0.0525385f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1186 N_VPWR_c_1954_n N_A_2185_397#_c_2175_n 0.0139102f $X=10.8 $Y=2.885 $X2=0
+ $Y2=0
cc_1187 N_VPWR_c_1960_n N_A_2185_397#_c_2175_n 0.0114622f $X=12.815 $Y=3.33
+ $X2=0 $Y2=0
cc_1188 N_VPWR_c_1950_n N_A_2185_397#_c_2175_n 0.00657784f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1955_n N_A_2185_397#_c_2176_n 0.0166412f $X=12.9 $Y=2.825 $X2=0
+ $Y2=0
cc_1190 N_VPWR_M1001_d N_A_2185_397#_c_2177_n 0.00724808f $X=12.615 $Y=1.985
+ $X2=0 $Y2=0
cc_1191 N_VPWR_c_1955_n N_A_2185_397#_c_2177_n 0.0127505f $X=12.9 $Y=2.825 $X2=0
+ $Y2=0
cc_1192 N_VPWR_c_1950_n N_A_2185_397#_c_2177_n 0.0120115f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1193 N_VPWR_c_1955_n N_A_2185_397#_c_2179_n 0.0125142f $X=12.9 $Y=2.825 $X2=0
+ $Y2=0
cc_1194 N_VPWR_c_1962_n N_A_2185_397#_c_2179_n 0.0151738f $X=14.715 $Y=3.33
+ $X2=0 $Y2=0
cc_1195 N_VPWR_c_1950_n N_A_2185_397#_c_2179_n 0.0120712f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1950_n A_3036_367# 0.00899413f $X=18 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1197 N_VPWR_c_1950_n N_Q_N_M1011_d 0.0023218f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1198 N_VPWR_c_1956_n N_Q_N_c_2228_n 0.0254541f $X=14.88 $Y=2.455 $X2=0 $Y2=0
cc_1199 N_VPWR_c_1967_n N_Q_N_c_2228_n 0.019758f $X=16.995 $Y=3.33 $X2=0 $Y2=0
cc_1200 N_VPWR_c_1950_n N_Q_N_c_2228_n 0.012508f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1201 N_VPWR_c_1950_n A_3490_367# 0.00899413f $X=18 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1202 N_VPWR_c_1950_n N_Q_M1046_d 0.0023218f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1203 N_VPWR_c_1957_n N_Q_c_2251_n 0.0418217f $X=17.16 $Y=1.98 $X2=0 $Y2=0
cc_1204 N_VPWR_c_1968_n N_Q_c_2251_n 0.019758f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1205 N_VPWR_c_1950_n N_Q_c_2251_n 0.012508f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1206 N_Q_N_c_2228_n N_VGND_c_2277_n 0.019758f $X=15.68 $Y=0.43 $X2=0 $Y2=0
cc_1207 N_Q_N_M1035_d N_VGND_c_2279_n 0.00230415f $X=15.54 $Y=0.24 $X2=0 $Y2=0
cc_1208 N_Q_N_c_2228_n N_VGND_c_2279_n 0.012508f $X=15.68 $Y=0.43 $X2=0 $Y2=0
cc_1209 N_Q_c_2251_n N_VGND_c_2272_n 0.0287733f $X=17.95 $Y=0.43 $X2=0 $Y2=0
cc_1210 N_Q_c_2251_n N_VGND_c_2278_n 0.019758f $X=17.95 $Y=0.43 $X2=0 $Y2=0
cc_1211 N_Q_c_2251_n N_VGND_c_2279_n 0.0125705f $X=17.95 $Y=0.43 $X2=0 $Y2=0
cc_1212 N_VGND_c_2279_n A_2825_48# 0.00312641f $X=18 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1213 N_VGND_c_2279_n A_3036_48# 0.00437243f $X=18 $Y=0 $X2=-0.19 $Y2=-0.245
