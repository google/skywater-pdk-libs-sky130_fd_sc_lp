* File: sky130_fd_sc_lp__invlp_4.spice
* Created: Fri Aug 28 10:40:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__invlp_4.pex.spice"
.subckt sky130_fd_sc_lp__invlp_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_114_53#_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.5 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_114_53#_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1764 AS=0.1176 PD=1.26 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1009_d N_A_M1011_g N_A_114_53#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1764 AS=0.1176 PD=1.26 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1003 N_A_114_53#_M1011_s N_A_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1006 N_A_114_53#_M1006_d N_A_M1006_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1007 N_A_114_53#_M1006_d N_A_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.5
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1014 N_A_114_53#_M1014_d N_A_M1014_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=9.996 NRS=0 M=1 R=5.6 SA=75003
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_A_M1015_g N_A_114_53#_M1014_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.147 PD=2.25 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75003.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_118_367#_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_118_367#_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1004_d N_A_M1005_g N_A_118_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1001 N_A_118_367#_M1005_s N_A_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2205 PD=1.54 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4 SA=75001.5
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1008 N_A_118_367#_M1008_d N_A_M1008_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75002
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1010 N_A_118_367#_M1008_d N_A_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4 SA=75002.5
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1013 N_A_118_367#_M1013_d N_A_M1013_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2205 PD=1.54 PS=1.61 NRD=0 NRS=0 M=1 R=8.4 SA=75003 SB=75000.7
+ A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g N_A_118_367#_M1013_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4473 AS=0.1764 PD=3.23 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75003.4
+ SB=75000.3 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__invlp_4.pxi.spice"
*
.ends
*
*
