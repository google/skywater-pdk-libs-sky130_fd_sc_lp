* NGSPICE file created from sky130_fd_sc_lp__o211ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 Y B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.1168e+12p pd=1.848e+07u as=2.9106e+12p ps=2.226e+07u
M1001 a_836_47# B1 a_57_47# VNB nshort w=840000u l=150000u
+  ad=1.4985e+12p pd=1.072e+07u as=1.6632e+12p ps=1.572e+07u
M1002 a_57_47# B1 a_836_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_836_47# C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.48e+06u
M1004 a_140_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.4112e+12p pd=1.232e+07u as=0p ps=0u
M1005 VPWR A1 a_140_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_57_47# VNB nshort w=840000u l=150000u
+  ad=9.492e+11p pd=8.98e+06u as=0p ps=0u
M1007 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_57_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y C1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_57_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_140_367# A2 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_140_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_836_47# B1 a_57_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_57_47# B1 a_836_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C1 a_836_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_57_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_140_367# A2 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A1 a_57_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A2 a_140_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_836_47# C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_57_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y C1 a_836_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A2 a_140_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_57_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_57_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y C1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_140_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

