* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand4bb_lp A_N B_N C D VGND VNB VPB VPWR Y
X0 a_114_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_47# A_N a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_456_47# C a_534_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_534_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND B_N a_708_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_384_47# a_332_352# a_456_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Y a_332_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VPWR B_N a_332_352# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_708_47# B_N a_332_352# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 Y a_27_47# a_384_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
