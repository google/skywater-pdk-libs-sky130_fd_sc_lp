* File: sky130_fd_sc_lp__o221a_lp.pxi.spice
* Created: Wed Sep  2 10:18:37 2020
* 
x_PM_SKY130_FD_SC_LP__O221A_LP%A_84_21# N_A_84_21#_M1012_d N_A_84_21#_M1001_d
+ N_A_84_21#_M1010_d N_A_84_21#_c_93_n N_A_84_21#_M1002_g N_A_84_21#_c_94_n
+ N_A_84_21#_M1000_g N_A_84_21#_c_95_n N_A_84_21#_c_96_n N_A_84_21#_M1009_g
+ N_A_84_21#_c_97_n N_A_84_21#_c_105_n N_A_84_21#_c_106_n N_A_84_21#_c_98_n
+ N_A_84_21#_c_99_n N_A_84_21#_c_108_n N_A_84_21#_c_117_p N_A_84_21#_c_109_n
+ N_A_84_21#_c_110_n N_A_84_21#_c_111_n N_A_84_21#_c_100_n N_A_84_21#_c_101_n
+ N_A_84_21#_c_102_n PM_SKY130_FD_SC_LP__O221A_LP%A_84_21#
x_PM_SKY130_FD_SC_LP__O221A_LP%A1 N_A1_M1005_g N_A1_M1003_g N_A1_c_202_n
+ N_A1_c_203_n N_A1_c_204_n N_A1_c_205_n N_A1_c_206_n A1 A1 N_A1_c_208_n
+ PM_SKY130_FD_SC_LP__O221A_LP%A1
x_PM_SKY130_FD_SC_LP__O221A_LP%A2 N_A2_M1001_g N_A2_M1006_g N_A2_c_254_n
+ N_A2_c_255_n A2 A2 N_A2_c_257_n PM_SKY130_FD_SC_LP__O221A_LP%A2
x_PM_SKY130_FD_SC_LP__O221A_LP%B2 N_B2_M1008_g N_B2_c_297_n N_B2_c_298_n
+ N_B2_c_299_n N_B2_M1007_g B2 B2 N_B2_c_301_n N_B2_c_302_n
+ PM_SKY130_FD_SC_LP__O221A_LP%B2
x_PM_SKY130_FD_SC_LP__O221A_LP%B1 N_B1_c_358_n N_B1_M1004_g N_B1_c_353_n
+ N_B1_c_354_n N_B1_M1011_g N_B1_c_360_n B1 N_B1_c_356_n N_B1_c_357_n
+ PM_SKY130_FD_SC_LP__O221A_LP%B1
x_PM_SKY130_FD_SC_LP__O221A_LP%C1 N_C1_c_409_n N_C1_M1010_g N_C1_c_410_n
+ N_C1_c_411_n N_C1_M1012_g N_C1_c_412_n C1 N_C1_c_407_n N_C1_c_408_n
+ PM_SKY130_FD_SC_LP__O221A_LP%C1
x_PM_SKY130_FD_SC_LP__O221A_LP%X N_X_M1002_s N_X_M1000_s N_X_c_452_n N_X_c_449_n
+ X X X PM_SKY130_FD_SC_LP__O221A_LP%X
x_PM_SKY130_FD_SC_LP__O221A_LP%VPWR N_VPWR_M1000_d N_VPWR_M1004_d N_VPWR_c_476_n
+ N_VPWR_c_477_n VPWR N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_475_n
+ N_VPWR_c_481_n N_VPWR_c_482_n PM_SKY130_FD_SC_LP__O221A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O221A_LP%VGND N_VGND_M1009_d N_VGND_M1006_d N_VGND_c_524_n
+ N_VGND_c_525_n N_VGND_c_526_n VGND N_VGND_c_527_n N_VGND_c_528_n
+ N_VGND_c_529_n N_VGND_c_530_n PM_SKY130_FD_SC_LP__O221A_LP%VGND
x_PM_SKY130_FD_SC_LP__O221A_LP%A_272_47# N_A_272_47#_M1003_d N_A_272_47#_M1007_d
+ N_A_272_47#_c_575_n N_A_272_47#_c_576_n N_A_272_47#_c_577_n
+ PM_SKY130_FD_SC_LP__O221A_LP%A_272_47#
x_PM_SKY130_FD_SC_LP__O221A_LP%A_490_141# N_A_490_141#_M1007_s
+ N_A_490_141#_M1011_d N_A_490_141#_c_612_n N_A_490_141#_c_632_n
+ N_A_490_141#_c_613_n PM_SKY130_FD_SC_LP__O221A_LP%A_490_141#
cc_1 VNB N_A_84_21#_c_93_n 0.0172354f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_2 VNB N_A_84_21#_c_94_n 0.0184061f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.715
cc_3 VNB N_A_84_21#_c_95_n 0.0204529f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_4 VNB N_A_84_21#_c_96_n 0.01359f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_5 VNB N_A_84_21#_c_97_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_6 VNB N_A_84_21#_c_98_n 0.00621681f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.39
cc_7 VNB N_A_84_21#_c_99_n 0.0166207f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.39
cc_8 VNB N_A_84_21#_c_100_n 0.030893f $X=-0.19 $Y=-0.245 $X2=3.82 $Y2=1.97
cc_9 VNB N_A_84_21#_c_101_n 0.0167284f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=0.85
cc_10 VNB N_A_84_21#_c_102_n 0.0205153f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.225
cc_11 VNB N_A1_c_202_n 0.0170898f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_12 VNB N_A1_c_203_n 0.0238816f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_13 VNB N_A1_c_204_n 0.00211967f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_14 VNB N_A1_c_205_n 0.0143983f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.225
cc_15 VNB N_A1_c_206_n 0.00916751f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.405
cc_16 VNB A1 0.00373964f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.715
cc_17 VNB N_A1_c_208_n 0.019875f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_18 VNB N_A2_M1006_g 0.0403591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_254_n 0.0220502f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_20 VNB N_A2_c_255_n 0.0019315f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_21 VNB A2 0.00562791f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_22 VNB N_A2_c_257_n 0.0163324f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.595
cc_23 VNB N_B2_c_297_n 0.030551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B2_c_298_n 0.0102342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B2_c_299_n 0.0138274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB B2 0.00970037f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_27 VNB N_B2_c_301_n 0.0223099f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.895
cc_28 VNB N_B2_c_302_n 0.0468882f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.595
cc_29 VNB N_B1_c_353_n 0.00748376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B1_c_354_n 0.00706981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B1_M1011_g 0.0290305f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_32 VNB N_B1_c_356_n 0.0259054f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.715
cc_33 VNB N_B1_c_357_n 0.00412367f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.895
cc_34 VNB N_C1_M1012_g 0.0319965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C1_c_407_n 0.0280924f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.405
cc_36 VNB N_C1_c_408_n 0.00303343f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.715
cc_37 VNB N_X_c_449_n 0.0289131f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_38 VNB X 0.0243904f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.225
cc_39 VNB X 0.0134386f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_40 VNB N_VPWR_c_475_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.39
cc_41 VNB N_VGND_c_524_n 0.00759122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_525_n 0.026731f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_43 VNB N_VGND_c_526_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_44 VNB N_VGND_c_527_n 0.0179305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_528_n 0.0621511f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_46 VNB N_VGND_c_529_n 0.255377f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.895
cc_47 VNB N_VGND_c_530_n 0.0158798f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.39
cc_48 VNB N_A_272_47#_c_575_n 0.0133811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_272_47#_c_576_n 0.00877209f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_50 VNB N_A_272_47#_c_577_n 0.00379004f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.225
cc_51 VNB N_A_490_141#_c_612_n 0.0077453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_490_141#_c_613_n 0.00610182f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.225
cc_53 VPB N_A_84_21#_c_94_n 0.00434968f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.715
cc_54 VPB N_A_84_21#_M1000_g 0.0331548f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.595
cc_55 VPB N_A_84_21#_c_105_n 0.0167238f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.895
cc_56 VPB N_A_84_21#_c_106_n 0.00266219f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.7
cc_57 VPB N_A_84_21#_c_98_n 2.74074e-19 $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.39
cc_58 VPB N_A_84_21#_c_108_n 0.0143311f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=2.055
cc_59 VPB N_A_84_21#_c_109_n 0.00447965f $X=-0.19 $Y=1.655 $X2=3.405 $Y2=2.055
cc_60 VPB N_A_84_21#_c_110_n 0.00667764f $X=-0.19 $Y=1.655 $X2=1.98 $Y2=2.055
cc_61 VPB N_A_84_21#_c_111_n 0.0729261f $X=-0.19 $Y=1.655 $X2=3.82 $Y2=2.055
cc_62 VPB N_A_84_21#_c_100_n 0.0153385f $X=-0.19 $Y=1.655 $X2=3.82 $Y2=1.97
cc_63 VPB N_A1_M1005_g 0.0344816f $X=-0.19 $Y=1.655 $X2=3.43 $Y2=2.095
cc_64 VPB N_A1_c_204_n 0.0117934f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.88
cc_65 VPB A1 7.56276e-19 $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.715
cc_66 VPB N_A2_M1001_g 0.033813f $X=-0.19 $Y=1.655 $X2=3.43 $Y2=2.095
cc_67 VPB N_A2_c_255_n 0.010854f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_68 VPB A2 0.00140835f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.88
cc_69 VPB N_B2_M1008_g 0.0381319f $X=-0.19 $Y=1.655 $X2=3.43 $Y2=2.095
cc_70 VPB B2 0.00486424f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.88
cc_71 VPB N_B2_c_301_n 0.00642472f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.895
cc_72 VPB N_B1_c_358_n 0.0244181f $X=-0.19 $Y=1.655 $X2=3.82 $Y2=0.61
cc_73 VPB N_B1_c_353_n 0.00476024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_B1_c_360_n 0.018882f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_75 VPB N_B1_c_356_n 0.00600421f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.715
cc_76 VPB N_B1_c_357_n 0.00418191f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.895
cc_77 VPB N_C1_c_409_n 0.0229078f $X=-0.19 $Y=1.655 $X2=3.82 $Y2=0.61
cc_78 VPB N_C1_c_410_n 0.0279317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_C1_c_411_n 0.0116596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_C1_c_412_n 0.0162813f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_81 VPB N_C1_c_407_n 0.00445132f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.405
cc_82 VPB N_C1_c_408_n 0.0040159f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.715
cc_83 VPB N_X_c_452_n 0.0477195f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_84 VPB N_X_c_449_n 0.0198276f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.88
cc_85 VPB N_VPWR_c_476_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_86 VPB N_VPWR_c_477_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.405
cc_87 VPB N_VPWR_c_478_n 0.0548934f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.595
cc_88 VPB N_VPWR_c_479_n 0.0289392f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.39
cc_89 VPB N_VPWR_c_475_n 0.0491228f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.39
cc_90 VPB N_VPWR_c_481_n 0.0245825f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=2.055
cc_91 VPB N_VPWR_c_482_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.98 $Y2=2.24
cc_92 N_A_84_21#_M1000_g N_A1_M1005_g 0.0275437f $X=0.59 $Y=2.595 $X2=0 $Y2=0
cc_93 N_A_84_21#_c_105_n N_A1_M1005_g 0.00375943f $X=0.6 $Y=1.895 $X2=0 $Y2=0
cc_94 N_A_84_21#_c_106_n N_A1_M1005_g 0.0038764f $X=0.645 $Y=1.7 $X2=0 $Y2=0
cc_95 N_A_84_21#_c_108_n N_A1_M1005_g 0.022761f $X=1.815 $Y=2.055 $X2=0 $Y2=0
cc_96 N_A_84_21#_c_117_p N_A1_M1005_g 0.0039963f $X=1.98 $Y=2.24 $X2=0 $Y2=0
cc_97 N_A_84_21#_c_102_n N_A1_c_202_n 0.00359595f $X=0.6 $Y=1.225 $X2=0 $Y2=0
cc_98 N_A_84_21#_c_94_n N_A1_c_203_n 0.0099089f $X=0.6 $Y=1.715 $X2=0 $Y2=0
cc_99 N_A_84_21#_c_105_n N_A1_c_204_n 0.0099089f $X=0.6 $Y=1.895 $X2=0 $Y2=0
cc_100 N_A_84_21#_c_106_n N_A1_c_204_n 5.54119e-19 $X=0.645 $Y=1.7 $X2=0 $Y2=0
cc_101 N_A_84_21#_c_108_n N_A1_c_204_n 5.43485e-19 $X=1.815 $Y=2.055 $X2=0 $Y2=0
cc_102 N_A_84_21#_c_96_n N_A1_c_205_n 0.010809f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_103 N_A_84_21#_c_95_n N_A1_c_206_n 0.0087141f $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_104 N_A_84_21#_c_106_n A1 0.00694705f $X=0.645 $Y=1.7 $X2=0 $Y2=0
cc_105 N_A_84_21#_c_98_n A1 0.0363845f $X=0.615 $Y=1.39 $X2=0 $Y2=0
cc_106 N_A_84_21#_c_99_n A1 6.38995e-19 $X=0.615 $Y=1.39 $X2=0 $Y2=0
cc_107 N_A_84_21#_c_108_n A1 0.0241279f $X=1.815 $Y=2.055 $X2=0 $Y2=0
cc_108 N_A_84_21#_c_98_n N_A1_c_208_n 0.00291435f $X=0.615 $Y=1.39 $X2=0 $Y2=0
cc_109 N_A_84_21#_c_99_n N_A1_c_208_n 0.0099089f $X=0.615 $Y=1.39 $X2=0 $Y2=0
cc_110 N_A_84_21#_c_102_n N_A1_c_208_n 4.39265e-19 $X=0.6 $Y=1.225 $X2=0 $Y2=0
cc_111 N_A_84_21#_c_108_n N_A2_M1001_g 0.0183235f $X=1.815 $Y=2.055 $X2=0 $Y2=0
cc_112 N_A_84_21#_c_117_p N_A2_M1001_g 0.0214638f $X=1.98 $Y=2.24 $X2=0 $Y2=0
cc_113 N_A_84_21#_c_110_n N_A2_M1001_g 0.0023941f $X=1.98 $Y=2.055 $X2=0 $Y2=0
cc_114 N_A_84_21#_c_110_n N_A2_c_255_n 0.00264669f $X=1.98 $Y=2.055 $X2=0 $Y2=0
cc_115 N_A_84_21#_c_108_n A2 0.0182583f $X=1.815 $Y=2.055 $X2=0 $Y2=0
cc_116 N_A_84_21#_c_110_n A2 0.00449095f $X=1.98 $Y=2.055 $X2=0 $Y2=0
cc_117 N_A_84_21#_c_109_n N_B2_M1008_g 0.0219258f $X=3.405 $Y=2.055 $X2=0 $Y2=0
cc_118 N_A_84_21#_c_109_n B2 0.0434595f $X=3.405 $Y=2.055 $X2=0 $Y2=0
cc_119 N_A_84_21#_c_110_n B2 0.00868118f $X=1.98 $Y=2.055 $X2=0 $Y2=0
cc_120 N_A_84_21#_c_109_n N_B2_c_301_n 4.79059e-19 $X=3.405 $Y=2.055 $X2=0 $Y2=0
cc_121 N_A_84_21#_c_109_n N_B1_c_358_n 0.0242371f $X=3.405 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_84_21#_c_111_n N_B1_c_358_n 9.80034e-19 $X=3.82 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_84_21#_c_109_n N_B1_c_353_n 0.00401082f $X=3.405 $Y=2.055 $X2=0 $Y2=0
cc_124 N_A_84_21#_c_109_n N_B1_c_356_n 5.91512e-19 $X=3.405 $Y=2.055 $X2=0 $Y2=0
cc_125 N_A_84_21#_c_109_n N_B1_c_357_n 0.0238034f $X=3.405 $Y=2.055 $X2=0 $Y2=0
cc_126 N_A_84_21#_c_109_n N_C1_c_409_n 0.0134873f $X=3.405 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_84_21#_c_111_n N_C1_c_409_n 0.0260163f $X=3.82 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_84_21#_c_111_n N_C1_c_410_n 0.0190449f $X=3.82 $Y=2.055 $X2=0 $Y2=0
cc_129 N_A_84_21#_c_109_n N_C1_c_411_n 0.00393921f $X=3.405 $Y=2.055 $X2=0 $Y2=0
cc_130 N_A_84_21#_c_111_n N_C1_c_411_n 0.00133018f $X=3.82 $Y=2.055 $X2=0 $Y2=0
cc_131 N_A_84_21#_c_100_n N_C1_M1012_g 0.00793322f $X=3.82 $Y=1.97 $X2=0 $Y2=0
cc_132 N_A_84_21#_c_100_n N_C1_c_412_n 0.00704815f $X=3.82 $Y=1.97 $X2=0 $Y2=0
cc_133 N_A_84_21#_c_111_n N_C1_c_407_n 0.00257951f $X=3.82 $Y=2.055 $X2=0 $Y2=0
cc_134 N_A_84_21#_c_100_n N_C1_c_407_n 0.00790613f $X=3.82 $Y=1.97 $X2=0 $Y2=0
cc_135 N_A_84_21#_c_101_n N_C1_c_407_n 0.00248562f $X=4.15 $Y=0.85 $X2=0 $Y2=0
cc_136 N_A_84_21#_c_111_n N_C1_c_408_n 0.0322105f $X=3.82 $Y=2.055 $X2=0 $Y2=0
cc_137 N_A_84_21#_c_100_n N_C1_c_408_n 0.0356132f $X=3.82 $Y=1.97 $X2=0 $Y2=0
cc_138 N_A_84_21#_c_101_n N_C1_c_408_n 0.00118166f $X=4.15 $Y=0.85 $X2=0 $Y2=0
cc_139 N_A_84_21#_M1000_g N_X_c_452_n 0.0244405f $X=0.59 $Y=2.595 $X2=0 $Y2=0
cc_140 N_A_84_21#_c_105_n N_X_c_452_n 0.00155244f $X=0.6 $Y=1.895 $X2=0 $Y2=0
cc_141 N_A_84_21#_c_106_n N_X_c_452_n 0.0082319f $X=0.645 $Y=1.7 $X2=0 $Y2=0
cc_142 N_A_84_21#_M1000_g N_X_c_449_n 0.00296539f $X=0.59 $Y=2.595 $X2=0 $Y2=0
cc_143 N_A_84_21#_c_106_n N_X_c_449_n 0.0193749f $X=0.645 $Y=1.7 $X2=0 $Y2=0
cc_144 N_A_84_21#_c_98_n N_X_c_449_n 0.0345603f $X=0.615 $Y=1.39 $X2=0 $Y2=0
cc_145 N_A_84_21#_c_102_n N_X_c_449_n 0.0210611f $X=0.6 $Y=1.225 $X2=0 $Y2=0
cc_146 N_A_84_21#_c_93_n X 0.00938353f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_147 N_A_84_21#_c_96_n X 0.00138622f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_148 N_A_84_21#_c_97_n X 0.00928413f $X=0.495 $Y=0.805 $X2=0 $Y2=0
cc_149 N_A_84_21#_c_97_n X 8.13208e-19 $X=0.495 $Y=0.805 $X2=0 $Y2=0
cc_150 N_A_84_21#_c_102_n X 0.0120203f $X=0.6 $Y=1.225 $X2=0 $Y2=0
cc_151 N_A_84_21#_c_106_n N_VPWR_M1000_d 7.70949e-19 $X=0.645 $Y=1.7 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_84_21#_c_108_n N_VPWR_M1000_d 0.00291474f $X=1.815 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A_84_21#_c_109_n N_VPWR_M1004_d 0.00180746f $X=3.405 $Y=2.055 $X2=0
+ $Y2=0
cc_154 N_A_84_21#_M1000_g N_VPWR_c_476_n 0.0205273f $X=0.59 $Y=2.595 $X2=0 $Y2=0
cc_155 N_A_84_21#_c_106_n N_VPWR_c_476_n 0.00777197f $X=0.645 $Y=1.7 $X2=0 $Y2=0
cc_156 N_A_84_21#_c_108_n N_VPWR_c_476_n 0.0139187f $X=1.815 $Y=2.055 $X2=0
+ $Y2=0
cc_157 N_A_84_21#_c_109_n N_VPWR_c_477_n 0.0163515f $X=3.405 $Y=2.055 $X2=0
+ $Y2=0
cc_158 N_A_84_21#_c_111_n N_VPWR_c_477_n 0.0519685f $X=3.82 $Y=2.055 $X2=0 $Y2=0
cc_159 N_A_84_21#_c_117_p N_VPWR_c_478_n 0.0183971f $X=1.98 $Y=2.24 $X2=0 $Y2=0
cc_160 N_A_84_21#_c_111_n N_VPWR_c_479_n 0.0534703f $X=3.82 $Y=2.055 $X2=0 $Y2=0
cc_161 N_A_84_21#_M1001_d N_VPWR_c_475_n 0.00308191f $X=1.84 $Y=2.095 $X2=0
+ $Y2=0
cc_162 N_A_84_21#_M1010_d N_VPWR_c_475_n 0.0023218f $X=3.43 $Y=2.095 $X2=0 $Y2=0
cc_163 N_A_84_21#_M1000_g N_VPWR_c_475_n 0.0145619f $X=0.59 $Y=2.595 $X2=0 $Y2=0
cc_164 N_A_84_21#_c_117_p N_VPWR_c_475_n 0.012508f $X=1.98 $Y=2.24 $X2=0 $Y2=0
cc_165 N_A_84_21#_c_111_n N_VPWR_c_475_n 0.0318546f $X=3.82 $Y=2.055 $X2=0 $Y2=0
cc_166 N_A_84_21#_M1000_g N_VPWR_c_481_n 0.00840199f $X=0.59 $Y=2.595 $X2=0
+ $Y2=0
cc_167 N_A_84_21#_c_108_n A_270_419# 0.0048076f $X=1.815 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_168 N_A_84_21#_c_109_n A_482_419# 0.0048076f $X=3.405 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_84_21#_c_93_n N_VGND_c_524_n 0.00237616f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_170 N_A_84_21#_c_96_n N_VGND_c_524_n 0.0130491f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_171 N_A_84_21#_c_93_n N_VGND_c_525_n 0.00549284f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_172 N_A_84_21#_c_95_n N_VGND_c_525_n 4.87571e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_173 N_A_84_21#_c_96_n N_VGND_c_525_n 0.00486043f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_174 N_A_84_21#_c_101_n N_VGND_c_528_n 0.0061111f $X=4.15 $Y=0.85 $X2=0 $Y2=0
cc_175 N_A_84_21#_c_93_n N_VGND_c_529_n 0.010905f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_176 N_A_84_21#_c_95_n N_VGND_c_529_n 6.51792e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_177 N_A_84_21#_c_96_n N_VGND_c_529_n 0.00814425f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_178 N_A_84_21#_c_101_n N_VGND_c_529_n 0.0104557f $X=4.15 $Y=0.85 $X2=0 $Y2=0
cc_179 N_A_84_21#_c_96_n N_A_272_47#_c_576_n 3.33295e-19 $X=0.855 $Y=0.73 $X2=0
+ $Y2=0
cc_180 N_A_84_21#_c_100_n N_A_490_141#_c_612_n 0.00642832f $X=3.82 $Y=1.97 $X2=0
+ $Y2=0
cc_181 N_A1_M1005_g N_A2_M1001_g 0.0294157f $X=1.225 $Y=2.595 $X2=0 $Y2=0
cc_182 N_A1_c_202_n N_A2_M1006_g 0.0117382f $X=1.185 $Y=1.12 $X2=0 $Y2=0
cc_183 N_A1_c_205_n N_A2_M1006_g 0.0194288f $X=1.28 $Y=0.73 $X2=0 $Y2=0
cc_184 N_A1_c_203_n N_A2_c_254_n 0.0294157f $X=1.185 $Y=1.625 $X2=0 $Y2=0
cc_185 N_A1_c_204_n N_A2_c_255_n 0.0294157f $X=1.185 $Y=1.79 $X2=0 $Y2=0
cc_186 A1 A2 0.0441456f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_187 N_A1_c_208_n A2 0.00403875f $X=1.185 $Y=1.285 $X2=0 $Y2=0
cc_188 A1 N_A2_c_257_n 8.15016e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A1_c_208_n N_A2_c_257_n 0.0294157f $X=1.185 $Y=1.285 $X2=0 $Y2=0
cc_190 N_A1_M1005_g N_X_c_452_n 9.36767e-19 $X=1.225 $Y=2.595 $X2=0 $Y2=0
cc_191 N_A1_M1005_g N_VPWR_c_476_n 0.0246622f $X=1.225 $Y=2.595 $X2=0 $Y2=0
cc_192 N_A1_M1005_g N_VPWR_c_478_n 0.00975641f $X=1.225 $Y=2.595 $X2=0 $Y2=0
cc_193 N_A1_M1005_g N_VPWR_c_475_n 0.0173141f $X=1.225 $Y=2.595 $X2=0 $Y2=0
cc_194 N_A1_c_205_n N_VGND_c_524_n 0.00309362f $X=1.28 $Y=0.73 $X2=0 $Y2=0
cc_195 A1 N_VGND_c_524_n 0.0057474f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A1_c_208_n N_VGND_c_524_n 9.09981e-19 $X=1.185 $Y=1.285 $X2=0 $Y2=0
cc_197 N_A1_c_205_n N_VGND_c_527_n 0.00549284f $X=1.28 $Y=0.73 $X2=0 $Y2=0
cc_198 N_A1_c_206_n N_VGND_c_527_n 2.07025e-19 $X=1.28 $Y=0.88 $X2=0 $Y2=0
cc_199 N_A1_c_205_n N_VGND_c_529_n 0.0100259f $X=1.28 $Y=0.73 $X2=0 $Y2=0
cc_200 N_A1_c_206_n N_VGND_c_529_n 2.72728e-19 $X=1.28 $Y=0.88 $X2=0 $Y2=0
cc_201 N_A1_c_205_n N_A_272_47#_c_576_n 0.00671522f $X=1.28 $Y=0.73 $X2=0 $Y2=0
cc_202 A1 N_A_272_47#_c_576_n 5.26502e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A2_M1001_g N_B2_M1008_g 0.0285443f $X=1.715 $Y=2.595 $X2=0 $Y2=0
cc_204 N_A2_c_255_n N_B2_M1008_g 0.0103374f $X=1.755 $Y=1.79 $X2=0 $Y2=0
cc_205 N_A2_M1006_g N_B2_c_298_n 0.0190009f $X=1.715 $Y=0.445 $X2=0 $Y2=0
cc_206 N_A2_c_254_n B2 0.00276239f $X=1.755 $Y=1.625 $X2=0 $Y2=0
cc_207 A2 B2 0.0320869f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_208 N_A2_c_254_n N_B2_c_301_n 0.0103374f $X=1.755 $Y=1.625 $X2=0 $Y2=0
cc_209 A2 N_B2_c_301_n 3.57277e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_210 A2 N_B2_c_302_n 0.00144111f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_211 N_A2_c_257_n N_B2_c_302_n 0.0118684f $X=1.755 $Y=1.285 $X2=0 $Y2=0
cc_212 N_A2_M1001_g N_VPWR_c_478_n 0.00939541f $X=1.715 $Y=2.595 $X2=0 $Y2=0
cc_213 N_A2_M1001_g N_VPWR_c_475_n 0.0162464f $X=1.715 $Y=2.595 $X2=0 $Y2=0
cc_214 N_A2_M1006_g N_VGND_c_527_n 0.00404158f $X=1.715 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A2_M1006_g N_VGND_c_529_n 0.00704786f $X=1.715 $Y=0.445 $X2=0 $Y2=0
cc_216 N_A2_M1006_g N_VGND_c_530_n 0.00704561f $X=1.715 $Y=0.445 $X2=0 $Y2=0
cc_217 N_A2_M1006_g N_A_272_47#_c_575_n 0.0104473f $X=1.715 $Y=0.445 $X2=0 $Y2=0
cc_218 A2 N_A_272_47#_c_575_n 0.00799001f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_219 N_A2_c_257_n N_A_272_47#_c_575_n 0.00208992f $X=1.755 $Y=1.285 $X2=0
+ $Y2=0
cc_220 N_A2_M1006_g N_A_272_47#_c_576_n 0.00989668f $X=1.715 $Y=0.445 $X2=0
+ $Y2=0
cc_221 A2 N_A_272_47#_c_576_n 0.00440685f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_222 N_A2_c_257_n N_A_272_47#_c_576_n 3.26907e-19 $X=1.755 $Y=1.285 $X2=0
+ $Y2=0
cc_223 A2 N_A_490_141#_c_613_n 0.00128369f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_224 N_B2_M1008_g N_B1_c_358_n 0.070789f $X=2.285 $Y=2.595 $X2=-0.19
+ $Y2=-0.245
cc_225 N_B2_c_299_n N_B1_c_358_n 2.09346e-19 $X=2.805 $Y=0.63 $X2=-0.19
+ $Y2=-0.245
cc_226 B2 N_B1_c_358_n 0.00238828f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_227 N_B2_c_299_n N_B1_c_354_n 0.00804921f $X=2.805 $Y=0.63 $X2=0 $Y2=0
cc_228 B2 N_B1_c_354_n 0.00459589f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_229 N_B2_c_301_n N_B1_c_354_n 0.0106977f $X=2.325 $Y=1.56 $X2=0 $Y2=0
cc_230 N_B2_c_297_n N_B1_M1011_g 0.020924f $X=2.73 $Y=0.555 $X2=0 $Y2=0
cc_231 N_B2_M1008_g N_B1_c_360_n 0.0100978f $X=2.285 $Y=2.595 $X2=0 $Y2=0
cc_232 B2 N_B1_c_360_n 0.00306869f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_233 B2 N_B1_c_356_n 4.86866e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_234 N_B2_c_301_n N_B1_c_356_n 0.00163382f $X=2.325 $Y=1.56 $X2=0 $Y2=0
cc_235 N_B2_c_302_n N_B1_c_356_n 6.94491e-19 $X=2.325 $Y=1.395 $X2=0 $Y2=0
cc_236 B2 N_B1_c_357_n 0.0246359f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_237 N_B2_c_301_n N_B1_c_357_n 3.76804e-19 $X=2.325 $Y=1.56 $X2=0 $Y2=0
cc_238 N_B2_c_302_n N_B1_c_357_n 0.00102635f $X=2.325 $Y=1.395 $X2=0 $Y2=0
cc_239 N_B2_M1008_g N_VPWR_c_477_n 0.00425608f $X=2.285 $Y=2.595 $X2=0 $Y2=0
cc_240 N_B2_M1008_g N_VPWR_c_478_n 0.00975641f $X=2.285 $Y=2.595 $X2=0 $Y2=0
cc_241 N_B2_M1008_g N_VPWR_c_475_n 0.0170985f $X=2.285 $Y=2.595 $X2=0 $Y2=0
cc_242 N_B2_c_298_n N_VGND_c_528_n 0.0129808f $X=2.375 $Y=0.555 $X2=0 $Y2=0
cc_243 N_B2_c_298_n N_VGND_c_529_n 0.0195233f $X=2.375 $Y=0.555 $X2=0 $Y2=0
cc_244 N_B2_c_297_n N_A_272_47#_c_575_n 0.0140468f $X=2.73 $Y=0.555 $X2=0 $Y2=0
cc_245 N_B2_c_298_n N_A_272_47#_c_575_n 0.00458948f $X=2.375 $Y=0.555 $X2=0
+ $Y2=0
cc_246 N_B2_c_299_n N_A_272_47#_c_575_n 0.00546043f $X=2.805 $Y=0.63 $X2=0 $Y2=0
cc_247 N_B2_c_301_n N_A_272_47#_c_575_n 0.00287046f $X=2.325 $Y=1.56 $X2=0 $Y2=0
cc_248 N_B2_c_302_n N_A_272_47#_c_575_n 0.0103161f $X=2.325 $Y=1.395 $X2=0 $Y2=0
cc_249 N_B2_c_298_n N_A_272_47#_c_576_n 4.39627e-19 $X=2.375 $Y=0.555 $X2=0
+ $Y2=0
cc_250 N_B2_c_297_n N_A_272_47#_c_577_n 4.0343e-19 $X=2.73 $Y=0.555 $X2=0 $Y2=0
cc_251 N_B2_c_299_n N_A_490_141#_c_612_n 0.00927174f $X=2.805 $Y=0.63 $X2=0
+ $Y2=0
cc_252 B2 N_A_490_141#_c_612_n 6.01221e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_253 N_B2_c_297_n N_A_490_141#_c_613_n 0.00103289f $X=2.73 $Y=0.555 $X2=0
+ $Y2=0
cc_254 N_B2_c_299_n N_A_490_141#_c_613_n 0.003715f $X=2.805 $Y=0.63 $X2=0 $Y2=0
cc_255 B2 N_A_490_141#_c_613_n 0.0213862f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_256 N_B2_c_301_n N_A_490_141#_c_613_n 0.0013927f $X=2.325 $Y=1.56 $X2=0 $Y2=0
cc_257 N_B2_c_302_n N_A_490_141#_c_613_n 0.00692472f $X=2.325 $Y=1.395 $X2=0
+ $Y2=0
cc_258 N_B1_c_358_n N_C1_c_409_n 0.015092f $X=2.775 $Y=2.09 $X2=-0.19 $Y2=-0.245
cc_259 N_B1_c_360_n N_C1_c_411_n 0.015092f $X=2.775 $Y=1.965 $X2=0 $Y2=0
cc_260 N_B1_c_356_n N_C1_c_411_n 0.0160097f $X=3.245 $Y=1.495 $X2=0 $Y2=0
cc_261 N_B1_c_357_n N_C1_c_411_n 0.00117742f $X=3.245 $Y=1.495 $X2=0 $Y2=0
cc_262 N_B1_M1011_g N_C1_M1012_g 0.0222589f $X=3.315 $Y=0.82 $X2=0 $Y2=0
cc_263 N_B1_c_357_n N_C1_c_412_n 5.96066e-19 $X=3.245 $Y=1.495 $X2=0 $Y2=0
cc_264 N_B1_c_356_n N_C1_c_407_n 0.020923f $X=3.245 $Y=1.495 $X2=0 $Y2=0
cc_265 N_B1_c_357_n N_C1_c_407_n 2.86728e-19 $X=3.245 $Y=1.495 $X2=0 $Y2=0
cc_266 N_B1_c_360_n N_C1_c_408_n 3.65371e-19 $X=2.775 $Y=1.965 $X2=0 $Y2=0
cc_267 N_B1_c_356_n N_C1_c_408_n 0.00231535f $X=3.245 $Y=1.495 $X2=0 $Y2=0
cc_268 N_B1_c_357_n N_C1_c_408_n 0.0366748f $X=3.245 $Y=1.495 $X2=0 $Y2=0
cc_269 N_B1_c_358_n N_VPWR_c_477_n 0.021443f $X=2.775 $Y=2.09 $X2=0 $Y2=0
cc_270 N_B1_c_358_n N_VPWR_c_478_n 0.008763f $X=2.775 $Y=2.09 $X2=0 $Y2=0
cc_271 N_B1_c_358_n N_VPWR_c_475_n 0.0144563f $X=2.775 $Y=2.09 $X2=0 $Y2=0
cc_272 N_B1_M1011_g N_VGND_c_528_n 0.00406951f $X=3.315 $Y=0.82 $X2=0 $Y2=0
cc_273 N_B1_M1011_g N_VGND_c_529_n 0.00473597f $X=3.315 $Y=0.82 $X2=0 $Y2=0
cc_274 N_B1_M1011_g N_A_272_47#_c_577_n 0.00536117f $X=3.315 $Y=0.82 $X2=0 $Y2=0
cc_275 N_B1_c_353_n N_A_490_141#_c_612_n 3.40597e-19 $X=3.08 $Y=1.585 $X2=0
+ $Y2=0
cc_276 N_B1_c_354_n N_A_490_141#_c_612_n 0.0043925f $X=2.9 $Y=1.585 $X2=0 $Y2=0
cc_277 N_B1_M1011_g N_A_490_141#_c_612_n 0.0155715f $X=3.315 $Y=0.82 $X2=0 $Y2=0
cc_278 N_B1_c_356_n N_A_490_141#_c_612_n 0.00187924f $X=3.245 $Y=1.495 $X2=0
+ $Y2=0
cc_279 N_B1_c_357_n N_A_490_141#_c_612_n 0.0249695f $X=3.245 $Y=1.495 $X2=0
+ $Y2=0
cc_280 N_B1_M1011_g N_A_490_141#_c_613_n 4.47088e-19 $X=3.315 $Y=0.82 $X2=0
+ $Y2=0
cc_281 N_C1_c_409_n N_VPWR_c_477_n 0.0203301f $X=3.305 $Y=2.02 $X2=0 $Y2=0
cc_282 N_C1_c_409_n N_VPWR_c_479_n 0.00840199f $X=3.305 $Y=2.02 $X2=0 $Y2=0
cc_283 N_C1_c_409_n N_VPWR_c_475_n 0.0148971f $X=3.305 $Y=2.02 $X2=0 $Y2=0
cc_284 N_C1_M1012_g N_VGND_c_528_n 0.00408363f $X=3.745 $Y=0.82 $X2=0 $Y2=0
cc_285 N_C1_M1012_g N_VGND_c_529_n 0.00473597f $X=3.745 $Y=0.82 $X2=0 $Y2=0
cc_286 N_C1_M1012_g N_A_272_47#_c_577_n 6.1786e-19 $X=3.745 $Y=0.82 $X2=0 $Y2=0
cc_287 N_C1_M1012_g N_A_490_141#_c_612_n 0.00441304f $X=3.745 $Y=0.82 $X2=0
+ $Y2=0
cc_288 N_C1_c_407_n N_A_490_141#_c_612_n 0.00115099f $X=3.785 $Y=1.495 $X2=0
+ $Y2=0
cc_289 N_C1_c_408_n N_A_490_141#_c_612_n 0.0167631f $X=3.785 $Y=1.495 $X2=0
+ $Y2=0
cc_290 N_C1_M1012_g N_A_490_141#_c_632_n 0.00367452f $X=3.745 $Y=0.82 $X2=0
+ $Y2=0
cc_291 N_X_c_452_n N_VPWR_c_476_n 0.0497241f $X=0.325 $Y=2.24 $X2=0 $Y2=0
cc_292 N_X_M1000_s N_VPWR_c_475_n 0.0023218f $X=0.18 $Y=2.095 $X2=0 $Y2=0
cc_293 N_X_c_452_n N_VPWR_c_475_n 0.0148296f $X=0.325 $Y=2.24 $X2=0 $Y2=0
cc_294 N_X_c_452_n N_VPWR_c_481_n 0.0238035f $X=0.325 $Y=2.24 $X2=0 $Y2=0
cc_295 X N_VGND_c_524_n 0.0134787f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_296 X N_VGND_c_525_n 0.0207998f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_297 N_X_M1002_s N_VGND_c_529_n 0.00232985f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_298 X N_VGND_c_529_n 0.0131612f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_299 N_VPWR_c_475_n A_270_419# 0.010279f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_300 N_VPWR_c_475_n A_482_419# 0.010279f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_301 A_114_47# N_VGND_c_529_n 0.00829524f $X=0.57 $Y=0.235 $X2=4.08 $Y2=0
cc_302 N_VGND_c_529_n N_A_272_47#_M1003_d 0.0022543f $X=4.08 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_303 N_VGND_M1006_d N_A_272_47#_c_575_n 0.00355566f $X=1.79 $Y=0.235 $X2=0
+ $Y2=0
cc_304 N_VGND_c_527_n N_A_272_47#_c_575_n 0.0032306f $X=1.845 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_c_528_n N_A_272_47#_c_575_n 0.0156678f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_c_529_n N_A_272_47#_c_575_n 0.0293367f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_530_n N_A_272_47#_c_575_n 0.0229917f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_308 N_VGND_c_524_n N_A_272_47#_c_576_n 0.0154229f $X=1.07 $Y=0.445 $X2=0
+ $Y2=0
cc_309 N_VGND_c_527_n N_A_272_47#_c_576_n 0.017446f $X=1.845 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_529_n N_A_272_47#_c_576_n 0.0123326f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_528_n N_A_272_47#_c_577_n 0.00754795f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_529_n N_A_272_47#_c_577_n 0.0102137f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_313 N_VGND_c_528_n N_A_490_141#_c_632_n 0.00367358f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_314 N_VGND_c_529_n N_A_490_141#_c_632_n 0.00708243f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_315 N_A_272_47#_c_575_n N_A_490_141#_M1007_s 0.00239779f $X=2.935 $Y=0.63
+ $X2=-0.19 $Y2=-0.245
cc_316 N_A_272_47#_M1007_d N_A_490_141#_c_612_n 0.00261503f $X=2.88 $Y=0.705
+ $X2=0 $Y2=0
cc_317 N_A_272_47#_c_575_n N_A_490_141#_c_612_n 0.00576904f $X=2.935 $Y=0.63
+ $X2=0 $Y2=0
cc_318 N_A_272_47#_c_577_n N_A_490_141#_c_612_n 0.0202883f $X=3.1 $Y=0.63 $X2=0
+ $Y2=0
cc_319 N_A_272_47#_c_575_n N_A_490_141#_c_613_n 0.0195191f $X=2.935 $Y=0.63
+ $X2=0 $Y2=0
