* File: sky130_fd_sc_lp__buf_16.pex.spice
* Created: Wed Sep  2 09:34:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUF_16%A 3 7 11 15 19 23 27 31 35 39 43 47 49 59 62
+ 76
c114 62 0 2.47794e-20 $X=2.16 $Y=1.295
c115 59 0 1.67963e-19 $X=2.57 $Y=1.48
r116 73 82 0.164635 $w=3.48e-07 $l=5e-09 $layer=LI1_cond $X=2.08 $Y=1.48
+ $X2=2.08 $Y2=1.485
r117 72 74 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=2.23 $Y=1.48
+ $X2=2.295 $Y2=1.48
r118 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.48 $X2=2.23 $Y2=1.48
r119 68 69 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.435 $Y=1.48
+ $X2=1.865 $Y2=1.48
r120 67 68 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.005 $Y=1.48
+ $X2=1.435 $Y2=1.48
r121 66 67 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.575 $Y=1.48
+ $X2=1.005 $Y2=1.48
r122 62 73 6.09148 $w=3.48e-07 $l=1.85e-07 $layer=LI1_cond $X=2.08 $Y=1.295
+ $X2=2.08 $Y2=1.48
r123 60 76 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.57 $Y=1.48
+ $X2=2.725 $Y2=1.48
r124 60 74 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=2.57 $Y=1.48
+ $X2=2.295 $Y2=1.48
r125 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.48 $X2=2.57 $Y2=1.48
r126 57 82 4.01183 $w=2e-07 $l=1.75e-07 $layer=LI1_cond $X=2.255 $Y=1.485
+ $X2=2.08 $Y2=1.485
r127 57 59 17.4682 $w=1.98e-07 $l=3.15e-07 $layer=LI1_cond $X=2.255 $Y=1.485
+ $X2=2.57 $Y2=1.485
r128 56 72 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.89 $Y=1.48
+ $X2=2.23 $Y2=1.48
r129 56 69 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.89 $Y=1.48
+ $X2=1.865 $Y2=1.48
r130 55 56 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.89
+ $Y=1.48 $X2=1.89 $Y2=1.48
r131 52 66 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=0.53 $Y=1.48
+ $X2=0.575 $Y2=1.48
r132 51 55 75.4182 $w=1.98e-07 $l=1.36e-06 $layer=LI1_cond $X=0.53 $Y=1.485
+ $X2=1.89 $Y2=1.485
r133 51 52 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.53
+ $Y=1.48 $X2=0.53 $Y2=1.48
r134 49 82 4.01183 $w=2e-07 $l=1.75e-07 $layer=LI1_cond $X=1.905 $Y=1.485
+ $X2=2.08 $Y2=1.485
r135 49 55 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.905 $Y=1.485
+ $X2=1.89 $Y2=1.485
r136 45 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.645
+ $X2=2.725 $Y2=1.48
r137 45 47 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.725 $Y=1.645
+ $X2=2.725 $Y2=2.465
r138 41 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.315
+ $X2=2.725 $Y2=1.48
r139 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.725 $Y=1.315
+ $X2=2.725 $Y2=0.655
r140 37 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.645
+ $X2=2.295 $Y2=1.48
r141 37 39 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.295 $Y=1.645
+ $X2=2.295 $Y2=2.465
r142 33 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.315
+ $X2=2.295 $Y2=1.48
r143 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.295 $Y=1.315
+ $X2=2.295 $Y2=0.655
r144 29 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.645
+ $X2=1.865 $Y2=1.48
r145 29 31 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.865 $Y=1.645
+ $X2=1.865 $Y2=2.465
r146 25 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.315
+ $X2=1.865 $Y2=1.48
r147 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.865 $Y=1.315
+ $X2=1.865 $Y2=0.655
r148 21 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.645
+ $X2=1.435 $Y2=1.48
r149 21 23 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.435 $Y=1.645
+ $X2=1.435 $Y2=2.465
r150 17 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.315
+ $X2=1.435 $Y2=1.48
r151 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.435 $Y=1.315
+ $X2=1.435 $Y2=0.655
r152 13 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.645
+ $X2=1.005 $Y2=1.48
r153 13 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.005 $Y=1.645
+ $X2=1.005 $Y2=2.465
r154 9 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.315
+ $X2=1.005 $Y2=1.48
r155 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.005 $Y=1.315
+ $X2=1.005 $Y2=0.655
r156 5 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.645
+ $X2=0.575 $Y2=1.48
r157 5 7 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.575 $Y=1.645
+ $X2=0.575 $Y2=2.465
r158 1 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.315
+ $X2=0.575 $Y2=1.48
r159 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.575 $Y=1.315
+ $X2=0.575 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_16%A_130_47# 1 2 3 4 5 6 21 23 25 28 30 32 35 39
+ 43 47 51 55 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 131
+ 135 139 141 143 147 151 155 156 157 158 161 167 169 171 175 181 183 185 187
+ 188 190 191 197 218 225 230 235 240 245 250 255
c375 218 0 2.47794e-20 $X=8.96 $Y=1.665
c376 185 0 1.55749e-19 $X=2.905 $Y=1.84
c377 141 0 1.67963e-19 $X=9.605 $Y=1.655
r378 254 255 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.96
+ $Y=1.49 $X2=8.96 $Y2=1.49
r379 249 250 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.1
+ $Y=1.49 $X2=8.1 $Y2=1.49
r380 244 245 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.24
+ $Y=1.49 $X2=7.24 $Y2=1.49
r381 239 240 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.38
+ $Y=1.49 $X2=6.38 $Y2=1.49
r382 234 235 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.52
+ $Y=1.49 $X2=5.52 $Y2=1.49
r383 229 230 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.66
+ $Y=1.49 $X2=4.66 $Y2=1.49
r384 224 225 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.8
+ $Y=1.49 $X2=3.8 $Y2=1.49
r385 222 224 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=3.585 $Y=1.525
+ $X2=3.8 $Y2=1.525
r386 221 222 61.8687 $w=3.35e-07 $l=4.3e-07 $layer=POLY_cond $X=3.155 $Y=1.525
+ $X2=3.585 $Y2=1.525
r387 219 255 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=8.96 $Y=1.665
+ $X2=8.96 $Y2=1.49
r388 218 219 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.96 $Y=1.665
+ $X2=8.96 $Y2=1.665
r389 216 250 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=8.1 $Y=1.665
+ $X2=8.1 $Y2=1.49
r390 215 218 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=8.1 $Y=1.665
+ $X2=8.96 $Y2=1.665
r391 215 216 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.1 $Y=1.665
+ $X2=8.1 $Y2=1.665
r392 213 245 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=7.24 $Y=1.665
+ $X2=7.24 $Y2=1.49
r393 212 215 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.24 $Y=1.665
+ $X2=8.1 $Y2=1.665
r394 212 213 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.24 $Y=1.665
+ $X2=7.24 $Y2=1.665
r395 210 240 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=6.38 $Y=1.665
+ $X2=6.38 $Y2=1.49
r396 209 212 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.38 $Y=1.665
+ $X2=7.24 $Y2=1.665
r397 209 210 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.38 $Y=1.665
+ $X2=6.38 $Y2=1.665
r398 207 235 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.49
r399 206 209 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=5.52 $Y=1.665
+ $X2=6.38 $Y2=1.665
r400 206 207 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r401 204 230 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=4.66 $Y=1.665
+ $X2=4.66 $Y2=1.49
r402 203 206 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=4.66 $Y=1.665
+ $X2=5.52 $Y2=1.665
r403 203 204 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.66 $Y=1.665
+ $X2=4.66 $Y2=1.665
r404 201 225 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=3.8 $Y=1.665
+ $X2=3.8 $Y2=1.49
r405 200 203 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=3.8 $Y=1.665
+ $X2=4.66 $Y2=1.665
r406 200 201 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.8 $Y=1.665
+ $X2=3.8 $Y2=1.665
r407 196 200 0.513283 $w=2.3e-07 $l=8e-07 $layer=MET1_cond $X=3 $Y=1.665 $X2=3.8
+ $Y2=1.665
r408 196 197 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3 $Y=1.665 $X2=3
+ $Y2=1.665
r409 194 197 5.25359 $w=1.88e-07 $l=9e-08 $layer=LI1_cond $X=3 $Y=1.755 $X2=3
+ $Y2=1.665
r410 193 197 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=3 $Y=1.215 $X2=3
+ $Y2=1.665
r411 191 192 10.0274 $w=2.19e-07 $l=1.8e-07 $layer=LI1_cond $X=2.527 $Y=0.95
+ $X2=2.527 $Y2=1.13
r412 188 189 10.5072 $w=2.09e-07 $l=1.8e-07 $layer=LI1_cond $X=1.637 $Y=0.95
+ $X2=1.637 $Y2=1.13
r413 186 190 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=1.84
+ $X2=2.51 $Y2=1.84
r414 185 194 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.905 $Y=1.84
+ $X2=3 $Y2=1.755
r415 185 186 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=1.84
+ $X2=2.64 $Y2=1.84
r416 184 192 2.22295 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=2.64 $Y=1.13
+ $X2=2.527 $Y2=1.13
r417 183 193 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.905 $Y=1.13
+ $X2=3 $Y2=1.215
r418 183 184 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=1.13
+ $X2=2.64 $Y2=1.13
r419 179 191 4.60889 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.527 $Y=0.865
+ $X2=2.527 $Y2=0.95
r420 179 181 14.0854 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=2.527 $Y=0.865
+ $X2=2.527 $Y2=0.59
r421 175 177 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=2.51 $Y=2.025
+ $X2=2.51 $Y2=2.865
r422 173 190 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.925
+ $X2=2.51 $Y2=1.84
r423 173 175 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=2.51 $Y=1.925
+ $X2=2.51 $Y2=2.025
r424 172 187 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.78 $Y=1.84
+ $X2=1.65 $Y2=1.84
r425 171 190 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.38 $Y=1.84
+ $X2=2.51 $Y2=1.84
r426 171 172 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.38 $Y=1.84
+ $X2=1.78 $Y2=1.84
r427 170 188 1.94907 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.745 $Y=0.95
+ $X2=1.637 $Y2=0.95
r428 169 191 2.22295 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=2.415 $Y=0.95
+ $X2=2.527 $Y2=0.95
r429 169 170 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.415 $Y=0.95
+ $X2=1.745 $Y2=0.95
r430 165 188 4.82326 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.637 $Y=0.865
+ $X2=1.637 $Y2=0.95
r431 165 167 14.7406 $w=2.13e-07 $l=2.75e-07 $layer=LI1_cond $X=1.637 $Y=0.865
+ $X2=1.637 $Y2=0.59
r432 161 163 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=1.65 $Y=2.025
+ $X2=1.65 $Y2=2.865
r433 159 187 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=1.925
+ $X2=1.65 $Y2=1.84
r434 159 161 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=1.65 $Y=1.925
+ $X2=1.65 $Y2=2.025
r435 157 187 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.52 $Y=1.84
+ $X2=1.65 $Y2=1.84
r436 157 158 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.52 $Y=1.84
+ $X2=0.92 $Y2=1.84
r437 155 189 1.94907 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.53 $Y=1.13
+ $X2=1.637 $Y2=1.13
r438 155 156 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.53 $Y=1.13
+ $X2=0.92 $Y2=1.13
r439 151 153 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=0.79 $Y=2.025
+ $X2=0.79 $Y2=2.865
r440 149 158 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.79 $Y=1.925
+ $X2=0.92 $Y2=1.84
r441 149 151 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=0.79 $Y=1.925
+ $X2=0.79 $Y2=2.025
r442 145 156 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.79 $Y=1.045
+ $X2=0.92 $Y2=1.13
r443 145 147 20.1678 $w=2.58e-07 $l=4.55e-07 $layer=LI1_cond $X=0.79 $Y=1.045
+ $X2=0.79 $Y2=0.59
r444 141 143 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.605 $Y=1.655
+ $X2=9.605 $Y2=2.465
r445 137 141 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=9.605 $Y=1.325
+ $X2=9.605 $Y2=1.525
r446 137 139 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=9.605 $Y=1.325
+ $X2=9.605 $Y2=0.655
r447 133 141 61.8687 $w=3.35e-07 $l=4.3e-07 $layer=POLY_cond $X=9.175 $Y=1.525
+ $X2=9.605 $Y2=1.525
r448 133 254 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=9.175 $Y=1.525
+ $X2=8.96 $Y2=1.525
r449 133 135 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.175 $Y=1.655
+ $X2=9.175 $Y2=2.465
r450 129 133 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=9.175 $Y=1.325
+ $X2=9.175 $Y2=1.525
r451 129 131 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=9.175 $Y=1.325
+ $X2=9.175 $Y2=0.655
r452 125 254 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=8.745 $Y=1.525
+ $X2=8.96 $Y2=1.525
r453 125 127 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=8.745 $Y=1.655
+ $X2=8.745 $Y2=2.465
r454 121 125 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=8.745 $Y=1.325
+ $X2=8.745 $Y2=1.525
r455 121 123 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=8.745 $Y=1.325
+ $X2=8.745 $Y2=0.655
r456 117 125 61.8687 $w=3.35e-07 $l=4.3e-07 $layer=POLY_cond $X=8.315 $Y=1.525
+ $X2=8.745 $Y2=1.525
r457 117 249 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=8.315 $Y=1.525
+ $X2=8.1 $Y2=1.525
r458 117 119 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=8.315 $Y=1.655
+ $X2=8.315 $Y2=2.465
r459 113 117 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=8.315 $Y=1.325
+ $X2=8.315 $Y2=1.525
r460 113 115 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=8.315 $Y=1.325
+ $X2=8.315 $Y2=0.655
r461 109 249 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=7.885 $Y=1.525
+ $X2=8.1 $Y2=1.525
r462 109 111 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.885 $Y=1.655
+ $X2=7.885 $Y2=2.465
r463 105 109 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.885 $Y=1.325
+ $X2=7.885 $Y2=1.525
r464 105 107 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.885 $Y=1.325
+ $X2=7.885 $Y2=0.655
r465 101 109 61.8687 $w=3.35e-07 $l=4.3e-07 $layer=POLY_cond $X=7.455 $Y=1.525
+ $X2=7.885 $Y2=1.525
r466 101 244 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=7.455 $Y=1.525
+ $X2=7.24 $Y2=1.525
r467 101 103 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.455 $Y=1.655
+ $X2=7.455 $Y2=2.465
r468 97 101 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.455 $Y=1.325
+ $X2=7.455 $Y2=1.525
r469 97 99 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.455 $Y=1.325
+ $X2=7.455 $Y2=0.655
r470 93 244 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=7.025 $Y=1.525
+ $X2=7.24 $Y2=1.525
r471 93 95 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.025 $Y=1.655
+ $X2=7.025 $Y2=2.465
r472 89 93 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.025 $Y=1.325
+ $X2=7.025 $Y2=1.525
r473 89 91 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.025 $Y=1.325
+ $X2=7.025 $Y2=0.655
r474 85 93 61.8687 $w=3.35e-07 $l=4.3e-07 $layer=POLY_cond $X=6.595 $Y=1.525
+ $X2=7.025 $Y2=1.525
r475 85 239 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=6.595 $Y=1.525
+ $X2=6.38 $Y2=1.525
r476 85 87 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.595 $Y=1.655
+ $X2=6.595 $Y2=2.465
r477 81 85 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=6.595 $Y=1.325
+ $X2=6.595 $Y2=1.525
r478 81 83 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.595 $Y=1.325
+ $X2=6.595 $Y2=0.655
r479 77 239 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=6.165 $Y=1.525
+ $X2=6.38 $Y2=1.525
r480 77 79 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.165 $Y=1.655
+ $X2=6.165 $Y2=2.465
r481 73 77 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=6.165 $Y=1.325
+ $X2=6.165 $Y2=1.525
r482 73 75 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.165 $Y=1.325
+ $X2=6.165 $Y2=0.655
r483 69 77 61.8687 $w=3.35e-07 $l=4.3e-07 $layer=POLY_cond $X=5.735 $Y=1.525
+ $X2=6.165 $Y2=1.525
r484 69 234 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=5.735 $Y=1.525
+ $X2=5.52 $Y2=1.525
r485 69 71 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.735 $Y=1.655
+ $X2=5.735 $Y2=2.465
r486 65 69 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.735 $Y=1.325
+ $X2=5.735 $Y2=1.525
r487 65 67 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.735 $Y=1.325
+ $X2=5.735 $Y2=0.655
r488 61 234 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=5.305 $Y=1.525
+ $X2=5.52 $Y2=1.525
r489 61 63 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.305 $Y=1.655
+ $X2=5.305 $Y2=2.465
r490 57 61 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.305 $Y=1.325
+ $X2=5.305 $Y2=1.525
r491 57 59 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.305 $Y=1.325
+ $X2=5.305 $Y2=0.655
r492 53 61 61.8687 $w=3.35e-07 $l=4.3e-07 $layer=POLY_cond $X=4.875 $Y=1.525
+ $X2=5.305 $Y2=1.525
r493 53 229 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=4.875 $Y=1.525
+ $X2=4.66 $Y2=1.525
r494 53 55 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.875 $Y=1.655
+ $X2=4.875 $Y2=2.465
r495 49 53 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=4.875 $Y=1.325
+ $X2=4.875 $Y2=1.525
r496 49 51 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=4.875 $Y=1.325
+ $X2=4.875 $Y2=0.655
r497 45 229 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=4.445 $Y=1.525
+ $X2=4.66 $Y2=1.525
r498 45 47 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.445 $Y=1.655
+ $X2=4.445 $Y2=2.465
r499 41 45 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=4.445 $Y=1.325
+ $X2=4.445 $Y2=1.525
r500 41 43 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=4.445 $Y=1.325
+ $X2=4.445 $Y2=0.655
r501 37 45 61.8687 $w=3.35e-07 $l=4.3e-07 $layer=POLY_cond $X=4.015 $Y=1.525
+ $X2=4.445 $Y2=1.525
r502 37 224 30.9343 $w=3.35e-07 $l=2.15e-07 $layer=POLY_cond $X=4.015 $Y=1.525
+ $X2=3.8 $Y2=1.525
r503 37 39 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.015 $Y=1.655
+ $X2=4.015 $Y2=2.465
r504 33 37 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=4.015 $Y=1.325
+ $X2=4.015 $Y2=1.525
r505 33 35 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=4.015 $Y=1.325
+ $X2=4.015 $Y2=0.655
r506 30 222 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.585 $Y=1.725
+ $X2=3.585 $Y2=1.525
r507 30 32 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.585 $Y=1.725
+ $X2=3.585 $Y2=2.465
r508 26 222 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.585 $Y=1.325
+ $X2=3.585 $Y2=1.525
r509 26 28 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=3.585 $Y=1.325
+ $X2=3.585 $Y2=0.655
r510 23 221 21.5811 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.155 $Y=1.725
+ $X2=3.155 $Y2=1.525
r511 23 25 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.155 $Y=1.725
+ $X2=3.155 $Y2=2.465
r512 19 221 21.5811 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.155 $Y=1.335
+ $X2=3.155 $Y2=1.525
r513 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.155 $Y=1.335
+ $X2=3.155 $Y2=0.655
r514 6 177 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.835 $X2=2.51 $Y2=2.865
r515 6 175 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.835 $X2=2.51 $Y2=2.025
r516 5 163 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.835 $X2=1.65 $Y2=2.865
r517 5 161 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.835 $X2=1.65 $Y2=2.025
r518 4 153 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.835 $X2=0.79 $Y2=2.865
r519 4 151 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.835 $X2=0.79 $Y2=2.025
r520 3 181 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=2.37
+ $Y=0.235 $X2=2.51 $Y2=0.59
r521 2 167 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.235 $X2=1.65 $Y2=0.59
r522 1 147 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=0.65
+ $Y=0.235 $X2=0.79 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 37 39 45 51
+ 57 63 67 71 77 83 89 95 99 103 107 109 114 115 117 118 119 120 122 123 125 126
+ 127 128 129 131 146 161 170 173 176 179 183
r199 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r200 179 180 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r201 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r202 173 174 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r203 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r204 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r205 165 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r206 165 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r207 164 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r208 162 179 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=8.96 $Y2=3.33
r209 162 164 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=9.36 $Y2=3.33
r210 161 182 4.44548 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=9.69 $Y=3.33
+ $X2=9.885 $Y2=3.33
r211 161 164 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.69 $Y=3.33
+ $X2=9.36 $Y2=3.33
r212 160 180 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r213 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r214 157 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r215 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r216 154 157 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r217 154 177 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r218 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r219 151 176 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.65 $Y=3.33
+ $X2=5.52 $Y2=3.33
r220 151 153 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.65 $Y=3.33
+ $X2=6 $Y2=3.33
r221 147 173 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.79 $Y=3.33
+ $X2=4.66 $Y2=3.33
r222 147 149 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.79 $Y=3.33
+ $X2=5.04 $Y2=3.33
r223 146 176 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.39 $Y=3.33
+ $X2=5.52 $Y2=3.33
r224 146 149 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.39 $Y=3.33
+ $X2=5.04 $Y2=3.33
r225 145 174 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r226 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r227 142 145 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r228 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r229 139 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r230 139 171 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r231 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r232 136 170 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.22 $Y2=3.33
r233 136 138 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.68 $Y2=3.33
r234 135 171 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r235 135 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r236 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r237 132 167 4.29038 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.49 $Y=3.33
+ $X2=0.245 $Y2=3.33
r238 132 134 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.49 $Y=3.33
+ $X2=0.72 $Y2=3.33
r239 131 170 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=1.22 $Y2=3.33
r240 131 134 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.72 $Y2=3.33
r241 129 177 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r242 129 174 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r243 129 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r244 127 159 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=7.97 $Y=3.33
+ $X2=7.92 $Y2=3.33
r245 127 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.97 $Y=3.33
+ $X2=8.1 $Y2=3.33
r246 125 156 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.11 $Y=3.33
+ $X2=6.96 $Y2=3.33
r247 125 126 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.11 $Y=3.33
+ $X2=7.24 $Y2=3.33
r248 124 159 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.37 $Y=3.33
+ $X2=7.92 $Y2=3.33
r249 124 126 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.37 $Y=3.33
+ $X2=7.24 $Y2=3.33
r250 122 153 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.25 $Y=3.33
+ $X2=6 $Y2=3.33
r251 122 123 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.25 $Y=3.33
+ $X2=6.38 $Y2=3.33
r252 121 156 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.51 $Y=3.33
+ $X2=6.96 $Y2=3.33
r253 121 123 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.51 $Y=3.33
+ $X2=6.38 $Y2=3.33
r254 119 144 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=3.33
+ $X2=3.6 $Y2=3.33
r255 119 120 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.67 $Y=3.33
+ $X2=3.8 $Y2=3.33
r256 117 141 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.81 $Y=3.33
+ $X2=2.64 $Y2=3.33
r257 117 118 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=2.81 $Y=3.33
+ $X2=2.952 $Y2=3.33
r258 116 144 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.6 $Y2=3.33
r259 116 118 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=2.952 $Y2=3.33
r260 114 138 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.95 $Y=3.33
+ $X2=1.68 $Y2=3.33
r261 114 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.95 $Y=3.33
+ $X2=2.08 $Y2=3.33
r262 113 141 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.21 $Y=3.33
+ $X2=2.64 $Y2=3.33
r263 113 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.21 $Y=3.33
+ $X2=2.08 $Y2=3.33
r264 109 112 31.448 $w=2.93e-07 $l=8.05e-07 $layer=LI1_cond $X=9.837 $Y=2.085
+ $X2=9.837 $Y2=2.89
r265 107 182 3.03205 $w=2.95e-07 $l=1.06325e-07 $layer=LI1_cond $X=9.837
+ $Y=3.245 $X2=9.885 $Y2=3.33
r266 107 112 13.8684 $w=2.93e-07 $l=3.55e-07 $layer=LI1_cond $X=9.837 $Y=3.245
+ $X2=9.837 $Y2=2.89
r267 103 106 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=8.96 $Y=2.085
+ $X2=8.96 $Y2=2.89
r268 101 179 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=3.245
+ $X2=8.96 $Y2=3.33
r269 101 106 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=8.96 $Y=3.245
+ $X2=8.96 $Y2=2.89
r270 100 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.23 $Y=3.33
+ $X2=8.1 $Y2=3.33
r271 99 179 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.83 $Y=3.33
+ $X2=8.96 $Y2=3.33
r272 99 100 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.83 $Y=3.33
+ $X2=8.23 $Y2=3.33
r273 95 98 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=8.1 $Y=2.085
+ $X2=8.1 $Y2=2.89
r274 93 128 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.1 $Y=3.245
+ $X2=8.1 $Y2=3.33
r275 93 98 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=8.1 $Y=3.245
+ $X2=8.1 $Y2=2.89
r276 89 92 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=7.24 $Y=2.085
+ $X2=7.24 $Y2=2.89
r277 87 126 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=3.245
+ $X2=7.24 $Y2=3.33
r278 87 92 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=7.24 $Y=3.245
+ $X2=7.24 $Y2=2.89
r279 83 86 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=6.38 $Y=2.085
+ $X2=6.38 $Y2=2.89
r280 81 123 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.38 $Y=3.245
+ $X2=6.38 $Y2=3.33
r281 81 86 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=6.38 $Y=3.245
+ $X2=6.38 $Y2=2.89
r282 77 80 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=5.52 $Y=2.085
+ $X2=5.52 $Y2=2.89
r283 75 176 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.52 $Y2=3.33
r284 75 80 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.52 $Y2=2.89
r285 71 74 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=4.66 $Y=2.085
+ $X2=4.66 $Y2=2.89
r286 69 173 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=3.245
+ $X2=4.66 $Y2=3.33
r287 69 74 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=4.66 $Y=3.245
+ $X2=4.66 $Y2=2.89
r288 68 120 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=3.8 $Y2=3.33
r289 67 173 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.53 $Y=3.33
+ $X2=4.66 $Y2=3.33
r290 67 68 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.53 $Y=3.33 $X2=3.93
+ $Y2=3.33
r291 63 66 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=3.8 $Y=2.085
+ $X2=3.8 $Y2=2.89
r292 61 120 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=3.245
+ $X2=3.8 $Y2=3.33
r293 61 66 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=3.8 $Y=3.245
+ $X2=3.8 $Y2=2.89
r294 57 60 27.4969 $w=2.83e-07 $l=6.8e-07 $layer=LI1_cond $X=2.952 $Y=2.26
+ $X2=2.952 $Y2=2.94
r295 55 118 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.952 $Y=3.245
+ $X2=2.952 $Y2=3.33
r296 55 60 12.3332 $w=2.83e-07 $l=3.05e-07 $layer=LI1_cond $X=2.952 $Y=3.245
+ $X2=2.952 $Y2=2.94
r297 51 54 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=2.08 $Y=2.26
+ $X2=2.08 $Y2=2.94
r298 49 115 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=3.33
r299 49 54 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=2.94
r300 45 48 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.22 $Y=2.26
+ $X2=1.22 $Y2=2.94
r301 43 170 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r302 43 48 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.94
r303 39 42 32.8153 $w=2.93e-07 $l=8.4e-07 $layer=LI1_cond $X=0.342 $Y=2.025
+ $X2=0.342 $Y2=2.865
r304 37 167 3.18714 $w=2.95e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.342 $Y=3.245
+ $X2=0.245 $Y2=3.33
r305 37 42 14.845 $w=2.93e-07 $l=3.8e-07 $layer=LI1_cond $X=0.342 $Y=3.245
+ $X2=0.342 $Y2=2.865
r306 12 112 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=2.89
r307 12 109 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=2.085
r308 11 106 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=8.82
+ $Y=1.835 $X2=8.96 $Y2=2.89
r309 11 103 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=8.82
+ $Y=1.835 $X2=8.96 $Y2=2.085
r310 10 98 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=7.96
+ $Y=1.835 $X2=8.1 $Y2=2.89
r311 10 95 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=7.96
+ $Y=1.835 $X2=8.1 $Y2=2.085
r312 9 92 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=1.835 $X2=7.24 $Y2=2.89
r313 9 89 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=1.835 $X2=7.24 $Y2=2.085
r314 8 86 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.835 $X2=6.38 $Y2=2.89
r315 8 83 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.835 $X2=6.38 $Y2=2.085
r316 7 80 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=5.38
+ $Y=1.835 $X2=5.52 $Y2=2.89
r317 7 77 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=5.38
+ $Y=1.835 $X2=5.52 $Y2=2.085
r318 6 74 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.835 $X2=4.66 $Y2=2.89
r319 6 71 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.835 $X2=4.66 $Y2=2.085
r320 5 66 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=1.835 $X2=3.8 $Y2=2.89
r321 5 63 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=1.835 $X2=3.8 $Y2=2.085
r322 4 60 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.835 $X2=2.94 $Y2=2.94
r323 4 57 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.835 $X2=2.94 $Y2=2.26
r324 3 54 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.08 $Y2=2.94
r325 3 51 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.08 $Y2=2.26
r326 2 48 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.22 $Y2=2.94
r327 2 45 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.22 $Y2=2.26
r328 1 42 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.835 $X2=0.36 $Y2=2.865
r329 1 39 400 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.835 $X2=0.36 $Y2=2.025
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 49
+ 52 62 72 82 92 102 112 122 127
c186 127 0 1.55749e-19 $X=9.39 $Y=2.035
r187 125 129 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=9.39 $Y=2.025
+ $X2=9.39 $Y2=2.865
r188 125 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.39 $Y=2.035
+ $X2=9.39 $Y2=2.035
r189 122 125 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=9.39 $Y=0.47
+ $X2=9.39 $Y2=2.025
r190 117 127 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=8.53 $Y=2.035
+ $X2=9.39 $Y2=2.035
r191 115 119 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=8.53 $Y=2.025
+ $X2=8.53 $Y2=2.865
r192 115 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.53 $Y=2.035
+ $X2=8.53 $Y2=2.035
r193 112 115 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=8.53 $Y=0.47
+ $X2=8.53 $Y2=2.025
r194 107 117 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.67 $Y=2.035
+ $X2=8.53 $Y2=2.035
r195 105 109 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=7.67 $Y=2.025
+ $X2=7.67 $Y2=2.865
r196 105 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.67 $Y=2.035
+ $X2=7.67 $Y2=2.035
r197 102 105 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=7.67 $Y=0.47
+ $X2=7.67 $Y2=2.025
r198 97 107 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.81 $Y=2.035
+ $X2=7.67 $Y2=2.035
r199 95 99 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=6.81 $Y=2.025
+ $X2=6.81 $Y2=2.865
r200 95 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.81 $Y=2.035
+ $X2=6.81 $Y2=2.035
r201 92 95 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=6.81 $Y=0.47
+ $X2=6.81 $Y2=2.025
r202 85 89 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=5.95 $Y=2.025
+ $X2=5.95 $Y2=2.865
r203 85 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.95 $Y=2.035
+ $X2=5.95 $Y2=2.035
r204 82 85 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=5.95 $Y=0.47
+ $X2=5.95 $Y2=2.025
r205 77 87 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=5.09 $Y=2.035
+ $X2=5.95 $Y2=2.035
r206 75 79 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=5.09 $Y=2.025
+ $X2=5.09 $Y2=2.865
r207 75 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.09 $Y=2.035
+ $X2=5.09 $Y2=2.035
r208 72 75 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=5.09 $Y=0.47
+ $X2=5.09 $Y2=2.025
r209 67 77 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=4.23 $Y=2.035
+ $X2=5.09 $Y2=2.035
r210 65 69 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=4.23 $Y=2.025
+ $X2=4.23 $Y2=2.865
r211 65 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.23 $Y=2.035
+ $X2=4.23 $Y2=2.035
r212 62 65 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=4.23 $Y=0.47
+ $X2=4.23 $Y2=2.025
r213 57 67 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=3.37 $Y=2.035
+ $X2=4.23 $Y2=2.035
r214 55 59 41.1937 $w=2.33e-07 $l=8.4e-07 $layer=LI1_cond $X=3.382 $Y=2.025
+ $X2=3.382 $Y2=2.865
r215 55 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.37 $Y=2.035
+ $X2=3.37 $Y2=2.035
r216 52 55 76.2574 $w=2.33e-07 $l=1.555e-06 $layer=LI1_cond $X=3.382 $Y=0.47
+ $X2=3.382 $Y2=2.025
r217 49 97 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=6.38 $Y=2.035
+ $X2=6.81 $Y2=2.035
r218 49 87 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=6.38 $Y=2.035
+ $X2=5.95 $Y2=2.035
r219 16 129 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=9.25
+ $Y=1.835 $X2=9.39 $Y2=2.865
r220 16 125 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=9.25
+ $Y=1.835 $X2=9.39 $Y2=2.025
r221 15 119 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=8.39
+ $Y=1.835 $X2=8.53 $Y2=2.865
r222 15 115 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=8.39
+ $Y=1.835 $X2=8.53 $Y2=2.025
r223 14 109 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=7.53
+ $Y=1.835 $X2=7.67 $Y2=2.865
r224 14 105 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=7.53
+ $Y=1.835 $X2=7.67 $Y2=2.025
r225 13 99 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=6.67
+ $Y=1.835 $X2=6.81 $Y2=2.865
r226 13 95 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=6.67
+ $Y=1.835 $X2=6.81 $Y2=2.025
r227 12 89 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=1.835 $X2=5.95 $Y2=2.865
r228 12 85 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=1.835 $X2=5.95 $Y2=2.025
r229 11 79 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.835 $X2=5.09 $Y2=2.865
r230 11 75 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.835 $X2=5.09 $Y2=2.025
r231 10 69 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=4.09
+ $Y=1.835 $X2=4.23 $Y2=2.865
r232 10 65 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=4.09
+ $Y=1.835 $X2=4.23 $Y2=2.025
r233 9 59 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.835 $X2=3.37 $Y2=2.865
r234 9 55 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.835 $X2=3.37 $Y2=2.025
r235 8 122 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=9.25
+ $Y=0.235 $X2=9.39 $Y2=0.47
r236 7 112 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=8.39
+ $Y=0.235 $X2=8.53 $Y2=0.47
r237 6 102 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=7.53
+ $Y=0.235 $X2=7.67 $Y2=0.47
r238 5 92 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=6.67
+ $Y=0.235 $X2=6.81 $Y2=0.47
r239 4 82 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.81
+ $Y=0.235 $X2=5.95 $Y2=0.47
r240 3 72 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.95
+ $Y=0.235 $X2=5.09 $Y2=0.47
r241 2 62 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.09
+ $Y=0.235 $X2=4.23 $Y2=0.47
r242 1 52 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=3.23
+ $Y=0.235 $X2=3.37 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 37 39 43 47
+ 51 55 57 61 65 69 73 77 79 83 85 87 90 91 92 93 95 96 98 99 100 101 102 104
+ 109 121 136 145 148 151 154 157 161
r167 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r168 157 158 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r169 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r170 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r171 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r172 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r173 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r174 140 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r175 140 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r176 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r177 137 157 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.09 $Y=0 $X2=8.96
+ $Y2=0
r178 137 139 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.09 $Y=0 $X2=9.36
+ $Y2=0
r179 136 160 4.44548 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=9.69 $Y=0
+ $X2=9.885 $Y2=0
r180 136 139 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.69 $Y=0
+ $X2=9.36 $Y2=0
r181 135 158 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.88 $Y2=0
r182 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r183 132 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.92 $Y2=0
r184 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r185 129 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r186 129 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r187 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r188 126 154 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.65 $Y=0 $X2=5.52
+ $Y2=0
r189 126 128 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.65 $Y=0 $X2=6
+ $Y2=0
r190 122 151 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.79 $Y=0 $X2=4.66
+ $Y2=0
r191 122 124 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.79 $Y=0
+ $X2=5.04 $Y2=0
r192 121 154 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.39 $Y=0 $X2=5.52
+ $Y2=0
r193 121 124 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.39 $Y=0
+ $X2=5.04 $Y2=0
r194 120 152 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.56 $Y2=0
r195 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r196 117 120 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r197 117 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r198 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r199 114 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.08 $Y2=0
r200 114 116 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.64 $Y2=0
r201 113 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r202 113 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=1.2 $Y2=0
r203 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r204 110 145 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.36 $Y=0
+ $X2=1.225 $Y2=0
r205 110 112 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.36 $Y=0 $X2=1.68
+ $Y2=0
r206 109 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=0
+ $X2=2.08 $Y2=0
r207 109 112 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=0
+ $X2=1.68 $Y2=0
r208 108 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.2 $Y2=0
r209 108 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r210 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r211 105 142 4.29038 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.49 $Y=0
+ $X2=0.245 $Y2=0
r212 105 107 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.49 $Y=0
+ $X2=0.72 $Y2=0
r213 104 145 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.09 $Y=0
+ $X2=1.225 $Y2=0
r214 104 107 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.72
+ $Y2=0
r215 102 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r216 102 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r217 102 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r218 100 134 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=7.97 $Y=0 $X2=7.92
+ $Y2=0
r219 100 101 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.97 $Y=0 $X2=8.1
+ $Y2=0
r220 98 131 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=6.96
+ $Y2=0
r221 98 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=7.24
+ $Y2=0
r222 97 134 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.37 $Y=0 $X2=7.92
+ $Y2=0
r223 97 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.37 $Y=0 $X2=7.24
+ $Y2=0
r224 95 128 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.25 $Y=0 $X2=6
+ $Y2=0
r225 95 96 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.25 $Y=0 $X2=6.38
+ $Y2=0
r226 94 131 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.51 $Y=0 $X2=6.96
+ $Y2=0
r227 94 96 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.51 $Y=0 $X2=6.38
+ $Y2=0
r228 92 119 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.6
+ $Y2=0
r229 92 93 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.8
+ $Y2=0
r230 90 116 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.64
+ $Y2=0
r231 90 91 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.952
+ $Y2=0
r232 89 119 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.095 $Y=0
+ $X2=3.6 $Y2=0
r233 89 91 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.095 $Y=0
+ $X2=2.952 $Y2=0
r234 85 160 3.03205 $w=2.95e-07 $l=1.06325e-07 $layer=LI1_cond $X=9.837 $Y=0.085
+ $X2=9.885 $Y2=0
r235 85 87 15.0404 $w=2.93e-07 $l=3.85e-07 $layer=LI1_cond $X=9.837 $Y=0.085
+ $X2=9.837 $Y2=0.47
r236 81 157 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0
r237 81 83 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0.47
r238 80 101 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.23 $Y=0 $X2=8.1
+ $Y2=0
r239 79 157 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.83 $Y=0 $X2=8.96
+ $Y2=0
r240 79 80 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.83 $Y=0 $X2=8.23
+ $Y2=0
r241 75 101 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.1 $Y=0.085
+ $X2=8.1 $Y2=0
r242 75 77 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=8.1 $Y=0.085
+ $X2=8.1 $Y2=0.47
r243 71 99 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0
r244 71 73 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0.47
r245 67 96 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.38 $Y=0.085
+ $X2=6.38 $Y2=0
r246 67 69 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=6.38 $Y=0.085
+ $X2=6.38 $Y2=0.47
r247 63 154 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.52 $Y2=0
r248 63 65 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.52 $Y2=0.47
r249 59 151 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.66 $Y2=0
r250 59 61 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.66 $Y2=0.47
r251 58 93 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.93 $Y=0 $X2=3.8
+ $Y2=0
r252 57 151 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.66
+ $Y2=0
r253 57 58 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=3.93
+ $Y2=0
r254 53 93 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=0.085
+ $X2=3.8 $Y2=0
r255 53 55 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=3.8 $Y=0.085
+ $X2=3.8 $Y2=0.47
r256 49 91 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.952 $Y=0.085
+ $X2=2.952 $Y2=0
r257 49 51 11.5244 $w=2.83e-07 $l=2.85e-07 $layer=LI1_cond $X=2.952 $Y=0.085
+ $X2=2.952 $Y2=0.37
r258 45 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0
r259 45 47 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0.56
r260 41 145 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0
r261 41 43 12.1647 $w=2.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0.37
r262 37 142 3.18714 $w=2.95e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.342 $Y=0.085
+ $X2=0.245 $Y2=0
r263 37 39 13.4777 $w=2.93e-07 $l=3.45e-07 $layer=LI1_cond $X=0.342 $Y=0.085
+ $X2=0.342 $Y2=0.43
r264 12 87 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=9.68
+ $Y=0.235 $X2=9.82 $Y2=0.47
r265 11 83 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=8.82
+ $Y=0.235 $X2=8.96 $Y2=0.47
r266 10 77 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=7.96
+ $Y=0.235 $X2=8.1 $Y2=0.47
r267 9 73 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=7.1
+ $Y=0.235 $X2=7.24 $Y2=0.47
r268 8 69 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=6.24
+ $Y=0.235 $X2=6.38 $Y2=0.47
r269 7 65 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.38
+ $Y=0.235 $X2=5.52 $Y2=0.47
r270 6 61 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.52
+ $Y=0.235 $X2=4.66 $Y2=0.47
r271 5 55 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=3.66
+ $Y=0.235 $X2=3.8 $Y2=0.47
r272 4 51 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=2.8
+ $Y=0.235 $X2=2.94 $Y2=0.37
r273 3 47 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.235 $X2=2.08 $Y2=0.56
r274 2 43 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.08
+ $Y=0.235 $X2=1.22 $Y2=0.37
r275 1 39 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=0.235
+ $Y=0.235 $X2=0.36 $Y2=0.43
.ends

