* File: sky130_fd_sc_lp__sdfstp_1.spice
* Created: Fri Aug 28 11:29:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfstp_1.pex.spice"
.subckt sky130_fd_sc_lp__sdfstp_1  VNB VPB SCD D SCE CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1014 A_124_128# N_SCD_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 N_A_196_128#_M1000_d N_SCE_M1000_g A_124_128# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 A_282_128# N_D_M1003_g N_A_196_128#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_A_324_102#_M1034_g A_282_128# VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0441 PD=0.74 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1038 N_A_324_102#_M1038_d N_SCE_M1038_g N_VGND_M1034_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=11.424 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_CLK_M1025_g N_A_702_47#_M1025_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1037 N_A_871_47#_M1037_d N_A_702_47#_M1037_g N_VGND_M1025_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_1135_57#_M1018_d N_A_702_47#_M1018_g N_A_196_128#_M1018_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.3135 PD=0.7 PS=2.35 NRD=0 NRS=101.424 M=1 R=2.8
+ SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1019 A_1221_57# N_A_871_47#_M1019_g N_A_1135_57#_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_1263_31#_M1022_g A_1221_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1039 A_1502_125# N_A_1135_57#_M1039_g N_A_1263_31#_M1039_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.1113 PD=0.78 PS=1.37 NRD=35.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.7 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_SET_B_M1021_g A_1502_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.199025 AS=0.0756 PD=1.35113 PS=0.78 NRD=151.428 NRS=35.712 M=1 R=2.8
+ SA=75000.7 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1007 A_1847_125# N_A_1135_57#_M1007_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.303275 PD=0.85 PS=2.05887 NRD=9.372 NRS=47.808 M=1 R=4.26667
+ SA=75001.3 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_1912_463#_M1002_d N_A_871_47#_M1002_g A_1847_125# VNB NSHORT L=0.15
+ W=0.64 AD=0.279487 AS=0.0672 PD=1.78113 PS=0.85 NRD=35.616 NRS=9.372 M=1
+ R=4.26667 SA=75001.7 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1006 A_2116_125# N_A_702_47#_M1006_g N_A_1912_463#_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.183413 PD=0.81 PS=1.16887 NRD=39.996 NRS=49.992 M=1
+ R=2.8 SA=75003.3 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1024 A_2224_125# N_A_2158_231#_M1024_g A_2116_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=39.996 M=1 R=2.8 SA=75003.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_SET_B_M1012_g A_2224_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=11.424 NRS=14.28 M=1 R=2.8 SA=75004.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1031 N_A_2158_231#_M1031_d N_A_1912_463#_M1031_g N_VGND_M1012_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75004.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1912_463#_M1005_g N_A_2598_153#_M1005_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0875 AS=0.1113 PD=0.8 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 N_Q_M1015_d N_A_2598_153#_M1015_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.175 PD=2.21 PS=1.6 NRD=0 NRS=4.284 M=1 R=5.6 SA=75000.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_SCD_M1013_g N_A_27_408#_M1013_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1033 A_196_408# N_SCE_M1033_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1036 N_A_196_128#_M1036_d N_D_M1036_g A_196_408# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=16.9223 NRS=15.3857 M=1 R=4.26667
+ SA=75001 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1009 N_A_27_408#_M1009_d N_A_324_102#_M1009_g N_A_196_128#_M1036_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1248 PD=1.81 PS=1.03 NRD=0 NRS=16.9223 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1026 N_A_324_102#_M1026_d N_SCE_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.39545 PD=1.81 PS=2.52 NRD=0 NRS=107.72 M=1 R=4.26667
+ SA=75000.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1027 N_VPWR_M1027_d N_CLK_M1027_g N_A_702_47#_M1027_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.3459 PD=0.92 PS=2.7 NRD=0 NRS=149.424 M=1 R=4.26667
+ SA=75000.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1016 N_A_871_47#_M1016_d N_A_702_47#_M1016_g N_VPWR_M1027_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1023 N_A_1135_57#_M1023_d N_A_871_47#_M1023_g N_A_196_128#_M1023_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1028 A_1221_463# N_A_702_47#_M1028_g N_A_1135_57#_M1023_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_1263_31#_M1032_g A_1221_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1281 AS=0.0441 PD=1.03 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_1263_31#_M1004_d N_A_1135_57#_M1004_g N_VPWR_M1032_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.06195 AS=0.1281 PD=0.715 PS=1.03 NRD=0 NRS=154.783 M=1
+ R=2.8 SA=75001.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_SET_B_M1020_g N_A_1263_31#_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1456 AS=0.06195 PD=1.02333 PS=0.715 NRD=143.042 NRS=7.0329 M=1
+ R=2.8 SA=75002.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1029 N_A_1703_379#_M1029_d N_A_1135_57#_M1029_g N_VPWR_M1020_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.2912 PD=2.21 PS=2.04667 NRD=0 NRS=26.3783 M=1
+ R=5.6 SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_1912_463#_M1001_d N_A_871_47#_M1001_g N_A_1810_463#_M1001_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0952 AS=0.1837 PD=0.823333 PS=1.82 NRD=80.5139
+ NRS=46.886 M=1 R=2.8 SA=75000.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_1703_379#_M1017_d N_A_702_47#_M1017_g N_A_1912_463#_M1001_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.221775 AS=0.1904 PD=2.21 PS=1.64667 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VPWR_M1010_d N_A_2158_231#_M1010_g N_A_1810_463#_M1010_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1035 N_A_1912_463#_M1035_d N_SET_B_M1035_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_2158_231#_M1011_d N_A_1912_463#_M1011_g N_VPWR_M1011_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_1912_463#_M1008_g N_A_2598_153#_M1008_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.14912 AS=0.1696 PD=1.14189 PS=1.81 NRD=24.625 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1030 N_Q_M1030_d N_A_2598_153#_M1030_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.29358 PD=3.05 PS=2.24811 NRD=0 NRS=8.077 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=27.5647 P=33.29
*
.include "sky130_fd_sc_lp__sdfstp_1.pxi.spice"
*
.ends
*
*
