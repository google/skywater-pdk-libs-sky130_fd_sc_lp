* NGSPICE file created from sky130_fd_sc_lp__nand4_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand4_lp A B C D VGND VNB VPB VPWR Y
M1000 VPWR C Y VPB phighvt w=1e+06u l=250000u
+  ad=9.25e+11p pd=7.85e+06u as=5.6e+11p ps=5.12e+06u
M1001 Y A a_324_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.764e+11p ps=1.68e+06u
M1002 a_132_47# D VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1003 a_324_47# B a_210_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
M1004 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y D VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_210_47# C a_132_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

