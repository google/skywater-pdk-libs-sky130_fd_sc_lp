* File: sky130_fd_sc_lp__invkapwr_4.pxi.spice
* Created: Fri Aug 28 10:39:16 2020
* 
x_PM_SKY130_FD_SC_LP__INVKAPWR_4%A N_A_M1001_g N_A_M1000_g N_A_M1002_g
+ N_A_M1004_g N_A_M1003_g N_A_M1007_g N_A_M1005_g N_A_M1008_g N_A_M1006_g
+ N_A_M1009_g A A A A A N_A_c_54_n N_A_c_55_n PM_SKY130_FD_SC_LP__INVKAPWR_4%A
x_PM_SKY130_FD_SC_LP__INVKAPWR_4%KAPWR N_KAPWR_M1001_d N_KAPWR_M1002_d
+ N_KAPWR_M1005_d N_KAPWR_M1009_d KAPWR N_KAPWR_c_153_p N_KAPWR_c_157_p
+ N_KAPWR_c_162_p N_KAPWR_c_167_p N_KAPWR_c_142_n KAPWR
+ PM_SKY130_FD_SC_LP__INVKAPWR_4%KAPWR
x_PM_SKY130_FD_SC_LP__INVKAPWR_4%Y N_Y_M1000_d N_Y_M1007_d N_Y_M1001_s
+ N_Y_M1003_s N_Y_M1006_s N_Y_c_187_n N_Y_c_188_n N_Y_c_189_n N_Y_c_199_n
+ N_Y_c_200_n N_Y_c_217_n N_Y_c_201_n N_Y_c_190_n N_Y_c_191_n N_Y_c_229_n
+ N_Y_c_202_n N_Y_c_192_n N_Y_c_237_n N_Y_c_203_n N_Y_c_193_n N_Y_c_204_n
+ N_Y_c_194_n N_Y_c_205_n Y Y Y N_Y_c_197_n N_Y_c_208_n Y
+ PM_SKY130_FD_SC_LP__INVKAPWR_4%Y
x_PM_SKY130_FD_SC_LP__INVKAPWR_4%VGND N_VGND_M1000_s N_VGND_M1004_s
+ N_VGND_M1008_s N_VGND_c_303_n N_VGND_c_304_n N_VGND_c_305_n VGND
+ N_VGND_c_306_n N_VGND_c_307_n N_VGND_c_308_n N_VGND_c_309_n N_VGND_c_310_n
+ N_VGND_c_311_n N_VGND_c_312_n PM_SKY130_FD_SC_LP__INVKAPWR_4%VGND
x_PM_SKY130_FD_SC_LP__INVKAPWR_4%VPWR VPWR N_VPWR_c_339_n VPWR
+ PM_SKY130_FD_SC_LP__INVKAPWR_4%VPWR
cc_1 VNB N_A_M1000_g 0.0452338f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=0.56
cc_2 VNB N_A_M1004_g 0.0357085f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=0.56
cc_3 VNB N_A_M1007_g 0.0357083f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=0.56
cc_4 VNB N_A_M1008_g 0.0452172f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=0.56
cc_5 VNB N_A_c_54_n 0.14785f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=1.46
cc_6 VNB N_A_c_55_n 0.0196611f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=1.46
cc_7 VNB N_Y_c_187_n 0.0302956f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.675
cc_8 VNB N_Y_c_188_n 0.0165372f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.465
cc_9 VNB N_Y_c_189_n 0.0128736f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.465
cc_10 VNB N_Y_c_190_n 0.00119645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_Y_c_191_n 0.00541162f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=2.465
cc_12 VNB N_Y_c_192_n 0.00119511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_Y_c_193_n 0.00212259f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.485
cc_14 VNB N_Y_c_194_n 0.00207568f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.46
cc_15 VNB Y 0.0159161f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.46
cc_16 VNB Y 0.0307643f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.46
cc_17 VNB N_Y_c_197_n 0.0132908f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=1.46
cc_18 VNB N_VGND_c_303_n 0.0235244f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=0.56
cc_19 VNB N_VGND_c_304_n 0.00697289f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.465
cc_20 VNB N_VGND_c_305_n 0.0235952f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=0.56
cc_21 VNB N_VGND_c_306_n 0.0171844f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=2.465
cc_22 VNB N_VGND_c_307_n 0.0170098f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=0.56
cc_23 VNB N_VGND_c_308_n 0.0217138f $X=-0.19 $Y=-0.245 $X2=2.795 $Y2=2.465
cc_24 VNB N_VGND_c_309_n 0.213186f $X=-0.19 $Y=-0.245 $X2=2.795 $Y2=2.465
cc_25 VNB N_VGND_c_310_n 0.0299338f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_26 VNB N_VGND_c_311_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.21
cc_27 VNB N_VGND_c_312_n 0.00577043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB VPWR 0.143779f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.675
cc_29 VPB N_A_M1001_g 0.0223406f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.465
cc_30 VPB N_A_M1002_g 0.0176925f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=2.465
cc_31 VPB N_A_M1003_g 0.0177107f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=2.465
cc_32 VPB N_A_M1005_g 0.0177107f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=2.465
cc_33 VPB N_A_M1006_g 0.0176925f $X=-0.19 $Y=1.655 $X2=2.365 $Y2=2.465
cc_34 VPB N_A_M1009_g 0.0223382f $X=-0.19 $Y=1.655 $X2=2.795 $Y2=2.465
cc_35 VPB N_A_c_54_n 0.0175902f $X=-0.19 $Y=1.655 $X2=2.7 $Y2=1.46
cc_36 VPB N_KAPWR_c_142_n 0.0379007f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_37 VPB N_Y_c_187_n 0.0029401f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=1.675
cc_38 VPB N_Y_c_199_n 0.00271023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_Y_c_200_n 0.0105735f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.295
cc_40 VPB N_Y_c_201_n 0.00244238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_Y_c_202_n 0.00239644f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_42 VPB N_Y_c_203_n 0.00204591f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.46
cc_43 VPB N_Y_c_204_n 0.00204591f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=1.485
cc_44 VPB N_Y_c_205_n 0.00209286f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.485
cc_45 VPB Y 0.00298715f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.46
cc_46 VPB Y 0.00199175f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.485
cc_47 VPB N_Y_c_208_n 0.0112565f $X=-0.19 $Y=1.655 $X2=2.795 $Y2=1.485
cc_48 VPB VPWR 0.0453892f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.675
cc_49 VPB N_VPWR_c_339_n 0.0948323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 N_A_M1001_g N_KAPWR_c_142_n 0.00731133f $X=0.645 $Y=2.465 $X2=0 $Y2=0
cc_51 N_A_M1002_g N_KAPWR_c_142_n 0.00731133f $X=1.075 $Y=2.465 $X2=0 $Y2=0
cc_52 N_A_M1003_g N_KAPWR_c_142_n 0.00731133f $X=1.505 $Y=2.465 $X2=0 $Y2=0
cc_53 N_A_M1005_g N_KAPWR_c_142_n 0.00731133f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_54 N_A_M1006_g N_KAPWR_c_142_n 0.00731133f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_55 N_A_M1009_g N_KAPWR_c_142_n 0.00731133f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_56 N_A_M1000_g N_Y_c_187_n 0.00398294f $X=1.075 $Y=0.56 $X2=0 $Y2=0
cc_57 N_A_c_54_n N_Y_c_187_n 0.00850442f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_58 N_A_c_55_n N_Y_c_187_n 0.0269937f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_59 N_A_M1000_g N_Y_c_188_n 0.0155371f $X=1.075 $Y=0.56 $X2=0 $Y2=0
cc_60 N_A_c_54_n N_Y_c_188_n 0.00243306f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_61 N_A_c_55_n N_Y_c_188_n 0.0461528f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_62 N_A_M1001_g N_Y_c_199_n 0.0159014f $X=0.645 $Y=2.465 $X2=0 $Y2=0
cc_63 N_A_c_55_n N_Y_c_199_n 0.0118161f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_64 N_A_M1001_g N_Y_c_217_n 8.21354e-19 $X=0.645 $Y=2.465 $X2=0 $Y2=0
cc_65 N_A_M1002_g N_Y_c_217_n 8.21794e-19 $X=1.075 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_M1002_g N_Y_c_201_n 0.0144277f $X=1.075 $Y=2.465 $X2=0 $Y2=0
cc_67 N_A_M1003_g N_Y_c_201_n 0.0144277f $X=1.505 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A_c_54_n N_Y_c_201_n 0.00269429f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_69 N_A_c_55_n N_Y_c_201_n 0.0443258f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_70 N_A_M1000_g N_Y_c_190_n 0.00194229f $X=1.075 $Y=0.56 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_Y_c_190_n 0.00105846f $X=1.505 $Y=0.56 $X2=0 $Y2=0
cc_72 N_A_M1004_g N_Y_c_191_n 0.0131322f $X=1.505 $Y=0.56 $X2=0 $Y2=0
cc_73 N_A_M1007_g N_Y_c_191_n 0.0131322f $X=1.935 $Y=0.56 $X2=0 $Y2=0
cc_74 N_A_c_54_n N_Y_c_191_n 5.70427e-19 $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_75 N_A_c_55_n N_Y_c_191_n 0.0457256f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_76 N_A_M1003_g N_Y_c_229_n 8.21354e-19 $X=1.505 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A_M1005_g N_Y_c_229_n 8.21794e-19 $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_M1005_g N_Y_c_202_n 0.0144277f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A_M1006_g N_Y_c_202_n 0.0144277f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A_c_54_n N_Y_c_202_n 0.00269429f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_81 N_A_c_55_n N_Y_c_202_n 0.0439495f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_82 N_A_M1007_g N_Y_c_192_n 0.00105549f $X=1.935 $Y=0.56 $X2=0 $Y2=0
cc_83 N_A_M1008_g N_Y_c_192_n 0.00192273f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_84 N_A_M1006_g N_Y_c_237_n 8.22659e-19 $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_M1009_g N_Y_c_237_n 8.22659e-19 $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A_c_54_n N_Y_c_203_n 0.0028086f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_87 N_A_c_55_n N_Y_c_203_n 0.0215289f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_88 N_A_c_54_n N_Y_c_193_n 6.30163e-19 $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_89 N_A_c_55_n N_Y_c_193_n 0.0229285f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_90 N_A_c_54_n N_Y_c_204_n 0.0028086f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_91 N_A_c_55_n N_Y_c_204_n 0.0215289f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_92 N_A_c_54_n N_Y_c_194_n 6.30163e-19 $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_93 N_A_c_55_n N_Y_c_194_n 0.0224875f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_94 N_A_c_54_n N_Y_c_205_n 0.0028086f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_95 N_A_c_55_n N_Y_c_205_n 0.0219511f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_96 N_A_M1008_g Y 0.0155371f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_97 N_A_c_54_n Y 0.00481111f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_98 N_A_c_55_n Y 0.0461529f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_99 N_A_M1008_g Y 0.00404256f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_100 N_A_c_54_n Y 0.0146731f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_101 N_A_c_55_n Y 0.0271544f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_102 N_A_M1009_g Y 0.0159821f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_c_54_n Y 0.00285842f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_104 N_A_c_55_n Y 0.0110823f $X=2.7 $Y=1.46 $X2=0 $Y2=0
cc_105 N_A_M1000_g N_VGND_c_303_n 0.0038152f $X=1.075 $Y=0.56 $X2=0 $Y2=0
cc_106 N_A_M1004_g N_VGND_c_304_n 0.00181038f $X=1.505 $Y=0.56 $X2=0 $Y2=0
cc_107 N_A_M1007_g N_VGND_c_304_n 0.00180279f $X=1.935 $Y=0.56 $X2=0 $Y2=0
cc_108 N_A_M1008_g N_VGND_c_305_n 0.00384067f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A_M1000_g N_VGND_c_306_n 0.00478016f $X=1.075 $Y=0.56 $X2=0 $Y2=0
cc_110 N_A_M1004_g N_VGND_c_306_n 0.00478016f $X=1.505 $Y=0.56 $X2=0 $Y2=0
cc_111 N_A_M1007_g N_VGND_c_307_n 0.00478016f $X=1.935 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A_M1008_g N_VGND_c_307_n 0.00478016f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_113 N_A_M1000_g N_VGND_c_309_n 0.0051579f $X=1.075 $Y=0.56 $X2=0 $Y2=0
cc_114 N_A_M1004_g N_VGND_c_309_n 0.00490796f $X=1.505 $Y=0.56 $X2=0 $Y2=0
cc_115 N_A_M1007_g N_VGND_c_309_n 0.00490796f $X=1.935 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A_M1008_g N_VGND_c_309_n 0.0051523f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_117 N_A_M1001_g VPWR 0.00638144f $X=0.645 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_118 N_A_M1002_g VPWR 0.0053229f $X=1.075 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_119 N_A_M1003_g VPWR 0.0053229f $X=1.505 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_120 N_A_M1005_g VPWR 0.0053229f $X=1.935 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_121 N_A_M1006_g VPWR 0.0053229f $X=2.365 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_122 N_A_M1009_g VPWR 0.00633019f $X=2.795 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_123 N_A_M1001_g N_VPWR_c_339_n 0.00585385f $X=0.645 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_M1002_g N_VPWR_c_339_n 0.00585385f $X=1.075 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_M1003_g N_VPWR_c_339_n 0.00585385f $X=1.505 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_M1005_g N_VPWR_c_339_n 0.00585385f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_M1006_g N_VPWR_c_339_n 0.00585385f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_M1009_g N_VPWR_c_339_n 0.00585385f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_129 N_KAPWR_c_142_n N_Y_M1001_s 9.4832e-19 $X=3.015 $Y=2.81 $X2=0 $Y2=0
cc_130 N_KAPWR_c_142_n N_Y_M1003_s 9.4832e-19 $X=3.015 $Y=2.81 $X2=0 $Y2=0
cc_131 N_KAPWR_c_142_n N_Y_M1006_s 7.22529e-19 $X=3.015 $Y=2.81 $X2=0 $Y2=0
cc_132 N_KAPWR_M1001_d N_Y_c_199_n 0.00119058f $X=0.3 $Y=1.835 $X2=0 $Y2=0
cc_133 N_KAPWR_c_153_p N_Y_c_199_n 0.00915704f $X=0.43 $Y=2.22 $X2=0 $Y2=0
cc_134 N_KAPWR_M1001_d N_Y_c_200_n 0.00134463f $X=0.3 $Y=1.835 $X2=0 $Y2=0
cc_135 N_KAPWR_c_153_p N_Y_c_200_n 0.00892602f $X=0.43 $Y=2.22 $X2=0 $Y2=0
cc_136 N_KAPWR_c_153_p N_Y_c_217_n 0.00885226f $X=0.43 $Y=2.22 $X2=0 $Y2=0
cc_137 N_KAPWR_c_157_p N_Y_c_217_n 0.0091127f $X=1.29 $Y=2.22 $X2=0 $Y2=0
cc_138 N_KAPWR_c_142_n N_Y_c_217_n 0.0284615f $X=3.015 $Y=2.81 $X2=0 $Y2=0
cc_139 N_KAPWR_M1002_d N_Y_c_201_n 0.00176461f $X=1.15 $Y=1.835 $X2=0 $Y2=0
cc_140 N_KAPWR_c_157_p N_Y_c_201_n 0.0135055f $X=1.29 $Y=2.22 $X2=0 $Y2=0
cc_141 N_KAPWR_c_157_p N_Y_c_229_n 0.00885226f $X=1.29 $Y=2.22 $X2=0 $Y2=0
cc_142 N_KAPWR_c_162_p N_Y_c_229_n 0.0091127f $X=2.15 $Y=2.22 $X2=0 $Y2=0
cc_143 N_KAPWR_c_142_n N_Y_c_229_n 0.0284615f $X=3.015 $Y=2.81 $X2=0 $Y2=0
cc_144 N_KAPWR_M1005_d N_Y_c_202_n 0.00176461f $X=2.01 $Y=1.835 $X2=0 $Y2=0
cc_145 N_KAPWR_c_162_p N_Y_c_202_n 0.0135055f $X=2.15 $Y=2.22 $X2=0 $Y2=0
cc_146 N_KAPWR_c_162_p N_Y_c_237_n 0.00911549f $X=2.15 $Y=2.22 $X2=0 $Y2=0
cc_147 N_KAPWR_c_167_p N_Y_c_237_n 0.0091127f $X=3.01 $Y=2.22 $X2=0 $Y2=0
cc_148 N_KAPWR_c_142_n N_Y_c_237_n 0.0288605f $X=3.015 $Y=2.81 $X2=0 $Y2=0
cc_149 N_KAPWR_M1009_d Y 0.00113743f $X=2.87 $Y=1.835 $X2=0 $Y2=0
cc_150 N_KAPWR_c_167_p Y 0.00875024f $X=3.01 $Y=2.22 $X2=0 $Y2=0
cc_151 N_KAPWR_M1009_d N_Y_c_208_n 0.0013308f $X=2.87 $Y=1.835 $X2=0 $Y2=0
cc_152 N_KAPWR_c_167_p N_Y_c_208_n 0.00892602f $X=3.01 $Y=2.22 $X2=0 $Y2=0
cc_153 N_KAPWR_M1001_d VPWR 0.00116402f $X=0.3 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_154 N_KAPWR_M1002_d VPWR 0.00121489f $X=1.15 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_155 N_KAPWR_M1005_d VPWR 0.00121489f $X=2.01 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_156 N_KAPWR_M1009_d VPWR 0.00114194f $X=2.87 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_157 N_KAPWR_c_153_p VPWR 0.00242444f $X=0.43 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_158 N_KAPWR_c_157_p VPWR 0.00242444f $X=1.29 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_159 N_KAPWR_c_162_p VPWR 0.00242444f $X=2.15 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_160 N_KAPWR_c_167_p VPWR 0.00237745f $X=3.01 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_161 N_KAPWR_c_142_n VPWR 0.335059f $X=3.015 $Y=2.81 $X2=-0.19 $Y2=1.655
cc_162 N_KAPWR_c_153_p N_VPWR_c_339_n 0.0165384f $X=0.43 $Y=2.22 $X2=0 $Y2=0
cc_163 N_KAPWR_c_157_p N_VPWR_c_339_n 0.0149362f $X=1.29 $Y=2.22 $X2=0 $Y2=0
cc_164 N_KAPWR_c_162_p N_VPWR_c_339_n 0.0149362f $X=2.15 $Y=2.22 $X2=0 $Y2=0
cc_165 N_KAPWR_c_167_p N_VPWR_c_339_n 0.0161868f $X=3.01 $Y=2.22 $X2=0 $Y2=0
cc_166 N_KAPWR_c_142_n N_VPWR_c_339_n 0.00847566f $X=3.015 $Y=2.81 $X2=0 $Y2=0
cc_167 N_Y_c_188_n N_VGND_c_303_n 0.0219547f $X=1.16 $Y=0.94 $X2=0 $Y2=0
cc_168 N_Y_c_191_n N_VGND_c_304_n 0.0169602f $X=2.02 $Y=0.94 $X2=0 $Y2=0
cc_169 Y N_VGND_c_305_n 0.022139f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_170 N_Y_c_190_n N_VGND_c_306_n 0.00786011f $X=1.29 $Y=0.56 $X2=0 $Y2=0
cc_171 N_Y_c_192_n N_VGND_c_307_n 0.0077623f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_172 N_Y_c_188_n N_VGND_c_309_n 0.0162091f $X=1.16 $Y=0.94 $X2=0 $Y2=0
cc_173 N_Y_c_189_n N_VGND_c_309_n 0.00670311f $X=0.4 $Y=0.94 $X2=0 $Y2=0
cc_174 N_Y_c_190_n N_VGND_c_309_n 0.00924776f $X=1.29 $Y=0.56 $X2=0 $Y2=0
cc_175 N_Y_c_191_n N_VGND_c_309_n 0.0106287f $X=2.02 $Y=0.94 $X2=0 $Y2=0
cc_176 N_Y_c_192_n N_VGND_c_309_n 0.00906853f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_177 Y N_VGND_c_309_n 0.0160501f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_178 N_Y_c_197_n N_VGND_c_309_n 0.00729456f $X=3.127 $Y=1.04 $X2=0 $Y2=0
cc_179 N_Y_M1001_s VPWR 0.00125588f $X=0.72 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_180 N_Y_M1003_s VPWR 0.00125588f $X=1.58 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_181 N_Y_M1006_s VPWR 0.0012358f $X=2.44 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_182 N_Y_c_217_n VPWR 0.0024325f $X=0.86 $Y=2 $X2=-0.19 $Y2=-0.245
cc_183 N_Y_c_229_n VPWR 0.0024325f $X=1.72 $Y=2 $X2=-0.19 $Y2=-0.245
cc_184 N_Y_c_237_n VPWR 0.00248057f $X=2.58 $Y=2 $X2=-0.19 $Y2=-0.245
cc_185 N_Y_c_217_n N_VPWR_c_339_n 0.0124051f $X=0.86 $Y=2 $X2=0 $Y2=0
cc_186 N_Y_c_229_n N_VPWR_c_339_n 0.0124051f $X=1.72 $Y=2 $X2=0 $Y2=0
cc_187 N_Y_c_237_n N_VPWR_c_339_n 0.012556f $X=2.58 $Y=2 $X2=0 $Y2=0
