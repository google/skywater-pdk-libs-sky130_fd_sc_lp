* File: sky130_fd_sc_lp__mux2i_0.spice
* Created: Wed Sep  2 10:00:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2i_0.pex.spice"
.subckt sky130_fd_sc_lp__mux2i_0  VNB VPB S A0 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_S_M1006_g N_A_47_48#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.1113 PD=0.84 PS=1.37 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1001 A_244_48# N_A_47_48#_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=17.136 M=1 R=2.8 SA=75000.8
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_A0_M1008_g A_244_48# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=21.42 NRS=18.564 M=1 R=2.8 SA=75001.1 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1005 A_436_48# N_A1_M1005_g N_Y_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.7
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_S_M1003_g A_436_48# VNB NSHORT L=0.15 W=0.42 AD=0.2205
+ AS=0.0504 PD=1.89 PS=0.66 NRD=74.28 NRS=18.564 M=1 R=2.8 SA=75002.1 SB=75000.4
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_S_M1002_g N_A_47_48#_M1002_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1536 AS=0.1696 PD=1.12 PS=1.81 NRD=29.2348 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1007 A_292_491# N_A_47_48#_M1007_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1536 PD=0.85 PS=1.12 NRD=15.3857 NRS=32.308 M=1 R=4.26667
+ SA=75000.8 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1009 N_Y_M1009_d N_A1_M1009_g A_292_491# VPB PHIGHVT L=0.15 W=0.64 AD=0.1136
+ AS=0.0672 PD=0.995 PS=0.85 NRD=13.8491 NRS=15.3857 M=1 R=4.26667 SA=75001.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 A_465_491# N_A0_M1000_g N_Y_M1009_d VPB PHIGHVT L=0.15 W=0.64 AD=0.088
+ AS=0.1136 PD=0.915 PS=0.995 NRD=25.3933 NRS=9.2196 M=1 R=4.26667 SA=75001.7
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1004_d N_S_M1004_g A_465_491# VPB PHIGHVT L=0.15 W=0.64 AD=0.1824
+ AS=0.088 PD=1.85 PS=0.915 NRD=0 NRS=25.3933 M=1 R=4.26667 SA=75002.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__mux2i_0.pxi.spice"
*
.ends
*
*
