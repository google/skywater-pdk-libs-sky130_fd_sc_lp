* File: sky130_fd_sc_lp__o2bb2a_1.pxi.spice
* Created: Fri Aug 28 11:11:41 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2A_1%A_80_21# N_A_80_21#_M1003_s N_A_80_21#_M1001_d
+ N_A_80_21#_M1005_g N_A_80_21#_M1011_g N_A_80_21#_c_82_n N_A_80_21#_c_83_n
+ N_A_80_21#_c_99_p N_A_80_21#_c_161_p N_A_80_21#_c_84_n N_A_80_21#_c_85_n
+ N_A_80_21#_c_86_n N_A_80_21#_c_87_n N_A_80_21#_c_88_n N_A_80_21#_c_89_n
+ N_A_80_21#_c_90_n N_A_80_21#_c_91_n N_A_80_21#_c_95_n N_A_80_21#_c_92_n
+ PM_SKY130_FD_SC_LP__O2BB2A_1%A_80_21#
x_PM_SKY130_FD_SC_LP__O2BB2A_1%A1_N N_A1_N_M1010_g N_A1_N_c_186_n N_A1_N_M1009_g
+ N_A1_N_c_188_n A1_N A1_N A1_N N_A1_N_c_185_n PM_SKY130_FD_SC_LP__O2BB2A_1%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2A_1%A2_N N_A2_N_c_228_n N_A2_N_M1007_g N_A2_N_M1004_g
+ N_A2_N_c_229_n A2_N N_A2_N_c_232_n N_A2_N_c_233_n N_A2_N_c_230_n
+ PM_SKY130_FD_SC_LP__O2BB2A_1%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2A_1%A_286_492# N_A_286_492#_M1007_d
+ N_A_286_492#_M1009_d N_A_286_492#_M1003_g N_A_286_492#_M1001_g
+ N_A_286_492#_c_279_n N_A_286_492#_c_287_n N_A_286_492#_c_346_p
+ N_A_286_492#_c_280_n N_A_286_492#_c_288_n N_A_286_492#_c_289_n
+ N_A_286_492#_c_281_n N_A_286_492#_c_282_n N_A_286_492#_c_283_n
+ N_A_286_492#_c_290_n N_A_286_492#_c_284_n
+ PM_SKY130_FD_SC_LP__O2BB2A_1%A_286_492#
x_PM_SKY130_FD_SC_LP__O2BB2A_1%B2 N_B2_M1006_g N_B2_M1008_g B2 B2 N_B2_c_359_n
+ PM_SKY130_FD_SC_LP__O2BB2A_1%B2
x_PM_SKY130_FD_SC_LP__O2BB2A_1%B1 N_B1_M1002_g N_B1_M1000_g N_B1_c_398_n
+ N_B1_c_399_n B1 B1 N_B1_c_403_n PM_SKY130_FD_SC_LP__O2BB2A_1%B1
x_PM_SKY130_FD_SC_LP__O2BB2A_1%X N_X_M1005_s N_X_M1011_s X X X X X X X
+ N_X_c_433_n PM_SKY130_FD_SC_LP__O2BB2A_1%X
x_PM_SKY130_FD_SC_LP__O2BB2A_1%VPWR N_VPWR_M1011_d N_VPWR_M1004_d N_VPWR_M1002_d
+ N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n VPWR
+ N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n
+ N_VPWR_c_444_n PM_SKY130_FD_SC_LP__O2BB2A_1%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2A_1%VGND N_VGND_M1005_d N_VGND_M1006_d N_VGND_c_498_n
+ N_VGND_c_499_n VGND N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n
+ N_VGND_c_503_n N_VGND_c_504_n N_VGND_c_505_n PM_SKY130_FD_SC_LP__O2BB2A_1%VGND
x_PM_SKY130_FD_SC_LP__O2BB2A_1%A_506_47# N_A_506_47#_M1003_d N_A_506_47#_M1000_d
+ N_A_506_47#_c_552_n N_A_506_47#_c_553_n N_A_506_47#_c_554_n
+ N_A_506_47#_c_555_n PM_SKY130_FD_SC_LP__O2BB2A_1%A_506_47#
cc_1 VNB N_A_80_21#_M1011_g 0.00875585f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB N_A_80_21#_c_82_n 0.00722204f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.35
cc_3 VNB N_A_80_21#_c_83_n 0.0394033f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.35
cc_4 VNB N_A_80_21#_c_84_n 0.0012164f $X=-0.19 $Y=-0.245 $X2=1.182 $Y2=0.86
cc_5 VNB N_A_80_21#_c_85_n 0.00454234f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=0.405
cc_6 VNB N_A_80_21#_c_86_n 0.00845934f $X=-0.19 $Y=-0.245 $X2=2.272 $Y2=1.055
cc_7 VNB N_A_80_21#_c_87_n 0.0069911f $X=-0.19 $Y=-0.245 $X2=2.67 $Y2=1.14
cc_8 VNB N_A_80_21#_c_88_n 0.00311314f $X=-0.19 $Y=-0.245 $X2=2.37 $Y2=1.14
cc_9 VNB N_A_80_21#_c_89_n 0.0031467f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.65
cc_10 VNB N_A_80_21#_c_90_n 0.0227929f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=0.45
cc_11 VNB N_A_80_21#_c_91_n 0.00351901f $X=-0.19 $Y=-0.245 $X2=2.272 $Y2=0.45
cc_12 VNB N_A_80_21#_c_92_n 0.0212839f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.185
cc_13 VNB N_A1_N_M1010_g 0.0376915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A1_N 0.00601693f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_15 VNB N_A1_N_c_185_n 0.015113f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.945
cc_16 VNB N_A2_N_c_228_n 0.0188298f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=0.235
cc_17 VNB N_A2_N_c_229_n 0.029373f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_18 VNB N_A2_N_c_230_n 0.017667f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.945
cc_19 VNB N_A_286_492#_M1003_g 0.0564667f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_20 VNB N_A_286_492#_c_279_n 0.00640394f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.35
cc_21 VNB N_A_286_492#_c_280_n 0.00831965f $X=-0.19 $Y=-0.245 $X2=2.272 $Y2=0.62
cc_22 VNB N_A_286_492#_c_281_n 0.0200579f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.225
cc_23 VNB N_A_286_492#_c_282_n 0.00270788f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.65
cc_24 VNB N_A_286_492#_c_283_n 0.00133818f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=0.45
cc_25 VNB N_A_286_492#_c_284_n 0.0167239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B2_M1006_g 0.0446114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B2_M1008_g 0.00129756f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_28 VNB B2 0.0304427f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_29 VNB N_B2_c_359_n 0.0410975f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.945
cc_30 VNB N_B1_M1000_g 0.0282968f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_31 VNB N_B1_c_398_n 0.0353597f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.515
cc_32 VNB N_B1_c_399_n 0.0298495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_433_n 0.0613903f $X=-0.19 $Y=-0.245 $X2=1.182 $Y2=0.86
cc_34 VNB N_VPWR_c_444_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_498_n 0.00824462f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_36 VNB N_VGND_c_499_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_500_n 0.0153759f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.35
cc_38 VNB N_VGND_c_501_n 0.0499357f $X=-0.19 $Y=-0.245 $X2=1.182 $Y2=0.86
cc_39 VNB N_VGND_c_502_n 0.0164297f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=0.445
cc_40 VNB N_VGND_c_503_n 0.222179f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=0.45
cc_41 VNB N_VGND_c_504_n 0.00551901f $X=-0.19 $Y=-0.245 $X2=2.67 $Y2=2.785
cc_42 VNB N_VGND_c_505_n 0.00436611f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.785
cc_43 VNB N_A_506_47#_c_552_n 0.00102632f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_44 VNB N_A_506_47#_c_553_n 0.0161118f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_45 VNB N_A_506_47#_c_554_n 0.00356759f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_46 VNB N_A_506_47#_c_555_n 0.0173143f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.35
cc_47 VPB N_A_80_21#_M1011_g 0.0262875f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_48 VPB N_A_80_21#_c_89_n 0.00473965f $X=-0.19 $Y=1.655 $X2=2.755 $Y2=2.65
cc_49 VPB N_A_80_21#_c_95_n 0.00261407f $X=-0.19 $Y=1.655 $X2=2.755 $Y2=2.785
cc_50 VPB N_A1_N_c_186_n 0.023531f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A1_N_M1009_g 0.0245765f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_52 VPB N_A1_N_c_188_n 0.0242054f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_53 VPB N_A1_N_c_185_n 0.0101482f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=0.945
cc_54 VPB N_A2_N_M1004_g 0.0261696f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_55 VPB N_A2_N_c_232_n 0.0300759f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.35
cc_56 VPB N_A2_N_c_233_n 0.00869846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A2_N_c_230_n 0.0109499f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=0.945
cc_58 VPB N_A_286_492#_M1001_g 0.0325619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_286_492#_c_279_n 0.0193406f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.35
cc_60 VPB N_A_286_492#_c_287_n 0.0170044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_286_492#_c_288_n 0.010072f $X=-0.19 $Y=1.655 $X2=2.67 $Y2=1.14
cc_62 VPB N_A_286_492#_c_289_n 0.00738484f $X=-0.19 $Y=1.655 $X2=2.37 $Y2=1.14
cc_63 VPB N_A_286_492#_c_290_n 0.00241673f $X=-0.19 $Y=1.655 $X2=2.24 $Y2=0.445
cc_64 VPB N_B2_M1008_g 0.0514133f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_65 VPB B2 0.0118767f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_66 VPB N_B1_M1002_g 0.0328021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_B1_c_398_n 0.0153409f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.515
cc_68 VPB B1 0.0254372f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.35
cc_69 VPB N_B1_c_403_n 0.0468665f $X=-0.19 $Y=1.655 $X2=1.32 $Y2=0.405
cc_70 VPB N_X_c_433_n 0.0567722f $X=-0.19 $Y=1.655 $X2=1.182 $Y2=0.86
cc_71 VPB N_VPWR_c_445_n 0.00916844f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_72 VPB N_VPWR_c_446_n 0.0165531f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.35
cc_73 VPB N_VPWR_c_447_n 0.0144238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_448_n 0.0312418f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.945
cc_75 VPB N_VPWR_c_449_n 0.0153973f $X=-0.19 $Y=1.655 $X2=1.32 $Y2=0.405
cc_76 VPB N_VPWR_c_450_n 0.0210047f $X=-0.19 $Y=1.655 $X2=2.755 $Y2=1.225
cc_77 VPB N_VPWR_c_451_n 0.0302263f $X=-0.19 $Y=1.655 $X2=2.272 $Y2=0.45
cc_78 VPB N_VPWR_c_452_n 0.0263103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_453_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_444_n 0.0777466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 N_A_80_21#_M1011_g N_A1_N_M1010_g 0.0114127f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_82_n N_A1_N_M1010_g 0.00621493f $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_83_n N_A1_N_M1010_g 0.0164699f $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_99_p N_A1_N_M1010_g 0.00871408f $X=1.045 $Y=0.945 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_84_n N_A1_N_M1010_g 0.00982005f $X=1.182 $Y=0.86 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_85_n N_A1_N_M1010_g 0.00283114f $X=1.32 $Y=0.405 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_92_n N_A1_N_M1010_g 0.0104328f $X=0.597 $Y=1.185 $X2=0 $Y2=0
cc_88 N_A_80_21#_M1011_g A1_N 0.00171143f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_82_n A1_N 0.0242731f $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_83_n A1_N 3.3658e-19 $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_99_p A1_N 0.021333f $X=1.045 $Y=0.945 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_99_p N_A1_N_c_185_n 4.04168e-19 $X=1.045 $Y=0.945 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_99_p N_A2_N_c_228_n 0.00134292f $X=1.045 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_80_21#_c_84_n N_A2_N_c_228_n 0.00519058f $X=1.182 $Y=0.86 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A_80_21#_c_86_n N_A2_N_c_228_n 0.00145694f $X=2.272 $Y=1.055 $X2=-0.19
+ $Y2=-0.245
cc_96 N_A_80_21#_c_88_n N_A2_N_c_228_n 5.43209e-19 $X=2.37 $Y=1.14 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_80_21#_c_90_n N_A2_N_c_228_n 0.00909667f $X=2.075 $Y=0.45 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_80_21#_c_91_n N_A2_N_c_228_n 0.00230776f $X=2.272 $Y=0.45 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_80_21#_c_90_n N_A2_N_c_229_n 6.76832e-19 $X=2.075 $Y=0.45 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_86_n N_A_286_492#_M1003_g 0.0126783f $X=2.272 $Y=1.055 $X2=0
+ $Y2=0
cc_101 N_A_80_21#_c_87_n N_A_286_492#_M1003_g 0.0168498f $X=2.67 $Y=1.14 $X2=0
+ $Y2=0
cc_102 N_A_80_21#_c_89_n N_A_286_492#_M1003_g 0.00384049f $X=2.755 $Y=2.65 $X2=0
+ $Y2=0
cc_103 N_A_80_21#_c_89_n N_A_286_492#_M1001_g 0.00570141f $X=2.755 $Y=2.65 $X2=0
+ $Y2=0
cc_104 N_A_80_21#_c_95_n N_A_286_492#_M1001_g 0.00487246f $X=2.755 $Y=2.785
+ $X2=0 $Y2=0
cc_105 N_A_80_21#_c_99_p N_A_286_492#_c_280_n 0.0111224f $X=1.045 $Y=0.945 $X2=0
+ $Y2=0
cc_106 N_A_80_21#_c_84_n N_A_286_492#_c_280_n 0.00967826f $X=1.182 $Y=0.86 $X2=0
+ $Y2=0
cc_107 N_A_80_21#_c_86_n N_A_286_492#_c_280_n 0.0193687f $X=2.272 $Y=1.055 $X2=0
+ $Y2=0
cc_108 N_A_80_21#_c_88_n N_A_286_492#_c_280_n 0.0102225f $X=2.37 $Y=1.14 $X2=0
+ $Y2=0
cc_109 N_A_80_21#_c_90_n N_A_286_492#_c_280_n 0.0241812f $X=2.075 $Y=0.45 $X2=0
+ $Y2=0
cc_110 N_A_80_21#_c_89_n N_A_286_492#_c_288_n 0.0135589f $X=2.755 $Y=2.65 $X2=0
+ $Y2=0
cc_111 N_A_80_21#_c_88_n N_A_286_492#_c_281_n 0.00518559f $X=2.37 $Y=1.14 $X2=0
+ $Y2=0
cc_112 N_A_80_21#_c_87_n N_A_286_492#_c_283_n 0.00945797f $X=2.67 $Y=1.14 $X2=0
+ $Y2=0
cc_113 N_A_80_21#_c_88_n N_A_286_492#_c_283_n 0.0109962f $X=2.37 $Y=1.14 $X2=0
+ $Y2=0
cc_114 N_A_80_21#_c_89_n N_A_286_492#_c_283_n 0.0135424f $X=2.755 $Y=2.65 $X2=0
+ $Y2=0
cc_115 N_A_80_21#_c_89_n N_A_286_492#_c_290_n 0.054102f $X=2.755 $Y=2.65 $X2=0
+ $Y2=0
cc_116 N_A_80_21#_c_87_n N_A_286_492#_c_284_n 0.00169339f $X=2.67 $Y=1.14 $X2=0
+ $Y2=0
cc_117 N_A_80_21#_c_88_n N_A_286_492#_c_284_n 9.94742e-19 $X=2.37 $Y=1.14 $X2=0
+ $Y2=0
cc_118 N_A_80_21#_c_89_n N_A_286_492#_c_284_n 0.00436594f $X=2.755 $Y=2.65 $X2=0
+ $Y2=0
cc_119 N_A_80_21#_c_87_n N_B2_M1006_g 0.00618999f $X=2.67 $Y=1.14 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_89_n N_B2_M1006_g 0.00131429f $X=2.755 $Y=2.65 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_89_n N_B2_M1008_g 0.0235135f $X=2.755 $Y=2.65 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_95_n N_B2_M1008_g 0.00537437f $X=2.755 $Y=2.785 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_87_n B2 0.0101458f $X=2.67 $Y=1.14 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_89_n B2 0.0406859f $X=2.755 $Y=2.65 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_89_n N_B2_c_359_n 0.00743212f $X=2.755 $Y=2.65 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_89_n N_B1_M1002_g 0.00192326f $X=2.755 $Y=2.65 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_95_n N_B1_M1002_g 7.65712e-19 $X=2.755 $Y=2.785 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_89_n N_B1_c_398_n 3.67934e-19 $X=2.755 $Y=2.65 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_89_n B1 0.0208817f $X=2.755 $Y=2.65 $X2=0 $Y2=0
cc_130 N_A_80_21#_c_89_n N_B1_c_403_n 5.18873e-19 $X=2.755 $Y=2.65 $X2=0 $Y2=0
cc_131 N_A_80_21#_c_82_n N_X_c_433_n 0.0358235f $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_92_n N_X_c_433_n 0.0294981f $X=0.597 $Y=1.185 $X2=0 $Y2=0
cc_133 N_A_80_21#_M1011_g N_VPWR_c_445_n 0.00902817f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_80_21#_c_82_n N_VPWR_c_445_n 0.0192117f $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_83_n N_VPWR_c_445_n 0.00180833f $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_95_n N_VPWR_c_446_n 0.0181691f $X=2.755 $Y=2.785 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_89_n N_VPWR_c_448_n 0.00425845f $X=2.755 $Y=2.65 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_95_n N_VPWR_c_448_n 0.00859568f $X=2.755 $Y=2.785 $X2=0
+ $Y2=0
cc_139 N_A_80_21#_M1011_g N_VPWR_c_449_n 0.00487821f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_80_21#_c_95_n N_VPWR_c_451_n 0.0110955f $X=2.755 $Y=2.785 $X2=0 $Y2=0
cc_141 N_A_80_21#_M1011_g N_VPWR_c_452_n 0.0160671f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_80_21#_M1011_g N_VPWR_c_444_n 0.00917991f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_80_21#_c_95_n N_VPWR_c_444_n 0.0114686f $X=2.755 $Y=2.785 $X2=0 $Y2=0
cc_144 N_A_80_21#_c_82_n N_VGND_M1005_d 5.54893e-19 $X=0.63 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_80_21#_c_99_p N_VGND_M1005_d 0.00648372f $X=1.045 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_80_21#_c_161_p N_VGND_M1005_d 0.00380942f $X=0.865 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_80_21#_c_83_n N_VGND_c_498_n 8.76527e-19 $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_148 N_A_80_21#_c_99_p N_VGND_c_498_n 6.82543e-19 $X=1.045 $Y=0.945 $X2=0
+ $Y2=0
cc_149 N_A_80_21#_c_161_p N_VGND_c_498_n 0.02462f $X=0.865 $Y=0.945 $X2=0 $Y2=0
cc_150 N_A_80_21#_c_84_n N_VGND_c_498_n 0.0124662f $X=1.182 $Y=0.86 $X2=0 $Y2=0
cc_151 N_A_80_21#_c_85_n N_VGND_c_498_n 0.0221859f $X=1.32 $Y=0.405 $X2=0 $Y2=0
cc_152 N_A_80_21#_c_92_n N_VGND_c_498_n 0.0141937f $X=0.597 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A_80_21#_c_92_n N_VGND_c_500_n 0.00486043f $X=0.597 $Y=1.185 $X2=0
+ $Y2=0
cc_154 N_A_80_21#_c_85_n N_VGND_c_501_n 0.0170186f $X=1.32 $Y=0.405 $X2=0 $Y2=0
cc_155 N_A_80_21#_c_90_n N_VGND_c_501_n 0.0588572f $X=2.075 $Y=0.45 $X2=0 $Y2=0
cc_156 N_A_80_21#_M1003_s N_VGND_c_503_n 0.00250893f $X=2.115 $Y=0.235 $X2=0
+ $Y2=0
cc_157 N_A_80_21#_c_99_p N_VGND_c_503_n 0.00578827f $X=1.045 $Y=0.945 $X2=0
+ $Y2=0
cc_158 N_A_80_21#_c_161_p N_VGND_c_503_n 0.00118545f $X=0.865 $Y=0.945 $X2=0
+ $Y2=0
cc_159 N_A_80_21#_c_85_n N_VGND_c_503_n 0.0105615f $X=1.32 $Y=0.405 $X2=0 $Y2=0
cc_160 N_A_80_21#_c_90_n N_VGND_c_503_n 0.0393163f $X=2.075 $Y=0.45 $X2=0 $Y2=0
cc_161 N_A_80_21#_c_92_n N_VGND_c_503_n 0.00917987f $X=0.597 $Y=1.185 $X2=0
+ $Y2=0
cc_162 N_A_80_21#_c_99_p A_237_131# 0.00242326f $X=1.045 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_80_21#_c_84_n A_237_131# 0.00202533f $X=1.182 $Y=0.86 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_80_21#_c_86_n N_A_506_47#_c_552_n 0.00454354f $X=2.272 $Y=1.055 $X2=0
+ $Y2=0
cc_165 N_A_80_21#_c_87_n N_A_506_47#_c_553_n 0.00604817f $X=2.67 $Y=1.14 $X2=0
+ $Y2=0
cc_166 N_A_80_21#_c_86_n N_A_506_47#_c_554_n 0.0144831f $X=2.272 $Y=1.055 $X2=0
+ $Y2=0
cc_167 N_A_80_21#_c_87_n N_A_506_47#_c_554_n 0.0196618f $X=2.67 $Y=1.14 $X2=0
+ $Y2=0
cc_168 N_A1_N_M1010_g N_A2_N_c_228_n 0.0405345f $X=1.11 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A1_N_c_188_n N_A2_N_M1004_g 0.0184021f $X=1.232 $Y=2.245 $X2=0 $Y2=0
cc_170 A1_N N_A2_N_c_229_n 0.00100168f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A1_N_c_185_n N_A2_N_c_229_n 3.7023e-19 $X=1.2 $Y=1.74 $X2=0 $Y2=0
cc_172 N_A1_N_c_186_n N_A2_N_c_232_n 0.0172256f $X=1.232 $Y=2.048 $X2=0 $Y2=0
cc_173 A1_N N_A2_N_c_233_n 0.0312452f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A1_N_c_185_n N_A2_N_c_233_n 0.00268871f $X=1.2 $Y=1.74 $X2=0 $Y2=0
cc_175 N_A1_N_M1010_g N_A2_N_c_230_n 0.00484323f $X=1.11 $Y=0.865 $X2=0 $Y2=0
cc_176 A1_N N_A2_N_c_230_n 0.0021412f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A1_N_c_185_n N_A2_N_c_230_n 0.0172256f $X=1.2 $Y=1.74 $X2=0 $Y2=0
cc_178 N_A1_N_M1010_g N_A_286_492#_c_280_n 0.00144759f $X=1.11 $Y=0.865 $X2=0
+ $Y2=0
cc_179 A1_N N_A_286_492#_c_280_n 0.0157322f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A1_N_M1009_g N_A_286_492#_c_289_n 0.00255261f $X=1.355 $Y=2.67 $X2=0
+ $Y2=0
cc_181 N_A1_N_M1010_g N_A_286_492#_c_282_n 4.96815e-19 $X=1.11 $Y=0.865 $X2=0
+ $Y2=0
cc_182 A1_N N_A_286_492#_c_282_n 0.0150846f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A1_N_c_186_n N_VPWR_c_445_n 0.00533645f $X=1.232 $Y=2.048 $X2=0 $Y2=0
cc_184 N_A1_N_M1009_g N_VPWR_c_445_n 0.00488921f $X=1.355 $Y=2.67 $X2=0 $Y2=0
cc_185 A1_N N_VPWR_c_445_n 0.0265844f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A1_N_M1009_g N_VPWR_c_450_n 0.00520566f $X=1.355 $Y=2.67 $X2=0 $Y2=0
cc_187 N_A1_N_M1009_g N_VPWR_c_452_n 0.00659649f $X=1.355 $Y=2.67 $X2=0 $Y2=0
cc_188 N_A1_N_c_188_n N_VPWR_c_452_n 0.00591997f $X=1.232 $Y=2.245 $X2=0 $Y2=0
cc_189 A1_N N_VPWR_c_452_n 0.0105515f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A1_N_M1009_g N_VPWR_c_444_n 0.00520574f $X=1.355 $Y=2.67 $X2=0 $Y2=0
cc_191 N_A1_N_M1010_g N_VGND_c_498_n 0.00133695f $X=1.11 $Y=0.865 $X2=0 $Y2=0
cc_192 N_A1_N_M1010_g N_VGND_c_501_n 7.51565e-19 $X=1.11 $Y=0.865 $X2=0 $Y2=0
cc_193 N_A1_N_M1010_g N_VGND_c_503_n 3.0748e-19 $X=1.11 $Y=0.865 $X2=0 $Y2=0
cc_194 N_A2_N_c_229_n N_A_286_492#_M1003_g 0.00345042f $X=1.745 $Y=1.26 $X2=0
+ $Y2=0
cc_195 N_A2_N_M1004_g N_A_286_492#_M1001_g 0.0147421f $X=1.785 $Y=2.67 $X2=0
+ $Y2=0
cc_196 N_A2_N_c_232_n N_A_286_492#_M1001_g 0.00363775f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_197 N_A2_N_c_232_n N_A_286_492#_c_279_n 0.0109159f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_198 N_A2_N_c_233_n N_A_286_492#_c_279_n 0.00169553f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_199 N_A2_N_c_228_n N_A_286_492#_c_280_n 0.00932704f $X=1.5 $Y=1.185 $X2=0
+ $Y2=0
cc_200 N_A2_N_c_229_n N_A_286_492#_c_280_n 0.0144158f $X=1.745 $Y=1.26 $X2=0
+ $Y2=0
cc_201 N_A2_N_c_230_n N_A_286_492#_c_280_n 0.00234991f $X=1.835 $Y=1.87 $X2=0
+ $Y2=0
cc_202 N_A2_N_M1004_g N_A_286_492#_c_288_n 0.0124766f $X=1.785 $Y=2.67 $X2=0
+ $Y2=0
cc_203 N_A2_N_c_232_n N_A_286_492#_c_288_n 0.00435618f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_204 N_A2_N_c_233_n N_A_286_492#_c_288_n 0.0241167f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_205 N_A2_N_c_233_n N_A_286_492#_c_289_n 0.0109391f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_206 N_A2_N_c_232_n N_A_286_492#_c_281_n 6.28147e-19 $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_207 N_A2_N_c_233_n N_A_286_492#_c_281_n 0.00921479f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_208 N_A2_N_c_232_n N_A_286_492#_c_282_n 3.55225e-19 $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_209 N_A2_N_c_233_n N_A_286_492#_c_282_n 0.0270233f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_210 N_A2_N_c_230_n N_A_286_492#_c_282_n 0.00912405f $X=1.835 $Y=1.87 $X2=0
+ $Y2=0
cc_211 N_A2_N_M1004_g N_A_286_492#_c_290_n 0.0020923f $X=1.785 $Y=2.67 $X2=0
+ $Y2=0
cc_212 N_A2_N_c_232_n N_A_286_492#_c_290_n 0.00186964f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_213 N_A2_N_c_233_n N_A_286_492#_c_290_n 0.0227771f $X=1.835 $Y=2.035 $X2=0
+ $Y2=0
cc_214 N_A2_N_c_230_n N_A_286_492#_c_290_n 0.00113885f $X=1.835 $Y=1.87 $X2=0
+ $Y2=0
cc_215 N_A2_N_c_230_n N_A_286_492#_c_284_n 0.0128293f $X=1.835 $Y=1.87 $X2=0
+ $Y2=0
cc_216 N_A2_N_M1004_g N_VPWR_c_446_n 0.00693691f $X=1.785 $Y=2.67 $X2=0 $Y2=0
cc_217 N_A2_N_M1004_g N_VPWR_c_450_n 0.00520566f $X=1.785 $Y=2.67 $X2=0 $Y2=0
cc_218 N_A2_N_M1004_g N_VPWR_c_444_n 0.00520574f $X=1.785 $Y=2.67 $X2=0 $Y2=0
cc_219 N_A2_N_c_228_n N_VGND_c_501_n 5.20335e-19 $X=1.5 $Y=1.185 $X2=0 $Y2=0
cc_220 N_A_286_492#_M1003_g N_B2_M1006_g 0.0393908f $X=2.455 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_286_492#_M1001_g N_B2_M1008_g 0.0255596f $X=2.455 $Y=2.67 $X2=0 $Y2=0
cc_222 N_A_286_492#_c_279_n N_B2_M1008_g 0.0173972f $X=2.405 $Y=1.91 $X2=0 $Y2=0
cc_223 N_A_286_492#_c_290_n N_B2_c_359_n 6.70921e-19 $X=2.37 $Y=2.31 $X2=0 $Y2=0
cc_224 N_A_286_492#_c_284_n N_B2_c_359_n 0.0173972f $X=2.405 $Y=1.57 $X2=0 $Y2=0
cc_225 N_A_286_492#_c_288_n N_VPWR_M1004_d 0.00529481f $X=2.24 $Y=2.395 $X2=0
+ $Y2=0
cc_226 N_A_286_492#_c_289_n N_VPWR_c_445_n 0.00580027f $X=1.675 $Y=2.395 $X2=0
+ $Y2=0
cc_227 N_A_286_492#_M1001_g N_VPWR_c_446_n 0.00544558f $X=2.455 $Y=2.67 $X2=0
+ $Y2=0
cc_228 N_A_286_492#_c_288_n N_VPWR_c_446_n 0.0265854f $X=2.24 $Y=2.395 $X2=0
+ $Y2=0
cc_229 N_A_286_492#_c_346_p N_VPWR_c_450_n 0.00543687f $X=1.57 $Y=2.67 $X2=0
+ $Y2=0
cc_230 N_A_286_492#_M1001_g N_VPWR_c_451_n 0.0049668f $X=2.455 $Y=2.67 $X2=0
+ $Y2=0
cc_231 N_A_286_492#_M1001_g N_VPWR_c_444_n 0.00520574f $X=2.455 $Y=2.67 $X2=0
+ $Y2=0
cc_232 N_A_286_492#_c_346_p N_VPWR_c_444_n 0.00790036f $X=1.57 $Y=2.67 $X2=0
+ $Y2=0
cc_233 N_A_286_492#_c_288_n N_VPWR_c_444_n 0.0180233f $X=2.24 $Y=2.395 $X2=0
+ $Y2=0
cc_234 N_A_286_492#_M1003_g N_VGND_c_499_n 0.00126049f $X=2.455 $Y=0.445 $X2=0
+ $Y2=0
cc_235 N_A_286_492#_M1003_g N_VGND_c_501_n 0.00585385f $X=2.455 $Y=0.445 $X2=0
+ $Y2=0
cc_236 N_A_286_492#_M1003_g N_VGND_c_503_n 0.0124078f $X=2.455 $Y=0.445 $X2=0
+ $Y2=0
cc_237 N_A_286_492#_M1003_g N_A_506_47#_c_552_n 5.36223e-19 $X=2.455 $Y=0.445
+ $X2=0 $Y2=0
cc_238 N_A_286_492#_M1003_g N_A_506_47#_c_554_n 0.00151072f $X=2.455 $Y=0.445
+ $X2=0 $Y2=0
cc_239 N_B2_M1006_g N_B1_M1000_g 0.0267985f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_240 N_B2_M1006_g N_B1_c_398_n 0.00212047f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_241 N_B2_M1008_g N_B1_c_398_n 0.00238731f $X=2.885 $Y=2.67 $X2=0 $Y2=0
cc_242 B2 N_B1_c_398_n 0.0313312f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_243 N_B2_c_359_n N_B1_c_398_n 0.018109f $X=3.105 $Y=1.465 $X2=0 $Y2=0
cc_244 B2 N_B1_c_399_n 0.00709945f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_245 N_B2_c_359_n N_B1_c_399_n 0.00164981f $X=3.105 $Y=1.465 $X2=0 $Y2=0
cc_246 N_B2_M1008_g B1 0.00219671f $X=2.885 $Y=2.67 $X2=0 $Y2=0
cc_247 B2 B1 0.0539061f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_248 N_B2_c_359_n B1 9.63288e-19 $X=3.105 $Y=1.465 $X2=0 $Y2=0
cc_249 N_B2_M1008_g N_B1_c_403_n 0.0578692f $X=2.885 $Y=2.67 $X2=0 $Y2=0
cc_250 B2 N_B1_c_403_n 0.00679929f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_251 N_B2_c_359_n N_B1_c_403_n 0.00387758f $X=3.105 $Y=1.465 $X2=0 $Y2=0
cc_252 N_B2_M1008_g N_VPWR_c_448_n 0.00160764f $X=2.885 $Y=2.67 $X2=0 $Y2=0
cc_253 N_B2_M1008_g N_VPWR_c_451_n 0.00491903f $X=2.885 $Y=2.67 $X2=0 $Y2=0
cc_254 N_B2_M1008_g N_VPWR_c_444_n 0.00520574f $X=2.885 $Y=2.67 $X2=0 $Y2=0
cc_255 N_B2_M1006_g N_VGND_c_499_n 0.00878665f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_256 N_B2_M1006_g N_VGND_c_501_n 0.00362954f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_257 N_B2_M1006_g N_VGND_c_503_n 0.00438424f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_258 N_B2_M1006_g N_A_506_47#_c_552_n 8.78457e-19 $X=2.885 $Y=0.445 $X2=0
+ $Y2=0
cc_259 N_B2_M1006_g N_A_506_47#_c_553_n 0.0151724f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_260 B2 N_A_506_47#_c_553_n 0.0475503f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_261 N_B2_c_359_n N_A_506_47#_c_553_n 0.00249734f $X=3.105 $Y=1.465 $X2=0
+ $Y2=0
cc_262 N_B1_M1002_g N_VPWR_c_448_n 0.0121489f $X=3.275 $Y=2.67 $X2=0 $Y2=0
cc_263 B1 N_VPWR_c_448_n 0.0169267f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_264 N_B1_c_403_n N_VPWR_c_448_n 0.00196913f $X=3.585 $Y=2.035 $X2=0 $Y2=0
cc_265 N_B1_M1002_g N_VPWR_c_451_n 0.00432588f $X=3.275 $Y=2.67 $X2=0 $Y2=0
cc_266 N_B1_M1002_g N_VPWR_c_444_n 0.00437282f $X=3.275 $Y=2.67 $X2=0 $Y2=0
cc_267 N_B1_M1000_g N_VGND_c_499_n 0.00981726f $X=3.315 $Y=0.445 $X2=0 $Y2=0
cc_268 N_B1_M1000_g N_VGND_c_502_n 0.00362954f $X=3.315 $Y=0.445 $X2=0 $Y2=0
cc_269 N_B1_M1000_g N_VGND_c_503_n 0.00540867f $X=3.315 $Y=0.445 $X2=0 $Y2=0
cc_270 N_B1_M1000_g N_A_506_47#_c_553_n 0.0128309f $X=3.315 $Y=0.445 $X2=0 $Y2=0
cc_271 N_B1_c_399_n N_A_506_47#_c_553_n 0.0079459f $X=3.585 $Y=0.985 $X2=0 $Y2=0
cc_272 N_B1_M1000_g N_A_506_47#_c_555_n 0.00202753f $X=3.315 $Y=0.445 $X2=0
+ $Y2=0
cc_273 N_X_c_433_n N_VPWR_c_445_n 0.0505127f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_274 N_X_c_433_n N_VPWR_c_449_n 0.0178111f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_275 N_X_M1011_s N_VPWR_c_444_n 0.00371702f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_276 N_X_c_433_n N_VPWR_c_444_n 0.0100304f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_277 N_X_c_433_n N_VGND_c_500_n 0.0178111f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_278 N_X_M1005_s N_VGND_c_503_n 0.00371702f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_279 N_X_c_433_n N_VGND_c_503_n 0.0100304f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_280 N_VGND_c_503_n N_A_506_47#_M1003_d 0.00284838f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_281 N_VGND_c_503_n N_A_506_47#_M1000_d 0.00237353f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_501_n N_A_506_47#_c_552_n 0.0117313f $X=2.935 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_503_n N_A_506_47#_c_552_n 0.00853596f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_499_n N_A_506_47#_c_553_n 0.0205535f $X=3.1 $Y=0.445 $X2=0 $Y2=0
cc_285 N_VGND_c_501_n N_A_506_47#_c_553_n 0.00238864f $X=2.935 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_502_n N_A_506_47#_c_553_n 0.00238864f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_c_503_n N_A_506_47#_c_553_n 0.00919325f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_288 N_VGND_c_502_n N_A_506_47#_c_555_n 0.015222f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_289 N_VGND_c_503_n N_A_506_47#_c_555_n 0.00987569f $X=3.6 $Y=0 $X2=0 $Y2=0
