* File: sky130_fd_sc_lp__o311a_1.spice
* Created: Fri Aug 28 11:13:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o311a_1.pex.spice"
.subckt sky130_fd_sc_lp__o311a_1  VNB VPB A1 A2 A3 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2667 AS=0.2226 PD=1.475 PS=2.21 NRD=8.568 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1011 N_A_267_47#_M1011_d N_A1_M1011_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1449 AS=0.2667 PD=1.185 PS=1.475 NRD=9.276 NRS=42.132 M=1 R=5.6 SA=75001
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_267_47#_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1827 AS=0.1449 PD=1.275 PS=1.185 NRD=11.424 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1005 N_A_267_47#_M1005_d N_A3_M1005_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1827 PD=1.23 PS=1.275 NRD=8.568 NRS=10.704 M=1 R=5.6 SA=75002.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1007 A_591_47# N_B1_M1007_g N_A_267_47#_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1638 PD=1.05 PS=1.23 NRD=7.14 NRS=7.14 M=1 R=5.6 SA=75002.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_A_80_21#_M1008_d N_C1_M1008_g A_591_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75003
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_80_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.3339 PD=1.65 PS=3.05 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1006 A_267_367# N_A1_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.18585 AS=0.2457 PD=1.555 PS=1.65 NRD=14.4598 NRS=6.2449 M=1 R=8.4
+ SA=75000.7 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1010 A_356_367# N_A2_M1010_g A_267_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.19215
+ AS=0.18585 PD=1.565 PS=1.555 NRD=15.2281 NRS=14.4598 M=1 R=8.4 SA=75001.2
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1000 N_A_80_21#_M1000_d N_A3_M1000_g A_356_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.19215 PD=1.65 PS=1.565 NRD=7.8012 NRS=15.2281 M=1 R=8.4
+ SA=75001.6 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_A_80_21#_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=7.8012 NRS=9.3772 M=1 R=8.4 SA=75002.2
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1009 N_A_80_21#_M1009_d N_C1_M1009_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3717 AS=0.2457 PD=3.11 PS=1.65 NRD=4.6886 NRS=9.3772 M=1 R=8.4 SA=75002.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o311a_1.pxi.spice"
*
.ends
*
*
