* File: sky130_fd_sc_lp__a2111o_2.pxi.spice
* Created: Fri Aug 28 09:45:57 2020
* 
x_PM_SKY130_FD_SC_LP__A2111O_2%A_86_275# N_A_86_275#_M1004_d N_A_86_275#_M1000_d
+ N_A_86_275#_M1008_s N_A_86_275#_M1005_g N_A_86_275#_c_75_n N_A_86_275#_M1003_g
+ N_A_86_275#_M1010_g N_A_86_275#_c_77_n N_A_86_275#_M1006_g N_A_86_275#_c_78_n
+ N_A_86_275#_c_79_n N_A_86_275#_c_145_p N_A_86_275#_c_86_n N_A_86_275#_c_87_n
+ N_A_86_275#_c_88_n N_A_86_275#_c_89_n N_A_86_275#_c_108_p N_A_86_275#_c_80_n
+ N_A_86_275#_c_121_p N_A_86_275#_c_81_n N_A_86_275#_c_82_n
+ PM_SKY130_FD_SC_LP__A2111O_2%A_86_275#
x_PM_SKY130_FD_SC_LP__A2111O_2%D1 N_D1_M1004_g N_D1_M1008_g D1 D1 N_D1_c_170_n
+ PM_SKY130_FD_SC_LP__A2111O_2%D1
x_PM_SKY130_FD_SC_LP__A2111O_2%C1 N_C1_M1011_g N_C1_M1009_g C1 C1 C1 C1
+ N_C1_c_204_n N_C1_c_205_n PM_SKY130_FD_SC_LP__A2111O_2%C1
x_PM_SKY130_FD_SC_LP__A2111O_2%B1 N_B1_M1001_g N_B1_M1000_g B1 N_B1_c_242_n
+ N_B1_c_243_n PM_SKY130_FD_SC_LP__A2111O_2%B1
x_PM_SKY130_FD_SC_LP__A2111O_2%A1 N_A1_M1013_g N_A1_M1007_g A1 A1 A1 A1
+ N_A1_c_273_n N_A1_c_274_n PM_SKY130_FD_SC_LP__A2111O_2%A1
x_PM_SKY130_FD_SC_LP__A2111O_2%A2 N_A2_M1002_g N_A2_M1012_g A2 A2 N_A2_c_312_n
+ N_A2_c_313_n PM_SKY130_FD_SC_LP__A2111O_2%A2
x_PM_SKY130_FD_SC_LP__A2111O_2%VPWR N_VPWR_M1005_s N_VPWR_M1010_s N_VPWR_M1007_d
+ N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n
+ N_VPWR_c_344_n VPWR N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_338_n
+ N_VPWR_c_348_n PM_SKY130_FD_SC_LP__A2111O_2%VPWR
x_PM_SKY130_FD_SC_LP__A2111O_2%X N_X_M1003_d N_X_M1005_d X X X X X X X
+ N_X_c_393_n X PM_SKY130_FD_SC_LP__A2111O_2%X
x_PM_SKY130_FD_SC_LP__A2111O_2%A_607_367# N_A_607_367#_M1001_d
+ N_A_607_367#_M1012_d N_A_607_367#_c_416_n N_A_607_367#_c_430_n
+ N_A_607_367#_c_418_n N_A_607_367#_c_414_n N_A_607_367#_c_415_n
+ PM_SKY130_FD_SC_LP__A2111O_2%A_607_367#
x_PM_SKY130_FD_SC_LP__A2111O_2%VGND N_VGND_M1003_s N_VGND_M1006_s N_VGND_M1009_d
+ N_VGND_M1002_d N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n N_VGND_c_439_n
+ N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n VGND N_VGND_c_443_n
+ N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_446_n N_VGND_c_447_n
+ PM_SKY130_FD_SC_LP__A2111O_2%VGND
cc_1 VNB N_A_86_275#_M1005_g 0.01034f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_2 VNB N_A_86_275#_c_75_n 0.0210923f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.195
cc_3 VNB N_A_86_275#_M1010_g 0.00651209f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_4 VNB N_A_86_275#_c_77_n 0.019138f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.195
cc_5 VNB N_A_86_275#_c_78_n 0.00193398f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.36
cc_6 VNB N_A_86_275#_c_79_n 0.00995373f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=1.09
cc_7 VNB N_A_86_275#_c_80_n 0.00886054f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=1.09
cc_8 VNB N_A_86_275#_c_81_n 0.00516572f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.09
cc_9 VNB N_A_86_275#_c_82_n 0.0916935f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.36
cc_10 VNB N_D1_M1004_g 0.0283801f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.835
cc_11 VNB D1 0.00744981f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.525
cc_12 VNB N_D1_c_170_n 0.0251558f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.195
cc_13 VNB N_C1_M1009_g 0.0250735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_C1_c_204_n 0.0240964f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_15 VNB N_C1_c_205_n 0.00398335f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_16 VNB N_B1_M1000_g 0.0258392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_242_n 0.0241338f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_18 VNB N_B1_c_243_n 0.00395826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1007_g 0.0063713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A1 0.0040074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_273_n 0.0314394f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.525
cc_22 VNB N_A1_c_274_n 0.0174156f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_23 VNB N_A2_M1012_g 0.00705037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB A2 0.0385266f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.525
cc_25 VNB N_A2_c_312_n 0.0339104f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.525
cc_26 VNB N_A2_c_313_n 0.0235354f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_27 VNB N_VPWR_c_338_n 0.203486f $X=-0.19 $Y=-0.245 $X2=3.212 $Y2=1.005
cc_28 VNB N_X_c_393_n 0.00188086f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.92
cc_29 VNB N_VGND_c_436_n 0.0135455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_437_n 0.0467451f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.665
cc_31 VNB N_VGND_c_438_n 0.0150365f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.525
cc_32 VNB N_VGND_c_439_n 0.00526884f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.195
cc_33 VNB N_VGND_c_440_n 0.0342778f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.92
cc_34 VNB N_VGND_c_441_n 0.0315793f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.36
cc_35 VNB N_VGND_c_442_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=1.09
cc_36 VNB N_VGND_c_443_n 0.0142356f $X=-0.19 $Y=-0.245 $X2=3.23 $Y2=0.42
cc_37 VNB N_VGND_c_444_n 0.26364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_445_n 0.0157126f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.36
cc_39 VNB N_VGND_c_446_n 0.0195555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_447_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_A_86_275#_M1005_g 0.0264709f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_42 VPB N_A_86_275#_M1010_g 0.0215129f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_43 VPB N_A_86_275#_c_78_n 0.00634092f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=1.36
cc_44 VPB N_A_86_275#_c_86_n 0.0175414f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=2.01
cc_45 VPB N_A_86_275#_c_87_n 0.00537031f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=2.01
cc_46 VPB N_A_86_275#_c_88_n 6.41923e-19 $X=-0.19 $Y=1.655 $X2=1.845 $Y2=2.1
cc_47 VPB N_A_86_275#_c_89_n 0.0127162f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=2.95
cc_48 VPB N_D1_M1008_g 0.0222863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB D1 0.00970561f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.525
cc_50 VPB N_D1_c_170_n 0.00662171f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.195
cc_51 VPB N_C1_M1011_g 0.0187356f $X=-0.19 $Y=1.655 $X2=1.72 $Y2=1.835
cc_52 VPB N_C1_c_204_n 0.00637715f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_53 VPB N_C1_c_205_n 0.00142082f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_54 VPB N_B1_M1001_g 0.0211385f $X=-0.19 $Y=1.655 $X2=1.72 $Y2=1.835
cc_55 VPB N_B1_c_242_n 0.0063779f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_56 VPB N_B1_c_243_n 0.00418555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A1_M1007_g 0.0222171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB A1 0.00251074f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A2_M1012_g 0.027094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB A2 0.0202751f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.525
cc_61 VPB N_VPWR_c_339_n 0.0112967f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.525
cc_62 VPB N_VPWR_c_340_n 0.0645061f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_63 VPB N_VPWR_c_341_n 0.0129119f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_64 VPB N_VPWR_c_342_n 0.0055721f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.665
cc_65 VPB N_VPWR_c_343_n 0.0637184f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=1.92
cc_66 VPB N_VPWR_c_344_n 0.00631825f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=1.36
cc_67 VPB N_VPWR_c_345_n 0.0131811f $X=-0.19 $Y=1.655 $X2=2.18 $Y2=1.09
cc_68 VPB N_VPWR_c_346_n 0.0266055f $X=-0.19 $Y=1.655 $X2=2.42 $Y2=1.09
cc_69 VPB N_VPWR_c_338_n 0.0730238f $X=-0.19 $Y=1.655 $X2=3.212 $Y2=1.005
cc_70 VPB N_VPWR_c_348_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.3 $Y2=1.09
cc_71 VPB N_X_c_393_n 0.00186627f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=1.92
cc_72 VPB N_A_607_367#_c_414_n 0.0075582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_607_367#_c_415_n 0.0377822f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.665
cc_74 N_A_86_275#_c_78_n N_D1_M1004_g 0.0012399f $X=1.25 $Y=1.36 $X2=0 $Y2=0
cc_75 N_A_86_275#_c_79_n N_D1_M1004_g 0.0153192f $X=2.18 $Y=1.09 $X2=0 $Y2=0
cc_76 N_A_86_275#_c_82_n N_D1_M1004_g 0.00372197f $X=1.015 $Y=1.36 $X2=0 $Y2=0
cc_77 N_A_86_275#_c_78_n N_D1_M1008_g 0.00349577f $X=1.25 $Y=1.36 $X2=0 $Y2=0
cc_78 N_A_86_275#_c_88_n N_D1_M1008_g 0.00307689f $X=1.845 $Y=2.1 $X2=0 $Y2=0
cc_79 N_A_86_275#_c_89_n N_D1_M1008_g 0.0185018f $X=1.845 $Y=2.95 $X2=0 $Y2=0
cc_80 N_A_86_275#_c_78_n D1 0.0350135f $X=1.25 $Y=1.36 $X2=0 $Y2=0
cc_81 N_A_86_275#_c_79_n D1 0.0459542f $X=2.18 $Y=1.09 $X2=0 $Y2=0
cc_82 N_A_86_275#_c_86_n D1 0.00764975f $X=1.68 $Y=2.01 $X2=0 $Y2=0
cc_83 N_A_86_275#_c_88_n D1 0.0263376f $X=1.845 $Y=2.1 $X2=0 $Y2=0
cc_84 N_A_86_275#_c_81_n D1 0.00673322f $X=2.3 $Y=1.09 $X2=0 $Y2=0
cc_85 N_A_86_275#_c_82_n D1 0.0016814f $X=1.015 $Y=1.36 $X2=0 $Y2=0
cc_86 N_A_86_275#_c_78_n N_D1_c_170_n 8.38487e-19 $X=1.25 $Y=1.36 $X2=0 $Y2=0
cc_87 N_A_86_275#_c_79_n N_D1_c_170_n 0.0040357f $X=2.18 $Y=1.09 $X2=0 $Y2=0
cc_88 N_A_86_275#_c_88_n N_D1_c_170_n 0.00102542f $X=1.845 $Y=2.1 $X2=0 $Y2=0
cc_89 N_A_86_275#_c_82_n N_D1_c_170_n 0.00515643f $X=1.015 $Y=1.36 $X2=0 $Y2=0
cc_90 N_A_86_275#_c_88_n N_C1_M1011_g 4.75178e-19 $X=1.845 $Y=2.1 $X2=0 $Y2=0
cc_91 N_A_86_275#_c_89_n N_C1_M1011_g 0.00284393f $X=1.845 $Y=2.95 $X2=0 $Y2=0
cc_92 N_A_86_275#_c_108_p N_C1_M1009_g 0.00972953f $X=2.275 $Y=0.42 $X2=0 $Y2=0
cc_93 N_A_86_275#_c_80_n N_C1_M1009_g 0.0132238f $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_94 N_A_86_275#_c_81_n N_C1_M1009_g 0.00137043f $X=2.3 $Y=1.09 $X2=0 $Y2=0
cc_95 N_A_86_275#_c_80_n N_C1_c_204_n 7.75442e-19 $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_96 N_A_86_275#_c_81_n N_C1_c_204_n 0.00338698f $X=2.3 $Y=1.09 $X2=0 $Y2=0
cc_97 N_A_86_275#_c_88_n N_C1_c_205_n 0.00703009f $X=1.845 $Y=2.1 $X2=0 $Y2=0
cc_98 N_A_86_275#_c_89_n N_C1_c_205_n 0.0318438f $X=1.845 $Y=2.95 $X2=0 $Y2=0
cc_99 N_A_86_275#_c_80_n N_C1_c_205_n 0.0294299f $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_100 N_A_86_275#_c_108_p N_B1_M1000_g 4.86841e-19 $X=2.275 $Y=0.42 $X2=0 $Y2=0
cc_101 N_A_86_275#_c_80_n N_B1_M1000_g 0.0151743f $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_102 N_A_86_275#_c_80_n N_B1_c_242_n 0.00327218f $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_103 N_A_86_275#_c_80_n N_B1_c_243_n 0.0282362f $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_104 N_A_86_275#_c_80_n A1 0.0140015f $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_105 N_A_86_275#_c_121_p A1 0.052656f $X=3.23 $Y=0.42 $X2=0 $Y2=0
cc_106 N_A_86_275#_c_80_n N_A1_c_274_n 0.00102292f $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_107 N_A_86_275#_c_121_p N_A1_c_274_n 0.00349894f $X=3.23 $Y=0.42 $X2=0 $Y2=0
cc_108 N_A_86_275#_c_78_n N_VPWR_M1010_s 9.34534e-19 $X=1.25 $Y=1.36 $X2=0 $Y2=0
cc_109 N_A_86_275#_c_87_n N_VPWR_M1010_s 0.0042407f $X=1.415 $Y=2.01 $X2=0 $Y2=0
cc_110 N_A_86_275#_M1005_g N_VPWR_c_340_n 0.0237276f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_111 N_A_86_275#_M1010_g N_VPWR_c_340_n 0.00105122f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_112 N_A_86_275#_M1005_g N_VPWR_c_341_n 9.1342e-19 $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_86_275#_M1010_g N_VPWR_c_341_n 0.0183734f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_86_275#_c_87_n N_VPWR_c_341_n 0.0224079f $X=1.415 $Y=2.01 $X2=0 $Y2=0
cc_115 N_A_86_275#_c_89_n N_VPWR_c_341_n 0.0395279f $X=1.845 $Y=2.95 $X2=0 $Y2=0
cc_116 N_A_86_275#_c_89_n N_VPWR_c_343_n 0.0210467f $X=1.845 $Y=2.95 $X2=0 $Y2=0
cc_117 N_A_86_275#_M1005_g N_VPWR_c_345_n 0.00486043f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_86_275#_M1010_g N_VPWR_c_345_n 0.00486043f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_A_86_275#_M1008_s N_VPWR_c_338_n 0.00215158f $X=1.72 $Y=1.835 $X2=0
+ $Y2=0
cc_120 N_A_86_275#_M1005_g N_VPWR_c_338_n 0.00835506f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_A_86_275#_M1010_g N_VPWR_c_338_n 0.00835506f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_A_86_275#_c_89_n N_VPWR_c_338_n 0.0125689f $X=1.845 $Y=2.95 $X2=0 $Y2=0
cc_123 N_A_86_275#_M1010_g X 0.00324005f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_86_275#_M1005_g N_X_c_393_n 0.0084223f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_86_275#_c_75_n N_X_c_393_n 0.0159788f $X=0.585 $Y=1.195 $X2=0 $Y2=0
cc_126 N_A_86_275#_M1010_g N_X_c_393_n 0.00784164f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_86_275#_c_77_n N_X_c_393_n 0.00136961f $X=1.015 $Y=1.195 $X2=0 $Y2=0
cc_128 N_A_86_275#_c_78_n N_X_c_393_n 0.053298f $X=1.25 $Y=1.36 $X2=0 $Y2=0
cc_129 N_A_86_275#_c_145_p N_X_c_393_n 0.0107682f $X=1.415 $Y=1.09 $X2=0 $Y2=0
cc_130 N_A_86_275#_c_82_n N_X_c_393_n 0.0313213f $X=1.015 $Y=1.36 $X2=0 $Y2=0
cc_131 N_A_86_275#_c_79_n N_VGND_M1006_s 0.00646723f $X=2.18 $Y=1.09 $X2=0 $Y2=0
cc_132 N_A_86_275#_c_145_p N_VGND_M1006_s 0.00305331f $X=1.415 $Y=1.09 $X2=0
+ $Y2=0
cc_133 N_A_86_275#_c_80_n N_VGND_M1009_d 0.00297421f $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_134 N_A_86_275#_c_75_n N_VGND_c_437_n 0.00659675f $X=0.585 $Y=1.195 $X2=0
+ $Y2=0
cc_135 N_A_86_275#_c_82_n N_VGND_c_437_n 0.00104326f $X=1.015 $Y=1.36 $X2=0
+ $Y2=0
cc_136 N_A_86_275#_c_108_p N_VGND_c_438_n 0.0143246f $X=2.275 $Y=0.42 $X2=0
+ $Y2=0
cc_137 N_A_86_275#_c_80_n N_VGND_c_439_n 0.0195425f $X=3.09 $Y=1.09 $X2=0 $Y2=0
cc_138 N_A_86_275#_c_121_p N_VGND_c_441_n 0.0151354f $X=3.23 $Y=0.42 $X2=0 $Y2=0
cc_139 N_A_86_275#_M1004_d N_VGND_c_444_n 0.00380103f $X=2.135 $Y=0.245 $X2=0
+ $Y2=0
cc_140 N_A_86_275#_M1000_d N_VGND_c_444_n 0.00580876f $X=3.09 $Y=0.245 $X2=0
+ $Y2=0
cc_141 N_A_86_275#_c_75_n N_VGND_c_444_n 0.0104567f $X=0.585 $Y=1.195 $X2=0
+ $Y2=0
cc_142 N_A_86_275#_c_77_n N_VGND_c_444_n 0.00820931f $X=1.015 $Y=1.195 $X2=0
+ $Y2=0
cc_143 N_A_86_275#_c_108_p N_VGND_c_444_n 0.00916141f $X=2.275 $Y=0.42 $X2=0
+ $Y2=0
cc_144 N_A_86_275#_c_121_p N_VGND_c_444_n 0.00944728f $X=3.23 $Y=0.42 $X2=0
+ $Y2=0
cc_145 N_A_86_275#_c_75_n N_VGND_c_445_n 0.00524356f $X=0.585 $Y=1.195 $X2=0
+ $Y2=0
cc_146 N_A_86_275#_c_77_n N_VGND_c_445_n 0.00477554f $X=1.015 $Y=1.195 $X2=0
+ $Y2=0
cc_147 N_A_86_275#_c_75_n N_VGND_c_446_n 7.01485e-19 $X=0.585 $Y=1.195 $X2=0
+ $Y2=0
cc_148 N_A_86_275#_c_77_n N_VGND_c_446_n 0.0118432f $X=1.015 $Y=1.195 $X2=0
+ $Y2=0
cc_149 N_A_86_275#_c_79_n N_VGND_c_446_n 0.043371f $X=2.18 $Y=1.09 $X2=0 $Y2=0
cc_150 N_A_86_275#_c_145_p N_VGND_c_446_n 0.0261207f $X=1.415 $Y=1.09 $X2=0
+ $Y2=0
cc_151 N_A_86_275#_c_82_n N_VGND_c_446_n 0.00152877f $X=1.015 $Y=1.36 $X2=0
+ $Y2=0
cc_152 N_D1_M1008_g N_C1_M1011_g 0.05543f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_153 N_D1_M1004_g N_C1_M1009_g 0.0243766f $X=2.06 $Y=0.665 $X2=0 $Y2=0
cc_154 D1 N_C1_c_204_n 0.0028362f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_155 N_D1_c_170_n N_C1_c_204_n 0.05543f $X=1.97 $Y=1.51 $X2=0 $Y2=0
cc_156 N_D1_M1008_g N_C1_c_205_n 0.00399641f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_157 D1 N_C1_c_205_n 0.0341707f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_158 N_D1_c_170_n N_C1_c_205_n 3.50526e-19 $X=1.97 $Y=1.51 $X2=0 $Y2=0
cc_159 N_D1_M1008_g N_VPWR_c_341_n 0.00358434f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_160 N_D1_M1008_g N_VPWR_c_343_n 0.0054895f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_161 N_D1_M1008_g N_VPWR_c_338_n 0.0111524f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_162 N_D1_M1004_g N_VGND_c_438_n 0.00477554f $X=2.06 $Y=0.665 $X2=0 $Y2=0
cc_163 N_D1_M1004_g N_VGND_c_444_n 0.00823465f $X=2.06 $Y=0.665 $X2=0 $Y2=0
cc_164 N_D1_M1004_g N_VGND_c_446_n 0.0117829f $X=2.06 $Y=0.665 $X2=0 $Y2=0
cc_165 N_C1_M1011_g N_B1_M1001_g 0.0412094f $X=2.42 $Y=2.465 $X2=0 $Y2=0
cc_166 N_C1_M1009_g N_B1_M1000_g 0.0193804f $X=2.49 $Y=0.665 $X2=0 $Y2=0
cc_167 N_C1_c_204_n N_B1_c_242_n 0.0204266f $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_168 N_C1_c_205_n N_B1_c_242_n 0.0181671f $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_169 N_C1_c_204_n N_B1_c_243_n 2.88118e-19 $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_170 N_C1_c_205_n N_B1_c_243_n 0.0324081f $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_171 N_C1_M1011_g N_VPWR_c_343_n 0.00490733f $X=2.42 $Y=2.465 $X2=0 $Y2=0
cc_172 N_C1_c_205_n N_VPWR_c_343_n 0.0138393f $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_173 N_C1_M1011_g N_VPWR_c_338_n 0.00857725f $X=2.42 $Y=2.465 $X2=0 $Y2=0
cc_174 N_C1_c_205_n N_VPWR_c_338_n 0.0131331f $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_175 N_C1_c_205_n A_499_367# 0.021893f $X=2.51 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_176 N_C1_M1009_g N_VGND_c_438_n 0.00569184f $X=2.49 $Y=0.665 $X2=0 $Y2=0
cc_177 N_C1_M1009_g N_VGND_c_439_n 0.0016792f $X=2.49 $Y=0.665 $X2=0 $Y2=0
cc_178 N_C1_M1009_g N_VGND_c_444_n 0.0107005f $X=2.49 $Y=0.665 $X2=0 $Y2=0
cc_179 N_C1_M1009_g N_VGND_c_446_n 6.89652e-19 $X=2.49 $Y=0.665 $X2=0 $Y2=0
cc_180 N_B1_M1001_g N_A1_M1007_g 0.0251159f $X=2.96 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B1_M1000_g A1 9.67021e-19 $X=3.015 $Y=0.665 $X2=0 $Y2=0
cc_182 N_B1_c_242_n A1 3.06284e-19 $X=3.05 $Y=1.51 $X2=0 $Y2=0
cc_183 N_B1_c_243_n A1 0.0285742f $X=3.05 $Y=1.51 $X2=0 $Y2=0
cc_184 N_B1_c_242_n N_A1_c_273_n 0.0199537f $X=3.05 $Y=1.51 $X2=0 $Y2=0
cc_185 N_B1_c_243_n N_A1_c_273_n 0.00274442f $X=3.05 $Y=1.51 $X2=0 $Y2=0
cc_186 N_B1_M1000_g N_A1_c_274_n 0.018437f $X=3.015 $Y=0.665 $X2=0 $Y2=0
cc_187 N_B1_M1001_g N_VPWR_c_343_n 0.00585385f $X=2.96 $Y=2.465 $X2=0 $Y2=0
cc_188 N_B1_M1001_g N_VPWR_c_338_n 0.011557f $X=2.96 $Y=2.465 $X2=0 $Y2=0
cc_189 N_B1_c_242_n N_A_607_367#_c_416_n 8.82341e-19 $X=3.05 $Y=1.51 $X2=0 $Y2=0
cc_190 N_B1_c_243_n N_A_607_367#_c_416_n 0.0193141f $X=3.05 $Y=1.51 $X2=0 $Y2=0
cc_191 N_B1_M1000_g N_VGND_c_439_n 0.00316453f $X=3.015 $Y=0.665 $X2=0 $Y2=0
cc_192 N_B1_M1000_g N_VGND_c_441_n 0.00575161f $X=3.015 $Y=0.665 $X2=0 $Y2=0
cc_193 N_B1_M1000_g N_VGND_c_444_n 0.0109524f $X=3.015 $Y=0.665 $X2=0 $Y2=0
cc_194 N_A1_M1007_g A2 6.16974e-19 $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_195 A1 A2 0.046905f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_196 N_A1_c_273_n A2 0.00113445f $X=3.59 $Y=1.36 $X2=0 $Y2=0
cc_197 N_A1_M1007_g N_A2_c_312_n 0.0288594f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_198 A1 N_A2_c_312_n 0.00173804f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_199 A1 N_A2_c_313_n 0.0101411f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_200 N_A1_c_273_n N_A2_c_313_n 0.0212998f $X=3.59 $Y=1.36 $X2=0 $Y2=0
cc_201 N_A1_c_274_n N_A2_c_313_n 0.0289656f $X=3.59 $Y=1.195 $X2=0 $Y2=0
cc_202 N_A1_M1007_g N_VPWR_c_342_n 0.00422051f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A1_M1007_g N_VPWR_c_343_n 0.00585385f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A1_M1007_g N_VPWR_c_338_n 0.0111121f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A1_M1007_g N_A_607_367#_c_418_n 0.0159822f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_206 A1 N_A_607_367#_c_418_n 0.0188972f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_207 N_A1_c_273_n N_A_607_367#_c_418_n 6.70567e-19 $X=3.59 $Y=1.36 $X2=0 $Y2=0
cc_208 N_A1_M1007_g N_A_607_367#_c_415_n 7.55964e-19 $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_209 A1 N_VGND_c_440_n 0.0352449f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_210 N_A1_c_274_n N_VGND_c_440_n 0.0017418f $X=3.59 $Y=1.195 $X2=0 $Y2=0
cc_211 A1 N_VGND_c_441_n 0.0129583f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_212 N_A1_c_274_n N_VGND_c_441_n 0.00476198f $X=3.59 $Y=1.195 $X2=0 $Y2=0
cc_213 A1 N_VGND_c_444_n 0.00986055f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_214 N_A1_c_274_n N_VGND_c_444_n 0.00869467f $X=3.59 $Y=1.195 $X2=0 $Y2=0
cc_215 A1 A_715_49# 0.0109871f $X=3.515 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_216 N_A2_M1012_g N_VPWR_c_342_n 0.00422051f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A2_M1012_g N_VPWR_c_346_n 0.00571722f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A2_M1012_g N_VPWR_c_338_n 0.0116614f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A2_M1012_g N_A_607_367#_c_418_n 0.012833f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_220 A2 N_A_607_367#_c_418_n 0.0107715f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_221 N_A2_M1012_g N_A_607_367#_c_414_n 2.78462e-19 $X=4.04 $Y=2.465 $X2=0
+ $Y2=0
cc_222 A2 N_A_607_367#_c_414_n 0.0246779f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_223 N_A2_c_312_n N_A_607_367#_c_414_n 7.65208e-19 $X=4.13 $Y=1.375 $X2=0
+ $Y2=0
cc_224 N_A2_M1012_g N_A_607_367#_c_415_n 0.0130023f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_225 A2 N_VGND_c_440_n 0.0260007f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_226 N_A2_c_312_n N_VGND_c_440_n 0.00401953f $X=4.13 $Y=1.375 $X2=0 $Y2=0
cc_227 N_A2_c_313_n N_VGND_c_440_n 0.0206311f $X=4.13 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A2_c_313_n N_VGND_c_441_n 0.00477554f $X=4.13 $Y=1.21 $X2=0 $Y2=0
cc_229 N_A2_c_313_n N_VGND_c_444_n 0.0085718f $X=4.13 $Y=1.21 $X2=0 $Y2=0
cc_230 N_VPWR_c_338_n N_X_M1005_d 0.00549325f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_231 N_VPWR_c_345_n X 0.00839145f $X=0.985 $Y=3.33 $X2=0 $Y2=0
cc_232 N_VPWR_c_338_n X 0.00702584f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_233 N_VPWR_c_340_n N_X_c_393_n 0.0452309f $X=0.29 $Y=1.98 $X2=0 $Y2=0
cc_234 N_VPWR_c_338_n A_427_367# 0.00899413f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_235 N_VPWR_c_338_n A_499_367# 0.00644098f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_236 N_VPWR_c_338_n N_A_607_367#_M1001_d 0.00526034f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_237 N_VPWR_c_338_n N_A_607_367#_M1012_d 0.00215158f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_343_n N_A_607_367#_c_430_n 0.0212513f $X=3.605 $Y=3.33 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_338_n N_A_607_367#_c_430_n 0.0127519f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_240 N_VPWR_M1007_d N_A_607_367#_c_418_n 0.00968267f $X=3.575 $Y=1.835 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_342_n N_A_607_367#_c_418_n 0.022455f $X=3.77 $Y=2.39 $X2=0 $Y2=0
cc_242 N_VPWR_c_346_n N_A_607_367#_c_415_n 0.0200241f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_338_n N_A_607_367#_c_415_n 0.0120544f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_244 N_X_c_393_n N_VGND_c_437_n 0.0316864f $X=0.8 $Y=0.42 $X2=0 $Y2=0
cc_245 N_X_M1003_d N_VGND_c_444_n 0.00380103f $X=0.66 $Y=0.245 $X2=0 $Y2=0
cc_246 N_X_c_393_n N_VGND_c_444_n 0.0101905f $X=0.8 $Y=0.42 $X2=0 $Y2=0
cc_247 N_X_c_393_n N_VGND_c_445_n 0.0163698f $X=0.8 $Y=0.42 $X2=0 $Y2=0
cc_248 N_VGND_c_444_n A_715_49# 0.00979873f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
