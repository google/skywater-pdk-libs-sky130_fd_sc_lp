* NGSPICE file created from sky130_fd_sc_lp__einvn_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__einvn_m A TE_B VGND VNB VPB VPWR Z
M1000 a_218_154# a_47_154# VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.218e+11p ps=1.42e+06u
M1001 Z A a_218_154# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1002 VPWR TE_B a_47_154# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.113e+11p ps=1.37e+06u
M1003 Z A a_232_535# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1004 VGND TE_B a_47_154# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 a_232_535# TE_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

