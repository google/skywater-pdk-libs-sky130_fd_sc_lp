* File: sky130_fd_sc_lp__buf_0.pxi.spice
* Created: Wed Sep  2 09:34:35 2020
* 
x_PM_SKY130_FD_SC_LP__BUF_0%A_70_157# N_A_70_157#_M1000_d N_A_70_157#_M1002_d
+ N_A_70_157#_M1003_g N_A_70_157#_M1001_g N_A_70_157#_c_42_n N_A_70_157#_c_43_n
+ N_A_70_157#_c_44_n N_A_70_157#_c_45_n N_A_70_157#_c_56_p N_A_70_157#_c_46_n
+ N_A_70_157#_c_47_n N_A_70_157#_c_52_n N_A_70_157#_c_53_n N_A_70_157#_c_54_n
+ N_A_70_157#_c_48_n N_A_70_157#_c_49_n N_A_70_157#_c_73_p
+ PM_SKY130_FD_SC_LP__BUF_0%A_70_157#
x_PM_SKY130_FD_SC_LP__BUF_0%A N_A_M1000_g N_A_M1002_g N_A_c_105_n N_A_c_110_n A
+ A N_A_c_107_n PM_SKY130_FD_SC_LP__BUF_0%A
x_PM_SKY130_FD_SC_LP__BUF_0%X N_X_M1003_s N_X_M1001_s N_X_c_137_n N_X_c_138_n
+ N_X_c_139_n X X X N_X_c_142_n X PM_SKY130_FD_SC_LP__BUF_0%X
x_PM_SKY130_FD_SC_LP__BUF_0%VPWR N_VPWR_M1001_d N_VPWR_c_161_n VPWR
+ N_VPWR_c_162_n N_VPWR_c_163_n N_VPWR_c_160_n N_VPWR_c_165_n
+ PM_SKY130_FD_SC_LP__BUF_0%VPWR
x_PM_SKY130_FD_SC_LP__BUF_0%VGND N_VGND_M1003_d N_VGND_c_180_n VGND
+ N_VGND_c_181_n N_VGND_c_182_n N_VGND_c_183_n N_VGND_c_184_n
+ PM_SKY130_FD_SC_LP__BUF_0%VGND
cc_1 VNB N_A_70_157#_M1001_g 0.0106151f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_2 VNB N_A_70_157#_c_42_n 0.0202868f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.785
cc_3 VNB N_A_70_157#_c_43_n 0.0252112f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.29
cc_4 VNB N_A_70_157#_c_44_n 0.0187856f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.455
cc_5 VNB N_A_70_157#_c_45_n 0.00126117f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.97
cc_6 VNB N_A_70_157#_c_46_n 0.00130162f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.055
cc_7 VNB N_A_70_157#_c_47_n 0.0200884f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=0.877
cc_8 VNB N_A_70_157#_c_48_n 0.0201034f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=0.465
cc_9 VNB N_A_70_157#_c_49_n 0.0164556f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.95
cc_10 VNB N_A_M1000_g 0.0484974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_105_n 0.0229627f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_12 VNB A 0.0224808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_c_107_n 0.0183728f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.97
cc_14 VNB N_X_c_137_n 0.013105f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_15 VNB N_X_c_138_n 0.00566523f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.95
cc_16 VNB N_X_c_139_n 0.0456001f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.785
cc_17 VNB N_VPWR_c_160_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.455
cc_18 VNB N_VGND_c_180_n 0.00631596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_181_n 0.0173033f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.455
cc_20 VNB N_VGND_c_182_n 0.0172072f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.455
cc_21 VNB N_VGND_c_183_n 0.112472f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.97
cc_22 VNB N_VGND_c_184_n 0.00632255f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.055
cc_23 VPB N_A_70_157#_M1001_g 0.0548539f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_24 VPB N_A_70_157#_c_46_n 0.00317422f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.055
cc_25 VPB N_A_70_157#_c_52_n 0.0206871f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=2.14
cc_26 VPB N_A_70_157#_c_53_n 0.00186744f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.14
cc_27 VPB N_A_70_157#_c_54_n 0.0366562f $X=-0.19 $Y=1.655 $X2=1.18 $Y2=2.845
cc_28 VPB N_A_M1002_g 0.065066f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.785
cc_29 VPB N_A_c_105_n 0.00544866f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_30 VPB N_A_c_110_n 0.0191852f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_31 VPB A 0.0117645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_X_c_138_n 0.00380479f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.95
cc_33 VPB X 0.0342248f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.29
cc_34 VPB N_X_c_142_n 0.0227712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB X 0.008666f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.877
cc_36 VPB N_VPWR_c_161_n 0.0101908f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_162_n 0.0173715f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_38 VPB N_VPWR_c_163_n 0.0183088f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.33
cc_39 VPB N_VPWR_c_160_n 0.0514514f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.455
cc_40 VPB N_VPWR_c_165_n 0.00487564f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.877
cc_41 N_A_70_157#_c_42_n N_A_M1000_g 0.00972807f $X=0.515 $Y=0.785 $X2=0 $Y2=0
cc_42 N_A_70_157#_c_56_p N_A_M1000_g 0.0011139f $X=0.555 $Y=1.33 $X2=0 $Y2=0
cc_43 N_A_70_157#_c_47_n N_A_M1000_g 0.0133867f $X=1.06 $Y=0.877 $X2=0 $Y2=0
cc_44 N_A_70_157#_c_48_n N_A_M1000_g 0.00497392f $X=1.18 $Y=0.465 $X2=0 $Y2=0
cc_45 N_A_70_157#_c_49_n N_A_M1000_g 0.0139175f $X=0.515 $Y=0.95 $X2=0 $Y2=0
cc_46 N_A_70_157#_c_52_n N_A_M1002_g 0.0147452f $X=0.995 $Y=2.14 $X2=0 $Y2=0
cc_47 N_A_70_157#_c_54_n N_A_M1002_g 0.0210628f $X=1.18 $Y=2.845 $X2=0 $Y2=0
cc_48 N_A_70_157#_M1001_g N_A_c_105_n 0.0448231f $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_49 N_A_70_157#_c_44_n N_A_c_105_n 0.0139175f $X=0.515 $Y=1.455 $X2=0 $Y2=0
cc_50 N_A_70_157#_c_46_n N_A_c_105_n 0.00636958f $X=0.595 $Y=2.055 $X2=0 $Y2=0
cc_51 N_A_70_157#_c_52_n N_A_c_110_n 0.0014092f $X=0.995 $Y=2.14 $X2=0 $Y2=0
cc_52 N_A_70_157#_M1001_g A 4.54057e-19 $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_53 N_A_70_157#_c_43_n A 0.00105662f $X=0.515 $Y=1.29 $X2=0 $Y2=0
cc_54 N_A_70_157#_c_56_p A 0.0474854f $X=0.555 $Y=1.33 $X2=0 $Y2=0
cc_55 N_A_70_157#_c_47_n A 0.0380128f $X=1.06 $Y=0.877 $X2=0 $Y2=0
cc_56 N_A_70_157#_c_52_n A 0.0393638f $X=0.995 $Y=2.14 $X2=0 $Y2=0
cc_57 N_A_70_157#_c_43_n N_A_c_107_n 0.0139175f $X=0.515 $Y=1.29 $X2=0 $Y2=0
cc_58 N_A_70_157#_c_47_n N_A_c_107_n 0.00116231f $X=1.06 $Y=0.877 $X2=0 $Y2=0
cc_59 N_A_70_157#_c_73_p N_A_c_107_n 0.0011139f $X=0.555 $Y=1.455 $X2=0 $Y2=0
cc_60 N_A_70_157#_M1001_g N_X_c_138_n 0.0184936f $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_61 N_A_70_157#_c_46_n N_X_c_138_n 0.0331288f $X=0.595 $Y=2.055 $X2=0 $Y2=0
cc_62 N_A_70_157#_M1001_g N_X_c_139_n 0.00309373f $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_63 N_A_70_157#_c_42_n N_X_c_139_n 0.00547137f $X=0.515 $Y=0.785 $X2=0 $Y2=0
cc_64 N_A_70_157#_c_45_n N_X_c_139_n 0.0147409f $X=0.555 $Y=0.97 $X2=0 $Y2=0
cc_65 N_A_70_157#_c_56_p N_X_c_139_n 0.0355813f $X=0.555 $Y=1.33 $X2=0 $Y2=0
cc_66 N_A_70_157#_c_46_n N_X_c_139_n 0.00799321f $X=0.595 $Y=2.055 $X2=0 $Y2=0
cc_67 N_A_70_157#_c_49_n N_X_c_139_n 0.0164669f $X=0.515 $Y=0.95 $X2=0 $Y2=0
cc_68 N_A_70_157#_c_53_n X 0.0139714f $X=0.68 $Y=2.14 $X2=0 $Y2=0
cc_69 N_A_70_157#_c_54_n X 0.00465459f $X=1.18 $Y=2.845 $X2=0 $Y2=0
cc_70 N_A_70_157#_M1001_g X 9.09997e-19 $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_71 N_A_70_157#_M1001_g N_VPWR_c_161_n 0.00295743f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_72 N_A_70_157#_c_52_n N_VPWR_c_161_n 0.0121245f $X=0.995 $Y=2.14 $X2=0 $Y2=0
cc_73 N_A_70_157#_c_53_n N_VPWR_c_161_n 0.0101662f $X=0.68 $Y=2.14 $X2=0 $Y2=0
cc_74 N_A_70_157#_c_54_n N_VPWR_c_161_n 0.0523563f $X=1.18 $Y=2.845 $X2=0 $Y2=0
cc_75 N_A_70_157#_M1001_g N_VPWR_c_162_n 0.00545548f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_76 N_A_70_157#_c_54_n N_VPWR_c_163_n 0.0247924f $X=1.18 $Y=2.845 $X2=0 $Y2=0
cc_77 N_A_70_157#_M1001_g N_VPWR_c_160_n 0.0111663f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_78 N_A_70_157#_c_54_n N_VPWR_c_160_n 0.0133281f $X=1.18 $Y=2.845 $X2=0 $Y2=0
cc_79 N_A_70_157#_c_42_n N_VGND_c_180_n 0.00329138f $X=0.515 $Y=0.785 $X2=0
+ $Y2=0
cc_80 N_A_70_157#_c_45_n N_VGND_c_180_n 0.0080426f $X=0.555 $Y=0.97 $X2=0 $Y2=0
cc_81 N_A_70_157#_c_47_n N_VGND_c_180_n 0.0143832f $X=1.06 $Y=0.877 $X2=0 $Y2=0
cc_82 N_A_70_157#_c_49_n N_VGND_c_180_n 7.90821e-19 $X=0.515 $Y=0.95 $X2=0 $Y2=0
cc_83 N_A_70_157#_c_42_n N_VGND_c_181_n 0.00565115f $X=0.515 $Y=0.785 $X2=0
+ $Y2=0
cc_84 N_A_70_157#_c_48_n N_VGND_c_182_n 0.0144999f $X=1.18 $Y=0.465 $X2=0 $Y2=0
cc_85 N_A_70_157#_c_42_n N_VGND_c_183_n 0.00785936f $X=0.515 $Y=0.785 $X2=0
+ $Y2=0
cc_86 N_A_70_157#_c_45_n N_VGND_c_183_n 0.00486696f $X=0.555 $Y=0.97 $X2=0 $Y2=0
cc_87 N_A_70_157#_c_47_n N_VGND_c_183_n 0.00585097f $X=1.06 $Y=0.877 $X2=0 $Y2=0
cc_88 N_A_70_157#_c_48_n N_VGND_c_183_n 0.0107504f $X=1.18 $Y=0.465 $X2=0 $Y2=0
cc_89 N_A_70_157#_c_49_n N_VGND_c_183_n 2.61071e-19 $X=0.515 $Y=0.95 $X2=0 $Y2=0
cc_90 N_A_M1002_g N_VPWR_c_161_n 0.0077567f $X=0.965 $Y=2.845 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_VPWR_c_163_n 0.00482865f $X=0.965 $Y=2.845 $X2=0 $Y2=0
cc_92 N_A_M1002_g N_VPWR_c_160_n 0.00965865f $X=0.965 $Y=2.845 $X2=0 $Y2=0
cc_93 N_A_M1000_g N_VGND_c_180_n 0.0033548f $X=0.965 $Y=0.465 $X2=0 $Y2=0
cc_94 N_A_M1000_g N_VGND_c_182_n 0.005634f $X=0.965 $Y=0.465 $X2=0 $Y2=0
cc_95 N_A_M1000_g N_VGND_c_183_n 0.00691709f $X=0.965 $Y=0.465 $X2=0 $Y2=0
cc_96 X N_VPWR_c_161_n 0.0294212f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_97 N_X_c_142_n N_VPWR_c_162_n 0.0220795f $X=0.26 $Y=2.56 $X2=0 $Y2=0
cc_98 N_X_c_142_n N_VPWR_c_160_n 0.0119743f $X=0.26 $Y=2.56 $X2=0 $Y2=0
cc_99 N_X_c_137_n N_VGND_c_181_n 0.0155464f $X=0.26 $Y=0.45 $X2=0 $Y2=0
cc_100 N_X_c_137_n N_VGND_c_183_n 0.0112574f $X=0.26 $Y=0.45 $X2=0 $Y2=0
