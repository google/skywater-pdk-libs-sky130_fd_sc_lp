# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__fa_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__fa_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 7.105000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 2.495000 1.920000 2.785000 1.965000 ;
        RECT 2.495000 2.105000 2.785000 2.150000 ;
        RECT 6.815000 1.920000 7.105000 1.965000 ;
        RECT 6.815000 2.105000 7.105000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.450000 1.095000 3.935000 1.165000 ;
        RECT 3.450000 1.165000 5.495000 1.185000 ;
        RECT 3.450000 1.185000 6.630000 1.355000 ;
        RECT 5.915000 1.355000 6.630000 1.825000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.865000 3.715000 2.120000 ;
        RECT 3.505000 2.120000 3.715000 2.940000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.365000 1.815000 ;
        RECT 0.085000 1.815000 0.375000 3.075000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.573300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.640000 0.255000 8.075000 1.020000 ;
        RECT 7.795000 1.815000 8.075000 3.075000 ;
        RECT 7.840000 1.020000 8.075000 1.815000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.535000  0.085000 1.200000 1.045000 ;
      RECT 0.535000  1.215000 0.795000 1.545000 ;
      RECT 0.555000  1.545000 0.795000 2.300000 ;
      RECT 0.555000  2.300000 1.920000 2.470000 ;
      RECT 0.555000  2.640000 0.885000 3.245000 ;
      RECT 1.005000  1.295000 1.345000 2.130000 ;
      RECT 1.630000  2.470000 1.920000 2.655000 ;
      RECT 1.700000  0.730000 1.985000 1.525000 ;
      RECT 1.700000  1.525000 5.700000 1.695000 ;
      RECT 1.700000  1.695000 1.920000 2.300000 ;
      RECT 2.090000  2.300000 3.335000 2.470000 ;
      RECT 2.090000  2.470000 2.390000 2.660000 ;
      RECT 2.155000  0.730000 2.390000 1.185000 ;
      RECT 2.155000  1.185000 3.280000 1.355000 ;
      RECT 2.365000  1.865000 2.785000 2.130000 ;
      RECT 2.560000  0.085000 2.890000 1.015000 ;
      RECT 2.570000  2.640000 2.900000 3.245000 ;
      RECT 3.060000  0.730000 3.280000 1.185000 ;
      RECT 3.080000  2.470000 3.335000 2.660000 ;
      RECT 3.635000  0.085000 3.935000 0.795000 ;
      RECT 3.885000  2.100000 4.120000 3.245000 ;
      RECT 4.105000  0.465000 4.345000 0.825000 ;
      RECT 4.105000  0.825000 5.495000 0.995000 ;
      RECT 4.290000  1.865000 5.435000 2.035000 ;
      RECT 4.290000  2.035000 4.535000 2.430000 ;
      RECT 4.515000  0.085000 4.845000 0.655000 ;
      RECT 4.705000  2.205000 5.035000 2.470000 ;
      RECT 4.845000  2.470000 5.035000 3.245000 ;
      RECT 5.015000  0.385000 5.495000 0.825000 ;
      RECT 5.205000  2.035000 5.435000 2.430000 ;
      RECT 5.605000  2.100000 5.875000 2.300000 ;
      RECT 5.605000  2.300000 7.625000 2.470000 ;
      RECT 5.665000  0.665000 6.970000 0.845000 ;
      RECT 5.665000  0.845000 7.470000 1.015000 ;
      RECT 6.820000  1.185000 7.120000 2.130000 ;
      RECT 7.140000  0.085000 7.470000 0.675000 ;
      RECT 7.285000  2.640000 7.615000 3.245000 ;
      RECT 7.290000  1.015000 7.470000 1.190000 ;
      RECT 7.290000  1.190000 7.660000 1.520000 ;
      RECT 7.290000  1.520000 7.625000 2.300000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  1.950000 1.285000 2.120000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.950000 2.725000 2.120000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  1.950000 7.045000 2.120000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__fa_1
