# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__buflp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__buflp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 1.055000 2.805000 2.890000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.646800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.550000 1.375000 2.735000 ;
        RECT 1.115000 0.595000 1.445000 1.095000 ;
        RECT 1.115000 1.095000 1.375000 1.550000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.095000 ;
      RECT 0.115000  1.815000 0.445000 3.245000 ;
      RECT 0.615000  0.255000 1.945000 0.425000 ;
      RECT 0.615000  0.425000 0.945000 1.095000 ;
      RECT 0.615000  1.815000 0.865000 2.905000 ;
      RECT 0.615000  2.905000 1.805000 3.075000 ;
      RECT 1.555000  1.815000 1.805000 2.905000 ;
      RECT 1.615000  0.425000 1.945000 1.095000 ;
      RECT 1.825000  1.265000 2.285000 1.595000 ;
      RECT 1.975000  1.815000 2.305000 3.245000 ;
      RECT 2.115000  0.085000 2.445000 0.545000 ;
      RECT 2.115000  0.715000 3.245000 0.885000 ;
      RECT 2.115000  0.885000 2.285000 1.265000 ;
      RECT 2.915000  0.255000 3.245000 0.715000 ;
      RECT 2.990000  0.885000 3.245000 2.545000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__buflp_2
END LIBRARY
