* File: sky130_fd_sc_lp__edfxbp_1.pxi.spice
* Created: Wed Sep  2 09:51:18 2020
* 
x_PM_SKY130_FD_SC_LP__EDFXBP_1%DE N_DE_M1007_g N_DE_M1001_g N_DE_c_272_n
+ N_DE_M1022_g N_DE_c_274_n N_DE_M1005_g N_DE_c_275_n N_DE_c_276_n DE DE DE
+ N_DE_c_278_n N_DE_c_279_n DE PM_SKY130_FD_SC_LP__EDFXBP_1%DE
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_120_179# N_A_120_179#_M1007_d
+ N_A_120_179#_M1001_d N_A_120_179#_M1002_g N_A_120_179#_M1026_g
+ N_A_120_179#_c_331_n N_A_120_179#_c_332_n N_A_120_179#_c_333_n
+ N_A_120_179#_c_334_n N_A_120_179#_c_335_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_120_179#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%D N_D_M1025_g N_D_M1029_g D N_D_c_395_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%D
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_587_350# N_A_587_350#_M1024_s
+ N_A_587_350#_M1034_s N_A_587_350#_M1003_g N_A_587_350#_c_446_n
+ N_A_587_350#_c_447_n N_A_587_350#_M1017_g N_A_587_350#_M1016_g
+ N_A_587_350#_M1019_g N_A_587_350#_c_435_n N_A_587_350#_c_436_n
+ N_A_587_350#_M1000_g N_A_587_350#_M1010_g N_A_587_350#_c_438_n
+ N_A_587_350#_c_439_n N_A_587_350#_c_440_n N_A_587_350#_c_441_n
+ N_A_587_350#_c_442_n N_A_587_350#_c_455_n N_A_587_350#_c_456_n
+ N_A_587_350#_c_457_n N_A_587_350#_c_520_p N_A_587_350#_c_443_n
+ N_A_587_350#_c_444_n PM_SKY130_FD_SC_LP__EDFXBP_1%A_587_350#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_958_290# N_A_958_290#_M1032_d
+ N_A_958_290#_M1021_d N_A_958_290#_M1033_g N_A_958_290#_M1011_g
+ N_A_958_290#_M1004_g N_A_958_290#_M1006_g N_A_958_290#_c_654_n
+ N_A_958_290#_c_641_n N_A_958_290#_c_642_n N_A_958_290#_c_643_n
+ N_A_958_290#_c_644_n N_A_958_290#_c_645_n N_A_958_290#_c_656_n
+ N_A_958_290#_c_646_n N_A_958_290#_c_647_n N_A_958_290#_c_648_n
+ N_A_958_290#_c_649_n N_A_958_290#_c_650_n N_A_958_290#_c_651_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_958_290#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_1067_65# N_A_1067_65#_M1035_d
+ N_A_1067_65#_M1015_d N_A_1067_65#_M1014_g N_A_1067_65#_c_785_n
+ N_A_1067_65#_M1027_g N_A_1067_65#_M1028_g N_A_1067_65#_M1009_g
+ N_A_1067_65#_c_787_n N_A_1067_65#_c_788_n N_A_1067_65#_c_798_n
+ N_A_1067_65#_c_789_n N_A_1067_65#_c_799_n N_A_1067_65#_c_800_n
+ N_A_1067_65#_c_801_n N_A_1067_65#_c_802_n N_A_1067_65#_c_803_n
+ N_A_1067_65#_c_887_p N_A_1067_65#_c_804_n N_A_1067_65#_c_805_n
+ N_A_1067_65#_c_823_n N_A_1067_65#_c_806_n N_A_1067_65#_c_807_n
+ N_A_1067_65#_c_790_n N_A_1067_65#_c_791_n N_A_1067_65#_c_792_n
+ N_A_1067_65#_c_793_n N_A_1067_65#_c_794_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_1067_65#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_902_396# N_A_902_396#_M1013_d
+ N_A_902_396#_M1008_d N_A_902_396#_c_981_n N_A_902_396#_M1035_g
+ N_A_902_396#_M1015_g N_A_902_396#_c_983_n N_A_902_396#_c_984_n
+ N_A_902_396#_c_985_n N_A_902_396#_c_1000_n N_A_902_396#_c_986_n
+ N_A_902_396#_c_987_n PM_SKY130_FD_SC_LP__EDFXBP_1%A_902_396#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%CLK N_CLK_c_1053_n N_CLK_M1023_g N_CLK_M1018_g
+ N_CLK_c_1055_n N_CLK_c_1061_n N_CLK_c_1056_n CLK N_CLK_c_1058_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%CLK
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_872_324# N_A_872_324#_M1018_s
+ N_A_872_324#_M1023_s N_A_872_324#_M1008_g N_A_872_324#_M1013_g
+ N_A_872_324#_c_1123_n N_A_872_324#_c_1124_n N_A_872_324#_M1032_g
+ N_A_872_324#_M1021_g N_A_872_324#_c_1109_n N_A_872_324#_c_1127_n
+ N_A_872_324#_M1030_g N_A_872_324#_M1020_g N_A_872_324#_c_1111_n
+ N_A_872_324#_c_1112_n N_A_872_324#_c_1113_n N_A_872_324#_c_1114_n
+ N_A_872_324#_c_1131_n N_A_872_324#_c_1115_n N_A_872_324#_c_1116_n
+ N_A_872_324#_c_1117_n N_A_872_324#_c_1118_n N_A_872_324#_c_1119_n
+ N_A_872_324#_c_1231_n N_A_872_324#_c_1120_n N_A_872_324#_c_1121_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_872_324#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_1865_367# N_A_1865_367#_M1020_d
+ N_A_1865_367#_M1030_d N_A_1865_367#_c_1280_n N_A_1865_367#_c_1281_n
+ N_A_1865_367#_c_1282_n N_A_1865_367#_c_1283_n N_A_1865_367#_M1024_g
+ N_A_1865_367#_M1034_g N_A_1865_367#_c_1285_n N_A_1865_367#_M1012_g
+ N_A_1865_367#_M1031_g N_A_1865_367#_c_1287_n N_A_1865_367#_c_1299_n
+ N_A_1865_367#_c_1300_n N_A_1865_367#_c_1301_n N_A_1865_367#_c_1288_n
+ N_A_1865_367#_c_1302_n N_A_1865_367#_c_1289_n N_A_1865_367#_c_1303_n
+ N_A_1865_367#_c_1304_n N_A_1865_367#_c_1305_n N_A_1865_367#_c_1290_n
+ N_A_1865_367#_c_1291_n N_A_1865_367#_c_1292_n N_A_1865_367#_c_1293_n
+ N_A_1865_367#_c_1307_n N_A_1865_367#_c_1294_n N_A_1865_367#_c_1295_n
+ N_A_1865_367#_c_1296_n PM_SKY130_FD_SC_LP__EDFXBP_1%A_1865_367#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%VPWR N_VPWR_M1001_s N_VPWR_M1005_d N_VPWR_M1027_d
+ N_VPWR_M1023_d N_VPWR_M1009_d N_VPWR_M1034_d N_VPWR_M1031_s N_VPWR_c_1463_n
+ N_VPWR_c_1464_n N_VPWR_c_1465_n N_VPWR_c_1466_n N_VPWR_c_1467_n
+ N_VPWR_c_1468_n N_VPWR_c_1469_n N_VPWR_c_1470_n N_VPWR_c_1471_n
+ N_VPWR_c_1472_n N_VPWR_c_1473_n N_VPWR_c_1474_n N_VPWR_c_1475_n
+ N_VPWR_c_1476_n VPWR N_VPWR_c_1477_n N_VPWR_c_1478_n N_VPWR_c_1479_n
+ N_VPWR_c_1480_n N_VPWR_c_1462_n N_VPWR_c_1482_n N_VPWR_c_1483_n
+ N_VPWR_c_1484_n PM_SKY130_FD_SC_LP__EDFXBP_1%VPWR
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_286_423# N_A_286_423#_M1005_s
+ N_A_286_423#_M1003_d N_A_286_423#_c_1602_n N_A_286_423#_c_1603_n
+ N_A_286_423#_c_1604_n N_A_286_423#_c_1605_n N_A_286_423#_c_1606_n
+ N_A_286_423#_c_1607_n N_A_286_423#_c_1608_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_286_423#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_531_423# N_A_531_423#_M1029_d
+ N_A_531_423#_M1013_s N_A_531_423#_M1025_d N_A_531_423#_M1033_d
+ N_A_531_423#_c_1658_n N_A_531_423#_c_1659_n N_A_531_423#_c_1660_n
+ N_A_531_423#_c_1652_n N_A_531_423#_c_1653_n N_A_531_423#_c_1654_n
+ N_A_531_423#_c_1655_n N_A_531_423#_c_1656_n N_A_531_423#_c_1663_n
+ N_A_531_423#_c_1664_n N_A_531_423#_c_1665_n N_A_531_423#_c_1657_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_531_423#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_761_396# N_A_761_396#_M1008_s
+ N_A_761_396#_M1027_s N_A_761_396#_c_1743_n N_A_761_396#_c_1744_n
+ N_A_761_396#_c_1745_n N_A_761_396#_c_1746_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_761_396#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_1781_367# N_A_1781_367#_M1030_s
+ N_A_1781_367#_M1009_s N_A_1781_367#_c_1776_n N_A_1781_367#_c_1777_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_1781_367#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_1971_388# N_A_1971_388#_M1004_d
+ N_A_1971_388#_M1019_d N_A_1971_388#_c_1799_n N_A_1971_388#_c_1800_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_1971_388#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%Q_N N_Q_N_M1000_d N_Q_N_M1010_d N_Q_N_c_1827_n
+ N_Q_N_c_1828_n Q_N Q_N N_Q_N_c_1836_n PM_SKY130_FD_SC_LP__EDFXBP_1%Q_N
x_PM_SKY130_FD_SC_LP__EDFXBP_1%Q N_Q_M1012_d N_Q_M1031_d N_Q_c_1855_n Q Q Q Q Q
+ N_Q_c_1854_n Q PM_SKY130_FD_SC_LP__EDFXBP_1%Q
x_PM_SKY130_FD_SC_LP__EDFXBP_1%VGND N_VGND_M1007_s N_VGND_M1022_d N_VGND_M1014_d
+ N_VGND_M1018_d N_VGND_M1028_d N_VGND_M1024_d N_VGND_M1012_s N_VGND_c_1867_n
+ N_VGND_c_1868_n N_VGND_c_1869_n N_VGND_c_1870_n N_VGND_c_1871_n
+ N_VGND_c_1872_n N_VGND_c_1873_n N_VGND_c_1874_n N_VGND_c_1875_n
+ N_VGND_c_1876_n N_VGND_c_1877_n VGND N_VGND_c_1878_n N_VGND_c_1879_n
+ N_VGND_c_1880_n N_VGND_c_1881_n N_VGND_c_1882_n N_VGND_c_1883_n
+ N_VGND_c_1884_n N_VGND_c_1885_n PM_SKY130_FD_SC_LP__EDFXBP_1%VGND
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_231_53# N_A_231_53#_M1022_s N_A_231_53#_M1029_s
+ N_A_231_53#_c_1992_n N_A_231_53#_c_1993_n N_A_231_53#_c_1994_n
+ N_A_231_53#_c_1995_n N_A_231_53#_c_1996_n N_A_231_53#_c_1997_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_231_53#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_404_53# N_A_404_53#_M1002_d N_A_404_53#_M1017_d
+ N_A_404_53#_c_2028_n N_A_404_53#_c_2029_n N_A_404_53#_c_2030_n
+ PM_SKY130_FD_SC_LP__EDFXBP_1%A_404_53#
x_PM_SKY130_FD_SC_LP__EDFXBP_1%A_1789_141# N_A_1789_141#_M1020_s
+ N_A_1789_141#_M1016_d N_A_1789_141#_c_2049_n N_A_1789_141#_c_2050_n
+ N_A_1789_141#_c_2056_n PM_SKY130_FD_SC_LP__EDFXBP_1%A_1789_141#
cc_1 VNB N_DE_M1007_g 0.0447182f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.105
cc_2 VNB N_DE_M1022_g 0.0714599f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.475
cc_3 VNB N_A_120_179#_M1002_g 0.049841f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.83
cc_4 VNB N_A_120_179#_M1026_g 0.00536619f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.755
cc_5 VNB N_A_120_179#_c_331_n 0.016729f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.005
cc_6 VNB N_A_120_179#_c_332_n 0.00131922f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.88
cc_7 VNB N_A_120_179#_c_333_n 0.029116f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.32
cc_8 VNB N_A_120_179#_c_334_n 0.0369867f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.69
cc_9 VNB N_A_120_179#_c_335_n 0.00121501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_D_M1025_g 0.00890604f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.105
cc_11 VNB N_D_M1029_g 0.0271957f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.725
cc_12 VNB D 0.0057881f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.83
cc_13 VNB N_D_c_395_n 0.0490812f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.755
cc_14 VNB N_A_587_350#_M1017_g 0.0427568f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.475
cc_15 VNB N_A_587_350#_M1016_g 0.0461012f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.325
cc_16 VNB N_A_587_350#_c_435_n 0.00699041f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.32
cc_17 VNB N_A_587_350#_c_436_n 0.00796765f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.69
cc_18 VNB N_A_587_350#_M1000_g 0.028328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_587_350#_c_438_n 0.00296031f $X=-0.19 $Y=-0.245 $X2=1.197
+ $Y2=2.405
cc_20 VNB N_A_587_350#_c_439_n 0.00341484f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.775
cc_21 VNB N_A_587_350#_c_440_n 0.0272115f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.735
cc_22 VNB N_A_587_350#_c_441_n 0.00311624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_587_350#_c_442_n 0.0325902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_587_350#_c_443_n 0.00798324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_587_350#_c_444_n 0.00832913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_958_290#_M1011_g 0.0421068f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.755
cc_27 VNB N_A_958_290#_M1004_g 0.0045641f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.005
cc_28 VNB N_A_958_290#_c_641_n 0.0141303f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.9
cc_29 VNB N_A_958_290#_c_642_n 0.00409609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_958_290#_c_643_n 0.028457f $X=-0.19 $Y=-0.245 $X2=1.197 $Y2=2.735
cc_31 VNB N_A_958_290#_c_644_n 0.0212552f $X=-0.19 $Y=-0.245 $X2=1.197 $Y2=2.035
cc_32 VNB N_A_958_290#_c_645_n 0.0156398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_958_290#_c_646_n 0.00133399f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.797
cc_34 VNB N_A_958_290#_c_647_n 0.0254659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_958_290#_c_648_n 0.00221907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_958_290#_c_649_n 0.020471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_958_290#_c_650_n 0.00717942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_958_290#_c_651_n 0.0130201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1067_65#_M1014_g 0.0226256f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.83
cc_40 VNB N_A_1067_65#_c_785_n 0.0222783f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.735
cc_41 VNB N_A_1067_65#_M1028_g 0.0273606f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.325
cc_42 VNB N_A_1067_65#_c_787_n 0.0175887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1067_65#_c_788_n 0.00308855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1067_65#_c_789_n 0.0243429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1067_65#_c_790_n 0.00202672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1067_65#_c_791_n 0.0421946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1067_65#_c_792_n 0.0244066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1067_65#_c_793_n 0.00447314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1067_65#_c_794_n 0.0149189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_902_396#_c_981_n 0.0233022f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.725
cc_51 VNB N_A_902_396#_M1015_g 0.0224637f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.735
cc_52 VNB N_A_902_396#_c_983_n 0.00529329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_902_396#_c_984_n 0.00764988f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.83
cc_54 VNB N_A_902_396#_c_985_n 0.00497623f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_55 VNB N_A_902_396#_c_986_n 0.0250386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_902_396#_c_987_n 0.047585f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.9
cc_57 VNB N_CLK_c_1053_n 0.0131931f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.755
cc_58 VNB N_CLK_M1018_g 0.0301679f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.83
cc_59 VNB N_CLK_c_1055_n 0.0212821f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.735
cc_60 VNB N_CLK_c_1056_n 0.00411239f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.005
cc_61 VNB CLK 0.00341997f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.325
cc_62 VNB N_CLK_c_1058_n 0.0397391f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.83
cc_63 VNB N_A_872_324#_M1013_g 0.0556742f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.755
cc_64 VNB N_A_872_324#_M1032_g 0.0284157f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.88
cc_65 VNB N_A_872_324#_c_1109_n 0.0256777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_872_324#_M1020_g 0.0422894f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.735
cc_67 VNB N_A_872_324#_c_1111_n 0.00362371f $X=-0.19 $Y=-0.245 $X2=1.197
+ $Y2=2.035
cc_68 VNB N_A_872_324#_c_1112_n 0.00723223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_872_324#_c_1113_n 0.0219211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_872_324#_c_1114_n 0.00348555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_872_324#_c_1115_n 0.00611493f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.9
cc_72 VNB N_A_872_324#_c_1116_n 0.00686318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_872_324#_c_1117_n 0.00950575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_872_324#_c_1118_n 0.00356563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_872_324#_c_1119_n 0.00823641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_872_324#_c_1120_n 0.00469396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_872_324#_c_1121_n 0.0285863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1865_367#_c_1280_n 0.0381744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1865_367#_c_1281_n 0.0191536f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.83
cc_80 VNB N_A_1865_367#_c_1282_n 0.00891301f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.83
cc_81 VNB N_A_1865_367#_c_1283_n 0.0169552f $X=-0.19 $Y=-0.245 $X2=1.16
+ $Y2=2.005
cc_82 VNB N_A_1865_367#_M1034_g 0.0132272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1865_367#_c_1285_n 0.0231018f $X=-0.19 $Y=-0.245 $X2=1.79
+ $Y2=2.325
cc_84 VNB N_A_1865_367#_M1031_g 0.00914772f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.88
cc_85 VNB N_A_1865_367#_c_1287_n 0.0172333f $X=-0.19 $Y=-0.245 $X2=1.115
+ $Y2=2.69
cc_86 VNB N_A_1865_367#_c_1288_n 0.0437001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1865_367#_c_1289_n 0.0141196f $X=-0.19 $Y=-0.245 $X2=1.197
+ $Y2=2.712
cc_88 VNB N_A_1865_367#_c_1290_n 0.00189055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1865_367#_c_1291_n 0.0154438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1865_367#_c_1292_n 0.00298648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1865_367#_c_1293_n 0.00582077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1865_367#_c_1294_n 0.00778697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1865_367#_c_1295_n 0.0118526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1865_367#_c_1296_n 0.0505773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VPWR_c_1462_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_531_423#_c_1652_n 0.00743154f $X=-0.19 $Y=-0.245 $X2=1.79
+ $Y2=2.325
cc_97 VNB N_A_531_423#_c_1653_n 0.00367435f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.83
cc_98 VNB N_A_531_423#_c_1654_n 0.0251607f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.88
cc_99 VNB N_A_531_423#_c_1655_n 0.0147758f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.32
cc_100 VNB N_A_531_423#_c_1656_n 0.011096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_531_423#_c_1657_n 0.00960878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_Q_N_c_1827_n 0.0122208f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.725
cc_103 VNB N_Q_N_c_1828_n 0.00998782f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.735
cc_104 VNB N_Q_c_1854_n 0.0603204f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_105 VNB N_VGND_c_1867_n 0.011635f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.88
cc_106 VNB N_VGND_c_1868_n 0.0813511f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_107 VNB N_VGND_c_1869_n 0.00550208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1870_n 0.0109069f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.9
cc_109 VNB N_VGND_c_1871_n 0.0220245f $X=-0.19 $Y=-0.245 $X2=1.197 $Y2=2.735
cc_110 VNB N_VGND_c_1872_n 0.0136026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1873_n 0.0665646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1874_n 0.0136687f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.735
cc_113 VNB N_VGND_c_1875_n 0.0386691f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.797
cc_114 VNB N_VGND_c_1876_n 0.0132033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1877_n 0.0190879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1878_n 0.0340309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1879_n 0.0947344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1880_n 0.0528521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1881_n 0.0199125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1882_n 0.823537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1883_n 0.003823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1884_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1885_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_231_53#_c_1992_n 0.0244913f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.83
cc_125 VNB N_A_231_53#_c_1993_n 0.00426494f $X=-0.19 $Y=-0.245 $X2=1.16
+ $Y2=2.735
cc_126 VNB N_A_231_53#_c_1994_n 0.0156249f $X=-0.19 $Y=-0.245 $X2=1.515
+ $Y2=1.755
cc_127 VNB N_A_231_53#_c_1995_n 0.0090008f $X=-0.19 $Y=-0.245 $X2=1.515
+ $Y2=0.475
cc_128 VNB N_A_231_53#_c_1996_n 0.00315214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_231_53#_c_1997_n 0.00543751f $X=-0.19 $Y=-0.245 $X2=1.79
+ $Y2=2.325
cc_130 VNB N_A_404_53#_c_2028_n 0.0297077f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=2.725
cc_131 VNB N_A_404_53#_c_2029_n 0.00656962f $X=-0.19 $Y=-0.245 $X2=1.16
+ $Y2=2.005
cc_132 VNB N_A_404_53#_c_2030_n 0.00562658f $X=-0.19 $Y=-0.245 $X2=1.515
+ $Y2=1.755
cc_133 VNB N_A_1789_141#_c_2049_n 0.0122867f $X=-0.19 $Y=-0.245 $X2=1.16
+ $Y2=2.735
cc_134 VNB N_A_1789_141#_c_2050_n 0.0079893f $X=-0.19 $Y=-0.245 $X2=1.515
+ $Y2=0.475
cc_135 VPB N_DE_M1007_g 0.00907286f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.105
cc_136 VPB N_DE_M1001_g 0.0562418f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.725
cc_137 VPB N_DE_c_272_n 0.0286191f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.83
cc_138 VPB N_DE_M1022_g 0.00715316f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=0.475
cc_139 VPB N_DE_c_274_n 0.0187656f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=2.005
cc_140 VPB N_DE_c_275_n 0.0106787f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.83
cc_141 VPB N_DE_c_276_n 0.0525378f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=1.88
cc_142 VPB DE 0.00616536f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.95
cc_143 VPB N_DE_c_278_n 0.0441364f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.9
cc_144 VPB N_DE_c_279_n 0.044139f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.735
cc_145 VPB DE 0.00629942f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.775
cc_146 VPB N_A_120_179#_M1026_g 0.0329505f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=1.755
cc_147 VPB N_A_120_179#_c_332_n 0.0129273f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.88
cc_148 VPB N_D_M1025_g 0.0326821f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.105
cc_149 VPB N_A_587_350#_M1003_g 0.0250867f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.83
cc_150 VPB N_A_587_350#_c_446_n 0.0148019f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.005
cc_151 VPB N_A_587_350#_c_447_n 0.00788147f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.735
cc_152 VPB N_A_587_350#_M1019_g 0.0329423f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=1.88
cc_153 VPB N_A_587_350#_c_435_n 0.00720438f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.32
cc_154 VPB N_A_587_350#_c_436_n 0.00893619f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.69
cc_155 VPB N_A_587_350#_M1010_g 0.0247823f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.9
cc_156 VPB N_A_587_350#_c_439_n 0.00560284f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.775
cc_157 VPB N_A_587_350#_c_440_n 0.00597573f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.735
cc_158 VPB N_A_587_350#_c_442_n 0.0432644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_587_350#_c_455_n 0.0575005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_587_350#_c_456_n 0.0151051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_587_350#_c_457_n 0.00615231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_587_350#_c_443_n 0.0256459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_587_350#_c_444_n 0.00744643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_958_290#_M1033_g 0.0259623f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.83
cc_165 VPB N_A_958_290#_M1004_g 0.0323711f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=2.005
cc_166 VPB N_A_958_290#_c_654_n 0.00726764f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.69
cc_167 VPB N_A_958_290#_c_645_n 0.00585997f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_958_290#_c_656_n 9.15619e-19 $X=-0.19 $Y=1.655 $X2=1.197
+ $Y2=2.405
cc_169 VPB N_A_958_290#_c_646_n 4.49516e-19 $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.797
cc_170 VPB N_A_958_290#_c_647_n 0.0187586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_958_290#_c_648_n 0.00132894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_958_290#_c_650_n 0.00123457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_1067_65#_M1027_g 0.0393145f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=0.475
cc_174 VPB N_A_1067_65#_M1009_g 0.0252773f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=1.88
cc_175 VPB N_A_1067_65#_c_788_n 0.00131041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_1067_65#_c_798_n 0.00332315f $X=-0.19 $Y=1.655 $X2=1.197
+ $Y2=2.035
cc_177 VPB N_A_1067_65#_c_799_n 0.0249119f $X=-0.19 $Y=1.655 $X2=1.197 $Y2=2.405
cc_178 VPB N_A_1067_65#_c_800_n 0.00307929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_1067_65#_c_801_n 0.00393533f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.775
cc_180 VPB N_A_1067_65#_c_802_n 0.00519948f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.775
cc_181 VPB N_A_1067_65#_c_803_n 7.61567e-19 $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.735
cc_182 VPB N_A_1067_65#_c_804_n 0.0124332f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_1067_65#_c_805_n 0.00223489f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1067_65#_c_806_n 0.0150337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1067_65#_c_807_n 0.00217114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_1067_65#_c_790_n 0.00130932f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_1067_65#_c_791_n 0.0153394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_1067_65#_c_793_n 0.00193737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1067_65#_c_794_n 0.0265986f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_902_396#_M1015_g 0.0240749f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.735
cc_191 VPB N_A_902_396#_c_984_n 0.00619965f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.83
cc_192 VPB N_CLK_M1023_g 0.0256916f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.905
cc_193 VPB N_CLK_c_1055_n 7.94199e-19 $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.735
cc_194 VPB N_CLK_c_1061_n 0.0187229f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=0.475
cc_195 VPB N_A_872_324#_M1008_g 0.0631452f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.83
cc_196 VPB N_A_872_324#_c_1123_n 0.285394f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=0.475
cc_197 VPB N_A_872_324#_c_1124_n 0.012806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_872_324#_M1021_g 0.0469794f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.69
cc_199 VPB N_A_872_324#_c_1109_n 0.0244318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_872_324#_c_1127_n 0.0226577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_872_324#_c_1111_n 0.00831888f $X=-0.19 $Y=1.655 $X2=1.197
+ $Y2=2.035
cc_202 VPB N_A_872_324#_c_1112_n 0.0223923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_872_324#_c_1114_n 0.00441527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_872_324#_c_1131_n 0.0128806f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.775
cc_205 VPB N_A_872_324#_c_1118_n 0.0026003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_872_324#_c_1120_n 0.00261552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_1865_367#_M1034_g 0.0234842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_1865_367#_M1031_g 0.0269061f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=1.88
cc_209 VPB N_A_1865_367#_c_1299_n 7.33434e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_1865_367#_c_1300_n 0.0166036f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.9
cc_211 VPB N_A_1865_367#_c_1301_n 0.0032951f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.9
cc_212 VPB N_A_1865_367#_c_1302_n 0.0271553f $X=-0.19 $Y=1.655 $X2=1.197
+ $Y2=2.405
cc_213 VPB N_A_1865_367#_c_1303_n 0.00772229f $X=-0.19 $Y=1.655 $X2=1.25
+ $Y2=2.735
cc_214 VPB N_A_1865_367#_c_1304_n 0.014412f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.797
cc_215 VPB N_A_1865_367#_c_1305_n 7.92214e-19 $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.9
cc_216 VPB N_A_1865_367#_c_1290_n 0.00742515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_1865_367#_c_1307_n 0.0113298f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1463_n 0.0116091f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=1.88
cc_219 VPB N_VPWR_c_1464_n 0.042274f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.95
cc_220 VPB N_VPWR_c_1465_n 0.0255434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1466_n 0.0134646f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.9
cc_222 VPB N_VPWR_c_1467_n 0.0150179f $X=-0.19 $Y=1.655 $X2=1.197 $Y2=2.735
cc_223 VPB N_VPWR_c_1468_n 0.00472864f $X=-0.19 $Y=1.655 $X2=1.197 $Y2=2.405
cc_224 VPB N_VPWR_c_1469_n 0.0132746f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.775
cc_225 VPB N_VPWR_c_1470_n 0.00722289f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1471_n 0.0424129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1472_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1473_n 0.0362568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1474_n 0.00223798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1475_n 0.0728107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1476_n 0.0032427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1477_n 0.0980584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1478_n 0.0402592f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1479_n 0.0197055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1480_n 0.0156742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1462_n 0.150543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1482_n 0.00330333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1483_n 0.00526199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1484_n 0.00511034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_286_423#_c_1602_n 0.00517629f $X=-0.19 $Y=1.655 $X2=1.085
+ $Y2=1.83
cc_241 VPB N_A_286_423#_c_1603_n 0.0152549f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.005
cc_242 VPB N_A_286_423#_c_1604_n 0.00143633f $X=-0.19 $Y=1.655 $X2=1.16
+ $Y2=2.735
cc_243 VPB N_A_286_423#_c_1605_n 0.00386981f $X=-0.19 $Y=1.655 $X2=1.515
+ $Y2=0.475
cc_244 VPB N_A_286_423#_c_1606_n 0.023327f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=0.475
cc_245 VPB N_A_286_423#_c_1607_n 0.00365847f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_286_423#_c_1608_n 0.00597824f $X=-0.19 $Y=1.655 $X2=1.79
+ $Y2=2.325
cc_247 VPB N_A_531_423#_c_1658_n 0.00375787f $X=-0.19 $Y=1.655 $X2=1.515
+ $Y2=0.475
cc_248 VPB N_A_531_423#_c_1659_n 0.0100711f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=2.005
cc_249 VPB N_A_531_423#_c_1660_n 0.00189106f $X=-0.19 $Y=1.655 $X2=1.79
+ $Y2=2.325
cc_250 VPB N_A_531_423#_c_1653_n 0.00112638f $X=-0.19 $Y=1.655 $X2=0.525
+ $Y2=1.83
cc_251 VPB N_A_531_423#_c_1656_n 0.00465374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_531_423#_c_1663_n 0.010693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_531_423#_c_1664_n 0.0028528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_531_423#_c_1665_n 0.00920775f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.9
cc_255 VPB N_A_761_396#_c_1743_n 0.0217956f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.83
cc_256 VPB N_A_761_396#_c_1744_n 0.0376224f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.005
cc_257 VPB N_A_761_396#_c_1745_n 0.00900204f $X=-0.19 $Y=1.655 $X2=1.16
+ $Y2=2.735
cc_258 VPB N_A_761_396#_c_1746_n 0.0148701f $X=-0.19 $Y=1.655 $X2=1.515
+ $Y2=0.475
cc_259 VPB N_A_1781_367#_c_1776_n 0.00389272f $X=-0.19 $Y=1.655 $X2=1.16
+ $Y2=2.735
cc_260 VPB N_A_1781_367#_c_1777_n 0.0227427f $X=-0.19 $Y=1.655 $X2=1.515
+ $Y2=1.755
cc_261 VPB N_A_1971_388#_c_1799_n 0.00517015f $X=-0.19 $Y=1.655 $X2=0.525
+ $Y2=2.725
cc_262 VPB N_A_1971_388#_c_1800_n 0.00861896f $X=-0.19 $Y=1.655 $X2=1.16
+ $Y2=2.005
cc_263 VPB N_Q_N_c_1828_n 0.00810101f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.735
cc_264 VPB N_Q_c_1855_n 0.034325f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.83
cc_265 VPB N_Q_c_1854_n 0.0162318f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.95
cc_266 VPB Q 0.00474557f $X=-0.19 $Y=1.655 $X2=1.197 $Y2=2.035
cc_267 N_DE_M1022_g N_A_120_179#_M1002_g 0.0478341f $X=1.515 $Y=0.475 $X2=0
+ $Y2=0
cc_268 N_DE_M1022_g N_A_120_179#_M1026_g 0.00662743f $X=1.515 $Y=0.475 $X2=0
+ $Y2=0
cc_269 N_DE_c_276_n N_A_120_179#_M1026_g 0.0167707f $X=1.515 $Y=1.88 $X2=0 $Y2=0
cc_270 N_DE_M1007_g N_A_120_179#_c_331_n 0.00569753f $X=0.525 $Y=1.105 $X2=0
+ $Y2=0
cc_271 N_DE_M1022_g N_A_120_179#_c_331_n 0.00524816f $X=1.515 $Y=0.475 $X2=0
+ $Y2=0
cc_272 N_DE_M1007_g N_A_120_179#_c_332_n 0.011961f $X=0.525 $Y=1.105 $X2=0 $Y2=0
cc_273 N_DE_M1001_g N_A_120_179#_c_332_n 0.035846f $X=0.525 $Y=2.725 $X2=0 $Y2=0
cc_274 N_DE_c_272_n N_A_120_179#_c_332_n 0.0187527f $X=1.085 $Y=1.83 $X2=0 $Y2=0
cc_275 N_DE_M1022_g N_A_120_179#_c_332_n 0.00468974f $X=1.515 $Y=0.475 $X2=0
+ $Y2=0
cc_276 N_DE_c_275_n N_A_120_179#_c_332_n 0.00651517f $X=0.525 $Y=1.83 $X2=0
+ $Y2=0
cc_277 N_DE_c_276_n N_A_120_179#_c_332_n 0.00979149f $X=1.515 $Y=1.88 $X2=0
+ $Y2=0
cc_278 DE N_A_120_179#_c_332_n 0.0850735f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_279 N_DE_c_272_n N_A_120_179#_c_333_n 0.0151611f $X=1.085 $Y=1.83 $X2=0 $Y2=0
cc_280 N_DE_M1022_g N_A_120_179#_c_333_n 0.0221954f $X=1.515 $Y=0.475 $X2=0
+ $Y2=0
cc_281 N_DE_c_276_n N_A_120_179#_c_333_n 0.00154526f $X=1.515 $Y=1.88 $X2=0
+ $Y2=0
cc_282 DE N_A_120_179#_c_333_n 0.0107668f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_283 N_DE_M1007_g N_A_120_179#_c_335_n 0.0183315f $X=0.525 $Y=1.105 $X2=0
+ $Y2=0
cc_284 N_DE_M1001_g N_VPWR_c_1464_n 0.00476117f $X=0.525 $Y=2.725 $X2=0 $Y2=0
cc_285 N_DE_c_274_n N_VPWR_c_1465_n 0.00177385f $X=1.79 $Y=2.005 $X2=0 $Y2=0
cc_286 DE N_VPWR_c_1465_n 0.00564123f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_287 N_DE_c_278_n N_VPWR_c_1465_n 0.00574368f $X=1.25 $Y=2.9 $X2=0 $Y2=0
cc_288 N_DE_c_279_n N_VPWR_c_1465_n 3.56704e-19 $X=1.25 $Y=2.735 $X2=0 $Y2=0
cc_289 DE N_VPWR_c_1465_n 0.010937f $X=1.2 $Y=2.775 $X2=0 $Y2=0
cc_290 N_DE_M1001_g N_VPWR_c_1471_n 0.00502664f $X=0.525 $Y=2.725 $X2=0 $Y2=0
cc_291 N_DE_c_274_n N_VPWR_c_1471_n 0.00336027f $X=1.79 $Y=2.005 $X2=0 $Y2=0
cc_292 N_DE_c_278_n N_VPWR_c_1471_n 0.00210846f $X=1.25 $Y=2.9 $X2=0 $Y2=0
cc_293 DE N_VPWR_c_1471_n 0.0206493f $X=1.2 $Y=2.775 $X2=0 $Y2=0
cc_294 N_DE_M1001_g N_VPWR_c_1462_n 0.0109943f $X=0.525 $Y=2.725 $X2=0 $Y2=0
cc_295 N_DE_c_274_n N_VPWR_c_1462_n 0.00424893f $X=1.79 $Y=2.005 $X2=0 $Y2=0
cc_296 DE N_VPWR_c_1462_n 0.0124157f $X=1.2 $Y=2.775 $X2=0 $Y2=0
cc_297 N_DE_c_274_n N_A_286_423#_c_1602_n 0.00891915f $X=1.79 $Y=2.005 $X2=0
+ $Y2=0
cc_298 N_DE_c_276_n N_A_286_423#_c_1602_n 0.00772932f $X=1.515 $Y=1.88 $X2=0
+ $Y2=0
cc_299 DE N_A_286_423#_c_1602_n 0.0470174f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_300 N_DE_c_279_n N_A_286_423#_c_1602_n 0.00180215f $X=1.25 $Y=2.735 $X2=0
+ $Y2=0
cc_301 N_DE_c_276_n N_A_286_423#_c_1603_n 0.00891893f $X=1.515 $Y=1.88 $X2=0
+ $Y2=0
cc_302 N_DE_M1022_g N_A_286_423#_c_1604_n 0.00189348f $X=1.515 $Y=0.475 $X2=0
+ $Y2=0
cc_303 N_DE_c_276_n N_A_286_423#_c_1604_n 0.0112694f $X=1.515 $Y=1.88 $X2=0
+ $Y2=0
cc_304 N_DE_c_276_n N_A_286_423#_c_1605_n 7.85943e-19 $X=1.515 $Y=1.88 $X2=0
+ $Y2=0
cc_305 N_DE_M1007_g N_VGND_c_1868_n 0.00593231f $X=0.525 $Y=1.105 $X2=0 $Y2=0
cc_306 N_DE_M1022_g N_VGND_c_1869_n 0.0104467f $X=1.515 $Y=0.475 $X2=0 $Y2=0
cc_307 N_DE_M1007_g N_VGND_c_1878_n 0.00297774f $X=0.525 $Y=1.105 $X2=0 $Y2=0
cc_308 N_DE_M1022_g N_VGND_c_1878_n 0.00461019f $X=1.515 $Y=0.475 $X2=0 $Y2=0
cc_309 N_DE_M1007_g N_VGND_c_1882_n 0.00400849f $X=0.525 $Y=1.105 $X2=0 $Y2=0
cc_310 N_DE_M1022_g N_VGND_c_1882_n 0.00930161f $X=1.515 $Y=0.475 $X2=0 $Y2=0
cc_311 N_DE_M1007_g N_A_231_53#_c_1992_n 0.00272943f $X=0.525 $Y=1.105 $X2=0
+ $Y2=0
cc_312 N_DE_M1022_g N_A_231_53#_c_1992_n 0.00764931f $X=1.515 $Y=0.475 $X2=0
+ $Y2=0
cc_313 N_DE_M1007_g N_A_231_53#_c_1993_n 4.07031e-19 $X=0.525 $Y=1.105 $X2=0
+ $Y2=0
cc_314 N_DE_M1022_g N_A_231_53#_c_1995_n 0.015752f $X=1.515 $Y=0.475 $X2=0 $Y2=0
cc_315 N_A_120_179#_M1026_g N_D_M1025_g 0.0375174f $X=2.22 $Y=2.325 $X2=0 $Y2=0
cc_316 N_A_120_179#_M1002_g D 2.94536e-19 $X=1.945 $Y=0.475 $X2=0 $Y2=0
cc_317 N_A_120_179#_c_333_n D 0.0136746f $X=2.035 $Y=1.4 $X2=0 $Y2=0
cc_318 N_A_120_179#_c_334_n D 6.00425e-19 $X=2.035 $Y=1.4 $X2=0 $Y2=0
cc_319 N_A_120_179#_M1002_g N_D_c_395_n 0.00154587f $X=1.945 $Y=0.475 $X2=0
+ $Y2=0
cc_320 N_A_120_179#_c_333_n N_D_c_395_n 0.00131466f $X=2.035 $Y=1.4 $X2=0 $Y2=0
cc_321 N_A_120_179#_c_334_n N_D_c_395_n 0.0447819f $X=2.035 $Y=1.4 $X2=0 $Y2=0
cc_322 N_A_120_179#_c_332_n N_VPWR_c_1464_n 0.025828f $X=0.74 $Y=2.55 $X2=0
+ $Y2=0
cc_323 N_A_120_179#_M1026_g N_VPWR_c_1465_n 0.00119082f $X=2.22 $Y=2.325 $X2=0
+ $Y2=0
cc_324 N_A_120_179#_c_332_n N_VPWR_c_1471_n 0.0220321f $X=0.74 $Y=2.55 $X2=0
+ $Y2=0
cc_325 N_A_120_179#_M1026_g N_VPWR_c_1477_n 0.00289174f $X=2.22 $Y=2.325 $X2=0
+ $Y2=0
cc_326 N_A_120_179#_M1026_g N_VPWR_c_1462_n 0.00355578f $X=2.22 $Y=2.325 $X2=0
+ $Y2=0
cc_327 N_A_120_179#_c_332_n N_VPWR_c_1462_n 0.0125808f $X=0.74 $Y=2.55 $X2=0
+ $Y2=0
cc_328 N_A_120_179#_M1026_g N_A_286_423#_c_1602_n 6.67538e-19 $X=2.22 $Y=2.325
+ $X2=0 $Y2=0
cc_329 N_A_120_179#_M1026_g N_A_286_423#_c_1603_n 0.0162417f $X=2.22 $Y=2.325
+ $X2=0 $Y2=0
cc_330 N_A_120_179#_c_333_n N_A_286_423#_c_1603_n 0.0334115f $X=2.035 $Y=1.4
+ $X2=0 $Y2=0
cc_331 N_A_120_179#_c_334_n N_A_286_423#_c_1603_n 0.0067107f $X=2.035 $Y=1.4
+ $X2=0 $Y2=0
cc_332 N_A_120_179#_c_332_n N_A_286_423#_c_1604_n 0.00494371f $X=0.74 $Y=2.55
+ $X2=0 $Y2=0
cc_333 N_A_120_179#_c_333_n N_A_286_423#_c_1604_n 0.0203637f $X=2.035 $Y=1.4
+ $X2=0 $Y2=0
cc_334 N_A_120_179#_M1026_g N_A_286_423#_c_1605_n 0.0136702f $X=2.22 $Y=2.325
+ $X2=0 $Y2=0
cc_335 N_A_120_179#_M1026_g N_A_531_423#_c_1658_n 5.18952e-19 $X=2.22 $Y=2.325
+ $X2=0 $Y2=0
cc_336 N_A_120_179#_c_331_n N_VGND_c_1868_n 0.013595f $X=0.74 $Y=1.105 $X2=0
+ $Y2=0
cc_337 N_A_120_179#_c_335_n N_VGND_c_1868_n 0.00475343f $X=0.74 $Y=1.4 $X2=0
+ $Y2=0
cc_338 N_A_120_179#_M1002_g N_VGND_c_1869_n 0.00343738f $X=1.945 $Y=0.475 $X2=0
+ $Y2=0
cc_339 N_A_120_179#_M1002_g N_VGND_c_1879_n 0.00520813f $X=1.945 $Y=0.475 $X2=0
+ $Y2=0
cc_340 N_A_120_179#_M1002_g N_VGND_c_1882_n 0.0107157f $X=1.945 $Y=0.475 $X2=0
+ $Y2=0
cc_341 N_A_120_179#_c_331_n N_A_231_53#_c_1992_n 6.27986e-19 $X=0.74 $Y=1.105
+ $X2=0 $Y2=0
cc_342 N_A_120_179#_c_331_n N_A_231_53#_c_1993_n 0.0121616f $X=0.74 $Y=1.105
+ $X2=0 $Y2=0
cc_343 N_A_120_179#_c_333_n N_A_231_53#_c_1993_n 0.0212368f $X=2.035 $Y=1.4
+ $X2=0 $Y2=0
cc_344 N_A_120_179#_c_333_n N_A_231_53#_c_1994_n 0.00203441f $X=2.035 $Y=1.4
+ $X2=0 $Y2=0
cc_345 N_A_120_179#_c_334_n N_A_231_53#_c_1994_n 0.00392049f $X=2.035 $Y=1.4
+ $X2=0 $Y2=0
cc_346 N_A_120_179#_M1002_g N_A_231_53#_c_1995_n 0.0111542f $X=1.945 $Y=0.475
+ $X2=0 $Y2=0
cc_347 N_A_120_179#_c_333_n N_A_231_53#_c_1995_n 0.0566093f $X=2.035 $Y=1.4
+ $X2=0 $Y2=0
cc_348 N_A_120_179#_M1002_g N_A_231_53#_c_1996_n 0.00687683f $X=1.945 $Y=0.475
+ $X2=0 $Y2=0
cc_349 N_A_120_179#_c_334_n N_A_231_53#_c_1996_n 0.00332999f $X=2.035 $Y=1.4
+ $X2=0 $Y2=0
cc_350 N_A_120_179#_M1002_g N_A_231_53#_c_1997_n 0.00480354f $X=1.945 $Y=0.475
+ $X2=0 $Y2=0
cc_351 N_A_120_179#_M1002_g N_A_404_53#_c_2030_n 0.00450548f $X=1.945 $Y=0.475
+ $X2=0 $Y2=0
cc_352 N_D_M1025_g N_A_587_350#_c_447_n 0.0220011f $X=2.58 $Y=2.325 $X2=0 $Y2=0
cc_353 N_D_c_395_n N_A_587_350#_c_447_n 0.00207777f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_354 N_D_M1029_g N_A_587_350#_M1017_g 0.0230652f $X=2.935 $Y=0.77 $X2=0 $Y2=0
cc_355 D N_A_587_350#_M1017_g 3.10518e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_356 N_D_c_395_n N_A_587_350#_M1017_g 0.00395895f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_357 N_D_M1025_g N_A_587_350#_c_442_n 0.00299748f $X=2.58 $Y=2.325 $X2=0 $Y2=0
cc_358 N_D_M1025_g N_A_286_423#_c_1603_n 0.00125061f $X=2.58 $Y=2.325 $X2=0
+ $Y2=0
cc_359 N_D_M1025_g N_A_286_423#_c_1605_n 0.00521133f $X=2.58 $Y=2.325 $X2=0
+ $Y2=0
cc_360 N_D_M1025_g N_A_286_423#_c_1606_n 0.00654616f $X=2.58 $Y=2.325 $X2=0
+ $Y2=0
cc_361 N_D_M1025_g N_A_286_423#_c_1608_n 5.06423e-19 $X=2.58 $Y=2.325 $X2=0
+ $Y2=0
cc_362 N_D_M1025_g N_A_531_423#_c_1658_n 0.00913736f $X=2.58 $Y=2.325 $X2=0
+ $Y2=0
cc_363 N_D_c_395_n N_A_531_423#_c_1659_n 0.00307955f $X=2.67 $Y=1.345 $X2=0
+ $Y2=0
cc_364 N_D_M1025_g N_A_531_423#_c_1660_n 0.00424622f $X=2.58 $Y=2.325 $X2=0
+ $Y2=0
cc_365 D N_A_531_423#_c_1660_n 0.0134392f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_366 N_D_c_395_n N_A_531_423#_c_1660_n 0.00290174f $X=2.67 $Y=1.345 $X2=0
+ $Y2=0
cc_367 N_D_M1029_g N_A_531_423#_c_1652_n 0.0113174f $X=2.935 $Y=0.77 $X2=0 $Y2=0
cc_368 D N_A_531_423#_c_1652_n 0.0049098f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_369 N_D_M1025_g N_A_531_423#_c_1653_n 0.0038163f $X=2.58 $Y=2.325 $X2=0 $Y2=0
cc_370 D N_A_531_423#_c_1653_n 0.0116363f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_371 N_D_c_395_n N_A_531_423#_c_1653_n 0.00189678f $X=2.67 $Y=1.345 $X2=0
+ $Y2=0
cc_372 N_D_M1029_g N_VGND_c_1879_n 6.24464e-19 $X=2.935 $Y=0.77 $X2=0 $Y2=0
cc_373 D N_A_231_53#_c_1994_n 0.00354389f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_374 N_D_c_395_n N_A_231_53#_c_1994_n 3.36691e-19 $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_375 N_D_M1029_g N_A_231_53#_c_1996_n 0.00129405f $X=2.935 $Y=0.77 $X2=0 $Y2=0
cc_376 N_D_M1029_g N_A_231_53#_c_1997_n 4.43583e-19 $X=2.935 $Y=0.77 $X2=0 $Y2=0
cc_377 D N_A_231_53#_c_1997_n 0.019212f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_378 N_D_c_395_n N_A_231_53#_c_1997_n 0.0018358f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_379 N_D_M1029_g N_A_404_53#_c_2028_n 0.00858539f $X=2.935 $Y=0.77 $X2=0 $Y2=0
cc_380 N_D_M1029_g N_A_404_53#_c_2030_n 0.00458834f $X=2.935 $Y=0.77 $X2=0 $Y2=0
cc_381 N_A_587_350#_c_455_n N_A_958_290#_M1021_d 5.6097e-19 $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_382 N_A_587_350#_c_455_n N_A_958_290#_M1033_g 0.00569996f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_383 N_A_587_350#_c_455_n N_A_958_290#_M1004_g 0.00387476f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_384 N_A_587_350#_c_455_n N_A_958_290#_c_654_n 0.0164094f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_385 N_A_587_350#_c_455_n N_A_958_290#_c_644_n 0.0108732f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_386 N_A_587_350#_c_455_n N_A_958_290#_c_645_n 0.22201f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_387 N_A_587_350#_c_455_n N_A_958_290#_c_656_n 0.023094f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_388 N_A_587_350#_c_455_n N_A_958_290#_c_646_n 0.0237183f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_389 N_A_587_350#_c_455_n N_A_958_290#_c_648_n 8.4675e-19 $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_390 N_A_587_350#_c_455_n N_A_958_290#_c_650_n 0.00177018f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_391 N_A_587_350#_c_455_n N_A_1067_65#_M1015_d 0.00218873f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_392 N_A_587_350#_c_455_n N_A_1067_65#_M1027_g 0.0105091f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_393 N_A_587_350#_M1016_g N_A_1067_65#_M1028_g 0.0126355f $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_394 N_A_587_350#_M1019_g N_A_1067_65#_M1009_g 0.0292916f $X=11.28 $Y=2.295
+ $X2=0 $Y2=0
cc_395 N_A_587_350#_c_436_n N_A_1067_65#_M1009_g 0.0070706f $X=11.355 $Y=1.67
+ $X2=0 $Y2=0
cc_396 N_A_587_350#_c_455_n N_A_1067_65#_M1009_g 0.00859438f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_397 N_A_587_350#_c_455_n N_A_1067_65#_c_788_n 0.0167178f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_398 N_A_587_350#_c_455_n N_A_1067_65#_c_798_n 0.0265013f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_399 N_A_587_350#_c_455_n N_A_1067_65#_c_802_n 0.0433646f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_400 N_A_587_350#_c_455_n N_A_1067_65#_c_803_n 0.0142355f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_401 N_A_587_350#_c_455_n N_A_1067_65#_c_804_n 0.0167926f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_402 N_A_587_350#_c_455_n N_A_1067_65#_c_823_n 0.0205044f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_403 N_A_587_350#_c_455_n N_A_1067_65#_c_806_n 0.0439573f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_404 N_A_587_350#_M1016_g N_A_1067_65#_c_790_n 0.00153696f $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_405 N_A_587_350#_M1016_g N_A_1067_65#_c_791_n 0.0114884f $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_406 N_A_587_350#_c_455_n N_A_1067_65#_c_791_n 0.00289105f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_407 N_A_587_350#_c_455_n N_A_1067_65#_c_794_n 0.0049331f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_408 N_A_587_350#_c_455_n N_A_902_396#_M1008_d 0.00116335f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_409 N_A_587_350#_c_455_n N_A_902_396#_M1015_g 0.0070675f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_410 N_A_587_350#_c_455_n N_A_902_396#_c_984_n 0.0172497f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_411 N_A_587_350#_c_455_n N_CLK_M1023_g 0.00614327f $X=12.095 $Y=2.035 $X2=0
+ $Y2=0
cc_412 N_A_587_350#_c_455_n N_A_872_324#_M1023_s 0.00201585f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_413 N_A_587_350#_c_455_n N_A_872_324#_M1008_g 0.00673877f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_414 N_A_587_350#_c_457_n N_A_872_324#_M1008_g 4.14098e-19 $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_415 N_A_587_350#_c_442_n N_A_872_324#_M1013_g 0.00236488f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_416 N_A_587_350#_c_455_n N_A_872_324#_M1021_g 0.00265443f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_417 N_A_587_350#_c_455_n N_A_872_324#_c_1109_n 0.00572224f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_418 N_A_587_350#_c_455_n N_A_872_324#_c_1127_n 0.00971387f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_419 N_A_587_350#_c_442_n N_A_872_324#_c_1111_n 0.00502855f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_420 N_A_587_350#_c_455_n N_A_872_324#_c_1111_n 0.00109795f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_421 N_A_587_350#_c_455_n N_A_872_324#_c_1131_n 0.0226245f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_422 N_A_587_350#_c_455_n N_A_872_324#_c_1118_n 0.00490897f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_423 N_A_587_350#_c_455_n N_A_872_324#_c_1120_n 0.00137775f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_424 N_A_587_350#_c_455_n N_A_1865_367#_M1030_d 0.00348341f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_425 N_A_587_350#_M1016_g N_A_1865_367#_c_1280_n 0.0185526f $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_426 N_A_587_350#_c_438_n N_A_1865_367#_c_1280_n 0.00499348f $X=12.025 $Y=0.98
+ $X2=0 $Y2=0
cc_427 N_A_587_350#_c_438_n N_A_1865_367#_c_1281_n 0.00786513f $X=12.025 $Y=0.98
+ $X2=0 $Y2=0
cc_428 N_A_587_350#_c_444_n N_A_1865_367#_c_1281_n 0.00975947f $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_429 N_A_587_350#_c_443_n N_A_1865_367#_c_1282_n 0.0152557f $X=11.73 $Y=1.67
+ $X2=0 $Y2=0
cc_430 N_A_587_350#_c_444_n N_A_1865_367#_c_1282_n 0.00150111f $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_431 N_A_587_350#_M1000_g N_A_1865_367#_c_1283_n 0.0179189f $X=12.83 $Y=0.705
+ $X2=0 $Y2=0
cc_432 N_A_587_350#_c_438_n N_A_1865_367#_c_1283_n 0.00865381f $X=12.025 $Y=0.98
+ $X2=0 $Y2=0
cc_433 N_A_587_350#_M1010_g N_A_1865_367#_M1034_g 0.0281169f $X=12.94 $Y=2.445
+ $X2=0 $Y2=0
cc_434 N_A_587_350#_c_439_n N_A_1865_367#_M1034_g 0.0102414f $X=12.85 $Y=1.49
+ $X2=0 $Y2=0
cc_435 N_A_587_350#_c_520_p N_A_1865_367#_M1034_g 0.00263219f $X=12.24 $Y=2.035
+ $X2=0 $Y2=0
cc_436 N_A_587_350#_c_443_n N_A_1865_367#_M1034_g 0.00681267f $X=11.73 $Y=1.67
+ $X2=0 $Y2=0
cc_437 N_A_587_350#_c_444_n N_A_1865_367#_M1034_g 0.0165224f $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_438 N_A_587_350#_M1000_g N_A_1865_367#_c_1287_n 0.00482387f $X=12.83 $Y=0.705
+ $X2=0 $Y2=0
cc_439 N_A_587_350#_c_438_n N_A_1865_367#_c_1287_n 0.001922f $X=12.025 $Y=0.98
+ $X2=0 $Y2=0
cc_440 N_A_587_350#_c_439_n N_A_1865_367#_c_1287_n 0.00335982f $X=12.85 $Y=1.49
+ $X2=0 $Y2=0
cc_441 N_A_587_350#_c_440_n N_A_1865_367#_c_1287_n 0.0213446f $X=12.85 $Y=1.49
+ $X2=0 $Y2=0
cc_442 N_A_587_350#_c_444_n N_A_1865_367#_c_1287_n 0.00947509f $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_443 N_A_587_350#_c_455_n N_A_1865_367#_c_1299_n 0.0206674f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_444 N_A_587_350#_M1019_g N_A_1865_367#_c_1300_n 0.00374811f $X=11.28 $Y=2.295
+ $X2=0 $Y2=0
cc_445 N_A_587_350#_c_455_n N_A_1865_367#_c_1300_n 0.0118741f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_446 N_A_587_350#_M1016_g N_A_1865_367#_c_1288_n 9.12839e-19 $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_447 N_A_587_350#_c_455_n N_A_1865_367#_c_1302_n 0.00835023f $X=12.095
+ $Y=2.035 $X2=0 $Y2=0
cc_448 N_A_587_350#_c_520_p N_A_1865_367#_c_1302_n 7.18054e-19 $X=12.24 $Y=2.035
+ $X2=0 $Y2=0
cc_449 N_A_587_350#_c_444_n N_A_1865_367#_c_1302_n 0.00560254f $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_450 N_A_587_350#_M1024_s N_A_1865_367#_c_1289_n 0.00137061f $X=11.89 $Y=0.705
+ $X2=0 $Y2=0
cc_451 N_A_587_350#_M1000_g N_A_1865_367#_c_1289_n 0.0160968f $X=12.83 $Y=0.705
+ $X2=0 $Y2=0
cc_452 N_A_587_350#_c_439_n N_A_1865_367#_c_1289_n 0.013704f $X=12.85 $Y=1.49
+ $X2=0 $Y2=0
cc_453 N_A_587_350#_c_440_n N_A_1865_367#_c_1289_n 9.37983e-19 $X=12.85 $Y=1.49
+ $X2=0 $Y2=0
cc_454 N_A_587_350#_c_444_n N_A_1865_367#_c_1289_n 0.00387689f $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_455 N_A_587_350#_M1010_g N_A_1865_367#_c_1303_n 0.00307078f $X=12.94 $Y=2.445
+ $X2=0 $Y2=0
cc_456 N_A_587_350#_M1010_g N_A_1865_367#_c_1304_n 0.0143654f $X=12.94 $Y=2.445
+ $X2=0 $Y2=0
cc_457 N_A_587_350#_M1034_s N_A_1865_367#_c_1305_n 0.0024164f $X=12.055 $Y=1.815
+ $X2=0 $Y2=0
cc_458 N_A_587_350#_c_520_p N_A_1865_367#_c_1305_n 0.00225291f $X=12.24 $Y=2.035
+ $X2=0 $Y2=0
cc_459 N_A_587_350#_c_444_n N_A_1865_367#_c_1305_n 0.00656127f $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_460 N_A_587_350#_M1000_g N_A_1865_367#_c_1290_n 0.00334104f $X=12.83 $Y=0.705
+ $X2=0 $Y2=0
cc_461 N_A_587_350#_M1010_g N_A_1865_367#_c_1290_n 0.00423519f $X=12.94 $Y=2.445
+ $X2=0 $Y2=0
cc_462 N_A_587_350#_M1016_g N_A_1865_367#_c_1293_n 0.00789042f $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_463 N_A_587_350#_M1019_g N_A_1865_367#_c_1307_n 0.0108902f $X=11.28 $Y=2.295
+ $X2=0 $Y2=0
cc_464 N_A_587_350#_c_455_n N_A_1865_367#_c_1307_n 9.28391e-19 $X=12.095
+ $Y=2.035 $X2=0 $Y2=0
cc_465 N_A_587_350#_M1016_g N_A_1865_367#_c_1294_n 0.0031575f $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_466 N_A_587_350#_M1024_s N_A_1865_367#_c_1295_n 8.19628e-19 $X=11.89 $Y=0.705
+ $X2=0 $Y2=0
cc_467 N_A_587_350#_M1016_g N_A_1865_367#_c_1295_n 5.17416e-19 $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_468 N_A_587_350#_c_438_n N_A_1865_367#_c_1295_n 0.0216217f $X=12.025 $Y=0.98
+ $X2=0 $Y2=0
cc_469 N_A_587_350#_M1000_g N_A_1865_367#_c_1296_n 0.00159804f $X=12.83 $Y=0.705
+ $X2=0 $Y2=0
cc_470 N_A_587_350#_c_440_n N_A_1865_367#_c_1296_n 0.00305588f $X=12.85 $Y=1.49
+ $X2=0 $Y2=0
cc_471 N_A_587_350#_c_455_n N_VPWR_M1027_d 0.00337103f $X=12.095 $Y=2.035 $X2=0
+ $Y2=0
cc_472 N_A_587_350#_c_455_n N_VPWR_M1009_d 0.00979196f $X=12.095 $Y=2.035 $X2=0
+ $Y2=0
cc_473 N_A_587_350#_c_455_n N_VPWR_c_1466_n 0.0174951f $X=12.095 $Y=2.035 $X2=0
+ $Y2=0
cc_474 N_A_587_350#_c_455_n N_VPWR_c_1467_n 0.00136648f $X=12.095 $Y=2.035 $X2=0
+ $Y2=0
cc_475 N_A_587_350#_M1010_g N_VPWR_c_1469_n 0.0138559f $X=12.94 $Y=2.445 $X2=0
+ $Y2=0
cc_476 N_A_587_350#_M1010_g N_VPWR_c_1470_n 0.00743142f $X=12.94 $Y=2.445 $X2=0
+ $Y2=0
cc_477 N_A_587_350#_M1003_g N_VPWR_c_1477_n 2.36211e-19 $X=3.01 $Y=2.325 $X2=0
+ $Y2=0
cc_478 N_A_587_350#_M1019_g N_VPWR_c_1478_n 6.84096e-19 $X=11.28 $Y=2.295 $X2=0
+ $Y2=0
cc_479 N_A_587_350#_M1010_g N_VPWR_c_1479_n 0.00469214f $X=12.94 $Y=2.445 $X2=0
+ $Y2=0
cc_480 N_A_587_350#_M1019_g N_VPWR_c_1462_n 4.45354e-19 $X=11.28 $Y=2.295 $X2=0
+ $Y2=0
cc_481 N_A_587_350#_M1010_g N_VPWR_c_1462_n 0.00566482f $X=12.94 $Y=2.445 $X2=0
+ $Y2=0
cc_482 N_A_587_350#_M1003_g N_A_286_423#_c_1606_n 0.00576606f $X=3.01 $Y=2.325
+ $X2=0 $Y2=0
cc_483 N_A_587_350#_M1003_g N_A_286_423#_c_1608_n 0.0110518f $X=3.01 $Y=2.325
+ $X2=0 $Y2=0
cc_484 N_A_587_350#_c_446_n N_A_286_423#_c_1608_n 0.00170987f $X=3.29 $Y=1.825
+ $X2=0 $Y2=0
cc_485 N_A_587_350#_c_456_n N_A_286_423#_c_1608_n 0.00168895f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_486 N_A_587_350#_c_457_n N_A_286_423#_c_1608_n 0.00345216f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_487 N_A_587_350#_M1003_g N_A_531_423#_c_1658_n 0.00278333f $X=3.01 $Y=2.325
+ $X2=0 $Y2=0
cc_488 N_A_587_350#_c_456_n N_A_531_423#_c_1658_n 0.00443662f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_489 N_A_587_350#_c_457_n N_A_531_423#_c_1658_n 0.00319744f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_490 N_A_587_350#_M1003_g N_A_531_423#_c_1659_n 0.00649069f $X=3.01 $Y=2.325
+ $X2=0 $Y2=0
cc_491 N_A_587_350#_c_446_n N_A_531_423#_c_1659_n 0.0100268f $X=3.29 $Y=1.825
+ $X2=0 $Y2=0
cc_492 N_A_587_350#_c_447_n N_A_531_423#_c_1659_n 0.00538562f $X=3.085 $Y=1.825
+ $X2=0 $Y2=0
cc_493 N_A_587_350#_c_441_n N_A_531_423#_c_1659_n 0.0126751f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_494 N_A_587_350#_c_442_n N_A_531_423#_c_1659_n 0.00297596f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_495 N_A_587_350#_M1017_g N_A_531_423#_c_1652_n 0.0141079f $X=3.365 $Y=0.77
+ $X2=0 $Y2=0
cc_496 N_A_587_350#_M1017_g N_A_531_423#_c_1653_n 0.00883697f $X=3.365 $Y=0.77
+ $X2=0 $Y2=0
cc_497 N_A_587_350#_c_441_n N_A_531_423#_c_1653_n 0.0200905f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_498 N_A_587_350#_c_442_n N_A_531_423#_c_1653_n 0.00843391f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_499 N_A_587_350#_M1017_g N_A_531_423#_c_1654_n 0.0148651f $X=3.365 $Y=0.77
+ $X2=0 $Y2=0
cc_500 N_A_587_350#_c_441_n N_A_531_423#_c_1654_n 0.0245697f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_501 N_A_587_350#_c_442_n N_A_531_423#_c_1654_n 0.00424181f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_502 N_A_587_350#_M1017_g N_A_531_423#_c_1655_n 0.00493497f $X=3.365 $Y=0.77
+ $X2=0 $Y2=0
cc_503 N_A_587_350#_c_441_n N_A_531_423#_c_1656_n 0.0132131f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_504 N_A_587_350#_c_442_n N_A_531_423#_c_1656_n 0.00395443f $X=3.655 $Y=1.615
+ $X2=0 $Y2=0
cc_505 N_A_587_350#_c_455_n N_A_531_423#_c_1656_n 0.0233684f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_506 N_A_587_350#_c_456_n N_A_531_423#_c_1656_n 9.70898e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_507 N_A_587_350#_c_457_n N_A_531_423#_c_1656_n 0.00516418f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_508 N_A_587_350#_c_455_n N_A_531_423#_c_1663_n 0.0119376f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_509 N_A_587_350#_c_455_n N_A_531_423#_c_1665_n 0.0306533f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_510 N_A_587_350#_c_455_n N_A_761_396#_M1008_s 0.00924249f $X=12.095 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_511 N_A_587_350#_c_455_n N_A_761_396#_c_1743_n 0.0214716f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_512 N_A_587_350#_c_456_n N_A_761_396#_c_1743_n 0.00152159f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_513 N_A_587_350#_c_457_n N_A_761_396#_c_1743_n 0.0122681f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_514 N_A_587_350#_c_455_n N_A_761_396#_c_1746_n 0.0115883f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_515 N_A_587_350#_c_455_n N_A_1781_367#_M1030_s 0.00340808f $X=12.095 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_516 N_A_587_350#_c_455_n N_A_1781_367#_M1009_s 0.00333504f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_517 N_A_587_350#_c_455_n N_A_1971_388#_M1004_d 0.00201864f $X=12.095 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_518 N_A_587_350#_M1019_g N_A_1971_388#_c_1799_n 0.0135623f $X=11.28 $Y=2.295
+ $X2=0 $Y2=0
cc_519 N_A_587_350#_c_435_n N_A_1971_388#_c_1799_n 0.00476826f $X=11.565 $Y=1.67
+ $X2=0 $Y2=0
cc_520 N_A_587_350#_c_436_n N_A_1971_388#_c_1799_n 0.00425361f $X=11.355 $Y=1.67
+ $X2=0 $Y2=0
cc_521 N_A_587_350#_c_455_n N_A_1971_388#_c_1799_n 0.0549751f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_522 N_A_587_350#_c_444_n N_A_1971_388#_c_1799_n 2.99177e-19 $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_523 N_A_587_350#_M1019_g N_A_1971_388#_c_1800_n 0.00750396f $X=11.28 $Y=2.295
+ $X2=0 $Y2=0
cc_524 N_A_587_350#_c_455_n N_A_1971_388#_c_1800_n 0.00718705f $X=12.095
+ $Y=2.035 $X2=0 $Y2=0
cc_525 N_A_587_350#_c_520_p N_A_1971_388#_c_1800_n 2.86915e-19 $X=12.24 $Y=2.035
+ $X2=0 $Y2=0
cc_526 N_A_587_350#_c_443_n N_A_1971_388#_c_1800_n 0.00559406f $X=11.73 $Y=1.67
+ $X2=0 $Y2=0
cc_527 N_A_587_350#_c_444_n N_A_1971_388#_c_1800_n 0.0204236f $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_528 N_A_587_350#_M1000_g N_Q_N_c_1827_n 0.00645152f $X=12.83 $Y=0.705 $X2=0
+ $Y2=0
cc_529 N_A_587_350#_c_439_n N_Q_N_c_1827_n 0.00954242f $X=12.85 $Y=1.49 $X2=0
+ $Y2=0
cc_530 N_A_587_350#_c_440_n N_Q_N_c_1827_n 0.00298368f $X=12.85 $Y=1.49 $X2=0
+ $Y2=0
cc_531 N_A_587_350#_M1000_g N_Q_N_c_1828_n 0.00409331f $X=12.83 $Y=0.705 $X2=0
+ $Y2=0
cc_532 N_A_587_350#_c_439_n N_Q_N_c_1828_n 0.0250968f $X=12.85 $Y=1.49 $X2=0
+ $Y2=0
cc_533 N_A_587_350#_c_440_n N_Q_N_c_1828_n 0.0106453f $X=12.85 $Y=1.49 $X2=0
+ $Y2=0
cc_534 N_A_587_350#_M1010_g N_Q_N_c_1836_n 0.0128168f $X=12.94 $Y=2.445 $X2=0
+ $Y2=0
cc_535 N_A_587_350#_c_439_n N_Q_N_c_1836_n 0.0278471f $X=12.85 $Y=1.49 $X2=0
+ $Y2=0
cc_536 N_A_587_350#_c_440_n N_Q_N_c_1836_n 0.00435527f $X=12.85 $Y=1.49 $X2=0
+ $Y2=0
cc_537 N_A_587_350#_c_520_p N_Q_N_c_1836_n 0.00646293f $X=12.24 $Y=2.035 $X2=0
+ $Y2=0
cc_538 N_A_587_350#_c_444_n N_Q_N_c_1836_n 0.0166545f $X=12.185 $Y=1.98 $X2=0
+ $Y2=0
cc_539 N_A_587_350#_M1000_g N_VGND_c_1874_n 0.00630741f $X=12.83 $Y=0.705 $X2=0
+ $Y2=0
cc_540 N_A_587_350#_M1016_g N_VGND_c_1875_n 4.7648e-19 $X=11.13 $Y=0.915 $X2=0
+ $Y2=0
cc_541 N_A_587_350#_M1000_g N_VGND_c_1876_n 0.00448732f $X=12.83 $Y=0.705 $X2=0
+ $Y2=0
cc_542 N_A_587_350#_M1000_g N_VGND_c_1877_n 0.00372834f $X=12.83 $Y=0.705 $X2=0
+ $Y2=0
cc_543 N_A_587_350#_M1017_g N_VGND_c_1879_n 6.24464e-19 $X=3.365 $Y=0.77 $X2=0
+ $Y2=0
cc_544 N_A_587_350#_M1000_g N_VGND_c_1882_n 0.00694202f $X=12.83 $Y=0.705 $X2=0
+ $Y2=0
cc_545 N_A_587_350#_M1017_g N_A_404_53#_c_2028_n 0.00665296f $X=3.365 $Y=0.77
+ $X2=0 $Y2=0
cc_546 N_A_587_350#_M1017_g N_A_404_53#_c_2029_n 0.0121066f $X=3.365 $Y=0.77
+ $X2=0 $Y2=0
cc_547 N_A_587_350#_M1016_g N_A_1789_141#_c_2050_n 0.00559654f $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_548 N_A_587_350#_c_436_n N_A_1789_141#_c_2050_n 0.00803165f $X=11.355 $Y=1.67
+ $X2=0 $Y2=0
cc_549 N_A_587_350#_c_438_n N_A_1789_141#_c_2050_n 0.0169705f $X=12.025 $Y=0.98
+ $X2=0 $Y2=0
cc_550 N_A_587_350#_c_443_n N_A_1789_141#_c_2050_n 3.43515e-19 $X=11.73 $Y=1.67
+ $X2=0 $Y2=0
cc_551 N_A_587_350#_c_444_n N_A_1789_141#_c_2050_n 0.00212142f $X=12.185 $Y=1.98
+ $X2=0 $Y2=0
cc_552 N_A_587_350#_M1016_g N_A_1789_141#_c_2056_n 0.018935f $X=11.13 $Y=0.915
+ $X2=0 $Y2=0
cc_553 N_A_587_350#_c_436_n N_A_1789_141#_c_2056_n 0.00185774f $X=11.355 $Y=1.67
+ $X2=0 $Y2=0
cc_554 N_A_958_290#_M1011_g N_A_1067_65#_M1014_g 0.0331672f $X=4.945 $Y=0.665
+ $X2=0 $Y2=0
cc_555 N_A_958_290#_M1011_g N_A_1067_65#_c_785_n 0.00731314f $X=4.945 $Y=0.665
+ $X2=0 $Y2=0
cc_556 N_A_958_290#_c_647_n N_A_1067_65#_c_785_n 0.0192688f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_557 N_A_958_290#_c_648_n N_A_1067_65#_c_785_n 0.00153963f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_558 N_A_958_290#_c_642_n N_A_1067_65#_M1028_g 0.00142274f $X=9.785 $Y=1.41
+ $X2=0 $Y2=0
cc_559 N_A_958_290#_c_643_n N_A_1067_65#_M1028_g 0.0175712f $X=9.785 $Y=1.41
+ $X2=0 $Y2=0
cc_560 N_A_958_290#_c_649_n N_A_1067_65#_M1028_g 0.0556546f $X=9.785 $Y=1.245
+ $X2=0 $Y2=0
cc_561 N_A_958_290#_M1033_g N_A_1067_65#_c_788_n 5.03415e-19 $X=4.865 $Y=2.19
+ $X2=0 $Y2=0
cc_562 N_A_958_290#_c_645_n N_A_1067_65#_c_788_n 0.0410489f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_563 N_A_958_290#_c_656_n N_A_1067_65#_c_788_n 5.58587e-19 $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_564 N_A_958_290#_c_647_n N_A_1067_65#_c_788_n 8.082e-19 $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_565 N_A_958_290#_c_648_n N_A_1067_65#_c_788_n 0.00923325f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_566 N_A_958_290#_c_654_n N_A_1067_65#_c_802_n 0.00834909f $X=8.505 $Y=2.145
+ $X2=0 $Y2=0
cc_567 N_A_958_290#_c_645_n N_A_1067_65#_c_802_n 0.0112965f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_568 N_A_958_290#_c_645_n N_A_1067_65#_c_803_n 0.00126206f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_569 N_A_958_290#_M1021_d N_A_1067_65#_c_804_n 0.00275315f $X=8.365 $Y=1.98
+ $X2=0 $Y2=0
cc_570 N_A_958_290#_c_654_n N_A_1067_65#_c_804_n 0.0184162f $X=8.505 $Y=2.145
+ $X2=0 $Y2=0
cc_571 N_A_958_290#_c_654_n N_A_1067_65#_c_823_n 0.0213904f $X=8.505 $Y=2.145
+ $X2=0 $Y2=0
cc_572 N_A_958_290#_M1004_g N_A_1067_65#_c_806_n 0.014081f $X=9.78 $Y=2.15 $X2=0
+ $Y2=0
cc_573 N_A_958_290#_c_643_n N_A_1067_65#_c_806_n 0.00440373f $X=9.785 $Y=1.41
+ $X2=0 $Y2=0
cc_574 N_A_958_290#_c_644_n N_A_1067_65#_c_806_n 0.0548094f $X=9.62 $Y=1.4 $X2=0
+ $Y2=0
cc_575 N_A_958_290#_c_644_n N_A_1067_65#_c_807_n 0.0131059f $X=9.62 $Y=1.4 $X2=0
+ $Y2=0
cc_576 N_A_958_290#_c_646_n N_A_1067_65#_c_807_n 2.93717e-19 $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_577 N_A_958_290#_c_650_n N_A_1067_65#_c_807_n 0.0099741f $X=8.477 $Y=1.47
+ $X2=0 $Y2=0
cc_578 N_A_958_290#_M1004_g N_A_1067_65#_c_790_n 0.00244859f $X=9.78 $Y=2.15
+ $X2=0 $Y2=0
cc_579 N_A_958_290#_c_642_n N_A_1067_65#_c_790_n 0.0125144f $X=9.785 $Y=1.41
+ $X2=0 $Y2=0
cc_580 N_A_958_290#_c_643_n N_A_1067_65#_c_790_n 4.13869e-19 $X=9.785 $Y=1.41
+ $X2=0 $Y2=0
cc_581 N_A_958_290#_M1004_g N_A_1067_65#_c_791_n 0.00419078f $X=9.78 $Y=2.15
+ $X2=0 $Y2=0
cc_582 N_A_958_290#_c_645_n N_A_1067_65#_c_793_n 0.023145f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_583 N_A_958_290#_M1033_g N_A_1067_65#_c_794_n 0.00260301f $X=4.865 $Y=2.19
+ $X2=0 $Y2=0
cc_584 N_A_958_290#_c_645_n N_A_1067_65#_c_794_n 0.00130835f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_585 N_A_958_290#_M1011_g N_A_902_396#_c_983_n 0.0148731f $X=4.945 $Y=0.665
+ $X2=0 $Y2=0
cc_586 N_A_958_290#_M1011_g N_A_902_396#_c_984_n 0.00449533f $X=4.945 $Y=0.665
+ $X2=0 $Y2=0
cc_587 N_A_958_290#_c_656_n N_A_902_396#_c_984_n 0.00642758f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_588 N_A_958_290#_c_647_n N_A_902_396#_c_984_n 0.00714797f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_589 N_A_958_290#_c_648_n N_A_902_396#_c_984_n 0.0207951f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_590 N_A_958_290#_M1011_g N_A_902_396#_c_985_n 0.0036341f $X=4.945 $Y=0.665
+ $X2=0 $Y2=0
cc_591 N_A_958_290#_c_647_n N_A_902_396#_c_985_n 0.00372758f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_592 N_A_958_290#_c_645_n N_A_902_396#_c_1000_n 0.0021863f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_593 N_A_958_290#_M1011_g N_A_902_396#_c_986_n 0.0116307f $X=4.945 $Y=0.665
+ $X2=0 $Y2=0
cc_594 N_A_958_290#_c_645_n N_A_902_396#_c_986_n 0.0134572f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_595 N_A_958_290#_c_656_n N_A_902_396#_c_986_n 0.00223745f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_596 N_A_958_290#_c_647_n N_A_902_396#_c_986_n 0.00151717f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_597 N_A_958_290#_c_648_n N_A_902_396#_c_986_n 0.0191806f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_598 N_A_958_290#_c_645_n N_CLK_c_1053_n 0.0026753f $X=8.255 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_599 N_A_958_290#_c_645_n N_CLK_c_1055_n 5.71356e-19 $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_600 N_A_958_290#_c_645_n N_CLK_c_1061_n 4.15227e-19 $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_601 N_A_958_290#_c_645_n CLK 0.0103455f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_602 N_A_958_290#_c_645_n N_CLK_c_1058_n 0.00798857f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_603 N_A_958_290#_c_647_n N_A_872_324#_M1008_g 0.0145878f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_604 N_A_958_290#_M1011_g N_A_872_324#_M1013_g 0.0248599f $X=4.945 $Y=0.665
+ $X2=0 $Y2=0
cc_605 N_A_958_290#_c_647_n N_A_872_324#_M1013_g 0.0152286f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_606 N_A_958_290#_M1033_g N_A_872_324#_c_1123_n 0.00211718f $X=4.865 $Y=2.19
+ $X2=0 $Y2=0
cc_607 N_A_958_290#_c_641_n N_A_872_324#_M1032_g 0.00782927f $X=8.375 $Y=0.69
+ $X2=0 $Y2=0
cc_608 N_A_958_290#_c_651_n N_A_872_324#_M1032_g 0.0103373f $X=8.477 $Y=1.385
+ $X2=0 $Y2=0
cc_609 N_A_958_290#_c_654_n N_A_872_324#_M1021_g 0.0085115f $X=8.505 $Y=2.145
+ $X2=0 $Y2=0
cc_610 N_A_958_290#_c_646_n N_A_872_324#_M1021_g 0.00147202f $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_611 N_A_958_290#_c_650_n N_A_872_324#_M1021_g 0.00234647f $X=8.477 $Y=1.47
+ $X2=0 $Y2=0
cc_612 N_A_958_290#_c_644_n N_A_872_324#_c_1109_n 0.0161458f $X=9.62 $Y=1.4
+ $X2=0 $Y2=0
cc_613 N_A_958_290#_c_650_n N_A_872_324#_c_1109_n 0.0231952f $X=8.477 $Y=1.47
+ $X2=0 $Y2=0
cc_614 N_A_958_290#_M1004_g N_A_872_324#_c_1127_n 0.0181897f $X=9.78 $Y=2.15
+ $X2=0 $Y2=0
cc_615 N_A_958_290#_c_654_n N_A_872_324#_c_1127_n 7.80089e-19 $X=8.505 $Y=2.145
+ $X2=0 $Y2=0
cc_616 N_A_958_290#_c_650_n N_A_872_324#_c_1127_n 0.00100665f $X=8.477 $Y=1.47
+ $X2=0 $Y2=0
cc_617 N_A_958_290#_c_641_n N_A_872_324#_M1020_g 0.00348688f $X=8.375 $Y=0.69
+ $X2=0 $Y2=0
cc_618 N_A_958_290#_c_642_n N_A_872_324#_M1020_g 9.02734e-19 $X=9.785 $Y=1.41
+ $X2=0 $Y2=0
cc_619 N_A_958_290#_c_643_n N_A_872_324#_M1020_g 0.0176121f $X=9.785 $Y=1.41
+ $X2=0 $Y2=0
cc_620 N_A_958_290#_c_644_n N_A_872_324#_M1020_g 0.0126309f $X=9.62 $Y=1.4 $X2=0
+ $Y2=0
cc_621 N_A_958_290#_c_649_n N_A_872_324#_M1020_g 0.0184761f $X=9.785 $Y=1.245
+ $X2=0 $Y2=0
cc_622 N_A_958_290#_c_650_n N_A_872_324#_M1020_g 8.71654e-19 $X=8.477 $Y=1.47
+ $X2=0 $Y2=0
cc_623 N_A_958_290#_c_651_n N_A_872_324#_M1020_g 0.00506239f $X=8.477 $Y=1.385
+ $X2=0 $Y2=0
cc_624 N_A_958_290#_c_645_n N_A_872_324#_c_1112_n 0.00761793f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_625 N_A_958_290#_c_646_n N_A_872_324#_c_1112_n 4.6293e-19 $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_626 N_A_958_290#_c_650_n N_A_872_324#_c_1112_n 0.00492348f $X=8.477 $Y=1.47
+ $X2=0 $Y2=0
cc_627 N_A_958_290#_c_646_n N_A_872_324#_c_1113_n 7.55481e-19 $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_628 N_A_958_290#_M1004_g N_A_872_324#_c_1114_n 0.00752949f $X=9.78 $Y=2.15
+ $X2=0 $Y2=0
cc_629 N_A_958_290#_c_645_n N_A_872_324#_c_1131_n 5.30708e-19 $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_630 N_A_958_290#_c_645_n N_A_872_324#_c_1116_n 0.00907554f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_631 N_A_958_290#_c_645_n N_A_872_324#_c_1117_n 0.00979834f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_632 N_A_958_290#_c_645_n N_A_872_324#_c_1118_n 0.019849f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_633 N_A_958_290#_c_645_n N_A_872_324#_c_1120_n 0.026932f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_634 N_A_958_290#_c_646_n N_A_872_324#_c_1120_n 0.0021298f $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_635 N_A_958_290#_c_651_n N_A_872_324#_c_1120_n 0.0478323f $X=8.477 $Y=1.385
+ $X2=0 $Y2=0
cc_636 N_A_958_290#_c_650_n N_A_872_324#_c_1121_n 0.0103373f $X=8.477 $Y=1.47
+ $X2=0 $Y2=0
cc_637 N_A_958_290#_M1004_g N_A_1865_367#_c_1299_n 0.00646144f $X=9.78 $Y=2.15
+ $X2=0 $Y2=0
cc_638 N_A_958_290#_M1004_g N_A_1865_367#_c_1300_n 0.00871135f $X=9.78 $Y=2.15
+ $X2=0 $Y2=0
cc_639 N_A_958_290#_c_649_n N_A_1865_367#_c_1291_n 0.00725155f $X=9.785 $Y=1.245
+ $X2=0 $Y2=0
cc_640 N_A_958_290#_c_649_n N_A_1865_367#_c_1292_n 0.00877168f $X=9.785 $Y=1.245
+ $X2=0 $Y2=0
cc_641 N_A_958_290#_M1033_g N_A_531_423#_c_1656_n 7.61817e-19 $X=4.865 $Y=2.19
+ $X2=0 $Y2=0
cc_642 N_A_958_290#_M1033_g N_A_531_423#_c_1663_n 0.00396687f $X=4.865 $Y=2.19
+ $X2=0 $Y2=0
cc_643 N_A_958_290#_M1033_g N_A_531_423#_c_1665_n 0.0109094f $X=4.865 $Y=2.19
+ $X2=0 $Y2=0
cc_644 N_A_958_290#_c_645_n N_A_531_423#_c_1665_n 2.50817e-19 $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_645 N_A_958_290#_c_656_n N_A_531_423#_c_1665_n 0.00121172f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_646 N_A_958_290#_c_647_n N_A_531_423#_c_1665_n 0.00238088f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_647 N_A_958_290#_c_648_n N_A_531_423#_c_1665_n 0.021804f $X=5.08 $Y=1.615
+ $X2=0 $Y2=0
cc_648 N_A_958_290#_M1033_g N_A_761_396#_c_1744_n 2.66192e-19 $X=4.865 $Y=2.19
+ $X2=0 $Y2=0
cc_649 N_A_958_290#_M1033_g N_A_761_396#_c_1746_n 7.59117e-19 $X=4.865 $Y=2.19
+ $X2=0 $Y2=0
cc_650 N_A_958_290#_M1004_g N_A_1781_367#_c_1777_n 7.66717e-19 $X=9.78 $Y=2.15
+ $X2=0 $Y2=0
cc_651 N_A_958_290#_M1004_g N_A_1971_388#_c_1799_n 0.00231324f $X=9.78 $Y=2.15
+ $X2=0 $Y2=0
cc_652 N_A_958_290#_M1011_g N_VGND_c_1870_n 0.00191638f $X=4.945 $Y=0.665 $X2=0
+ $Y2=0
cc_653 N_A_958_290#_c_641_n N_VGND_c_1871_n 0.0180055f $X=8.375 $Y=0.69 $X2=0
+ $Y2=0
cc_654 N_A_958_290#_c_641_n N_VGND_c_1873_n 0.00999358f $X=8.375 $Y=0.69 $X2=0
+ $Y2=0
cc_655 N_A_958_290#_c_649_n N_VGND_c_1873_n 0.00368186f $X=9.785 $Y=1.245 $X2=0
+ $Y2=0
cc_656 N_A_958_290#_M1011_g N_VGND_c_1879_n 0.00494808f $X=4.945 $Y=0.665 $X2=0
+ $Y2=0
cc_657 N_A_958_290#_M1011_g N_VGND_c_1882_n 0.00519032f $X=4.945 $Y=0.665 $X2=0
+ $Y2=0
cc_658 N_A_958_290#_c_641_n N_VGND_c_1882_n 0.0112197f $X=8.375 $Y=0.69 $X2=0
+ $Y2=0
cc_659 N_A_958_290#_c_649_n N_VGND_c_1882_n 0.00608439f $X=9.785 $Y=1.245 $X2=0
+ $Y2=0
cc_660 N_A_958_290#_c_641_n N_A_1789_141#_c_2049_n 0.0219659f $X=8.375 $Y=0.69
+ $X2=0 $Y2=0
cc_661 N_A_958_290#_c_644_n N_A_1789_141#_c_2049_n 0.0209177f $X=9.62 $Y=1.4
+ $X2=0 $Y2=0
cc_662 N_A_958_290#_c_649_n N_A_1789_141#_c_2049_n 0.0012171f $X=9.785 $Y=1.245
+ $X2=0 $Y2=0
cc_663 N_A_958_290#_c_642_n N_A_1789_141#_c_2056_n 0.0201555f $X=9.785 $Y=1.41
+ $X2=0 $Y2=0
cc_664 N_A_958_290#_c_643_n N_A_1789_141#_c_2056_n 0.00372735f $X=9.785 $Y=1.41
+ $X2=0 $Y2=0
cc_665 N_A_958_290#_c_644_n N_A_1789_141#_c_2056_n 0.0153055f $X=9.62 $Y=1.4
+ $X2=0 $Y2=0
cc_666 N_A_958_290#_c_649_n N_A_1789_141#_c_2056_n 0.0109961f $X=9.785 $Y=1.245
+ $X2=0 $Y2=0
cc_667 N_A_1067_65#_M1014_g N_A_902_396#_c_981_n 0.0115061f $X=5.41 $Y=0.665
+ $X2=0 $Y2=0
cc_668 N_A_1067_65#_c_789_n N_A_902_396#_c_981_n 0.00491856f $X=6.575 $Y=1.555
+ $X2=0 $Y2=0
cc_669 N_A_1067_65#_c_792_n N_A_902_396#_c_981_n 0.0112592f $X=6.575 $Y=0.535
+ $X2=0 $Y2=0
cc_670 N_A_1067_65#_c_785_n N_A_902_396#_M1015_g 0.00557668f $X=5.56 $Y=1.555
+ $X2=0 $Y2=0
cc_671 N_A_1067_65#_c_788_n N_A_902_396#_M1015_g 0.0158838f $X=6.41 $Y=1.72
+ $X2=0 $Y2=0
cc_672 N_A_1067_65#_c_798_n N_A_902_396#_M1015_g 0.0166172f $X=6.575 $Y=2.01
+ $X2=0 $Y2=0
cc_673 N_A_1067_65#_c_800_n N_A_902_396#_M1015_g 6.85188e-19 $X=6.66 $Y=2.905
+ $X2=0 $Y2=0
cc_674 N_A_1067_65#_c_793_n N_A_902_396#_M1015_g 0.00781599f $X=6.535 $Y=1.72
+ $X2=0 $Y2=0
cc_675 N_A_1067_65#_c_794_n N_A_902_396#_M1015_g 0.0289495f $X=5.825 $Y=1.72
+ $X2=0 $Y2=0
cc_676 N_A_1067_65#_M1014_g N_A_902_396#_c_983_n 0.00225357f $X=5.41 $Y=0.665
+ $X2=0 $Y2=0
cc_677 N_A_1067_65#_M1014_g N_A_902_396#_c_1000_n 3.94001e-19 $X=5.41 $Y=0.665
+ $X2=0 $Y2=0
cc_678 N_A_1067_65#_c_785_n N_A_902_396#_c_1000_n 4.10433e-19 $X=5.56 $Y=1.555
+ $X2=0 $Y2=0
cc_679 N_A_1067_65#_c_788_n N_A_902_396#_c_1000_n 0.0177462f $X=6.41 $Y=1.72
+ $X2=0 $Y2=0
cc_680 N_A_1067_65#_c_789_n N_A_902_396#_c_1000_n 0.0234506f $X=6.575 $Y=1.555
+ $X2=0 $Y2=0
cc_681 N_A_1067_65#_c_792_n N_A_902_396#_c_1000_n 0.0141731f $X=6.575 $Y=0.535
+ $X2=0 $Y2=0
cc_682 N_A_1067_65#_c_785_n N_A_902_396#_c_986_n 0.00421904f $X=5.56 $Y=1.555
+ $X2=0 $Y2=0
cc_683 N_A_1067_65#_c_787_n N_A_902_396#_c_986_n 0.0162383f $X=5.56 $Y=1.135
+ $X2=0 $Y2=0
cc_684 N_A_1067_65#_c_788_n N_A_902_396#_c_986_n 0.0181201f $X=6.41 $Y=1.72
+ $X2=0 $Y2=0
cc_685 N_A_1067_65#_c_794_n N_A_902_396#_c_986_n 0.00589322f $X=5.825 $Y=1.72
+ $X2=0 $Y2=0
cc_686 N_A_1067_65#_c_787_n N_A_902_396#_c_987_n 0.0100004f $X=5.56 $Y=1.135
+ $X2=0 $Y2=0
cc_687 N_A_1067_65#_c_788_n N_A_902_396#_c_987_n 0.0076472f $X=6.41 $Y=1.72
+ $X2=0 $Y2=0
cc_688 N_A_1067_65#_c_789_n N_A_902_396#_c_987_n 0.0132745f $X=6.575 $Y=1.555
+ $X2=0 $Y2=0
cc_689 N_A_1067_65#_c_792_n N_A_902_396#_c_987_n 0.0105008f $X=6.575 $Y=0.535
+ $X2=0 $Y2=0
cc_690 N_A_1067_65#_c_798_n N_CLK_M1023_g 0.0038055f $X=6.575 $Y=2.01 $X2=0
+ $Y2=0
cc_691 N_A_1067_65#_c_799_n N_CLK_M1023_g 0.00322857f $X=7.37 $Y=2.905 $X2=0
+ $Y2=0
cc_692 N_A_1067_65#_c_801_n N_CLK_M1023_g 0.0209582f $X=7.455 $Y=2.82 $X2=0
+ $Y2=0
cc_693 N_A_1067_65#_c_803_n N_CLK_M1023_g 0.00579311f $X=7.54 $Y=2.045 $X2=0
+ $Y2=0
cc_694 N_A_1067_65#_c_887_p N_CLK_M1023_g 9.66074e-19 $X=8.155 $Y=2.515 $X2=0
+ $Y2=0
cc_695 N_A_1067_65#_c_803_n N_CLK_c_1061_n 0.00430028f $X=7.54 $Y=2.045 $X2=0
+ $Y2=0
cc_696 N_A_1067_65#_c_793_n N_CLK_c_1061_n 6.5957e-19 $X=6.535 $Y=1.72 $X2=0
+ $Y2=0
cc_697 N_A_1067_65#_c_789_n CLK 0.0237223f $X=6.575 $Y=1.555 $X2=0 $Y2=0
cc_698 N_A_1067_65#_c_789_n N_CLK_c_1058_n 0.00115395f $X=6.575 $Y=1.555 $X2=0
+ $Y2=0
cc_699 N_A_1067_65#_M1027_g N_A_872_324#_c_1123_n 0.00879826f $X=5.825 $Y=2.495
+ $X2=0 $Y2=0
cc_700 N_A_1067_65#_c_799_n N_A_872_324#_c_1123_n 0.0177638f $X=7.37 $Y=2.905
+ $X2=0 $Y2=0
cc_701 N_A_1067_65#_c_800_n N_A_872_324#_c_1123_n 0.00557034f $X=6.66 $Y=2.905
+ $X2=0 $Y2=0
cc_702 N_A_1067_65#_c_805_n N_A_872_324#_c_1123_n 0.00105798f $X=8.24 $Y=2.6
+ $X2=0 $Y2=0
cc_703 N_A_1067_65#_c_801_n N_A_872_324#_M1021_g 0.00112716f $X=7.455 $Y=2.82
+ $X2=0 $Y2=0
cc_704 N_A_1067_65#_c_802_n N_A_872_324#_M1021_g 0.00591549f $X=8.07 $Y=2.045
+ $X2=0 $Y2=0
cc_705 N_A_1067_65#_c_887_p N_A_872_324#_M1021_g 0.0160705f $X=8.155 $Y=2.515
+ $X2=0 $Y2=0
cc_706 N_A_1067_65#_c_804_n N_A_872_324#_M1021_g 0.011385f $X=8.95 $Y=2.6 $X2=0
+ $Y2=0
cc_707 N_A_1067_65#_c_805_n N_A_872_324#_M1021_g 0.00391163f $X=8.24 $Y=2.6
+ $X2=0 $Y2=0
cc_708 N_A_1067_65#_c_823_n N_A_872_324#_M1021_g 0.00454626f $X=9.035 $Y=2.515
+ $X2=0 $Y2=0
cc_709 N_A_1067_65#_c_807_n N_A_872_324#_c_1109_n 0.00332551f $X=9.12 $Y=1.82
+ $X2=0 $Y2=0
cc_710 N_A_1067_65#_c_823_n N_A_872_324#_c_1127_n 0.0123373f $X=9.035 $Y=2.515
+ $X2=0 $Y2=0
cc_711 N_A_1067_65#_c_806_n N_A_872_324#_c_1127_n 0.0122759f $X=10.19 $Y=1.82
+ $X2=0 $Y2=0
cc_712 N_A_1067_65#_c_802_n N_A_872_324#_c_1112_n 0.00751605f $X=8.07 $Y=2.045
+ $X2=0 $Y2=0
cc_713 N_A_1067_65#_c_806_n N_A_872_324#_c_1114_n 0.00176086f $X=10.19 $Y=1.82
+ $X2=0 $Y2=0
cc_714 N_A_1067_65#_c_798_n N_A_872_324#_c_1131_n 0.0396791f $X=6.575 $Y=2.01
+ $X2=0 $Y2=0
cc_715 N_A_1067_65#_c_799_n N_A_872_324#_c_1131_n 0.0190301f $X=7.37 $Y=2.905
+ $X2=0 $Y2=0
cc_716 N_A_1067_65#_c_801_n N_A_872_324#_c_1131_n 0.0172052f $X=7.455 $Y=2.82
+ $X2=0 $Y2=0
cc_717 N_A_1067_65#_c_803_n N_A_872_324#_c_1131_n 0.00834909f $X=7.54 $Y=2.045
+ $X2=0 $Y2=0
cc_718 N_A_1067_65#_c_793_n N_A_872_324#_c_1131_n 0.00639112f $X=6.535 $Y=1.72
+ $X2=0 $Y2=0
cc_719 N_A_1067_65#_c_803_n N_A_872_324#_c_1118_n 0.00929286f $X=7.54 $Y=2.045
+ $X2=0 $Y2=0
cc_720 N_A_1067_65#_c_793_n N_A_872_324#_c_1118_n 0.00849742f $X=6.535 $Y=1.72
+ $X2=0 $Y2=0
cc_721 N_A_1067_65#_c_789_n N_A_872_324#_c_1119_n 0.00635775f $X=6.575 $Y=1.555
+ $X2=0 $Y2=0
cc_722 N_A_1067_65#_c_792_n N_A_872_324#_c_1119_n 0.0155047f $X=6.575 $Y=0.535
+ $X2=0 $Y2=0
cc_723 N_A_1067_65#_c_802_n N_A_872_324#_c_1120_n 0.0192812f $X=8.07 $Y=2.045
+ $X2=0 $Y2=0
cc_724 N_A_1067_65#_c_806_n N_A_1865_367#_M1030_d 0.00212484f $X=10.19 $Y=1.82
+ $X2=0 $Y2=0
cc_725 N_A_1067_65#_c_823_n N_A_1865_367#_c_1299_n 0.0127373f $X=9.035 $Y=2.515
+ $X2=0 $Y2=0
cc_726 N_A_1067_65#_c_806_n N_A_1865_367#_c_1299_n 0.0171928f $X=10.19 $Y=1.82
+ $X2=0 $Y2=0
cc_727 N_A_1067_65#_M1009_g N_A_1865_367#_c_1300_n 0.0145389f $X=10.74 $Y=2.465
+ $X2=0 $Y2=0
cc_728 N_A_1067_65#_c_806_n N_A_1865_367#_c_1300_n 0.00257747f $X=10.19 $Y=1.82
+ $X2=0 $Y2=0
cc_729 N_A_1067_65#_M1028_g N_A_1865_367#_c_1291_n 0.00125731f $X=10.265
+ $Y=0.705 $X2=0 $Y2=0
cc_730 N_A_1067_65#_M1028_g N_A_1865_367#_c_1292_n 0.0128277f $X=10.265 $Y=0.705
+ $X2=0 $Y2=0
cc_731 N_A_1067_65#_M1028_g N_A_1865_367#_c_1293_n 0.00488118f $X=10.265
+ $Y=0.705 $X2=0 $Y2=0
cc_732 N_A_1067_65#_M1009_g N_A_1865_367#_c_1307_n 0.00402206f $X=10.74 $Y=2.465
+ $X2=0 $Y2=0
cc_733 N_A_1067_65#_c_788_n N_VPWR_M1027_d 0.00217331f $X=6.41 $Y=1.72 $X2=0
+ $Y2=0
cc_734 N_A_1067_65#_c_801_n N_VPWR_M1023_d 0.00590291f $X=7.455 $Y=2.82 $X2=0
+ $Y2=0
cc_735 N_A_1067_65#_c_802_n N_VPWR_M1023_d 0.0193589f $X=8.07 $Y=2.045 $X2=0
+ $Y2=0
cc_736 N_A_1067_65#_c_887_p N_VPWR_M1023_d 0.00482776f $X=8.155 $Y=2.515 $X2=0
+ $Y2=0
cc_737 N_A_1067_65#_c_805_n N_VPWR_M1023_d 0.00110885f $X=8.24 $Y=2.6 $X2=0
+ $Y2=0
cc_738 N_A_1067_65#_M1027_g N_VPWR_c_1466_n 0.00998424f $X=5.825 $Y=2.495 $X2=0
+ $Y2=0
cc_739 N_A_1067_65#_c_788_n N_VPWR_c_1466_n 0.0156832f $X=6.41 $Y=1.72 $X2=0
+ $Y2=0
cc_740 N_A_1067_65#_c_798_n N_VPWR_c_1466_n 0.0307889f $X=6.575 $Y=2.01 $X2=0
+ $Y2=0
cc_741 N_A_1067_65#_c_800_n N_VPWR_c_1466_n 0.014091f $X=6.66 $Y=2.905 $X2=0
+ $Y2=0
cc_742 N_A_1067_65#_c_799_n N_VPWR_c_1467_n 0.0137879f $X=7.37 $Y=2.905 $X2=0
+ $Y2=0
cc_743 N_A_1067_65#_c_801_n N_VPWR_c_1467_n 0.0360082f $X=7.455 $Y=2.82 $X2=0
+ $Y2=0
cc_744 N_A_1067_65#_c_802_n N_VPWR_c_1467_n 0.0117089f $X=8.07 $Y=2.045 $X2=0
+ $Y2=0
cc_745 N_A_1067_65#_c_887_p N_VPWR_c_1467_n 0.0142355f $X=8.155 $Y=2.515 $X2=0
+ $Y2=0
cc_746 N_A_1067_65#_c_805_n N_VPWR_c_1467_n 0.0134566f $X=8.24 $Y=2.6 $X2=0
+ $Y2=0
cc_747 N_A_1067_65#_M1009_g N_VPWR_c_1468_n 0.00438959f $X=10.74 $Y=2.465 $X2=0
+ $Y2=0
cc_748 N_A_1067_65#_c_799_n N_VPWR_c_1473_n 0.0376646f $X=7.37 $Y=2.905 $X2=0
+ $Y2=0
cc_749 N_A_1067_65#_c_800_n N_VPWR_c_1473_n 0.0116114f $X=6.66 $Y=2.905 $X2=0
+ $Y2=0
cc_750 N_A_1067_65#_M1009_g N_VPWR_c_1475_n 0.00424871f $X=10.74 $Y=2.465 $X2=0
+ $Y2=0
cc_751 N_A_1067_65#_c_804_n N_VPWR_c_1475_n 0.0110037f $X=8.95 $Y=2.6 $X2=0
+ $Y2=0
cc_752 N_A_1067_65#_c_805_n N_VPWR_c_1475_n 0.00331292f $X=8.24 $Y=2.6 $X2=0
+ $Y2=0
cc_753 N_A_1067_65#_M1027_g N_VPWR_c_1462_n 7.94319e-19 $X=5.825 $Y=2.495 $X2=0
+ $Y2=0
cc_754 N_A_1067_65#_M1009_g N_VPWR_c_1462_n 0.00861229f $X=10.74 $Y=2.465 $X2=0
+ $Y2=0
cc_755 N_A_1067_65#_c_799_n N_VPWR_c_1462_n 0.028058f $X=7.37 $Y=2.905 $X2=0
+ $Y2=0
cc_756 N_A_1067_65#_c_800_n N_VPWR_c_1462_n 0.00828634f $X=6.66 $Y=2.905 $X2=0
+ $Y2=0
cc_757 N_A_1067_65#_c_804_n N_VPWR_c_1462_n 0.0173927f $X=8.95 $Y=2.6 $X2=0
+ $Y2=0
cc_758 N_A_1067_65#_c_805_n N_VPWR_c_1462_n 0.00440399f $X=8.24 $Y=2.6 $X2=0
+ $Y2=0
cc_759 N_A_1067_65#_M1027_g N_A_531_423#_c_1663_n 3.82952e-19 $X=5.825 $Y=2.495
+ $X2=0 $Y2=0
cc_760 N_A_1067_65#_M1027_g N_A_531_423#_c_1665_n 0.00703002f $X=5.825 $Y=2.495
+ $X2=0 $Y2=0
cc_761 N_A_1067_65#_M1027_g N_A_761_396#_c_1746_n 0.010677f $X=5.825 $Y=2.495
+ $X2=0 $Y2=0
cc_762 N_A_1067_65#_c_788_n N_A_761_396#_c_1746_n 0.0059837f $X=6.41 $Y=1.72
+ $X2=0 $Y2=0
cc_763 N_A_1067_65#_c_794_n N_A_761_396#_c_1746_n 0.00642633f $X=5.825 $Y=1.72
+ $X2=0 $Y2=0
cc_764 N_A_1067_65#_c_804_n N_A_1781_367#_M1030_s 0.0050287f $X=8.95 $Y=2.6
+ $X2=-0.19 $Y2=-0.245
cc_765 N_A_1067_65#_c_823_n N_A_1781_367#_M1030_s 0.0118888f $X=9.035 $Y=2.515
+ $X2=-0.19 $Y2=-0.245
cc_766 N_A_1067_65#_c_807_n N_A_1781_367#_M1030_s 0.00105069f $X=9.12 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_767 N_A_1067_65#_c_806_n N_A_1781_367#_M1009_s 0.00252745f $X=10.19 $Y=1.82
+ $X2=0 $Y2=0
cc_768 N_A_1067_65#_M1009_g N_A_1781_367#_c_1776_n 0.00360852f $X=10.74 $Y=2.465
+ $X2=0 $Y2=0
cc_769 N_A_1067_65#_c_804_n N_A_1781_367#_c_1777_n 0.017807f $X=8.95 $Y=2.6
+ $X2=0 $Y2=0
cc_770 N_A_1067_65#_M1009_g N_A_1971_388#_c_1799_n 0.014538f $X=10.74 $Y=2.465
+ $X2=0 $Y2=0
cc_771 N_A_1067_65#_c_806_n N_A_1971_388#_c_1799_n 0.0423301f $X=10.19 $Y=1.82
+ $X2=0 $Y2=0
cc_772 N_A_1067_65#_c_791_n N_A_1971_388#_c_1799_n 0.00415249f $X=10.355 $Y=1.51
+ $X2=0 $Y2=0
cc_773 N_A_1067_65#_M1014_g N_VGND_c_1870_n 0.0138896f $X=5.41 $Y=0.665 $X2=0
+ $Y2=0
cc_774 N_A_1067_65#_c_787_n N_VGND_c_1870_n 0.00413535f $X=5.56 $Y=1.135 $X2=0
+ $Y2=0
cc_775 N_A_1067_65#_c_792_n N_VGND_c_1870_n 0.0286067f $X=6.575 $Y=0.535 $X2=0
+ $Y2=0
cc_776 N_A_1067_65#_M1028_g N_VGND_c_1872_n 0.00650051f $X=10.265 $Y=0.705 $X2=0
+ $Y2=0
cc_777 N_A_1067_65#_M1028_g N_VGND_c_1873_n 0.00372834f $X=10.265 $Y=0.705 $X2=0
+ $Y2=0
cc_778 N_A_1067_65#_M1014_g N_VGND_c_1879_n 0.00429764f $X=5.41 $Y=0.665 $X2=0
+ $Y2=0
cc_779 N_A_1067_65#_c_792_n N_VGND_c_1880_n 0.0356346f $X=6.575 $Y=0.535 $X2=0
+ $Y2=0
cc_780 N_A_1067_65#_M1035_d N_VGND_c_1882_n 0.00233022f $X=6.11 $Y=0.235 $X2=0
+ $Y2=0
cc_781 N_A_1067_65#_M1014_g N_VGND_c_1882_n 0.00435987f $X=5.41 $Y=0.665 $X2=0
+ $Y2=0
cc_782 N_A_1067_65#_M1028_g N_VGND_c_1882_n 0.00612119f $X=10.265 $Y=0.705 $X2=0
+ $Y2=0
cc_783 N_A_1067_65#_c_792_n N_VGND_c_1882_n 0.0219827f $X=6.575 $Y=0.535 $X2=0
+ $Y2=0
cc_784 N_A_1067_65#_M1028_g N_A_1789_141#_c_2056_n 0.012489f $X=10.265 $Y=0.705
+ $X2=0 $Y2=0
cc_785 N_A_1067_65#_c_806_n N_A_1789_141#_c_2056_n 0.00533944f $X=10.19 $Y=1.82
+ $X2=0 $Y2=0
cc_786 N_A_1067_65#_c_790_n N_A_1789_141#_c_2056_n 0.0154619f $X=10.355 $Y=1.51
+ $X2=0 $Y2=0
cc_787 N_A_1067_65#_c_791_n N_A_1789_141#_c_2056_n 0.00922349f $X=10.355 $Y=1.51
+ $X2=0 $Y2=0
cc_788 N_A_902_396#_c_987_n N_CLK_c_1058_n 0.00826696f $X=6.36 $Y=1.15 $X2=0
+ $Y2=0
cc_789 N_A_902_396#_c_984_n N_A_872_324#_M1008_g 0.00167535f $X=4.65 $Y=2.16
+ $X2=0 $Y2=0
cc_790 N_A_902_396#_c_983_n N_A_872_324#_M1013_g 0.00209069f $X=4.73 $Y=0.665
+ $X2=0 $Y2=0
cc_791 N_A_902_396#_c_984_n N_A_872_324#_M1013_g 0.00403091f $X=4.65 $Y=2.16
+ $X2=0 $Y2=0
cc_792 N_A_902_396#_c_985_n N_A_872_324#_M1013_g 0.00162548f $X=4.73 $Y=1.16
+ $X2=0 $Y2=0
cc_793 N_A_902_396#_M1015_g N_A_872_324#_c_1123_n 0.00879951f $X=6.36 $Y=2.285
+ $X2=0 $Y2=0
cc_794 N_A_902_396#_M1015_g N_A_872_324#_c_1131_n 0.0022126f $X=6.36 $Y=2.285
+ $X2=0 $Y2=0
cc_795 N_A_902_396#_M1015_g N_A_872_324#_c_1118_n 6.64198e-19 $X=6.36 $Y=2.285
+ $X2=0 $Y2=0
cc_796 N_A_902_396#_M1015_g N_VPWR_c_1466_n 0.00253761f $X=6.36 $Y=2.285 $X2=0
+ $Y2=0
cc_797 N_A_902_396#_M1015_g N_VPWR_c_1462_n 7.91655e-19 $X=6.36 $Y=2.285 $X2=0
+ $Y2=0
cc_798 N_A_902_396#_c_983_n N_A_531_423#_c_1655_n 0.0173815f $X=4.73 $Y=0.665
+ $X2=0 $Y2=0
cc_799 N_A_902_396#_c_985_n N_A_531_423#_c_1655_n 0.00208181f $X=4.73 $Y=1.16
+ $X2=0 $Y2=0
cc_800 N_A_902_396#_c_984_n N_A_531_423#_c_1656_n 0.0634971f $X=4.65 $Y=2.16
+ $X2=0 $Y2=0
cc_801 N_A_902_396#_c_984_n N_A_531_423#_c_1663_n 0.0126352f $X=4.65 $Y=2.16
+ $X2=0 $Y2=0
cc_802 N_A_902_396#_c_984_n N_A_531_423#_c_1665_n 0.0165303f $X=4.65 $Y=2.16
+ $X2=0 $Y2=0
cc_803 N_A_902_396#_c_984_n N_A_531_423#_c_1657_n 0.00198967f $X=4.65 $Y=2.16
+ $X2=0 $Y2=0
cc_804 N_A_902_396#_c_985_n N_A_531_423#_c_1657_n 0.0130324f $X=4.73 $Y=1.16
+ $X2=0 $Y2=0
cc_805 N_A_902_396#_c_981_n N_VGND_c_1870_n 0.0128311f $X=6.035 $Y=0.985 $X2=0
+ $Y2=0
cc_806 N_A_902_396#_c_983_n N_VGND_c_1870_n 0.0128446f $X=4.73 $Y=0.665 $X2=0
+ $Y2=0
cc_807 N_A_902_396#_c_986_n N_VGND_c_1870_n 0.02583f $X=5.97 $Y=1.15 $X2=0 $Y2=0
cc_808 N_A_902_396#_c_983_n N_VGND_c_1879_n 0.010825f $X=4.73 $Y=0.665 $X2=0
+ $Y2=0
cc_809 N_A_902_396#_c_981_n N_VGND_c_1880_n 0.00547815f $X=6.035 $Y=0.985 $X2=0
+ $Y2=0
cc_810 N_A_902_396#_c_981_n N_VGND_c_1882_n 0.012854f $X=6.035 $Y=0.985 $X2=0
+ $Y2=0
cc_811 N_A_902_396#_c_983_n N_VGND_c_1882_n 0.0114514f $X=4.73 $Y=0.665 $X2=0
+ $Y2=0
cc_812 N_CLK_M1023_g N_A_872_324#_c_1123_n 0.00483219f $X=7.32 $Y=2.3 $X2=0
+ $Y2=0
cc_813 N_CLK_M1018_g N_A_872_324#_M1032_g 0.0111171f $X=7.46 $Y=0.69 $X2=0 $Y2=0
cc_814 N_CLK_c_1061_n N_A_872_324#_c_1112_n 0.012058f $X=7.46 $Y=1.745 $X2=0
+ $Y2=0
cc_815 N_CLK_c_1055_n N_A_872_324#_c_1113_n 0.012058f $X=7.46 $Y=1.67 $X2=0
+ $Y2=0
cc_816 N_CLK_c_1061_n N_A_872_324#_c_1131_n 0.00842279f $X=7.46 $Y=1.745 $X2=0
+ $Y2=0
cc_817 N_CLK_M1018_g N_A_872_324#_c_1115_n 0.00777802f $X=7.46 $Y=0.69 $X2=0
+ $Y2=0
cc_818 N_CLK_c_1055_n N_A_872_324#_c_1116_n 0.00948295f $X=7.46 $Y=1.67 $X2=0
+ $Y2=0
cc_819 CLK N_A_872_324#_c_1116_n 0.0114632f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_820 N_CLK_c_1058_n N_A_872_324#_c_1116_n 4.71756e-19 $X=7.005 $Y=1.175 $X2=0
+ $Y2=0
cc_821 N_CLK_c_1055_n N_A_872_324#_c_1117_n 4.52736e-19 $X=7.46 $Y=1.67 $X2=0
+ $Y2=0
cc_822 N_CLK_c_1056_n N_A_872_324#_c_1117_n 0.00236916f $X=7.46 $Y=1.175 $X2=0
+ $Y2=0
cc_823 N_CLK_c_1053_n N_A_872_324#_c_1118_n 0.00316666f $X=7.385 $Y=1.175 $X2=0
+ $Y2=0
cc_824 N_CLK_c_1055_n N_A_872_324#_c_1118_n 0.00215255f $X=7.46 $Y=1.67 $X2=0
+ $Y2=0
cc_825 N_CLK_c_1061_n N_A_872_324#_c_1118_n 0.00995163f $X=7.46 $Y=1.745 $X2=0
+ $Y2=0
cc_826 CLK N_A_872_324#_c_1118_n 0.014181f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_827 N_CLK_c_1058_n N_A_872_324#_c_1118_n 0.00500971f $X=7.005 $Y=1.175 $X2=0
+ $Y2=0
cc_828 N_CLK_M1018_g N_A_872_324#_c_1119_n 0.0152091f $X=7.46 $Y=0.69 $X2=0
+ $Y2=0
cc_829 CLK N_A_872_324#_c_1119_n 0.0157909f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_830 N_CLK_c_1058_n N_A_872_324#_c_1119_n 0.0111926f $X=7.005 $Y=1.175 $X2=0
+ $Y2=0
cc_831 N_CLK_c_1053_n N_A_872_324#_c_1231_n 0.00385352f $X=7.385 $Y=1.175 $X2=0
+ $Y2=0
cc_832 N_CLK_c_1055_n N_A_872_324#_c_1231_n 2.88146e-19 $X=7.46 $Y=1.67 $X2=0
+ $Y2=0
cc_833 N_CLK_c_1056_n N_A_872_324#_c_1231_n 0.00190683f $X=7.46 $Y=1.175 $X2=0
+ $Y2=0
cc_834 CLK N_A_872_324#_c_1231_n 0.013037f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_835 N_CLK_c_1055_n N_A_872_324#_c_1120_n 0.00166089f $X=7.46 $Y=1.67 $X2=0
+ $Y2=0
cc_836 N_CLK_c_1056_n N_A_872_324#_c_1121_n 0.012058f $X=7.46 $Y=1.175 $X2=0
+ $Y2=0
cc_837 N_CLK_M1023_g N_VPWR_c_1467_n 0.00219462f $X=7.32 $Y=2.3 $X2=0 $Y2=0
cc_838 N_CLK_M1018_g N_VGND_c_1871_n 0.00890308f $X=7.46 $Y=0.69 $X2=0 $Y2=0
cc_839 N_CLK_M1018_g N_VGND_c_1880_n 0.00404051f $X=7.46 $Y=0.69 $X2=0 $Y2=0
cc_840 N_CLK_M1018_g N_VGND_c_1882_n 0.00511399f $X=7.46 $Y=0.69 $X2=0 $Y2=0
cc_841 N_A_872_324#_c_1127_n N_A_1865_367#_c_1299_n 0.00524051f $X=9.25 $Y=1.725
+ $X2=0 $Y2=0
cc_842 N_A_872_324#_c_1127_n N_A_1865_367#_c_1301_n 0.00531474f $X=9.25 $Y=1.725
+ $X2=0 $Y2=0
cc_843 N_A_872_324#_M1020_g N_A_1865_367#_c_1291_n 0.00329957f $X=9.305 $Y=0.915
+ $X2=0 $Y2=0
cc_844 N_A_872_324#_c_1123_n N_VPWR_c_1466_n 0.0216291f $X=8.215 $Y=3.15 $X2=0
+ $Y2=0
cc_845 N_A_872_324#_c_1123_n N_VPWR_c_1467_n 0.0168923f $X=8.215 $Y=3.15 $X2=0
+ $Y2=0
cc_846 N_A_872_324#_M1021_g N_VPWR_c_1467_n 0.0105866f $X=8.29 $Y=2.3 $X2=0
+ $Y2=0
cc_847 N_A_872_324#_c_1123_n N_VPWR_c_1473_n 0.0367066f $X=8.215 $Y=3.15 $X2=0
+ $Y2=0
cc_848 N_A_872_324#_c_1123_n N_VPWR_c_1475_n 0.0144972f $X=8.215 $Y=3.15 $X2=0
+ $Y2=0
cc_849 N_A_872_324#_c_1127_n N_VPWR_c_1475_n 0.00359964f $X=9.25 $Y=1.725 $X2=0
+ $Y2=0
cc_850 N_A_872_324#_c_1124_n N_VPWR_c_1477_n 0.0367702f $X=4.51 $Y=3.15 $X2=0
+ $Y2=0
cc_851 N_A_872_324#_c_1123_n N_VPWR_c_1462_n 0.101233f $X=8.215 $Y=3.15 $X2=0
+ $Y2=0
cc_852 N_A_872_324#_c_1124_n N_VPWR_c_1462_n 0.00604685f $X=4.51 $Y=3.15 $X2=0
+ $Y2=0
cc_853 N_A_872_324#_c_1127_n N_VPWR_c_1462_n 0.00805223f $X=9.25 $Y=1.725 $X2=0
+ $Y2=0
cc_854 N_A_872_324#_M1013_g N_A_531_423#_c_1655_n 0.00640399f $X=4.475 $Y=0.665
+ $X2=0 $Y2=0
cc_855 N_A_872_324#_M1008_g N_A_531_423#_c_1656_n 0.0215457f $X=4.435 $Y=2.19
+ $X2=0 $Y2=0
cc_856 N_A_872_324#_M1013_g N_A_531_423#_c_1656_n 0.00612348f $X=4.475 $Y=0.665
+ $X2=0 $Y2=0
cc_857 N_A_872_324#_c_1111_n N_A_531_423#_c_1656_n 0.00409437f $X=4.455 $Y=1.77
+ $X2=0 $Y2=0
cc_858 N_A_872_324#_M1008_g N_A_531_423#_c_1663_n 0.0103167f $X=4.435 $Y=2.19
+ $X2=0 $Y2=0
cc_859 N_A_872_324#_M1008_g N_A_531_423#_c_1664_n 0.00368691f $X=4.435 $Y=2.19
+ $X2=0 $Y2=0
cc_860 N_A_872_324#_M1008_g N_A_531_423#_c_1665_n 9.22276e-19 $X=4.435 $Y=2.19
+ $X2=0 $Y2=0
cc_861 N_A_872_324#_M1013_g N_A_531_423#_c_1657_n 0.00415728f $X=4.475 $Y=0.665
+ $X2=0 $Y2=0
cc_862 N_A_872_324#_M1008_g N_A_761_396#_c_1743_n 0.00891401f $X=4.435 $Y=2.19
+ $X2=0 $Y2=0
cc_863 N_A_872_324#_M1008_g N_A_761_396#_c_1744_n 0.0136556f $X=4.435 $Y=2.19
+ $X2=0 $Y2=0
cc_864 N_A_872_324#_c_1123_n N_A_761_396#_c_1744_n 0.0256411f $X=8.215 $Y=3.15
+ $X2=0 $Y2=0
cc_865 N_A_872_324#_M1021_g N_A_1781_367#_c_1777_n 0.00613377f $X=8.29 $Y=2.3
+ $X2=0 $Y2=0
cc_866 N_A_872_324#_c_1127_n N_A_1781_367#_c_1777_n 0.0148413f $X=9.25 $Y=1.725
+ $X2=0 $Y2=0
cc_867 N_A_872_324#_M1032_g N_VGND_c_1871_n 0.00685995f $X=8.16 $Y=0.69 $X2=0
+ $Y2=0
cc_868 N_A_872_324#_c_1117_n N_VGND_c_1871_n 0.00596548f $X=7.775 $Y=1.185 $X2=0
+ $Y2=0
cc_869 N_A_872_324#_c_1119_n N_VGND_c_1871_n 0.0221168f $X=7.13 $Y=0.69 $X2=0
+ $Y2=0
cc_870 N_A_872_324#_c_1120_n N_VGND_c_1871_n 0.0216591f $X=7.94 $Y=1.265 $X2=0
+ $Y2=0
cc_871 N_A_872_324#_c_1121_n N_VGND_c_1871_n 0.00197431f $X=7.94 $Y=1.265 $X2=0
+ $Y2=0
cc_872 N_A_872_324#_M1032_g N_VGND_c_1873_n 0.00479399f $X=8.16 $Y=0.69 $X2=0
+ $Y2=0
cc_873 N_A_872_324#_M1020_g N_VGND_c_1873_n 0.00362015f $X=9.305 $Y=0.915 $X2=0
+ $Y2=0
cc_874 N_A_872_324#_M1013_g N_VGND_c_1879_n 0.00517164f $X=4.475 $Y=0.665 $X2=0
+ $Y2=0
cc_875 N_A_872_324#_c_1119_n N_VGND_c_1880_n 0.0103911f $X=7.13 $Y=0.69 $X2=0
+ $Y2=0
cc_876 N_A_872_324#_M1013_g N_VGND_c_1882_n 0.00519032f $X=4.475 $Y=0.665 $X2=0
+ $Y2=0
cc_877 N_A_872_324#_M1032_g N_VGND_c_1882_n 0.00511399f $X=8.16 $Y=0.69 $X2=0
+ $Y2=0
cc_878 N_A_872_324#_M1020_g N_VGND_c_1882_n 0.00447875f $X=9.305 $Y=0.915 $X2=0
+ $Y2=0
cc_879 N_A_872_324#_c_1119_n N_VGND_c_1882_n 0.0164735f $X=7.13 $Y=0.69 $X2=0
+ $Y2=0
cc_880 N_A_872_324#_M1013_g N_A_404_53#_c_2028_n 0.00296645f $X=4.475 $Y=0.665
+ $X2=0 $Y2=0
cc_881 N_A_872_324#_M1032_g N_A_1789_141#_c_2049_n 5.76812e-19 $X=8.16 $Y=0.69
+ $X2=0 $Y2=0
cc_882 N_A_872_324#_M1020_g N_A_1789_141#_c_2049_n 0.00817419f $X=9.305 $Y=0.915
+ $X2=0 $Y2=0
cc_883 N_A_872_324#_M1020_g N_A_1789_141#_c_2056_n 0.0100043f $X=9.305 $Y=0.915
+ $X2=0 $Y2=0
cc_884 N_A_1865_367#_c_1300_n N_VPWR_M1009_d 0.00589424f $X=11.22 $Y=2.52 $X2=0
+ $Y2=0
cc_885 N_A_1865_367#_c_1304_n N_VPWR_M1034_d 0.00757803f $X=13.54 $Y=2.43 $X2=0
+ $Y2=0
cc_886 N_A_1865_367#_c_1304_n N_VPWR_M1031_s 0.00342855f $X=13.54 $Y=2.43 $X2=0
+ $Y2=0
cc_887 N_A_1865_367#_c_1290_n N_VPWR_M1031_s 0.00281733f $X=13.705 $Y=1.35 $X2=0
+ $Y2=0
cc_888 N_A_1865_367#_c_1300_n N_VPWR_c_1468_n 0.0124328f $X=11.22 $Y=2.52 $X2=0
+ $Y2=0
cc_889 N_A_1865_367#_c_1307_n N_VPWR_c_1468_n 0.00638707f $X=11.305 $Y=2.52
+ $X2=0 $Y2=0
cc_890 N_A_1865_367#_c_1302_n N_VPWR_c_1469_n 0.0144409f $X=12.21 $Y=2.79 $X2=0
+ $Y2=0
cc_891 N_A_1865_367#_c_1303_n N_VPWR_c_1469_n 7.25377e-19 $X=12.295 $Y=2.705
+ $X2=0 $Y2=0
cc_892 N_A_1865_367#_c_1304_n N_VPWR_c_1469_n 0.0205787f $X=13.54 $Y=2.43 $X2=0
+ $Y2=0
cc_893 N_A_1865_367#_M1031_g N_VPWR_c_1470_n 0.011548f $X=13.92 $Y=2.465 $X2=0
+ $Y2=0
cc_894 N_A_1865_367#_c_1304_n N_VPWR_c_1470_n 0.0223762f $X=13.54 $Y=2.43 $X2=0
+ $Y2=0
cc_895 N_A_1865_367#_c_1300_n N_VPWR_c_1475_n 0.00208901f $X=11.22 $Y=2.52 $X2=0
+ $Y2=0
cc_896 N_A_1865_367#_M1034_g N_VPWR_c_1478_n 0.00209575f $X=12.4 $Y=2.135 $X2=0
+ $Y2=0
cc_897 N_A_1865_367#_c_1300_n N_VPWR_c_1478_n 0.00265985f $X=11.22 $Y=2.52 $X2=0
+ $Y2=0
cc_898 N_A_1865_367#_c_1302_n N_VPWR_c_1478_n 0.0284513f $X=12.21 $Y=2.79 $X2=0
+ $Y2=0
cc_899 N_A_1865_367#_c_1307_n N_VPWR_c_1478_n 0.00509529f $X=11.305 $Y=2.52
+ $X2=0 $Y2=0
cc_900 N_A_1865_367#_M1031_g N_VPWR_c_1480_n 0.00486043f $X=13.92 $Y=2.465 $X2=0
+ $Y2=0
cc_901 N_A_1865_367#_M1030_d N_VPWR_c_1462_n 0.00220439f $X=9.325 $Y=1.835 $X2=0
+ $Y2=0
cc_902 N_A_1865_367#_M1034_g N_VPWR_c_1462_n 0.00258272f $X=12.4 $Y=2.135 $X2=0
+ $Y2=0
cc_903 N_A_1865_367#_M1031_g N_VPWR_c_1462_n 0.00918457f $X=13.92 $Y=2.465 $X2=0
+ $Y2=0
cc_904 N_A_1865_367#_c_1300_n N_VPWR_c_1462_n 0.0120167f $X=11.22 $Y=2.52 $X2=0
+ $Y2=0
cc_905 N_A_1865_367#_c_1302_n N_VPWR_c_1462_n 0.0326909f $X=12.21 $Y=2.79 $X2=0
+ $Y2=0
cc_906 N_A_1865_367#_c_1304_n N_VPWR_c_1462_n 0.0304888f $X=13.54 $Y=2.43 $X2=0
+ $Y2=0
cc_907 N_A_1865_367#_c_1307_n N_VPWR_c_1462_n 0.00570094f $X=11.305 $Y=2.52
+ $X2=0 $Y2=0
cc_908 N_A_1865_367#_c_1300_n N_A_1781_367#_M1009_s 0.00530448f $X=11.22 $Y=2.52
+ $X2=0 $Y2=0
cc_909 N_A_1865_367#_c_1300_n N_A_1781_367#_c_1776_n 0.01885f $X=11.22 $Y=2.52
+ $X2=0 $Y2=0
cc_910 N_A_1865_367#_M1030_d N_A_1781_367#_c_1777_n 0.00537218f $X=9.325
+ $Y=1.835 $X2=0 $Y2=0
cc_911 N_A_1865_367#_c_1300_n N_A_1781_367#_c_1777_n 0.0375904f $X=11.22 $Y=2.52
+ $X2=0 $Y2=0
cc_912 N_A_1865_367#_c_1301_n N_A_1781_367#_c_1777_n 0.0199827f $X=9.63 $Y=2.52
+ $X2=0 $Y2=0
cc_913 N_A_1865_367#_c_1299_n N_A_1971_388#_c_1799_n 0.0119097f $X=9.465
+ $Y=2.435 $X2=0 $Y2=0
cc_914 N_A_1865_367#_c_1300_n N_A_1971_388#_c_1799_n 0.0770089f $X=11.22 $Y=2.52
+ $X2=0 $Y2=0
cc_915 N_A_1865_367#_c_1302_n N_A_1971_388#_c_1799_n 0.0051604f $X=12.21 $Y=2.79
+ $X2=0 $Y2=0
cc_916 N_A_1865_367#_c_1307_n N_A_1971_388#_c_1799_n 0.00869797f $X=11.305
+ $Y=2.52 $X2=0 $Y2=0
cc_917 N_A_1865_367#_M1034_g N_A_1971_388#_c_1800_n 0.0053441f $X=12.4 $Y=2.135
+ $X2=0 $Y2=0
cc_918 N_A_1865_367#_c_1302_n N_A_1971_388#_c_1800_n 0.0182161f $X=12.21 $Y=2.79
+ $X2=0 $Y2=0
cc_919 N_A_1865_367#_c_1303_n N_A_1971_388#_c_1800_n 4.15802e-19 $X=12.295
+ $Y=2.705 $X2=0 $Y2=0
cc_920 N_A_1865_367#_c_1305_n N_A_1971_388#_c_1800_n 0.00807641f $X=12.38
+ $Y=2.43 $X2=0 $Y2=0
cc_921 N_A_1865_367#_c_1307_n N_A_1971_388#_c_1800_n 0.00403492f $X=11.305
+ $Y=2.52 $X2=0 $Y2=0
cc_922 N_A_1865_367#_c_1289_n N_Q_N_M1000_d 0.00660287f $X=13.54 $Y=0.63
+ $X2=-0.19 $Y2=-0.245
cc_923 N_A_1865_367#_c_1304_n N_Q_N_M1010_d 0.00773754f $X=13.54 $Y=2.43 $X2=0
+ $Y2=0
cc_924 N_A_1865_367#_c_1283_n N_Q_N_c_1827_n 0.00111676f $X=12.24 $Y=1.235 $X2=0
+ $Y2=0
cc_925 N_A_1865_367#_c_1285_n N_Q_N_c_1827_n 0.0010157f $X=13.915 $Y=1.185 $X2=0
+ $Y2=0
cc_926 N_A_1865_367#_c_1289_n N_Q_N_c_1827_n 0.0317548f $X=13.54 $Y=0.63 $X2=0
+ $Y2=0
cc_927 N_A_1865_367#_c_1290_n N_Q_N_c_1827_n 0.0203681f $X=13.705 $Y=1.35 $X2=0
+ $Y2=0
cc_928 N_A_1865_367#_M1031_g N_Q_N_c_1828_n 0.00255411f $X=13.92 $Y=2.465 $X2=0
+ $Y2=0
cc_929 N_A_1865_367#_c_1304_n N_Q_N_c_1828_n 0.0133692f $X=13.54 $Y=2.43 $X2=0
+ $Y2=0
cc_930 N_A_1865_367#_c_1290_n N_Q_N_c_1828_n 0.0790399f $X=13.705 $Y=1.35 $X2=0
+ $Y2=0
cc_931 N_A_1865_367#_c_1296_n N_Q_N_c_1828_n 0.00329721f $X=13.92 $Y=1.35 $X2=0
+ $Y2=0
cc_932 N_A_1865_367#_M1034_g N_Q_N_c_1836_n 0.00311959f $X=12.4 $Y=2.135 $X2=0
+ $Y2=0
cc_933 N_A_1865_367#_c_1304_n N_Q_N_c_1836_n 0.0336685f $X=13.54 $Y=2.43 $X2=0
+ $Y2=0
cc_934 N_A_1865_367#_c_1285_n N_Q_c_1854_n 0.00454529f $X=13.915 $Y=1.185 $X2=0
+ $Y2=0
cc_935 N_A_1865_367#_c_1290_n N_Q_c_1854_n 0.0803342f $X=13.705 $Y=1.35 $X2=0
+ $Y2=0
cc_936 N_A_1865_367#_c_1296_n N_Q_c_1854_n 0.0164393f $X=13.92 $Y=1.35 $X2=0
+ $Y2=0
cc_937 N_A_1865_367#_c_1292_n N_VGND_M1028_d 0.0115995f $X=10.94 $Y=0.49 $X2=0
+ $Y2=0
cc_938 N_A_1865_367#_c_1293_n N_VGND_M1028_d 6.52315e-19 $X=11.11 $Y=0.49 $X2=0
+ $Y2=0
cc_939 N_A_1865_367#_c_1289_n N_VGND_M1024_d 0.0100696f $X=13.54 $Y=0.63 $X2=0
+ $Y2=0
cc_940 N_A_1865_367#_c_1289_n N_VGND_M1012_s 0.00902952f $X=13.54 $Y=0.63 $X2=0
+ $Y2=0
cc_941 N_A_1865_367#_c_1290_n N_VGND_M1012_s 0.00707283f $X=13.705 $Y=1.35 $X2=0
+ $Y2=0
cc_942 N_A_1865_367#_c_1291_n N_VGND_c_1872_n 0.0027804f $X=9.635 $Y=0.49 $X2=0
+ $Y2=0
cc_943 N_A_1865_367#_c_1292_n N_VGND_c_1872_n 0.0230478f $X=10.94 $Y=0.49 $X2=0
+ $Y2=0
cc_944 N_A_1865_367#_c_1293_n N_VGND_c_1872_n 0.00840977f $X=11.11 $Y=0.49 $X2=0
+ $Y2=0
cc_945 N_A_1865_367#_c_1291_n N_VGND_c_1873_n 0.0213833f $X=9.635 $Y=0.49 $X2=0
+ $Y2=0
cc_946 N_A_1865_367#_c_1292_n N_VGND_c_1873_n 0.011692f $X=10.94 $Y=0.49 $X2=0
+ $Y2=0
cc_947 N_A_1865_367#_c_1288_n N_VGND_c_1874_n 4.79526e-19 $X=11.65 $Y=0.43 $X2=0
+ $Y2=0
cc_948 N_A_1865_367#_c_1289_n N_VGND_c_1874_n 0.0229777f $X=13.54 $Y=0.63 $X2=0
+ $Y2=0
cc_949 N_A_1865_367#_c_1295_n N_VGND_c_1874_n 0.00483704f $X=11.97 $Y=0.49 $X2=0
+ $Y2=0
cc_950 N_A_1865_367#_c_1283_n N_VGND_c_1875_n 6.22765e-19 $X=12.24 $Y=1.235
+ $X2=0 $Y2=0
cc_951 N_A_1865_367#_c_1288_n N_VGND_c_1875_n 0.00777248f $X=11.65 $Y=0.43 $X2=0
+ $Y2=0
cc_952 N_A_1865_367#_c_1289_n N_VGND_c_1875_n 0.00893096f $X=13.54 $Y=0.63 $X2=0
+ $Y2=0
cc_953 N_A_1865_367#_c_1292_n N_VGND_c_1875_n 0.00401349f $X=10.94 $Y=0.49 $X2=0
+ $Y2=0
cc_954 N_A_1865_367#_c_1293_n N_VGND_c_1875_n 0.0651577f $X=11.11 $Y=0.49 $X2=0
+ $Y2=0
cc_955 N_A_1865_367#_c_1285_n N_VGND_c_1876_n 0.00770281f $X=13.915 $Y=1.185
+ $X2=0 $Y2=0
cc_956 N_A_1865_367#_c_1289_n N_VGND_c_1876_n 0.0245519f $X=13.54 $Y=0.63 $X2=0
+ $Y2=0
cc_957 N_A_1865_367#_c_1289_n N_VGND_c_1877_n 0.0145152f $X=13.54 $Y=0.63 $X2=0
+ $Y2=0
cc_958 N_A_1865_367#_c_1285_n N_VGND_c_1881_n 0.00556333f $X=13.915 $Y=1.185
+ $X2=0 $Y2=0
cc_959 N_A_1865_367#_c_1289_n N_VGND_c_1881_n 0.00205231f $X=13.54 $Y=0.63 $X2=0
+ $Y2=0
cc_960 N_A_1865_367#_c_1285_n N_VGND_c_1882_n 0.0123288f $X=13.915 $Y=1.185
+ $X2=0 $Y2=0
cc_961 N_A_1865_367#_c_1288_n N_VGND_c_1882_n 0.0111008f $X=11.65 $Y=0.43 $X2=0
+ $Y2=0
cc_962 N_A_1865_367#_c_1289_n N_VGND_c_1882_n 0.0410815f $X=13.54 $Y=0.63 $X2=0
+ $Y2=0
cc_963 N_A_1865_367#_c_1291_n N_VGND_c_1882_n 0.012466f $X=9.635 $Y=0.49 $X2=0
+ $Y2=0
cc_964 N_A_1865_367#_c_1292_n N_VGND_c_1882_n 0.0252944f $X=10.94 $Y=0.49 $X2=0
+ $Y2=0
cc_965 N_A_1865_367#_c_1293_n N_VGND_c_1882_n 0.0390518f $X=11.11 $Y=0.49 $X2=0
+ $Y2=0
cc_966 N_A_1865_367#_c_1291_n N_A_1789_141#_c_2049_n 0.00191683f $X=9.635
+ $Y=0.49 $X2=0 $Y2=0
cc_967 N_A_1865_367#_c_1280_n N_A_1789_141#_c_2050_n 0.00644674f $X=11.74
+ $Y=1.235 $X2=0 $Y2=0
cc_968 N_A_1865_367#_c_1288_n N_A_1789_141#_c_2050_n 0.00306728f $X=11.65
+ $Y=0.43 $X2=0 $Y2=0
cc_969 N_A_1865_367#_c_1294_n N_A_1789_141#_c_2050_n 0.0246304f $X=11.8 $Y=0.49
+ $X2=0 $Y2=0
cc_970 N_A_1865_367#_M1020_d N_A_1789_141#_c_2056_n 0.00791266f $X=9.38 $Y=0.705
+ $X2=0 $Y2=0
cc_971 N_A_1865_367#_c_1291_n N_A_1789_141#_c_2056_n 0.0203362f $X=9.635 $Y=0.49
+ $X2=0 $Y2=0
cc_972 N_A_1865_367#_c_1292_n N_A_1789_141#_c_2056_n 0.0742569f $X=10.94 $Y=0.49
+ $X2=0 $Y2=0
cc_973 N_A_1865_367#_c_1294_n N_A_1789_141#_c_2056_n 0.00302334f $X=11.8 $Y=0.49
+ $X2=0 $Y2=0
cc_974 N_A_1865_367#_c_1292_n A_1986_57# 0.0038632f $X=10.94 $Y=0.49 $X2=-0.19
+ $Y2=-0.245
cc_975 N_VPWR_c_1465_n N_A_286_423#_c_1602_n 0.0171734f $X=2.005 $Y=2.325 $X2=0
+ $Y2=0
cc_976 N_VPWR_c_1462_n N_A_286_423#_c_1602_n 0.0102628f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_977 N_VPWR_c_1465_n N_A_286_423#_c_1603_n 0.0136256f $X=2.005 $Y=2.325 $X2=0
+ $Y2=0
cc_978 N_VPWR_c_1465_n N_A_286_423#_c_1605_n 0.0288267f $X=2.005 $Y=2.325 $X2=0
+ $Y2=0
cc_979 N_VPWR_c_1477_n N_A_286_423#_c_1606_n 0.027763f $X=5.98 $Y=3.33 $X2=0
+ $Y2=0
cc_980 N_VPWR_c_1462_n N_A_286_423#_c_1606_n 0.0295777f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_981 N_VPWR_c_1465_n N_A_286_423#_c_1607_n 0.0137879f $X=2.005 $Y=2.325 $X2=0
+ $Y2=0
cc_982 N_VPWR_c_1477_n N_A_286_423#_c_1607_n 0.00582061f $X=5.98 $Y=3.33 $X2=0
+ $Y2=0
cc_983 N_VPWR_c_1462_n N_A_286_423#_c_1607_n 0.005987f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_984 N_VPWR_c_1466_n N_A_761_396#_c_1744_n 0.0129217f $X=6.145 $Y=2.395 $X2=0
+ $Y2=0
cc_985 N_VPWR_c_1477_n N_A_761_396#_c_1744_n 0.107232f $X=5.98 $Y=3.33 $X2=0
+ $Y2=0
cc_986 N_VPWR_c_1462_n N_A_761_396#_c_1744_n 0.0596947f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_987 N_VPWR_c_1477_n N_A_761_396#_c_1745_n 0.0114622f $X=5.98 $Y=3.33 $X2=0
+ $Y2=0
cc_988 N_VPWR_c_1462_n N_A_761_396#_c_1745_n 0.00657784f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_989 N_VPWR_c_1466_n N_A_761_396#_c_1746_n 0.0419791f $X=6.145 $Y=2.395 $X2=0
+ $Y2=0
cc_990 N_VPWR_c_1462_n N_A_1781_367#_M1030_s 0.00219634f $X=14.16 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_991 N_VPWR_c_1462_n N_A_1781_367#_M1009_s 0.00220439f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_992 N_VPWR_c_1475_n N_A_1781_367#_c_1777_n 0.105921f $X=10.87 $Y=3.33 $X2=0
+ $Y2=0
cc_993 N_VPWR_c_1462_n N_A_1781_367#_c_1777_n 0.0674764f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_994 N_VPWR_M1009_d N_A_1971_388#_c_1799_n 0.00799374f $X=10.815 $Y=1.835
+ $X2=0 $Y2=0
cc_995 N_VPWR_M1034_d N_Q_N_c_1836_n 0.00875838f $X=12.475 $Y=1.815 $X2=0 $Y2=0
cc_996 N_VPWR_c_1462_n N_Q_M1031_d 0.00410879f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_997 N_VPWR_c_1480_n N_Q_c_1855_n 0.0163977f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_998 N_VPWR_c_1462_n N_Q_c_1855_n 0.00959046f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_999 N_A_286_423#_c_1605_n A_459_423# 0.00356941f $X=2.355 $Y=2.735 $X2=-0.19
+ $Y2=1.655
cc_1000 N_A_286_423#_c_1605_n N_A_531_423#_c_1658_n 0.0426803f $X=2.355 $Y=2.735
+ $X2=0 $Y2=0
cc_1001 N_A_286_423#_c_1606_n N_A_531_423#_c_1658_n 0.0192005f $X=3.06 $Y=2.82
+ $X2=0 $Y2=0
cc_1002 N_A_286_423#_c_1608_n N_A_531_423#_c_1658_n 0.0172103f $X=3.225 $Y=2.325
+ $X2=0 $Y2=0
cc_1003 N_A_286_423#_c_1608_n N_A_531_423#_c_1659_n 0.0213232f $X=3.225 $Y=2.325
+ $X2=0 $Y2=0
cc_1004 N_A_286_423#_c_1603_n N_A_531_423#_c_1660_n 0.0139268f $X=2.27 $Y=1.83
+ $X2=0 $Y2=0
cc_1005 N_A_286_423#_c_1606_n N_A_761_396#_c_1743_n 0.00591519f $X=3.06 $Y=2.82
+ $X2=0 $Y2=0
cc_1006 N_A_286_423#_c_1608_n N_A_761_396#_c_1743_n 0.0189549f $X=3.225 $Y=2.325
+ $X2=0 $Y2=0
cc_1007 N_A_286_423#_c_1606_n N_A_761_396#_c_1745_n 4.10092e-19 $X=3.06 $Y=2.82
+ $X2=0 $Y2=0
cc_1008 N_A_531_423#_c_1656_n N_A_761_396#_M1008_s 0.00383379f $X=4.3 $Y=2.545
+ $X2=-0.19 $Y2=-0.245
cc_1009 N_A_531_423#_c_1656_n N_A_761_396#_c_1743_n 0.040302f $X=4.3 $Y=2.545
+ $X2=0 $Y2=0
cc_1010 N_A_531_423#_c_1664_n N_A_761_396#_c_1743_n 0.013787f $X=4.385 $Y=2.63
+ $X2=0 $Y2=0
cc_1011 N_A_531_423#_c_1663_n N_A_761_396#_c_1744_n 0.0599212f $X=4.915 $Y=2.63
+ $X2=0 $Y2=0
cc_1012 N_A_531_423#_c_1664_n N_A_761_396#_c_1744_n 0.0125751f $X=4.385 $Y=2.63
+ $X2=0 $Y2=0
cc_1013 N_A_531_423#_c_1663_n N_A_761_396#_c_1746_n 0.0134079f $X=4.915 $Y=2.63
+ $X2=0 $Y2=0
cc_1014 N_A_531_423#_c_1665_n N_A_761_396#_c_1746_n 0.0207642f $X=5.08 $Y=2.19
+ $X2=0 $Y2=0
cc_1015 N_A_531_423#_c_1655_n N_VGND_c_1879_n 0.0108889f $X=4.22 $Y=0.665 $X2=0
+ $Y2=0
cc_1016 N_A_531_423#_c_1655_n N_VGND_c_1882_n 0.0114747f $X=4.22 $Y=0.665 $X2=0
+ $Y2=0
cc_1017 N_A_531_423#_c_1652_n N_A_231_53#_c_1997_n 0.0146043f $X=3.225 $Y=1.27
+ $X2=0 $Y2=0
cc_1018 N_A_531_423#_c_1652_n N_A_404_53#_c_2028_n 0.0194437f $X=3.225 $Y=1.27
+ $X2=0 $Y2=0
cc_1019 N_A_531_423#_c_1654_n N_A_404_53#_c_2028_n 0.00428399f $X=4.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1020 N_A_531_423#_c_1654_n N_A_404_53#_c_2029_n 0.0259264f $X=4.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1021 N_A_531_423#_c_1655_n N_A_404_53#_c_2029_n 0.0326647f $X=4.22 $Y=0.665
+ $X2=0 $Y2=0
cc_1022 N_A_1781_367#_M1009_s N_A_1971_388#_c_1799_n 0.00527995f $X=10.395
+ $Y=1.835 $X2=0 $Y2=0
cc_1023 N_Q_c_1854_n N_VGND_c_1881_n 0.016728f $X=14.13 $Y=0.43 $X2=0 $Y2=0
cc_1024 N_Q_M1012_d N_VGND_c_1882_n 0.00415073f $X=13.99 $Y=0.235 $X2=0 $Y2=0
cc_1025 N_Q_c_1854_n N_VGND_c_1882_n 0.00978392f $X=14.13 $Y=0.43 $X2=0 $Y2=0
cc_1026 N_VGND_c_1869_n N_A_231_53#_c_1992_n 0.0158413f $X=1.73 $Y=0.475 $X2=0
+ $Y2=0
cc_1027 N_VGND_c_1878_n N_A_231_53#_c_1992_n 0.0163773f $X=1.565 $Y=0 $X2=0
+ $Y2=0
cc_1028 N_VGND_c_1882_n N_A_231_53#_c_1992_n 0.00959046f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1029 N_VGND_c_1869_n N_A_231_53#_c_1995_n 0.0199134f $X=1.73 $Y=0.475 $X2=0
+ $Y2=0
cc_1030 N_VGND_c_1882_n N_A_231_53#_c_1996_n 0.00127743f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1031 N_VGND_c_1879_n N_A_404_53#_c_2028_n 0.0931028f $X=5.46 $Y=0 $X2=0 $Y2=0
cc_1032 N_VGND_c_1882_n N_A_404_53#_c_2028_n 0.0564782f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1033 N_VGND_c_1879_n N_A_404_53#_c_2030_n 0.0190464f $X=5.46 $Y=0 $X2=0 $Y2=0
cc_1034 N_VGND_c_1882_n N_A_404_53#_c_2030_n 0.0123847f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1035 N_VGND_c_1873_n N_A_1789_141#_c_2049_n 0.00579524f $X=10.43 $Y=0 $X2=0
+ $Y2=0
cc_1036 N_VGND_c_1882_n N_A_1789_141#_c_2049_n 0.00943528f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1037 N_VGND_M1028_d N_A_1789_141#_c_2056_n 0.0225316f $X=10.34 $Y=0.285 $X2=0
+ $Y2=0
cc_1038 N_A_231_53#_c_1994_n N_A_404_53#_c_2028_n 0.00833393f $X=2.555 $Y=0.915
+ $X2=0 $Y2=0
cc_1039 N_A_231_53#_c_1997_n N_A_404_53#_c_2028_n 0.0175837f $X=2.72 $Y=0.805
+ $X2=0 $Y2=0
cc_1040 N_A_231_53#_c_1996_n N_A_404_53#_c_2030_n 0.0219649f $X=2.165 $Y=0.942
+ $X2=0 $Y2=0
cc_1041 N_A_231_53#_c_1997_n N_A_404_53#_c_2030_n 0.00231108f $X=2.72 $Y=0.805
+ $X2=0 $Y2=0
cc_1042 N_A_1789_141#_c_2056_n A_1986_57# 0.0046747f $X=11.29 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
