* File: sky130_fd_sc_lp__a22oi_0.spice
* Created: Wed Sep  2 09:22:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22oi_0.pex.spice"
.subckt sky130_fd_sc_lp__a22oi_0  VNB VPB B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1006 A_121_47# N_B2_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1218 PD=0.63 PS=1.42 NRD=14.28 NRS=7.14 M=1 R=2.8 SA=75000.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g A_121_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0441 PD=0.84 PS=0.63 NRD=7.14 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1007 A_307_47# N_A1_M1007_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0882 PD=0.63 PS=0.84 NRD=14.28 NRS=32.856 M=1 R=2.8 SA=75001.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_307_47# VNB NSHORT L=0.15 W=0.42 AD=0.1239
+ AS=0.0441 PD=1.43 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_B2_M1004_g N_A_45_405#_M1004_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.192 PD=0.92 PS=1.88 NRD=0 NRS=10.7562 M=1 R=4.26667 SA=75000.2
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1005 N_A_45_405#_M1005_d N_B1_M1005_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_45_405#_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_45_405#_M1000_d N_A2_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
c_52 VPB 0 9.10919e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a22oi_0.pxi.spice"
*
.ends
*
*
