* File: sky130_fd_sc_lp__einvn_lp.pxi.spice
* Created: Fri Aug 28 10:33:12 2020
* 
x_PM_SKY130_FD_SC_LP__EINVN_LP%TE_B N_TE_B_M1003_g N_TE_B_c_40_n N_TE_B_M1004_g
+ N_TE_B_M1001_g N_TE_B_c_41_n N_TE_B_M1002_g TE_B N_TE_B_c_38_n N_TE_B_c_39_n
+ PM_SKY130_FD_SC_LP__EINVN_LP%TE_B
x_PM_SKY130_FD_SC_LP__EINVN_LP%A_28_148# N_A_28_148#_M1003_s N_A_28_148#_M1004_s
+ N_A_28_148#_M1000_g N_A_28_148#_c_79_n N_A_28_148#_c_80_n N_A_28_148#_c_81_n
+ N_A_28_148#_c_82_n N_A_28_148#_c_83_n N_A_28_148#_c_84_n N_A_28_148#_c_85_n
+ PM_SKY130_FD_SC_LP__EINVN_LP%A_28_148#
x_PM_SKY130_FD_SC_LP__EINVN_LP%A N_A_c_127_n N_A_M1006_g N_A_M1005_g N_A_c_129_n
+ A A N_A_c_126_n PM_SKY130_FD_SC_LP__EINVN_LP%A
x_PM_SKY130_FD_SC_LP__EINVN_LP%VPWR N_VPWR_M1004_d N_VPWR_c_154_n VPWR
+ N_VPWR_c_155_n N_VPWR_c_153_n N_VPWR_c_157_n PM_SKY130_FD_SC_LP__EINVN_LP%VPWR
x_PM_SKY130_FD_SC_LP__EINVN_LP%Z N_Z_M1005_d N_Z_M1006_d Z Z Z Z Z N_Z_c_175_n
+ PM_SKY130_FD_SC_LP__EINVN_LP%Z
x_PM_SKY130_FD_SC_LP__EINVN_LP%VGND N_VGND_M1001_d N_VGND_c_191_n VGND
+ N_VGND_c_192_n N_VGND_c_193_n N_VGND_c_194_n N_VGND_c_195_n
+ PM_SKY130_FD_SC_LP__EINVN_LP%VGND
cc_1 VNB N_TE_B_M1003_g 0.0372965f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.95
cc_2 VNB N_TE_B_M1001_g 0.029527f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.95
cc_3 VNB N_TE_B_c_38_n 2.86395e-19 $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.745
cc_4 VNB N_TE_B_c_39_n 0.0100087f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.787
cc_5 VNB N_A_28_148#_c_79_n 0.0241253f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.995
cc_6 VNB N_A_28_148#_c_80_n 0.0132148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_28_148#_c_81_n 0.0151008f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.745
cc_8 VNB N_A_28_148#_c_82_n 0.00770964f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.787
cc_9 VNB N_A_28_148#_c_83_n 0.0154629f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.995
cc_10 VNB N_A_28_148#_c_84_n 0.0354887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_28_148#_c_85_n 0.0183452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_M1005_g 0.0372064f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.57
cc_13 VNB A 0.0329741f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=2.57
cc_14 VNB N_A_c_126_n 0.0482368f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.787
cc_15 VNB N_VPWR_c_153_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.787
cc_16 VNB Z 0.0125231f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.58
cc_17 VNB N_Z_c_175_n 0.0298333f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.787
cc_18 VNB N_VGND_c_191_n 0.0295777f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.57
cc_19 VNB N_VGND_c_192_n 0.0298687f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.95
cc_20 VNB N_VGND_c_193_n 0.0337261f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.787
cc_21 VNB N_VGND_c_194_n 0.183573f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.787
cc_22 VNB N_VGND_c_195_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.745
cc_23 VPB N_TE_B_c_40_n 0.0227167f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.995
cc_24 VPB N_TE_B_c_41_n 0.0197177f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=1.995
cc_25 VPB N_TE_B_c_38_n 7.43345e-19 $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.745
cc_26 VPB N_TE_B_c_39_n 0.0592311f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=1.787
cc_27 VPB N_A_28_148#_c_80_n 0.0624214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_A_c_127_n 0.0239203f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.58
cc_29 VPB N_A_M1005_g 0.0134684f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.57
cc_30 VPB N_A_c_129_n 0.030327f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=0.95
cc_31 VPB N_VPWR_c_154_n 0.00113276f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=1.58
cc_32 VPB N_VPWR_c_155_n 0.0396425f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.787
cc_33 VPB N_VPWR_c_153_n 0.0644005f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.787
cc_34 VPB N_VPWR_c_157_n 0.025574f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.745
cc_35 VPB Z 0.0767489f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=1.58
cc_36 N_TE_B_M1003_g N_A_28_148#_c_79_n 0.011203f $X=0.5 $Y=0.95 $X2=0 $Y2=0
cc_37 N_TE_B_M1001_g N_A_28_148#_c_79_n 0.00179788f $X=0.86 $Y=0.95 $X2=0 $Y2=0
cc_38 N_TE_B_M1003_g N_A_28_148#_c_80_n 0.0181885f $X=0.5 $Y=0.95 $X2=0 $Y2=0
cc_39 N_TE_B_c_38_n N_A_28_148#_c_80_n 0.0397016f $X=0.77 $Y=1.745 $X2=0 $Y2=0
cc_40 N_TE_B_c_39_n N_A_28_148#_c_80_n 0.00445382f $X=0.86 $Y=1.787 $X2=0 $Y2=0
cc_41 N_TE_B_M1003_g N_A_28_148#_c_81_n 0.014163f $X=0.5 $Y=0.95 $X2=0 $Y2=0
cc_42 N_TE_B_M1001_g N_A_28_148#_c_81_n 0.0134019f $X=0.86 $Y=0.95 $X2=0 $Y2=0
cc_43 N_TE_B_c_38_n N_A_28_148#_c_81_n 0.0241878f $X=0.77 $Y=1.745 $X2=0 $Y2=0
cc_44 N_TE_B_c_39_n N_A_28_148#_c_81_n 0.00766073f $X=0.86 $Y=1.787 $X2=0 $Y2=0
cc_45 N_TE_B_M1003_g N_A_28_148#_c_82_n 0.0050081f $X=0.5 $Y=0.95 $X2=0 $Y2=0
cc_46 N_TE_B_M1001_g N_A_28_148#_c_83_n 0.00136939f $X=0.86 $Y=0.95 $X2=0 $Y2=0
cc_47 N_TE_B_c_38_n N_A_28_148#_c_83_n 0.00113941f $X=0.77 $Y=1.745 $X2=0 $Y2=0
cc_48 N_TE_B_c_39_n N_A_28_148#_c_83_n 6.34951e-19 $X=0.86 $Y=1.787 $X2=0 $Y2=0
cc_49 N_TE_B_M1001_g N_A_28_148#_c_84_n 0.0182282f $X=0.86 $Y=0.95 $X2=0 $Y2=0
cc_50 N_TE_B_c_39_n N_A_28_148#_c_84_n 0.00470494f $X=0.86 $Y=1.787 $X2=0 $Y2=0
cc_51 N_TE_B_M1001_g N_A_28_148#_c_85_n 0.0119472f $X=0.86 $Y=0.95 $X2=0 $Y2=0
cc_52 N_TE_B_c_41_n N_A_c_127_n 0.0382892f $X=1.135 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_53 N_TE_B_c_38_n N_A_c_129_n 5.99741e-19 $X=0.77 $Y=1.745 $X2=0 $Y2=0
cc_54 N_TE_B_c_39_n N_A_c_129_n 0.0384168f $X=0.86 $Y=1.787 $X2=0 $Y2=0
cc_55 N_TE_B_c_38_n N_VPWR_M1004_d 0.00261538f $X=0.77 $Y=1.745 $X2=-0.19
+ $Y2=-0.245
cc_56 N_TE_B_c_40_n N_VPWR_c_154_n 0.0179465f $X=0.605 $Y=1.995 $X2=0 $Y2=0
cc_57 N_TE_B_c_41_n N_VPWR_c_154_n 0.0210774f $X=1.135 $Y=1.995 $X2=0 $Y2=0
cc_58 N_TE_B_c_38_n N_VPWR_c_154_n 0.0144051f $X=0.77 $Y=1.745 $X2=0 $Y2=0
cc_59 N_TE_B_c_39_n N_VPWR_c_154_n 5.41299e-19 $X=0.86 $Y=1.787 $X2=0 $Y2=0
cc_60 N_TE_B_c_41_n N_VPWR_c_155_n 0.00838537f $X=1.135 $Y=1.995 $X2=0 $Y2=0
cc_61 N_TE_B_c_40_n N_VPWR_c_153_n 0.0153108f $X=0.605 $Y=1.995 $X2=0 $Y2=0
cc_62 N_TE_B_c_41_n N_VPWR_c_153_n 0.014363f $X=1.135 $Y=1.995 $X2=0 $Y2=0
cc_63 N_TE_B_c_40_n N_VPWR_c_157_n 0.00838537f $X=0.605 $Y=1.995 $X2=0 $Y2=0
cc_64 N_TE_B_c_39_n Z 0.00530957f $X=0.86 $Y=1.787 $X2=0 $Y2=0
cc_65 N_TE_B_M1003_g N_VGND_c_191_n 0.00144992f $X=0.5 $Y=0.95 $X2=0 $Y2=0
cc_66 N_TE_B_M1001_g N_VGND_c_191_n 0.00958992f $X=0.86 $Y=0.95 $X2=0 $Y2=0
cc_67 N_TE_B_M1003_g N_VGND_c_192_n 0.00347474f $X=0.5 $Y=0.95 $X2=0 $Y2=0
cc_68 N_TE_B_M1001_g N_VGND_c_192_n 0.00298903f $X=0.86 $Y=0.95 $X2=0 $Y2=0
cc_69 N_TE_B_M1003_g N_VGND_c_194_n 0.00438782f $X=0.5 $Y=0.95 $X2=0 $Y2=0
cc_70 N_TE_B_M1001_g N_VGND_c_194_n 0.00368577f $X=0.86 $Y=0.95 $X2=0 $Y2=0
cc_71 N_A_28_148#_c_83_n N_A_M1005_g 5.59058e-19 $X=1.34 $Y=1.315 $X2=0 $Y2=0
cc_72 N_A_28_148#_c_84_n N_A_M1005_g 0.0174678f $X=1.34 $Y=1.435 $X2=0 $Y2=0
cc_73 N_A_28_148#_c_84_n N_A_c_129_n 3.28026e-19 $X=1.34 $Y=1.435 $X2=0 $Y2=0
cc_74 N_A_28_148#_c_85_n A 5.8445e-19 $X=1.34 $Y=1.27 $X2=0 $Y2=0
cc_75 N_A_28_148#_c_85_n N_A_c_126_n 0.0235569f $X=1.34 $Y=1.27 $X2=0 $Y2=0
cc_76 N_A_28_148#_c_80_n N_VPWR_c_153_n 0.0117186f $X=0.34 $Y=2.215 $X2=0 $Y2=0
cc_77 N_A_28_148#_c_80_n N_VPWR_c_157_n 0.0200856f $X=0.34 $Y=2.215 $X2=0 $Y2=0
cc_78 N_A_28_148#_c_83_n Z 0.00983164f $X=1.34 $Y=1.315 $X2=0 $Y2=0
cc_79 N_A_28_148#_c_84_n Z 9.32903e-19 $X=1.34 $Y=1.435 $X2=0 $Y2=0
cc_80 N_A_28_148#_c_83_n N_Z_c_175_n 0.0155396f $X=1.34 $Y=1.315 $X2=0 $Y2=0
cc_81 N_A_28_148#_c_84_n N_Z_c_175_n 0.00119474f $X=1.34 $Y=1.435 $X2=0 $Y2=0
cc_82 N_A_28_148#_c_85_n N_Z_c_175_n 0.00261167f $X=1.34 $Y=1.27 $X2=0 $Y2=0
cc_83 N_A_28_148#_c_79_n N_VGND_c_191_n 0.0110409f $X=0.285 $Y=0.95 $X2=0 $Y2=0
cc_84 N_A_28_148#_c_81_n N_VGND_c_191_n 0.0182886f $X=1.175 $Y=1.315 $X2=0 $Y2=0
cc_85 N_A_28_148#_c_83_n N_VGND_c_191_n 0.00418345f $X=1.34 $Y=1.315 $X2=0 $Y2=0
cc_86 N_A_28_148#_c_84_n N_VGND_c_191_n 3.70349e-19 $X=1.34 $Y=1.435 $X2=0 $Y2=0
cc_87 N_A_28_148#_c_85_n N_VGND_c_191_n 0.00266036f $X=1.34 $Y=1.27 $X2=0 $Y2=0
cc_88 N_A_28_148#_c_79_n N_VGND_c_192_n 0.00556708f $X=0.285 $Y=0.95 $X2=0 $Y2=0
cc_89 N_A_28_148#_c_85_n N_VGND_c_193_n 0.00359559f $X=1.34 $Y=1.27 $X2=0 $Y2=0
cc_90 N_A_28_148#_c_79_n N_VGND_c_194_n 0.00931589f $X=0.285 $Y=0.95 $X2=0 $Y2=0
cc_91 N_A_28_148#_c_85_n N_VGND_c_194_n 0.00438782f $X=1.34 $Y=1.27 $X2=0 $Y2=0
cc_92 N_A_c_127_n N_VPWR_c_154_n 0.00404338f $X=1.625 $Y=1.99 $X2=0 $Y2=0
cc_93 N_A_c_127_n N_VPWR_c_155_n 0.00898892f $X=1.625 $Y=1.99 $X2=0 $Y2=0
cc_94 N_A_c_127_n N_VPWR_c_153_n 0.0169236f $X=1.625 $Y=1.99 $X2=0 $Y2=0
cc_95 N_A_c_127_n Z 0.0242274f $X=1.625 $Y=1.99 $X2=0 $Y2=0
cc_96 N_A_M1005_g Z 0.0173083f $X=1.82 $Y=0.95 $X2=0 $Y2=0
cc_97 N_A_c_129_n Z 0.01261f $X=1.82 $Y=1.915 $X2=0 $Y2=0
cc_98 N_A_M1005_g N_Z_c_175_n 0.0193358f $X=1.82 $Y=0.95 $X2=0 $Y2=0
cc_99 A N_Z_c_175_n 0.0373274f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_100 N_A_c_126_n N_Z_c_175_n 0.00135581f $X=1.945 $Y=0.465 $X2=0 $Y2=0
cc_101 A N_VGND_c_191_n 0.0176573f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_102 N_A_c_126_n N_VGND_c_191_n 0.00341686f $X=1.945 $Y=0.465 $X2=0 $Y2=0
cc_103 A N_VGND_c_193_n 0.0280571f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_104 N_A_c_126_n N_VGND_c_193_n 0.00291928f $X=1.945 $Y=0.465 $X2=0 $Y2=0
cc_105 A N_VGND_c_194_n 0.0247997f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_106 N_A_c_126_n N_VGND_c_194_n 0.00122917f $X=1.945 $Y=0.465 $X2=0 $Y2=0
cc_107 N_VPWR_c_155_n Z 0.0345914f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_108 N_VPWR_c_153_n Z 0.021083f $X=2.16 $Y=3.33 $X2=0 $Y2=0
