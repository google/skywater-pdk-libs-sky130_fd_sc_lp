* File: sky130_fd_sc_lp__nand4bb_m.pxi.spice
* Created: Fri Aug 28 10:52:55 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4BB_M%B_N N_B_N_M1005_g N_B_N_M1003_g B_N B_N
+ N_B_N_c_76_n N_B_N_c_77_n PM_SKY130_FD_SC_LP__NAND4BB_M%B_N
x_PM_SKY130_FD_SC_LP__NAND4BB_M%D N_D_M1000_g N_D_M1009_g D D D N_D_c_111_n
+ N_D_c_112_n PM_SKY130_FD_SC_LP__NAND4BB_M%D
x_PM_SKY130_FD_SC_LP__NAND4BB_M%C N_C_M1011_g N_C_M1002_g C C C N_C_c_150_n
+ N_C_c_151_n PM_SKY130_FD_SC_LP__NAND4BB_M%C
x_PM_SKY130_FD_SC_LP__NAND4BB_M%A_27_151# N_A_27_151#_M1005_s
+ N_A_27_151#_M1003_s N_A_27_151#_c_188_n N_A_27_151#_M1006_g
+ N_A_27_151#_M1010_g N_A_27_151#_c_190_n N_A_27_151#_c_186_n
+ N_A_27_151#_c_191_n N_A_27_151#_c_187_n N_A_27_151#_c_193_n
+ N_A_27_151#_c_194_n PM_SKY130_FD_SC_LP__NAND4BB_M%A_27_151#
x_PM_SKY130_FD_SC_LP__NAND4BB_M%A_469_125# N_A_469_125#_M1007_d
+ N_A_469_125#_M1008_d N_A_469_125#_M1001_g N_A_469_125#_c_242_n
+ N_A_469_125#_M1004_g N_A_469_125#_c_243_n N_A_469_125#_c_249_n
+ N_A_469_125#_c_244_n N_A_469_125#_c_245_n
+ PM_SKY130_FD_SC_LP__NAND4BB_M%A_469_125#
x_PM_SKY130_FD_SC_LP__NAND4BB_M%A_N N_A_N_M1008_g N_A_N_M1007_g N_A_N_c_294_n
+ N_A_N_c_295_n A_N A_N N_A_N_c_297_n PM_SKY130_FD_SC_LP__NAND4BB_M%A_N
x_PM_SKY130_FD_SC_LP__NAND4BB_M%VPWR N_VPWR_M1003_d N_VPWR_M1002_d
+ N_VPWR_M1004_d N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n
+ N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n VPWR
+ N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_325_n N_VPWR_c_337_n
+ PM_SKY130_FD_SC_LP__NAND4BB_M%VPWR
x_PM_SKY130_FD_SC_LP__NAND4BB_M%Y N_Y_M1001_d N_Y_M1009_d N_Y_M1010_d
+ N_Y_c_379_n N_Y_c_376_n N_Y_c_388_n N_Y_c_380_n N_Y_c_377_n Y Y Y Y
+ PM_SKY130_FD_SC_LP__NAND4BB_M%Y
x_PM_SKY130_FD_SC_LP__NAND4BB_M%VGND N_VGND_M1005_d N_VGND_M1007_s
+ N_VGND_c_423_n N_VGND_c_424_n VGND N_VGND_c_425_n N_VGND_c_426_n
+ N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n
+ PM_SKY130_FD_SC_LP__NAND4BB_M%VGND
cc_1 VNB N_B_N_M1003_g 0.0024985f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.225
cc_2 VNB B_N 0.00759902f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_B_N_c_76_n 0.0331926f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.45
cc_4 VNB N_B_N_c_77_n 0.0233361f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.285
cc_5 VNB N_D_M1009_g 0.00234628f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.225
cc_6 VNB D 0.00756004f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB D 0.00380107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_D_c_111_n 0.0370303f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.615
cc_9 VNB N_D_c_112_n 0.0170182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_C_M1002_g 0.00216995f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.225
cc_11 VNB C 0.0151809f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_C_c_150_n 0.0328422f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.285
cc_13 VNB N_C_c_151_n 0.016489f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.295
cc_14 VNB N_A_27_151#_M1006_g 0.0337119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_151#_c_186_n 0.0088718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_151#_c_187_n 0.0277123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_469_125#_M1001_g 0.0280609f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB N_A_469_125#_c_242_n 0.02998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_469_125#_c_243_n 0.00792343f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.285
cc_20 VNB N_A_469_125#_c_244_n 0.0441604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_469_125#_c_245_n 0.00883216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_N_M1008_g 0.00696326f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.965
cc_23 VNB N_A_N_M1007_g 0.0293655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_N_c_294_n 0.0099121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_N_c_295_n 0.0199691f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.45
cc_26 VNB A_N 0.0102242f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.285
cc_27 VNB N_A_N_c_297_n 0.037183f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.45
cc_28 VNB N_VPWR_c_325_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_376_n 0.00136085f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.45
cc_30 VNB N_Y_c_377_n 0.00710371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB Y 6.15562e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_423_n 0.0369034f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_33 VNB N_VGND_c_424_n 0.0138343f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.45
cc_34 VNB N_VGND_c_425_n 0.0213956f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.295
cc_35 VNB N_VGND_c_426_n 0.0620888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_427_n 0.0165789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_428_n 0.28068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_429_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_430_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_B_N_M1003_g 0.0340363f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.225
cc_41 VPB B_N 0.00820146f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_42 VPB N_D_M1009_g 0.0348834f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.225
cc_43 VPB N_C_M1002_g 0.0308357f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.225
cc_44 VPB N_A_27_151#_c_188_n 0.109145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_27_151#_M1006_g 0.047992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_27_151#_c_190_n 0.0160323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_27_151#_c_191_n 0.0131836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_27_151#_c_187_n 0.0242475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_27_151#_c_193_n 0.015436f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_27_151#_c_194_n 0.0475761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_469_125#_c_242_n 0.0234411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_469_125#_M1004_g 0.0225053f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.45
cc_53 VPB N_A_469_125#_c_243_n 0.00882177f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.285
cc_54 VPB N_A_469_125#_c_249_n 0.0181303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_469_125#_c_245_n 0.0175761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_N_M1008_g 0.0424516f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.965
cc_57 VPB N_VPWR_c_326_n 0.00306214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_327_n 0.0112443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_328_n 0.0144472f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.45
cc_60 VPB N_VPWR_c_329_n 0.0346547f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_330_n 0.0251973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_331_n 0.00334761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_332_n 0.0191525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_333_n 0.00299251f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_334_n 0.0203639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_335_n 0.0330106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_325_n 0.0905106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_337_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_Y_c_379_n 0.00134272f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.45
cc_70 VPB N_Y_c_380_n 0.00909498f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.615
cc_71 VPB Y 0.00107157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB Y 0.0180099f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB Y 0.00562654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 N_B_N_M1003_g N_D_M1009_g 0.0211471f $X=0.54 $Y=2.225 $X2=0 $Y2=0
cc_75 B_N N_D_M1009_g 0.003044f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 B_N D 0.0036354f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_B_N_c_77_n D 0.00116915f $X=0.53 $Y=1.285 $X2=0 $Y2=0
cc_78 B_N D 0.0249831f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B_N_c_76_n D 2.94137e-19 $X=0.53 $Y=1.45 $X2=0 $Y2=0
cc_80 B_N N_D_c_111_n 0.00224802f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_81 N_B_N_c_76_n N_D_c_111_n 0.0204463f $X=0.53 $Y=1.45 $X2=0 $Y2=0
cc_82 B_N N_D_c_112_n 6.24354e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 N_B_N_c_77_n N_D_c_112_n 0.0107193f $X=0.53 $Y=1.285 $X2=0 $Y2=0
cc_84 N_B_N_M1003_g N_A_27_151#_c_190_n 0.00578621f $X=0.54 $Y=2.225 $X2=0 $Y2=0
cc_85 N_B_N_c_77_n N_A_27_151#_c_186_n 0.00405812f $X=0.53 $Y=1.285 $X2=0 $Y2=0
cc_86 N_B_N_M1003_g N_A_27_151#_c_191_n 0.00514826f $X=0.54 $Y=2.225 $X2=0 $Y2=0
cc_87 B_N N_A_27_151#_c_191_n 0.00364259f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B_N_c_76_n N_A_27_151#_c_191_n 0.00185637f $X=0.53 $Y=1.45 $X2=0 $Y2=0
cc_89 N_B_N_M1003_g N_A_27_151#_c_187_n 0.0136072f $X=0.54 $Y=2.225 $X2=0 $Y2=0
cc_90 B_N N_A_27_151#_c_187_n 0.0396609f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B_N_c_76_n N_A_27_151#_c_187_n 0.00808178f $X=0.53 $Y=1.45 $X2=0 $Y2=0
cc_92 N_B_N_c_77_n N_A_27_151#_c_187_n 0.00630608f $X=0.53 $Y=1.285 $X2=0 $Y2=0
cc_93 N_B_N_M1003_g N_A_27_151#_c_193_n 5.60406e-19 $X=0.54 $Y=2.225 $X2=0 $Y2=0
cc_94 N_B_N_M1003_g N_A_27_151#_c_194_n 0.0101874f $X=0.54 $Y=2.225 $X2=0 $Y2=0
cc_95 N_B_N_M1003_g N_VPWR_c_326_n 0.00351907f $X=0.54 $Y=2.225 $X2=0 $Y2=0
cc_96 B_N N_VPWR_c_326_n 0.00271962f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_97 B_N N_VGND_c_423_n 0.0155644f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_98 N_B_N_c_76_n N_VGND_c_423_n 5.73431e-19 $X=0.53 $Y=1.45 $X2=0 $Y2=0
cc_99 N_B_N_c_77_n N_VGND_c_423_n 0.00570173f $X=0.53 $Y=1.285 $X2=0 $Y2=0
cc_100 N_B_N_c_77_n N_VGND_c_425_n 0.00352953f $X=0.53 $Y=1.285 $X2=0 $Y2=0
cc_101 N_B_N_c_77_n N_VGND_c_428_n 0.00434946f $X=0.53 $Y=1.285 $X2=0 $Y2=0
cc_102 N_D_M1009_g N_C_M1002_g 0.0280093f $X=1.16 $Y=2.265 $X2=0 $Y2=0
cc_103 D C 0.037378f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_104 D C 0.0195407f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_D_c_111_n C 3.35817e-19 $X=1.07 $Y=1.45 $X2=0 $Y2=0
cc_106 N_D_c_112_n C 6.82347e-19 $X=1.07 $Y=1.285 $X2=0 $Y2=0
cc_107 D N_C_c_150_n 0.00217778f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_108 N_D_c_111_n N_C_c_150_n 0.029679f $X=1.07 $Y=1.45 $X2=0 $Y2=0
cc_109 D N_C_c_151_n 0.00245869f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_110 N_D_c_112_n N_C_c_151_n 0.029679f $X=1.07 $Y=1.285 $X2=0 $Y2=0
cc_111 N_D_M1009_g N_A_27_151#_c_188_n 0.00619064f $X=1.16 $Y=2.265 $X2=0 $Y2=0
cc_112 N_D_M1009_g N_A_27_151#_c_190_n 2.74487e-19 $X=1.16 $Y=2.265 $X2=0 $Y2=0
cc_113 N_D_M1009_g N_VPWR_c_326_n 0.0109042f $X=1.16 $Y=2.265 $X2=0 $Y2=0
cc_114 N_D_c_111_n N_VPWR_c_326_n 0.001486f $X=1.07 $Y=1.45 $X2=0 $Y2=0
cc_115 N_D_M1009_g N_VPWR_c_325_n 7.64857e-19 $X=1.16 $Y=2.265 $X2=0 $Y2=0
cc_116 N_D_M1009_g N_Y_c_379_n 0.0017418f $X=1.16 $Y=2.265 $X2=0 $Y2=0
cc_117 N_D_M1009_g N_Y_c_380_n 0.00551383f $X=1.16 $Y=2.265 $X2=0 $Y2=0
cc_118 D N_Y_c_380_n 0.00116478f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_119 D N_VGND_c_423_n 0.0427176f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_120 N_D_c_111_n N_VGND_c_423_n 0.00114563f $X=1.07 $Y=1.45 $X2=0 $Y2=0
cc_121 N_D_c_112_n N_VGND_c_423_n 0.00335495f $X=1.07 $Y=1.285 $X2=0 $Y2=0
cc_122 D N_VGND_c_426_n 0.00584355f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_123 N_D_c_112_n N_VGND_c_426_n 0.00112698f $X=1.07 $Y=1.285 $X2=0 $Y2=0
cc_124 D N_VGND_c_428_n 0.00593617f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_125 N_D_c_112_n N_VGND_c_428_n 8.98888e-19 $X=1.07 $Y=1.285 $X2=0 $Y2=0
cc_126 N_C_M1002_g N_A_27_151#_c_188_n 0.00631055f $X=1.59 $Y=2.265 $X2=0 $Y2=0
cc_127 N_C_M1002_g N_A_27_151#_M1006_g 0.0232983f $X=1.59 $Y=2.265 $X2=0 $Y2=0
cc_128 C N_A_27_151#_M1006_g 0.0120993f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_129 N_C_c_150_n N_A_27_151#_M1006_g 0.019346f $X=1.61 $Y=1.45 $X2=0 $Y2=0
cc_130 N_C_c_151_n N_A_27_151#_M1006_g 0.016996f $X=1.61 $Y=1.285 $X2=0 $Y2=0
cc_131 N_C_M1002_g N_VPWR_c_326_n 6.28877e-19 $X=1.59 $Y=2.265 $X2=0 $Y2=0
cc_132 N_C_M1002_g N_VPWR_c_328_n 0.00168787f $X=1.59 $Y=2.265 $X2=0 $Y2=0
cc_133 N_C_M1002_g N_VPWR_c_325_n 8.46637e-19 $X=1.59 $Y=2.265 $X2=0 $Y2=0
cc_134 N_C_M1002_g N_Y_c_379_n 9.06486e-19 $X=1.59 $Y=2.265 $X2=0 $Y2=0
cc_135 C N_Y_c_388_n 0.00855366f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 N_C_c_150_n N_Y_c_380_n 0.00159214f $X=1.61 $Y=1.45 $X2=0 $Y2=0
cc_137 N_C_M1002_g Y 0.00101827f $X=1.59 $Y=2.265 $X2=0 $Y2=0
cc_138 C Y 0.0181726f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_139 N_C_c_150_n Y 0.00101177f $X=1.61 $Y=1.45 $X2=0 $Y2=0
cc_140 N_C_M1002_g Y 0.0150873f $X=1.59 $Y=2.265 $X2=0 $Y2=0
cc_141 C Y 0.0162843f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_142 N_C_c_150_n Y 0.0024638f $X=1.61 $Y=1.45 $X2=0 $Y2=0
cc_143 N_C_M1002_g Y 6.29185e-19 $X=1.59 $Y=2.265 $X2=0 $Y2=0
cc_144 C N_VGND_c_426_n 0.00827836f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_145 N_C_c_151_n N_VGND_c_426_n 0.00213646f $X=1.61 $Y=1.285 $X2=0 $Y2=0
cc_146 C N_VGND_c_428_n 0.00840958f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_147 N_C_c_151_n N_VGND_c_428_n 0.00234871f $X=1.61 $Y=1.285 $X2=0 $Y2=0
cc_148 C A_319_151# 0.00506696f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_149 N_A_27_151#_M1006_g N_A_469_125#_M1001_g 0.0590246f $X=2.06 $Y=0.965
+ $X2=0 $Y2=0
cc_150 N_A_27_151#_M1006_g N_A_469_125#_c_242_n 0.0293419f $X=2.06 $Y=0.965
+ $X2=0 $Y2=0
cc_151 N_A_27_151#_M1006_g N_A_469_125#_c_243_n 2.46672e-19 $X=2.06 $Y=0.965
+ $X2=0 $Y2=0
cc_152 N_A_27_151#_c_188_n N_VPWR_c_326_n 0.00333245f $X=1.985 $Y=3.03 $X2=0
+ $Y2=0
cc_153 N_A_27_151#_c_191_n N_VPWR_c_326_n 0.0297479f $X=0.325 $Y=2.29 $X2=0
+ $Y2=0
cc_154 N_A_27_151#_c_187_n N_VPWR_c_326_n 6.67855e-19 $X=0.322 $Y=2.185 $X2=0
+ $Y2=0
cc_155 N_A_27_151#_c_188_n N_VPWR_c_327_n 0.0171967f $X=1.985 $Y=3.03 $X2=0
+ $Y2=0
cc_156 N_A_27_151#_c_190_n N_VPWR_c_327_n 0.00806623f $X=0.385 $Y=2.775 $X2=0
+ $Y2=0
cc_157 N_A_27_151#_c_193_n N_VPWR_c_327_n 0.023053f $X=0.575 $Y=2.94 $X2=0 $Y2=0
cc_158 N_A_27_151#_c_194_n N_VPWR_c_327_n 0.00127201f $X=0.575 $Y=2.94 $X2=0
+ $Y2=0
cc_159 N_A_27_151#_c_188_n N_VPWR_c_328_n 0.0169454f $X=1.985 $Y=3.03 $X2=0
+ $Y2=0
cc_160 N_A_27_151#_M1006_g N_VPWR_c_328_n 0.011318f $X=2.06 $Y=0.965 $X2=0 $Y2=0
cc_161 N_A_27_151#_M1006_g N_VPWR_c_329_n 0.0102335f $X=2.06 $Y=0.965 $X2=0
+ $Y2=0
cc_162 N_A_27_151#_c_193_n N_VPWR_c_330_n 0.0338243f $X=0.575 $Y=2.94 $X2=0
+ $Y2=0
cc_163 N_A_27_151#_c_194_n N_VPWR_c_330_n 0.00920052f $X=0.575 $Y=2.94 $X2=0
+ $Y2=0
cc_164 N_A_27_151#_c_188_n N_VPWR_c_332_n 0.0176856f $X=1.985 $Y=3.03 $X2=0
+ $Y2=0
cc_165 N_A_27_151#_c_188_n N_VPWR_c_334_n 0.00742396f $X=1.985 $Y=3.03 $X2=0
+ $Y2=0
cc_166 N_A_27_151#_c_188_n N_VPWR_c_325_n 0.0446884f $X=1.985 $Y=3.03 $X2=0
+ $Y2=0
cc_167 N_A_27_151#_c_193_n N_VPWR_c_325_n 0.0182917f $X=0.575 $Y=2.94 $X2=0
+ $Y2=0
cc_168 N_A_27_151#_c_194_n N_VPWR_c_325_n 0.00772789f $X=0.575 $Y=2.94 $X2=0
+ $Y2=0
cc_169 N_A_27_151#_c_188_n N_Y_c_379_n 0.00471472f $X=1.985 $Y=3.03 $X2=0 $Y2=0
cc_170 N_A_27_151#_M1006_g N_Y_c_388_n 0.00709875f $X=2.06 $Y=0.965 $X2=0 $Y2=0
cc_171 N_A_27_151#_M1006_g Y 0.0158347f $X=2.06 $Y=0.965 $X2=0 $Y2=0
cc_172 N_A_27_151#_M1006_g Y 0.013969f $X=2.06 $Y=0.965 $X2=0 $Y2=0
cc_173 N_A_27_151#_M1006_g Y 0.0120593f $X=2.06 $Y=0.965 $X2=0 $Y2=0
cc_174 N_A_27_151#_M1006_g N_VGND_c_426_n 0.00352953f $X=2.06 $Y=0.965 $X2=0
+ $Y2=0
cc_175 N_A_27_151#_M1006_g N_VGND_c_428_n 0.00434946f $X=2.06 $Y=0.965 $X2=0
+ $Y2=0
cc_176 N_A_27_151#_c_186_n N_VGND_c_428_n 0.0117098f $X=0.26 $Y=0.925 $X2=0
+ $Y2=0
cc_177 N_A_469_125#_M1004_g N_A_N_M1008_g 0.0112537f $X=2.49 $Y=2.265 $X2=0
+ $Y2=0
cc_178 N_A_469_125#_c_243_n N_A_N_M1008_g 0.0148391f $X=3.205 $Y=1.725 $X2=0
+ $Y2=0
cc_179 N_A_469_125#_c_249_n N_A_N_M1008_g 0.0128151f $X=3.37 $Y=2.2 $X2=0 $Y2=0
cc_180 N_A_469_125#_c_244_n N_A_N_M1008_g 7.59948e-19 $X=3.57 $Y=0.49 $X2=0
+ $Y2=0
cc_181 N_A_469_125#_c_245_n N_A_N_M1008_g 0.00826472f $X=3.44 $Y=1.725 $X2=0
+ $Y2=0
cc_182 N_A_469_125#_c_244_n N_A_N_M1007_g 0.0279486f $X=3.57 $Y=0.49 $X2=0 $Y2=0
cc_183 N_A_469_125#_M1001_g N_A_N_c_295_n 5.38997e-19 $X=2.42 $Y=0.965 $X2=0
+ $Y2=0
cc_184 N_A_469_125#_c_242_n N_A_N_c_295_n 0.0224749f $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_185 N_A_469_125#_c_245_n N_A_N_c_295_n 0.00913473f $X=3.44 $Y=1.725 $X2=0
+ $Y2=0
cc_186 N_A_469_125#_M1001_g A_N 0.00473812f $X=2.42 $Y=0.965 $X2=0 $Y2=0
cc_187 N_A_469_125#_c_243_n A_N 0.0136373f $X=3.205 $Y=1.725 $X2=0 $Y2=0
cc_188 N_A_469_125#_c_244_n A_N 0.04212f $X=3.57 $Y=0.49 $X2=0 $Y2=0
cc_189 N_A_469_125#_c_245_n A_N 0.00858401f $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_190 N_A_469_125#_M1001_g N_A_N_c_297_n 0.00491828f $X=2.42 $Y=0.965 $X2=0
+ $Y2=0
cc_191 N_A_469_125#_c_242_n N_VPWR_c_329_n 0.00486684f $X=2.49 $Y=1.89 $X2=0
+ $Y2=0
cc_192 N_A_469_125#_M1004_g N_VPWR_c_329_n 0.00751743f $X=2.49 $Y=2.265 $X2=0
+ $Y2=0
cc_193 N_A_469_125#_c_243_n N_VPWR_c_329_n 0.0147797f $X=3.205 $Y=1.725 $X2=0
+ $Y2=0
cc_194 N_A_469_125#_c_249_n N_VPWR_c_329_n 0.00369102f $X=3.37 $Y=2.2 $X2=0
+ $Y2=0
cc_195 N_A_469_125#_M1004_g N_VPWR_c_334_n 0.00259749f $X=2.49 $Y=2.265 $X2=0
+ $Y2=0
cc_196 N_A_469_125#_M1004_g N_VPWR_c_325_n 0.00344639f $X=2.49 $Y=2.265 $X2=0
+ $Y2=0
cc_197 N_A_469_125#_M1001_g N_Y_c_376_n 0.0156809f $X=2.42 $Y=0.965 $X2=0 $Y2=0
cc_198 N_A_469_125#_c_242_n N_Y_c_376_n 0.00456662f $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_199 N_A_469_125#_c_243_n N_Y_c_376_n 0.00465092f $X=3.205 $Y=1.725 $X2=0
+ $Y2=0
cc_200 N_A_469_125#_M1001_g N_Y_c_388_n 0.0024849f $X=2.42 $Y=0.965 $X2=0 $Y2=0
cc_201 N_A_469_125#_M1001_g N_Y_c_377_n 0.00449476f $X=2.42 $Y=0.965 $X2=0 $Y2=0
cc_202 N_A_469_125#_c_242_n N_Y_c_377_n 0.00378455f $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_203 N_A_469_125#_c_243_n N_Y_c_377_n 0.0100217f $X=3.205 $Y=1.725 $X2=0 $Y2=0
cc_204 N_A_469_125#_M1001_g Y 0.00626945f $X=2.42 $Y=0.965 $X2=0 $Y2=0
cc_205 N_A_469_125#_c_242_n Y 0.0107813f $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_206 N_A_469_125#_c_243_n Y 0.0201441f $X=3.205 $Y=1.725 $X2=0 $Y2=0
cc_207 N_A_469_125#_c_242_n Y 0.00371868f $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_208 N_A_469_125#_c_243_n Y 0.00631577f $X=3.205 $Y=1.725 $X2=0 $Y2=0
cc_209 N_A_469_125#_M1004_g Y 0.00262139f $X=2.49 $Y=2.265 $X2=0 $Y2=0
cc_210 N_A_469_125#_M1001_g N_VGND_c_426_n 0.00352953f $X=2.42 $Y=0.965 $X2=0
+ $Y2=0
cc_211 N_A_469_125#_c_244_n N_VGND_c_427_n 0.00906426f $X=3.57 $Y=0.49 $X2=0
+ $Y2=0
cc_212 N_A_469_125#_M1007_d N_VGND_c_428_n 0.0048747f $X=3.43 $Y=0.235 $X2=0
+ $Y2=0
cc_213 N_A_469_125#_M1001_g N_VGND_c_428_n 0.00434946f $X=2.42 $Y=0.965 $X2=0
+ $Y2=0
cc_214 N_A_469_125#_c_244_n N_VGND_c_428_n 0.00703984f $X=3.57 $Y=0.49 $X2=0
+ $Y2=0
cc_215 N_A_N_M1008_g N_VPWR_c_329_n 0.00813791f $X=3.155 $Y=2.265 $X2=0 $Y2=0
cc_216 N_A_N_M1008_g N_VPWR_c_335_n 0.00312414f $X=3.155 $Y=2.265 $X2=0 $Y2=0
cc_217 N_A_N_M1008_g N_VPWR_c_325_n 0.00410284f $X=3.155 $Y=2.265 $X2=0 $Y2=0
cc_218 A_N N_Y_c_377_n 0.0247701f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_219 N_A_N_c_297_n N_Y_c_377_n 0.00107f $X=3.22 $Y=1 $X2=0 $Y2=0
cc_220 A_N Y 0.00443526f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_221 N_A_N_M1007_g N_VGND_c_424_n 0.0117237f $X=3.355 $Y=0.445 $X2=0 $Y2=0
cc_222 A_N N_VGND_c_424_n 0.0123156f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_223 N_A_N_c_297_n N_VGND_c_424_n 0.00127228f $X=3.22 $Y=1 $X2=0 $Y2=0
cc_224 N_A_N_M1007_g N_VGND_c_427_n 0.00486043f $X=3.355 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A_N_M1007_g N_VGND_c_428_n 0.00936946f $X=3.355 $Y=0.445 $X2=0 $Y2=0
cc_226 A_N N_VGND_c_428_n 0.00139836f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_227 N_VPWR_c_328_n Y 0.013281f $X=1.805 $Y=2.33 $X2=0 $Y2=0
cc_228 N_VPWR_c_328_n Y 0.0257328f $X=1.805 $Y=2.33 $X2=0 $Y2=0
cc_229 N_VPWR_c_329_n Y 0.0137913f $X=2.705 $Y=2.33 $X2=0 $Y2=0
cc_230 N_VPWR_c_325_n Y 0.0112034f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_231 N_Y_c_388_n A_427_151# 0.00433061f $X=2.36 $Y=1.13 $X2=-0.19 $Y2=-0.245
