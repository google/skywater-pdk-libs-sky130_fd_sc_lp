* NGSPICE file created from sky130_fd_sc_lp__a21oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.56e+11p pd=6.24e+06u as=1.3734e+12p ps=1.226e+07u
M1001 a_27_367# B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1002 Y B1 VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=7.14e+11p ps=6.74e+06u
M1003 a_110_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1004 a_27_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B1 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_110_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A1 a_110_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A2 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_110_47# A1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

