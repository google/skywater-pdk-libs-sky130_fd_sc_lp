* NGSPICE file created from sky130_fd_sc_lp__a21oi_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21oi_lp A1 A2 B1 VGND VNB VPB VPWR Y
M1000 Y B1 a_31_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=5.65e+11p ps=5.13e+06u
M1001 a_31_409# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1002 a_132_47# A2 VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.394e+11p ps=2.82e+06u
M1003 a_324_47# B1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.764e+11p ps=1.68e+06u
M1004 VGND B1 a_324_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_31_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A1 a_132_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

