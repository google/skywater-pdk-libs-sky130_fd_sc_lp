* File: sky130_fd_sc_lp__iso1n_lp2.pex.spice
* Created: Wed Sep  2 09:58:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__ISO1N_LP2%SLEEP_B 1 3 5 6 10 12 14 15 16 23
c43 16 0 4.55941e-20 $X=0.72 $Y=1.665
r44 21 23 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.67 $Y=1.68
+ $X2=0.805 $Y2=1.68
r45 18 21 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.495 $Y=1.68
+ $X2=0.67 $Y2=1.68
r46 16 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.68 $X2=0.67 $Y2=1.68
r47 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.855 $Y=1.04
+ $X2=0.855 $Y2=0.755
r48 8 23 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.805 $Y=1.845
+ $X2=0.805 $Y2=1.68
r49 8 10 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.805 $Y=1.845
+ $X2=0.805 $Y2=2.545
r50 7 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.57 $Y=1.115
+ $X2=0.495 $Y2=1.115
r51 6 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.78 $Y=1.115
+ $X2=0.855 $Y2=1.04
r52 6 7 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.78 $Y=1.115 $X2=0.57
+ $Y2=1.115
r53 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.495 $Y2=1.68
r54 4 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.19
+ $X2=0.495 $Y2=1.115
r55 4 5 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.495 $Y=1.19
+ $X2=0.495 $Y2=1.515
r56 1 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.04
+ $X2=0.495 $Y2=1.115
r57 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.04 $X2=0.495
+ $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP2%A_27_109# 1 2 9 13 17 23 26 29 35 37 41 43
+ 44 46 47
c79 23 0 3.36635e-19 $X=1.675 $Y=1.24
c80 13 0 4.55941e-20 $X=1.375 $Y=2.545
r81 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.335
+ $Y=1.33 $X2=1.335 $Y2=1.33
r82 43 44 9.57885 $w=5.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.37 $Y=2.19
+ $X2=0.37 $Y2=2.025
r83 38 41 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.25
+ $X2=0.28 $Y2=1.25
r84 37 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=1.25
+ $X2=1.335 $Y2=1.25
r85 37 38 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.17 $Y=1.25
+ $X2=0.445 $Y2=1.25
r86 33 43 2.11073 $w=5.08e-07 $l=9e-08 $layer=LI1_cond $X=0.37 $Y=2.28 $X2=0.37
+ $Y2=2.19
r87 33 35 14.5406 $w=5.08e-07 $l=6.2e-07 $layer=LI1_cond $X=0.37 $Y=2.28
+ $X2=0.37 $Y2=2.9
r88 31 41 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=1.335
+ $X2=0.28 $Y2=1.25
r89 31 44 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.2 $Y=1.335 $X2=0.2
+ $Y2=2.025
r90 27 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=1.165
+ $X2=0.28 $Y2=1.25
r91 27 29 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=1.165
+ $X2=0.28 $Y2=0.755
r92 25 47 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.335 $Y=1.67
+ $X2=1.335 $Y2=1.33
r93 25 26 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.67
+ $X2=1.335 $Y2=1.835
r94 22 47 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.335 $Y=1.315
+ $X2=1.335 $Y2=1.33
r95 22 23 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.335 $Y=1.24
+ $X2=1.675 $Y2=1.24
r96 19 22 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=1.285 $Y=1.24
+ $X2=1.335 $Y2=1.24
r97 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.675 $Y=1.165
+ $X2=1.675 $Y2=1.24
r98 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.675 $Y=1.165
+ $X2=1.675 $Y2=0.755
r99 13 26 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.375 $Y=2.545
+ $X2=1.375 $Y2=1.835
r100 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.285 $Y=1.165
+ $X2=1.285 $Y2=1.24
r101 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.285 $Y=1.165
+ $X2=1.285 $Y2=0.755
r102 2 43 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=2.045 $X2=0.54 $Y2=2.19
r103 2 35 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=2.045 $X2=0.54 $Y2=2.9
r104 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.545 $X2=0.28 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP2%A 3 7 11 13 14 20
c41 14 0 1.47195e-19 $X=2.64 $Y=1.295
r42 20 22 2.92121 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.525 $Y=1.435
+ $X2=2.545 $Y2=1.435
r43 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.525
+ $Y=1.33 $X2=2.525 $Y2=1.33
r44 18 20 49.6606 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.185 $Y=1.435
+ $X2=2.525 $Y2=1.435
r45 14 21 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.33
+ $X2=2.525 $Y2=1.33
r46 13 21 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.16 $Y=1.33
+ $X2=2.525 $Y2=1.33
r47 9 22 21.2229 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.545 $Y=1.165
+ $X2=2.545 $Y2=1.435
r48 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.545 $Y=1.165
+ $X2=2.545 $Y2=0.755
r49 5 18 21.2229 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.185 $Y=1.165
+ $X2=2.185 $Y2=1.435
r50 5 7 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.185 $Y=1.165
+ $X2=2.185 $Y2=0.755
r51 1 18 46.7394 $w=3.3e-07 $l=4.34511e-07 $layer=POLY_cond $X=1.865 $Y=1.705
+ $X2=2.185 $Y2=1.435
r52 1 3 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.865 $Y=1.705
+ $X2=1.865 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP2%A_350_109# 1 2 9 13 17 20 23 27 31 32 37
+ 39
c69 20 0 1.20445e-19 $X=1.78 $Y=1.675
r70 34 37 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.78 $Y=0.8 $X2=1.89
+ $Y2=0.8
r71 32 41 66.9034 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=3.155 $Y=1.34
+ $X2=3.155 $Y2=1.845
r72 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.1 $Y=1.34
+ $X2=3.1 $Y2=1.34
r73 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.1 $Y=1.675 $X2=3.1
+ $Y2=1.34
r74 28 39 4.39717 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=2.295 $Y=1.76 $X2=1.995
+ $Y2=1.76
r75 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.935 $Y=1.76
+ $X2=3.1 $Y2=1.675
r76 27 28 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.935 $Y=1.76
+ $X2=2.295 $Y2=1.76
r77 23 25 14.1536 $w=5.98e-07 $l=7.1e-07 $layer=LI1_cond $X=1.995 $Y=2.19
+ $X2=1.995 $Y2=2.9
r78 21 39 2.50573 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=1.845
+ $X2=1.995 $Y2=1.76
r79 21 23 6.87745 $w=5.98e-07 $l=3.45e-07 $layer=LI1_cond $X=1.995 $Y=1.845
+ $X2=1.995 $Y2=2.19
r80 20 39 2.50573 $w=3.85e-07 $l=2.53969e-07 $layer=LI1_cond $X=1.78 $Y=1.675
+ $X2=1.995 $Y2=1.76
r81 19 34 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.78 $Y=0.985
+ $X2=1.78 $Y2=0.8
r82 19 20 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.78 $Y=0.985
+ $X2=1.78 $Y2=1.675
r83 15 32 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=3.335 $Y=1.175
+ $X2=3.155 $Y2=1.34
r84 15 17 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.335 $Y=1.175
+ $X2=3.335 $Y2=0.755
r85 13 41 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.285 $Y=2.545
+ $X2=3.285 $Y2=1.845
r86 7 32 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=2.975 $Y=1.175
+ $X2=3.155 $Y2=1.34
r87 7 9 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.975 $Y=1.175
+ $X2=2.975 $Y2=0.755
r88 2 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=2.045 $X2=2.13 $Y2=2.9
r89 2 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=2.045 $X2=2.13 $Y2=2.19
r90 1 37 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.545 $X2=1.89 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP2%VPWR 1 2 9 15 20 21 22 24 34 35 38
r34 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r36 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r37 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=3.33
+ $X2=1.07 $Y2=3.33
r39 29 31 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=1.235 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 27 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.07 $Y2=3.33
r43 24 26 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 22 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 22 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 20 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.02 $Y2=3.33
r48 19 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.02 $Y2=3.33
r50 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.02 $Y=2.19 $X2=3.02
+ $Y2=2.9
r51 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=3.33
r52 13 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=2.9
r53 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.07 $Y=2.19 $X2=1.07
+ $Y2=2.9
r54 7 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245 $X2=1.07
+ $Y2=3.33
r55 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.9
r56 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=2.045 $X2=3.02 $Y2=2.9
r57 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=2.045 $X2=3.02 $Y2=2.19
r58 1 12 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=2.045 $X2=1.07 $Y2=2.9
r59 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=2.045 $X2=1.07 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP2%X 1 2 7 8 9 10 11 36 40 43
r19 43 44 0.646955 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=3.55 $Y=2.035
+ $X2=3.55 $Y2=2.025
r20 40 41 2.39308 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=3.55 $Y=0.925 $X2=3.55
+ $Y2=0.985
r21 11 33 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.55 $Y=2.405
+ $X2=3.55 $Y2=2.9
r22 11 29 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.55 $Y=2.405
+ $X2=3.55 $Y2=2.19
r23 10 29 4.12086 $w=3.28e-07 $l=1.18e-07 $layer=LI1_cond $X=3.55 $Y=2.072
+ $X2=3.55 $Y2=2.19
r24 10 43 1.29213 $w=3.28e-07 $l=3.7e-08 $layer=LI1_cond $X=3.55 $Y=2.072
+ $X2=3.55 $Y2=2.035
r25 10 44 1.56403 $w=2.78e-07 $l=3.8e-08 $layer=LI1_cond $X=3.575 $Y=1.987
+ $X2=3.575 $Y2=2.025
r26 9 10 13.2531 $w=2.78e-07 $l=3.22e-07 $layer=LI1_cond $X=3.575 $Y=1.665
+ $X2=3.575 $Y2=1.987
r27 8 9 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.575 $Y=1.295
+ $X2=3.575 $Y2=1.665
r28 7 40 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=3.55 $Y=0.912
+ $X2=3.55 $Y2=0.925
r29 7 36 5.48283 $w=3.28e-07 $l=1.57e-07 $layer=LI1_cond $X=3.55 $Y=0.912
+ $X2=3.55 $Y2=0.755
r30 7 8 12.2653 $w=2.78e-07 $l=2.98e-07 $layer=LI1_cond $X=3.575 $Y=0.997
+ $X2=3.575 $Y2=1.295
r31 7 41 0.493904 $w=2.78e-07 $l=1.2e-08 $layer=LI1_cond $X=3.575 $Y=0.997
+ $X2=3.575 $Y2=0.985
r32 2 33 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.045 $X2=3.55 $Y2=2.9
r33 2 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.045 $X2=3.55 $Y2=2.19
r34 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.545 $X2=3.55 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP2%KAGND 1 2 9 17 20 22 23
c48 23 0 1.8944e-19 $X=2.94 $Y=0.555
r49 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.94 $Y=0.555
+ $X2=2.94 $Y2=0.555
r50 19 22 2.9902 $w=7.18e-07 $l=1.8e-07 $layer=LI1_cond $X=2.76 $Y=0.625
+ $X2=2.94 $Y2=0.625
r51 19 20 13.4248 $w=7.18e-07 $l=3.15e-07 $layer=LI1_cond $X=2.76 $Y=0.625
+ $X2=2.445 $Y2=0.625
r52 17 20 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=1.385 $Y=0.35
+ $X2=2.445 $Y2=0.35
r53 15 17 10.4346 $w=7.18e-07 $l=1.35e-07 $layer=LI1_cond $X=1.25 $Y=0.625
+ $X2=1.385 $Y2=0.625
r54 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.25 $Y=0.555
+ $X2=1.25 $Y2=0.555
r55 12 15 2.9902 $w=7.18e-07 $l=1.8e-07 $layer=LI1_cond $X=1.07 $Y=0.625
+ $X2=1.25 $Y2=0.625
r56 9 23 0.654436 $w=2.3e-07 $l=1.02e-06 $layer=MET1_cond $X=1.92 $Y=0.555
+ $X2=2.94 $Y2=0.555
r57 9 16 0.429875 $w=2.3e-07 $l=6.7e-07 $layer=MET1_cond $X=1.92 $Y=0.555
+ $X2=1.25 $Y2=0.555
r58 2 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.545 $X2=2.76 $Y2=0.755
r59 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.545 $X2=1.07 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1N_LP2%VGND 1 5 8 15
r20 5 8 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r21 4 8 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r22 4 5 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r23 1 15 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=0.122
+ $X2=1.92 $Y2=0.123
r24 1 5 0.00397135 $w=3.84e-06 $l=1.22e-07 $layer=MET1_cond $X=1.92 $Y=0.122
+ $X2=1.92 $Y2=0
.ends

