* File: sky130_fd_sc_lp__ebufn_8.pxi.spice
* Created: Wed Sep  2 09:50:58 2020
* 
x_PM_SKY130_FD_SC_LP__EBUFN_8%A_84_21# N_A_84_21#_M1008_s N_A_84_21#_M1019_s
+ N_A_84_21#_M1003_g N_A_84_21#_M1006_g N_A_84_21#_M1005_g N_A_84_21#_M1011_g
+ N_A_84_21#_M1009_g N_A_84_21#_M1016_g N_A_84_21#_M1010_g N_A_84_21#_M1021_g
+ N_A_84_21#_M1017_g N_A_84_21#_M1022_g N_A_84_21#_M1025_g N_A_84_21#_M1024_g
+ N_A_84_21#_M1028_g N_A_84_21#_M1035_g N_A_84_21#_M1031_g N_A_84_21#_M1036_g
+ N_A_84_21#_c_208_n N_A_84_21#_c_219_n N_A_84_21#_c_220_n N_A_84_21#_c_253_p
+ N_A_84_21#_c_221_n N_A_84_21#_c_237_p N_A_84_21#_c_238_p N_A_84_21#_c_276_p
+ N_A_84_21#_c_325_p N_A_84_21#_c_222_n N_A_84_21#_c_223_n N_A_84_21#_c_209_n
+ N_A_84_21#_c_210_n PM_SKY130_FD_SC_LP__EBUFN_8%A_84_21#
x_PM_SKY130_FD_SC_LP__EBUFN_8%A_772_21# N_A_772_21#_M1020_s N_A_772_21#_M1012_s
+ N_A_772_21#_c_468_n N_A_772_21#_M1001_g N_A_772_21#_c_469_n
+ N_A_772_21#_c_470_n N_A_772_21#_c_471_n N_A_772_21#_M1004_g
+ N_A_772_21#_c_472_n N_A_772_21#_c_473_n N_A_772_21#_M1007_g
+ N_A_772_21#_c_474_n N_A_772_21#_c_475_n N_A_772_21#_M1015_g
+ N_A_772_21#_c_476_n N_A_772_21#_c_477_n N_A_772_21#_M1023_g
+ N_A_772_21#_c_478_n N_A_772_21#_c_479_n N_A_772_21#_M1026_g
+ N_A_772_21#_c_480_n N_A_772_21#_c_481_n N_A_772_21#_M1029_g
+ N_A_772_21#_c_482_n N_A_772_21#_c_483_n N_A_772_21#_M1037_g
+ N_A_772_21#_c_484_n N_A_772_21#_c_485_n N_A_772_21#_c_486_n
+ N_A_772_21#_c_487_n N_A_772_21#_c_488_n N_A_772_21#_c_489_n
+ N_A_772_21#_c_490_n N_A_772_21#_c_491_n N_A_772_21#_c_492_n
+ N_A_772_21#_c_493_n N_A_772_21#_c_494_n N_A_772_21#_c_497_n
+ N_A_772_21#_c_498_n N_A_772_21#_c_495_n N_A_772_21#_c_496_n
+ N_A_772_21#_c_499_n PM_SKY130_FD_SC_LP__EBUFN_8%A_772_21#
x_PM_SKY130_FD_SC_LP__EBUFN_8%TE_B N_TE_B_c_664_n N_TE_B_M1000_g N_TE_B_c_645_n
+ N_TE_B_c_646_n N_TE_B_c_667_n N_TE_B_M1002_g N_TE_B_c_647_n N_TE_B_c_669_n
+ N_TE_B_M1013_g N_TE_B_c_648_n N_TE_B_c_671_n N_TE_B_M1014_g N_TE_B_c_649_n
+ N_TE_B_c_673_n N_TE_B_M1018_g N_TE_B_c_650_n N_TE_B_c_675_n N_TE_B_M1027_g
+ N_TE_B_c_651_n N_TE_B_c_677_n N_TE_B_M1030_g N_TE_B_c_652_n N_TE_B_c_679_n
+ N_TE_B_M1034_g N_TE_B_c_653_n N_TE_B_M1020_g N_TE_B_M1012_g N_TE_B_c_654_n
+ N_TE_B_c_655_n N_TE_B_c_656_n N_TE_B_c_657_n N_TE_B_c_658_n N_TE_B_c_659_n
+ N_TE_B_c_660_n TE_B N_TE_B_c_661_n N_TE_B_c_662_n N_TE_B_c_663_n
+ N_TE_B_c_689_n PM_SKY130_FD_SC_LP__EBUFN_8%TE_B
x_PM_SKY130_FD_SC_LP__EBUFN_8%A N_A_c_841_n N_A_M1008_g N_A_M1019_g N_A_c_843_n
+ N_A_M1032_g N_A_M1033_g A N_A_c_846_n PM_SKY130_FD_SC_LP__EBUFN_8%A
x_PM_SKY130_FD_SC_LP__EBUFN_8%A_27_367# N_A_27_367#_M1006_s N_A_27_367#_M1011_s
+ N_A_27_367#_M1021_s N_A_27_367#_M1024_s N_A_27_367#_M1036_s
+ N_A_27_367#_M1002_s N_A_27_367#_M1014_s N_A_27_367#_M1027_s
+ N_A_27_367#_M1034_s N_A_27_367#_c_880_n N_A_27_367#_c_881_n
+ N_A_27_367#_c_894_n N_A_27_367#_c_896_n N_A_27_367#_c_898_n
+ N_A_27_367#_c_957_p N_A_27_367#_c_900_n N_A_27_367#_c_959_p
+ N_A_27_367#_c_902_n N_A_27_367#_c_882_n N_A_27_367#_c_983_p
+ N_A_27_367#_c_883_n N_A_27_367#_c_920_n N_A_27_367#_c_884_n
+ N_A_27_367#_c_927_n N_A_27_367#_c_885_n N_A_27_367#_c_886_n
+ N_A_27_367#_c_936_n N_A_27_367#_c_938_n N_A_27_367#_c_910_n
+ N_A_27_367#_c_912_n N_A_27_367#_c_985_p N_A_27_367#_c_986_p
+ N_A_27_367#_c_887_n N_A_27_367#_c_888_n N_A_27_367#_c_947_n
+ N_A_27_367#_c_889_n PM_SKY130_FD_SC_LP__EBUFN_8%A_27_367#
x_PM_SKY130_FD_SC_LP__EBUFN_8%Z N_Z_M1003_s N_Z_M1009_s N_Z_M1017_s N_Z_M1028_s
+ N_Z_M1006_d N_Z_M1016_d N_Z_M1022_d N_Z_M1035_d N_Z_c_1025_n N_Z_c_1011_n
+ N_Z_c_1018_n N_Z_c_1019_n N_Z_c_1012_n N_Z_c_1044_n N_Z_c_1013_n N_Z_c_1020_n
+ N_Z_c_1056_n N_Z_c_1014_n N_Z_c_1021_n N_Z_c_1069_n N_Z_c_1109_n N_Z_c_1015_n
+ N_Z_c_1022_n N_Z_c_1016_n N_Z_c_1023_n N_Z_c_1024_n Z Z N_Z_c_1017_n
+ PM_SKY130_FD_SC_LP__EBUFN_8%Z
x_PM_SKY130_FD_SC_LP__EBUFN_8%VPWR N_VPWR_M1000_d N_VPWR_M1013_d N_VPWR_M1018_d
+ N_VPWR_M1030_d N_VPWR_M1012_d N_VPWR_M1033_d N_VPWR_c_1148_n N_VPWR_c_1149_n
+ N_VPWR_c_1150_n N_VPWR_c_1151_n N_VPWR_c_1152_n N_VPWR_c_1153_n
+ N_VPWR_c_1154_n N_VPWR_c_1155_n N_VPWR_c_1156_n N_VPWR_c_1157_n
+ N_VPWR_c_1158_n N_VPWR_c_1159_n N_VPWR_c_1160_n VPWR N_VPWR_c_1161_n
+ N_VPWR_c_1162_n N_VPWR_c_1163_n N_VPWR_c_1164_n N_VPWR_c_1165_n
+ N_VPWR_c_1147_n PM_SKY130_FD_SC_LP__EBUFN_8%VPWR
x_PM_SKY130_FD_SC_LP__EBUFN_8%A_27_47# N_A_27_47#_M1003_d N_A_27_47#_M1005_d
+ N_A_27_47#_M1010_d N_A_27_47#_M1025_d N_A_27_47#_M1031_d N_A_27_47#_M1004_s
+ N_A_27_47#_M1015_s N_A_27_47#_M1026_s N_A_27_47#_M1037_s N_A_27_47#_c_1289_n
+ N_A_27_47#_c_1377_n N_A_27_47#_c_1291_n N_A_27_47#_c_1382_n
+ N_A_27_47#_c_1293_n N_A_27_47#_c_1387_n N_A_27_47#_c_1295_n
+ N_A_27_47#_c_1405_p N_A_27_47#_c_1281_n N_A_27_47#_c_1282_n
+ N_A_27_47#_c_1283_n N_A_27_47#_c_1313_n N_A_27_47#_c_1284_n
+ N_A_27_47#_c_1322_n N_A_27_47#_c_1285_n N_A_27_47#_c_1331_n
+ N_A_27_47#_c_1286_n N_A_27_47#_c_1287_n N_A_27_47#_c_1288_n
+ N_A_27_47#_c_1407_p N_A_27_47#_c_1408_p N_A_27_47#_c_1409_p
+ N_A_27_47#_c_1304_n N_A_27_47#_c_1305_n N_A_27_47#_c_1306_n
+ PM_SKY130_FD_SC_LP__EBUFN_8%A_27_47#
x_PM_SKY130_FD_SC_LP__EBUFN_8%VGND N_VGND_M1001_d N_VGND_M1007_d N_VGND_M1023_d
+ N_VGND_M1029_d N_VGND_M1020_d N_VGND_M1032_d N_VGND_c_1433_n N_VGND_c_1434_n
+ N_VGND_c_1435_n N_VGND_c_1436_n N_VGND_c_1437_n N_VGND_c_1438_n
+ N_VGND_c_1439_n N_VGND_c_1440_n N_VGND_c_1441_n N_VGND_c_1442_n
+ N_VGND_c_1443_n N_VGND_c_1444_n N_VGND_c_1445_n VGND N_VGND_c_1446_n
+ N_VGND_c_1447_n N_VGND_c_1448_n N_VGND_c_1449_n N_VGND_c_1450_n
+ N_VGND_c_1451_n PM_SKY130_FD_SC_LP__EBUFN_8%VGND
cc_1 VNB N_A_84_21#_M1003_g 0.0290743f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_2 VNB N_A_84_21#_M1006_g 7.21425e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_3 VNB N_A_84_21#_M1005_g 0.022138f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_4 VNB N_A_84_21#_M1011_g 4.54864e-19 $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_5 VNB N_A_84_21#_M1009_g 0.022166f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_6 VNB N_A_84_21#_M1016_g 4.5732e-19 $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=2.465
cc_7 VNB N_A_84_21#_M1010_g 0.0221931f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.655
cc_8 VNB N_A_84_21#_M1021_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=2.465
cc_9 VNB N_A_84_21#_M1017_g 0.0221931f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.655
cc_10 VNB N_A_84_21#_M1022_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_11 VNB N_A_84_21#_M1025_g 0.0221931f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_12 VNB N_A_84_21#_M1024_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_13 VNB N_A_84_21#_M1028_g 0.0221862f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=0.655
cc_14 VNB N_A_84_21#_M1035_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=2.465
cc_15 VNB N_A_84_21#_M1031_g 0.0228877f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=0.655
cc_16 VNB N_A_84_21#_M1036_g 4.7301e-19 $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=2.465
cc_17 VNB N_A_84_21#_c_208_n 0.0289829f $X=-0.19 $Y=-0.245 $X2=6.555 $Y2=1.56
cc_18 VNB N_A_84_21#_c_209_n 0.0109021f $X=-0.19 $Y=-0.245 $X2=8.695 $Y2=1.815
cc_19 VNB N_A_84_21#_c_210_n 0.173045f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.48
cc_20 VNB N_A_772_21#_c_468_n 0.0157034f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.315
cc_21 VNB N_A_772_21#_c_469_n 0.0122626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_772_21#_c_470_n 0.00729667f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.645
cc_23 VNB N_A_772_21#_c_471_n 0.0154996f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_24 VNB N_A_772_21#_c_472_n 0.0122626f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.315
cc_25 VNB N_A_772_21#_c_473_n 0.0154978f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_26 VNB N_A_772_21#_c_474_n 0.0122626f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_27 VNB N_A_772_21#_c_475_n 0.0154978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_772_21#_c_476_n 0.0122626f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_29 VNB N_A_772_21#_c_477_n 0.0154978f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.645
cc_30 VNB N_A_772_21#_c_478_n 0.0122626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_772_21#_c_479_n 0.0154978f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.655
cc_32 VNB N_A_772_21#_c_480_n 0.0122626f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.645
cc_33 VNB N_A_772_21#_c_481_n 0.0154978f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=2.465
cc_34 VNB N_A_772_21#_c_482_n 0.0122936f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.655
cc_35 VNB N_A_772_21#_c_483_n 0.0185886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_772_21#_c_484_n 0.0271614f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_37 VNB N_A_772_21#_c_485_n 0.0151555f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_38 VNB N_A_772_21#_c_486_n 0.00511394f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_39 VNB N_A_772_21#_c_487_n 0.00511394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_772_21#_c_488_n 0.00511394f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.645
cc_41 VNB N_A_772_21#_c_489_n 0.00511394f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_42 VNB N_A_772_21#_c_490_n 0.00511394f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_43 VNB N_A_772_21#_c_491_n 0.00511391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_772_21#_c_492_n 0.00514684f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.315
cc_45 VNB N_A_772_21#_c_493_n 0.0163188f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=0.655
cc_46 VNB N_A_772_21#_c_494_n 0.0134452f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.645
cc_47 VNB N_A_772_21#_c_495_n 0.00549712f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.315
cc_48 VNB N_A_772_21#_c_496_n 0.0465852f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=0.655
cc_49 VNB N_TE_B_c_645_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_TE_B_c_646_n 0.00412776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_TE_B_c_647_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_52 VNB N_TE_B_c_648_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_TE_B_c_649_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.645
cc_54 VNB N_TE_B_c_650_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_55 VNB N_TE_B_c_651_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=2.465
cc_56 VNB N_TE_B_c_652_n 0.00650026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_TE_B_c_653_n 0.0238096f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.315
cc_58 VNB N_TE_B_c_654_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.315
cc_59 VNB N_TE_B_c_655_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_60 VNB N_TE_B_c_656_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_61 VNB N_TE_B_c_657_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_TE_B_c_658_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.645
cc_63 VNB N_TE_B_c_659_n 0.00299786f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_64 VNB N_TE_B_c_660_n 0.00401376f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_65 VNB N_TE_B_c_661_n 0.0469976f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=0.655
cc_66 VNB N_TE_B_c_662_n 0.00608781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_TE_B_c_663_n 0.0200678f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.645
cc_68 VNB N_A_c_841_n 0.0162781f $X=-0.19 $Y=-0.245 $X2=8.72 $Y2=0.235
cc_69 VNB N_A_M1019_g 0.00725623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_c_843_n 0.0214901f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_71 VNB N_A_M1033_g 0.0111791f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_72 VNB A 0.00375127f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.315
cc_73 VNB N_A_c_846_n 0.0503072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_Z_c_1011_n 0.002006f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=2.465
cc_75 VNB N_Z_c_1012_n 0.00281069f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.645
cc_76 VNB N_Z_c_1013_n 0.00225436f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.645
cc_77 VNB N_Z_c_1014_n 0.00455029f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_78 VNB N_Z_c_1015_n 0.00229592f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=0.655
cc_79 VNB N_Z_c_1016_n 0.00229592f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=2.465
cc_80 VNB N_Z_c_1017_n 0.0183836f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=1.56
cc_81 VNB N_VPWR_c_1147_n 0.40251f $X=-0.19 $Y=-0.245 $X2=3.3 $Y2=1.48
cc_82 VNB N_A_27_47#_c_1281_n 9.12681e-19 $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.645
cc_83 VNB N_A_27_47#_c_1282_n 0.00632873f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_84 VNB N_A_27_47#_c_1283_n 0.00358753f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_85 VNB N_A_27_47#_c_1284_n 0.00538792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_27_47#_c_1285_n 0.00538792f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=0.655
cc_87 VNB N_A_27_47#_c_1286_n 0.00567035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_27_47#_c_1287_n 3.56834e-19 $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.48
cc_89 VNB N_A_27_47#_c_1288_n 0.0291024f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=1.56
cc_90 VNB N_VGND_c_1433_n 0.00238736f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_91 VNB N_VGND_c_1434_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_92 VNB N_VGND_c_1435_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=2.465
cc_93 VNB N_VGND_c_1436_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.655
cc_94 VNB N_VGND_c_1437_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=2.465
cc_95 VNB N_VGND_c_1438_n 0.011635f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.315
cc_96 VNB N_VGND_c_1439_n 0.0469785f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.655
cc_97 VNB N_VGND_c_1440_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_98 VNB N_VGND_c_1441_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_99 VNB N_VGND_c_1442_n 0.0190399f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.315
cc_100 VNB N_VGND_c_1443_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_101 VNB N_VGND_c_1444_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1445_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.645
cc_103 VNB N_VGND_c_1446_n 0.0922026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1447_n 0.0387696f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.48
cc_105 VNB N_VGND_c_1448_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=6.555 $Y2=1.56
cc_106 VNB N_VGND_c_1449_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=8.365 $Y2=2.4
cc_107 VNB N_VGND_c_1450_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=8.45 $Y2=1.815
cc_108 VNB N_VGND_c_1451_n 0.458857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VPB N_A_84_21#_M1006_g 0.0273379f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_110 VPB N_A_84_21#_M1011_g 0.0195468f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_111 VPB N_A_84_21#_M1016_g 0.0195863f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_112 VPB N_A_84_21#_M1021_g 0.0196107f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_113 VPB N_A_84_21#_M1022_g 0.0196107f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.465
cc_114 VPB N_A_84_21#_M1024_g 0.0196107f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_115 VPB N_A_84_21#_M1035_g 0.0196107f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=2.465
cc_116 VPB N_A_84_21#_M1036_g 0.0200687f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=2.465
cc_117 VPB N_A_84_21#_c_219_n 0.00103903f $X=-0.19 $Y=1.655 $X2=6.64 $Y2=2.025
cc_118 VPB N_A_84_21#_c_220_n 0.00929231f $X=-0.19 $Y=1.655 $X2=7.495 $Y2=2.11
cc_119 VPB N_A_84_21#_c_221_n 0.00686109f $X=-0.19 $Y=1.655 $X2=8.365 $Y2=2.4
cc_120 VPB N_A_84_21#_c_222_n 0.0139846f $X=-0.19 $Y=1.655 $X2=7.58 $Y2=2.11
cc_121 VPB N_A_84_21#_c_223_n 0.00446747f $X=-0.19 $Y=1.655 $X2=8.86 $Y2=1.98
cc_122 VPB N_A_84_21#_c_209_n 0.00262201f $X=-0.19 $Y=1.655 $X2=8.695 $Y2=1.815
cc_123 VPB N_A_772_21#_c_497_n 0.00288909f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=2.465
cc_124 VPB N_A_772_21#_c_498_n 0.0037317f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=2.465
cc_125 VPB N_A_772_21#_c_499_n 0.00819292f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=2.465
cc_126 VPB N_TE_B_c_664_n 0.0160123f $X=-0.19 $Y=1.655 $X2=8.72 $Y2=0.235
cc_127 VPB N_TE_B_c_645_n 0.00421372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_TE_B_c_646_n 0.00251798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_TE_B_c_667_n 0.0159999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_TE_B_c_647_n 0.00421299f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.655
cc_131 VPB N_TE_B_c_669_n 0.0159999f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.645
cc_132 VPB N_TE_B_c_648_n 0.00421372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_TE_B_c_671_n 0.0159999f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_134 VPB N_TE_B_c_649_n 0.00421299f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.645
cc_135 VPB N_TE_B_c_673_n 0.0159999f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_136 VPB N_TE_B_c_650_n 0.00421372f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=0.655
cc_137 VPB N_TE_B_c_675_n 0.0159929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_TE_B_c_651_n 0.00421299f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_139 VPB N_TE_B_c_677_n 0.0155272f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=1.315
cc_140 VPB N_TE_B_c_652_n 0.00466425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_TE_B_c_679_n 0.0197687f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_142 VPB N_TE_B_c_653_n 0.0264317f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=1.315
cc_143 VPB N_TE_B_c_654_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=1.315
cc_144 VPB N_TE_B_c_655_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=0.655
cc_145 VPB N_TE_B_c_656_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=0.655
cc_146 VPB N_TE_B_c_657_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_TE_B_c_658_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=1.645
cc_148 VPB N_TE_B_c_659_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_149 VPB N_TE_B_c_660_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_150 VPB N_TE_B_c_661_n 0.00981938f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=0.655
cc_151 VPB N_TE_B_c_689_n 0.0199981f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=2.465
cc_152 VPB N_A_M1019_g 0.0198764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_M1033_g 0.0271713f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_154 VPB N_A_27_367#_c_880_n 0.00719502f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_155 VPB N_A_27_367#_c_881_n 0.0457612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_27_367#_c_882_n 0.00172881f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_157 VPB N_A_27_367#_c_883_n 0.00235654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_27_367#_c_884_n 0.00186047f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=2.465
cc_159 VPB N_A_27_367#_c_885_n 0.00186047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_27_367#_c_886_n 0.00162958f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=2.465
cc_161 VPB N_A_27_367#_c_887_n 0.0019013f $X=-0.19 $Y=1.655 $X2=8.86 $Y2=0.42
cc_162 VPB N_A_27_367#_c_888_n 0.0019013f $X=-0.19 $Y=1.655 $X2=8.86 $Y2=2.485
cc_163 VPB N_A_27_367#_c_889_n 0.0240327f $X=-0.19 $Y=1.655 $X2=3.3 $Y2=1.48
cc_164 VPB N_Z_c_1018_n 0.00288801f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_Z_c_1019_n 0.003467f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=0.655
cc_166 VPB N_Z_c_1020_n 0.00225436f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.465
cc_167 VPB N_Z_c_1021_n 0.00225436f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=1.315
cc_168 VPB N_Z_c_1022_n 0.00230427f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=1.645
cc_169 VPB N_Z_c_1023_n 0.00230427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_Z_c_1024_n 0.00230427f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=1.48
cc_171 VPB N_VPWR_c_1148_n 0.00238736f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_172 VPB N_VPWR_c_1149_n 0.0047158f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=0.655
cc_173 VPB N_VPWR_c_1150_n 0.00412866f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_174 VPB N_VPWR_c_1151_n 0.00231123f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=0.655
cc_175 VPB N_VPWR_c_1152_n 0.00238736f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_176 VPB N_VPWR_c_1153_n 0.0116091f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=1.315
cc_177 VPB N_VPWR_c_1154_n 0.062339f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=0.655
cc_178 VPB N_VPWR_c_1155_n 0.0185788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1156_n 0.00324402f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=1.315
cc_180 VPB N_VPWR_c_1157_n 0.0185788f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=0.655
cc_181 VPB N_VPWR_c_1158_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1159_n 0.0158404f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_183 VPB N_VPWR_c_1160_n 0.00357074f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_184 VPB N_VPWR_c_1161_n 0.0921713f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=0.655
cc_185 VPB N_VPWR_c_1162_n 0.0418183f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=1.48
cc_186 VPB N_VPWR_c_1163_n 0.0185788f $X=-0.19 $Y=1.655 $X2=6.725 $Y2=2.11
cc_187 VPB N_VPWR_c_1164_n 0.00356964f $X=-0.19 $Y=1.655 $X2=8.86 $Y2=0.42
cc_188 VPB N_VPWR_c_1165_n 0.00356964f $X=-0.19 $Y=1.655 $X2=8.86 $Y2=2.485
cc_189 VPB N_VPWR_c_1147_n 0.0605132f $X=-0.19 $Y=1.655 $X2=3.3 $Y2=1.48
cc_190 N_A_84_21#_c_221_n N_A_772_21#_M1012_s 0.00782136f $X=8.365 $Y=2.4 $X2=0
+ $Y2=0
cc_191 N_A_84_21#_M1031_g N_A_772_21#_c_468_n 0.0106849f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_192 N_A_84_21#_c_208_n N_A_772_21#_c_470_n 0.0173052f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_193 N_A_84_21#_c_210_n N_A_772_21#_c_470_n 0.0106849f $X=3.505 $Y=1.48 $X2=0
+ $Y2=0
cc_194 N_A_84_21#_c_220_n N_A_772_21#_c_482_n 5.47511e-19 $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_195 N_A_84_21#_c_220_n N_A_772_21#_c_484_n 8.83737e-19 $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_196 N_A_84_21#_c_208_n N_A_772_21#_c_491_n 0.00123744f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_197 N_A_84_21#_c_220_n N_A_772_21#_c_492_n 5.05532e-19 $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_198 N_A_84_21#_c_221_n N_A_772_21#_c_497_n 0.00643308f $X=8.365 $Y=2.4 $X2=0
+ $Y2=0
cc_199 N_A_84_21#_c_222_n N_A_772_21#_c_497_n 0.00233413f $X=7.58 $Y=2.11 $X2=0
+ $Y2=0
cc_200 N_A_84_21#_c_220_n N_A_772_21#_c_498_n 0.00675638f $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_201 N_A_84_21#_c_222_n N_A_772_21#_c_498_n 0.0126514f $X=7.58 $Y=2.11 $X2=0
+ $Y2=0
cc_202 N_A_84_21#_c_237_p N_A_772_21#_c_495_n 0.0128586f $X=8.86 $Y=0.84 $X2=0
+ $Y2=0
cc_203 N_A_84_21#_c_238_p N_A_772_21#_c_495_n 0.00532173f $X=8.86 $Y=0.42 $X2=0
+ $Y2=0
cc_204 N_A_84_21#_c_221_n N_A_772_21#_c_499_n 0.0212577f $X=8.365 $Y=2.4 $X2=0
+ $Y2=0
cc_205 N_A_84_21#_c_222_n N_A_772_21#_c_499_n 0.00951416f $X=7.58 $Y=2.11 $X2=0
+ $Y2=0
cc_206 N_A_84_21#_c_209_n N_A_772_21#_c_499_n 0.0324943f $X=8.695 $Y=1.815 $X2=0
+ $Y2=0
cc_207 N_A_84_21#_M1036_g N_TE_B_c_664_n 0.0124689f $X=3.505 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_208 N_A_84_21#_c_208_n N_TE_B_c_645_n 0.00638796f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_209 N_A_84_21#_c_208_n N_TE_B_c_646_n 0.00461801f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_210 N_A_84_21#_c_210_n N_TE_B_c_646_n 0.0124689f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_211 N_A_84_21#_c_208_n N_TE_B_c_647_n 0.00637806f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_212 N_A_84_21#_c_208_n N_TE_B_c_648_n 0.00638796f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_213 N_A_84_21#_c_208_n N_TE_B_c_649_n 0.00637806f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_214 N_A_84_21#_c_208_n N_TE_B_c_650_n 0.00638796f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_215 N_A_84_21#_c_219_n N_TE_B_c_675_n 5.17212e-19 $X=6.64 $Y=2.025 $X2=0
+ $Y2=0
cc_216 N_A_84_21#_c_208_n N_TE_B_c_651_n 0.00802952f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_217 N_A_84_21#_c_219_n N_TE_B_c_677_n 0.00594207f $X=6.64 $Y=2.025 $X2=0
+ $Y2=0
cc_218 N_A_84_21#_c_253_p N_TE_B_c_677_n 0.00438212f $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_219 N_A_84_21#_c_208_n N_TE_B_c_652_n 0.0052046f $X=6.555 $Y=1.56 $X2=0 $Y2=0
cc_220 N_A_84_21#_c_219_n N_TE_B_c_652_n 0.00546227f $X=6.64 $Y=2.025 $X2=0
+ $Y2=0
cc_221 N_A_84_21#_c_220_n N_TE_B_c_652_n 0.00162374f $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_222 N_A_84_21#_c_219_n N_TE_B_c_679_n 0.00637569f $X=6.64 $Y=2.025 $X2=0
+ $Y2=0
cc_223 N_A_84_21#_c_220_n N_TE_B_c_679_n 0.0132484f $X=7.495 $Y=2.11 $X2=0 $Y2=0
cc_224 N_A_84_21#_c_222_n N_TE_B_c_679_n 0.00429029f $X=7.58 $Y=2.11 $X2=0 $Y2=0
cc_225 N_A_84_21#_c_220_n N_TE_B_c_653_n 0.00950068f $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_226 N_A_84_21#_c_221_n N_TE_B_c_653_n 0.00140449f $X=8.365 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_84_21#_c_222_n N_TE_B_c_653_n 9.51866e-19 $X=7.58 $Y=2.11 $X2=0 $Y2=0
cc_228 N_A_84_21#_c_208_n N_TE_B_c_654_n 0.00379186f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_229 N_A_84_21#_c_208_n N_TE_B_c_655_n 0.00379186f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_230 N_A_84_21#_c_208_n N_TE_B_c_656_n 0.00379186f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_231 N_A_84_21#_c_208_n N_TE_B_c_657_n 0.00379186f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_232 N_A_84_21#_c_208_n N_TE_B_c_658_n 0.00379186f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_233 N_A_84_21#_c_208_n N_TE_B_c_659_n 0.00677453f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_234 N_A_84_21#_c_219_n N_TE_B_c_659_n 0.00374706f $X=6.64 $Y=2.025 $X2=0
+ $Y2=0
cc_235 N_A_84_21#_c_223_n N_TE_B_c_661_n 0.00984425f $X=8.86 $Y=1.98 $X2=0 $Y2=0
cc_236 N_A_84_21#_c_209_n N_TE_B_c_662_n 0.0254324f $X=8.695 $Y=1.815 $X2=0
+ $Y2=0
cc_237 N_A_84_21#_c_237_p N_TE_B_c_663_n 0.00138727f $X=8.86 $Y=0.84 $X2=0 $Y2=0
cc_238 N_A_84_21#_c_238_p N_TE_B_c_663_n 6.24294e-19 $X=8.86 $Y=0.42 $X2=0 $Y2=0
cc_239 N_A_84_21#_c_209_n N_TE_B_c_663_n 0.00984425f $X=8.695 $Y=1.815 $X2=0
+ $Y2=0
cc_240 N_A_84_21#_c_221_n N_TE_B_c_689_n 0.0162905f $X=8.365 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A_84_21#_c_276_p N_TE_B_c_689_n 9.67478e-19 $X=8.86 $Y=2.91 $X2=0 $Y2=0
cc_242 N_A_84_21#_c_222_n N_TE_B_c_689_n 0.00429029f $X=7.58 $Y=2.11 $X2=0 $Y2=0
cc_243 N_A_84_21#_c_223_n N_TE_B_c_689_n 2.82164e-19 $X=8.86 $Y=1.98 $X2=0 $Y2=0
cc_244 N_A_84_21#_c_237_p N_A_c_841_n 0.01311f $X=8.86 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_245 N_A_84_21#_c_238_p N_A_c_841_n 0.00794586f $X=8.86 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_246 N_A_84_21#_c_209_n N_A_c_841_n 0.0129084f $X=8.695 $Y=1.815 $X2=-0.19
+ $Y2=-0.245
cc_247 N_A_84_21#_c_276_p N_A_M1019_g 0.00852789f $X=8.86 $Y=2.91 $X2=0 $Y2=0
cc_248 N_A_84_21#_c_223_n N_A_M1019_g 0.0271786f $X=8.86 $Y=1.98 $X2=0 $Y2=0
cc_249 N_A_84_21#_c_237_p N_A_c_843_n 0.00224022f $X=8.86 $Y=0.84 $X2=0 $Y2=0
cc_250 N_A_84_21#_c_238_p N_A_c_843_n 0.00707388f $X=8.86 $Y=0.42 $X2=0 $Y2=0
cc_251 N_A_84_21#_c_276_p N_A_M1033_g 0.00752654f $X=8.86 $Y=2.91 $X2=0 $Y2=0
cc_252 N_A_84_21#_c_223_n N_A_M1033_g 0.00888948f $X=8.86 $Y=1.98 $X2=0 $Y2=0
cc_253 N_A_84_21#_c_237_p A 0.0205336f $X=8.86 $Y=0.84 $X2=0 $Y2=0
cc_254 N_A_84_21#_c_223_n A 0.0174707f $X=8.86 $Y=1.98 $X2=0 $Y2=0
cc_255 N_A_84_21#_c_209_n A 0.0251362f $X=8.695 $Y=1.815 $X2=0 $Y2=0
cc_256 N_A_84_21#_c_237_p N_A_c_846_n 6.94598e-19 $X=8.86 $Y=0.84 $X2=0 $Y2=0
cc_257 N_A_84_21#_c_223_n N_A_c_846_n 7.38095e-19 $X=8.86 $Y=1.98 $X2=0 $Y2=0
cc_258 N_A_84_21#_c_220_n N_A_27_367#_M1034_s 0.00650122f $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_259 N_A_84_21#_M1006_g N_A_27_367#_c_880_n 5.89773e-19 $X=0.495 $Y=2.465
+ $X2=0 $Y2=0
cc_260 N_A_84_21#_M1006_g N_A_27_367#_c_881_n 0.0164264f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_261 N_A_84_21#_M1011_g N_A_27_367#_c_881_n 7.17462e-19 $X=0.925 $Y=2.465
+ $X2=0 $Y2=0
cc_262 N_A_84_21#_M1006_g N_A_27_367#_c_894_n 0.0105205f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_263 N_A_84_21#_M1011_g N_A_27_367#_c_894_n 0.0105205f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A_84_21#_M1006_g N_A_27_367#_c_896_n 6.10078e-19 $X=0.495 $Y=2.465
+ $X2=0 $Y2=0
cc_265 N_A_84_21#_M1011_g N_A_27_367#_c_896_n 0.0111058f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_266 N_A_84_21#_M1016_g N_A_27_367#_c_898_n 0.0115031f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_267 N_A_84_21#_M1021_g N_A_27_367#_c_898_n 0.0115031f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_268 N_A_84_21#_M1022_g N_A_27_367#_c_900_n 0.0115031f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_269 N_A_84_21#_M1024_g N_A_27_367#_c_900_n 0.0115031f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_A_84_21#_M1035_g N_A_27_367#_c_902_n 0.0114565f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_84_21#_M1036_g N_A_27_367#_c_902_n 0.0115031f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_272 N_A_84_21#_c_208_n N_A_27_367#_c_882_n 0.0143583f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_273 N_A_84_21#_c_208_n N_A_27_367#_c_883_n 0.0426707f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_274 N_A_84_21#_c_208_n N_A_27_367#_c_884_n 0.0368384f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_275 N_A_84_21#_c_208_n N_A_27_367#_c_885_n 0.0368384f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_276 N_A_84_21#_c_208_n N_A_27_367#_c_886_n 0.0200256f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_277 N_A_84_21#_c_219_n N_A_27_367#_c_886_n 0.00667447f $X=6.64 $Y=2.025 $X2=0
+ $Y2=0
cc_278 N_A_84_21#_c_220_n N_A_27_367#_c_910_n 0.0147941f $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_279 N_A_84_21#_c_253_p N_A_27_367#_c_910_n 0.00896703f $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_280 N_A_84_21#_M1011_g N_A_27_367#_c_912_n 5.89773e-19 $X=0.925 $Y=2.465
+ $X2=0 $Y2=0
cc_281 N_A_84_21#_c_208_n N_A_27_367#_c_887_n 0.0263346f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_282 N_A_84_21#_c_208_n N_A_27_367#_c_888_n 0.0263346f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_283 N_A_84_21#_c_220_n N_A_27_367#_c_889_n 0.0221791f $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_284 N_A_84_21#_c_222_n N_A_27_367#_c_889_n 0.0101352f $X=7.58 $Y=2.11 $X2=0
+ $Y2=0
cc_285 N_A_84_21#_M1003_g N_Z_c_1025_n 0.00465849f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_286 N_A_84_21#_M1005_g N_Z_c_1025_n 0.00563901f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_287 N_A_84_21#_M1009_g N_Z_c_1025_n 5.62335e-19 $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_288 N_A_84_21#_M1003_g N_Z_c_1011_n 0.0119611f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_289 N_A_84_21#_M1005_g N_Z_c_1011_n 0.00825926f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_290 N_A_84_21#_c_325_p N_Z_c_1011_n 0.0056664f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_291 N_A_84_21#_c_210_n N_Z_c_1011_n 0.0117416f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_292 N_A_84_21#_M1006_g N_Z_c_1018_n 0.00403324f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A_84_21#_M1011_g N_Z_c_1018_n 0.00403324f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A_84_21#_c_325_p N_Z_c_1018_n 0.0112733f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_295 N_A_84_21#_c_210_n N_Z_c_1018_n 0.0196292f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_296 N_A_84_21#_M1011_g N_Z_c_1019_n 0.0146489f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A_84_21#_M1016_g N_Z_c_1019_n 0.0111034f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A_84_21#_c_325_p N_Z_c_1019_n 0.0227981f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_299 N_A_84_21#_c_210_n N_Z_c_1019_n 0.00226668f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_300 N_A_84_21#_M1005_g N_Z_c_1012_n 0.0107261f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_301 N_A_84_21#_M1009_g N_Z_c_1012_n 0.00889811f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_302 N_A_84_21#_c_325_p N_Z_c_1012_n 0.0227981f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_303 N_A_84_21#_c_210_n N_Z_c_1012_n 0.00226668f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_304 N_A_84_21#_M1005_g N_Z_c_1044_n 5.62335e-19 $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_305 N_A_84_21#_M1009_g N_Z_c_1044_n 0.00563901f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_306 N_A_84_21#_M1010_g N_Z_c_1044_n 0.00563901f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_307 N_A_84_21#_M1017_g N_Z_c_1044_n 5.62335e-19 $X=2.215 $Y=0.655 $X2=0 $Y2=0
cc_308 N_A_84_21#_M1010_g N_Z_c_1013_n 0.00889811f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_309 N_A_84_21#_M1017_g N_Z_c_1013_n 0.00889811f $X=2.215 $Y=0.655 $X2=0 $Y2=0
cc_310 N_A_84_21#_c_325_p N_Z_c_1013_n 0.0388321f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_311 N_A_84_21#_c_210_n N_Z_c_1013_n 0.00224206f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_312 N_A_84_21#_M1021_g N_Z_c_1020_n 0.01115f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_313 N_A_84_21#_M1022_g N_Z_c_1020_n 0.01115f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A_84_21#_c_325_p N_Z_c_1020_n 0.0388321f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_315 N_A_84_21#_c_210_n N_Z_c_1020_n 0.00224206f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_316 N_A_84_21#_M1010_g N_Z_c_1056_n 5.62335e-19 $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_317 N_A_84_21#_M1017_g N_Z_c_1056_n 0.00563901f $X=2.215 $Y=0.655 $X2=0 $Y2=0
cc_318 N_A_84_21#_M1025_g N_Z_c_1056_n 0.00563901f $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_319 N_A_84_21#_M1028_g N_Z_c_1056_n 5.62335e-19 $X=3.075 $Y=0.655 $X2=0 $Y2=0
cc_320 N_A_84_21#_M1025_g N_Z_c_1014_n 0.00889811f $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_321 N_A_84_21#_M1028_g N_Z_c_1014_n 0.0113726f $X=3.075 $Y=0.655 $X2=0 $Y2=0
cc_322 N_A_84_21#_M1031_g N_Z_c_1014_n 0.00384654f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_323 N_A_84_21#_c_325_p N_Z_c_1014_n 0.0659283f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_324 N_A_84_21#_c_210_n N_Z_c_1014_n 0.00455346f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_325 N_A_84_21#_M1024_g N_Z_c_1021_n 0.01115f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_326 N_A_84_21#_M1035_g N_Z_c_1021_n 0.01115f $X=3.075 $Y=2.465 $X2=0 $Y2=0
cc_327 N_A_84_21#_c_325_p N_Z_c_1021_n 0.0388321f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_328 N_A_84_21#_c_210_n N_Z_c_1021_n 0.00224206f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_329 N_A_84_21#_M1025_g N_Z_c_1069_n 5.62335e-19 $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_330 N_A_84_21#_M1028_g N_Z_c_1069_n 0.00563901f $X=3.075 $Y=0.655 $X2=0 $Y2=0
cc_331 N_A_84_21#_M1031_g N_Z_c_1069_n 0.00443684f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_332 N_A_84_21#_M1009_g N_Z_c_1015_n 0.00247446f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_333 N_A_84_21#_M1010_g N_Z_c_1015_n 0.00247446f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_334 N_A_84_21#_c_325_p N_Z_c_1015_n 0.0271338f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_335 N_A_84_21#_c_210_n N_Z_c_1015_n 0.00231141f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_336 N_A_84_21#_M1011_g N_Z_c_1022_n 7.15041e-19 $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_337 N_A_84_21#_M1016_g N_Z_c_1022_n 0.0128652f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_338 N_A_84_21#_M1021_g N_Z_c_1022_n 0.0126541f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_339 N_A_84_21#_M1022_g N_Z_c_1022_n 6.07933e-19 $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_340 N_A_84_21#_c_325_p N_Z_c_1022_n 0.0276081f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_341 N_A_84_21#_c_210_n N_Z_c_1022_n 0.00232957f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_342 N_A_84_21#_M1017_g N_Z_c_1016_n 0.00247446f $X=2.215 $Y=0.655 $X2=0 $Y2=0
cc_343 N_A_84_21#_M1025_g N_Z_c_1016_n 0.00247446f $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_344 N_A_84_21#_c_325_p N_Z_c_1016_n 0.0271338f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_345 N_A_84_21#_c_210_n N_Z_c_1016_n 0.00231141f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_346 N_A_84_21#_M1021_g N_Z_c_1023_n 6.07933e-19 $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_347 N_A_84_21#_M1022_g N_Z_c_1023_n 0.0126541f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_348 N_A_84_21#_M1024_g N_Z_c_1023_n 0.0126541f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_349 N_A_84_21#_M1035_g N_Z_c_1023_n 6.07933e-19 $X=3.075 $Y=2.465 $X2=0 $Y2=0
cc_350 N_A_84_21#_c_325_p N_Z_c_1023_n 0.0276081f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_351 N_A_84_21#_c_210_n N_Z_c_1023_n 0.00232957f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_352 N_A_84_21#_M1024_g N_Z_c_1024_n 6.07933e-19 $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_353 N_A_84_21#_M1035_g N_Z_c_1024_n 0.0126541f $X=3.075 $Y=2.465 $X2=0 $Y2=0
cc_354 N_A_84_21#_M1036_g N_Z_c_1024_n 0.0128123f $X=3.505 $Y=2.465 $X2=0 $Y2=0
cc_355 N_A_84_21#_c_325_p N_Z_c_1024_n 0.0275704f $X=3.3 $Y=1.48 $X2=0 $Y2=0
cc_356 N_A_84_21#_c_210_n N_Z_c_1024_n 0.00232957f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_357 N_A_84_21#_M1003_g N_Z_c_1017_n 0.00989921f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_358 N_A_84_21#_c_210_n N_Z_c_1017_n 0.00809811f $X=3.505 $Y=1.48 $X2=0 $Y2=0
cc_359 N_A_84_21#_c_219_n N_VPWR_M1030_d 0.00215798f $X=6.64 $Y=2.025 $X2=0
+ $Y2=0
cc_360 N_A_84_21#_c_220_n N_VPWR_M1030_d 0.00221499f $X=7.495 $Y=2.11 $X2=0
+ $Y2=0
cc_361 N_A_84_21#_c_253_p N_VPWR_M1030_d 8.55688e-19 $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_362 N_A_84_21#_c_221_n N_VPWR_M1012_d 0.00128614f $X=8.365 $Y=2.4 $X2=0 $Y2=0
cc_363 N_A_84_21#_c_223_n N_VPWR_M1012_d 0.00743519f $X=8.86 $Y=1.98 $X2=0 $Y2=0
cc_364 N_A_84_21#_M1036_g N_VPWR_c_1148_n 0.00107091f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_A_84_21#_c_221_n N_VPWR_c_1152_n 0.003222f $X=8.365 $Y=2.4 $X2=0 $Y2=0
cc_366 N_A_84_21#_c_223_n N_VPWR_c_1152_n 0.0129405f $X=8.86 $Y=1.98 $X2=0 $Y2=0
cc_367 N_A_84_21#_c_223_n N_VPWR_c_1154_n 0.0485359f $X=8.86 $Y=1.98 $X2=0 $Y2=0
cc_368 N_A_84_21#_M1006_g N_VPWR_c_1161_n 0.00357842f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_369 N_A_84_21#_M1011_g N_VPWR_c_1161_n 0.00357842f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_370 N_A_84_21#_M1016_g N_VPWR_c_1161_n 0.00357877f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_371 N_A_84_21#_M1021_g N_VPWR_c_1161_n 0.00357877f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_372 N_A_84_21#_M1022_g N_VPWR_c_1161_n 0.00357877f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_373 N_A_84_21#_M1024_g N_VPWR_c_1161_n 0.00357877f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_374 N_A_84_21#_M1035_g N_VPWR_c_1161_n 0.00357877f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_375 N_A_84_21#_M1036_g N_VPWR_c_1161_n 0.00357877f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_376 N_A_84_21#_c_276_p N_VPWR_c_1163_n 0.0189236f $X=8.86 $Y=2.91 $X2=0 $Y2=0
cc_377 N_A_84_21#_M1019_s N_VPWR_c_1147_n 0.00223559f $X=8.72 $Y=1.835 $X2=0
+ $Y2=0
cc_378 N_A_84_21#_M1006_g N_VPWR_c_1147_n 0.00630218f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_379 N_A_84_21#_M1011_g N_VPWR_c_1147_n 0.00535118f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_380 N_A_84_21#_M1016_g N_VPWR_c_1147_n 0.0053512f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_381 N_A_84_21#_M1021_g N_VPWR_c_1147_n 0.0053512f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_382 N_A_84_21#_M1022_g N_VPWR_c_1147_n 0.0053512f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_383 N_A_84_21#_M1024_g N_VPWR_c_1147_n 0.0053512f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_384 N_A_84_21#_M1035_g N_VPWR_c_1147_n 0.0053512f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_385 N_A_84_21#_M1036_g N_VPWR_c_1147_n 0.00537654f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_386 N_A_84_21#_c_221_n N_VPWR_c_1147_n 0.0200838f $X=8.365 $Y=2.4 $X2=0 $Y2=0
cc_387 N_A_84_21#_c_276_p N_VPWR_c_1147_n 0.0123859f $X=8.86 $Y=2.91 $X2=0 $Y2=0
cc_388 N_A_84_21#_c_222_n N_VPWR_c_1147_n 0.00634627f $X=7.58 $Y=2.11 $X2=0
+ $Y2=0
cc_389 N_A_84_21#_c_223_n N_VPWR_c_1147_n 0.00663174f $X=8.86 $Y=1.98 $X2=0
+ $Y2=0
cc_390 N_A_84_21#_M1003_g N_A_27_47#_c_1289_n 0.0115031f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_391 N_A_84_21#_M1005_g N_A_27_47#_c_1289_n 0.0101666f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_392 N_A_84_21#_M1009_g N_A_27_47#_c_1291_n 0.0101666f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_393 N_A_84_21#_M1010_g N_A_27_47#_c_1291_n 0.0101666f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_394 N_A_84_21#_M1017_g N_A_27_47#_c_1293_n 0.0101666f $X=2.215 $Y=0.655 $X2=0
+ $Y2=0
cc_395 N_A_84_21#_M1025_g N_A_27_47#_c_1293_n 0.0101666f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_396 N_A_84_21#_M1028_g N_A_27_47#_c_1295_n 0.01012f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_397 N_A_84_21#_M1031_g N_A_27_47#_c_1295_n 0.0115031f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_398 N_A_84_21#_M1031_g N_A_27_47#_c_1281_n 9.26489e-19 $X=3.505 $Y=0.655
+ $X2=0 $Y2=0
cc_399 N_A_84_21#_c_208_n N_A_27_47#_c_1282_n 0.0436966f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_400 N_A_84_21#_M1031_g N_A_27_47#_c_1283_n 0.00514561f $X=3.505 $Y=0.655
+ $X2=0 $Y2=0
cc_401 N_A_84_21#_c_208_n N_A_27_47#_c_1283_n 0.0143583f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_402 N_A_84_21#_c_208_n N_A_27_47#_c_1284_n 0.0377708f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_403 N_A_84_21#_c_208_n N_A_27_47#_c_1285_n 0.0377708f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_404 N_A_84_21#_c_208_n N_A_27_47#_c_1286_n 0.0201154f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_405 N_A_84_21#_c_208_n N_A_27_47#_c_1304_n 0.026287f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_406 N_A_84_21#_c_208_n N_A_27_47#_c_1305_n 0.026287f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_407 N_A_84_21#_c_208_n N_A_27_47#_c_1306_n 0.026287f $X=6.555 $Y=1.56 $X2=0
+ $Y2=0
cc_408 N_A_84_21#_c_237_p N_VGND_M1020_d 0.00373324f $X=8.86 $Y=0.84 $X2=0 $Y2=0
cc_409 N_A_84_21#_c_209_n N_VGND_M1020_d 0.00120688f $X=8.695 $Y=1.815 $X2=0
+ $Y2=0
cc_410 N_A_84_21#_M1031_g N_VGND_c_1433_n 0.00107091f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_411 N_A_84_21#_c_237_p N_VGND_c_1437_n 0.0117772f $X=8.86 $Y=0.84 $X2=0 $Y2=0
cc_412 N_A_84_21#_c_209_n N_VGND_c_1439_n 5.53166e-19 $X=8.695 $Y=1.815 $X2=0
+ $Y2=0
cc_413 N_A_84_21#_M1003_g N_VGND_c_1446_n 0.00357877f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_414 N_A_84_21#_M1005_g N_VGND_c_1446_n 0.00357877f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_415 N_A_84_21#_M1009_g N_VGND_c_1446_n 0.00357877f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_416 N_A_84_21#_M1010_g N_VGND_c_1446_n 0.00357877f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_417 N_A_84_21#_M1017_g N_VGND_c_1446_n 0.00357877f $X=2.215 $Y=0.655 $X2=0
+ $Y2=0
cc_418 N_A_84_21#_M1025_g N_VGND_c_1446_n 0.00357877f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_419 N_A_84_21#_M1028_g N_VGND_c_1446_n 0.00357877f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_420 N_A_84_21#_M1031_g N_VGND_c_1446_n 0.00357877f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_421 N_A_84_21#_c_238_p N_VGND_c_1448_n 0.018762f $X=8.86 $Y=0.42 $X2=0 $Y2=0
cc_422 N_A_84_21#_M1008_s N_VGND_c_1451_n 0.00223559f $X=8.72 $Y=0.235 $X2=0
+ $Y2=0
cc_423 N_A_84_21#_M1003_g N_VGND_c_1451_n 0.0063022f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_424 N_A_84_21#_M1005_g N_VGND_c_1451_n 0.00542194f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_425 N_A_84_21#_M1009_g N_VGND_c_1451_n 0.00542194f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_426 N_A_84_21#_M1010_g N_VGND_c_1451_n 0.00542194f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_427 N_A_84_21#_M1017_g N_VGND_c_1451_n 0.00542194f $X=2.215 $Y=0.655 $X2=0
+ $Y2=0
cc_428 N_A_84_21#_M1025_g N_VGND_c_1451_n 0.00542194f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_429 N_A_84_21#_M1028_g N_VGND_c_1451_n 0.00542194f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_430 N_A_84_21#_M1031_g N_VGND_c_1451_n 0.00537654f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_431 N_A_84_21#_c_237_p N_VGND_c_1451_n 0.00582163f $X=8.86 $Y=0.84 $X2=0
+ $Y2=0
cc_432 N_A_84_21#_c_238_p N_VGND_c_1451_n 0.0123366f $X=8.86 $Y=0.42 $X2=0 $Y2=0
cc_433 N_A_772_21#_c_469_n N_TE_B_c_645_n 0.0127375f $X=4.29 $Y=1.26 $X2=0 $Y2=0
cc_434 N_A_772_21#_c_470_n N_TE_B_c_646_n 0.0127375f $X=4.01 $Y=1.26 $X2=0 $Y2=0
cc_435 N_A_772_21#_c_472_n N_TE_B_c_647_n 0.0127375f $X=4.72 $Y=1.26 $X2=0 $Y2=0
cc_436 N_A_772_21#_c_474_n N_TE_B_c_648_n 0.0127375f $X=5.15 $Y=1.26 $X2=0 $Y2=0
cc_437 N_A_772_21#_c_476_n N_TE_B_c_649_n 0.0127375f $X=5.58 $Y=1.26 $X2=0 $Y2=0
cc_438 N_A_772_21#_c_478_n N_TE_B_c_650_n 0.0127375f $X=6.01 $Y=1.26 $X2=0 $Y2=0
cc_439 N_A_772_21#_c_480_n N_TE_B_c_651_n 0.0127375f $X=6.44 $Y=1.26 $X2=0 $Y2=0
cc_440 N_A_772_21#_c_482_n N_TE_B_c_652_n 0.0127375f $X=6.87 $Y=1.26 $X2=0 $Y2=0
cc_441 N_A_772_21#_c_498_n N_TE_B_c_679_n 0.00391286f $X=7.635 $Y=1.77 $X2=0
+ $Y2=0
cc_442 N_A_772_21#_c_484_n N_TE_B_c_653_n 0.0127375f $X=7.415 $Y=1.26 $X2=0
+ $Y2=0
cc_443 N_A_772_21#_c_493_n N_TE_B_c_653_n 0.00216828f $X=7.58 $Y=0.925 $X2=0
+ $Y2=0
cc_444 N_A_772_21#_c_494_n N_TE_B_c_653_n 0.0149027f $X=7.525 $Y=1.685 $X2=0
+ $Y2=0
cc_445 N_A_772_21#_c_497_n N_TE_B_c_653_n 0.0079199f $X=7.835 $Y=1.77 $X2=0
+ $Y2=0
cc_446 N_A_772_21#_c_498_n N_TE_B_c_653_n 0.00645153f $X=7.635 $Y=1.77 $X2=0
+ $Y2=0
cc_447 N_A_772_21#_c_495_n N_TE_B_c_653_n 0.00201073f $X=7.58 $Y=0.42 $X2=0
+ $Y2=0
cc_448 N_A_772_21#_c_499_n N_TE_B_c_653_n 0.00106189f $X=8 $Y=1.77 $X2=0 $Y2=0
cc_449 N_A_772_21#_c_486_n N_TE_B_c_654_n 0.0127375f $X=4.365 $Y=1.26 $X2=0
+ $Y2=0
cc_450 N_A_772_21#_c_487_n N_TE_B_c_655_n 0.0127375f $X=4.795 $Y=1.26 $X2=0
+ $Y2=0
cc_451 N_A_772_21#_c_488_n N_TE_B_c_656_n 0.0127375f $X=5.225 $Y=1.26 $X2=0
+ $Y2=0
cc_452 N_A_772_21#_c_489_n N_TE_B_c_657_n 0.0127375f $X=5.655 $Y=1.26 $X2=0
+ $Y2=0
cc_453 N_A_772_21#_c_490_n N_TE_B_c_658_n 0.0127375f $X=6.085 $Y=1.26 $X2=0
+ $Y2=0
cc_454 N_A_772_21#_c_491_n N_TE_B_c_659_n 0.0127375f $X=6.515 $Y=1.26 $X2=0
+ $Y2=0
cc_455 N_A_772_21#_c_492_n N_TE_B_c_660_n 0.0127375f $X=6.945 $Y=1.26 $X2=0
+ $Y2=0
cc_456 N_A_772_21#_c_484_n N_TE_B_c_661_n 0.00626584f $X=7.415 $Y=1.26 $X2=0
+ $Y2=0
cc_457 N_A_772_21#_c_494_n N_TE_B_c_661_n 0.00379592f $X=7.525 $Y=1.685 $X2=0
+ $Y2=0
cc_458 N_A_772_21#_c_495_n N_TE_B_c_661_n 0.00195893f $X=7.58 $Y=0.42 $X2=0
+ $Y2=0
cc_459 N_A_772_21#_c_499_n N_TE_B_c_661_n 0.00975186f $X=8 $Y=1.77 $X2=0 $Y2=0
cc_460 N_A_772_21#_c_485_n N_TE_B_c_662_n 4.75143e-19 $X=7.49 $Y=1.185 $X2=0
+ $Y2=0
cc_461 N_A_772_21#_c_494_n N_TE_B_c_662_n 0.0273772f $X=7.525 $Y=1.685 $X2=0
+ $Y2=0
cc_462 N_A_772_21#_c_497_n N_TE_B_c_662_n 0.00226773f $X=7.835 $Y=1.77 $X2=0
+ $Y2=0
cc_463 N_A_772_21#_c_495_n N_TE_B_c_662_n 0.0284789f $X=7.58 $Y=0.42 $X2=0 $Y2=0
cc_464 N_A_772_21#_c_499_n N_TE_B_c_662_n 0.025492f $X=8 $Y=1.77 $X2=0 $Y2=0
cc_465 N_A_772_21#_c_485_n N_TE_B_c_663_n 0.00300863f $X=7.49 $Y=1.185 $X2=0
+ $Y2=0
cc_466 N_A_772_21#_c_494_n N_TE_B_c_663_n 0.00268624f $X=7.525 $Y=1.685 $X2=0
+ $Y2=0
cc_467 N_A_772_21#_c_495_n N_TE_B_c_663_n 0.0101337f $X=7.58 $Y=0.42 $X2=0 $Y2=0
cc_468 N_A_772_21#_c_496_n N_TE_B_c_663_n 0.00999764f $X=7.58 $Y=0.42 $X2=0
+ $Y2=0
cc_469 N_A_772_21#_c_497_n N_TE_B_c_689_n 3.75382e-19 $X=7.835 $Y=1.77 $X2=0
+ $Y2=0
cc_470 N_A_772_21#_c_499_n N_TE_B_c_689_n 0.00704156f $X=8 $Y=1.77 $X2=0 $Y2=0
cc_471 N_A_772_21#_c_495_n N_A_c_841_n 7.54362e-19 $X=7.58 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_472 N_A_772_21#_c_499_n N_A_M1019_g 2.58466e-19 $X=8 $Y=1.77 $X2=0 $Y2=0
cc_473 N_A_772_21#_M1012_s N_VPWR_c_1147_n 0.00423886f $X=7.855 $Y=1.835 $X2=0
+ $Y2=0
cc_474 N_A_772_21#_c_468_n N_A_27_47#_c_1281_n 0.00123476f $X=3.935 $Y=1.185
+ $X2=0 $Y2=0
cc_475 N_A_772_21#_c_468_n N_A_27_47#_c_1282_n 0.00758729f $X=3.935 $Y=1.185
+ $X2=0 $Y2=0
cc_476 N_A_772_21#_c_469_n N_A_27_47#_c_1282_n 0.00606528f $X=4.29 $Y=1.26 $X2=0
+ $Y2=0
cc_477 N_A_772_21#_c_470_n N_A_27_47#_c_1282_n 0.00354297f $X=4.01 $Y=1.26 $X2=0
+ $Y2=0
cc_478 N_A_772_21#_c_471_n N_A_27_47#_c_1282_n 0.00660493f $X=4.365 $Y=1.185
+ $X2=0 $Y2=0
cc_479 N_A_772_21#_c_486_n N_A_27_47#_c_1282_n 0.00203622f $X=4.365 $Y=1.26
+ $X2=0 $Y2=0
cc_480 N_A_772_21#_c_468_n N_A_27_47#_c_1313_n 6.7664e-19 $X=3.935 $Y=1.185
+ $X2=0 $Y2=0
cc_481 N_A_772_21#_c_471_n N_A_27_47#_c_1313_n 0.0128372f $X=4.365 $Y=1.185
+ $X2=0 $Y2=0
cc_482 N_A_772_21#_c_473_n N_A_27_47#_c_1313_n 0.0126262f $X=4.795 $Y=1.185
+ $X2=0 $Y2=0
cc_483 N_A_772_21#_c_475_n N_A_27_47#_c_1313_n 6.46727e-19 $X=5.225 $Y=1.185
+ $X2=0 $Y2=0
cc_484 N_A_772_21#_c_473_n N_A_27_47#_c_1284_n 0.00661824f $X=4.795 $Y=1.185
+ $X2=0 $Y2=0
cc_485 N_A_772_21#_c_474_n N_A_27_47#_c_1284_n 0.00606528f $X=5.15 $Y=1.26 $X2=0
+ $Y2=0
cc_486 N_A_772_21#_c_475_n N_A_27_47#_c_1284_n 0.00661824f $X=5.225 $Y=1.185
+ $X2=0 $Y2=0
cc_487 N_A_772_21#_c_487_n N_A_27_47#_c_1284_n 0.00203622f $X=4.795 $Y=1.26
+ $X2=0 $Y2=0
cc_488 N_A_772_21#_c_488_n N_A_27_47#_c_1284_n 0.00203622f $X=5.225 $Y=1.26
+ $X2=0 $Y2=0
cc_489 N_A_772_21#_c_473_n N_A_27_47#_c_1322_n 6.3479e-19 $X=4.795 $Y=1.185
+ $X2=0 $Y2=0
cc_490 N_A_772_21#_c_475_n N_A_27_47#_c_1322_n 0.0127355f $X=5.225 $Y=1.185
+ $X2=0 $Y2=0
cc_491 N_A_772_21#_c_477_n N_A_27_47#_c_1322_n 0.0127355f $X=5.655 $Y=1.185
+ $X2=0 $Y2=0
cc_492 N_A_772_21#_c_479_n N_A_27_47#_c_1322_n 6.3479e-19 $X=6.085 $Y=1.185
+ $X2=0 $Y2=0
cc_493 N_A_772_21#_c_477_n N_A_27_47#_c_1285_n 0.00661824f $X=5.655 $Y=1.185
+ $X2=0 $Y2=0
cc_494 N_A_772_21#_c_478_n N_A_27_47#_c_1285_n 0.00606528f $X=6.01 $Y=1.26 $X2=0
+ $Y2=0
cc_495 N_A_772_21#_c_479_n N_A_27_47#_c_1285_n 0.00661824f $X=6.085 $Y=1.185
+ $X2=0 $Y2=0
cc_496 N_A_772_21#_c_489_n N_A_27_47#_c_1285_n 0.00203622f $X=5.655 $Y=1.26
+ $X2=0 $Y2=0
cc_497 N_A_772_21#_c_490_n N_A_27_47#_c_1285_n 0.00203622f $X=6.085 $Y=1.26
+ $X2=0 $Y2=0
cc_498 N_A_772_21#_c_477_n N_A_27_47#_c_1331_n 6.46727e-19 $X=5.655 $Y=1.185
+ $X2=0 $Y2=0
cc_499 N_A_772_21#_c_479_n N_A_27_47#_c_1331_n 0.0126262f $X=6.085 $Y=1.185
+ $X2=0 $Y2=0
cc_500 N_A_772_21#_c_481_n N_A_27_47#_c_1331_n 0.0126262f $X=6.515 $Y=1.185
+ $X2=0 $Y2=0
cc_501 N_A_772_21#_c_483_n N_A_27_47#_c_1331_n 6.46727e-19 $X=6.945 $Y=1.185
+ $X2=0 $Y2=0
cc_502 N_A_772_21#_c_481_n N_A_27_47#_c_1286_n 0.00660493f $X=6.515 $Y=1.185
+ $X2=0 $Y2=0
cc_503 N_A_772_21#_c_482_n N_A_27_47#_c_1286_n 0.00715351f $X=6.87 $Y=1.26 $X2=0
+ $Y2=0
cc_504 N_A_772_21#_c_483_n N_A_27_47#_c_1286_n 0.00729562f $X=6.945 $Y=1.185
+ $X2=0 $Y2=0
cc_505 N_A_772_21#_c_484_n N_A_27_47#_c_1286_n 0.0108434f $X=7.415 $Y=1.26 $X2=0
+ $Y2=0
cc_506 N_A_772_21#_c_485_n N_A_27_47#_c_1286_n 3.73873e-19 $X=7.49 $Y=1.185
+ $X2=0 $Y2=0
cc_507 N_A_772_21#_c_491_n N_A_27_47#_c_1286_n 0.00203544f $X=6.515 $Y=1.26
+ $X2=0 $Y2=0
cc_508 N_A_772_21#_c_492_n N_A_27_47#_c_1286_n 0.00363484f $X=6.945 $Y=1.26
+ $X2=0 $Y2=0
cc_509 N_A_772_21#_c_494_n N_A_27_47#_c_1286_n 0.0133739f $X=7.525 $Y=1.685
+ $X2=0 $Y2=0
cc_510 N_A_772_21#_c_481_n N_A_27_47#_c_1287_n 6.49145e-19 $X=6.515 $Y=1.185
+ $X2=0 $Y2=0
cc_511 N_A_772_21#_c_483_n N_A_27_47#_c_1287_n 0.0125382f $X=6.945 $Y=1.185
+ $X2=0 $Y2=0
cc_512 N_A_772_21#_c_495_n N_A_27_47#_c_1287_n 0.0698454f $X=7.58 $Y=0.42 $X2=0
+ $Y2=0
cc_513 N_A_772_21#_c_496_n N_A_27_47#_c_1287_n 0.00666405f $X=7.58 $Y=0.42 $X2=0
+ $Y2=0
cc_514 N_A_772_21#_c_471_n N_A_27_47#_c_1304_n 7.00608e-19 $X=4.365 $Y=1.185
+ $X2=0 $Y2=0
cc_515 N_A_772_21#_c_472_n N_A_27_47#_c_1304_n 0.00698564f $X=4.72 $Y=1.26 $X2=0
+ $Y2=0
cc_516 N_A_772_21#_c_473_n N_A_27_47#_c_1304_n 7.00608e-19 $X=4.795 $Y=1.185
+ $X2=0 $Y2=0
cc_517 N_A_772_21#_c_486_n N_A_27_47#_c_1304_n 4.11567e-19 $X=4.365 $Y=1.26
+ $X2=0 $Y2=0
cc_518 N_A_772_21#_c_487_n N_A_27_47#_c_1304_n 4.11567e-19 $X=4.795 $Y=1.26
+ $X2=0 $Y2=0
cc_519 N_A_772_21#_c_475_n N_A_27_47#_c_1305_n 7.00608e-19 $X=5.225 $Y=1.185
+ $X2=0 $Y2=0
cc_520 N_A_772_21#_c_476_n N_A_27_47#_c_1305_n 0.00698564f $X=5.58 $Y=1.26 $X2=0
+ $Y2=0
cc_521 N_A_772_21#_c_477_n N_A_27_47#_c_1305_n 7.00608e-19 $X=5.655 $Y=1.185
+ $X2=0 $Y2=0
cc_522 N_A_772_21#_c_488_n N_A_27_47#_c_1305_n 4.11567e-19 $X=5.225 $Y=1.26
+ $X2=0 $Y2=0
cc_523 N_A_772_21#_c_489_n N_A_27_47#_c_1305_n 4.11567e-19 $X=5.655 $Y=1.26
+ $X2=0 $Y2=0
cc_524 N_A_772_21#_c_479_n N_A_27_47#_c_1306_n 7.00608e-19 $X=6.085 $Y=1.185
+ $X2=0 $Y2=0
cc_525 N_A_772_21#_c_480_n N_A_27_47#_c_1306_n 0.00698564f $X=6.44 $Y=1.26 $X2=0
+ $Y2=0
cc_526 N_A_772_21#_c_481_n N_A_27_47#_c_1306_n 7.00608e-19 $X=6.515 $Y=1.185
+ $X2=0 $Y2=0
cc_527 N_A_772_21#_c_490_n N_A_27_47#_c_1306_n 4.11567e-19 $X=6.085 $Y=1.26
+ $X2=0 $Y2=0
cc_528 N_A_772_21#_c_491_n N_A_27_47#_c_1306_n 4.11567e-19 $X=6.515 $Y=1.26
+ $X2=0 $Y2=0
cc_529 N_A_772_21#_c_468_n N_VGND_c_1433_n 0.0127113f $X=3.935 $Y=1.185 $X2=0
+ $Y2=0
cc_530 N_A_772_21#_c_469_n N_VGND_c_1433_n 7.02169e-19 $X=4.29 $Y=1.26 $X2=0
+ $Y2=0
cc_531 N_A_772_21#_c_471_n N_VGND_c_1433_n 0.00295454f $X=4.365 $Y=1.185 $X2=0
+ $Y2=0
cc_532 N_A_772_21#_c_473_n N_VGND_c_1434_n 0.00284434f $X=4.795 $Y=1.185 $X2=0
+ $Y2=0
cc_533 N_A_772_21#_c_474_n N_VGND_c_1434_n 7.02169e-19 $X=5.15 $Y=1.26 $X2=0
+ $Y2=0
cc_534 N_A_772_21#_c_475_n N_VGND_c_1434_n 0.00284434f $X=5.225 $Y=1.185 $X2=0
+ $Y2=0
cc_535 N_A_772_21#_c_477_n N_VGND_c_1435_n 0.00284434f $X=5.655 $Y=1.185 $X2=0
+ $Y2=0
cc_536 N_A_772_21#_c_478_n N_VGND_c_1435_n 7.02169e-19 $X=6.01 $Y=1.26 $X2=0
+ $Y2=0
cc_537 N_A_772_21#_c_479_n N_VGND_c_1435_n 0.00284434f $X=6.085 $Y=1.185 $X2=0
+ $Y2=0
cc_538 N_A_772_21#_c_481_n N_VGND_c_1436_n 0.00284434f $X=6.515 $Y=1.185 $X2=0
+ $Y2=0
cc_539 N_A_772_21#_c_482_n N_VGND_c_1436_n 7.02169e-19 $X=6.87 $Y=1.26 $X2=0
+ $Y2=0
cc_540 N_A_772_21#_c_483_n N_VGND_c_1436_n 0.00284434f $X=6.945 $Y=1.185 $X2=0
+ $Y2=0
cc_541 N_A_772_21#_c_471_n N_VGND_c_1440_n 0.0054895f $X=4.365 $Y=1.185 $X2=0
+ $Y2=0
cc_542 N_A_772_21#_c_473_n N_VGND_c_1440_n 0.0054895f $X=4.795 $Y=1.185 $X2=0
+ $Y2=0
cc_543 N_A_772_21#_c_475_n N_VGND_c_1442_n 0.00550269f $X=5.225 $Y=1.185 $X2=0
+ $Y2=0
cc_544 N_A_772_21#_c_477_n N_VGND_c_1442_n 0.00550269f $X=5.655 $Y=1.185 $X2=0
+ $Y2=0
cc_545 N_A_772_21#_c_479_n N_VGND_c_1444_n 0.0054895f $X=6.085 $Y=1.185 $X2=0
+ $Y2=0
cc_546 N_A_772_21#_c_481_n N_VGND_c_1444_n 0.0054895f $X=6.515 $Y=1.185 $X2=0
+ $Y2=0
cc_547 N_A_772_21#_c_468_n N_VGND_c_1446_n 0.00486043f $X=3.935 $Y=1.185 $X2=0
+ $Y2=0
cc_548 N_A_772_21#_c_483_n N_VGND_c_1447_n 0.0054895f $X=6.945 $Y=1.185 $X2=0
+ $Y2=0
cc_549 N_A_772_21#_c_495_n N_VGND_c_1447_n 0.0499714f $X=7.58 $Y=0.42 $X2=0
+ $Y2=0
cc_550 N_A_772_21#_c_496_n N_VGND_c_1447_n 0.00213688f $X=7.58 $Y=0.42 $X2=0
+ $Y2=0
cc_551 N_A_772_21#_M1020_s N_VGND_c_1451_n 0.00231914f $X=7.855 $Y=0.235 $X2=0
+ $Y2=0
cc_552 N_A_772_21#_c_468_n N_VGND_c_1451_n 0.0082726f $X=3.935 $Y=1.185 $X2=0
+ $Y2=0
cc_553 N_A_772_21#_c_471_n N_VGND_c_1451_n 0.00979301f $X=4.365 $Y=1.185 $X2=0
+ $Y2=0
cc_554 N_A_772_21#_c_473_n N_VGND_c_1451_n 0.00979301f $X=4.795 $Y=1.185 $X2=0
+ $Y2=0
cc_555 N_A_772_21#_c_475_n N_VGND_c_1451_n 0.00979494f $X=5.225 $Y=1.185 $X2=0
+ $Y2=0
cc_556 N_A_772_21#_c_477_n N_VGND_c_1451_n 0.00979494f $X=5.655 $Y=1.185 $X2=0
+ $Y2=0
cc_557 N_A_772_21#_c_479_n N_VGND_c_1451_n 0.00979301f $X=6.085 $Y=1.185 $X2=0
+ $Y2=0
cc_558 N_A_772_21#_c_481_n N_VGND_c_1451_n 0.00979301f $X=6.515 $Y=1.185 $X2=0
+ $Y2=0
cc_559 N_A_772_21#_c_483_n N_VGND_c_1451_n 0.0110927f $X=6.945 $Y=1.185 $X2=0
+ $Y2=0
cc_560 N_A_772_21#_c_495_n N_VGND_c_1451_n 0.028703f $X=7.58 $Y=0.42 $X2=0 $Y2=0
cc_561 N_TE_B_c_663_n N_A_c_841_n 0.032309f $X=8.077 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_562 N_TE_B_c_689_n N_A_M1019_g 0.032309f $X=8.077 $Y=1.725 $X2=0 $Y2=0
cc_563 N_TE_B_c_661_n N_A_c_846_n 0.032309f $X=8.03 $Y=1.35 $X2=0 $Y2=0
cc_564 N_TE_B_c_664_n N_A_27_367#_c_883_n 0.012335f $X=3.935 $Y=1.725 $X2=0
+ $Y2=0
cc_565 N_TE_B_c_645_n N_A_27_367#_c_883_n 0.00210149f $X=4.29 $Y=1.65 $X2=0
+ $Y2=0
cc_566 N_TE_B_c_667_n N_A_27_367#_c_883_n 0.0110181f $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_567 N_TE_B_c_664_n N_A_27_367#_c_920_n 8.34666e-19 $X=3.935 $Y=1.725 $X2=0
+ $Y2=0
cc_568 N_TE_B_c_667_n N_A_27_367#_c_920_n 0.0146703f $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_569 N_TE_B_c_669_n N_A_27_367#_c_920_n 0.0144592f $X=4.795 $Y=1.725 $X2=0
+ $Y2=0
cc_570 N_TE_B_c_671_n N_A_27_367#_c_920_n 7.09394e-19 $X=5.225 $Y=1.725 $X2=0
+ $Y2=0
cc_571 N_TE_B_c_669_n N_A_27_367#_c_884_n 0.0110646f $X=4.795 $Y=1.725 $X2=0
+ $Y2=0
cc_572 N_TE_B_c_648_n N_A_27_367#_c_884_n 0.00210149f $X=5.15 $Y=1.65 $X2=0
+ $Y2=0
cc_573 N_TE_B_c_671_n N_A_27_367#_c_884_n 0.0110646f $X=5.225 $Y=1.725 $X2=0
+ $Y2=0
cc_574 N_TE_B_c_669_n N_A_27_367#_c_927_n 7.09394e-19 $X=4.795 $Y=1.725 $X2=0
+ $Y2=0
cc_575 N_TE_B_c_671_n N_A_27_367#_c_927_n 0.0144592f $X=5.225 $Y=1.725 $X2=0
+ $Y2=0
cc_576 N_TE_B_c_673_n N_A_27_367#_c_927_n 0.0144592f $X=5.655 $Y=1.725 $X2=0
+ $Y2=0
cc_577 N_TE_B_c_675_n N_A_27_367#_c_927_n 7.09394e-19 $X=6.085 $Y=1.725 $X2=0
+ $Y2=0
cc_578 N_TE_B_c_673_n N_A_27_367#_c_885_n 0.0110181f $X=5.655 $Y=1.725 $X2=0
+ $Y2=0
cc_579 N_TE_B_c_650_n N_A_27_367#_c_885_n 0.00210149f $X=6.01 $Y=1.65 $X2=0
+ $Y2=0
cc_580 N_TE_B_c_675_n N_A_27_367#_c_885_n 0.0110646f $X=6.085 $Y=1.725 $X2=0
+ $Y2=0
cc_581 N_TE_B_c_675_n N_A_27_367#_c_886_n 9.02626e-19 $X=6.085 $Y=1.725 $X2=0
+ $Y2=0
cc_582 N_TE_B_c_651_n N_A_27_367#_c_886_n 0.00220396f $X=6.44 $Y=1.65 $X2=0
+ $Y2=0
cc_583 N_TE_B_c_673_n N_A_27_367#_c_936_n 4.98588e-19 $X=5.655 $Y=1.725 $X2=0
+ $Y2=0
cc_584 N_TE_B_c_675_n N_A_27_367#_c_936_n 0.00579476f $X=6.085 $Y=1.725 $X2=0
+ $Y2=0
cc_585 N_TE_B_c_675_n N_A_27_367#_c_938_n 0.00645347f $X=6.085 $Y=1.725 $X2=0
+ $Y2=0
cc_586 N_TE_B_c_677_n N_A_27_367#_c_910_n 0.0130894f $X=6.515 $Y=1.725 $X2=0
+ $Y2=0
cc_587 N_TE_B_c_679_n N_A_27_367#_c_910_n 0.00853569f $X=6.945 $Y=1.725 $X2=0
+ $Y2=0
cc_588 N_TE_B_c_667_n N_A_27_367#_c_887_n 9.57158e-19 $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_589 N_TE_B_c_647_n N_A_27_367#_c_887_n 0.00220396f $X=4.72 $Y=1.65 $X2=0
+ $Y2=0
cc_590 N_TE_B_c_669_n N_A_27_367#_c_887_n 9.57158e-19 $X=4.795 $Y=1.725 $X2=0
+ $Y2=0
cc_591 N_TE_B_c_671_n N_A_27_367#_c_888_n 9.57158e-19 $X=5.225 $Y=1.725 $X2=0
+ $Y2=0
cc_592 N_TE_B_c_649_n N_A_27_367#_c_888_n 0.00220396f $X=5.58 $Y=1.65 $X2=0
+ $Y2=0
cc_593 N_TE_B_c_673_n N_A_27_367#_c_888_n 9.57158e-19 $X=5.655 $Y=1.725 $X2=0
+ $Y2=0
cc_594 N_TE_B_c_675_n N_A_27_367#_c_947_n 0.0017646f $X=6.085 $Y=1.725 $X2=0
+ $Y2=0
cc_595 N_TE_B_c_677_n N_A_27_367#_c_889_n 6.30913e-19 $X=6.515 $Y=1.725 $X2=0
+ $Y2=0
cc_596 N_TE_B_c_679_n N_A_27_367#_c_889_n 0.00789881f $X=6.945 $Y=1.725 $X2=0
+ $Y2=0
cc_597 N_TE_B_c_664_n N_VPWR_c_1148_n 0.0168132f $X=3.935 $Y=1.725 $X2=0 $Y2=0
cc_598 N_TE_B_c_667_n N_VPWR_c_1148_n 0.00383836f $X=4.365 $Y=1.725 $X2=0 $Y2=0
cc_599 N_TE_B_c_669_n N_VPWR_c_1149_n 0.00372815f $X=4.795 $Y=1.725 $X2=0 $Y2=0
cc_600 N_TE_B_c_671_n N_VPWR_c_1149_n 0.00372815f $X=5.225 $Y=1.725 $X2=0 $Y2=0
cc_601 N_TE_B_c_673_n N_VPWR_c_1150_n 0.00372815f $X=5.655 $Y=1.725 $X2=0 $Y2=0
cc_602 N_TE_B_c_675_n N_VPWR_c_1150_n 0.00242144f $X=6.085 $Y=1.725 $X2=0 $Y2=0
cc_603 N_TE_B_c_675_n N_VPWR_c_1151_n 5.90687e-19 $X=6.085 $Y=1.725 $X2=0 $Y2=0
cc_604 N_TE_B_c_677_n N_VPWR_c_1151_n 0.00805364f $X=6.515 $Y=1.725 $X2=0 $Y2=0
cc_605 N_TE_B_c_679_n N_VPWR_c_1151_n 0.00287037f $X=6.945 $Y=1.725 $X2=0 $Y2=0
cc_606 N_TE_B_c_689_n N_VPWR_c_1152_n 0.0235043f $X=8.077 $Y=1.725 $X2=0 $Y2=0
cc_607 N_TE_B_c_667_n N_VPWR_c_1155_n 0.0054895f $X=4.365 $Y=1.725 $X2=0 $Y2=0
cc_608 N_TE_B_c_669_n N_VPWR_c_1155_n 0.0054895f $X=4.795 $Y=1.725 $X2=0 $Y2=0
cc_609 N_TE_B_c_671_n N_VPWR_c_1157_n 0.0054895f $X=5.225 $Y=1.725 $X2=0 $Y2=0
cc_610 N_TE_B_c_673_n N_VPWR_c_1157_n 0.0054895f $X=5.655 $Y=1.725 $X2=0 $Y2=0
cc_611 N_TE_B_c_675_n N_VPWR_c_1159_n 0.0054895f $X=6.085 $Y=1.725 $X2=0 $Y2=0
cc_612 N_TE_B_c_677_n N_VPWR_c_1159_n 0.00486043f $X=6.515 $Y=1.725 $X2=0 $Y2=0
cc_613 N_TE_B_c_664_n N_VPWR_c_1161_n 0.00486043f $X=3.935 $Y=1.725 $X2=0 $Y2=0
cc_614 N_TE_B_c_679_n N_VPWR_c_1162_n 0.0054895f $X=6.945 $Y=1.725 $X2=0 $Y2=0
cc_615 N_TE_B_c_689_n N_VPWR_c_1162_n 0.00486043f $X=8.077 $Y=1.725 $X2=0 $Y2=0
cc_616 N_TE_B_c_664_n N_VPWR_c_1147_n 0.0082726f $X=3.935 $Y=1.725 $X2=0 $Y2=0
cc_617 N_TE_B_c_667_n N_VPWR_c_1147_n 0.00979301f $X=4.365 $Y=1.725 $X2=0 $Y2=0
cc_618 N_TE_B_c_669_n N_VPWR_c_1147_n 0.00979301f $X=4.795 $Y=1.725 $X2=0 $Y2=0
cc_619 N_TE_B_c_671_n N_VPWR_c_1147_n 0.00979301f $X=5.225 $Y=1.725 $X2=0 $Y2=0
cc_620 N_TE_B_c_673_n N_VPWR_c_1147_n 0.00979301f $X=5.655 $Y=1.725 $X2=0 $Y2=0
cc_621 N_TE_B_c_675_n N_VPWR_c_1147_n 0.00979301f $X=6.085 $Y=1.725 $X2=0 $Y2=0
cc_622 N_TE_B_c_677_n N_VPWR_c_1147_n 0.00444753f $X=6.515 $Y=1.725 $X2=0 $Y2=0
cc_623 N_TE_B_c_679_n N_VPWR_c_1147_n 0.00727721f $X=6.945 $Y=1.725 $X2=0 $Y2=0
cc_624 N_TE_B_c_689_n N_VPWR_c_1147_n 0.00602946f $X=8.077 $Y=1.725 $X2=0 $Y2=0
cc_625 N_TE_B_c_646_n N_A_27_47#_c_1282_n 5.52071e-19 $X=4.01 $Y=1.65 $X2=0
+ $Y2=0
cc_626 N_TE_B_c_655_n N_A_27_47#_c_1284_n 5.26766e-19 $X=4.795 $Y=1.65 $X2=0
+ $Y2=0
cc_627 N_TE_B_c_657_n N_A_27_47#_c_1285_n 5.26766e-19 $X=5.655 $Y=1.65 $X2=0
+ $Y2=0
cc_628 N_TE_B_c_652_n N_A_27_47#_c_1286_n 0.00185993f $X=6.87 $Y=1.65 $X2=0
+ $Y2=0
cc_629 N_TE_B_c_659_n N_A_27_47#_c_1286_n 2.60763e-19 $X=6.515 $Y=1.65 $X2=0
+ $Y2=0
cc_630 N_TE_B_c_660_n N_A_27_47#_c_1286_n 0.00160884f $X=6.945 $Y=1.65 $X2=0
+ $Y2=0
cc_631 N_TE_B_c_654_n N_A_27_47#_c_1304_n 3.23907e-19 $X=4.365 $Y=1.65 $X2=0
+ $Y2=0
cc_632 N_TE_B_c_656_n N_A_27_47#_c_1305_n 3.23907e-19 $X=5.225 $Y=1.65 $X2=0
+ $Y2=0
cc_633 N_TE_B_c_658_n N_A_27_47#_c_1306_n 3.23907e-19 $X=6.085 $Y=1.65 $X2=0
+ $Y2=0
cc_634 N_TE_B_c_663_n N_VGND_c_1437_n 0.00290159f $X=8.077 $Y=1.185 $X2=0 $Y2=0
cc_635 N_TE_B_c_663_n N_VGND_c_1447_n 0.0054895f $X=8.077 $Y=1.185 $X2=0 $Y2=0
cc_636 N_TE_B_c_663_n N_VGND_c_1451_n 0.0111812f $X=8.077 $Y=1.185 $X2=0 $Y2=0
cc_637 N_A_M1019_g N_VPWR_c_1152_n 0.00303283f $X=8.645 $Y=2.465 $X2=0 $Y2=0
cc_638 N_A_M1033_g N_VPWR_c_1154_n 0.00858314f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_639 N_A_M1019_g N_VPWR_c_1163_n 0.0054895f $X=8.645 $Y=2.465 $X2=0 $Y2=0
cc_640 N_A_M1033_g N_VPWR_c_1163_n 0.0054895f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_641 N_A_M1019_g N_VPWR_c_1147_n 0.00618371f $X=8.645 $Y=2.465 $X2=0 $Y2=0
cc_642 N_A_M1033_g N_VPWR_c_1147_n 0.0107696f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_643 N_A_c_841_n N_VGND_c_1437_n 0.00290159f $X=8.645 $Y=1.185 $X2=0 $Y2=0
cc_644 N_A_c_843_n N_VGND_c_1439_n 0.00813084f $X=9.075 $Y=1.185 $X2=0 $Y2=0
cc_645 N_A_c_841_n N_VGND_c_1448_n 0.0054895f $X=8.645 $Y=1.185 $X2=0 $Y2=0
cc_646 N_A_c_843_n N_VGND_c_1448_n 0.0054895f $X=9.075 $Y=1.185 $X2=0 $Y2=0
cc_647 N_A_c_841_n N_VGND_c_1451_n 0.00617541f $X=8.645 $Y=1.185 $X2=0 $Y2=0
cc_648 N_A_c_843_n N_VGND_c_1451_n 0.0107235f $X=9.075 $Y=1.185 $X2=0 $Y2=0
cc_649 N_A_27_367#_c_894_n N_Z_M1006_d 0.00332344f $X=0.975 $Y=2.99 $X2=0 $Y2=0
cc_650 N_A_27_367#_c_898_n N_Z_M1016_d 0.00332344f $X=1.915 $Y=2.99 $X2=0 $Y2=0
cc_651 N_A_27_367#_c_900_n N_Z_M1022_d 0.00332344f $X=2.775 $Y=2.99 $X2=0 $Y2=0
cc_652 N_A_27_367#_c_902_n N_Z_M1035_d 0.00332344f $X=3.635 $Y=2.99 $X2=0 $Y2=0
cc_653 N_A_27_367#_M1011_s N_Z_c_1019_n 0.00176461f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_654 N_A_27_367#_c_896_n N_Z_c_1019_n 0.0152916f $X=1.14 $Y=2.32 $X2=0 $Y2=0
cc_655 N_A_27_367#_M1021_s N_Z_c_1020_n 0.00176461f $X=1.86 $Y=1.835 $X2=0 $Y2=0
cc_656 N_A_27_367#_c_957_p N_Z_c_1020_n 0.0135055f $X=2 $Y=2.32 $X2=0 $Y2=0
cc_657 N_A_27_367#_M1024_s N_Z_c_1021_n 0.00176461f $X=2.72 $Y=1.835 $X2=0 $Y2=0
cc_658 N_A_27_367#_c_959_p N_Z_c_1021_n 0.0135055f $X=2.86 $Y=2.32 $X2=0 $Y2=0
cc_659 N_A_27_367#_c_881_n N_Z_c_1109_n 0.00697079f $X=0.28 $Y=1.98 $X2=0 $Y2=0
cc_660 N_A_27_367#_c_894_n N_Z_c_1109_n 0.0126348f $X=0.975 $Y=2.99 $X2=0 $Y2=0
cc_661 N_A_27_367#_c_898_n N_Z_c_1022_n 0.0159805f $X=1.915 $Y=2.99 $X2=0 $Y2=0
cc_662 N_A_27_367#_c_900_n N_Z_c_1023_n 0.0159805f $X=2.775 $Y=2.99 $X2=0 $Y2=0
cc_663 N_A_27_367#_c_902_n N_Z_c_1024_n 0.0159805f $X=3.635 $Y=2.99 $X2=0 $Y2=0
cc_664 N_A_27_367#_c_882_n N_Z_c_1024_n 0.00772305f $X=3.72 $Y=1.985 $X2=0 $Y2=0
cc_665 N_A_27_367#_c_881_n N_Z_c_1017_n 0.0148572f $X=0.28 $Y=1.98 $X2=0 $Y2=0
cc_666 N_A_27_367#_c_883_n N_VPWR_M1000_d 0.00176461f $X=4.415 $Y=1.9 $X2=-0.19
+ $Y2=1.655
cc_667 N_A_27_367#_c_884_n N_VPWR_M1013_d 0.00176461f $X=5.275 $Y=1.9 $X2=0
+ $Y2=0
cc_668 N_A_27_367#_c_885_n N_VPWR_M1018_d 0.00176461f $X=6.135 $Y=1.9 $X2=0
+ $Y2=0
cc_669 N_A_27_367#_c_910_n N_VPWR_M1030_d 0.00340956f $X=6.995 $Y=2.45 $X2=0
+ $Y2=0
cc_670 N_A_27_367#_c_883_n N_VPWR_c_1148_n 0.0152916f $X=4.415 $Y=1.9 $X2=0
+ $Y2=0
cc_671 N_A_27_367#_c_884_n N_VPWR_c_1149_n 0.0135055f $X=5.275 $Y=1.9 $X2=0
+ $Y2=0
cc_672 N_A_27_367#_c_885_n N_VPWR_c_1150_n 0.0135055f $X=6.135 $Y=1.9 $X2=0
+ $Y2=0
cc_673 N_A_27_367#_c_910_n N_VPWR_c_1151_n 0.0149901f $X=6.995 $Y=2.45 $X2=0
+ $Y2=0
cc_674 N_A_27_367#_c_920_n N_VPWR_c_1155_n 0.0189236f $X=4.58 $Y=2.91 $X2=0
+ $Y2=0
cc_675 N_A_27_367#_c_927_n N_VPWR_c_1157_n 0.0189236f $X=5.44 $Y=2.91 $X2=0
+ $Y2=0
cc_676 N_A_27_367#_c_938_n N_VPWR_c_1159_n 0.0153332f $X=6.3 $Y=2.91 $X2=0 $Y2=0
cc_677 N_A_27_367#_c_880_n N_VPWR_c_1161_n 0.021159f $X=0.28 $Y=2.905 $X2=0
+ $Y2=0
cc_678 N_A_27_367#_c_894_n N_VPWR_c_1161_n 0.0298674f $X=0.975 $Y=2.99 $X2=0
+ $Y2=0
cc_679 N_A_27_367#_c_898_n N_VPWR_c_1161_n 0.0368226f $X=1.915 $Y=2.99 $X2=0
+ $Y2=0
cc_680 N_A_27_367#_c_900_n N_VPWR_c_1161_n 0.0368226f $X=2.775 $Y=2.99 $X2=0
+ $Y2=0
cc_681 N_A_27_367#_c_902_n N_VPWR_c_1161_n 0.0368226f $X=3.635 $Y=2.99 $X2=0
+ $Y2=0
cc_682 N_A_27_367#_c_983_p N_VPWR_c_1161_n 0.0118138f $X=3.72 $Y=2.905 $X2=0
+ $Y2=0
cc_683 N_A_27_367#_c_912_n N_VPWR_c_1161_n 0.0154369f $X=1.1 $Y=2.99 $X2=0 $Y2=0
cc_684 N_A_27_367#_c_985_p N_VPWR_c_1161_n 0.0118138f $X=2 $Y=2.99 $X2=0 $Y2=0
cc_685 N_A_27_367#_c_986_p N_VPWR_c_1161_n 0.0118138f $X=2.86 $Y=2.99 $X2=0
+ $Y2=0
cc_686 N_A_27_367#_c_889_n N_VPWR_c_1162_n 0.0210796f $X=7.16 $Y=2.53 $X2=0
+ $Y2=0
cc_687 N_A_27_367#_M1006_s N_VPWR_c_1147_n 0.00231914f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_688 N_A_27_367#_M1011_s N_VPWR_c_1147_n 0.00223562f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_689 N_A_27_367#_M1021_s N_VPWR_c_1147_n 0.00223566f $X=1.86 $Y=1.835 $X2=0
+ $Y2=0
cc_690 N_A_27_367#_M1024_s N_VPWR_c_1147_n 0.00223566f $X=2.72 $Y=1.835 $X2=0
+ $Y2=0
cc_691 N_A_27_367#_M1036_s N_VPWR_c_1147_n 0.00411415f $X=3.58 $Y=1.835 $X2=0
+ $Y2=0
cc_692 N_A_27_367#_M1002_s N_VPWR_c_1147_n 0.00223559f $X=4.44 $Y=1.835 $X2=0
+ $Y2=0
cc_693 N_A_27_367#_M1014_s N_VPWR_c_1147_n 0.00223559f $X=5.3 $Y=1.835 $X2=0
+ $Y2=0
cc_694 N_A_27_367#_M1027_s N_VPWR_c_1147_n 0.00254932f $X=6.16 $Y=1.835 $X2=0
+ $Y2=0
cc_695 N_A_27_367#_M1034_s N_VPWR_c_1147_n 0.00231914f $X=7.02 $Y=1.835 $X2=0
+ $Y2=0
cc_696 N_A_27_367#_c_880_n N_VPWR_c_1147_n 0.0126421f $X=0.28 $Y=2.905 $X2=0
+ $Y2=0
cc_697 N_A_27_367#_c_894_n N_VPWR_c_1147_n 0.0187823f $X=0.975 $Y=2.99 $X2=0
+ $Y2=0
cc_698 N_A_27_367#_c_898_n N_VPWR_c_1147_n 0.024428f $X=1.915 $Y=2.99 $X2=0
+ $Y2=0
cc_699 N_A_27_367#_c_900_n N_VPWR_c_1147_n 0.024428f $X=2.775 $Y=2.99 $X2=0
+ $Y2=0
cc_700 N_A_27_367#_c_902_n N_VPWR_c_1147_n 0.024428f $X=3.635 $Y=2.99 $X2=0
+ $Y2=0
cc_701 N_A_27_367#_c_983_p N_VPWR_c_1147_n 0.00658808f $X=3.72 $Y=2.905 $X2=0
+ $Y2=0
cc_702 N_A_27_367#_c_920_n N_VPWR_c_1147_n 0.0123859f $X=4.58 $Y=2.91 $X2=0
+ $Y2=0
cc_703 N_A_27_367#_c_927_n N_VPWR_c_1147_n 0.0123859f $X=5.44 $Y=2.91 $X2=0
+ $Y2=0
cc_704 N_A_27_367#_c_938_n N_VPWR_c_1147_n 0.00945339f $X=6.3 $Y=2.91 $X2=0
+ $Y2=0
cc_705 N_A_27_367#_c_910_n N_VPWR_c_1147_n 0.0118711f $X=6.995 $Y=2.45 $X2=0
+ $Y2=0
cc_706 N_A_27_367#_c_912_n N_VPWR_c_1147_n 0.00952129f $X=1.1 $Y=2.99 $X2=0
+ $Y2=0
cc_707 N_A_27_367#_c_985_p N_VPWR_c_1147_n 0.00658808f $X=2 $Y=2.99 $X2=0 $Y2=0
cc_708 N_A_27_367#_c_986_p N_VPWR_c_1147_n 0.00658808f $X=2.86 $Y=2.99 $X2=0
+ $Y2=0
cc_709 N_A_27_367#_c_889_n N_VPWR_c_1147_n 0.0125834f $X=7.16 $Y=2.53 $X2=0
+ $Y2=0
cc_710 N_Z_M1006_d N_VPWR_c_1147_n 0.00225186f $X=0.57 $Y=1.835 $X2=0 $Y2=0
cc_711 N_Z_M1016_d N_VPWR_c_1147_n 0.00225186f $X=1.43 $Y=1.835 $X2=0 $Y2=0
cc_712 N_Z_M1022_d N_VPWR_c_1147_n 0.00225186f $X=2.29 $Y=1.835 $X2=0 $Y2=0
cc_713 N_Z_M1035_d N_VPWR_c_1147_n 0.00225186f $X=3.15 $Y=1.835 $X2=0 $Y2=0
cc_714 N_Z_c_1012_n N_A_27_47#_M1005_d 0.00176461f $X=1.405 $Y=1.06 $X2=0 $Y2=0
cc_715 N_Z_c_1013_n N_A_27_47#_M1010_d 0.00176461f $X=2.265 $Y=1.06 $X2=0 $Y2=0
cc_716 N_Z_c_1014_n N_A_27_47#_M1025_d 0.00176461f $X=3.125 $Y=1.06 $X2=0 $Y2=0
cc_717 N_Z_M1003_s N_A_27_47#_c_1289_n 0.00332344f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_718 N_Z_c_1025_n N_A_27_47#_c_1289_n 0.0160265f $X=0.71 $Y=0.805 $X2=0 $Y2=0
cc_719 N_Z_c_1012_n N_A_27_47#_c_1289_n 0.00320534f $X=1.405 $Y=1.06 $X2=0 $Y2=0
cc_720 N_Z_c_1012_n N_A_27_47#_c_1377_n 0.0132747f $X=1.405 $Y=1.06 $X2=0 $Y2=0
cc_721 N_Z_M1009_s N_A_27_47#_c_1291_n 0.00332344f $X=1.43 $Y=0.235 $X2=0 $Y2=0
cc_722 N_Z_c_1012_n N_A_27_47#_c_1291_n 0.00320534f $X=1.405 $Y=1.06 $X2=0 $Y2=0
cc_723 N_Z_c_1044_n N_A_27_47#_c_1291_n 0.0157943f $X=1.57 $Y=0.805 $X2=0 $Y2=0
cc_724 N_Z_c_1013_n N_A_27_47#_c_1291_n 0.00320534f $X=2.265 $Y=1.06 $X2=0 $Y2=0
cc_725 N_Z_c_1013_n N_A_27_47#_c_1382_n 0.0132747f $X=2.265 $Y=1.06 $X2=0 $Y2=0
cc_726 N_Z_M1017_s N_A_27_47#_c_1293_n 0.00332344f $X=2.29 $Y=0.235 $X2=0 $Y2=0
cc_727 N_Z_c_1013_n N_A_27_47#_c_1293_n 0.00320534f $X=2.265 $Y=1.06 $X2=0 $Y2=0
cc_728 N_Z_c_1056_n N_A_27_47#_c_1293_n 0.0157943f $X=2.43 $Y=0.805 $X2=0 $Y2=0
cc_729 N_Z_c_1014_n N_A_27_47#_c_1293_n 0.00320534f $X=3.125 $Y=1.06 $X2=0 $Y2=0
cc_730 N_Z_c_1014_n N_A_27_47#_c_1387_n 0.0132747f $X=3.125 $Y=1.06 $X2=0 $Y2=0
cc_731 N_Z_M1028_s N_A_27_47#_c_1295_n 0.00332344f $X=3.15 $Y=0.235 $X2=0 $Y2=0
cc_732 N_Z_c_1014_n N_A_27_47#_c_1295_n 0.00320534f $X=3.125 $Y=1.06 $X2=0 $Y2=0
cc_733 N_Z_c_1069_n N_A_27_47#_c_1295_n 0.0157943f $X=3.29 $Y=0.805 $X2=0 $Y2=0
cc_734 N_Z_c_1014_n N_A_27_47#_c_1281_n 0.00854023f $X=3.125 $Y=1.06 $X2=0 $Y2=0
cc_735 N_Z_c_1014_n N_A_27_47#_c_1283_n 8.53482e-19 $X=3.125 $Y=1.06 $X2=0 $Y2=0
cc_736 N_Z_c_1017_n N_A_27_47#_c_1288_n 0.0201602f $X=0.545 $Y=1.295 $X2=0 $Y2=0
cc_737 N_Z_M1003_s N_VGND_c_1451_n 0.00225186f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_738 N_Z_M1009_s N_VGND_c_1451_n 0.00225186f $X=1.43 $Y=0.235 $X2=0 $Y2=0
cc_739 N_Z_M1017_s N_VGND_c_1451_n 0.00225186f $X=2.29 $Y=0.235 $X2=0 $Y2=0
cc_740 N_Z_M1028_s N_VGND_c_1451_n 0.00225186f $X=3.15 $Y=0.235 $X2=0 $Y2=0
cc_741 N_A_27_47#_c_1282_n N_VGND_c_1433_n 0.0177053f $X=4.415 $Y=1.22 $X2=0
+ $Y2=0
cc_742 N_A_27_47#_c_1284_n N_VGND_c_1434_n 0.013802f $X=5.275 $Y=1.22 $X2=0
+ $Y2=0
cc_743 N_A_27_47#_c_1285_n N_VGND_c_1435_n 0.013802f $X=6.135 $Y=1.22 $X2=0
+ $Y2=0
cc_744 N_A_27_47#_c_1286_n N_VGND_c_1436_n 0.013802f $X=6.995 $Y=1.22 $X2=0
+ $Y2=0
cc_745 N_A_27_47#_c_1313_n N_VGND_c_1440_n 0.0189236f $X=4.58 $Y=0.42 $X2=0
+ $Y2=0
cc_746 N_A_27_47#_c_1322_n N_VGND_c_1442_n 0.015091f $X=5.44 $Y=0.38 $X2=0 $Y2=0
cc_747 N_A_27_47#_c_1331_n N_VGND_c_1444_n 0.0189236f $X=6.3 $Y=0.42 $X2=0 $Y2=0
cc_748 N_A_27_47#_c_1289_n N_VGND_c_1446_n 0.0368488f $X=1.055 $Y=0.34 $X2=0
+ $Y2=0
cc_749 N_A_27_47#_c_1291_n N_VGND_c_1446_n 0.0368751f $X=1.915 $Y=0.34 $X2=0
+ $Y2=0
cc_750 N_A_27_47#_c_1293_n N_VGND_c_1446_n 0.0368751f $X=2.775 $Y=0.34 $X2=0
+ $Y2=0
cc_751 N_A_27_47#_c_1295_n N_VGND_c_1446_n 0.0368488f $X=3.635 $Y=0.34 $X2=0
+ $Y2=0
cc_752 N_A_27_47#_c_1405_p N_VGND_c_1446_n 0.0118138f $X=3.72 $Y=0.425 $X2=0
+ $Y2=0
cc_753 N_A_27_47#_c_1288_n N_VGND_c_1446_n 0.017536f $X=0.28 $Y=0.42 $X2=0 $Y2=0
cc_754 N_A_27_47#_c_1407_p N_VGND_c_1446_n 0.0116347f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_755 N_A_27_47#_c_1408_p N_VGND_c_1446_n 0.0116347f $X=2 $Y=0.34 $X2=0 $Y2=0
cc_756 N_A_27_47#_c_1409_p N_VGND_c_1446_n 0.0116347f $X=2.86 $Y=0.34 $X2=0
+ $Y2=0
cc_757 N_A_27_47#_c_1287_n N_VGND_c_1447_n 0.0153681f $X=7.16 $Y=0.42 $X2=0
+ $Y2=0
cc_758 N_A_27_47#_M1003_d N_VGND_c_1451_n 0.00231918f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_759 N_A_27_47#_M1005_d N_VGND_c_1451_n 0.00225174f $X=1 $Y=0.235 $X2=0 $Y2=0
cc_760 N_A_27_47#_M1010_d N_VGND_c_1451_n 0.00225174f $X=1.86 $Y=0.235 $X2=0
+ $Y2=0
cc_761 N_A_27_47#_M1025_d N_VGND_c_1451_n 0.00225174f $X=2.72 $Y=0.235 $X2=0
+ $Y2=0
cc_762 N_A_27_47#_M1031_d N_VGND_c_1451_n 0.00411415f $X=3.58 $Y=0.235 $X2=0
+ $Y2=0
cc_763 N_A_27_47#_M1004_s N_VGND_c_1451_n 0.00223559f $X=4.44 $Y=0.235 $X2=0
+ $Y2=0
cc_764 N_A_27_47#_M1015_s N_VGND_c_1451_n 0.00225632f $X=5.3 $Y=0.235 $X2=0
+ $Y2=0
cc_765 N_A_27_47#_M1026_s N_VGND_c_1451_n 0.00223559f $X=6.16 $Y=0.235 $X2=0
+ $Y2=0
cc_766 N_A_27_47#_M1037_s N_VGND_c_1451_n 0.00444118f $X=7.02 $Y=0.235 $X2=0
+ $Y2=0
cc_767 N_A_27_47#_c_1289_n N_VGND_c_1451_n 0.0244986f $X=1.055 $Y=0.34 $X2=0
+ $Y2=0
cc_768 N_A_27_47#_c_1291_n N_VGND_c_1451_n 0.0245693f $X=1.915 $Y=0.34 $X2=0
+ $Y2=0
cc_769 N_A_27_47#_c_1293_n N_VGND_c_1451_n 0.0245693f $X=2.775 $Y=0.34 $X2=0
+ $Y2=0
cc_770 N_A_27_47#_c_1295_n N_VGND_c_1451_n 0.0244986f $X=3.635 $Y=0.34 $X2=0
+ $Y2=0
cc_771 N_A_27_47#_c_1405_p N_VGND_c_1451_n 0.00658808f $X=3.72 $Y=0.425 $X2=0
+ $Y2=0
cc_772 N_A_27_47#_c_1313_n N_VGND_c_1451_n 0.0123859f $X=4.58 $Y=0.42 $X2=0
+ $Y2=0
cc_773 N_A_27_47#_c_1322_n N_VGND_c_1451_n 0.0121307f $X=5.44 $Y=0.38 $X2=0
+ $Y2=0
cc_774 N_A_27_47#_c_1331_n N_VGND_c_1451_n 0.0123859f $X=6.3 $Y=0.42 $X2=0 $Y2=0
cc_775 N_A_27_47#_c_1287_n N_VGND_c_1451_n 0.00945867f $X=7.16 $Y=0.42 $X2=0
+ $Y2=0
cc_776 N_A_27_47#_c_1288_n N_VGND_c_1451_n 0.00970886f $X=0.28 $Y=0.42 $X2=0
+ $Y2=0
cc_777 N_A_27_47#_c_1407_p N_VGND_c_1451_n 0.00655263f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_778 N_A_27_47#_c_1408_p N_VGND_c_1451_n 0.00655263f $X=2 $Y=0.34 $X2=0 $Y2=0
cc_779 N_A_27_47#_c_1409_p N_VGND_c_1451_n 0.00655263f $X=2.86 $Y=0.34 $X2=0
+ $Y2=0
