* File: sky130_fd_sc_lp__or2_1.pxi.spice
* Created: Wed Sep  2 10:28:57 2020
* 
x_PM_SKY130_FD_SC_LP__OR2_1%B N_B_c_43_n N_B_c_44_n N_B_c_45_n N_B_M1001_g
+ N_B_c_49_n N_B_M1003_g B N_B_c_47_n PM_SKY130_FD_SC_LP__OR2_1%B
x_PM_SKY130_FD_SC_LP__OR2_1%A N_A_M1005_g N_A_M1002_g A A N_A_c_76_n N_A_c_77_n
+ PM_SKY130_FD_SC_LP__OR2_1%A
x_PM_SKY130_FD_SC_LP__OR2_1%A_76_367# N_A_76_367#_M1001_d N_A_76_367#_M1003_s
+ N_A_76_367#_M1000_g N_A_76_367#_M1004_g N_A_76_367#_c_121_n
+ N_A_76_367#_c_122_n N_A_76_367#_c_123_n N_A_76_367#_c_141_n
+ N_A_76_367#_c_116_n N_A_76_367#_c_117_n N_A_76_367#_c_118_n
+ N_A_76_367#_c_148_n N_A_76_367#_c_119_n PM_SKY130_FD_SC_LP__OR2_1%A_76_367#
x_PM_SKY130_FD_SC_LP__OR2_1%VPWR N_VPWR_M1005_d N_VPWR_c_180_n VPWR
+ N_VPWR_c_181_n N_VPWR_c_182_n N_VPWR_c_179_n N_VPWR_c_184_n
+ PM_SKY130_FD_SC_LP__OR2_1%VPWR
x_PM_SKY130_FD_SC_LP__OR2_1%X N_X_M1000_d N_X_M1004_d X X X X X X X N_X_c_199_n
+ PM_SKY130_FD_SC_LP__OR2_1%X
x_PM_SKY130_FD_SC_LP__OR2_1%VGND N_VGND_M1001_s N_VGND_M1002_d N_VGND_c_213_n
+ N_VGND_c_214_n N_VGND_c_215_n N_VGND_c_216_n N_VGND_c_217_n N_VGND_c_218_n
+ VGND N_VGND_c_219_n N_VGND_c_220_n PM_SKY130_FD_SC_LP__OR2_1%VGND
cc_1 VNB N_B_c_43_n 0.0171225f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.26
cc_2 VNB N_B_c_44_n 0.0100967f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.65
cc_3 VNB N_B_c_45_n 0.020915f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.185
cc_4 VNB B 0.0323535f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_B_c_47_n 0.047052f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.35
cc_6 VNB N_A_M1005_g 0.0104039f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.65
cc_7 VNB A 0.0103566f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.045
cc_8 VNB N_A_c_76_n 0.0309721f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.26
cc_9 VNB N_A_c_77_n 0.0192035f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.35
cc_10 VNB N_A_76_367#_M1000_g 0.0227833f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.045
cc_11 VNB N_A_76_367#_M1004_g 0.00689153f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.26
cc_12 VNB N_A_76_367#_c_116_n 0.00256721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_76_367#_c_117_n 0.00158959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_76_367#_c_118_n 0.0401612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_76_367#_c_119_n 0.00139819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_179_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB X 0.00927881f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.725
cc_18 VNB X 0.0317616f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.045
cc_19 VNB N_X_c_199_n 0.0275828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_213_n 0.0470037f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.045
cc_21 VNB N_VGND_c_214_n 0.0153786f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.26
cc_22 VNB N_VGND_c_215_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.35
cc_23 VNB N_VGND_c_216_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.65
cc_24 VNB N_VGND_c_217_n 0.0223165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_218_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_219_n 0.0184198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_220_n 0.17053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_B_c_44_n 0.00963318f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.65
cc_29 VPB N_B_c_49_n 0.0248277f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.725
cc_30 VPB N_B_c_47_n 0.0104857f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.35
cc_31 VPB N_A_M1005_g 0.0244695f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.65
cc_32 VPB N_A_76_367#_M1004_g 0.025923f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.26
cc_33 VPB N_A_76_367#_c_121_n 0.0151722f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.65
cc_34 VPB N_A_76_367#_c_122_n 0.00731948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_76_367#_c_123_n 0.00529457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A_76_367#_c_116_n 3.54537e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_180_n 0.0446188f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.865
cc_38 VPB N_VPWR_c_181_n 0.0390568f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.26
cc_39 VPB N_VPWR_c_182_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_179_n 0.0879129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_184_n 0.0125138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB X 0.0570052f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.045
cc_43 N_B_c_44_n N_A_M1005_g 0.0437529f $X=0.645 $Y=1.65 $X2=0 $Y2=0
cc_44 N_B_c_43_n A 0.0135077f $X=0.645 $Y=1.26 $X2=0 $Y2=0
cc_45 N_B_c_44_n A 0.0015216f $X=0.645 $Y=1.65 $X2=0 $Y2=0
cc_46 B A 0.0259013f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_B_c_47_n A 6.40197e-19 $X=0.27 $Y=1.35 $X2=0 $Y2=0
cc_48 N_B_c_43_n N_A_c_76_n 0.00846166f $X=0.645 $Y=1.26 $X2=0 $Y2=0
cc_49 B N_A_c_76_n 4.053e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_50 N_B_c_47_n N_A_c_76_n 7.84747e-19 $X=0.27 $Y=1.35 $X2=0 $Y2=0
cc_51 N_B_c_45_n N_A_c_77_n 0.0122943f $X=0.72 $Y=1.185 $X2=0 $Y2=0
cc_52 N_B_c_49_n N_A_76_367#_c_121_n 0.0070736f $X=0.72 $Y=1.725 $X2=0 $Y2=0
cc_53 N_B_c_44_n N_A_76_367#_c_122_n 0.00178734f $X=0.645 $Y=1.65 $X2=0 $Y2=0
cc_54 N_B_c_49_n N_A_76_367#_c_122_n 0.0080044f $X=0.72 $Y=1.725 $X2=0 $Y2=0
cc_55 N_B_c_43_n N_A_76_367#_c_123_n 9.08509e-19 $X=0.645 $Y=1.26 $X2=0 $Y2=0
cc_56 N_B_c_44_n N_A_76_367#_c_123_n 0.0087221f $X=0.645 $Y=1.65 $X2=0 $Y2=0
cc_57 N_B_c_49_n N_A_76_367#_c_123_n 0.00280843f $X=0.72 $Y=1.725 $X2=0 $Y2=0
cc_58 B N_A_76_367#_c_123_n 0.00745332f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_59 N_B_c_47_n N_A_76_367#_c_123_n 0.00554335f $X=0.27 $Y=1.35 $X2=0 $Y2=0
cc_60 N_B_c_49_n N_VPWR_c_180_n 0.00137829f $X=0.72 $Y=1.725 $X2=0 $Y2=0
cc_61 N_B_c_45_n N_VGND_c_213_n 0.00984937f $X=0.72 $Y=1.185 $X2=0 $Y2=0
cc_62 B N_VGND_c_213_n 0.00823677f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_63 N_B_c_47_n N_VGND_c_213_n 0.00761577f $X=0.27 $Y=1.35 $X2=0 $Y2=0
cc_64 N_B_c_45_n N_VGND_c_217_n 0.00332367f $X=0.72 $Y=1.185 $X2=0 $Y2=0
cc_65 N_B_c_45_n N_VGND_c_220_n 0.00387424f $X=0.72 $Y=1.185 $X2=0 $Y2=0
cc_66 N_A_c_76_n N_A_76_367#_M1000_g 8.0778e-19 $X=1.2 $Y=1.35 $X2=0 $Y2=0
cc_67 N_A_c_77_n N_A_76_367#_M1000_g 0.0110212f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_68 N_A_M1005_g N_A_76_367#_M1004_g 0.00568549f $X=1.11 $Y=2.045 $X2=0 $Y2=0
cc_69 N_A_M1005_g N_A_76_367#_c_121_n 0.00136338f $X=1.11 $Y=2.045 $X2=0 $Y2=0
cc_70 N_A_M1005_g N_A_76_367#_c_122_n 0.0151393f $X=1.11 $Y=2.045 $X2=0 $Y2=0
cc_71 A N_A_76_367#_c_122_n 0.0524773f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_c_76_n N_A_76_367#_c_122_n 0.0041933f $X=1.2 $Y=1.35 $X2=0 $Y2=0
cc_73 A N_A_76_367#_c_123_n 0.00529018f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_74 A N_A_76_367#_c_141_n 0.0171233f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_c_76_n N_A_76_367#_c_141_n 0.0030657f $X=1.2 $Y=1.35 $X2=0 $Y2=0
cc_76 N_A_c_77_n N_A_76_367#_c_141_n 0.00987855f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_77 N_A_M1005_g N_A_76_367#_c_116_n 0.00358419f $X=1.11 $Y=2.045 $X2=0 $Y2=0
cc_78 N_A_M1005_g N_A_76_367#_c_118_n 5.91761e-19 $X=1.11 $Y=2.045 $X2=0 $Y2=0
cc_79 A N_A_76_367#_c_118_n 3.43432e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A_c_76_n N_A_76_367#_c_118_n 0.0167961f $X=1.2 $Y=1.35 $X2=0 $Y2=0
cc_81 A N_A_76_367#_c_148_n 0.0180105f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_c_77_n N_A_76_367#_c_148_n 0.00498747f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_83 A N_A_76_367#_c_119_n 0.0250403f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_84 N_A_c_76_n N_A_76_367#_c_119_n 0.00141797f $X=1.2 $Y=1.35 $X2=0 $Y2=0
cc_85 N_A_c_77_n N_A_76_367#_c_119_n 0.00290307f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_86 N_A_M1005_g N_VPWR_c_180_n 0.00998093f $X=1.11 $Y=2.045 $X2=0 $Y2=0
cc_87 A N_VGND_c_213_n 0.00265613f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A_c_77_n N_VGND_c_213_n 7.88529e-19 $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_89 N_A_c_77_n N_VGND_c_214_n 0.00416468f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_90 N_A_c_77_n N_VGND_c_217_n 0.00385987f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_91 N_A_c_77_n N_VGND_c_220_n 0.0046122f $X=1.2 $Y=1.185 $X2=0 $Y2=0
cc_92 N_A_76_367#_c_122_n A_159_367# 0.0048076f $X=1.545 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_76_367#_c_122_n N_VPWR_M1005_d 0.00627998f $X=1.545 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_76_367#_M1004_g N_VPWR_c_180_n 0.0198153f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_95 N_A_76_367#_c_121_n N_VPWR_c_180_n 0.00622847f $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_96 N_A_76_367#_c_122_n N_VPWR_c_180_n 0.0507151f $X=1.545 $Y=1.77 $X2=0 $Y2=0
cc_97 N_A_76_367#_c_118_n N_VPWR_c_180_n 8.85682e-19 $X=1.77 $Y=1.375 $X2=0
+ $Y2=0
cc_98 N_A_76_367#_M1004_g N_VPWR_c_182_n 0.00486043f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_99 N_A_76_367#_M1004_g N_VPWR_c_179_n 0.00917987f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_100 N_A_76_367#_c_118_n X 0.00428211f $X=1.77 $Y=1.375 $X2=0 $Y2=0
cc_101 N_A_76_367#_M1000_g X 0.00303874f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_102 N_A_76_367#_c_122_n X 0.0132f $X=1.545 $Y=1.77 $X2=0 $Y2=0
cc_103 N_A_76_367#_c_117_n X 0.0368818f $X=1.77 $Y=1.375 $X2=0 $Y2=0
cc_104 N_A_76_367#_c_118_n X 0.0185376f $X=1.77 $Y=1.375 $X2=0 $Y2=0
cc_105 N_A_76_367#_c_119_n X 0.0076169f $X=1.71 $Y=1.21 $X2=0 $Y2=0
cc_106 N_A_76_367#_c_141_n N_VGND_M1002_d 0.0105003f $X=1.545 $Y=0.945 $X2=0
+ $Y2=0
cc_107 N_A_76_367#_c_119_n N_VGND_M1002_d 5.76007e-19 $X=1.71 $Y=1.21 $X2=0
+ $Y2=0
cc_108 N_A_76_367#_M1000_g N_VGND_c_214_n 0.0135817f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_109 N_A_76_367#_c_141_n N_VGND_c_214_n 0.0209363f $X=1.545 $Y=0.945 $X2=0
+ $Y2=0
cc_110 N_A_76_367#_c_117_n N_VGND_c_214_n 6.38284e-19 $X=1.77 $Y=1.375 $X2=0
+ $Y2=0
cc_111 N_A_76_367#_c_118_n N_VGND_c_214_n 3.07924e-19 $X=1.77 $Y=1.375 $X2=0
+ $Y2=0
cc_112 N_A_76_367#_c_148_n N_VGND_c_217_n 0.00356195f $X=0.935 $Y=0.865 $X2=0
+ $Y2=0
cc_113 N_A_76_367#_M1000_g N_VGND_c_219_n 0.00486043f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_114 N_A_76_367#_M1000_g N_VGND_c_220_n 0.00928803f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_115 N_A_76_367#_c_141_n N_VGND_c_220_n 0.0110023f $X=1.545 $Y=0.945 $X2=0
+ $Y2=0
cc_116 N_A_76_367#_c_148_n N_VGND_c_220_n 0.00717557f $X=0.935 $Y=0.865 $X2=0
+ $Y2=0
cc_117 N_VPWR_c_179_n N_X_M1004_d 0.00371702f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_118 N_VPWR_c_182_n X 0.018528f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_119 N_VPWR_c_179_n X 0.0104192f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_120 N_X_c_199_n N_VGND_c_219_n 0.0285641f $X=2 $Y=0.42 $X2=0 $Y2=0
cc_121 N_X_M1000_d N_VGND_c_220_n 0.00371702f $X=1.86 $Y=0.235 $X2=0 $Y2=0
cc_122 N_X_c_199_n N_VGND_c_220_n 0.0158621f $X=2 $Y=0.42 $X2=0 $Y2=0
