* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor2_4 A B VGND VNB VPB VPWR X
X0 VPWR A a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_110_47# B X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 X B a_110_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VPWR A a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_110_47# B X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_27_367# a_776_255# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_27_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_1199_367# B a_776_255# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_27_367# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VPWR A a_1199_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_27_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VPWR B a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_1199_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 X a_776_255# a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_27_367# a_776_255# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 X a_776_255# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_776_255# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 X a_776_255# a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VGND B a_776_255# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_1199_367# B a_776_255# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 VGND a_776_255# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_1199_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_776_255# B a_1199_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_27_367# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 VGND A a_776_255# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_776_255# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 VGND A a_776_255# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 a_776_255# B a_1199_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_776_255# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 X B a_110_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 X a_776_255# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 VGND B a_776_255# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 VPWR B a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 VPWR A a_1199_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 VGND a_776_255# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 a_776_255# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
