* File: sky130_fd_sc_lp__clkdlybuf4s50_2.spice
* Created: Wed Sep  2 09:40:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkdlybuf4s50_2.pex.spice"
.subckt sky130_fd_sc_lp__clkdlybuf4s50_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_27_52#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0876085 AS=0.1113 PD=0.804507 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_A_282_52#_M1004_d N_A_27_52#_M1004_g N_VGND_M1005_d VNB NSHORT L=0.5
+ W=1 AD=0.265 AS=0.208592 PD=2.53 PS=1.91549 NRD=0 NRS=2.988 M=1 R=2 SA=250000
+ SB=250000 A=0.5 P=3 MULT=1
MM1008 N_VGND_M1008_d N_A_282_52#_M1008_g N_A_394_52#_M1008_s VNB NSHORT L=0.5
+ W=1 AD=0.208592 AS=0.265 PD=1.91549 PS=2.53 NRD=0 NRS=0 M=1 R=2 SA=250000
+ SB=250000 A=0.5 P=3 MULT=1
MM1001 N_VGND_M1008_d N_A_394_52#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0876085 AS=0.0588 PD=0.804507 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_394_52#_M1006_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1722 AS=0.0588 PD=1.66 PS=0.7 NRD=41.424 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_A_27_52#_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.236947 AS=0.3339 PD=1.80637 PS=3.05 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1000 N_A_282_52#_M1000_d N_A_27_52#_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.5
+ W=1 AD=0.265 AS=0.188053 PD=2.53 PS=1.43363 NRD=0 NRS=1.9503 M=1 R=2 SA=250001
+ SB=250000 A=0.5 P=3 MULT=1
MM1003 N_VPWR_M1003_d N_A_282_52#_M1003_g N_A_394_52#_M1003_s VPB PHIGHVT L=0.5
+ W=1 AD=0.188053 AS=0.265 PD=1.43363 PS=2.53 NRD=0 NRS=0 M=1 R=2 SA=250000
+ SB=250001 A=0.5 P=3 MULT=1
MM1002 N_X_M1002_d N_A_394_52#_M1002_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.236947 PD=1.54 PS=1.80637 NRD=0 NRS=12.4898 M=1 R=8.4
+ SA=75000.9 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1007 N_X_M1002_d N_A_394_52#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.5166 PD=1.54 PS=3.34 NRD=0 NRS=22.655 M=1 R=8.4 SA=75001.3
+ SB=75000.3 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__clkdlybuf4s50_2.pxi.spice"
*
.ends
*
*
