* File: sky130_fd_sc_lp__iso0p_lp.pxi.spice
* Created: Fri Aug 28 10:40:56 2020
* 
x_PM_SKY130_FD_SC_LP__ISO0P_LP%SLEEP N_SLEEP_M1012_g N_SLEEP_M1005_g
+ N_SLEEP_M1006_g N_SLEEP_M1002_g SLEEP SLEEP N_SLEEP_c_62_n
+ PM_SKY130_FD_SC_LP__ISO0P_LP%SLEEP
x_PM_SKY130_FD_SC_LP__ISO0P_LP%A_27_93# N_A_27_93#_M1012_s N_A_27_93#_M1005_s
+ N_A_27_93#_M1011_g N_A_27_93#_M1007_g N_A_27_93#_M1013_g N_A_27_93#_c_96_n
+ N_A_27_93#_c_101_n N_A_27_93#_c_102_n N_A_27_93#_c_115_n N_A_27_93#_c_97_n
+ N_A_27_93#_c_104_n PM_SKY130_FD_SC_LP__ISO0P_LP%A_27_93#
x_PM_SKY130_FD_SC_LP__ISO0P_LP%A N_A_M1001_g N_A_c_156_n N_A_M1000_g N_A_M1010_g
+ N_A_c_159_n N_A_c_160_n A N_A_c_161_n N_A_c_164_n
+ PM_SKY130_FD_SC_LP__ISO0P_LP%A
x_PM_SKY130_FD_SC_LP__ISO0P_LP%A_342_489# N_A_342_489#_M1001_d
+ N_A_342_489#_M1013_d N_A_342_489#_c_204_n N_A_342_489#_M1003_g
+ N_A_342_489#_M1008_g N_A_342_489#_c_205_n N_A_342_489#_M1004_g
+ N_A_342_489#_M1009_g N_A_342_489#_c_214_n N_A_342_489#_c_215_n
+ N_A_342_489#_c_216_n N_A_342_489#_c_206_n N_A_342_489#_c_207_n
+ N_A_342_489#_c_208_n N_A_342_489#_c_209_n N_A_342_489#_c_210_n
+ N_A_342_489#_c_211_n PM_SKY130_FD_SC_LP__ISO0P_LP%A_342_489#
x_PM_SKY130_FD_SC_LP__ISO0P_LP%KAPWR N_KAPWR_M1002_d N_KAPWR_M1010_d KAPWR
+ N_KAPWR_c_279_n N_KAPWR_c_280_n N_KAPWR_c_281_n
+ PM_SKY130_FD_SC_LP__ISO0P_LP%KAPWR
x_PM_SKY130_FD_SC_LP__ISO0P_LP%X N_X_M1004_d N_X_M1009_d X X X X X N_X_c_328_n
+ PM_SKY130_FD_SC_LP__ISO0P_LP%X
x_PM_SKY130_FD_SC_LP__ISO0P_LP%VGND N_VGND_M1006_d N_VGND_M1003_s N_VGND_c_341_n
+ N_VGND_c_342_n VGND N_VGND_c_343_n N_VGND_c_344_n N_VGND_c_345_n
+ N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n PM_SKY130_FD_SC_LP__ISO0P_LP%VGND
x_PM_SKY130_FD_SC_LP__ISO0P_LP%VPWR VPWR N_VPWR_c_384_n VPWR
+ PM_SKY130_FD_SC_LP__ISO0P_LP%VPWR
cc_1 VNB N_SLEEP_M1012_g 0.0340203f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.675
cc_2 VNB N_SLEEP_M1006_g 0.035339f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.675
cc_3 VNB SLEEP 0.00855277f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_SLEEP_c_62_n 0.0357139f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.465
cc_5 VNB N_A_27_93#_M1007_g 0.0380418f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.985
cc_6 VNB N_A_27_93#_c_96_n 0.0426945f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.465
cc_7 VNB N_A_27_93#_c_97_n 0.0440266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_c_156_n 0.0109922f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.985
cc_9 VNB N_A_M1000_g 3.61206e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_M1010_g 3.74535e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_159_n 0.017557f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.655
cc_12 VNB N_A_c_160_n 0.0170764f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.655
cc_13 VNB N_A_c_161_n 0.0536741f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.465
cc_14 VNB N_A_342_489#_c_204_n 0.0188631f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.655
cc_15 VNB N_A_342_489#_c_205_n 0.020326f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.655
cc_16 VNB N_A_342_489#_c_206_n 0.00555058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_342_489#_c_207_n 0.0220155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_342_489#_c_208_n 0.0010417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_342_489#_c_209_n 0.0015967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_342_489#_c_210_n 0.00393769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_342_489#_c_211_n 0.0639765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_X_c_328_n 0.0647669f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_23 VNB N_VGND_c_341_n 0.0162715f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.3
cc_24 VNB N_VGND_c_342_n 0.0186777f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.985
cc_25 VNB N_VGND_c_343_n 0.0291685f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_26 VNB N_VGND_c_344_n 0.0295741f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.465
cc_27 VNB N_VGND_c_345_n 0.0303334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_346_n 0.271448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_347_n 0.0130796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_348_n 0.00644364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB VPWR 0.163682f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.465
cc_32 VPB N_SLEEP_M1005_g 0.0378818f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.655
cc_33 VPB N_SLEEP_M1002_g 0.0310565f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.655
cc_34 VPB N_SLEEP_c_62_n 0.0330344f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.465
cc_35 VPB N_A_27_93#_M1011_g 0.0307453f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.3
cc_36 VPB N_A_27_93#_M1013_g 0.032226f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_37 VPB N_A_27_93#_c_96_n 0.0197538f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.465
cc_38 VPB N_A_27_93#_c_101_n 0.0100893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_93#_c_102_n 0.0222599f $X=-0.19 $Y=1.655 $X2=0.732 $Y2=1.465
cc_40 VPB N_A_27_93#_c_97_n 0.0320078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_27_93#_c_104_n 0.00739525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_M1000_g 0.0472892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_M1010_g 0.0486001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_c_164_n 0.00506862f $X=-0.19 $Y=1.655 $X2=0.732 $Y2=1.295
cc_45 VPB N_A_342_489#_M1008_g 0.0190615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_342_489#_M1009_g 0.0199177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_342_489#_c_214_n 0.00687382f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.465
cc_48 VPB N_A_342_489#_c_215_n 0.00752427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_342_489#_c_216_n 0.00990386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_342_489#_c_210_n 0.00161812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_342_489#_c_211_n 0.00366798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_KAPWR_c_279_n 0.00430848f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.675
cc_53 VPB N_KAPWR_c_280_n 0.00765914f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_KAPWR_c_281_n 0.0274865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_X_c_328_n 0.0573741f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_56 VPB VPWR 0.062193f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.465
cc_57 VPB N_VPWR_c_384_n 0.114606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 N_SLEEP_M1002_g N_A_27_93#_M1011_g 0.0314794f $X=0.845 $Y=2.655 $X2=0
+ $Y2=0
cc_59 N_SLEEP_M1006_g N_A_27_93#_M1007_g 0.0116365f $X=0.845 $Y=0.675 $X2=0
+ $Y2=0
cc_60 SLEEP N_A_27_93#_M1007_g 7.25913e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_61 N_SLEEP_M1012_g N_A_27_93#_c_96_n 0.0412295f $X=0.485 $Y=0.675 $X2=0 $Y2=0
cc_62 SLEEP N_A_27_93#_c_96_n 0.0568433f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_63 N_SLEEP_M1005_g N_A_27_93#_c_101_n 0.010058f $X=0.485 $Y=2.655 $X2=0 $Y2=0
cc_64 N_SLEEP_M1005_g N_A_27_93#_c_102_n 0.0164476f $X=0.485 $Y=2.655 $X2=0
+ $Y2=0
cc_65 N_SLEEP_M1002_g N_A_27_93#_c_102_n 0.0108193f $X=0.845 $Y=2.655 $X2=0
+ $Y2=0
cc_66 SLEEP N_A_27_93#_c_102_n 0.0292015f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_SLEEP_c_62_n N_A_27_93#_c_102_n 8.69237e-19 $X=0.71 $Y=1.465 $X2=0 $Y2=0
cc_68 SLEEP N_A_27_93#_c_115_n 0.0260401f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_SLEEP_c_62_n N_A_27_93#_c_115_n 0.0032643f $X=0.71 $Y=1.465 $X2=0 $Y2=0
cc_70 SLEEP N_A_27_93#_c_97_n 0.00270332f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_SLEEP_c_62_n N_A_27_93#_c_97_n 0.0314794f $X=0.71 $Y=1.465 $X2=0 $Y2=0
cc_72 N_SLEEP_M1005_g N_KAPWR_c_279_n 0.00172352f $X=0.485 $Y=2.655 $X2=0 $Y2=0
cc_73 N_SLEEP_M1002_g N_KAPWR_c_279_n 0.00936957f $X=0.845 $Y=2.655 $X2=0 $Y2=0
cc_74 N_SLEEP_M1005_g N_KAPWR_c_281_n 0.00549309f $X=0.485 $Y=2.655 $X2=0 $Y2=0
cc_75 N_SLEEP_M1002_g N_KAPWR_c_281_n 0.00347368f $X=0.845 $Y=2.655 $X2=0 $Y2=0
cc_76 N_SLEEP_M1012_g N_VGND_c_341_n 0.00161762f $X=0.485 $Y=0.675 $X2=0 $Y2=0
cc_77 N_SLEEP_M1006_g N_VGND_c_341_n 0.0125781f $X=0.845 $Y=0.675 $X2=0 $Y2=0
cc_78 SLEEP N_VGND_c_341_n 0.00116827f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_SLEEP_M1012_g N_VGND_c_343_n 0.00510437f $X=0.485 $Y=0.675 $X2=0 $Y2=0
cc_80 N_SLEEP_M1006_g N_VGND_c_343_n 0.00424179f $X=0.845 $Y=0.675 $X2=0 $Y2=0
cc_81 N_SLEEP_M1012_g N_VGND_c_346_n 0.00515964f $X=0.485 $Y=0.675 $X2=0 $Y2=0
cc_82 N_SLEEP_M1006_g N_VGND_c_346_n 0.0043341f $X=0.845 $Y=0.675 $X2=0 $Y2=0
cc_83 N_SLEEP_M1005_g VPWR 0.00310524f $X=0.485 $Y=2.655 $X2=-0.19 $Y2=-0.245
cc_84 N_SLEEP_M1002_g VPWR 0.00310524f $X=0.845 $Y=2.655 $X2=-0.19 $Y2=-0.245
cc_85 N_SLEEP_M1005_g N_VPWR_c_384_n 0.00510437f $X=0.485 $Y=2.655 $X2=0 $Y2=0
cc_86 N_SLEEP_M1002_g N_VPWR_c_384_n 0.00488015f $X=0.845 $Y=2.655 $X2=0 $Y2=0
cc_87 N_A_27_93#_M1007_g N_A_c_156_n 0.00439272f $X=1.625 $Y=0.675 $X2=0 $Y2=0
cc_88 N_A_27_93#_c_115_n N_A_M1000_g 0.0011996f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_89 N_A_27_93#_c_97_n N_A_M1000_g 0.0393575f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_90 N_A_27_93#_M1007_g N_A_c_159_n 0.0484202f $X=1.625 $Y=0.675 $X2=0 $Y2=0
cc_91 N_A_27_93#_c_115_n N_A_c_161_n 9.47243e-19 $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_92 N_A_27_93#_c_97_n N_A_c_161_n 0.021439f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_93 N_A_27_93#_c_115_n N_A_c_164_n 0.0152671f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_94 N_A_27_93#_c_97_n N_A_c_164_n 0.0020496f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_95 N_A_27_93#_M1013_g N_A_342_489#_c_214_n 0.00689056f $X=1.635 $Y=2.655
+ $X2=0 $Y2=0
cc_96 N_A_27_93#_c_102_n N_A_342_489#_c_214_n 0.00888624f $X=1.2 $Y=2.15 $X2=0
+ $Y2=0
cc_97 N_A_27_93#_c_102_n N_A_342_489#_c_216_n 0.00534853f $X=1.2 $Y=2.15 $X2=0
+ $Y2=0
cc_98 N_A_27_93#_c_115_n N_A_342_489#_c_216_n 0.00931347f $X=1.43 $Y=1.475 $X2=0
+ $Y2=0
cc_99 N_A_27_93#_c_97_n N_A_342_489#_c_216_n 0.0014554f $X=1.43 $Y=1.475 $X2=0
+ $Y2=0
cc_100 N_A_27_93#_M1007_g N_A_342_489#_c_208_n 0.00100859f $X=1.625 $Y=0.675
+ $X2=0 $Y2=0
cc_101 N_A_27_93#_M1011_g N_KAPWR_c_279_n 0.00949732f $X=1.275 $Y=2.655 $X2=0
+ $Y2=0
cc_102 N_A_27_93#_M1013_g N_KAPWR_c_279_n 0.00174298f $X=1.635 $Y=2.655 $X2=0
+ $Y2=0
cc_103 N_A_27_93#_c_101_n N_KAPWR_c_279_n 0.00568038f $X=0.27 $Y=2.61 $X2=0
+ $Y2=0
cc_104 N_A_27_93#_c_102_n N_KAPWR_c_279_n 0.0166689f $X=1.2 $Y=2.15 $X2=0 $Y2=0
cc_105 N_A_27_93#_M1005_s N_KAPWR_c_281_n 0.00121005f $X=0.135 $Y=2.445 $X2=0
+ $Y2=0
cc_106 N_A_27_93#_M1011_g N_KAPWR_c_281_n 0.00340134f $X=1.275 $Y=2.655 $X2=0
+ $Y2=0
cc_107 N_A_27_93#_M1013_g N_KAPWR_c_281_n 0.0086286f $X=1.635 $Y=2.655 $X2=0
+ $Y2=0
cc_108 N_A_27_93#_c_101_n N_KAPWR_c_281_n 0.0269979f $X=0.27 $Y=2.61 $X2=0 $Y2=0
cc_109 N_A_27_93#_c_102_n N_KAPWR_c_281_n 0.03356f $X=1.2 $Y=2.15 $X2=0 $Y2=0
cc_110 N_A_27_93#_M1007_g N_VGND_c_341_n 0.0127454f $X=1.625 $Y=0.675 $X2=0
+ $Y2=0
cc_111 N_A_27_93#_c_96_n N_VGND_c_341_n 0.00748999f $X=0.27 $Y=0.72 $X2=0 $Y2=0
cc_112 N_A_27_93#_c_115_n N_VGND_c_341_n 0.0118129f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_113 N_A_27_93#_c_97_n N_VGND_c_341_n 0.00765182f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_114 N_A_27_93#_c_96_n N_VGND_c_343_n 0.00734893f $X=0.27 $Y=0.72 $X2=0 $Y2=0
cc_115 N_A_27_93#_M1007_g N_VGND_c_344_n 0.00424179f $X=1.625 $Y=0.675 $X2=0
+ $Y2=0
cc_116 N_A_27_93#_M1007_g N_VGND_c_346_n 0.0043341f $X=1.625 $Y=0.675 $X2=0
+ $Y2=0
cc_117 N_A_27_93#_c_96_n N_VGND_c_346_n 0.00765198f $X=0.27 $Y=0.72 $X2=0 $Y2=0
cc_118 N_A_27_93#_M1011_g VPWR 0.00310524f $X=1.275 $Y=2.655 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_27_93#_M1013_g VPWR 0.00310524f $X=1.635 $Y=2.655 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_27_93#_c_101_n VPWR 9.87876e-19 $X=0.27 $Y=2.61 $X2=-0.19 $Y2=-0.245
cc_121 N_A_27_93#_M1011_g N_VPWR_c_384_n 0.00488015f $X=1.275 $Y=2.655 $X2=0
+ $Y2=0
cc_122 N_A_27_93#_M1013_g N_VPWR_c_384_n 0.00510437f $X=1.635 $Y=2.655 $X2=0
+ $Y2=0
cc_123 N_A_27_93#_c_101_n N_VPWR_c_384_n 0.00631118f $X=0.27 $Y=2.61 $X2=0 $Y2=0
cc_124 N_A_M1000_g N_A_342_489#_c_214_n 0.00717896f $X=2.085 $Y=2.655 $X2=0
+ $Y2=0
cc_125 N_A_M1000_g N_A_342_489#_c_215_n 0.0112555f $X=2.085 $Y=2.655 $X2=0 $Y2=0
cc_126 N_A_M1010_g N_A_342_489#_c_215_n 0.0118511f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_127 N_A_c_161_n N_A_342_489#_c_215_n 9.9437e-19 $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_128 N_A_c_164_n N_A_342_489#_c_215_n 0.0443923f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_129 N_A_c_159_n N_A_342_489#_c_206_n 0.00656473f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_160_n N_A_342_489#_c_206_n 0.00111161f $X=2.02 $Y=1.145 $X2=0 $Y2=0
cc_131 N_A_c_161_n N_A_342_489#_c_207_n 0.00949144f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_132 N_A_c_164_n N_A_342_489#_c_207_n 0.0266037f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_133 N_A_c_156_n N_A_342_489#_c_208_n 0.00403612f $X=2.055 $Y=1.315 $X2=0
+ $Y2=0
cc_134 N_A_c_160_n N_A_342_489#_c_208_n 0.00634201f $X=2.02 $Y=1.145 $X2=0 $Y2=0
cc_135 N_A_c_161_n N_A_342_489#_c_208_n 0.00511378f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_136 N_A_c_164_n N_A_342_489#_c_208_n 0.0177261f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_137 N_A_c_156_n N_A_342_489#_c_210_n 0.00198796f $X=2.055 $Y=1.315 $X2=0
+ $Y2=0
cc_138 N_A_M1010_g N_A_342_489#_c_210_n 0.00248423f $X=2.445 $Y=2.655 $X2=0
+ $Y2=0
cc_139 N_A_c_161_n N_A_342_489#_c_210_n 0.00356425f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_140 N_A_c_164_n N_A_342_489#_c_210_n 0.0305846f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_141 N_A_M1010_g N_A_342_489#_c_211_n 0.032745f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_142 N_A_c_161_n N_A_342_489#_c_211_n 0.0217991f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_143 N_A_c_164_n N_A_342_489#_c_211_n 6.78031e-19 $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_144 N_A_M1010_g N_KAPWR_c_280_n 0.00925984f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_145 N_A_M1000_g N_KAPWR_c_281_n 0.00522532f $X=2.085 $Y=2.655 $X2=0 $Y2=0
cc_146 N_A_M1010_g N_KAPWR_c_281_n 0.00605929f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_147 N_A_c_159_n N_VGND_c_341_n 0.00161762f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_c_159_n N_VGND_c_342_n 0.00333051f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_c_159_n N_VGND_c_344_n 0.00510437f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_c_159_n N_VGND_c_346_n 0.00515964f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_M1000_g VPWR 0.00310524f $X=2.085 $Y=2.655 $X2=-0.19 $Y2=-0.245
cc_152 N_A_M1010_g VPWR 0.00310524f $X=2.445 $Y=2.655 $X2=-0.19 $Y2=-0.245
cc_153 N_A_M1000_g N_VPWR_c_384_n 0.00510437f $X=2.085 $Y=2.655 $X2=0 $Y2=0
cc_154 N_A_M1010_g N_VPWR_c_384_n 0.00510437f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_155 N_A_342_489#_c_215_n N_KAPWR_M1010_d 0.00855785f $X=2.82 $Y=2.04 $X2=0
+ $Y2=0
cc_156 N_A_342_489#_c_214_n N_KAPWR_c_279_n 0.00541814f $X=1.87 $Y=2.61 $X2=0
+ $Y2=0
cc_157 N_A_342_489#_M1008_g N_KAPWR_c_280_n 0.0161766f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A_342_489#_M1009_g N_KAPWR_c_280_n 0.00243443f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A_342_489#_c_214_n N_KAPWR_c_280_n 0.00724646f $X=1.87 $Y=2.61 $X2=0
+ $Y2=0
cc_160 N_A_342_489#_c_215_n N_KAPWR_c_280_n 0.0261057f $X=2.82 $Y=2.04 $X2=0
+ $Y2=0
cc_161 N_A_342_489#_M1013_d N_KAPWR_c_281_n 0.0025361f $X=1.71 $Y=2.445 $X2=0
+ $Y2=0
cc_162 N_A_342_489#_M1008_g N_KAPWR_c_281_n 0.0032244f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_342_489#_M1009_g N_KAPWR_c_281_n 0.00939325f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_342_489#_c_214_n N_KAPWR_c_281_n 0.0265285f $X=1.87 $Y=2.61 $X2=0
+ $Y2=0
cc_165 N_A_342_489#_c_215_n N_KAPWR_c_281_n 0.0293845f $X=2.82 $Y=2.04 $X2=0
+ $Y2=0
cc_166 N_A_342_489#_c_215_n A_602_367# 0.00216169f $X=2.82 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_167 N_A_342_489#_c_205_n N_X_c_328_n 0.032978f $X=3.295 $Y=1.005 $X2=0 $Y2=0
cc_168 N_A_342_489#_c_209_n N_X_c_328_n 0.0185607f $X=3.025 $Y=1.225 $X2=0 $Y2=0
cc_169 N_A_342_489#_c_210_n N_X_c_328_n 0.0538185f $X=3.025 $Y=1.955 $X2=0 $Y2=0
cc_170 N_A_342_489#_c_206_n N_VGND_c_341_n 0.00748572f $X=2.2 $Y=0.72 $X2=0
+ $Y2=0
cc_171 N_A_342_489#_c_204_n N_VGND_c_342_n 0.0132046f $X=2.935 $Y=1.17 $X2=0
+ $Y2=0
cc_172 N_A_342_489#_c_205_n N_VGND_c_342_n 0.00168986f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_173 N_A_342_489#_c_206_n N_VGND_c_342_n 0.0247472f $X=2.2 $Y=0.72 $X2=0 $Y2=0
cc_174 N_A_342_489#_c_207_n N_VGND_c_342_n 0.0219254f $X=2.82 $Y=1.115 $X2=0
+ $Y2=0
cc_175 N_A_342_489#_c_209_n N_VGND_c_342_n 0.00386325f $X=3.025 $Y=1.225 $X2=0
+ $Y2=0
cc_176 N_A_342_489#_c_206_n N_VGND_c_344_n 0.00701182f $X=2.2 $Y=0.72 $X2=0
+ $Y2=0
cc_177 N_A_342_489#_c_204_n N_VGND_c_345_n 0.00424179f $X=2.935 $Y=1.17 $X2=0
+ $Y2=0
cc_178 N_A_342_489#_c_205_n N_VGND_c_345_n 0.00510437f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_179 N_A_342_489#_c_204_n N_VGND_c_346_n 0.0043341f $X=2.935 $Y=1.17 $X2=0
+ $Y2=0
cc_180 N_A_342_489#_c_205_n N_VGND_c_346_n 0.00515964f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_181 N_A_342_489#_c_206_n N_VGND_c_346_n 0.00730097f $X=2.2 $Y=0.72 $X2=0
+ $Y2=0
cc_182 N_A_342_489#_M1008_g VPWR 0.00654919f $X=2.935 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_342_489#_M1009_g VPWR 0.00628702f $X=3.295 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_342_489#_c_214_n VPWR 9.42561e-19 $X=1.87 $Y=2.61 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_342_489#_M1008_g N_VPWR_c_384_n 0.00510997f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A_342_489#_M1009_g N_VPWR_c_384_n 0.00585385f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_342_489#_c_214_n N_VPWR_c_384_n 0.00601718f $X=1.87 $Y=2.61 $X2=0
+ $Y2=0
cc_188 A_112_489# N_KAPWR_c_281_n 0.00237263f $X=0.56 $Y=2.445 $X2=2.7 $Y2=2.775
cc_189 N_KAPWR_c_281_n A_270_489# 0.00236976f $X=2.7 $Y=2.775 $X2=-0.19
+ $Y2=1.655
cc_190 N_KAPWR_c_281_n A_432_489# 0.00269277f $X=2.7 $Y=2.775 $X2=-0.19
+ $Y2=1.655
cc_191 N_KAPWR_c_281_n A_602_367# 0.00387996f $X=2.7 $Y=2.775 $X2=-0.19
+ $Y2=1.655
cc_192 N_KAPWR_c_281_n N_X_M1009_d 0.00127496f $X=2.7 $Y=2.775 $X2=0 $Y2=0
cc_193 N_KAPWR_c_280_n N_X_c_328_n 0.0121272f $X=2.72 $Y=2.38 $X2=0 $Y2=0
cc_194 N_KAPWR_c_281_n N_X_c_328_n 0.0420519f $X=2.7 $Y=2.775 $X2=0 $Y2=0
cc_195 N_KAPWR_M1010_d VPWR 0.00121973f $X=2.52 $Y=2.445 $X2=-0.19 $Y2=1.655
cc_196 N_KAPWR_c_279_n VPWR 0.00340959f $X=1.06 $Y=2.61 $X2=-0.19 $Y2=1.655
cc_197 N_KAPWR_c_280_n VPWR 0.00410258f $X=2.72 $Y=2.38 $X2=-0.19 $Y2=1.655
cc_198 N_KAPWR_c_281_n VPWR 0.340095f $X=2.7 $Y=2.775 $X2=-0.19 $Y2=1.655
cc_199 N_KAPWR_c_279_n N_VPWR_c_384_n 0.0113319f $X=1.06 $Y=2.61 $X2=0 $Y2=0
cc_200 N_KAPWR_c_280_n N_VPWR_c_384_n 0.0249343f $X=2.72 $Y=2.38 $X2=0 $Y2=0
cc_201 N_KAPWR_c_281_n N_VPWR_c_384_n 0.013598f $X=2.7 $Y=2.775 $X2=0 $Y2=0
cc_202 A_602_367# VPWR 0.00190157f $X=3.01 $Y=1.835 $X2=2.06 $Y2=0.465
cc_203 N_X_c_328_n N_VGND_c_345_n 0.0101312f $X=3.51 $Y=0.72 $X2=0 $Y2=0
cc_204 N_X_c_328_n N_VGND_c_346_n 0.0121005f $X=3.51 $Y=0.72 $X2=0 $Y2=0
cc_205 N_X_M1009_d VPWR 0.00135204f $X=3.37 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_206 N_X_c_328_n VPWR 0.00383788f $X=3.51 $Y=0.72 $X2=-0.19 $Y2=-0.245
cc_207 N_X_c_328_n N_VPWR_c_384_n 0.0240782f $X=3.51 $Y=0.72 $X2=0 $Y2=0
