* NGSPICE file created from sky130_fd_sc_lp__invlp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__invlp_2 A VGND VNB VPB VPWR Y
M1000 VPWR A a_116_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=8.064e+11p pd=6.32e+06u as=7.056e+11p ps=6.16e+06u
M1001 VGND A a_116_55# VNB nshort w=840000u l=150000u
+  ad=4.788e+11p pd=4.5e+06u as=5.292e+11p ps=4.62e+06u
M1002 a_116_55# A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1003 a_116_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_116_367# A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1005 Y A a_116_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_116_55# A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A a_116_55# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

