* File: sky130_fd_sc_lp__dfrtp_1.pex.spice
* Created: Wed Sep  2 09:43:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFRTP_1%CLK 3 7 11 12 13 14 18 19
r37 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r38 13 14 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.282 $Y=1.665
+ $X2=0.282 $Y2=2.035
r39 13 19 1.53659 $w=3.73e-07 $l=5e-08 $layer=LI1_cond $X=0.282 $Y=1.665
+ $X2=0.282 $Y2=1.615
r40 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.955
+ $X2=0.385 $Y2=1.615
r41 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.955
+ $X2=0.385 $Y2=2.12
r42 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.45
+ $X2=0.385 $Y2=1.615
r43 7 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.475 $Y=2.63
+ $X2=0.475 $Y2=2.12
r44 3 10 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.475 $Y=0.78
+ $X2=0.475 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%A_27_114# 1 2 8 11 15 18 21 25 27 29 30 33
+ 37 39 40 42 44 46 47 48 50 51 52 54 55 56 59 60 66 67 72 73 76 78 79 80 81 82
+ 83 84 86 87 88 90 92 94
c269 87 0 1.84213e-19 $X=6.2 $Y=1.92
c270 86 0 1.81739e-19 $X=6.2 $Y=1.92
c271 83 0 1.78624e-19 $X=4.835 $Y=0.587
c272 47 0 5.32993e-20 $X=1.655 $Y=0.365
c273 27 0 1.17665e-19 $X=7.01 $Y=0.555
c274 21 0 9.07137e-20 $X=3.19 $Y=2.875
r275 87 97 14.0031 $w=3.27e-07 $l=9.5e-08 $layer=POLY_cond $X=6.2 $Y=1.92
+ $X2=6.295 $Y2=1.92
r276 86 88 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=1.92
+ $X2=6.225 $Y2=1.755
r277 86 87 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.2
+ $Y=1.92 $X2=6.2 $Y2=1.92
r278 83 84 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.835 $Y=0.615
+ $X2=5.505 $Y2=0.615
r279 82 83 22.5367 $w=1.78e-07 $l=3.65e-07 $layer=LI1_cond $X=4.47 $Y=0.587
+ $X2=4.835 $Y2=0.587
r280 79 92 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.265
+ $X2=1.04 $Y2=1.1
r281 78 79 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.995
+ $Y=1.265 $X2=0.995 $Y2=1.265
r282 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.01
+ $Y=0.39 $X2=7.01 $Y2=0.39
r283 70 90 2.66603 $w=3.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.345 $Y=0.39
+ $X2=6.26 $Y2=0.48
r284 70 72 28.3842 $w=2.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.345 $Y=0.39
+ $X2=7.01 $Y2=0.39
r285 68 90 4.14084 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=6.26 $Y=0.705
+ $X2=6.26 $Y2=0.48
r286 68 88 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=6.26 $Y=0.705
+ $X2=6.26 $Y2=1.755
r287 67 84 10.429 $w=4.48e-07 $l=2.25e-07 $layer=LI1_cond $X=5.73 $Y=0.48
+ $X2=5.505 $Y2=0.48
r288 66 90 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.48
+ $X2=6.26 $Y2=0.48
r289 66 67 11.8279 $w=4.48e-07 $l=4.45e-07 $layer=LI1_cond $X=6.175 $Y=0.48
+ $X2=5.73 $Y2=0.48
r290 63 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.395 $Y=0.555
+ $X2=3.31 $Y2=0.555
r291 63 82 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=3.395 $Y=0.555
+ $X2=4.47 $Y2=0.555
r292 60 95 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.287 $Y=1.44
+ $X2=3.287 $Y2=1.605
r293 60 94 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.287 $Y=1.44
+ $X2=3.287 $Y2=1.275
r294 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.31
+ $Y=1.44 $X2=3.31 $Y2=1.44
r295 57 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=0.64
+ $X2=3.31 $Y2=0.555
r296 57 59 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.31 $Y=0.64 $X2=3.31
+ $Y2=1.44
r297 55 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=0.555
+ $X2=3.31 $Y2=0.555
r298 55 56 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.225 $Y=0.555
+ $X2=2.685 $Y2=0.555
r299 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.6 $Y=0.64
+ $X2=2.685 $Y2=0.555
r300 53 54 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.6 $Y=0.64
+ $X2=2.6 $Y2=1.175
r301 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.515 $Y=1.26
+ $X2=2.6 $Y2=1.175
r302 51 52 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.515 $Y=1.26
+ $X2=1.825 $Y2=1.26
r303 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.74 $Y=1.175
+ $X2=1.825 $Y2=1.26
r304 49 50 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.74 $Y=0.45
+ $X2=1.74 $Y2=1.175
r305 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.655 $Y=0.365
+ $X2=1.74 $Y2=0.45
r306 47 48 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.655 $Y=0.365
+ $X2=1.125 $Y2=0.365
r307 46 78 3.17288 $w=3.15e-07 $l=1.84594e-07 $layer=LI1_cond $X=1.04 $Y=1.1
+ $X2=0.895 $Y2=1.19
r308 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.04 $Y=0.45
+ $X2=1.125 $Y2=0.365
r309 45 46 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.04 $Y=0.45
+ $X2=1.04 $Y2=1.1
r310 44 80 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.75 $Y=2.3
+ $X2=0.75 $Y2=1.77
r311 42 80 10.9702 $w=4.58e-07 $l=2.3e-07 $layer=LI1_cond $X=0.895 $Y=1.54
+ $X2=0.895 $Y2=1.77
r312 41 78 3.17288 $w=3.15e-07 $l=9e-08 $layer=LI1_cond $X=0.895 $Y=1.28
+ $X2=0.895 $Y2=1.19
r313 41 42 6.76044 $w=4.58e-07 $l=2.6e-07 $layer=LI1_cond $X=0.895 $Y=1.28
+ $X2=0.895 $Y2=1.54
r314 39 78 3.41642 $w=1.8e-07 $l=2.3e-07 $layer=LI1_cond $X=0.665 $Y=1.19
+ $X2=0.895 $Y2=1.19
r315 39 40 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=0.665 $Y=1.19
+ $X2=0.425 $Y2=1.19
r316 38 76 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.355 $Y=2.385
+ $X2=0.225 $Y2=2.385
r317 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=2.385
+ $X2=0.75 $Y2=2.3
r318 37 38 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.665 $Y=2.385
+ $X2=0.355 $Y2=2.385
r319 31 40 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.26 $Y=1.1
+ $X2=0.425 $Y2=1.19
r320 31 33 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=1.1
+ $X2=0.26 $Y2=0.785
r321 27 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.01 $Y=0.555
+ $X2=7.01 $Y2=0.39
r322 27 29 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.01 $Y=0.555
+ $X2=7.01 $Y2=0.875
r323 23 97 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.295 $Y=2.085
+ $X2=6.295 $Y2=1.92
r324 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.295 $Y=2.085
+ $X2=6.295 $Y2=2.665
r325 21 95 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=3.19 $Y=2.875
+ $X2=3.19 $Y2=1.605
r326 18 94 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.175 $Y=0.955
+ $X2=3.175 $Y2=1.275
r327 15 92 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.175 $Y=0.78
+ $X2=1.175 $Y2=1.1
r328 11 30 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.905 $Y=2.63
+ $X2=0.905 $Y2=1.77
r329 8 30 52.1105 $w=4.2e-07 $l=2.1e-07 $layer=POLY_cond $X=1.04 $Y=1.56
+ $X2=1.04 $Y2=1.77
r330 7 79 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=1.04 $Y=1.31
+ $X2=1.04 $Y2=1.265
r331 7 8 33.1044 $w=4.2e-07 $l=2.5e-07 $layer=POLY_cond $X=1.04 $Y=1.31 $X2=1.04
+ $Y2=1.56
r332 2 76 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.31 $X2=0.26 $Y2=2.465
r333 1 33 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.57 $X2=0.26 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%D 3 7 9 13 14
c42 14 0 2.5562e-19 $X=2.38 $Y=1.67
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.67 $X2=2.38 $Y2=1.67
r44 11 13 17.4919 $w=2.48e-07 $l=9e-08 $layer=POLY_cond $X=2.29 $Y=1.67 $X2=2.38
+ $Y2=1.67
r45 9 14 7.80115 $w=3.23e-07 $l=2.2e-07 $layer=LI1_cond $X=2.16 $Y=1.677
+ $X2=2.38 $Y2=1.677
r46 5 13 70.9395 $w=2.48e-07 $l=4.39829e-07 $layer=POLY_cond $X=2.745 $Y=1.505
+ $X2=2.38 $Y2=1.67
r47 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.745 $Y=1.505
+ $X2=2.745 $Y2=0.955
r48 1 11 14.534 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.835
+ $X2=2.29 $Y2=1.67
r49 1 3 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.29 $Y=1.835
+ $X2=2.29 $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%A_196_462# 1 2 9 13 17 19 20 23 28 31 35 39
+ 40 42 44 45 47 48 49 50 59 63 64 79
c198 64 0 2.50656e-19 $X=6.96 $Y=1.71
c199 50 0 2.63988e-19 $X=3.745 $Y=2.035
c200 47 0 2.57019e-20 $X=3.455 $Y=2.035
c201 42 0 4.17781e-20 $X=3.85 $Y=1.875
c202 19 0 1.84213e-19 $X=6.575 $Y=1.44
r203 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.96
+ $Y=1.71 $X2=6.96 $Y2=1.71
r204 60 64 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=6.96 $Y=2.035
+ $X2=6.96 $Y2=1.71
r205 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=2.035
+ $X2=6.96 $Y2=2.035
r206 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=2.035
+ $X2=3.6 $Y2=2.035
r207 53 75 1.31291 $w=3.93e-07 $l=4.5e-08 $layer=LI1_cond $X=1.2 $Y=2.137
+ $X2=1.155 $Y2=2.137
r208 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r209 50 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=2.035
+ $X2=3.6 $Y2=2.035
r210 49 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=6.96 $Y2=2.035
r211 49 50 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=3.745 $Y2=2.035
r212 48 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r213 47 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.455 $Y=2.035
+ $X2=3.6 $Y2=2.035
r214 47 48 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=3.455 $Y=2.035
+ $X2=1.345 $Y2=2.035
r215 45 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.85 $Y=1.47
+ $X2=3.85 $Y2=1.305
r216 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.85
+ $Y=1.47 $X2=3.85 $Y2=1.47
r217 42 57 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.85 $Y=2.027
+ $X2=3.6 $Y2=2.027
r218 42 44 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.85 $Y=1.875
+ $X2=3.85 $Y2=1.47
r219 40 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=2.24
+ $X2=2.74 $Y2=2.405
r220 39 79 69.5955 $w=1.98e-07 $l=1.255e-06 $layer=LI1_cond $X=2.74 $Y=2.235
+ $X2=1.485 $Y2=2.235
r221 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=2.24 $X2=2.74 $Y2=2.24
r222 33 79 5.57506 $w=3.93e-07 $l=9.5e-08 $layer=LI1_cond $X=1.39 $Y=2.137
+ $X2=1.485 $Y2=2.137
r223 33 53 5.5434 $w=3.93e-07 $l=1.9e-07 $layer=LI1_cond $X=1.39 $Y=2.137
+ $X2=1.2 $Y2=2.137
r224 33 35 67.4211 $w=1.88e-07 $l=1.155e-06 $layer=LI1_cond $X=1.39 $Y=1.94
+ $X2=1.39 $Y2=0.785
r225 29 75 3.18482 $w=2.6e-07 $l=1.98e-07 $layer=LI1_cond $X=1.155 $Y=2.335
+ $X2=1.155 $Y2=2.137
r226 29 31 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=1.155 $Y=2.335
+ $X2=1.155 $Y2=2.455
r227 27 63 46.1022 $w=3.8e-07 $l=3.15e-07 $layer=POLY_cond $X=6.935 $Y=2.025
+ $X2=6.935 $Y2=1.71
r228 27 28 48.9106 $w=3.8e-07 $l=1.9e-07 $layer=POLY_cond $X=6.935 $Y=2.025
+ $X2=6.935 $Y2=2.215
r229 26 63 2.19534 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=6.935 $Y=1.695
+ $X2=6.935 $Y2=1.71
r230 23 28 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.82 $Y=2.795
+ $X2=6.82 $Y2=2.215
r231 19 26 90.2297 $w=1.99e-07 $l=4.09145e-07 $layer=POLY_cond $X=6.575 $Y=1.44
+ $X2=6.935 $Y2=1.545
r232 19 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.575 $Y=1.44
+ $X2=6.235 $Y2=1.44
r233 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.16 $Y=1.365
+ $X2=6.235 $Y2=1.44
r234 15 17 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.16 $Y=1.365 $X2=6.16
+ $Y2=0.765
r235 13 69 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.94 $Y=0.955
+ $X2=3.94 $Y2=1.305
r236 9 67 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.72 $Y=2.875 $X2=2.72
+ $Y2=2.405
r237 2 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.31 $X2=1.12 $Y2=2.455
r238 1 35 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.25
+ $Y=0.57 $X2=1.39 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%A_695_375# 1 2 9 11 12 15 19 20 23 25 27 28
+ 33 36 40
c107 27 0 3.29571e-19 $X=4.39 $Y=1.52
c108 12 0 9.05148e-20 $X=3.625 $Y=1.95
c109 9 0 1.84048e-19 $X=3.55 $Y=2.875
r110 37 40 10.2591 $w=1.98e-07 $l=1.85e-07 $layer=LI1_cond $X=5.85 $Y=2.365
+ $X2=6.035 $Y2=2.365
r111 33 35 4.08188 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=5.83 $Y=0.96
+ $X2=5.83 $Y2=1.065
r112 27 30 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=4.39 $Y=1.52 $X2=4.39
+ $Y2=1.58
r113 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.39
+ $Y=1.52 $X2=4.39 $Y2=1.52
r114 25 37 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.85 $Y=2.265 $X2=5.85
+ $Y2=2.365
r115 24 36 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=5.85 $Y=1.665
+ $X2=5.8 $Y2=1.58
r116 24 25 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.85 $Y=1.665
+ $X2=5.85 $Y2=2.265
r117 23 36 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=1.495 $X2=5.8
+ $Y2=1.58
r118 23 35 18.3537 $w=2.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.8 $Y=1.495
+ $X2=5.8 $Y2=1.065
r119 21 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.555 $Y=1.58
+ $X2=4.39 $Y2=1.58
r120 20 36 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.665 $Y=1.58
+ $X2=5.8 $Y2=1.58
r121 20 21 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=5.665 $Y=1.58
+ $X2=4.555 $Y2=1.58
r122 19 28 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.39 $Y=1.875
+ $X2=4.39 $Y2=1.52
r123 18 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.39 $Y=1.355
+ $X2=4.39 $Y2=1.52
r124 15 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.3 $Y=0.955 $X2=4.3
+ $Y2=1.355
r125 11 19 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.225 $Y=1.95
+ $X2=4.39 $Y2=1.875
r126 11 12 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.225 $Y=1.95
+ $X2=3.625 $Y2=1.95
r127 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.55 $Y=2.025
+ $X2=3.625 $Y2=1.95
r128 7 9 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=3.55 $Y=2.025
+ $X2=3.55 $Y2=2.875
r129 2 40 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=5.825
+ $Y=2.255 $X2=6.035 $Y2=2.38
r130 1 33 182 $w=1.7e-07 $l=7.61906e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.315 $X2=5.83 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%RESET_B 3 5 6 9 11 13 15 16 17 21 24 28 30
+ 32 33 35 37 38 40 41 45 49 58 59 63
c187 58 0 1.05907e-19 $X=7.98 $Y=1.72
c188 17 0 4.17781e-20 $X=4.16 $Y=2.47
c189 16 0 1.85329e-19 $X=4.585 $Y=2.47
c190 9 0 2.18205e-19 $X=2.385 $Y=0.955
r191 61 63 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=7.395 $Y=1.72
+ $X2=7.44 $Y2=1.72
r192 57 59 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=7.98 $Y=1.72
+ $X2=8.11 $Y2=1.72
r193 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.98
+ $Y=1.72 $X2=7.98 $Y2=1.72
r194 54 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.89 $Y=1.72 $X2=7.98
+ $Y2=1.72
r195 49 61 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=1.72
+ $X2=7.395 $Y2=1.72
r196 49 58 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=7.46 $Y=1.72
+ $X2=7.98 $Y2=1.72
r197 49 63 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=7.46 $Y=1.72 $X2=7.44
+ $Y2=1.72
r198 45 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.85 $Y=2.72
+ $X2=5.85 $Y2=2.99
r199 40 43 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.75 $Y=2.56
+ $X2=4.75 $Y2=2.72
r200 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.75
+ $Y=2.56 $X2=4.75 $Y2=2.56
r201 37 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.31 $Y=1.885
+ $X2=7.31 $Y2=1.72
r202 37 38 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.31 $Y=1.885
+ $X2=7.31 $Y2=2.905
r203 36 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.935 $Y=2.99
+ $X2=5.85 $Y2=2.99
r204 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.225 $Y=2.99
+ $X2=7.31 $Y2=2.905
r205 35 36 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=7.225 $Y=2.99
+ $X2=5.935 $Y2=2.99
r206 34 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.915 $Y=2.72
+ $X2=4.75 $Y2=2.72
r207 33 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=5.85 $Y2=2.72
r208 33 34 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=4.915 $Y2=2.72
r209 31 41 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.75 $Y=2.545
+ $X2=4.75 $Y2=2.56
r210 31 32 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.75 $Y=2.545
+ $X2=4.75 $Y2=2.47
r211 26 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.11 $Y=1.885
+ $X2=8.11 $Y2=1.72
r212 26 28 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=8.11 $Y=1.885
+ $X2=8.11 $Y2=2.795
r213 22 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.89 $Y=1.555
+ $X2=7.89 $Y2=1.72
r214 22 24 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.89 $Y=1.555
+ $X2=7.89 $Y2=0.875
r215 19 32 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.84 $Y=2.395
+ $X2=4.75 $Y2=2.47
r216 19 21 846.064 $w=1.5e-07 $l=1.65e-06 $layer=POLY_cond $X=4.84 $Y=2.395
+ $X2=4.84 $Y2=0.745
r217 18 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.84 $Y=0.375
+ $X2=4.84 $Y2=0.745
r218 16 32 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.585 $Y=2.47
+ $X2=4.75 $Y2=2.47
r219 16 17 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.585 $Y=2.47
+ $X2=4.16 $Y2=2.47
r220 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.085 $Y=2.545
+ $X2=4.16 $Y2=2.47
r221 13 15 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.085 $Y=2.545
+ $X2=4.085 $Y2=2.875
r222 12 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.46 $Y=0.3
+ $X2=2.385 $Y2=0.3
r223 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.765 $Y=0.3
+ $X2=4.84 $Y2=0.375
r224 11 12 1181.93 $w=1.5e-07 $l=2.305e-06 $layer=POLY_cond $X=4.765 $Y=0.3
+ $X2=2.46 $Y2=0.3
r225 7 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.385 $Y=0.375
+ $X2=2.385 $Y2=0.3
r226 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.385 $Y=0.375
+ $X2=2.385 $Y2=0.955
r227 5 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.31 $Y=0.3
+ $X2=2.385 $Y2=0.3
r228 5 6 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.31 $Y=0.3
+ $X2=1.935 $Y2=0.3
r229 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.86 $Y=0.375
+ $X2=1.935 $Y2=0.3
r230 1 3 1281.91 $w=1.5e-07 $l=2.5e-06 $layer=POLY_cond $X=1.86 $Y=0.375
+ $X2=1.86 $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%A_559_533# 1 2 3 12 14 15 19 21 26 27 31 32
+ 33 37 40 41 42 43 44 45 52 53 60 63
c151 42 0 1.19746e-19 $X=4.415 $Y=2.21
c152 15 0 1.81739e-19 $X=5.675 $Y=2.02
c153 12 0 1.78624e-19 $X=5.5 $Y=1.065
r154 53 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.32 $Y=1.93 $X2=5.32
+ $Y2=2.02
r155 53 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=1.93
+ $X2=5.32 $Y2=1.765
r156 52 55 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=5.32 $Y=1.93
+ $X2=5.32 $Y2=2.21
r157 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.32
+ $Y=1.93 $X2=5.32 $Y2=1.93
r158 49 60 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.32 $Y=1.23 $X2=5.5
+ $Y2=1.23
r159 49 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.32 $Y=1.23 $X2=5.23
+ $Y2=1.23
r160 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.32
+ $Y=1.23 $X2=5.32 $Y2=1.23
r161 45 48 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=5.32 $Y=1.035
+ $X2=5.32 $Y2=1.23
r162 41 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=2.21
+ $X2=5.32 $Y2=2.21
r163 41 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.155 $Y=2.21
+ $X2=4.415 $Y2=2.21
r164 40 44 3.77418 $w=2.45e-07 $l=9.66954e-08 $layer=LI1_cond $X=4.305 $Y=2.445
+ $X2=4.28 $Y2=2.53
r165 39 42 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.305 $Y=2.295
+ $X2=4.415 $Y2=2.21
r166 39 40 7.85757 $w=2.18e-07 $l=1.5e-07 $layer=LI1_cond $X=4.305 $Y=2.295
+ $X2=4.305 $Y2=2.445
r167 35 44 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=2.615
+ $X2=4.28 $Y2=2.53
r168 35 37 10.8842 $w=2.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.28 $Y=2.615
+ $X2=4.28 $Y2=2.87
r169 33 45 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=1.035
+ $X2=5.32 $Y2=1.035
r170 33 43 53.342 $w=2.08e-07 $l=1.01e-06 $layer=LI1_cond $X=5.155 $Y=1.035
+ $X2=4.145 $Y2=1.035
r171 31 44 2.68609 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.145 $Y=2.53
+ $X2=4.28 $Y2=2.53
r172 31 32 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.145 $Y=2.53
+ $X2=3.585 $Y2=2.53
r173 27 43 7.28026 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.98 $Y=0.975
+ $X2=4.145 $Y2=0.975
r174 27 29 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.98 $Y=0.975
+ $X2=3.68 $Y2=0.975
r175 25 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.5 $Y=2.615
+ $X2=3.585 $Y2=2.53
r176 25 26 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.5 $Y=2.615
+ $X2=3.5 $Y2=2.845
r177 21 26 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.415 $Y=2.96
+ $X2=3.5 $Y2=2.845
r178 21 23 22.0467 $w=2.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.415 $Y=2.96
+ $X2=2.975 $Y2=2.96
r179 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.75 $Y=2.095
+ $X2=5.75 $Y2=2.675
r180 16 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.485 $Y=2.02
+ $X2=5.32 $Y2=2.02
r181 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.675 $Y=2.02
+ $X2=5.75 $Y2=2.095
r182 15 16 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.675 $Y=2.02
+ $X2=5.485 $Y2=2.02
r183 12 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.5 $Y=1.065
+ $X2=5.5 $Y2=1.23
r184 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.5 $Y=1.065
+ $X2=5.5 $Y2=0.635
r185 10 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.23 $Y=1.395
+ $X2=5.23 $Y2=1.23
r186 10 63 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.23 $Y=1.395
+ $X2=5.23 $Y2=1.765
r187 3 37 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=2.665 $X2=4.3 $Y2=2.87
r188 2 23 600 $w=1.7e-07 $l=3.6404e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=2.665 $X2=2.975 $Y2=2.95
r189 1 29 182 $w=1.7e-07 $l=5.32729e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.745 $X2=3.68 $Y2=0.975
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%A_1467_419# 1 2 9 13 15 18 22 24 28 31 32
c78 18 0 1.32991e-19 $X=7.66 $Y=2.26
r79 33 35 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=7.41 $Y=2.26 $X2=7.46
+ $Y2=2.26
r80 30 31 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=8.91 $Y=1.025
+ $X2=8.91 $Y2=2.095
r81 29 32 6.07544 $w=2.5e-07 $l=1.88809e-07 $layer=LI1_cond $X=8.465 $Y=2.18
+ $X2=8.312 $Y2=2.26
r82 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.825 $Y=2.18
+ $X2=8.91 $Y2=2.095
r83 28 29 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.825 $Y=2.18
+ $X2=8.465 $Y2=2.18
r84 24 30 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.825 $Y=0.86
+ $X2=8.91 $Y2=1.025
r85 24 26 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=8.825 $Y=0.86
+ $X2=8.465 $Y2=0.86
r86 20 32 0.637292 $w=3.05e-07 $l=1.65e-07 $layer=LI1_cond $X=8.312 $Y=2.425
+ $X2=8.312 $Y2=2.26
r87 20 22 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=8.312 $Y=2.425
+ $X2=8.312 $Y2=2.795
r88 18 35 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=7.66 $Y=2.26 $X2=7.46
+ $Y2=2.26
r89 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.66
+ $Y=2.26 $X2=7.66 $Y2=2.26
r90 15 32 6.07544 $w=2.5e-07 $l=1.52e-07 $layer=LI1_cond $X=8.16 $Y=2.26
+ $X2=8.312 $Y2=2.26
r91 15 17 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=8.16 $Y=2.26 $X2=7.66
+ $Y2=2.26
r92 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=2.095
+ $X2=7.46 $Y2=2.26
r93 11 13 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=7.46 $Y=2.095
+ $X2=7.46 $Y2=0.875
r94 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.41 $Y=2.425
+ $X2=7.41 $Y2=2.26
r95 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.41 $Y=2.425 $X2=7.41
+ $Y2=2.795
r96 2 22 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.185
+ $Y=2.585 $X2=8.325 $Y2=2.795
r97 1 26 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=8.325
+ $Y=0.665 $X2=8.465 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%A_1247_89# 1 2 7 9 12 14 16 18 22 25 27 31
+ 35 40 41 43 45 46
c115 16 0 9.41644e-20 $X=9.5 $Y=1.345
c116 12 0 1.05907e-19 $X=8.54 $Y=2.795
r117 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.56
+ $Y=1.36 $X2=8.56 $Y2=1.36
r118 40 41 13.0916 $w=3.23e-07 $l=3.05e-07 $layer=LI1_cond $X=6.532 $Y=2.57
+ $X2=6.532 $Y2=2.265
r119 36 43 2.28545 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.775 $Y=1.28
+ $X2=6.645 $Y2=1.28
r120 35 45 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.395 $Y=1.28
+ $X2=8.525 $Y2=1.28
r121 35 36 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=8.395 $Y=1.28
+ $X2=6.775 $Y2=1.28
r122 33 43 4.14756 $w=2.2e-07 $l=1.03078e-07 $layer=LI1_cond $X=6.605 $Y=1.365
+ $X2=6.645 $Y2=1.28
r123 33 41 55.4545 $w=1.78e-07 $l=9e-07 $layer=LI1_cond $X=6.605 $Y=1.365
+ $X2=6.605 $Y2=2.265
r124 29 43 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=1.195
+ $X2=6.645 $Y2=1.28
r125 29 31 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=6.645 $Y=1.195
+ $X2=6.645 $Y2=0.86
r126 26 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.56 $Y=1.7
+ $X2=8.56 $Y2=1.36
r127 26 27 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.56 $Y=1.7
+ $X2=8.56 $Y2=1.865
r128 24 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.56 $Y=1.345
+ $X2=8.56 $Y2=1.36
r129 24 25 13.5877 $w=2.4e-07 $l=1.42653e-07 $layer=POLY_cond $X=8.56 $Y=1.345
+ $X2=8.45 $Y2=1.27
r130 20 28 89.3387 $w=1.78e-07 $l=3.43475e-07 $layer=POLY_cond $X=9.575 $Y=0.945
+ $X2=9.537 $Y2=1.27
r131 20 22 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.575 $Y=0.945
+ $X2=9.575 $Y2=0.595
r132 16 28 21.642 $w=1.78e-07 $l=9.16515e-08 $layer=POLY_cond $X=9.5 $Y=1.345
+ $X2=9.537 $Y2=1.27
r133 16 18 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.5 $Y=1.345 $X2=9.5
+ $Y2=2.155
r134 15 25 12.1617 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=8.725 $Y=1.27
+ $X2=8.45 $Y2=1.27
r135 14 28 6.87779 $w=1.5e-07 $l=1.12e-07 $layer=POLY_cond $X=9.425 $Y=1.27
+ $X2=9.537 $Y2=1.27
r136 14 15 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=9.425 $Y=1.27
+ $X2=8.725 $Y2=1.27
r137 12 27 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=8.54 $Y=2.795
+ $X2=8.54 $Y2=1.865
r138 7 25 13.5877 $w=2.4e-07 $l=2.34521e-07 $layer=POLY_cond $X=8.25 $Y=1.195
+ $X2=8.45 $Y2=1.27
r139 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.25 $Y=1.195
+ $X2=8.25 $Y2=0.875
r140 2 40 600 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_PDIFF $count=1 $X=6.37
+ $Y=2.245 $X2=6.51 $Y2=2.57
r141 1 31 182 $w=1.7e-07 $l=5.72582e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.445 $X2=6.61 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%A_1832_367# 1 2 9 13 16 20 24 25 27 29
c47 27 0 9.41644e-20 $X=9.345 $Y=1.5
r48 25 30 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.972 $Y=1.5
+ $X2=9.972 $Y2=1.665
r49 25 29 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.972 $Y=1.5
+ $X2=9.972 $Y2=1.335
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.95
+ $Y=1.5 $X2=9.95 $Y2=1.5
r51 22 27 0.911997 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=9.525 $Y=1.5
+ $X2=9.345 $Y2=1.5
r52 22 24 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=9.525 $Y=1.5
+ $X2=9.95 $Y2=1.5
r53 18 27 5.7047 $w=2.92e-07 $l=1.96074e-07 $layer=LI1_cond $X=9.277 $Y=1.665
+ $X2=9.345 $Y2=1.5
r54 18 20 16.3903 $w=2.23e-07 $l=3.2e-07 $layer=LI1_cond $X=9.277 $Y=1.665
+ $X2=9.277 $Y2=1.985
r55 14 27 5.7047 $w=2.92e-07 $l=1.65e-07 $layer=LI1_cond $X=9.345 $Y=1.335
+ $X2=9.345 $Y2=1.5
r56 14 16 23.6891 $w=3.58e-07 $l=7.4e-07 $layer=LI1_cond $X=9.345 $Y=1.335
+ $X2=9.345 $Y2=0.595
r57 13 29 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.085 $Y=0.805
+ $X2=10.085 $Y2=1.335
r58 9 30 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=10.01 $Y=2.465
+ $X2=10.01 $Y2=1.665
r59 2 20 300 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=2 $X=9.16
+ $Y=1.835 $X2=9.285 $Y2=1.985
r60 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.235
+ $Y=0.385 $X2=9.36 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 49 50
+ 52 53 55 56 57 59 64 73 87 93 94 97 100 103 110
r139 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r140 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r141 103 106 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.42 $Y=3.07
+ $X2=5.42 $Y2=3.33
r142 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r143 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r144 94 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r145 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r146 91 110 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=9.96 $Y=3.33
+ $X2=9.772 $Y2=3.33
r147 91 93 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.96 $Y=3.33
+ $X2=10.32 $Y2=3.33
r148 90 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r149 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r150 87 110 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=9.585 $Y=3.33
+ $X2=9.772 $Y2=3.33
r151 87 89 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=9.585 $Y=3.33
+ $X2=9.36 $Y2=3.33
r152 86 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r153 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r154 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 83 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=5.52 $Y2=3.33
r156 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r157 80 106 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.585 $Y=3.33
+ $X2=5.42 $Y2=3.33
r158 80 82 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=5.585 $Y=3.33
+ $X2=7.44 $Y2=3.33
r159 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r160 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r161 75 78 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r162 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r163 73 106 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.255 $Y=3.33
+ $X2=5.42 $Y2=3.33
r164 73 78 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.255 $Y=3.33
+ $X2=5.04 $Y2=3.33
r165 72 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r166 72 101 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.16 $Y2=3.33
r167 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r168 69 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=3.33
+ $X2=2.075 $Y2=3.33
r169 69 71 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.24 $Y=3.33
+ $X2=3.6 $Y2=3.33
r170 68 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r171 68 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r172 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r173 65 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r174 65 67 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r175 64 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=3.33
+ $X2=2.075 $Y2=3.33
r176 64 67 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.91 $Y=3.33
+ $X2=1.68 $Y2=3.33
r177 62 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r178 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r179 59 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r180 59 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r181 57 107 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r182 57 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r183 55 85 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.635 $Y=3.33
+ $X2=8.4 $Y2=3.33
r184 55 56 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=8.635 $Y=3.33
+ $X2=8.777 $Y2=3.33
r185 54 89 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=8.92 $Y=3.33
+ $X2=9.36 $Y2=3.33
r186 54 56 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=8.92 $Y=3.33
+ $X2=8.777 $Y2=3.33
r187 52 82 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.565 $Y=3.33
+ $X2=7.44 $Y2=3.33
r188 52 53 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.565 $Y=3.33
+ $X2=7.735 $Y2=3.33
r189 51 85 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=8.4 $Y2=3.33
r190 51 53 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=7.735 $Y2=3.33
r191 49 71 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.6 $Y2=3.33
r192 49 50 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.865 $Y2=3.33
r193 48 75 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.975 $Y=3.33
+ $X2=4.08 $Y2=3.33
r194 48 50 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.975 $Y=3.33
+ $X2=3.865 $Y2=3.33
r195 44 47 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=9.772 $Y=2.01
+ $X2=9.772 $Y2=2.49
r196 42 110 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.772 $Y=3.245
+ $X2=9.772 $Y2=3.33
r197 42 47 23.2025 $w=3.73e-07 $l=7.55e-07 $layer=LI1_cond $X=9.772 $Y=3.245
+ $X2=9.772 $Y2=2.49
r198 38 56 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=8.777 $Y=3.245
+ $X2=8.777 $Y2=3.33
r199 38 40 18.1965 $w=2.83e-07 $l=4.5e-07 $layer=LI1_cond $X=8.777 $Y=3.245
+ $X2=8.777 $Y2=2.795
r200 34 53 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.735 $Y=3.245
+ $X2=7.735 $Y2=3.33
r201 34 36 15.2529 $w=3.38e-07 $l=4.5e-07 $layer=LI1_cond $X=7.735 $Y=3.245
+ $X2=7.735 $Y2=2.795
r202 30 50 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=3.245
+ $X2=3.865 $Y2=3.33
r203 30 32 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=3.865 $Y=3.245
+ $X2=3.865 $Y2=2.96
r204 26 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=3.245
+ $X2=2.075 $Y2=3.33
r205 26 28 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.075 $Y=3.245
+ $X2=2.075 $Y2=2.96
r206 22 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r207 22 24 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.76
r208 7 47 300 $w=1.7e-07 $l=7.5705e-07 $layer=licon1_PDIFF $count=2 $X=9.575
+ $Y=1.835 $X2=9.795 $Y2=2.49
r209 7 44 600 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=9.575
+ $Y=1.835 $X2=9.75 $Y2=2.01
r210 6 40 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.615
+ $Y=2.585 $X2=8.755 $Y2=2.795
r211 5 36 600 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_PDIFF $count=1 $X=7.485
+ $Y=2.585 $X2=7.74 $Y2=2.795
r212 4 103 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.275
+ $Y=2.255 $X2=5.42 $Y2=3.07
r213 3 32 600 $w=1.7e-07 $l=3.89776e-07 $layer=licon1_PDIFF $count=1 $X=3.625
+ $Y=2.665 $X2=3.845 $Y2=2.96
r214 2 28 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=2.665 $X2=2.075 $Y2=2.96
r215 1 24 600 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.31 $X2=0.69 $Y2=2.76
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%A_304_533# 1 2 3 12 14 15 18 20 24 27 28 31
c73 31 0 9.05148e-20 $X=3.16 $Y=1.87
c74 20 0 1.84048e-19 $X=3.075 $Y=2.59
c75 15 0 2.57019e-20 $X=1.74 $Y=2.59
r76 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=1.955
+ $X2=3.16 $Y2=1.87
r77 26 27 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.16 $Y=1.955
+ $X2=3.16 $Y2=2.505
r78 22 31 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.955 $Y=1.87
+ $X2=3.16 $Y2=1.87
r79 22 24 44.9182 $w=1.98e-07 $l=8.1e-07 $layer=LI1_cond $X=2.955 $Y=1.785
+ $X2=2.955 $Y2=0.975
r80 21 28 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=2.59
+ $X2=2.525 $Y2=2.59
r81 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.075 $Y=2.59
+ $X2=3.16 $Y2=2.505
r82 20 21 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.075 $Y=2.59
+ $X2=2.64 $Y2=2.59
r83 16 28 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=2.675
+ $X2=2.525 $Y2=2.59
r84 16 18 9.77071 $w=2.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.525 $Y=2.675
+ $X2=2.525 $Y2=2.87
r85 14 28 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.41 $Y=2.59
+ $X2=2.525 $Y2=2.59
r86 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.41 $Y=2.59
+ $X2=1.74 $Y2=2.59
r87 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.61 $Y=2.675
+ $X2=1.74 $Y2=2.59
r88 10 12 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=1.61 $Y=2.675
+ $X2=1.61 $Y2=2.87
r89 3 18 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=2.665 $X2=2.505 $Y2=2.87
r90 2 12 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=2.665 $X2=1.645 $Y2=2.87
r91 1 24 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.745 $X2=2.96 $Y2=0.975
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%Q 1 2 9 13 15 16 17 18
r14 17 18 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.34 $Y=1.295
+ $X2=10.34 $Y2=1.665
r15 16 17 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.34 $Y=0.925
+ $X2=10.34 $Y2=1.295
r16 15 16 16.8598 $w=2.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.34 $Y=0.53
+ $X2=10.34 $Y2=0.925
r17 14 18 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.34 $Y=1.845
+ $X2=10.34 $Y2=1.665
r18 13 14 6.08772 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=10.302 $Y=2.01
+ $X2=10.302 $Y2=1.845
r19 7 13 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=10.302 $Y=2.017
+ $X2=10.302 $Y2=2.01
r20 7 9 29.8299 $w=3.43e-07 $l=8.93e-07 $layer=LI1_cond $X=10.302 $Y=2.017
+ $X2=10.302 $Y2=2.91
r21 2 13 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=10.085
+ $Y=1.835 $X2=10.225 $Y2=2.01
r22 2 9 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.085
+ $Y=1.835 $X2=10.225 $Y2=2.91
r23 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.16
+ $Y=0.385 $X2=10.3 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_1%VGND 1 2 3 4 5 18 22 26 30 35 36 37 39 44 49
+ 61 70 71 74 77 81 87
r108 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r109 81 84 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.17 $Y=0 $X2=5.17
+ $Y2=0.26
r110 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r111 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r112 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r113 71 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r114 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r115 68 87 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=10.035 $Y=0
+ $X2=9.865 $Y2=0
r116 68 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.035 $Y=0
+ $X2=10.32 $Y2=0
r117 67 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r118 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r119 64 67 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.36 $Y2=0
r120 63 66 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.36
+ $Y2=0
r121 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r122 61 87 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.695 $Y=0 $X2=9.865
+ $Y2=0
r123 61 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.695 $Y=0
+ $X2=9.36 $Y2=0
r124 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r125 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r126 57 60 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=7.44 $Y2=0
r127 56 59 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r128 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r129 54 81 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.17
+ $Y2=0
r130 54 56 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.335 $Y=0
+ $X2=5.52 $Y2=0
r131 53 82 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r132 53 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r133 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r134 50 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.17
+ $Y2=0
r135 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.335 $Y=0
+ $X2=2.64 $Y2=0
r136 49 81 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.005 $Y=0 $X2=5.17
+ $Y2=0
r137 49 52 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=5.005 $Y=0
+ $X2=2.64 $Y2=0
r138 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r139 48 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r140 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r141 45 74 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.69
+ $Y2=0
r142 45 47 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=0.785 $Y=0
+ $X2=1.68 $Y2=0
r143 44 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.17
+ $Y2=0
r144 44 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=1.68 $Y2=0
r145 42 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r146 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r147 39 74 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.69
+ $Y2=0
r148 39 41 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.24 $Y2=0
r149 37 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.52 $Y2=0
r150 37 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.04 $Y2=0
r151 35 59 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=7.51 $Y=0 $X2=7.44
+ $Y2=0
r152 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.51 $Y=0 $X2=7.675
+ $Y2=0
r153 34 63 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.84 $Y=0 $X2=7.92
+ $Y2=0
r154 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.84 $Y=0 $X2=7.675
+ $Y2=0
r155 30 32 18.473 $w=3.38e-07 $l=5.45e-07 $layer=LI1_cond $X=9.865 $Y=0.51
+ $X2=9.865 $Y2=1.055
r156 28 87 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=9.865 $Y=0.085
+ $X2=9.865 $Y2=0
r157 28 30 14.4055 $w=3.38e-07 $l=4.25e-07 $layer=LI1_cond $X=9.865 $Y=0.085
+ $X2=9.865 $Y2=0.51
r158 24 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.675 $Y=0.085
+ $X2=7.675 $Y2=0
r159 24 26 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=7.675 $Y=0.085
+ $X2=7.675 $Y2=0.86
r160 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=0.085
+ $X2=2.17 $Y2=0
r161 20 22 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=2.17 $Y=0.085
+ $X2=2.17 $Y2=0.91
r162 16 74 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r163 16 18 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.765
r164 5 32 182 $w=1.7e-07 $l=7.72205e-07 $layer=licon1_NDIFF $count=1 $X=9.65
+ $Y=0.385 $X2=9.87 $Y2=1.055
r165 5 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.65
+ $Y=0.385 $X2=9.86 $Y2=0.51
r166 4 26 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=7.535
+ $Y=0.665 $X2=7.675 $Y2=0.86
r167 3 84 182 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_NDIFF $count=1 $X=4.915
+ $Y=0.535 $X2=5.17 $Y2=0.26
r168 2 22 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.745 $X2=2.17 $Y2=0.91
r169 1 18 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.57 $X2=0.69 $Y2=0.765
.ends

