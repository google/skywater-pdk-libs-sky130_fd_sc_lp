* File: sky130_fd_sc_lp__dlxbp_lp.spice
* Created: Wed Sep  2 09:48:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxbp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dlxbp_lp  VNB VPB D GATE VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1021 A_114_111# N_D_M1021_g N_A_27_111#_M1021_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_D_M1010_g A_114_111# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1011 A_272_111# N_GATE_M1011_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_A_350_111#_M1033_d N_GATE_M1033_g A_272_111# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_556_47# N_A_350_111#_M1007_g N_A_469_47#_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_350_111#_M1008_g A_556_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1009 A_720_47# N_A_27_111#_M1009_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1019 N_A_798_47#_M1019_d N_A_469_47#_M1019_g A_720_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1020 A_900_47# N_A_350_111#_M1020_g N_A_798_47#_M1019_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0756 PD=0.81 PS=0.78 NRD=39.996 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_969_407#_M1001_g A_900_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1064 AS=0.0819 PD=0.876667 PS=0.81 NRD=55.704 NRS=39.996 M=1 R=2.8
+ SA=75002.5 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1031 A_1133_47# N_A_798_47#_M1031_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2128 PD=1.05 PS=1.75333 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1022 N_A_969_407#_M1022_d N_A_798_47#_M1022_g A_1133_47# VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75002
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1034 A_1403_47# N_A_969_407#_M1034_g N_Q_M1034_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2394 PD=1.05 PS=2.25 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A_969_407#_M1002_g A_1403_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1904 AS=0.0882 PD=1.64667 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1035 A_1584_131# N_A_969_407#_M1035_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0952 PD=0.66 PS=0.823333 NRD=18.564 NRS=49.044 M=1 R=2.8
+ SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_A_1662_131#_M1024_d N_A_969_407#_M1024_g A_1584_131# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 A_1860_53# N_A_1662_131#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2394 PD=1.05 PS=2.25 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1030 N_Q_N_M1030_d N_A_1662_131#_M1030_g A_1860_53# VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1032 A_112_481# N_D_M1032_g N_A_27_111#_M1032_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.176 PD=0.85 PS=1.83 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1028 N_VPWR_M1028_d N_D_M1028_g A_112_481# VPB PHIGHVT L=0.15 W=0.64 AD=0.1024
+ AS=0.0672 PD=0.96 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1025 A_278_481# N_GATE_M1025_g N_VPWR_M1028_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1024 PD=0.85 PS=0.96 NRD=15.3857 NRS=12.2928 M=1 R=4.26667
+ SA=75001 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1023 N_A_350_111#_M1023_d N_GATE_M1023_g A_278_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.4904 AS=0.0672 PD=3.78 PS=0.85 NRD=218.926 NRS=15.3857 M=1 R=4.26667
+ SA=75001.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1012 A_567_475# N_A_350_111#_M1012_g N_A_469_47#_M1012_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0672 AS=0.176 PD=0.85 PS=1.83 NRD=15.3857 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1015 N_VPWR_M1015_d N_A_350_111#_M1015_g A_567_475# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1152 AS=0.0672 PD=1 PS=0.85 NRD=24.6053 NRS=15.3857 M=1 R=4.26667
+ SA=75000.6 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1013 A_741_475# N_A_27_111#_M1013_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1152 PD=0.88 PS=1 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1017 N_A_798_47#_M1017_d N_A_350_111#_M1017_g A_741_475# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.136091 AS=0.0768 PD=1.24377 PS=0.88 NRD=0 NRS=19.9955 M=1
+ R=4.26667 SA=75001.5 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1029 A_927_519# N_A_469_47#_M1029_g N_A_798_47#_M1017_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0893094 PD=0.66 PS=0.816226 NRD=30.4759 NRS=51.5943 M=1
+ R=2.8 SA=75002 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_969_407#_M1005_g A_927_519# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.119175 AS=0.0504 PD=0.9225 PS=0.66 NRD=143.042 NRS=30.4759 M=1 R=2.8
+ SA=75002.4 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1026 A_1152_361# N_A_798_47#_M1026_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.357525 PD=1.47 PS=2.7675 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_A_969_407#_M1014_d N_A_798_47#_M1014_g A_1152_361# VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3465 AS=0.1323 PD=3.07 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1018 A_1418_361# N_A_969_407#_M1018_g N_Q_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3465 PD=1.47 PS=3.07 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_A_969_407#_M1016_g A_1418_361# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.276471 AS=0.1323 PD=2.18179 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1000 A_1597_361# N_A_969_407#_M1000_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.140429 PD=0.85 PS=1.10821 NRD=15.3857 NRS=32.308 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1003 N_A_1662_131#_M1003_d N_A_969_407#_M1003_g A_1597_361# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.176 AS=0.0672 PD=1.83 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 A_1863_367# N_A_1662_131#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.3465 PD=1.47 PS=3.07 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_Q_N_M1006_d N_A_1662_131#_M1006_g A_1863_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3402 AS=0.1323 PD=3.06 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX36_noxref VNB VPB NWDIODE A=19.9849 P=25.23
c_182 VPB 0 4.62333e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlxbp_lp.pxi.spice"
*
.ends
*
*
