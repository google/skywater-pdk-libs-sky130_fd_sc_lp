* File: sky130_fd_sc_lp__o22a_1.pxi.spice
* Created: Wed Sep  2 10:19:48 2020
* 
x_PM_SKY130_FD_SC_LP__O22A_1%A_80_21# N_A_80_21#_M1000_d N_A_80_21#_M1009_d
+ N_A_80_21#_c_60_n N_A_80_21#_M1004_g N_A_80_21#_M1006_g N_A_80_21#_c_62_n
+ N_A_80_21#_c_63_n N_A_80_21#_c_64_n N_A_80_21#_c_65_n N_A_80_21#_c_66_n
+ N_A_80_21#_c_76_p N_A_80_21#_c_107_p N_A_80_21#_c_126_p N_A_80_21#_c_89_p
+ N_A_80_21#_c_94_p N_A_80_21#_c_67_n N_A_80_21#_c_68_n
+ PM_SKY130_FD_SC_LP__O22A_1%A_80_21#
x_PM_SKY130_FD_SC_LP__O22A_1%B1 N_B1_M1000_g N_B1_M1008_g B1 N_B1_c_130_n
+ N_B1_c_131_n PM_SKY130_FD_SC_LP__O22A_1%B1
x_PM_SKY130_FD_SC_LP__O22A_1%B2 N_B2_M1009_g N_B2_M1001_g B2 N_B2_c_164_n
+ N_B2_c_167_n PM_SKY130_FD_SC_LP__O22A_1%B2
x_PM_SKY130_FD_SC_LP__O22A_1%A2 N_A2_M1007_g N_A2_M1005_g A2 A2 A2 A2
+ N_A2_c_200_n N_A2_c_201_n PM_SKY130_FD_SC_LP__O22A_1%A2
x_PM_SKY130_FD_SC_LP__O22A_1%A1 N_A1_M1002_g N_A1_M1003_g A1 N_A1_c_238_n
+ N_A1_c_239_n PM_SKY130_FD_SC_LP__O22A_1%A1
x_PM_SKY130_FD_SC_LP__O22A_1%X N_X_M1004_s N_X_M1006_s N_X_c_261_n N_X_c_262_n
+ N_X_c_276_p X X X X X X X X PM_SKY130_FD_SC_LP__O22A_1%X
x_PM_SKY130_FD_SC_LP__O22A_1%VPWR N_VPWR_M1006_d N_VPWR_M1003_d N_VPWR_c_285_n
+ N_VPWR_c_286_n N_VPWR_c_287_n VPWR N_VPWR_c_288_n N_VPWR_c_289_n
+ N_VPWR_c_290_n N_VPWR_c_284_n PM_SKY130_FD_SC_LP__O22A_1%VPWR
x_PM_SKY130_FD_SC_LP__O22A_1%VGND N_VGND_M1004_d N_VGND_M1007_d N_VGND_c_329_n
+ N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n VGND N_VGND_c_333_n
+ N_VGND_c_334_n N_VGND_c_335_n N_VGND_c_336_n PM_SKY130_FD_SC_LP__O22A_1%VGND
x_PM_SKY130_FD_SC_LP__O22A_1%A_265_47# N_A_265_47#_M1000_s N_A_265_47#_M1001_d
+ N_A_265_47#_M1002_d N_A_265_47#_c_377_n N_A_265_47#_c_389_n
+ N_A_265_47#_c_390_n N_A_265_47#_c_374_n N_A_265_47#_c_375_n
+ N_A_265_47#_c_408_n N_A_265_47#_c_376_n PM_SKY130_FD_SC_LP__O22A_1%A_265_47#
cc_1 VNB N_A_80_21#_c_60_n 0.0222867f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_A_80_21#_M1006_g 0.00847289f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.465
cc_3 VNB N_A_80_21#_c_62_n 0.0176846f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.35
cc_4 VNB N_A_80_21#_c_63_n 0.0489518f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.35
cc_5 VNB N_A_80_21#_c_64_n 0.00637824f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.16
cc_6 VNB N_A_80_21#_c_65_n 0.0033009f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.93
cc_7 VNB N_A_80_21#_c_66_n 0.0242844f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.16
cc_8 VNB N_A_80_21#_c_67_n 0.003381f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.16
cc_9 VNB N_A_80_21#_c_68_n 0.00692367f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.16
cc_10 VNB N_B1_M1000_g 0.0291094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_c_130_n 0.0258836f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.465
cc_12 VNB N_B1_c_131_n 0.00176698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B2_M1001_g 0.0270358f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_14 VNB N_B2_c_164_n 0.0286568f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.465
cc_15 VNB N_A2_M1007_g 0.0273486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_200_n 0.0237554f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.93
cc_17 VNB N_A2_c_201_n 0.00446163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1002_g 0.0305946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1003_g 0.00142184f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_20 VNB N_A1_c_238_n 0.0715261f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.35
cc_21 VNB N_A1_c_239_n 0.00129815f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.35
cc_22 VNB X 0.0297138f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.35
cc_23 VNB N_VPWR_c_284_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_329_n 0.00495479f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_25 VNB N_VGND_c_330_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_331_n 0.0504477f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.16
cc_27 VNB N_VGND_c_332_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.16
cc_28 VNB N_VGND_c_333_n 0.0193567f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.16
cc_29 VNB N_VGND_c_334_n 0.0265167f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=2.775
cc_30 VNB N_VGND_c_335_n 0.236974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_336_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.35
cc_32 VNB N_A_265_47#_c_374_n 0.0145233f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.16
cc_33 VNB N_A_265_47#_c_375_n 0.00693609f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.16
cc_34 VNB N_A_265_47#_c_376_n 0.00975526f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.015
cc_35 VPB N_A_80_21#_M1006_g 0.0259574f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.465
cc_36 VPB N_A_80_21#_c_65_n 0.00158832f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.93
cc_37 VPB N_B1_M1008_g 0.0202572f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_38 VPB N_B1_c_130_n 0.00648288f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.465
cc_39 VPB N_B1_c_131_n 0.00306523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_B2_M1009_g 0.0200896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_B2_c_164_n 0.00654814f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.465
cc_42 VPB N_B2_c_167_n 0.00222856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A2_M1005_g 0.0205026f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_44 VPB N_A2_c_200_n 0.00633246f $X=-0.19 $Y=1.655 $X2=1.9 $Y2=0.93
cc_45 VPB N_A2_c_201_n 0.00192701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A1_M1003_g 0.0260229f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_47 VPB N_A1_c_239_n 0.0112502f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.35
cc_48 VPB N_X_c_261_n 0.0153183f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_49 VPB N_X_c_262_n 0.00209686f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_50 VPB X 0.00901783f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.35
cc_51 VPB X 0.00824409f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.93
cc_52 VPB X 0.0462376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_285_n 0.00495479f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_54 VPB N_VPWR_c_286_n 0.0140295f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.465
cc_55 VPB N_VPWR_c_287_n 0.00496839f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_288_n 0.034666f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.93
cc_57 VPB N_VPWR_c_289_n 0.0604661f $X=-0.19 $Y=1.655 $X2=1.9 $Y2=1.075
cc_58 VPB N_VPWR_c_290_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_284_n 0.0658358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 N_A_80_21#_c_63_n N_B1_M1000_g 0.00275425f $X=0.915 $Y=1.35 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_65_n N_B1_M1000_g 0.00180478f $X=1.145 $Y=1.93 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_66_n N_B1_M1000_g 0.0134991f $X=1.795 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_80_21#_M1006_g N_B1_M1008_g 0.0247077f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_65_n N_B1_M1008_g 0.00345409f $X=1.145 $Y=1.93 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_76_p N_B1_M1008_g 0.0158583f $X=2.165 $Y=2.015 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_63_n N_B1_c_130_n 0.0106646f $X=0.915 $Y=1.35 $X2=0 $Y2=0
cc_67 N_A_80_21#_c_65_n N_B1_c_130_n 0.00349497f $X=1.145 $Y=1.93 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_66_n N_B1_c_130_n 0.00442186f $X=1.795 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_76_p N_B1_c_130_n 9.15918e-19 $X=2.165 $Y=2.015 $X2=0 $Y2=0
cc_70 N_A_80_21#_M1006_g N_B1_c_131_n 2.16893e-19 $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_63_n N_B1_c_131_n 2.47205e-19 $X=0.915 $Y=1.35 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_65_n N_B1_c_131_n 0.0238421f $X=1.145 $Y=1.93 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_66_n N_B1_c_131_n 0.0250333f $X=1.795 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_76_p N_B1_c_131_n 0.0226728f $X=2.165 $Y=2.015 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_76_p N_B2_M1009_g 0.0126936f $X=2.165 $Y=2.015 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_66_n N_B2_M1001_g 0.00325867f $X=1.795 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_66_n N_B2_c_164_n 7.57358e-19 $X=1.795 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_89_p N_B2_c_164_n 8.75467e-19 $X=2.27 $Y=2.1 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_66_n N_B2_c_167_n 0.00189267f $X=1.795 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_76_p N_B2_c_167_n 0.0115725f $X=2.165 $Y=2.015 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_89_p N_B2_c_167_n 0.0110643f $X=2.27 $Y=2.1 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_89_p N_A2_M1005_g 7.36419e-19 $X=2.27 $Y=2.1 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_94_p N_A2_M1005_g 0.0045113f $X=2.27 $Y=2.775 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_62_n N_X_c_261_n 0.00794421f $X=0.55 $Y=1.35 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_67_n N_X_c_261_n 0.00492585f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_80_21#_M1006_g N_X_c_262_n 4.72727e-19 $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_63_n N_X_c_262_n 0.0047475f $X=0.915 $Y=1.35 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_65_n N_X_c_262_n 0.00455739f $X=1.145 $Y=1.93 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_67_n N_X_c_262_n 0.00976464f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_60_n X 0.0140789f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_91 N_A_80_21#_M1006_g X 0.00706031f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_67_n X 0.0262166f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_80_21#_M1006_g X 0.00214421f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_65_n N_VPWR_M1006_d 0.00127597f $X=1.145 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A_80_21#_c_76_p N_VPWR_M1006_d 0.0191808f $X=2.165 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_96 N_A_80_21#_c_107_p N_VPWR_M1006_d 0.00165788f $X=1.23 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_80_21#_M1006_g N_VPWR_c_285_n 0.00322989f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_76_p N_VPWR_c_285_n 0.00379027f $X=2.165 $Y=2.015 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_107_p N_VPWR_c_285_n 0.00573525f $X=1.23 $Y=2.015 $X2=0 $Y2=0
cc_100 N_A_80_21#_M1006_g N_VPWR_c_288_n 0.00585385f $X=0.99 $Y=2.465 $X2=0
+ $Y2=0
cc_101 N_A_80_21#_c_94_p N_VPWR_c_289_n 0.00739149f $X=2.27 $Y=2.775 $X2=0 $Y2=0
cc_102 N_A_80_21#_M1009_d N_VPWR_c_284_n 0.0113468f $X=2.13 $Y=1.835 $X2=0 $Y2=0
cc_103 N_A_80_21#_M1006_g N_VPWR_c_284_n 0.0126037f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_94_p N_VPWR_c_284_n 0.00749404f $X=2.27 $Y=2.775 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_76_p A_348_367# 0.0096152f $X=2.165 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_106 N_A_80_21#_c_67_n N_VGND_M1004_d 0.00470837f $X=0.715 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_107 N_A_80_21#_c_60_n N_VGND_c_329_n 0.00460896f $X=0.475 $Y=1.185 $X2=0
+ $Y2=0
cc_108 N_A_80_21#_c_63_n N_VGND_c_329_n 0.00119668f $X=0.915 $Y=1.35 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_67_n N_VGND_c_329_n 0.0156033f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_60_n N_VGND_c_333_n 0.00585385f $X=0.475 $Y=1.185 $X2=0
+ $Y2=0
cc_111 N_A_80_21#_M1000_d N_VGND_c_335_n 0.00250485f $X=1.74 $Y=0.235 $X2=0
+ $Y2=0
cc_112 N_A_80_21#_c_60_n N_VGND_c_335_n 0.0130026f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_113 N_A_80_21#_M1000_d N_A_265_47#_c_377_n 0.00444564f $X=1.74 $Y=0.235 $X2=0
+ $Y2=0
cc_114 N_A_80_21#_c_66_n N_A_265_47#_c_377_n 0.00405582f $X=1.795 $Y=1.16 $X2=0
+ $Y2=0
cc_115 N_A_80_21#_c_126_p N_A_265_47#_c_377_n 0.0101306f $X=1.9 $Y=0.93 $X2=0
+ $Y2=0
cc_116 N_A_80_21#_c_66_n N_A_265_47#_c_375_n 0.00771956f $X=1.795 $Y=1.16 $X2=0
+ $Y2=0
cc_117 N_A_80_21#_c_66_n N_A_265_47#_c_376_n 0.0230731f $X=1.795 $Y=1.16 $X2=0
+ $Y2=0
cc_118 N_B1_M1008_g N_B2_M1009_g 0.0513539f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B1_M1000_g N_B2_M1001_g 0.0375513f $X=1.665 $Y=0.655 $X2=0 $Y2=0
cc_120 N_B1_c_130_n N_B2_c_164_n 0.0513539f $X=1.575 $Y=1.51 $X2=0 $Y2=0
cc_121 N_B1_c_131_n N_B2_c_164_n 0.00195302f $X=1.575 $Y=1.51 $X2=0 $Y2=0
cc_122 N_B1_c_130_n N_B2_c_167_n 3.96249e-19 $X=1.575 $Y=1.51 $X2=0 $Y2=0
cc_123 N_B1_c_131_n N_B2_c_167_n 0.0216763f $X=1.575 $Y=1.51 $X2=0 $Y2=0
cc_124 N_B1_M1008_g N_VPWR_c_285_n 0.0154475f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B1_M1008_g N_VPWR_c_289_n 0.00585385f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B1_M1008_g N_VPWR_c_284_n 0.011444f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B1_M1000_g N_VGND_c_331_n 0.00375954f $X=1.665 $Y=0.655 $X2=0 $Y2=0
cc_128 N_B1_M1000_g N_VGND_c_335_n 0.00695185f $X=1.665 $Y=0.655 $X2=0 $Y2=0
cc_129 N_B1_M1000_g N_A_265_47#_c_377_n 0.00885601f $X=1.665 $Y=0.655 $X2=0
+ $Y2=0
cc_130 N_B1_M1000_g N_A_265_47#_c_376_n 0.00704444f $X=1.665 $Y=0.655 $X2=0
+ $Y2=0
cc_131 N_B2_M1001_g N_A2_M1007_g 0.0251618f $X=2.115 $Y=0.655 $X2=0 $Y2=0
cc_132 N_B2_M1009_g N_A2_M1005_g 0.0255106f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_133 N_B2_c_167_n N_A2_M1005_g 2.99202e-19 $X=2.145 $Y=1.51 $X2=0 $Y2=0
cc_134 N_B2_c_164_n N_A2_c_200_n 0.0165688f $X=2.145 $Y=1.51 $X2=0 $Y2=0
cc_135 N_B2_c_167_n N_A2_c_200_n 3.10661e-19 $X=2.145 $Y=1.51 $X2=0 $Y2=0
cc_136 N_B2_M1009_g N_A2_c_201_n 0.0022298f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_137 N_B2_c_164_n N_A2_c_201_n 0.00172438f $X=2.145 $Y=1.51 $X2=0 $Y2=0
cc_138 N_B2_c_167_n N_A2_c_201_n 0.0210368f $X=2.145 $Y=1.51 $X2=0 $Y2=0
cc_139 N_B2_M1009_g N_VPWR_c_289_n 0.00585385f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_140 N_B2_M1009_g N_VPWR_c_284_n 0.0112998f $X=2.055 $Y=2.465 $X2=0 $Y2=0
cc_141 N_B2_M1001_g N_VGND_c_330_n 0.00132955f $X=2.115 $Y=0.655 $X2=0 $Y2=0
cc_142 N_B2_M1001_g N_VGND_c_331_n 0.00375986f $X=2.115 $Y=0.655 $X2=0 $Y2=0
cc_143 N_B2_M1001_g N_VGND_c_335_n 0.00582967f $X=2.115 $Y=0.655 $X2=0 $Y2=0
cc_144 N_B2_M1001_g N_A_265_47#_c_377_n 0.0128915f $X=2.115 $Y=0.655 $X2=0 $Y2=0
cc_145 N_B2_M1001_g N_A_265_47#_c_375_n 0.00125328f $X=2.115 $Y=0.655 $X2=0
+ $Y2=0
cc_146 N_B2_c_164_n N_A_265_47#_c_375_n 0.00210838f $X=2.145 $Y=1.51 $X2=0 $Y2=0
cc_147 N_B2_c_167_n N_A_265_47#_c_375_n 0.00532403f $X=2.145 $Y=1.51 $X2=0 $Y2=0
cc_148 N_B2_M1001_g N_A_265_47#_c_376_n 7.3356e-19 $X=2.115 $Y=0.655 $X2=0 $Y2=0
cc_149 N_A2_M1007_g N_A1_M1002_g 0.024338f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_150 N_A2_M1005_g N_A1_M1003_g 0.0417717f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A2_c_201_n N_A1_M1003_g 0.0496246f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_152 N_A2_c_200_n N_A1_c_238_n 0.0190171f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_153 N_A2_c_201_n N_A1_c_238_n 0.00723124f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_154 N_A2_c_200_n N_A1_c_239_n 3.29354e-19 $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A2_c_201_n N_A1_c_239_n 0.0250439f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_156 N_A2_c_201_n N_VPWR_c_287_n 0.0571361f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A2_M1005_g N_VPWR_c_289_n 0.00398598f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A2_c_201_n N_VPWR_c_289_n 0.0166396f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A2_M1005_g N_VPWR_c_284_n 0.00640958f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A2_c_201_n N_VPWR_c_284_n 0.0210869f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_161 N_A2_c_201_n A_545_367# 0.0077965f $X=2.74 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_162 N_A2_M1007_g N_VGND_c_330_n 0.0134783f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_163 N_A2_M1007_g N_VGND_c_331_n 0.00486043f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_164 N_A2_M1007_g N_VGND_c_335_n 0.00863238f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_165 N_A2_M1007_g N_A_265_47#_c_389_n 0.00162119f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_166 N_A2_M1007_g N_A_265_47#_c_390_n 0.00678885f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_167 N_A2_M1007_g N_A_265_47#_c_374_n 0.0156881f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A2_c_200_n N_A_265_47#_c_374_n 0.00419993f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A2_c_201_n N_A_265_47#_c_374_n 0.039131f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A1_M1003_g N_VPWR_c_287_n 0.0108971f $X=3.22 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A1_c_238_n N_VPWR_c_287_n 0.00119317f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_172 N_A1_c_239_n N_VPWR_c_287_n 0.0107636f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_173 N_A1_M1003_g N_VPWR_c_289_n 0.00511915f $X=3.22 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A1_M1003_g N_VPWR_c_284_n 0.01015f $X=3.22 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A1_M1002_g N_VGND_c_330_n 0.0117253f $X=3.22 $Y=0.655 $X2=0 $Y2=0
cc_176 N_A1_M1002_g N_VGND_c_334_n 0.00585385f $X=3.22 $Y=0.655 $X2=0 $Y2=0
cc_177 N_A1_M1002_g N_VGND_c_335_n 0.0124556f $X=3.22 $Y=0.655 $X2=0 $Y2=0
cc_178 N_A1_M1002_g N_A_265_47#_c_374_n 0.0185097f $X=3.22 $Y=0.655 $X2=0 $Y2=0
cc_179 N_A1_c_238_n N_A_265_47#_c_374_n 0.00788955f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_180 N_A1_c_239_n N_A_265_47#_c_374_n 0.0116428f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_181 N_X_c_276_p N_VPWR_c_288_n 0.00520647f $X=0.775 $Y=2.66 $X2=0 $Y2=0
cc_182 X N_VPWR_c_288_n 0.00623633f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_183 N_X_M1006_s N_VPWR_c_284_n 0.00452099f $X=0.65 $Y=1.835 $X2=0 $Y2=0
cc_184 N_X_c_276_p N_VPWR_c_284_n 0.00693435f $X=0.775 $Y=2.66 $X2=0 $Y2=0
cc_185 X N_VPWR_c_284_n 0.00710559f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_186 X N_VGND_c_333_n 0.00657075f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_187 N_X_M1004_s N_VGND_c_335_n 0.00433698f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_188 X N_VGND_c_335_n 0.00732528f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_189 N_VPWR_c_284_n A_348_367# 0.010279f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_190 N_VPWR_c_284_n A_545_367# 0.00398889f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_191 N_VGND_c_335_n N_A_265_47#_M1000_s 0.00223961f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_192 N_VGND_c_335_n N_A_265_47#_M1001_d 0.00804887f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_193 N_VGND_c_335_n N_A_265_47#_M1002_d 0.00433698f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_c_331_n N_A_265_47#_c_377_n 0.021557f $X=2.7 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_c_335_n N_A_265_47#_c_377_n 0.0203177f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_c_330_n N_A_265_47#_c_389_n 0.00997958f $X=2.865 $Y=0.38 $X2=0
+ $Y2=0
cc_197 N_VGND_c_331_n N_A_265_47#_c_389_n 0.00884692f $X=2.7 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_335_n N_A_265_47#_c_389_n 0.00777922f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_330_n N_A_265_47#_c_390_n 0.0165095f $X=2.865 $Y=0.38 $X2=0
+ $Y2=0
cc_200 N_VGND_M1007_d N_A_265_47#_c_374_n 0.00516974f $X=2.725 $Y=0.235 $X2=0
+ $Y2=0
cc_201 N_VGND_c_330_n N_A_265_47#_c_374_n 0.0209601f $X=2.865 $Y=0.38 $X2=0
+ $Y2=0
cc_202 N_VGND_c_334_n N_A_265_47#_c_408_n 0.00657075f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_c_335_n N_A_265_47#_c_408_n 0.00732528f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_204 N_VGND_c_329_n N_A_265_47#_c_376_n 0.0204434f $X=0.69 $Y=0.38 $X2=0 $Y2=0
cc_205 N_VGND_c_331_n N_A_265_47#_c_376_n 0.0132397f $X=2.7 $Y=0 $X2=0 $Y2=0
cc_206 N_VGND_c_335_n N_A_265_47#_c_376_n 0.0120072f $X=3.6 $Y=0 $X2=0 $Y2=0
