* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtp_lp D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_566_73# D a_638_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_408_73# a_186_57# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_384_345# a_186_57# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_1208_75# a_887_343# a_1420_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR a_1208_75# a_1949_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND a_1208_75# a_1857_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_862_101# a_186_57# a_887_343# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1949_367# a_1208_75# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND D a_566_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1857_47# a_1208_75# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR a_1208_75# a_996_343# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_1510_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_887_343# a_294_547# a_996_343# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_800_343# a_638_73# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_800_343# a_186_57# a_887_343# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_1208_75# a_887_343# a_1510_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_887_343# a_294_547# a_1058_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_114_470# GATE a_186_57# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_1420_367# a_887_343# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_294_547# a_186_57# a_408_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_1208_75# a_862_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR GATE a_114_470# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 VPWR D a_617_345# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_617_345# D a_638_73# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_114_57# GATE a_186_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND GATE a_114_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_294_547# a_186_57# a_384_345# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_1058_101# a_638_73# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR RESET_B a_1593_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_1593_367# RESET_B a_1208_75# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
