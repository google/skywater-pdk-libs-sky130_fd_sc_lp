* File: sky130_fd_sc_lp__nand4_2.spice
* Created: Wed Sep  2 10:05:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4_2.pex.spice"
.subckt sky130_fd_sc_lp__nand4_2  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1004 N_A_69_47#_M1004_d N_D_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1011 N_A_69_47#_M1011_d N_D_M1011_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1302 AS=0.1176 PD=1.15 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1009 N_A_330_47#_M1009_d N_C_M1009_g N_A_69_47#_M1011_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1302 PD=1.12 PS=1.15 NRD=0 NRS=4.284 M=1 R=5.6
+ SA=75001.1 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1014 N_A_330_47#_M1009_d N_C_M1014_g N_A_69_47#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_523_67#_M1007_d N_B_M1007_g N_A_330_47#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1013 N_A_523_67#_M1013_d N_B_M1013_g N_A_330_47#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1006 N_A_523_67#_M1013_d N_A_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1012 N_A_523_67#_M1012_d N_A_M1012_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.7623 AS=0.1764 PD=3.73 PS=1.54 NRD=17.7103 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_D_M1005_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001 SB=75003.1
+ A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1005_d N_C_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.4
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_C_M1010_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=7.0329 NRS=0 M=1 R=8.4 SA=75001.8
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2268 PD=1.54 PS=1.62 NRD=0 NRS=5.4569 M=1 R=8.4 SA=75002.3
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1015 N_Y_M1003_d N_B_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=1.79 NRD=0 NRS=19.5424 M=1 R=8.4 SA=75002.8
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1015_s N_A_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=1.79 PS=1.54 NRD=19.5424 NRS=0 M=1 R=8.4 SA=75003.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__nand4_2.pxi.spice"
*
.ends
*
*
