* File: sky130_fd_sc_lp__a221o_lp.pex.spice
* Created: Fri Aug 28 09:52:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221O_LP%A_96_183# 1 2 3 12 17 18 19 20 22 25 26 29
+ 32 33 34 37 39 40 42 50 51 52 55 56 59 60
c135 40 0 1.26285e-19 $X=2.785 $Y=0.905
c136 12 0 1.85134e-20 $X=0.685 $Y=2.595
r137 59 60 8.71334 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=4.502 $Y=2.185
+ $X2=4.502 $Y2=2.02
r138 54 56 5.36476 $w=6.78e-07 $l=3.05e-07 $layer=LI1_cond $X=4.32 $Y=0.65
+ $X2=4.625 $Y2=0.65
r139 54 55 10.6764 $w=6.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=0.65
+ $X2=4.155 $Y2=0.65
r140 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.645
+ $Y=1.08 $X2=0.645 $Y2=1.08
r141 47 56 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=4.625 $Y=0.99
+ $X2=4.625 $Y2=0.65
r142 47 60 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=4.625 $Y=0.99
+ $X2=4.625 $Y2=2.02
r143 44 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=0.905
+ $X2=3.095 $Y2=0.905
r144 44 55 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=3.18 $Y=0.905
+ $X2=4.155 $Y2=0.905
r145 41 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.99
+ $X2=3.095 $Y2=0.905
r146 41 42 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.095 $Y=0.99
+ $X2=3.095 $Y2=1.71
r147 39 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=0.905
+ $X2=3.095 $Y2=0.905
r148 39 40 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.01 $Y=0.905
+ $X2=2.785 $Y2=0.905
r149 35 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.62 $Y=0.82
+ $X2=2.785 $Y2=0.905
r150 35 37 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.62 $Y=0.82
+ $X2=2.62 $Y2=0.54
r151 33 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.01 $Y=1.795
+ $X2=3.095 $Y2=1.71
r152 33 34 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=3.01 $Y=1.795
+ $X2=1.75 $Y2=1.795
r153 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.665 $Y=1.71
+ $X2=1.75 $Y2=1.795
r154 31 32 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.665 $Y=1.085
+ $X2=1.665 $Y2=1.71
r155 30 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=1 $X2=0.645
+ $Y2=1
r156 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=1
+ $X2=1.665 $Y2=1.085
r157 29 30 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.58 $Y=1 $X2=0.81
+ $Y2=1
r158 25 51 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.645 $Y=1.42
+ $X2=0.645 $Y2=1.08
r159 25 26 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=1.42
+ $X2=0.645 $Y2=1.585
r160 24 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=0.915
+ $X2=0.645 $Y2=1.08
r161 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.095 $Y=0.255
+ $X2=1.095 $Y2=0.54
r162 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.02 $Y=0.18
+ $X2=1.095 $Y2=0.255
r163 18 19 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.02 $Y=0.18
+ $X2=0.81 $Y2=0.18
r164 17 24 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.735 $Y=0.54
+ $X2=0.735 $Y2=0.915
r165 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.735 $Y=0.255
+ $X2=0.81 $Y2=0.18
r166 14 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.735 $Y=0.255
+ $X2=0.735 $Y2=0.54
r167 12 26 250.938 $w=2.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.685 $Y=2.595
+ $X2=0.685 $Y2=1.585
r168 3 59 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=4.32
+ $Y=2 $X2=4.46 $Y2=2.185
r169 2 54 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.18
+ $Y=0.33 $X2=4.32 $Y2=0.54
r170 1 37 182 $w=1.7e-07 $l=6.46529e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.33 $X2=2.62 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%A2 3 7 9 12 13
c42 13 0 1.85134e-20 $X=1.235 $Y=1.43
c43 12 0 1.11072e-19 $X=1.235 $Y=1.43
r44 12 15 63.4589 $w=6.1e-07 $l=5.05e-07 $layer=POLY_cond $X=1.375 $Y=1.43
+ $X2=1.375 $Y2=1.935
r45 12 14 49.7869 $w=6.1e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.43
+ $X2=1.375 $Y2=1.265
r46 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.235
+ $Y=1.43 $X2=1.235 $Y2=1.43
r47 9 13 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.235 $Y=1.665
+ $X2=1.235 $Y2=1.43
r48 7 14 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=1.605 $Y=0.54
+ $X2=1.605 $Y2=1.265
r49 3 15 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.485 $Y=2.595
+ $X2=1.485 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%A1 3 7 9 10 11 12 17 19
c44 19 0 1.26285e-19 $X=2.09 $Y=0.86
r45 17 19 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.025
+ $X2=2.09 $Y2=0.86
r46 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.095
+ $Y=1.025 $X2=2.095 $Y2=1.025
r47 12 18 9.01912 $w=3.43e-07 $l=2.7e-07 $layer=LI1_cond $X=2.102 $Y=1.295
+ $X2=2.102 $Y2=1.025
r48 11 18 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=2.102 $Y=0.925
+ $X2=2.102 $Y2=1.025
r49 10 11 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.102 $Y=0.555
+ $X2=2.102 $Y2=0.925
r50 8 17 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=2.09 $Y=1.03 $X2=2.09
+ $Y2=1.025
r51 8 9 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=2.09 $Y=1.03 $X2=2.09
+ $Y2=1.36
r52 7 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.995 $Y=0.54
+ $X2=1.995 $Y2=0.86
r53 1 9 47.2392 $w=3.01e-07 $l=3.30379e-07 $layer=POLY_cond $X=2.015 $Y=1.655
+ $X2=2.09 $Y2=1.36
r54 1 3 233.546 $w=2.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.015 $Y=1.655
+ $X2=2.015 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%B1 2 3 4 7 9 11 12 19
r54 17 19 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.665 $Y=1.345
+ $X2=2.835 $Y2=1.345
r55 14 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.575 $Y=1.345
+ $X2=2.665 $Y2=1.345
r56 12 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.345 $X2=2.665 $Y2=1.345
r57 9 11 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.135 $Y=3.075
+ $X2=3.135 $Y2=2.5
r58 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.18
+ $X2=2.835 $Y2=1.345
r59 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.835 $Y=1.18 $X2=2.835
+ $Y2=0.54
r60 3 9 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=3.01 $Y=3.15
+ $X2=3.135 $Y2=3.075
r61 3 4 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.01 $Y=3.15 $X2=2.65
+ $Y2=3.15
r62 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.575 $Y=3.075
+ $X2=2.65 $Y2=3.15
r63 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.51
+ $X2=2.575 $Y2=1.345
r64 1 2 802.479 $w=1.5e-07 $l=1.565e-06 $layer=POLY_cond $X=2.575 $Y=1.51
+ $X2=2.575 $Y2=3.075
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%B2 3 7 9 10 18
c44 9 0 1.64503e-19 $X=3.6 $Y=1.295
r45 16 18 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.55 $Y=1.38
+ $X2=3.665 $Y2=1.38
r46 13 16 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=3.225 $Y=1.38
+ $X2=3.55 $Y2=1.38
r47 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.55 $Y=1.295
+ $X2=3.55 $Y2=1.665
r48 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.38 $X2=3.55 $Y2=1.38
r49 5 18 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.545
+ $X2=3.665 $Y2=1.38
r50 5 7 237.273 $w=2.5e-07 $l=9.55e-07 $layer=POLY_cond $X=3.665 $Y=1.545
+ $X2=3.665 $Y2=2.5
r51 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=1.215
+ $X2=3.225 $Y2=1.38
r52 1 3 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.225 $Y=1.215
+ $X2=3.225 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%C1 1 3 4 5 6 8 11 13 15 17 18 19 20 24
c51 5 0 1.64503e-19 $X=3.82 $Y=0.9
r52 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.195
+ $Y=1.335 $X2=4.195 $Y2=1.335
r53 20 25 9.62801 $w=3.93e-07 $l=3.3e-07 $layer=LI1_cond $X=4.162 $Y=1.665
+ $X2=4.162 $Y2=1.335
r54 19 25 1.16703 $w=3.93e-07 $l=4e-08 $layer=LI1_cond $X=4.162 $Y=1.295
+ $X2=4.162 $Y2=1.335
r55 18 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.195 $Y=1.675
+ $X2=4.195 $Y2=1.335
r56 17 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.195 $Y=1.17
+ $X2=4.195 $Y2=1.335
r57 11 18 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.195 $Y=1.84
+ $X2=4.195 $Y2=1.675
r58 11 13 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.195 $Y=1.84
+ $X2=4.195 $Y2=2.5
r59 9 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.105 $Y=0.975
+ $X2=4.105 $Y2=0.9
r60 9 17 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.105 $Y=0.975
+ $X2=4.105 $Y2=1.17
r61 6 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.105 $Y=0.825
+ $X2=4.105 $Y2=0.9
r62 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.105 $Y=0.825
+ $X2=4.105 $Y2=0.54
r63 4 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.03 $Y=0.9 $X2=4.105
+ $Y2=0.9
r64 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.03 $Y=0.9 $X2=3.82
+ $Y2=0.9
r65 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.745 $Y=0.825
+ $X2=3.82 $Y2=0.9
r66 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.745 $Y=0.825
+ $X2=3.745 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%X 1 2 7 12 13 14 33
c26 12 0 1.11072e-19 $X=0.72 $Y=2.035
r27 24 37 0.589616 $w=7.08e-07 $l=3.5e-08 $layer=LI1_cond $X=0.48 $Y=2.275
+ $X2=0.48 $Y2=2.24
r28 13 14 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.48 $Y=2.405
+ $X2=0.48 $Y2=2.775
r29 13 24 2.19 $w=7.08e-07 $l=1.3e-07 $layer=LI1_cond $X=0.48 $Y=2.405 $X2=0.48
+ $Y2=2.275
r30 12 37 3.45347 $w=7.08e-07 $l=2.05e-07 $layer=LI1_cond $X=0.48 $Y=2.035
+ $X2=0.48 $Y2=2.24
r31 12 33 10.0269 $w=7.08e-07 $l=1.15e-07 $layer=LI1_cond $X=0.48 $Y=2.035
+ $X2=0.48 $Y2=1.92
r32 7 11 11.8188 $w=3.2e-07 $l=4.02654e-07 $layer=LI1_cond $X=0.21 $Y=0.735
+ $X2=0.52 $Y2=0.522
r33 7 33 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=0.21 $Y=0.735
+ $X2=0.21 $Y2=1.92
r34 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.275
+ $Y=2.095 $X2=0.42 $Y2=2.24
r35 1 11 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=0.375
+ $Y=0.33 $X2=0.52 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%VPWR 1 2 9 11 15 17 19 29 30 33 36
r46 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r50 27 30 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 26 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r52 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.28 $Y2=3.33
r54 24 26 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r58 19 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 17 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 17 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=3.33
r62 13 15 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=2.575
r63 12 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r64 11 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.28 $Y2=3.33
r65 11 12 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.345 $Y2=3.33
r66 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245 $X2=1.18
+ $Y2=3.33
r67 7 9 33.7002 $w=3.28e-07 $l=9.65e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.28
r68 2 15 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=2.14
+ $Y=2.095 $X2=2.28 $Y2=2.575
r69 1 9 300 $w=1.7e-07 $l=4.53156e-07 $layer=licon1_PDIFF $count=2 $X=0.81
+ $Y=2.095 $X2=1.18 $Y2=2.28
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%A_322_419# 1 2 9 11 12 13
r35 13 15 5.7303 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=3.4 $Y=2.23 $X2=3.4
+ $Y2=2.385
r36 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.235 $Y=2.145
+ $X2=3.4 $Y2=2.23
r37 11 12 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=3.235 $Y=2.145
+ $X2=1.915 $Y2=2.145
r38 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.75 $Y=2.23
+ $X2=1.915 $Y2=2.145
r39 7 9 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.75 $Y=2.23 $X2=1.75
+ $Y2=2.24
r40 2 15 600 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=3.26 $Y=2
+ $X2=3.4 $Y2=2.385
r41 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.61
+ $Y=2.095 $X2=1.75 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%A_545_400# 1 2 9 11 12 15
r32 13 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.93 $Y=2.895
+ $X2=3.93 $Y2=2.185
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.765 $Y=2.98
+ $X2=3.93 $Y2=2.895
r34 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.765 $Y=2.98
+ $X2=3.035 $Y2=2.98
r35 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.87 $Y=2.895
+ $X2=3.035 $Y2=2.98
r36 7 9 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=2.87 $Y=2.895 $X2=2.87
+ $Y2=2.715
r37 2 15 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=3.79 $Y=2
+ $X2=3.93 $Y2=2.185
r38 1 9 600 $w=1.7e-07 $l=7.84156e-07 $layer=licon1_PDIFF $count=1 $X=2.725 $Y=2
+ $X2=2.87 $Y2=2.715
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_LP%VGND 1 2 9 13 16 17 18 27 36 37 40
r46 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r47 37 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r48 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r49 34 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=0 $X2=3.44
+ $Y2=0
r50 34 36 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.605 $Y=0 $X2=4.56
+ $Y2=0
r51 33 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r52 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r53 29 32 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r54 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 27 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=0 $X2=3.44
+ $Y2=0
r56 27 32 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=0 $X2=3.12
+ $Y2=0
r57 26 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r58 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 22 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r60 21 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r61 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r62 18 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r63 18 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r64 16 25 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.2
+ $Y2=0
r65 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.39
+ $Y2=0
r66 15 29 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=0 $X2=1.68
+ $Y2=0
r67 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=0 $X2=1.39
+ $Y2=0
r68 11 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=0.085
+ $X2=3.44 $Y2=0
r69 11 13 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.44 $Y=0.085
+ $X2=3.44 $Y2=0.475
r70 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.39 $Y=0.085 $X2=1.39
+ $Y2=0
r71 7 9 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.39 $Y=0.085
+ $X2=1.39 $Y2=0.52
r72 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.3
+ $Y=0.33 $X2=3.44 $Y2=0.475
r73 1 9 182 $w=1.7e-07 $l=3.00333e-07 $layer=licon1_NDIFF $count=1 $X=1.17
+ $Y=0.33 $X2=1.39 $Y2=0.52
.ends

