# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a211oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a211oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.835000 1.180000 3.205000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 1.345000 1.645000 1.615000 ;
        RECT 0.120000 1.615000 3.555000 1.785000 ;
        RECT 3.385000 1.270000 3.760000 1.535000 ;
        RECT 3.385000 1.535000 3.555000 1.615000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.980000 1.210000 7.240000 1.255000 ;
        RECT 3.980000 1.255000 5.180000 1.515000 ;
        RECT 4.895000 1.085000 7.240000 1.210000 ;
        RECT 6.980000 1.255000 7.240000 1.515000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.350000 1.425000 6.710000 1.645000 ;
        RECT 5.350000 1.645000 6.145000 1.765000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.116800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.835000 0.755000 7.580000 0.915000 ;
        RECT 1.835000 0.915000 4.725000 1.010000 ;
        RECT 4.055000 0.255000 4.355000 0.725000 ;
        RECT 4.055000 0.725000 5.285000 0.745000 ;
        RECT 4.055000 0.745000 7.580000 0.755000 ;
        RECT 4.955000 0.255000 5.285000 0.725000 ;
        RECT 5.395000 1.935000 7.580000 1.985000 ;
        RECT 5.395000 1.985000 6.615000 2.145000 ;
        RECT 5.815000 0.255000 6.145000 0.745000 ;
        RECT 6.315000 1.815000 7.580000 1.935000 ;
        RECT 6.675000 0.255000 7.005000 0.745000 ;
        RECT 7.410000 0.915000 7.580000 1.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  0.085000 0.415000 1.095000 ;
      RECT 0.185000  1.955000 3.945000 2.125000 ;
      RECT 0.185000  2.125000 0.445000 3.075000 ;
      RECT 0.585000  0.255000 0.805000 1.005000 ;
      RECT 0.585000  1.005000 1.665000 1.175000 ;
      RECT 0.615000  2.295000 0.945000 3.245000 ;
      RECT 0.975000  0.085000 1.305000 0.835000 ;
      RECT 1.115000  2.125000 1.305000 3.075000 ;
      RECT 1.475000  0.255000 3.385000 0.585000 ;
      RECT 1.475000  0.585000 1.665000 1.005000 ;
      RECT 1.475000  2.295000 1.805000 3.245000 ;
      RECT 1.975000  2.125000 2.165000 3.075000 ;
      RECT 2.335000  2.295000 2.665000 3.245000 ;
      RECT 2.835000  2.125000 3.025000 3.075000 ;
      RECT 3.195000  2.295000 3.525000 3.245000 ;
      RECT 3.555000  0.085000 3.885000 0.585000 ;
      RECT 3.695000  2.125000 3.945000 3.075000 ;
      RECT 3.735000  1.705000 4.805000 1.875000 ;
      RECT 3.735000  1.875000 3.945000 1.955000 ;
      RECT 4.165000  2.045000 4.375000 2.745000 ;
      RECT 4.165000  2.745000 6.965000 3.075000 ;
      RECT 4.525000  0.085000 4.785000 0.555000 ;
      RECT 4.595000  1.875000 4.805000 2.325000 ;
      RECT 4.595000  2.325000 7.465000 2.575000 ;
      RECT 5.455000  0.085000 5.645000 0.575000 ;
      RECT 6.315000  0.085000 6.505000 0.575000 ;
      RECT 7.135000  2.165000 7.465000 2.325000 ;
      RECT 7.135000  2.575000 7.465000 3.055000 ;
      RECT 7.175000  0.085000 7.435000 0.575000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__a211oi_4
END LIBRARY
