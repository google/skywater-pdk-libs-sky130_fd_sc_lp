* File: sky130_fd_sc_lp__and2b_4.spice
* Created: Fri Aug 28 10:05:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and2b_4.pex.spice"
.subckt sky130_fd_sc_lp__and2b_4  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_N_M1006_g N_A_43_367#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=28.56 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_213_23#_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1001_d N_A_213_23#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9 SB=75002
+ A=0.126 P=1.98 MULT=1
MM1008 N_X_M1008_d N_A_213_23#_M1008_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.3
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1012 N_X_M1008_d N_A_213_23#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1785 PD=1.12 PS=1.265 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1010 A_616_49# N_B_M1010_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.1785 PD=1.05 PS=1.265 NRD=7.14 NRS=10.704 M=1 R=5.6 SA=75002.3 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1011 N_A_213_23#_M1011_d N_A_43_367#_M1011_g A_616_49# VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75002.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_A_N_M1004_g N_A_43_367#_M1004_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.101325 AS=0.1113 PD=0.8475 PS=1.37 NRD=87.3498 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_213_23#_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.303975 PD=1.54 PS=2.5425 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1002 N_X_M1000_d N_A_213_23#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8 SB=75002
+ A=0.189 P=2.82 MULT=1
MM1005 N_X_M1005_d N_A_213_23#_M1005_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.2
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1013 N_X_M1005_d N_A_213_23#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.22365 PD=1.54 PS=1.615 NRD=0 NRS=5.4569 M=1 R=8.4 SA=75001.7
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1009 N_A_213_23#_M1009_d N_B_M1009_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.22365 PD=1.54 PS=1.615 NRD=0 NRS=6.2449 M=1 R=8.4 SA=75002.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A_43_367#_M1003_g N_A_213_23#_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_39 VNB 0 5.24654e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__and2b_4.pxi.spice"
*
.ends
*
*
