* File: sky130_fd_sc_lp__a2bb2o_4.pex.spice
* Created: Fri Aug 28 09:56:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%B1 3 7 11 15 17 20 23 24 26 27 30 31 43
c82 31 0 5.42069e-20 $X=0.635 $Y=1.95
c83 27 0 1.87504e-19 $X=1.805 $Y=1.51
c84 23 0 1.33101e-19 $X=1.55 $Y=1.95
r85 41 43 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.715 $Y=2.035
+ $X2=0.72 $Y2=2.035
r86 31 41 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=2.035
+ $X2=0.715 $Y2=2.035
r87 31 43 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.76 $Y=2.035 $X2=0.72
+ $Y2=2.035
r88 30 31 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=0.76 $Y2=2.035
r89 29 31 15.247 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.63 $Y=1.645
+ $X2=0.63 $Y2=1.95
r90 27 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.51
+ $X2=1.805 $Y2=1.675
r91 27 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.51
+ $X2=1.805 $Y2=1.345
r92 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.805
+ $Y=1.51 $X2=1.805 $Y2=1.51
r93 24 26 8.16314 $w=2.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.635 $Y=1.525
+ $X2=1.805 $Y2=1.525
r94 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.55 $Y=1.95
+ $X2=1.465 $Y2=2.035
r95 22 24 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.55 $Y=1.645
+ $X2=1.635 $Y2=1.525
r96 22 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.55 $Y=1.645
+ $X2=1.55 $Y2=1.95
r97 20 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.405 $Y=1.51
+ $X2=0.405 $Y2=1.675
r98 20 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.405 $Y=1.51
+ $X2=0.405 $Y2=1.345
r99 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.51 $X2=0.405 $Y2=1.51
r100 17 29 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.545 $Y=1.495
+ $X2=0.63 $Y2=1.645
r101 17 19 5.37807 $w=2.98e-07 $l=1.4e-07 $layer=LI1_cond $X=0.545 $Y=1.495
+ $X2=0.405 $Y2=1.495
r102 15 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.825 $Y=2.465
+ $X2=1.825 $Y2=1.675
r103 11 39 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.785 $Y=0.655
+ $X2=1.785 $Y2=1.345
r104 7 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.495 $Y=2.465
+ $X2=0.495 $Y2=1.675
r105 3 36 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=0.655
+ $X2=0.495 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%B2 3 7 11 15 17 23 24
c50 23 0 1.87504e-19 $X=1.06 $Y=1.51
r51 22 24 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=1.06 $Y=1.51
+ $X2=1.355 $Y2=1.51
r52 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.51 $X2=1.06 $Y2=1.51
r53 19 22 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=1.06 $Y2=1.51
r54 17 23 4.46572 $w=3.98e-07 $l=1.55e-07 $layer=LI1_cond $X=1.095 $Y=1.665
+ $X2=1.095 $Y2=1.51
r55 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.675
+ $X2=1.355 $Y2=1.51
r56 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.355 $Y=1.675
+ $X2=1.355 $Y2=2.465
r57 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.345
+ $X2=1.355 $Y2=1.51
r58 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.355 $Y=1.345
+ $X2=1.355 $Y2=0.655
r59 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.675
+ $X2=0.925 $Y2=1.51
r60 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.925 $Y=1.675
+ $X2=0.925 $Y2=2.465
r61 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=1.51
r62 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%A_436_21# 1 2 3 12 16 18 22 26 28 32 34 35
+ 36 37 40 44 46 50 52 53
r117 48 50 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.69 $Y=0.725
+ $X2=4.69 $Y2=0.42
r118 47 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.835 $Y=0.81
+ $X2=3.705 $Y2=0.81
r119 46 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.525 $Y=0.81
+ $X2=4.69 $Y2=0.725
r120 46 47 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.525 $Y=0.81
+ $X2=3.835 $Y2=0.81
r121 42 53 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.66 $Y=2.035
+ $X2=3.66 $Y2=1.845
r122 42 44 28.2554 $w=2.08e-07 $l=5.35e-07 $layer=LI1_cond $X=3.745 $Y=2.035
+ $X2=4.28 $Y2=2.035
r123 38 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=0.725
+ $X2=3.705 $Y2=0.81
r124 38 40 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=3.705 $Y=0.725
+ $X2=3.705 $Y2=0.42
r125 36 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=1.845
+ $X2=3.66 $Y2=1.845
r126 36 37 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.575 $Y=1.845
+ $X2=2.925 $Y2=1.845
r127 34 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.575 $Y=0.81
+ $X2=3.705 $Y2=0.81
r128 34 35 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.575 $Y=0.81
+ $X2=2.925 $Y2=0.81
r129 33 60 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.807 $Y=1.44
+ $X2=2.807 $Y2=1.605
r130 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.44 $X2=2.84 $Y2=1.44
r131 30 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.84 $Y=1.76
+ $X2=2.925 $Y2=1.845
r132 30 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.84 $Y=1.76
+ $X2=2.84 $Y2=1.44
r133 29 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.84 $Y=0.895
+ $X2=2.925 $Y2=0.81
r134 29 32 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.84 $Y=0.895
+ $X2=2.84 $Y2=1.44
r135 26 60 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.685 $Y=2.465
+ $X2=2.685 $Y2=1.605
r136 22 58 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.685 $Y=0.655
+ $X2=2.685 $Y2=1.275
r137 19 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.33 $Y=1.35
+ $X2=2.255 $Y2=1.35
r138 18 33 12.6719 $w=3.95e-07 $l=9e-08 $layer=POLY_cond $X=2.807 $Y=1.35
+ $X2=2.807 $Y2=1.44
r139 18 58 32.8921 $w=3.95e-07 $l=7.5e-08 $layer=POLY_cond $X=2.807 $Y=1.35
+ $X2=2.807 $Y2=1.275
r140 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.61 $Y=1.35
+ $X2=2.33 $Y2=1.35
r141 14 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.255 $Y=1.425
+ $X2=2.255 $Y2=1.35
r142 14 16 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.255 $Y=1.425
+ $X2=2.255 $Y2=2.465
r143 10 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.255 $Y=1.275
+ $X2=2.255 $Y2=1.35
r144 10 12 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.255 $Y=1.275
+ $X2=2.255 $Y2=0.655
r145 3 44 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=4.14
+ $Y=1.835 $X2=4.28 $Y2=2.035
r146 2 50 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.55
+ $Y=0.235 $X2=4.69 $Y2=0.42
r147 1 40 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.53
+ $Y=0.235 $X2=3.67 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%A1_N 1 3 4 6 9 12 14 21 26 27 28
c82 27 0 2.17925e-19 $X=4.945 $Y=1.35
c83 26 0 5.38188e-20 $X=4.945 $Y=1.35
c84 14 0 9.12621e-20 $X=3.41 $Y=1.15
r85 26 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.945 $Y=1.35
+ $X2=4.945 $Y2=1.515
r86 26 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.945 $Y=1.35
+ $X2=4.945 $Y2=1.185
r87 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.945
+ $Y=1.35 $X2=4.945 $Y2=1.35
r88 21 27 10.2331 $w=4.48e-07 $l=3.85e-07 $layer=LI1_cond $X=4.56 $Y=1.29
+ $X2=4.945 $Y2=1.29
r89 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.41
+ $Y=1.35 $X2=3.41 $Y2=1.35
r90 15 21 51.4005 $w=1.93e-07 $l=9e-07 $layer=LI1_cond $X=3.575 $Y=1.15
+ $X2=4.475 $Y2=1.15
r91 14 18 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.41 $Y=1.15 $X2=3.41
+ $Y2=1.35
r92 14 15 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=1.15
+ $X2=3.575 $Y2=1.15
r93 12 29 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.925 $Y=2.465
+ $X2=4.925 $Y2=1.515
r94 9 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.905 $Y=0.655
+ $X2=4.905 $Y2=1.185
r95 4 19 72.647 $w=2.97e-07 $l=4.47074e-07 $layer=POLY_cond $X=3.635 $Y=1.725
+ $X2=3.477 $Y2=1.35
r96 4 6 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.635 $Y=1.725
+ $X2=3.635 $Y2=2.465
r97 1 19 38.5662 $w=2.97e-07 $l=1.75656e-07 $layer=POLY_cond $X=3.455 $Y=1.185
+ $X2=3.477 $Y2=1.35
r98 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.455 $Y=1.185
+ $X2=3.455 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%A2_N 1 3 6 8 10 13 15 21 22
c53 21 0 5.38188e-20 $X=4.13 $Y=1.5
c54 1 0 9.12621e-20 $X=3.89 $Y=1.185
r55 22 23 2.38025 $w=4.05e-07 $l=2e-08 $layer=POLY_cond $X=4.475 $Y=1.425
+ $X2=4.495 $Y2=1.425
r56 20 22 41.0593 $w=4.05e-07 $l=3.45e-07 $layer=POLY_cond $X=4.13 $Y=1.425
+ $X2=4.475 $Y2=1.425
r57 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.13
+ $Y=1.5 $X2=4.13 $Y2=1.5
r58 18 20 7.7358 $w=4.05e-07 $l=6.5e-08 $layer=POLY_cond $X=4.065 $Y=1.425
+ $X2=4.13 $Y2=1.425
r59 15 21 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.13 $Y=1.665
+ $X2=4.13 $Y2=1.5
r60 11 23 26.1659 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.495 $Y=1.665
+ $X2=4.495 $Y2=1.425
r61 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.495 $Y=1.665
+ $X2=4.495 $Y2=2.465
r62 8 22 26.1659 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.475 $Y=1.185
+ $X2=4.475 $Y2=1.425
r63 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.475 $Y=1.185
+ $X2=4.475 $Y2=0.655
r64 4 18 26.1659 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.065 $Y=1.665
+ $X2=4.065 $Y2=1.425
r65 4 6 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.065 $Y=1.665 $X2=4.065
+ $Y2=2.465
r66 1 18 20.8272 $w=4.05e-07 $l=3.15595e-07 $layer=POLY_cond $X=3.89 $Y=1.185
+ $X2=4.065 $Y2=1.425
r67 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.89 $Y=1.185 $X2=3.89
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%A_200_47# 1 2 3 12 16 20 24 28 32 36 40 44
+ 46 47 51 54 58 60 62 65 66 71 74 76 88
c157 88 0 9.57946e-20 $X=6.685 $Y=1.49
r158 88 89 5.17485 $w=3.26e-07 $l=3.5e-08 $layer=POLY_cond $X=6.685 $Y=1.49
+ $X2=6.72 $Y2=1.49
r159 85 86 5.17485 $w=3.26e-07 $l=3.5e-08 $layer=POLY_cond $X=6.255 $Y=1.49
+ $X2=6.29 $Y2=1.49
r160 84 85 58.4018 $w=3.26e-07 $l=3.95e-07 $layer=POLY_cond $X=5.86 $Y=1.49
+ $X2=6.255 $Y2=1.49
r161 83 84 5.17485 $w=3.26e-07 $l=3.5e-08 $layer=POLY_cond $X=5.825 $Y=1.49
+ $X2=5.86 $Y2=1.49
r162 80 81 3.69632 $w=3.26e-07 $l=2.5e-08 $layer=POLY_cond $X=5.395 $Y=1.49
+ $X2=5.42 $Y2=1.49
r163 76 78 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.32 $Y=2.185
+ $X2=3.32 $Y2=2.395
r164 72 88 22.9172 $w=3.26e-07 $l=1.55e-07 $layer=POLY_cond $X=6.53 $Y=1.49
+ $X2=6.685 $Y2=1.49
r165 72 86 35.4847 $w=3.26e-07 $l=2.4e-07 $layer=POLY_cond $X=6.53 $Y=1.49
+ $X2=6.29 $Y2=1.49
r166 71 72 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.53
+ $Y=1.49 $X2=6.53 $Y2=1.49
r167 69 83 46.5736 $w=3.26e-07 $l=3.15e-07 $layer=POLY_cond $X=5.51 $Y=1.49
+ $X2=5.825 $Y2=1.49
r168 69 81 13.3067 $w=3.26e-07 $l=9e-08 $layer=POLY_cond $X=5.51 $Y=1.49
+ $X2=5.42 $Y2=1.49
r169 68 71 62.8485 $w=1.78e-07 $l=1.02e-06 $layer=LI1_cond $X=5.51 $Y=1.495
+ $X2=6.53 $Y2=1.495
r170 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.51
+ $Y=1.49 $X2=5.51 $Y2=1.49
r171 66 68 8.0101 $w=1.78e-07 $l=1.3e-07 $layer=LI1_cond $X=5.38 $Y=1.495
+ $X2=5.51 $Y2=1.495
r172 64 66 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.295 $Y=1.585
+ $X2=5.38 $Y2=1.495
r173 64 65 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=5.295 $Y=1.585
+ $X2=5.295 $Y2=2.31
r174 63 78 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=2.395
+ $X2=3.32 $Y2=2.395
r175 62 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.21 $Y=2.395
+ $X2=5.295 $Y2=2.31
r176 62 63 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=5.21 $Y=2.395
+ $X2=3.405 $Y2=2.395
r177 61 75 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.565 $Y=2.185
+ $X2=2.455 $Y2=2.185
r178 60 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=2.185
+ $X2=3.32 $Y2=2.185
r179 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.235 $Y=2.185
+ $X2=2.565 $Y2=2.185
r180 56 74 4.3182 $w=2.1e-07 $l=8.9861e-08 $layer=LI1_cond $X=2.465 $Y=1.065
+ $X2=2.455 $Y2=1.15
r181 56 58 35.7682 $w=1.98e-07 $l=6.45e-07 $layer=LI1_cond $X=2.465 $Y=1.065
+ $X2=2.465 $Y2=0.42
r182 52 75 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=2.27
+ $X2=2.455 $Y2=2.185
r183 52 54 15.7151 $w=2.18e-07 $l=3e-07 $layer=LI1_cond $X=2.455 $Y=2.27
+ $X2=2.455 $Y2=2.57
r184 49 75 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=2.1
+ $X2=2.455 $Y2=2.185
r185 49 51 6.28605 $w=2.18e-07 $l=1.2e-07 $layer=LI1_cond $X=2.455 $Y=2.1
+ $X2=2.455 $Y2=1.98
r186 48 74 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=1.235
+ $X2=2.455 $Y2=1.15
r187 48 51 39.0259 $w=2.18e-07 $l=7.45e-07 $layer=LI1_cond $X=2.455 $Y=1.235
+ $X2=2.455 $Y2=1.98
r188 46 74 2.11342 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.345 $Y=1.15
+ $X2=2.455 $Y2=1.15
r189 46 47 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=2.345 $Y=1.15
+ $X2=1.235 $Y2=1.15
r190 42 47 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=1.127 $Y=1.065
+ $X2=1.235 $Y2=1.15
r191 42 44 16.3486 $w=2.13e-07 $l=3.05e-07 $layer=LI1_cond $X=1.127 $Y=1.065
+ $X2=1.127 $Y2=0.76
r192 38 89 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.72 $Y=1.655
+ $X2=6.72 $Y2=1.49
r193 38 40 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.72 $Y=1.655
+ $X2=6.72 $Y2=2.465
r194 34 88 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.685 $Y=1.325
+ $X2=6.685 $Y2=1.49
r195 34 36 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.685 $Y=1.325
+ $X2=6.685 $Y2=0.655
r196 30 86 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.29 $Y=1.655
+ $X2=6.29 $Y2=1.49
r197 30 32 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.29 $Y=1.655
+ $X2=6.29 $Y2=2.465
r198 26 85 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.255 $Y=1.325
+ $X2=6.255 $Y2=1.49
r199 26 28 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.255 $Y=1.325
+ $X2=6.255 $Y2=0.655
r200 22 84 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.86 $Y=1.655
+ $X2=5.86 $Y2=1.49
r201 22 24 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.86 $Y=1.655
+ $X2=5.86 $Y2=2.465
r202 18 83 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=1.325
+ $X2=5.825 $Y2=1.49
r203 18 20 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.825 $Y=1.325
+ $X2=5.825 $Y2=0.655
r204 14 81 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.42 $Y=1.655
+ $X2=5.42 $Y2=1.49
r205 14 16 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.42 $Y=1.655
+ $X2=5.42 $Y2=2.465
r206 10 80 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.325
+ $X2=5.395 $Y2=1.49
r207 10 12 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.395 $Y=1.325
+ $X2=5.395 $Y2=0.655
r208 3 54 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=1.835 $X2=2.47 $Y2=2.57
r209 3 51 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=1.835 $X2=2.47 $Y2=1.98
r210 2 58 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.33
+ $Y=0.235 $X2=2.47 $Y2=0.42
r211 1 44 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.14 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%A_27_367# 1 2 3 4 15 19 23 25 29 33 34 37
+ 40 41
r60 35 37 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.9 $Y=2.905 $X2=2.9
+ $Y2=2.535
r61 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.735 $Y=2.99
+ $X2=2.9 $Y2=2.905
r62 33 34 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.735 $Y=2.99
+ $X2=2.175 $Y2=2.99
r63 32 34 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.055 $Y=2.905
+ $X2=2.175 $Y2=2.99
r64 31 43 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.46
+ $X2=2.055 $Y2=2.375
r65 31 32 21.3682 $w=2.38e-07 $l=4.45e-07 $layer=LI1_cond $X=2.055 $Y=2.46
+ $X2=2.055 $Y2=2.905
r66 27 43 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.29
+ $X2=2.055 $Y2=2.375
r67 27 29 14.8857 $w=2.38e-07 $l=3.1e-07 $layer=LI1_cond $X=2.055 $Y=2.29
+ $X2=2.055 $Y2=1.98
r68 26 41 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.255 $Y=2.375
+ $X2=1.15 $Y2=2.375
r69 25 43 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.935 $Y=2.375
+ $X2=2.055 $Y2=2.375
r70 25 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.935 $Y=2.375
+ $X2=1.255 $Y2=2.375
r71 21 41 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=2.46
+ $X2=1.15 $Y2=2.375
r72 21 23 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=2.46 $X2=1.15
+ $Y2=2.465
r73 20 40 3.18746 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.375 $Y=2.375
+ $X2=0.235 $Y2=2.375
r74 19 41 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.045 $Y=2.375
+ $X2=1.15 $Y2=2.375
r75 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.045 $Y=2.375
+ $X2=0.375 $Y2=2.375
r76 13 40 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=2.29 $X2=0.235
+ $Y2=2.375
r77 13 15 12.7592 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=0.235 $Y=2.29
+ $X2=0.235 $Y2=1.98
r78 4 37 300 $w=1.7e-07 $l=7.66812e-07 $layer=licon1_PDIFF $count=2 $X=2.76
+ $Y=1.835 $X2=2.9 $Y2=2.535
r79 3 43 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=1.9
+ $Y=1.835 $X2=2.04 $Y2=2.45
r80 3 29 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.835 $X2=2.04 $Y2=1.98
r81 2 23 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2.465
r82 1 40 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.45
r83 1 15 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 43 48 49
+ 50 52 57 66 70 75 81 84 87 90 94
r114 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r116 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r118 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r119 79 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r120 79 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r121 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 76 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.24 $Y=3.33
+ $X2=6.075 $Y2=3.33
r123 76 78 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r124 75 93 4.48816 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.8 $Y=3.33 $X2=7
+ $Y2=3.33
r125 75 78 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.8 $Y=3.33 $X2=6.48
+ $Y2=3.33
r126 74 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r127 74 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r128 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r129 71 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=3.33
+ $X2=5.185 $Y2=3.33
r130 71 73 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.35 $Y=3.33
+ $X2=5.52 $Y2=3.33
r131 70 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.91 $Y=3.33
+ $X2=6.075 $Y2=3.33
r132 70 73 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.91 $Y=3.33
+ $X2=5.52 $Y2=3.33
r133 66 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=5.185 $Y2=3.33
r134 66 68 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=3.6 $Y2=3.33
r135 65 85 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=1.68 $Y2=3.33
r136 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r137 62 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=1.59 $Y2=3.33
r138 62 64 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=3.12 $Y2=3.33
r139 61 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r140 61 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r141 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r142 58 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.71 $Y2=3.33
r143 58 60 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=1.2 $Y2=3.33
r144 57 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.59 $Y2=3.33
r145 57 60 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r146 55 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r148 52 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.71 $Y2=3.33
r149 52 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.24 $Y2=3.33
r150 50 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r151 50 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r152 50 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r153 48 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=3.33
+ $X2=3.12 $Y2=3.33
r154 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=3.33
+ $X2=3.42 $Y2=3.33
r155 47 68 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=3.6 $Y2=3.33
r156 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=3.42 $Y2=3.33
r157 43 46 26.5062 $w=2.98e-07 $l=6.9e-07 $layer=LI1_cond $X=6.95 $Y=2.26
+ $X2=6.95 $Y2=2.95
r158 41 93 3.02951 $w=3e-07 $l=1.07121e-07 $layer=LI1_cond $X=6.95 $Y=3.245
+ $X2=7 $Y2=3.33
r159 41 46 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=6.95 $Y=3.245
+ $X2=6.95 $Y2=2.95
r160 37 40 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=6.075 $Y=2.26
+ $X2=6.075 $Y2=2.95
r161 35 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=3.245
+ $X2=6.075 $Y2=3.33
r162 35 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.075 $Y=3.245
+ $X2=6.075 $Y2=2.95
r163 31 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.185 $Y=3.245
+ $X2=5.185 $Y2=3.33
r164 31 33 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=5.185 $Y=3.245
+ $X2=5.185 $Y2=2.775
r165 27 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=3.245
+ $X2=3.42 $Y2=3.33
r166 27 29 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=3.42 $Y=3.245
+ $X2=3.42 $Y2=2.775
r167 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.59 $Y2=3.33
r168 23 25 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.59 $Y2=2.755
r169 19 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=3.245
+ $X2=0.71 $Y2=3.33
r170 19 21 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.71 $Y=3.245
+ $X2=0.71 $Y2=2.755
r171 6 46 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.835 $X2=6.935 $Y2=2.95
r172 6 43 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.835 $X2=6.935 $Y2=2.26
r173 5 40 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.935
+ $Y=1.835 $X2=6.075 $Y2=2.95
r174 5 37 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=5.935
+ $Y=1.835 $X2=6.075 $Y2=2.26
r175 4 33 600 $w=1.7e-07 $l=1.02835e-06 $layer=licon1_PDIFF $count=1 $X=5
+ $Y=1.835 $X2=5.185 $Y2=2.775
r176 3 29 600 $w=1.7e-07 $l=1.00055e-06 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.835 $X2=3.42 $Y2=2.775
r177 2 25 600 $w=1.7e-07 $l=9.96795e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.59 $Y2=2.755
r178 1 21 600 $w=1.7e-07 $l=9.87522e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%A_742_367# 1 2 11
r11 8 11 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=3.85 $Y=2.835
+ $X2=4.71 $Y2=2.835
r12 2 11 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=4.57
+ $Y=1.835 $X2=4.71 $Y2=2.835
r13 1 8 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.835 $X2=3.85 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 40 41
+ 43 44 49 51
r61 49 51 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=6.96 $Y=1.235 $X2=6.96
+ $Y2=1.295
r62 43 49 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.96 $Y=1.15 $X2=6.96
+ $Y2=1.235
r63 43 44 23.3561 $w=1.68e-07 $l=3.58e-07 $layer=LI1_cond $X=6.96 $Y=1.307
+ $X2=6.96 $Y2=1.665
r64 43 51 0.782888 $w=1.68e-07 $l=1.2e-08 $layer=LI1_cond $X=6.96 $Y=1.307
+ $X2=6.96 $Y2=1.295
r65 42 44 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.96 $Y=1.755 $X2=6.96
+ $Y2=1.665
r66 39 43 17.8434 $w=1.93e-07 $l=3.1e-07 $layer=LI1_cond $X=6.565 $Y=1.15
+ $X2=6.875 $Y2=1.15
r67 39 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.565 $Y=1.15
+ $X2=6.47 $Y2=1.15
r68 38 41 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.63 $Y=1.84 $X2=6.52
+ $Y2=1.84
r69 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.875 $Y=1.84
+ $X2=6.96 $Y2=1.755
r70 37 38 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.875 $Y=1.84
+ $X2=6.63 $Y2=1.84
r71 33 35 49.7646 $w=2.18e-07 $l=9.5e-07 $layer=LI1_cond $X=6.52 $Y=1.96
+ $X2=6.52 $Y2=2.91
r72 31 41 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.925
+ $X2=6.52 $Y2=1.84
r73 31 33 1.83343 $w=2.18e-07 $l=3.5e-08 $layer=LI1_cond $X=6.52 $Y=1.925
+ $X2=6.52 $Y2=1.96
r74 27 40 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=1.065
+ $X2=6.47 $Y2=1.15
r75 27 29 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=6.47 $Y=1.065
+ $X2=6.47 $Y2=0.42
r76 25 41 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.41 $Y=1.84 $X2=6.52
+ $Y2=1.84
r77 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.41 $Y=1.84
+ $X2=5.74 $Y2=1.84
r78 23 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.375 $Y=1.15
+ $X2=6.47 $Y2=1.15
r79 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.375 $Y=1.15
+ $X2=5.705 $Y2=1.15
r80 19 21 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=5.645 $Y=1.96
+ $X2=5.645 $Y2=2.91
r81 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.645 $Y=1.925
+ $X2=5.74 $Y2=1.84
r82 17 19 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=5.645 $Y=1.925
+ $X2=5.645 $Y2=1.96
r83 13 24 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.59 $Y=1.065
+ $X2=5.705 $Y2=1.15
r84 13 15 32.3185 $w=2.28e-07 $l=6.45e-07 $layer=LI1_cond $X=5.59 $Y=1.065
+ $X2=5.59 $Y2=0.42
r85 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.365
+ $Y=1.835 $X2=6.505 $Y2=2.91
r86 4 33 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=6.365
+ $Y=1.835 $X2=6.505 $Y2=1.96
r87 3 21 400 $w=1.7e-07 $l=1.14755e-06 $layer=licon1_PDIFF $count=1 $X=5.495
+ $Y=1.835 $X2=5.645 $Y2=2.91
r88 3 19 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=5.495
+ $Y=1.835 $X2=5.645 $Y2=1.96
r89 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.33
+ $Y=0.235 $X2=6.47 $Y2=0.42
r90 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.47
+ $Y=0.235 $X2=5.61 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%VGND 1 2 3 4 5 6 7 22 24 28 30 34 36 40 44
+ 46 48 51 52 53 66 71 82 85 87 90 93 97
c119 5 0 1.22131e-19 $X=4.98 $Y=0.235
r120 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r121 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r122 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r123 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r124 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r125 84 85 10.4169 $w=6.38e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0.235
+ $X2=3.405 $Y2=0.235
r126 80 84 2.24265 $w=6.38e-07 $l=1.2e-07 $layer=LI1_cond $X=3.12 $Y=0.235
+ $X2=3.24 $Y2=0.235
r127 80 82 14.5284 $w=6.38e-07 $l=3.85e-07 $layer=LI1_cond $X=3.12 $Y=0.235
+ $X2=2.735 $Y2=0.235
r128 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r129 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r130 75 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r131 75 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r132 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r133 72 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6.04
+ $Y2=0
r134 72 74 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.205 $Y=0
+ $X2=6.48 $Y2=0
r135 71 96 4.69206 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=6.735 $Y=0
+ $X2=6.967 $Y2=0
r136 71 74 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.735 $Y=0
+ $X2=6.48 $Y2=0
r137 70 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r138 70 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r139 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r140 67 90 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.305 $Y=0 $X2=5.165
+ $Y2=0
r141 67 69 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.305 $Y=0
+ $X2=5.52 $Y2=0
r142 66 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=0 $X2=6.04
+ $Y2=0
r143 66 69 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.875 $Y=0
+ $X2=5.52 $Y2=0
r144 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r145 64 82 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.735
+ $Y2=0
r146 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r147 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r148 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r149 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r150 58 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r151 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r152 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r153 55 77 4.32671 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.2 $Y2=0
r154 55 57 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.72
+ $Y2=0
r155 53 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r156 53 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r157 51 60 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.905 $Y=0
+ $X2=1.68 $Y2=0
r158 51 52 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=2.045
+ $Y2=0
r159 50 64 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=2.64 $Y2=0
r160 50 52 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.045
+ $Y2=0
r161 46 96 3.07411 $w=3.3e-07 $l=1.13666e-07 $layer=LI1_cond $X=6.9 $Y=0.085
+ $X2=6.967 $Y2=0
r162 46 48 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.9 $Y=0.085
+ $X2=6.9 $Y2=0.36
r163 42 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.04 $Y=0.085
+ $X2=6.04 $Y2=0
r164 42 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.04 $Y=0.085
+ $X2=6.04 $Y2=0.36
r165 38 90 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.085
+ $X2=5.165 $Y2=0
r166 38 40 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=5.165 $Y=0.085
+ $X2=5.165 $Y2=0.38
r167 37 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=0 $X2=4.18
+ $Y2=0
r168 36 90 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.025 $Y=0 $X2=5.165
+ $Y2=0
r169 36 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.025 $Y=0
+ $X2=4.345 $Y2=0
r170 32 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=0.085
+ $X2=4.18 $Y2=0
r171 32 34 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.18 $Y=0.085
+ $X2=4.18 $Y2=0.39
r172 30 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.18
+ $Y2=0
r173 30 85 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.015 $Y=0
+ $X2=3.405 $Y2=0
r174 26 52 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0
r175 26 28 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0.38
r176 22 77 3.07196 $w=2.85e-07 $l=1.09864e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.2 $Y2=0
r177 22 24 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r178 7 48 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.76
+ $Y=0.235 $X2=6.9 $Y2=0.36
r179 6 44 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.9
+ $Y=0.235 $X2=6.04 $Y2=0.36
r180 5 40 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=4.98
+ $Y=0.235 $X2=5.14 $Y2=0.38
r181 4 34 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=3.965
+ $Y=0.235 $X2=4.18 $Y2=0.39
r182 3 84 91 $w=1.7e-07 $l=5.71314e-07 $layer=licon1_NDIFF $count=2 $X=2.76
+ $Y=0.235 $X2=3.24 $Y2=0.435
r183 2 28 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.86
+ $Y=0.235 $X2=2.02 $Y2=0.38
r184 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.235 $X2=0.28 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_4%A_114_47# 1 2 9 14 16
r24 10 14 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.85 $Y=0.34 $X2=0.71
+ $Y2=0.34
r25 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0.34
+ $X2=1.57 $Y2=0.34
r26 9 10 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.405 $Y=0.34
+ $X2=0.85 $Y2=0.34
r27 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.38
r28 1 14 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.42
.ends

