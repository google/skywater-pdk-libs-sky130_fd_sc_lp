* File: sky130_fd_sc_lp__einvn_2.pxi.spice
* Created: Wed Sep  2 09:51:39 2020
* 
x_PM_SKY130_FD_SC_LP__EINVN_2%TE_B N_TE_B_M1002_g N_TE_B_c_61_n N_TE_B_c_67_n
+ N_TE_B_M1006_g N_TE_B_c_68_n N_TE_B_M1007_g N_TE_B_c_62_n N_TE_B_c_63_n
+ N_TE_B_c_71_n N_TE_B_M1009_g TE_B TE_B N_TE_B_c_65_n N_TE_B_c_66_n
+ PM_SKY130_FD_SC_LP__EINVN_2%TE_B
x_PM_SKY130_FD_SC_LP__EINVN_2%A_28_62# N_A_28_62#_M1002_s N_A_28_62#_M1006_s
+ N_A_28_62#_c_119_n N_A_28_62#_M1004_g N_A_28_62#_c_120_n N_A_28_62#_M1005_g
+ N_A_28_62#_c_121_n N_A_28_62#_c_126_n N_A_28_62#_c_127_n N_A_28_62#_c_122_n
+ N_A_28_62#_c_129_n N_A_28_62#_c_123_n N_A_28_62#_c_124_n
+ PM_SKY130_FD_SC_LP__EINVN_2%A_28_62#
x_PM_SKY130_FD_SC_LP__EINVN_2%A N_A_M1001_g N_A_M1000_g N_A_c_183_n N_A_M1003_g
+ N_A_M1008_g N_A_c_185_n A N_A_c_187_n N_A_c_188_n
+ PM_SKY130_FD_SC_LP__EINVN_2%A
x_PM_SKY130_FD_SC_LP__EINVN_2%VPWR N_VPWR_M1006_d N_VPWR_M1009_d N_VPWR_c_229_n
+ N_VPWR_c_230_n VPWR N_VPWR_c_231_n N_VPWR_c_232_n N_VPWR_c_233_n
+ N_VPWR_c_228_n N_VPWR_c_235_n N_VPWR_c_236_n PM_SKY130_FD_SC_LP__EINVN_2%VPWR
x_PM_SKY130_FD_SC_LP__EINVN_2%A_220_367# N_A_220_367#_M1007_s
+ N_A_220_367#_M1000_d N_A_220_367#_c_285_n N_A_220_367#_c_273_n
+ N_A_220_367#_c_281_n N_A_220_367#_c_298_p N_A_220_367#_c_275_n
+ N_A_220_367#_c_282_n PM_SKY130_FD_SC_LP__EINVN_2%A_220_367#
x_PM_SKY130_FD_SC_LP__EINVN_2%Z N_Z_M1001_d N_Z_M1000_s N_Z_M1008_s N_Z_c_301_n
+ N_Z_c_302_n N_Z_c_303_n N_Z_c_304_n Z Z Z Z Z N_Z_c_327_n
+ PM_SKY130_FD_SC_LP__EINVN_2%Z
x_PM_SKY130_FD_SC_LP__EINVN_2%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_c_344_n
+ N_VGND_c_345_n N_VGND_c_346_n VGND N_VGND_c_347_n N_VGND_c_348_n
+ N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n PM_SKY130_FD_SC_LP__EINVN_2%VGND
x_PM_SKY130_FD_SC_LP__EINVN_2%A_251_47# N_A_251_47#_M1004_s N_A_251_47#_M1005_s
+ N_A_251_47#_M1003_s N_A_251_47#_c_387_n N_A_251_47#_c_388_n
+ N_A_251_47#_c_389_n N_A_251_47#_c_421_n N_A_251_47#_c_405_n
+ N_A_251_47#_c_390_n PM_SKY130_FD_SC_LP__EINVN_2%A_251_47#
cc_1 VNB N_TE_B_c_61_n 0.0501725f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.575
cc_2 VNB N_TE_B_c_62_n 0.0208478f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.65
cc_3 VNB N_TE_B_c_63_n 0.0197324f $X=-0.19 $Y=-0.245 $X2=1.1 $Y2=1.65
cc_4 VNB TE_B 0.0174589f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_5 VNB N_TE_B_c_65_n 0.0227251f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.005
cc_6 VNB N_TE_B_c_66_n 0.0233818f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=0.84
cc_7 VNB N_A_28_62#_c_119_n 0.0189804f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.155
cc_8 VNB N_A_28_62#_c_120_n 0.0152123f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.465
cc_9 VNB N_A_28_62#_c_121_n 0.0630269f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.465
cc_10 VNB N_A_28_62#_c_122_n 0.00104648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_28_62#_c_123_n 0.00864023f $X=-0.19 $Y=-0.245 $X2=0.747 $Y2=0.925
cc_12 VNB N_A_28_62#_c_124_n 0.0625408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_M1001_g 0.025123f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.52
cc_14 VNB N_A_M1000_g 0.00660908f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.155
cc_15 VNB N_A_c_183_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.725
cc_16 VNB N_A_M1008_g 0.0103416f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.465
cc_17 VNB N_A_c_185_n 0.00536961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A 0.0152384f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.65
cc_19 VNB N_A_c_187_n 0.0352249f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_A_c_188_n 0.0228496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_228_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Z 0.00350375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_344_n 0.00824677f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.725
cc_24 VNB N_VGND_c_345_n 0.0208062f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.465
cc_25 VNB N_VGND_c_346_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.465
cc_26 VNB N_VGND_c_347_n 0.0170192f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.65
cc_27 VNB N_VGND_c_348_n 0.0343683f $X=-0.19 $Y=-0.245 $X2=0.747 $Y2=0.925
cc_28 VNB N_VGND_c_349_n 0.205153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_350_n 0.0056753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_351_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_251_47#_c_387_n 0.00994485f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.65
cc_32 VNB N_A_251_47#_c_388_n 0.00751802f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.725
cc_33 VNB N_A_251_47#_c_389_n 0.00467732f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.465
cc_34 VNB N_A_251_47#_c_390_n 0.0303646f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.005
cc_35 VPB N_TE_B_c_67_n 0.0227252f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.725
cc_36 VPB N_TE_B_c_68_n 0.0182783f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=1.725
cc_37 VPB N_TE_B_c_62_n 0.00798339f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=1.65
cc_38 VPB N_TE_B_c_63_n 0.0124943f $X=-0.19 $Y=1.655 $X2=1.1 $Y2=1.65
cc_39 VPB N_TE_B_c_71_n 0.0186908f $X=-0.19 $Y=1.655 $X2=1.455 $Y2=1.725
cc_40 VPB N_A_28_62#_c_121_n 0.00123126f $X=-0.19 $Y=1.655 $X2=1.455 $Y2=2.465
cc_41 VPB N_A_28_62#_c_126_n 0.0316867f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=1.65
cc_42 VPB N_A_28_62#_c_127_n 0.0062101f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_43 VPB N_A_28_62#_c_122_n 5.0231e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_28_62#_c_129_n 0.0100282f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=1.005
cc_45 VPB N_A_M1000_g 0.0235689f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.155
cc_46 VPB N_A_M1008_g 0.0247854f $X=-0.19 $Y=1.655 $X2=1.455 $Y2=2.465
cc_47 VPB N_VPWR_c_229_n 0.0261036f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=1.725
cc_48 VPB N_VPWR_c_230_n 0.00918301f $X=-0.19 $Y=1.655 $X2=1.455 $Y2=2.465
cc_49 VPB N_VPWR_c_231_n 0.0212365f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=1.65
cc_50 VPB N_VPWR_c_232_n 0.0149824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_233_n 0.0450315f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_228_n 0.0567881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_235_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_236_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_220_367#_c_273_n 0.0150229f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=2.465
cc_56 VPB N_Z_c_301_n 0.00410146f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=1.65
cc_57 VPB N_Z_c_302_n 0.0123854f $X=-0.19 $Y=1.655 $X2=1.455 $Y2=1.725
cc_58 VPB N_Z_c_303_n 0.00744853f $X=-0.19 $Y=1.655 $X2=1.455 $Y2=2.465
cc_59 VPB N_Z_c_304_n 0.0459966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB Z 0.00105618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 TE_B N_A_28_62#_c_119_n 0.00339959f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_62 N_TE_B_c_65_n N_A_28_62#_c_119_n 0.00188589f $X=0.635 $Y=1.005 $X2=0 $Y2=0
cc_63 TE_B N_A_28_62#_c_121_n 0.0506183f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_64 N_TE_B_c_66_n N_A_28_62#_c_121_n 0.0308173f $X=0.612 $Y=0.84 $X2=0 $Y2=0
cc_65 N_TE_B_c_67_n N_A_28_62#_c_126_n 0.00738917f $X=0.5 $Y=1.725 $X2=0 $Y2=0
cc_66 N_TE_B_c_68_n N_A_28_62#_c_126_n 6.08913e-19 $X=1.025 $Y=1.725 $X2=0 $Y2=0
cc_67 N_TE_B_c_67_n N_A_28_62#_c_127_n 0.00988431f $X=0.5 $Y=1.725 $X2=0 $Y2=0
cc_68 N_TE_B_c_68_n N_A_28_62#_c_127_n 0.0116883f $X=1.025 $Y=1.725 $X2=0 $Y2=0
cc_69 N_TE_B_c_62_n N_A_28_62#_c_127_n 0.0137998f $X=1.38 $Y=1.65 $X2=0 $Y2=0
cc_70 N_TE_B_c_63_n N_A_28_62#_c_127_n 0.0218f $X=1.1 $Y=1.65 $X2=0 $Y2=0
cc_71 N_TE_B_c_71_n N_A_28_62#_c_127_n 0.00920173f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_72 TE_B N_A_28_62#_c_127_n 0.0305459f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_73 N_TE_B_c_62_n N_A_28_62#_c_122_n 0.00310056f $X=1.38 $Y=1.65 $X2=0 $Y2=0
cc_74 N_TE_B_c_67_n N_A_28_62#_c_129_n 0.00227117f $X=0.5 $Y=1.725 $X2=0 $Y2=0
cc_75 N_TE_B_c_63_n N_A_28_62#_c_129_n 0.00118216f $X=1.1 $Y=1.65 $X2=0 $Y2=0
cc_76 N_TE_B_c_61_n N_A_28_62#_c_124_n 0.00188589f $X=0.612 $Y=1.575 $X2=0 $Y2=0
cc_77 N_TE_B_c_62_n N_A_28_62#_c_124_n 0.00247699f $X=1.38 $Y=1.65 $X2=0 $Y2=0
cc_78 N_TE_B_c_67_n N_VPWR_c_229_n 0.00462735f $X=0.5 $Y=1.725 $X2=0 $Y2=0
cc_79 N_TE_B_c_68_n N_VPWR_c_229_n 0.00422012f $X=1.025 $Y=1.725 $X2=0 $Y2=0
cc_80 N_TE_B_c_63_n N_VPWR_c_229_n 0.00113268f $X=1.1 $Y=1.65 $X2=0 $Y2=0
cc_81 N_TE_B_c_68_n N_VPWR_c_230_n 5.84138e-19 $X=1.025 $Y=1.725 $X2=0 $Y2=0
cc_82 N_TE_B_c_71_n N_VPWR_c_230_n 0.011877f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_83 N_TE_B_c_67_n N_VPWR_c_231_n 0.00312414f $X=0.5 $Y=1.725 $X2=0 $Y2=0
cc_84 N_TE_B_c_68_n N_VPWR_c_232_n 0.00585385f $X=1.025 $Y=1.725 $X2=0 $Y2=0
cc_85 N_TE_B_c_71_n N_VPWR_c_232_n 0.00486043f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_86 N_TE_B_c_67_n N_VPWR_c_228_n 0.00410284f $X=0.5 $Y=1.725 $X2=0 $Y2=0
cc_87 N_TE_B_c_68_n N_VPWR_c_228_n 0.0118494f $X=1.025 $Y=1.725 $X2=0 $Y2=0
cc_88 N_TE_B_c_71_n N_VPWR_c_228_n 0.004514f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_89 N_TE_B_c_71_n N_A_220_367#_c_273_n 0.0127564f $X=1.455 $Y=1.725 $X2=0
+ $Y2=0
cc_90 N_TE_B_c_62_n N_A_220_367#_c_275_n 5.90216e-19 $X=1.38 $Y=1.65 $X2=0 $Y2=0
cc_91 N_TE_B_c_71_n N_A_220_367#_c_275_n 0.0149908f $X=1.455 $Y=1.725 $X2=0
+ $Y2=0
cc_92 N_TE_B_c_71_n N_Z_c_301_n 0.00658387f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_93 N_TE_B_c_62_n N_Z_c_303_n 4.93109e-19 $X=1.38 $Y=1.65 $X2=0 $Y2=0
cc_94 N_TE_B_c_71_n N_Z_c_303_n 6.56485e-19 $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_95 TE_B N_VGND_c_344_n 0.0164494f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_96 N_TE_B_c_65_n N_VGND_c_344_n 0.00142286f $X=0.635 $Y=1.005 $X2=0 $Y2=0
cc_97 N_TE_B_c_66_n N_VGND_c_344_n 0.0119198f $X=0.612 $Y=0.84 $X2=0 $Y2=0
cc_98 N_TE_B_c_66_n N_VGND_c_347_n 0.00425877f $X=0.612 $Y=0.84 $X2=0 $Y2=0
cc_99 TE_B N_VGND_c_349_n 0.00397f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_100 N_TE_B_c_66_n N_VGND_c_349_n 0.00844494f $X=0.612 $Y=0.84 $X2=0 $Y2=0
cc_101 TE_B N_A_251_47#_c_387_n 0.00989172f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_102 N_TE_B_c_65_n N_A_251_47#_c_387_n 5.44337e-19 $X=0.635 $Y=1.005 $X2=0
+ $Y2=0
cc_103 N_TE_B_c_66_n N_A_251_47#_c_387_n 0.00595579f $X=0.612 $Y=0.84 $X2=0
+ $Y2=0
cc_104 N_TE_B_c_62_n N_A_251_47#_c_388_n 0.00105347f $X=1.38 $Y=1.65 $X2=0 $Y2=0
cc_105 N_TE_B_c_62_n N_A_251_47#_c_389_n 0.00585243f $X=1.38 $Y=1.65 $X2=0 $Y2=0
cc_106 TE_B N_A_251_47#_c_389_n 0.0110258f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_107 N_TE_B_c_65_n N_A_251_47#_c_389_n 6.66796e-19 $X=0.635 $Y=1.005 $X2=0
+ $Y2=0
cc_108 N_A_28_62#_c_120_n N_A_M1001_g 0.0174207f $X=2.025 $Y=1.185 $X2=0 $Y2=0
cc_109 N_A_28_62#_c_123_n N_A_M1001_g 8.44325e-19 $X=1.935 $Y=1.44 $X2=0 $Y2=0
cc_110 N_A_28_62#_c_127_n N_A_M1000_g 0.00108015f $X=1.77 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_28_62#_c_122_n N_A_M1000_g 0.00143119f $X=1.855 $Y=1.68 $X2=0 $Y2=0
cc_112 N_A_28_62#_c_124_n N_A_c_185_n 0.0174207f $X=1.935 $Y=1.44 $X2=0 $Y2=0
cc_113 N_A_28_62#_c_127_n N_VPWR_M1006_d 0.00277448f $X=1.77 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_28_62#_c_127_n N_VPWR_M1009_d 0.00369536f $X=1.77 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_28_62#_c_126_n N_VPWR_c_229_n 0.0178223f $X=0.285 $Y=1.98 $X2=0 $Y2=0
cc_116 N_A_28_62#_c_127_n N_VPWR_c_229_n 0.0212345f $X=1.77 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_28_62#_c_126_n N_VPWR_c_228_n 0.012861f $X=0.285 $Y=1.98 $X2=0 $Y2=0
cc_118 N_A_28_62#_c_127_n N_A_220_367#_M1007_s 0.00176461f $X=1.77 $Y=1.765
+ $X2=-0.19 $Y2=-0.245
cc_119 N_A_28_62#_c_127_n N_A_220_367#_c_273_n 0.0163927f $X=1.77 $Y=1.765 $X2=0
+ $Y2=0
cc_120 N_A_28_62#_c_127_n N_A_220_367#_c_275_n 0.0152401f $X=1.77 $Y=1.765 $X2=0
+ $Y2=0
cc_121 N_A_28_62#_c_127_n N_Z_c_303_n 0.0134922f $X=1.77 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_28_62#_c_120_n Z 0.00107287f $X=2.025 $Y=1.185 $X2=0 $Y2=0
cc_123 N_A_28_62#_c_127_n Z 8.4932e-19 $X=1.77 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_28_62#_c_122_n Z 0.00408042f $X=1.855 $Y=1.68 $X2=0 $Y2=0
cc_125 N_A_28_62#_c_123_n Z 0.00696543f $X=1.935 $Y=1.44 $X2=0 $Y2=0
cc_126 N_A_28_62#_c_124_n Z 4.5165e-19 $X=1.935 $Y=1.44 $X2=0 $Y2=0
cc_127 N_A_28_62#_c_119_n N_VGND_c_344_n 0.00242395f $X=1.595 $Y=1.185 $X2=0
+ $Y2=0
cc_128 N_A_28_62#_c_119_n N_VGND_c_345_n 0.00486043f $X=1.595 $Y=1.185 $X2=0
+ $Y2=0
cc_129 N_A_28_62#_c_119_n N_VGND_c_346_n 0.0119381f $X=1.595 $Y=1.185 $X2=0
+ $Y2=0
cc_130 N_A_28_62#_c_120_n N_VGND_c_346_n 0.0113499f $X=2.025 $Y=1.185 $X2=0
+ $Y2=0
cc_131 N_A_28_62#_c_121_n N_VGND_c_347_n 0.0114303f $X=0.265 $Y=0.52 $X2=0 $Y2=0
cc_132 N_A_28_62#_c_120_n N_VGND_c_348_n 0.00486043f $X=2.025 $Y=1.185 $X2=0
+ $Y2=0
cc_133 N_A_28_62#_c_119_n N_VGND_c_349_n 0.00954696f $X=1.595 $Y=1.185 $X2=0
+ $Y2=0
cc_134 N_A_28_62#_c_120_n N_VGND_c_349_n 0.0082726f $X=2.025 $Y=1.185 $X2=0
+ $Y2=0
cc_135 N_A_28_62#_c_121_n N_VGND_c_349_n 0.00986179f $X=0.265 $Y=0.52 $X2=0
+ $Y2=0
cc_136 N_A_28_62#_c_119_n N_A_251_47#_c_388_n 0.0144827f $X=1.595 $Y=1.185 $X2=0
+ $Y2=0
cc_137 N_A_28_62#_c_120_n N_A_251_47#_c_388_n 0.0131717f $X=2.025 $Y=1.185 $X2=0
+ $Y2=0
cc_138 N_A_28_62#_c_127_n N_A_251_47#_c_388_n 0.00962964f $X=1.77 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_28_62#_c_123_n N_A_251_47#_c_388_n 0.0232349f $X=1.935 $Y=1.44 $X2=0
+ $Y2=0
cc_140 N_A_28_62#_c_124_n N_A_251_47#_c_388_n 0.00284602f $X=1.935 $Y=1.44 $X2=0
+ $Y2=0
cc_141 N_A_28_62#_c_127_n N_A_251_47#_c_389_n 0.00929937f $X=1.77 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A_M1000_g N_VPWR_c_230_n 0.00877449f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_M1000_g N_VPWR_c_233_n 0.0054895f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_M1008_g N_VPWR_c_233_n 0.00585385f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1000_g N_VPWR_c_228_n 0.00765772f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_M1008_g N_VPWR_c_228_n 0.0116979f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_M1000_g N_A_220_367#_c_273_n 0.0118778f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_M1000_g N_A_220_367#_c_281_n 0.0166062f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_M1000_g N_A_220_367#_c_282_n 9.80814e-19 $X=2.455 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_M1008_g N_Z_c_302_n 0.0184827f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_151 A N_Z_c_302_n 0.0286801f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A_c_187_n N_Z_c_302_n 0.00450443f $X=2.99 $Y=1.36 $X2=0 $Y2=0
cc_153 N_A_M1000_g N_Z_c_303_n 0.0156099f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_c_183_n N_Z_c_303_n 4.81398e-19 $X=2.81 $Y=1.45 $X2=0 $Y2=0
cc_155 N_A_M1001_g Z 0.0107017f $X=2.455 $Y=0.655 $X2=0 $Y2=0
cc_156 N_A_M1000_g Z 0.00516846f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_c_183_n Z 0.00913923f $X=2.81 $Y=1.45 $X2=0 $Y2=0
cc_158 N_A_M1008_g Z 0.00447048f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A_c_185_n Z 0.00236416f $X=2.455 $Y=1.45 $X2=0 $Y2=0
cc_160 A Z 0.0250712f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_161 N_A_c_188_n Z 0.0066875f $X=2.982 $Y=1.195 $X2=0 $Y2=0
cc_162 N_A_M1001_g N_Z_c_327_n 0.00359944f $X=2.455 $Y=0.655 $X2=0 $Y2=0
cc_163 N_A_c_188_n N_Z_c_327_n 0.00448868f $X=2.982 $Y=1.195 $X2=0 $Y2=0
cc_164 N_A_M1001_g N_VGND_c_346_n 0.00109252f $X=2.455 $Y=0.655 $X2=0 $Y2=0
cc_165 N_A_M1001_g N_VGND_c_348_n 0.00357877f $X=2.455 $Y=0.655 $X2=0 $Y2=0
cc_166 N_A_c_188_n N_VGND_c_348_n 0.00357877f $X=2.982 $Y=1.195 $X2=0 $Y2=0
cc_167 N_A_M1001_g N_VGND_c_349_n 0.00537654f $X=2.455 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A_c_188_n N_VGND_c_349_n 0.00628381f $X=2.982 $Y=1.195 $X2=0 $Y2=0
cc_169 N_A_M1001_g N_A_251_47#_c_388_n 8.03868e-19 $X=2.455 $Y=0.655 $X2=0 $Y2=0
cc_170 N_A_M1001_g N_A_251_47#_c_405_n 0.0111972f $X=2.455 $Y=0.655 $X2=0 $Y2=0
cc_171 N_A_c_188_n N_A_251_47#_c_405_n 0.0114565f $X=2.982 $Y=1.195 $X2=0 $Y2=0
cc_172 A N_A_251_47#_c_390_n 0.0213292f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A_c_187_n N_A_251_47#_c_390_n 0.00343753f $X=2.99 $Y=1.36 $X2=0 $Y2=0
cc_174 N_VPWR_c_228_n N_A_220_367#_M1007_s 0.00251545f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_175 N_VPWR_c_228_n N_A_220_367#_M1000_d 0.00240953f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_232_n N_A_220_367#_c_285_n 0.0140491f $X=1.505 $Y=3.33 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_228_n N_A_220_367#_c_285_n 0.0090585f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_178 N_VPWR_M1009_d N_A_220_367#_c_273_n 0.00662568f $X=1.53 $Y=1.835 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_230_n N_A_220_367#_c_273_n 0.0215105f $X=1.67 $Y=2.79 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_228_n N_A_220_367#_c_273_n 0.0262128f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_230_n N_A_220_367#_c_281_n 0.0113528f $X=1.67 $Y=2.79 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_233_n N_A_220_367#_c_281_n 0.0171073f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_228_n N_A_220_367#_c_281_n 0.0114026f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_228_n N_A_220_367#_c_275_n 0.00238693f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_228_n N_Z_M1000_s 0.00389753f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_186 N_VPWR_c_228_n N_Z_M1008_s 0.0026734f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_187 N_VPWR_c_233_n N_Z_c_304_n 0.0188755f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_188 N_VPWR_c_228_n N_Z_c_304_n 0.0111968f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_189 N_A_220_367#_c_273_n N_Z_M1000_s 0.00716549f $X=2.505 $Y=2.41 $X2=0 $Y2=0
cc_190 N_A_220_367#_c_273_n N_Z_c_301_n 0.016086f $X=2.505 $Y=2.41 $X2=0 $Y2=0
cc_191 N_A_220_367#_M1000_d N_Z_c_303_n 0.00157327f $X=2.53 $Y=1.835 $X2=0 $Y2=0
cc_192 N_A_220_367#_c_273_n N_Z_c_303_n 0.00385789f $X=2.505 $Y=2.41 $X2=0 $Y2=0
cc_193 N_A_220_367#_c_298_p N_Z_c_303_n 0.013469f $X=2.67 $Y=2.21 $X2=0 $Y2=0
cc_194 N_A_220_367#_c_282_n N_Z_c_303_n 8.43884e-19 $X=2.655 $Y=2.41 $X2=0 $Y2=0
cc_195 N_Z_M1001_d N_VGND_c_349_n 0.00225186f $X=2.53 $Y=0.235 $X2=0 $Y2=0
cc_196 N_Z_c_303_n N_A_251_47#_c_388_n 0.00807861f $X=2.735 $Y=1.79 $X2=0 $Y2=0
cc_197 Z N_A_251_47#_c_388_n 0.0107192f $X=2.64 $Y=0.925 $X2=0 $Y2=0
cc_198 N_Z_M1001_d N_A_251_47#_c_405_n 0.00332344f $X=2.53 $Y=0.235 $X2=0 $Y2=0
cc_199 N_Z_c_327_n N_A_251_47#_c_405_n 0.0165042f $X=2.67 $Y=0.72 $X2=0 $Y2=0
cc_200 N_VGND_c_349_n N_A_251_47#_M1004_s 0.00371702f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_201 N_VGND_c_349_n N_A_251_47#_M1005_s 0.00376627f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_349_n N_A_251_47#_M1003_s 0.00215161f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_c_344_n N_A_251_47#_c_387_n 0.0156017f $X=0.715 $Y=0.455 $X2=0
+ $Y2=0
cc_204 N_VGND_c_345_n N_A_251_47#_c_387_n 0.0178111f $X=1.645 $Y=0 $X2=0 $Y2=0
cc_205 N_VGND_c_349_n N_A_251_47#_c_387_n 0.0100304f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_206 N_VGND_M1004_d N_A_251_47#_c_388_n 0.00176461f $X=1.67 $Y=0.235 $X2=0
+ $Y2=0
cc_207 N_VGND_c_346_n N_A_251_47#_c_388_n 0.0170777f $X=1.81 $Y=0.38 $X2=0 $Y2=0
cc_208 N_VGND_c_348_n N_A_251_47#_c_421_n 0.0121686f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_209 N_VGND_c_349_n N_A_251_47#_c_421_n 0.00698742f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_348_n N_A_251_47#_c_405_n 0.0364699f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_349_n N_A_251_47#_c_405_n 0.024052f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_212 N_VGND_c_348_n N_A_251_47#_c_390_n 0.0179183f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_c_349_n N_A_251_47#_c_390_n 0.0101082f $X=3.12 $Y=0 $X2=0 $Y2=0
