* NGSPICE file created from sky130_fd_sc_lp__clkinvlp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__clkinvlp_2 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.8e+11p pd=2.56e+06u as=5.3e+11p ps=5.06e+06u
M1001 a_185_67# A VGND VNB nshort w=550000u l=150000u
+  ad=1.32e+11p pd=1.58e+06u as=1.5675e+11p ps=1.67e+06u
M1002 Y A a_185_67# VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1003 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

