* File: sky130_fd_sc_lp__srsdfstp_1.pex.spice
* Created: Wed Sep  2 10:39:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%SCD 3 7 11 12 13 14 18
r35 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.39
+ $Y=1.37 $X2=0.39 $Y2=1.37
r36 14 19 5.89113 $w=6.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=0.39 $Y2=1.54
r37 13 19 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=1.54
+ $X2=0.39 $Y2=1.54
r38 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.39 $Y=1.71
+ $X2=0.39 $Y2=1.37
r39 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.39 $Y=1.71
+ $X2=0.39 $Y2=1.875
r40 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.39 $Y=1.205
+ $X2=0.39 $Y2=1.37
r41 7 12 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=0.48 $Y=2.725
+ $X2=0.48 $Y2=1.875
r42 3 10 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.48 $Y=0.805 $X2=0.48
+ $Y2=1.205
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%D 3 7 9 12 13
c39 7 0 9.92106e-20 $X=1.38 $Y=2.725
r40 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.71
+ $X2=1.29 $Y2=1.875
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.71
+ $X2=1.29 $Y2=1.545
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.29
+ $Y=1.71 $X2=1.29 $Y2=1.71
r43 9 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.71 $X2=1.29
+ $Y2=1.71
r44 7 15 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.38 $Y=2.725
+ $X2=1.38 $Y2=1.875
r45 3 14 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.3 $Y=0.805 $X2=1.3
+ $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_339_93# 1 2 9 13 16 18 19 25
c50 19 0 1.99409e-19 $X=2.1 $Y=1.47
r51 22 25 6.36424 $w=3.33e-07 $l=1.85e-07 $layer=LI1_cond $X=2.47 $Y=0.842
+ $X2=2.655 $Y2=0.842
r52 19 29 80.5075 $w=5.7e-07 $l=5.05e-07 $layer=POLY_cond $X=1.98 $Y=1.47
+ $X2=1.98 $Y2=1.975
r53 19 28 48.5934 $w=5.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=1.47
+ $X2=1.98 $Y2=1.305
r54 18 21 8.34643 $w=6.87e-07 $l=4.7e-07 $layer=LI1_cond $X=2.33 $Y=1.47
+ $X2=2.33 $Y2=1.94
r55 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.1 $Y=1.47
+ $X2=2.1 $Y2=1.47
r56 16 18 10.936 $w=6.87e-07 $l=2.24332e-07 $layer=LI1_cond $X=2.47 $Y=1.305
+ $X2=2.33 $Y2=1.47
r57 15 22 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.47 $Y=1.01
+ $X2=2.47 $Y2=0.842
r58 15 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.47 $Y=1.01
+ $X2=2.47 $Y2=1.305
r59 13 29 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.81 $Y=2.725
+ $X2=1.81 $Y2=1.975
r60 9 28 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.77 $Y=0.805 $X2=1.77
+ $Y2=1.305
r61 2 21 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.795 $X2=2.555 $Y2=1.94
r62 1 25 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.51
+ $Y=0.695 $X2=2.655 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%SCE 2 6 9 11 12 15 20 22 25 27 30
c84 27 0 1.99409e-19 $X=3.12 $Y=1.295
c85 25 0 6.37051e-20 $X=0.99 $Y=2.16
c86 6 0 2.10137e-20 $X=0.87 $Y=0.805
r87 30 33 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.39
+ $X2=2.875 $Y2=1.555
r88 30 32 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.39
+ $X2=2.875 $Y2=1.225
r89 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.89
+ $Y=1.39 $X2=2.89 $Y2=1.39
r90 27 31 7.06832 $w=3.73e-07 $l=2.3e-07 $layer=LI1_cond $X=3.12 $Y=1.367
+ $X2=2.89 $Y2=1.367
r91 23 25 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.84 $Y=2.16
+ $X2=0.99 $Y2=2.16
r92 21 22 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.855 $Y=1.125
+ $X2=0.855 $Y2=1.275
r93 20 32 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.87 $Y=0.905
+ $X2=2.87 $Y2=1.225
r94 17 20 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.87 $Y=0.255
+ $X2=2.87 $Y2=0.905
r95 15 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.77 $Y=2.115
+ $X2=2.77 $Y2=1.555
r96 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.795 $Y=0.18
+ $X2=2.87 $Y2=0.255
r97 11 12 948.617 $w=1.5e-07 $l=1.85e-06 $layer=POLY_cond $X=2.795 $Y=0.18
+ $X2=0.945 $Y2=0.18
r98 7 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.99 $Y=2.235
+ $X2=0.99 $Y2=2.16
r99 7 9 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.99 $Y=2.235 $X2=0.99
+ $Y2=2.725
r100 6 21 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.87 $Y=0.805
+ $X2=0.87 $Y2=1.125
r101 3 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.87 $Y=0.255
+ $X2=0.945 $Y2=0.18
r102 3 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.87 $Y=0.255
+ $X2=0.87 $Y2=0.805
r103 2 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.84 $Y=2.085
+ $X2=0.84 $Y2=2.16
r104 2 22 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.84 $Y=2.085
+ $X2=0.84 $Y2=1.275
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_689_139# 1 2 7 9 10 11 13 16 20 24 28
+ 34 37 40 42 43 46 47 48 52 53 54 56 59 60 61 63 70 75 77 78 80 81 83 84 85 87
+ 88 89 93 98 99 103
c329 99 0 1.61775e-19 $X=14.205 $Y=1.745
c330 98 0 1.90565e-19 $X=14.205 $Y=1.745
c331 70 0 1.1927e-19 $X=4.015 $Y=0.42
c332 20 0 1.29262e-19 $X=8.205 $Y=0.945
c333 11 0 2.36741e-19 $X=4.905 $Y=0.255
r334 107 109 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=8.205 $Y=1.575
+ $X2=8.565 $Y2=1.575
r335 99 114 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=14.205 $Y=1.745
+ $X2=14.205 $Y2=1.91
r336 98 100 16.5504 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=14.205 $Y=1.745
+ $X2=14.205 $Y2=2.095
r337 98 99 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.205
+ $Y=1.745 $X2=14.205 $Y2=1.745
r338 93 95 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=13.27 $Y=2.095
+ $X2=13.27 $Y2=2.31
r339 89 91 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=12.06 $Y=2.31
+ $X2=12.06 $Y2=2.49
r340 87 88 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=9.425 $Y=1.885
+ $X2=9.425 $Y2=2.135
r341 84 109 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=8.645 $Y=1.575
+ $X2=8.565 $Y2=1.575
r342 83 86 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.64 $Y=1.575
+ $X2=8.64 $Y2=1.74
r343 83 85 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.64 $Y=1.575
+ $X2=8.64 $Y2=1.41
r344 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.645
+ $Y=1.575 $X2=8.645 $Y2=1.575
r345 80 81 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=5.95 $Y=1.592
+ $X2=6.12 $Y2=1.592
r346 77 78 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.17
+ $Y=1.89 $X2=4.17 $Y2=1.89
r347 75 77 1.32706 $w=3.28e-07 $l=3.8e-08 $layer=LI1_cond $X=4.132 $Y=1.89
+ $X2=4.17 $Y2=1.89
r348 74 75 14.5627 $w=3.28e-07 $l=4.17e-07 $layer=LI1_cond $X=3.715 $Y=1.89
+ $X2=4.132 $Y2=1.89
r349 71 74 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.585 $Y=1.89
+ $X2=3.715 $Y2=1.89
r350 69 103 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.85 $Y=0.42
+ $X2=3.85 $Y2=0.18
r351 68 70 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.85 $Y=0.42
+ $X2=4.015 $Y2=0.42
r352 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.85
+ $Y=0.42 $X2=3.85 $Y2=0.42
r353 65 68 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.585 $Y=0.42
+ $X2=3.85 $Y2=0.42
r354 64 93 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.355 $Y=2.095
+ $X2=13.27 $Y2=2.095
r355 63 100 3.17874 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.04 $Y=2.095
+ $X2=14.205 $Y2=2.095
r356 63 64 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=14.04 $Y=2.095
+ $X2=13.355 $Y2=2.095
r357 62 89 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.145 $Y=2.31
+ $X2=12.06 $Y2=2.31
r358 61 95 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.185 $Y=2.31
+ $X2=13.27 $Y2=2.31
r359 61 62 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=13.185 $Y=2.31
+ $X2=12.145 $Y2=2.31
r360 59 91 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.975 $Y=2.49
+ $X2=12.06 $Y2=2.49
r361 59 60 162.449 $w=1.68e-07 $l=2.49e-06 $layer=LI1_cond $X=11.975 $Y=2.49
+ $X2=9.485 $Y2=2.49
r362 57 87 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=9.45 $Y=0.765
+ $X2=9.45 $Y2=1.885
r363 56 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.4 $Y=2.405
+ $X2=9.485 $Y2=2.49
r364 56 88 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.4 $Y=2.405 $X2=9.4
+ $Y2=2.135
r365 53 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.365 $Y=0.68
+ $X2=9.45 $Y2=0.765
r366 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.365 $Y=0.68
+ $X2=8.695 $Y2=0.68
r367 52 86 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=8.61 $Y=2.905
+ $X2=8.61 $Y2=1.74
r368 49 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.61 $Y=0.765
+ $X2=8.695 $Y2=0.68
r369 49 85 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=8.61 $Y=0.765
+ $X2=8.61 $Y2=1.41
r370 47 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.525 $Y=2.99
+ $X2=8.61 $Y2=2.905
r371 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.525 $Y=2.99
+ $X2=8.015 $Y2=2.99
r372 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=2.905
+ $X2=8.015 $Y2=2.99
r373 45 46 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=7.93 $Y=1.64
+ $X2=7.93 $Y2=2.905
r374 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.845 $Y=1.555
+ $X2=7.93 $Y2=1.64
r375 43 81 112.54 $w=1.68e-07 $l=1.725e-06 $layer=LI1_cond $X=7.845 $Y=1.555
+ $X2=6.12 $Y2=1.555
r376 42 80 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.28 $Y=1.63
+ $X2=5.95 $Y2=1.63
r377 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.195 $Y=1.545
+ $X2=5.28 $Y2=1.63
r378 39 40 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=5.195 $Y=0.425
+ $X2=5.195 $Y2=1.545
r379 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.11 $Y=0.34
+ $X2=5.195 $Y2=0.425
r380 37 70 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=5.11 $Y=0.34
+ $X2=4.015 $Y2=0.34
r381 32 71 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=1.725
+ $X2=3.585 $Y2=1.89
r382 32 34 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=3.585 $Y=1.725
+ $X2=3.585 $Y2=0.905
r383 31 65 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0.585
+ $X2=3.585 $Y2=0.42
r384 31 34 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.585 $Y=0.585
+ $X2=3.585 $Y2=0.905
r385 30 78 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.17 $Y=2.245
+ $X2=4.17 $Y2=1.89
r386 28 114 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.185 $Y=2.57
+ $X2=14.185 $Y2=1.91
r387 22 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.41
+ $X2=8.565 $Y2=1.575
r388 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.565 $Y=1.41
+ $X2=8.565 $Y2=0.945
r389 18 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.205 $Y=1.41
+ $X2=8.205 $Y2=1.575
r390 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.205 $Y=1.41
+ $X2=8.205 $Y2=0.945
r391 14 16 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=5.155 $Y=2.395
+ $X2=5.155 $Y2=2.885
r392 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.905 $Y=0.255
+ $X2=4.905 $Y2=0.575
r393 10 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.335 $Y=2.32
+ $X2=4.17 $Y2=2.245
r394 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.08 $Y=2.32
+ $X2=5.155 $Y2=2.395
r395 9 10 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=5.08 $Y=2.32
+ $X2=4.335 $Y2=2.32
r396 8 103 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=0.18
+ $X2=3.85 $Y2=0.18
r397 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.83 $Y=0.18
+ $X2=4.905 $Y2=0.255
r398 7 8 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.83 $Y=0.18
+ $X2=4.015 $Y2=0.18
r399 2 74 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.575
+ $Y=1.795 $X2=3.715 $Y2=1.94
r400 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.695 $X2=3.585 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_659_113# 1 2 7 9 10 12 13 14 15 17 18
+ 22 24 26 27 28 29 31 32 36 38 43 44 45 48 49 51 52 54 55 56 58 59 60 62 63 64
+ 66 69 70 72 75 76 77 78 80 81 85 86 87 98
c352 85 0 9.34843e-20 $X=15.49 $Y=1.9
c353 81 0 1.58197e-19 $X=14.255 $Y=0.72
c354 75 0 3.92185e-19 $X=12.59 $Y=1.545
c355 59 0 1.29262e-19 $X=7.535 $Y=1.215
c356 49 0 8.63062e-21 $X=5.615 $Y=1.29
c357 48 0 1.82358e-19 $X=5.615 $Y=1.29
c358 24 0 1.37287e-19 $X=8.485 $Y=2.145
c359 15 0 1.1927e-19 $X=4.36 $Y=1.225
c360 10 0 4.32663e-20 $X=3.5 $Y=1.375
r361 102 103 44.4629 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=5.615 $Y=1.3
+ $X2=5.615 $Y2=1.455
r362 95 98 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=15.49 $Y=2.025
+ $X2=15.6 $Y2=2.025
r363 87 89 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13.27 $Y=0.68
+ $X2=13.27 $Y2=0.985
r364 85 95 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.49 $Y=1.9
+ $X2=15.49 $Y2=2.025
r365 84 85 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=15.49 $Y=0.845
+ $X2=15.49 $Y2=1.9
r366 81 93 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=14.17 $Y=0.72
+ $X2=14.17 $Y2=0.985
r367 81 83 28.5806 $w=2.48e-07 $l=6.2e-07 $layer=LI1_cond $X=14.255 $Y=0.72
+ $X2=14.875 $Y2=0.72
r368 80 84 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=15.405 $Y=0.72
+ $X2=15.49 $Y2=0.845
r369 80 83 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=15.405 $Y=0.72
+ $X2=14.875 $Y2=0.72
r370 79 89 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.355 $Y=0.985
+ $X2=13.27 $Y2=0.985
r371 78 93 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.085 $Y=0.985
+ $X2=14.17 $Y2=0.985
r372 78 79 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=14.085 $Y=0.985
+ $X2=13.355 $Y2=0.985
r373 76 87 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.185 $Y=0.68
+ $X2=13.27 $Y2=0.68
r374 76 77 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=13.185 $Y=0.68
+ $X2=12.675 $Y2=0.68
r375 74 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.59 $Y=0.765
+ $X2=12.675 $Y2=0.68
r376 74 75 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=12.59 $Y=0.765
+ $X2=12.59 $Y2=1.545
r377 73 86 2.11342 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=1.63
+ $X2=10.25 $Y2=1.63
r378 72 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.505 $Y=1.63
+ $X2=12.59 $Y2=1.545
r379 72 73 136.353 $w=1.68e-07 $l=2.09e-06 $layer=LI1_cond $X=12.505 $Y=1.63
+ $X2=10.415 $Y2=1.63
r380 70 106 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.25 $Y=1.98
+ $X2=10.25 $Y2=2.07
r381 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.25
+ $Y=1.98 $X2=10.25 $Y2=1.98
r382 67 86 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=10.29 $Y=1.715
+ $X2=10.25 $Y2=1.63
r383 67 69 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=10.29 $Y=1.715
+ $X2=10.29 $Y2=1.98
r384 66 86 4.3182 $w=2.1e-07 $l=1.18427e-07 $layer=LI1_cond $X=10.17 $Y=1.545
+ $X2=10.25 $Y2=1.63
r385 65 66 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=10.17 $Y=0.425
+ $X2=10.17 $Y2=1.545
r386 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.085 $Y=0.34
+ $X2=10.17 $Y2=0.425
r387 63 64 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=10.085 $Y=0.34
+ $X2=7.705 $Y2=0.34
r388 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.62 $Y=0.425
+ $X2=7.705 $Y2=0.34
r389 61 62 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.62 $Y=0.425
+ $X2=7.62 $Y2=1.13
r390 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.535 $Y=1.215
+ $X2=7.62 $Y2=1.13
r391 59 60 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=7.535 $Y=1.215
+ $X2=6.895 $Y2=1.215
r392 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.81 $Y=1.13
+ $X2=6.895 $Y2=1.215
r393 57 58 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.81 $Y=0.425
+ $X2=6.81 $Y2=1.13
r394 55 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.725 $Y=0.34
+ $X2=6.81 $Y2=0.425
r395 55 56 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.725 $Y=0.34
+ $X2=6.135 $Y2=0.34
r396 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.05 $Y=0.425
+ $X2=6.135 $Y2=0.34
r397 53 54 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.05 $Y=0.425
+ $X2=6.05 $Y2=0.675
r398 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.965 $Y=0.76
+ $X2=6.05 $Y2=0.675
r399 51 52 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.965 $Y=0.76
+ $X2=5.78 $Y2=0.76
r400 49 102 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.615 $Y=1.29
+ $X2=5.615 $Y2=1.3
r401 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.615
+ $Y=1.29 $X2=5.615 $Y2=1.29
r402 46 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.615 $Y=0.845
+ $X2=5.78 $Y2=0.76
r403 46 48 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.615 $Y=0.845
+ $X2=5.615 $Y2=1.29
r404 40 42 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=3.37 $Y=1.3 $X2=3.5
+ $Y2=1.3
r405 39 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.65 $Y=2.07
+ $X2=9.575 $Y2=2.07
r406 38 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.085 $Y=2.07
+ $X2=10.25 $Y2=2.07
r407 38 39 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.085 $Y=2.07
+ $X2=9.65 $Y2=2.07
r408 34 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.575 $Y=1.995
+ $X2=9.575 $Y2=2.07
r409 34 36 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=9.575 $Y=1.995
+ $X2=9.575 $Y2=0.835
r410 33 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.92 $Y=2.07
+ $X2=8.845 $Y2=2.07
r411 32 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.5 $Y=2.07
+ $X2=9.575 $Y2=2.07
r412 32 33 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.5 $Y=2.07
+ $X2=8.92 $Y2=2.07
r413 29 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.845 $Y=2.145
+ $X2=8.845 $Y2=2.07
r414 29 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.845 $Y=2.145
+ $X2=8.845 $Y2=2.675
r415 27 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.77 $Y=2.07
+ $X2=8.845 $Y2=2.07
r416 27 28 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.77 $Y=2.07
+ $X2=8.56 $Y2=2.07
r417 24 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.485 $Y=2.145
+ $X2=8.56 $Y2=2.07
r418 24 26 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.485 $Y=2.145
+ $X2=8.485 $Y2=2.675
r419 22 103 733.255 $w=1.5e-07 $l=1.43e-06 $layer=POLY_cond $X=5.585 $Y=2.885
+ $X2=5.585 $Y2=1.455
r420 19 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.435 $Y=1.3
+ $X2=4.36 $Y2=1.3
r421 18 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.45 $Y=1.3
+ $X2=5.615 $Y2=1.3
r422 18 19 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=5.45 $Y=1.3
+ $X2=4.435 $Y2=1.3
r423 15 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.36 $Y=1.225
+ $X2=4.36 $Y2=1.3
r424 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.36 $Y=1.225
+ $X2=4.36 $Y2=0.905
r425 14 42 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.575 $Y=1.3
+ $X2=3.5 $Y2=1.3
r426 13 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.285 $Y=1.3
+ $X2=4.36 $Y2=1.3
r427 13 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.285 $Y=1.3
+ $X2=3.575 $Y2=1.3
r428 10 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.5 $Y=1.375
+ $X2=3.5 $Y2=1.3
r429 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.5 $Y=1.375
+ $X2=3.5 $Y2=2.115
r430 7 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.37 $Y=1.225
+ $X2=3.37 $Y2=1.3
r431 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.37 $Y=1.225
+ $X2=3.37 $Y2=0.905
r432 2 98 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.46
+ $Y=1.92 $X2=15.6 $Y2=2.065
r433 1 83 182 $w=1.7e-07 $l=3.85746e-07 $layer=licon1_NDIFF $count=1 $X=14.73
+ $Y=0.36 $X2=14.875 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1068_21# 1 2 7 9 10 11 14 16 18 23 27
+ 31 33 34 40
c95 40 0 1.82358e-19 $X=6.065 $Y=2.185
c96 34 0 1.6215e-19 $X=6.845 $Y=2.375
c97 33 0 1.26986e-19 $X=6.23 $Y=2.365
c98 23 0 1.88211e-20 $X=6.68 $Y=2.375
c99 18 0 1.63324e-19 $X=6.305 $Y=1.157
r100 34 37 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=6.845 $Y=2.375
+ $X2=6.845 $Y2=2.48
r101 31 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=2.35
+ $X2=6.065 $Y2=2.515
r102 31 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=2.35
+ $X2=6.065 $Y2=2.185
r103 30 33 8.02406 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=2.365
+ $X2=6.23 $Y2=2.365
r104 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=2.35 $X2=6.065 $Y2=2.35
r105 25 27 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.43 $Y=1.015
+ $X2=6.43 $Y2=0.76
r106 23 34 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.68 $Y=2.375
+ $X2=6.845 $Y2=2.375
r107 23 33 23.5727 $w=2.18e-07 $l=4.5e-07 $layer=LI1_cond $X=6.68 $Y=2.375
+ $X2=6.23 $Y2=2.375
r108 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.155
+ $Y=1.18 $X2=6.155 $Y2=1.18
r109 18 25 6.85451 $w=2.85e-07 $l=1.94715e-07 $layer=LI1_cond $X=6.305 $Y=1.157
+ $X2=6.43 $Y2=1.015
r110 18 20 6.06549 $w=2.83e-07 $l=1.5e-07 $layer=LI1_cond $X=6.305 $Y=1.157
+ $X2=6.155 $Y2=1.157
r111 16 21 39.393 $w=2.52e-07 $l=1.65e-07 $layer=POLY_cond $X=6.155 $Y=1.345
+ $X2=6.155 $Y2=1.18
r112 16 40 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.155 $Y=1.345
+ $X2=6.155 $Y2=2.185
r113 14 41 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.975 $Y=2.885
+ $X2=5.975 $Y2=2.515
r114 10 21 65.0317 $w=2.52e-07 $l=4.14367e-07 $layer=POLY_cond $X=5.99 $Y=0.84
+ $X2=6.155 $Y2=1.18
r115 10 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=5.99 $Y=0.84 $X2=5.49
+ $Y2=0.84
r116 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.415 $Y=0.765
+ $X2=5.49 $Y2=0.84
r117 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.415 $Y=0.765
+ $X2=5.415 $Y2=0.445
r118 2 37 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=6.59
+ $Y=2.675 $X2=6.845 $Y2=2.48
r119 1 27 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.245
+ $Y=0.485 $X2=6.39 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_887_139# 1 2 9 13 17 21 24 25 26 29 33
+ 36 38 39 44 46 47
c130 39 0 2.7285e-20 $X=7.51 $Y=1.93
c131 36 0 2.08416e-20 $X=6.605 $Y=1.93
c132 24 0 9.456e-20 $X=4.855 $Y=1.905
c133 21 0 1.6215e-19 $X=7.63 $Y=2.675
c134 9 0 1.26986e-19 $X=6.515 $Y=2.885
r135 42 44 7.28048 $w=4.58e-07 $l=2.8e-07 $layer=LI1_cond $X=4.575 $Y=0.905
+ $X2=4.855 $Y2=0.905
r136 39 52 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.525 $Y=1.93
+ $X2=7.525 $Y2=2.095
r137 39 51 72.229 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=7.525 $Y=1.93
+ $X2=7.525 $Y2=1.605
r138 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.51
+ $Y=1.93 $X2=7.51 $Y2=1.93
r139 36 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.605 $Y=1.93
+ $X2=6.605 $Y2=2.095
r140 35 38 36.5951 $w=2.83e-07 $l=9.05e-07 $layer=LI1_cond $X=6.605 $Y=1.952
+ $X2=7.51 $Y2=1.952
r141 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.605
+ $Y=1.93 $X2=6.605 $Y2=1.93
r142 33 47 7.14116 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=6.582 $Y=1.952
+ $X2=6.44 $Y2=1.952
r143 33 35 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=6.582 $Y=1.952
+ $X2=6.605 $Y2=1.952
r144 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.535 $Y=1.99
+ $X2=5.37 $Y2=1.99
r145 32 47 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=5.535 $Y=1.99
+ $X2=6.44 $Y2=1.99
r146 27 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.37 $Y=2.075
+ $X2=5.37 $Y2=1.99
r147 27 29 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5.37 $Y=2.075
+ $X2=5.37 $Y2=2.865
r148 25 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=1.99
+ $X2=5.37 $Y2=1.99
r149 25 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.205 $Y=1.99
+ $X2=4.94 $Y2=1.99
r150 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.855 $Y=1.905
+ $X2=4.94 $Y2=1.99
r151 23 44 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.855 $Y=1.135
+ $X2=4.855 $Y2=0.905
r152 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.855 $Y=1.135
+ $X2=4.855 $Y2=1.905
r153 21 52 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.63 $Y=2.675
+ $X2=7.63 $Y2=2.095
r154 17 51 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.63 $Y=0.945
+ $X2=7.63 $Y2=1.605
r155 11 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.605 $Y=1.765
+ $X2=6.605 $Y2=1.93
r156 11 13 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=6.605 $Y=1.765
+ $X2=6.605 $Y2=0.695
r157 9 49 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.515 $Y=2.885
+ $X2=6.515 $Y2=2.095
r158 2 29 600 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=5.23
+ $Y=2.675 $X2=5.37 $Y2=2.865
r159 1 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.435
+ $Y=0.695 $X2=4.575 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1972_99# 1 2 9 11 12 15 17 23 25 26 27
+ 28 30 34 37 38 40 44 46 51 53 54 59
c143 54 0 1.58197e-19 $X=14.59 $Y=1.205
c144 53 0 1.55755e-19 $X=14.59 $Y=1.205
c145 40 0 1.08965e-19 $X=10.82 $Y=1.97
r146 54 63 41.5123 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=14.59 $Y=1.205
+ $X2=14.59 $Y2=1.37
r147 53 56 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=14.59 $Y=1.205
+ $X2=14.59 $Y2=1.325
r148 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.59
+ $Y=1.205 $X2=14.59 $Y2=1.205
r149 46 49 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=11.64 $Y=1.97
+ $X2=11.64 $Y2=2.15
r150 44 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.82 $Y=2.05
+ $X2=10.82 $Y2=1.885
r151 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.82
+ $Y=2.05 $X2=10.82 $Y2=2.05
r152 40 43 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.82 $Y=1.97
+ $X2=10.82 $Y2=2.05
r153 39 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.015 $Y=1.325
+ $X2=12.93 $Y2=1.325
r154 38 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.425 $Y=1.325
+ $X2=14.59 $Y2=1.325
r155 38 39 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=14.425 $Y=1.325
+ $X2=13.015 $Y2=1.325
r156 36 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.93 $Y=1.41
+ $X2=12.93 $Y2=1.325
r157 36 37 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=12.93 $Y=1.41
+ $X2=12.93 $Y2=1.885
r158 32 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.93 $Y=1.24
+ $X2=12.93 $Y2=1.325
r159 32 34 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=12.93 $Y=1.24
+ $X2=12.93 $Y2=1.1
r160 31 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.805 $Y=1.97
+ $X2=11.64 $Y2=1.97
r161 30 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.845 $Y=1.97
+ $X2=12.93 $Y2=1.885
r162 30 31 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=12.845 $Y=1.97
+ $X2=11.805 $Y2=1.97
r163 29 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.985 $Y=1.97
+ $X2=10.82 $Y2=1.97
r164 28 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.475 $Y=1.97
+ $X2=11.64 $Y2=1.97
r165 28 29 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=11.475 $Y=1.97
+ $X2=10.985 $Y2=1.97
r166 27 63 227.895 $w=1.75e-07 $l=5.7e-07 $layer=POLY_cond $X=14.667 $Y=1.94
+ $X2=14.667 $Y2=1.37
r167 23 27 36.7171 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=14.705 $Y=2.065
+ $X2=14.705 $Y2=1.94
r168 23 25 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=14.705 $Y=2.065
+ $X2=14.705 $Y2=2.57
r169 19 59 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=10.73 $Y=1.575
+ $X2=10.73 $Y2=1.885
r170 18 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.37 $Y=1.5
+ $X2=10.295 $Y2=1.5
r171 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.655 $Y=1.5
+ $X2=10.73 $Y2=1.575
r172 17 18 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.655 $Y=1.5
+ $X2=10.37 $Y2=1.5
r173 13 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.295 $Y=1.425
+ $X2=10.295 $Y2=1.5
r174 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=10.295 $Y=1.425
+ $X2=10.295 $Y2=0.835
r175 11 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.22 $Y=1.5
+ $X2=10.295 $Y2=1.5
r176 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.22 $Y=1.5
+ $X2=10.01 $Y2=1.5
r177 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.935 $Y=1.425
+ $X2=10.01 $Y2=1.5
r178 7 9 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=9.935 $Y=1.425
+ $X2=9.935 $Y2=0.835
r179 2 49 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.495
+ $Y=2.005 $X2=11.64 $Y2=2.15
r180 1 34 182 $w=1.7e-07 $l=6.19516e-07 $layer=licon1_NDIFF $count=1 $X=12.675
+ $Y=0.595 $X2=12.93 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_2216_99# 1 2 7 9 11 12 14 17 20 23 26
+ 27 28 29 32 33 34 35 37 39 43 49
c166 43 0 1.97565e-19 $X=13.69 $Y=0.63
c167 29 0 9.74383e-20 $X=15.745 $Y=0.34
c168 23 0 1.0685e-19 $X=11.79 $Y=1.29
c169 14 0 4.66987e-20 $X=13.165 $Y=2.57
c170 12 0 1.59391e-19 $X=13.165 $Y=1.37
r171 43 51 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=13.69 $Y=0.63
+ $X2=13.395 $Y2=0.63
r172 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.69
+ $Y=0.63 $X2=13.69 $Y2=0.63
r173 39 42 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=13.69 $Y=0.34
+ $X2=13.69 $Y2=0.63
r174 35 47 11.4375 $w=3.36e-07 $l=4.45477e-07 $layer=LI1_cond $X=16.645 $Y=1.05
+ $X2=16.96 $Y2=0.735
r175 35 37 30.7824 $w=3.78e-07 $l=1.015e-06 $layer=LI1_cond $X=16.645 $Y=1.05
+ $X2=16.645 $Y2=2.065
r176 33 35 9.87124 $w=3.36e-07 $l=2.28583e-07 $layer=LI1_cond $X=16.455 $Y=0.965
+ $X2=16.645 $Y2=1.05
r177 33 34 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=16.455 $Y=0.965
+ $X2=15.915 $Y2=0.965
r178 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.83 $Y=0.88
+ $X2=15.915 $Y2=0.965
r179 31 32 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=15.83 $Y=0.425
+ $X2=15.83 $Y2=0.88
r180 30 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.855 $Y=0.34
+ $X2=13.69 $Y2=0.34
r181 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.745 $Y=0.34
+ $X2=15.83 $Y2=0.425
r182 29 30 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=15.745 $Y=0.34
+ $X2=13.855 $Y2=0.34
r183 27 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.525 $Y=0.34
+ $X2=13.69 $Y2=0.34
r184 27 28 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=13.525 $Y=0.34
+ $X2=12.335 $Y2=0.34
r185 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.25 $Y=0.425
+ $X2=12.335 $Y2=0.34
r186 25 26 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=12.25 $Y=0.425
+ $X2=12.25 $Y2=1.125
r187 23 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.79 $Y=1.29
+ $X2=11.625 $Y2=1.29
r188 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.79
+ $Y=1.29 $X2=11.79 $Y2=1.29
r189 20 26 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.165 $Y=1.25
+ $X2=12.25 $Y2=1.125
r190 20 22 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=12.165 $Y=1.25
+ $X2=11.79 $Y2=1.25
r191 16 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.395 $Y=0.795
+ $X2=13.395 $Y2=0.63
r192 16 17 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=13.395 $Y=0.795
+ $X2=13.395 $Y2=1.22
r193 12 17 87.9841 $w=1.26e-07 $l=2.3e-07 $layer=POLY_cond $X=13.165 $Y=1.295
+ $X2=13.395 $Y2=1.295
r194 12 14 298.144 $w=2.5e-07 $l=1.2e-06 $layer=POLY_cond $X=13.165 $Y=1.37
+ $X2=13.165 $Y2=2.57
r195 11 49 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=11.23 $Y=1.23
+ $X2=11.625 $Y2=1.23
r196 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.155 $Y=1.155
+ $X2=11.23 $Y2=1.23
r197 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.155 $Y=1.155
+ $X2=11.155 $Y2=0.835
r198 2 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=16.53
+ $Y=1.92 $X2=16.67 $Y2=2.065
r199 1 47 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=16.82
+ $Y=0.36 $X2=16.96 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1728_125# 1 2 3 11 12 13 16 18 20 23 26
+ 27 28 29 31 33 36 40 42 43 45 48 53 57 60 63 65 68 72 78 79 81 82 87
c217 81 0 1.37034e-20 $X=17.17 $Y=1.66
c218 78 0 1.61775e-19 $X=14.425 $Y=2.42
c219 43 0 1.37287e-19 $X=9.02 $Y=2.62
c220 13 0 1.08965e-19 $X=11.375 $Y=1.82
r221 81 84 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=17.17 $Y=1.66
+ $X2=17.17 $Y2=1.825
r222 81 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.17
+ $Y=1.66 $X2=17.17 $Y2=1.66
r223 78 79 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=14.425 $Y=2.42
+ $X2=14.595 $Y2=2.42
r224 75 76 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=13.965 $Y=2.54
+ $X2=13.965 $Y2=2.65
r225 72 75 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=13.965 $Y=2.435
+ $X2=13.965 $Y2=2.54
r226 60 84 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=17.135 $Y=2.32
+ $X2=17.135 $Y2=1.825
r227 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.05 $Y=2.405
+ $X2=17.135 $Y2=2.32
r228 57 79 160.166 $w=1.68e-07 $l=2.455e-06 $layer=LI1_cond $X=17.05 $Y=2.405
+ $X2=14.595 $Y2=2.405
r229 56 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.13 $Y=2.435
+ $X2=13.965 $Y2=2.435
r230 56 78 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=14.13 $Y=2.435
+ $X2=14.425 $Y2=2.435
r231 54 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.485 $Y=2.65
+ $X2=12.4 $Y2=2.65
r232 53 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.8 $Y=2.65
+ $X2=13.965 $Y2=2.65
r233 53 54 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=13.8 $Y=2.65
+ $X2=12.485 $Y2=2.65
r234 52 87 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=11.17 $Y=2.91
+ $X2=11.3 $Y2=2.91
r235 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.17
+ $Y=2.91 $X2=11.17 $Y2=2.91
r236 49 67 3.16498 $w=3.3e-07 $l=1.53297e-07 $layer=LI1_cond $X=9.145 $Y=2.91
+ $X2=9.02 $Y2=2.847
r237 49 51 70.7181 $w=3.28e-07 $l=2.025e-06 $layer=LI1_cond $X=9.145 $Y=2.91
+ $X2=11.17 $Y2=2.91
r238 48 68 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.4 $Y=2.91
+ $X2=12.4 $Y2=2.65
r239 48 51 39.9863 $w=3.28e-07 $l=1.145e-06 $layer=LI1_cond $X=12.315 $Y=2.91
+ $X2=11.17 $Y2=2.91
r240 46 63 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.01 $Y=1.225
+ $X2=9.01 $Y2=1.08
r241 46 65 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=9.01 $Y=1.225
+ $X2=9.01 $Y2=2.235
r242 43 67 3.82155 $w=2.5e-07 $l=2.27e-07 $layer=LI1_cond $X=9.02 $Y=2.62
+ $X2=9.02 $Y2=2.847
r243 43 45 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=9.02 $Y=2.62
+ $X2=9.02 $Y2=2.4
r244 42 65 6.44059 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=9.02 $Y=2.36
+ $X2=9.02 $Y2=2.235
r245 42 45 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=9.02 $Y=2.36 $X2=9.02
+ $Y2=2.4
r246 34 36 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=17.705 $Y=0.795
+ $X2=17.705 $Y2=0.445
r247 31 33 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=17.69 $Y=1.905
+ $X2=17.69 $Y2=2.335
r248 30 82 27.8707 $w=2.94e-07 $l=2.38642e-07 $layer=POLY_cond $X=17.335 $Y=1.83
+ $X2=17.17 $Y2=1.66
r249 29 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.615 $Y=1.83
+ $X2=17.69 $Y2=1.905
r250 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=17.615 $Y=1.83
+ $X2=17.335 $Y2=1.83
r251 27 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.63 $Y=0.87
+ $X2=17.705 $Y2=0.795
r252 27 28 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=17.63 $Y=0.87
+ $X2=17.335 $Y2=0.87
r253 26 82 38.5845 $w=2.94e-07 $l=2.05122e-07 $layer=POLY_cond $X=17.26 $Y=1.495
+ $X2=17.17 $Y2=1.66
r254 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.26 $Y=0.945
+ $X2=17.335 $Y2=0.87
r255 25 26 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=17.26 $Y=0.945
+ $X2=17.26 $Y2=1.495
r256 21 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.6 $Y=1.745
+ $X2=12.6 $Y2=1.82
r257 21 23 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=12.6 $Y=1.745 $X2=12.6
+ $Y2=0.805
r258 18 40 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=12.475 $Y=1.82
+ $X2=12.6 $Y2=1.82
r259 18 38 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=12.475 $Y=1.82
+ $X2=12.24 $Y2=1.82
r260 18 20 117.608 $w=2.5e-07 $l=6.1e-07 $layer=POLY_cond $X=12.475 $Y=1.895
+ $X2=12.475 $Y2=2.505
r261 14 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.24 $Y=1.745
+ $X2=12.24 $Y2=1.82
r262 14 16 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=12.24 $Y=1.745
+ $X2=12.24 $Y2=0.805
r263 12 38 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.165 $Y=1.82
+ $X2=12.24 $Y2=1.82
r264 12 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=12.165 $Y=1.82
+ $X2=11.375 $Y2=1.82
r265 11 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.3 $Y=2.745
+ $X2=11.3 $Y2=2.91
r266 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.3 $Y=1.895
+ $X2=11.375 $Y2=1.82
r267 10 11 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=11.3 $Y=1.895
+ $X2=11.3 $Y2=2.745
r268 3 75 600 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_PDIFF $count=1 $X=13.78
+ $Y=2.07 $X2=13.92 $Y2=2.54
r269 2 67 600 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=1 $X=8.92
+ $Y=2.255 $X2=9.06 $Y2=2.865
r270 2 45 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.92
+ $Y=2.255 $X2=9.06 $Y2=2.4
r271 1 63 182 $w=1.7e-07 $l=6.82697e-07 $layer=licon1_NDIFF $count=1 $X=8.64
+ $Y=0.625 $X2=9.03 $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%SET_B 4 7 9 10 13 15 19 23 24 26 28 29 30
+ 33 35
c122 35 0 9.38031e-20 $X=13.665 $Y=1.58
c123 23 0 2.52517e-19 $X=14.065 $Y=1.265
c124 7 0 1.88211e-20 $X=7.06 $Y=2.465
c125 4 0 1.63324e-19 $X=7 $Y=0.695
r126 33 36 34.1291 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=13.665 $Y=1.745
+ $X2=13.665 $Y2=1.92
r127 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.665 $Y=1.745
+ $X2=13.665 $Y2=1.58
r128 30 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.665
+ $Y=1.745 $X2=13.665 $Y2=1.745
r129 27 28 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=7.03 $Y=1.34
+ $X2=7.03 $Y2=1.49
r130 25 26 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=14.14 $Y=0.255
+ $X2=14.14 $Y2=1.19
r131 23 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.065 $Y=1.265
+ $X2=14.14 $Y2=1.19
r132 23 24 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=14.065 $Y=1.265
+ $X2=13.83 $Y2=1.265
r133 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.755 $Y=1.34
+ $X2=13.83 $Y2=1.265
r134 21 35 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=13.755 $Y=1.34
+ $X2=13.755 $Y2=1.58
r135 19 36 161.495 $w=2.5e-07 $l=6.5e-07 $layer=POLY_cond $X=13.655 $Y=2.57
+ $X2=13.655 $Y2=1.92
r136 16 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.8 $Y=0.18
+ $X2=10.725 $Y2=0.18
r137 15 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.065 $Y=0.18
+ $X2=14.14 $Y2=0.255
r138 15 16 1674.18 $w=1.5e-07 $l=3.265e-06 $layer=POLY_cond $X=14.065 $Y=0.18
+ $X2=10.8 $Y2=0.18
r139 11 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.725 $Y=0.255
+ $X2=10.725 $Y2=0.18
r140 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.725 $Y=0.255
+ $X2=10.725 $Y2=0.835
r141 9 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.65 $Y=0.18
+ $X2=10.725 $Y2=0.18
r142 9 10 1833.14 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=10.65 $Y=0.18
+ $X2=7.075 $Y2=0.18
r143 7 28 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=7.06 $Y=2.465
+ $X2=7.06 $Y2=1.49
r144 4 27 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=7 $Y=0.695 $X2=7
+ $Y2=1.34
r145 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7 $Y=0.255
+ $X2=7.075 $Y2=0.18
r146 1 4 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7 $Y=0.255 $X2=7
+ $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%CLK 3 7 9 10 11 20
c41 20 0 1.53981e-19 $X=15.385 $Y=1.51
r42 19 20 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=15.205 $Y=1.51
+ $X2=15.385 $Y2=1.51
r43 16 19 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=15.13 $Y=1.51
+ $X2=15.205 $Y2=1.51
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.13
+ $Y=1.51 $X2=15.13 $Y2=1.51
r45 10 11 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=15.1 $Y=1.665
+ $X2=15.1 $Y2=2.035
r46 10 17 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=15.1 $Y=1.665
+ $X2=15.1 $Y2=1.51
r47 9 17 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=15.1 $Y=1.295
+ $X2=15.1 $Y2=1.51
r48 5 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.385 $Y=1.675
+ $X2=15.385 $Y2=1.51
r49 5 7 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=15.385 $Y=1.675
+ $X2=15.385 $Y2=2.24
r50 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.205 $Y=1.345
+ $X2=15.205 $Y2=1.51
r51 1 3 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=15.205 $Y=1.345
+ $X2=15.205 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%SLEEP_B 3 7 11 13 15 18 24 26 27 28 36 38
c76 36 0 1.53981e-19 $X=16.095 $Y=1.385
c77 18 0 9.74383e-20 $X=16.385 $Y=0.57
c78 11 0 9.34843e-20 $X=15.955 $Y=0.57
r79 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.095
+ $Y=1.385 $X2=16.095 $Y2=1.385
r80 33 35 17.4819 $w=3.86e-07 $l=1.4e-07 $layer=POLY_cond $X=15.955 $Y=1.252
+ $X2=16.095 $Y2=1.252
r81 32 33 17.4819 $w=3.86e-07 $l=1.4e-07 $layer=POLY_cond $X=15.815 $Y=1.252
+ $X2=15.955 $Y2=1.252
r82 27 28 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=16.097 $Y=1.665
+ $X2=16.097 $Y2=2.035
r83 27 36 9.92874 $w=3.23e-07 $l=2.8e-07 $layer=LI1_cond $X=16.097 $Y=1.665
+ $X2=16.097 $Y2=1.385
r84 22 38 36.2124 $w=3.86e-07 $l=2.9e-07 $layer=POLY_cond $X=16.745 $Y=1.252
+ $X2=16.455 $Y2=1.252
r85 22 24 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=16.745 $Y=1.105
+ $X2=16.745 $Y2=0.57
r86 20 38 24.9932 $w=1.5e-07 $l=2.98e-07 $layer=POLY_cond $X=16.455 $Y=1.55
+ $X2=16.455 $Y2=1.252
r87 20 26 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=16.455 $Y=1.55
+ $X2=16.455 $Y2=1.79
r88 16 38 8.74093 $w=3.86e-07 $l=7e-08 $layer=POLY_cond $X=16.385 $Y=1.252
+ $X2=16.455 $Y2=1.252
r89 16 35 36.2124 $w=3.86e-07 $l=2.9e-07 $layer=POLY_cond $X=16.385 $Y=1.252
+ $X2=16.095 $Y2=1.252
r90 16 18 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=16.385 $Y=1.105
+ $X2=16.385 $Y2=0.57
r91 13 26 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=16.405 $Y=1.915
+ $X2=16.405 $Y2=1.79
r92 13 15 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=16.405 $Y=1.915
+ $X2=16.405 $Y2=2.42
r93 9 33 24.9932 $w=1.5e-07 $l=2.97e-07 $layer=POLY_cond $X=15.955 $Y=0.955
+ $X2=15.955 $Y2=1.252
r94 9 11 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=15.955 $Y=0.955
+ $X2=15.955 $Y2=0.57
r95 5 32 24.9932 $w=1.5e-07 $l=2.98e-07 $layer=POLY_cond $X=15.815 $Y=1.55
+ $X2=15.815 $Y2=1.252
r96 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=15.815 $Y=1.55
+ $X2=15.815 $Y2=2.24
r97 1 32 27.4715 $w=3.86e-07 $l=3.91853e-07 $layer=POLY_cond $X=15.595 $Y=0.955
+ $X2=15.815 $Y2=1.252
r98 1 3 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=15.595 $Y=0.955
+ $X2=15.595 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_3466_403# 1 2 9 13 14 16 19 24 25 28 31
+ 32 34
c62 25 0 1.37034e-20 $X=18.095 $Y=1.35
r63 28 30 10.6287 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=17.5 $Y=0.445
+ $X2=17.5 $Y2=0.675
r64 25 35 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=18.122 $Y=1.35
+ $X2=18.122 $Y2=1.515
r65 25 34 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=18.122 $Y=1.35
+ $X2=18.122 $Y2=1.185
r66 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.095
+ $Y=1.35 $X2=18.095 $Y2=1.35
r67 22 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.675 $Y=1.35
+ $X2=17.59 $Y2=1.35
r68 22 24 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=17.675 $Y=1.35
+ $X2=18.095 $Y2=1.35
r69 20 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.59 $Y=1.515
+ $X2=17.59 $Y2=1.35
r70 20 31 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=17.59 $Y=1.515
+ $X2=17.59 $Y2=1.995
r71 19 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.59 $Y=1.185
+ $X2=17.59 $Y2=1.35
r72 19 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=17.59 $Y=1.185
+ $X2=17.59 $Y2=0.675
r73 14 31 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=17.532 $Y=2.137
+ $X2=17.532 $Y2=1.995
r74 14 16 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=17.532 $Y=2.137
+ $X2=17.532 $Y2=2.16
r75 13 34 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=18.24 $Y=0.655
+ $X2=18.24 $Y2=1.185
r76 9 35 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=18.235 $Y=2.465
+ $X2=18.235 $Y2=1.515
r77 2 16 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=17.33
+ $Y=2.015 $X2=17.475 $Y2=2.16
r78 1 28 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=17.36
+ $Y=0.235 $X2=17.49 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_27_481# 1 2 9 11 12 14 15 16 19
c54 9 0 6.37051e-20 $X=0.265 $Y=2.55
r55 17 19 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.065 $Y=2.905
+ $X2=2.065 $Y2=2.815
r56 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.94 $Y=2.99
+ $X2=2.065 $Y2=2.905
r57 15 16 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.94 $Y=2.99
+ $X2=1.19 $Y2=2.99
r58 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.105 $Y=2.905
+ $X2=1.19 $Y2=2.99
r59 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.105 $Y=2.215
+ $X2=1.105 $Y2=2.905
r60 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.02 $Y=2.13
+ $X2=1.105 $Y2=2.215
r61 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.02 $Y=2.13 $X2=0.43
+ $Y2=2.13
r62 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.265 $Y=2.215
+ $X2=0.43 $Y2=2.13
r63 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.265 $Y=2.215
+ $X2=0.265 $Y2=2.55
r64 2 19 600 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_PDIFF $count=1 $X=1.885
+ $Y=2.405 $X2=2.025 $Y2=2.815
r65 1 9 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.405 $X2=0.265 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%VPWR 1 2 3 4 5 18 22 26 30 36 43 44 45 47
+ 52 67 71 81 82 85 88 91 94
r162 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=3.33 $X2=18
+ $Y2=3.33
r163 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r164 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r165 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r166 82 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=18.48 $Y=3.33
+ $X2=18 $Y2=3.33
r167 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.48 $Y=3.33
+ $X2=18.48 $Y2=3.33
r168 79 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.185 $Y=3.33
+ $X2=18.02 $Y2=3.33
r169 79 81 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=18.185 $Y=3.33
+ $X2=18.48 $Y2=3.33
r170 78 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=3.33
+ $X2=18 $Y2=3.33
r171 77 78 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=17.52
+ $Y=3.33 $X2=17.52 $Y2=3.33
r172 75 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r173 74 77 626.31 $w=1.68e-07 $l=9.6e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=17.52 $Y2=3.33
r174 74 75 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=7.92
+ $Y=3.33 $X2=7.92 $Y2=3.33
r175 72 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.58 $Y=3.33
+ $X2=7.415 $Y2=3.33
r176 72 74 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.58 $Y=3.33
+ $X2=7.92 $Y2=3.33
r177 71 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.855 $Y=3.33
+ $X2=18.02 $Y2=3.33
r178 71 77 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=17.855 $Y=3.33
+ $X2=17.52 $Y2=3.33
r179 70 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r180 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r181 67 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.25 $Y=3.33
+ $X2=7.415 $Y2=3.33
r182 67 69 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.25 $Y=3.33
+ $X2=6.96 $Y2=3.33
r183 66 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r184 65 66 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r185 63 66 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r186 63 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r187 62 65 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r188 62 63 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r189 60 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=3.33
+ $X2=3.085 $Y2=3.33
r190 60 62 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=3.33
+ $X2=3.6 $Y2=3.33
r191 59 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r192 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r193 56 59 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r194 56 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 55 58 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r196 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r197 53 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.85 $Y=3.33
+ $X2=0.725 $Y2=3.33
r198 53 55 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.85 $Y=3.33
+ $X2=1.2 $Y2=3.33
r199 52 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=3.33
+ $X2=3.085 $Y2=3.33
r200 52 58 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r201 50 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r202 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r203 47 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.725 $Y2=3.33
r204 47 49 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.24 $Y2=3.33
r205 45 78 2.27448 $w=4.9e-07 $l=8.16e-06 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=17.52 $Y2=3.33
r206 45 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=7.92 $Y2=3.33
r207 43 65 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=6.025 $Y=3.33 $X2=6
+ $Y2=3.33
r208 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.025 $Y=3.33
+ $X2=6.19 $Y2=3.33
r209 42 69 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.355 $Y=3.33
+ $X2=6.96 $Y2=3.33
r210 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.355 $Y=3.33
+ $X2=6.19 $Y2=3.33
r211 39 41 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=18.02 $Y=2.465
+ $X2=18.02 $Y2=2.95
r212 36 39 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=18.02 $Y=1.98
+ $X2=18.02 $Y2=2.465
r213 34 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.02 $Y=3.245
+ $X2=18.02 $Y2=3.33
r214 34 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=18.02 $Y=3.245
+ $X2=18.02 $Y2=2.95
r215 30 33 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.415 $Y=2.42
+ $X2=7.415 $Y2=2.95
r216 28 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=3.245
+ $X2=7.415 $Y2=3.33
r217 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.415 $Y=3.245
+ $X2=7.415 $Y2=2.95
r218 24 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=3.245
+ $X2=6.19 $Y2=3.33
r219 24 26 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.19 $Y=3.245
+ $X2=6.19 $Y2=2.885
r220 20 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=3.245
+ $X2=3.085 $Y2=3.33
r221 20 22 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=3.085 $Y=3.245
+ $X2=3.085 $Y2=2.73
r222 16 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r223 16 18 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.55
r224 5 41 600 $w=1.7e-07 $l=1.05482e-06 $layer=licon1_PDIFF $count=1 $X=17.765
+ $Y=2.015 $X2=18.02 $Y2=2.95
r225 5 39 600 $w=1.7e-07 $l=5.6325e-07 $layer=licon1_PDIFF $count=1 $X=17.765
+ $Y=2.015 $X2=18.02 $Y2=2.465
r226 5 36 600 $w=1.7e-07 $l=2.71937e-07 $layer=licon1_PDIFF $count=1 $X=17.765
+ $Y=2.015 $X2=18.02 $Y2=1.98
r227 4 33 600 $w=1.7e-07 $l=8.2318e-07 $layer=licon1_PDIFF $count=1 $X=7.135
+ $Y=2.255 $X2=7.415 $Y2=2.95
r228 4 30 600 $w=1.7e-07 $l=3.52987e-07 $layer=licon1_PDIFF $count=1 $X=7.135
+ $Y=2.255 $X2=7.415 $Y2=2.42
r229 3 26 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.05
+ $Y=2.675 $X2=6.19 $Y2=2.885
r230 2 22 600 $w=1.7e-07 $l=1.04815e-06 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.795 $X2=3.085 $Y2=2.73
r231 1 18 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=2.405 $X2=0.765 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_189_119# 1 2 3 4 13 17 20 21 22 25 27
+ 28 30 32 36 37
c115 25 0 4.32663e-20 $X=4.145 $Y=0.945
c116 17 0 9.92106e-20 $X=3.665 $Y=2.31
c117 13 0 2.10137e-20 $X=1.6 $Y=0.95
r118 36 39 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=1.6 $Y=2.31 $X2=1.6
+ $Y2=2.6
r119 36 37 5.76029 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=2.31 $X2=1.6
+ $Y2=2.225
r120 32 34 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.085 $Y=0.805
+ $X2=1.085 $Y2=0.95
r121 30 43 12.4097 $w=3.49e-07 $l=4.47856e-07 $layer=LI1_cond $X=4.515 $Y=2.655
+ $X2=4.87 $Y2=2.865
r122 29 30 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=4.515 $Y=1.555
+ $X2=4.515 $Y2=2.655
r123 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.43 $Y=1.47
+ $X2=4.515 $Y2=1.555
r124 27 28 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.43 $Y=1.47 $X2=4.23
+ $Y2=1.47
r125 23 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.105 $Y=1.385
+ $X2=4.23 $Y2=1.47
r126 23 25 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=4.105 $Y=1.385
+ $X2=4.105 $Y2=0.945
r127 21 30 6.18747 $w=3.49e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.43 $Y=2.74
+ $X2=4.515 $Y2=2.655
r128 21 22 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.43 $Y=2.74
+ $X2=3.835 $Y2=2.74
r129 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.75 $Y=2.655
+ $X2=3.835 $Y2=2.74
r130 19 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.75 $Y=2.395
+ $X2=3.75 $Y2=2.655
r131 18 36 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.77 $Y=2.31 $X2=1.6
+ $Y2=2.31
r132 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.665 $Y=2.31
+ $X2=3.75 $Y2=2.395
r133 17 18 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=3.665 $Y=2.31
+ $X2=1.77 $Y2=2.31
r134 15 37 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=1.685 $Y=1.035
+ $X2=1.685 $Y2=2.225
r135 14 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=0.95
+ $X2=1.085 $Y2=0.95
r136 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=0.95
+ $X2=1.685 $Y2=1.035
r137 13 14 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.6 $Y=0.95
+ $X2=1.25 $Y2=0.95
r138 4 43 600 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=4.725
+ $Y=2.675 $X2=4.87 $Y2=2.865
r139 3 39 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.455
+ $Y=2.405 $X2=1.595 $Y2=2.6
r140 2 25 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=4
+ $Y=0.695 $X2=4.145 $Y2=0.945
r141 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.945
+ $Y=0.595 $X2=1.085 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1541_125# 1 2 9 13 17
c35 13 0 7.75523e-20 $X=8.27 $Y=2.4
r36 11 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.27 $Y=1.265
+ $X2=8.27 $Y2=1.18
r37 11 13 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=8.27 $Y=1.265
+ $X2=8.27 $Y2=2.4
r38 7 17 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.01 $Y=1.18 $X2=8.27
+ $Y2=1.18
r39 7 9 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.01 $Y=1.095
+ $X2=8.01 $Y2=0.76
r40 2 13 600 $w=1.7e-07 $l=6.33364e-07 $layer=licon1_PDIFF $count=1 $X=7.705
+ $Y=2.255 $X2=8.27 $Y2=2.4
r41 1 9 91 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_NDIFF $count=2 $X=7.705
+ $Y=0.625 $X2=7.99 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%KAPWR 1 2 3 10 14 17 18 23
c135 18 0 2.08416e-20 $X=16.08 $Y=2.82
r136 23 27 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=15.07 $Y=2.82
+ $X2=15.07 $Y2=2.99
r137 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=2.82
+ $X2=15.12 $Y2=2.82
r138 18 24 0.52469 $w=2.7e-07 $l=9.6e-07 $layer=MET1_cond $X=16.08 $Y=2.81
+ $X2=15.12 $Y2=2.81
r139 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=2.82
+ $X2=16.08 $Y2=2.82
r140 14 24 3.14814 $w=2.7e-07 $l=5.76e-06 $layer=MET1_cond $X=9.36 $Y=2.81
+ $X2=15.12 $Y2=2.81
r141 10 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.905 $Y=2.99
+ $X2=15.07 $Y2=2.99
r142 10 12 136.027 $w=1.68e-07 $l=2.085e-06 $layer=LI1_cond $X=14.905 $Y=2.99
+ $X2=12.82 $Y2=2.99
r143 3 17 600 $w=1.7e-07 $l=9.5687e-07 $layer=licon1_PDIFF $count=1 $X=15.89
+ $Y=1.92 $X2=16.14 $Y2=2.76
r144 2 23 600 $w=1.7e-07 $l=9.07097e-07 $layer=licon1_PDIFF $count=1 $X=14.83
+ $Y=2.07 $X2=15.07 $Y2=2.865
r145 1 12 600 $w=1.7e-07 $l=1.08946e-06 $layer=licon1_PDIFF $count=1 $X=12.6
+ $Y=2.005 $X2=12.82 $Y2=2.99
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%Q 1 2 7 8 9 10 11 12 13 22
r14 13 40 6.10117 $w=2.53e-07 $l=1.35e-07 $layer=LI1_cond $X=18.492 $Y=2.775
+ $X2=18.492 $Y2=2.91
r15 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=18.492 $Y=2.405
+ $X2=18.492 $Y2=2.775
r16 11 12 19.2074 $w=2.53e-07 $l=4.25e-07 $layer=LI1_cond $X=18.492 $Y=1.98
+ $X2=18.492 $Y2=2.405
r17 10 11 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=18.492 $Y=1.665
+ $X2=18.492 $Y2=1.98
r18 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=18.492 $Y=1.295
+ $X2=18.492 $Y2=1.665
r19 8 9 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=18.492 $Y=0.925
+ $X2=18.492 $Y2=1.295
r20 7 8 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=18.492 $Y=0.555
+ $X2=18.492 $Y2=0.925
r21 7 22 6.10117 $w=2.53e-07 $l=1.35e-07 $layer=LI1_cond $X=18.492 $Y=0.555
+ $X2=18.492 $Y2=0.42
r22 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=18.31
+ $Y=1.835 $X2=18.45 $Y2=2.91
r23 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=18.31
+ $Y=1.835 $X2=18.45 $Y2=1.98
r24 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=18.315
+ $Y=0.235 $X2=18.455 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46
+ 50 52 56 60 64 69 70 72 73 75 76 77 86 90 102 113 122 123 129 132 135 138 141
c182 123 0 1.14697e-20 $X=18.48 $Y=0
c183 42 0 1.50811e-19 $X=5.63 $Y=0.4
r184 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=0 $X2=18
+ $Y2=0
r185 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r186 136 139 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r187 135 136 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r188 132 133 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r189 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r190 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r191 123 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=18.48 $Y=0
+ $X2=18 $Y2=0
r192 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.48 $Y=0
+ $X2=18.48 $Y2=0
r193 120 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.19 $Y=0
+ $X2=18.025 $Y2=0
r194 120 122 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=18.19 $Y=0
+ $X2=18.48 $Y2=0
r195 119 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=0
+ $X2=18 $Y2=0
r196 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r197 116 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=17.52 $Y2=0
r198 115 118 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=16.56 $Y=0
+ $X2=17.52 $Y2=0
r199 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r200 113 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.86 $Y=0
+ $X2=18.025 $Y2=0
r201 113 118 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=17.86 $Y=0
+ $X2=17.52 $Y2=0
r202 112 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=16.56 $Y2=0
r203 111 112 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r204 109 112 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=16.08 $Y2=0
r205 109 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r206 108 111 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=16.08 $Y2=0
r207 108 109 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r208 106 138 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.995 $Y=0
+ $X2=11.87 $Y2=0
r209 106 108 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.995 $Y=0
+ $X2=12.24 $Y2=0
r210 104 105 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r211 102 135 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.775 $Y=0
+ $X2=10.9 $Y2=0
r212 102 104 217.578 $w=1.68e-07 $l=3.335e-06 $layer=LI1_cond $X=10.775 $Y=0
+ $X2=7.44 $Y2=0
r213 101 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r214 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r215 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r216 98 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r217 97 100 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r218 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r219 95 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.795 $Y=0
+ $X2=5.63 $Y2=0
r220 95 97 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=6
+ $Y2=0
r221 94 133 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=5.52 $Y2=0
r222 94 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r223 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r224 91 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=0
+ $X2=3.085 $Y2=0
r225 91 93 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.6
+ $Y2=0
r226 90 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=5.63 $Y2=0
r227 90 93 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=3.6 $Y2=0
r228 89 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.12 $Y2=0
r229 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r230 86 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=0
+ $X2=3.085 $Y2=0
r231 86 88 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=2.64
+ $Y2=0
r232 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r233 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r234 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r235 82 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r236 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r237 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r238 79 126 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0
+ $X2=0.215 $Y2=0
r239 79 81 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r240 77 136 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r241 77 105 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=7.44 $Y2=0
r242 75 111 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=16.085 $Y=0
+ $X2=16.08 $Y2=0
r243 75 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.085 $Y=0
+ $X2=16.21 $Y2=0
r244 74 115 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=16.335 $Y=0
+ $X2=16.56 $Y2=0
r245 74 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.335 $Y=0
+ $X2=16.21 $Y2=0
r246 72 100 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.115 $Y=0
+ $X2=6.96 $Y2=0
r247 72 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.115 $Y=0 $X2=7.24
+ $Y2=0
r248 71 104 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.365 $Y=0
+ $X2=7.44 $Y2=0
r249 71 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.365 $Y=0 $X2=7.24
+ $Y2=0
r250 69 84 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.68
+ $Y2=0
r251 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.065
+ $Y2=0
r252 68 88 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.64
+ $Y2=0
r253 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.065
+ $Y2=0
r254 64 66 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=18.025 $Y=0.38
+ $X2=18.025 $Y2=0.85
r255 62 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.025 $Y=0.085
+ $X2=18.025 $Y2=0
r256 62 64 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=18.025 $Y=0.085
+ $X2=18.025 $Y2=0.38
r257 58 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.21 $Y=0.085
+ $X2=16.21 $Y2=0
r258 58 60 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=16.21 $Y=0.085
+ $X2=16.21 $Y2=0.525
r259 54 138 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.87 $Y=0.085
+ $X2=11.87 $Y2=0
r260 54 56 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=11.87 $Y=0.085
+ $X2=11.87 $Y2=0.765
r261 53 135 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.025 $Y=0
+ $X2=10.9 $Y2=0
r262 52 138 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.745 $Y=0
+ $X2=11.87 $Y2=0
r263 52 53 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=11.745 $Y=0
+ $X2=11.025 $Y2=0
r264 48 135 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.9 $Y=0.085
+ $X2=10.9 $Y2=0
r265 48 50 33.8818 $w=2.48e-07 $l=7.35e-07 $layer=LI1_cond $X=10.9 $Y=0.085
+ $X2=10.9 $Y2=0.82
r266 44 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0
r267 44 46 28.8111 $w=2.48e-07 $l=6.25e-07 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0.71
r268 40 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.63 $Y=0.085
+ $X2=5.63 $Y2=0
r269 40 42 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.63 $Y=0.085
+ $X2=5.63 $Y2=0.4
r270 36 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.085
+ $X2=3.085 $Y2=0
r271 36 38 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=3.085 $Y=0.085
+ $X2=3.085 $Y2=0.84
r272 32 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.085
+ $X2=2.065 $Y2=0
r273 32 34 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=2.065 $Y=0.085
+ $X2=2.065 $Y2=0.805
r274 28 126 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.215 $Y2=0
r275 28 30 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.805
r276 9 66 182 $w=1.7e-07 $l=7.27255e-07 $layer=licon1_NDIFF $count=1 $X=17.78
+ $Y=0.235 $X2=18.025 $Y2=0.85
r277 9 64 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=17.78
+ $Y=0.235 $X2=18.025 $Y2=0.38
r278 8 60 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=16.03
+ $Y=0.36 $X2=16.17 $Y2=0.525
r279 7 56 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=11.775
+ $Y=0.595 $X2=11.91 $Y2=0.765
r280 6 50 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=10.8
+ $Y=0.625 $X2=10.94 $Y2=0.82
r281 5 46 182 $w=1.7e-07 $l=3.11047e-07 $layer=licon1_NDIFF $count=1 $X=7.075
+ $Y=0.485 $X2=7.28 $Y2=0.71
r282 4 42 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.49
+ $Y=0.235 $X2=5.63 $Y2=0.4
r283 3 38 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.695 $X2=3.085 $Y2=0.84
r284 2 34 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.595 $X2=2.025 $Y2=0.805
r285 1 30 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.595 $X2=0.265 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_2074_125# 1 2 9 11 12 15
c34 15 0 1.0685e-19 $X=11.37 $Y=0.835
r35 13 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=11.33 $Y=1.205
+ $X2=11.33 $Y2=0.835
r36 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.205 $Y=1.29
+ $X2=11.33 $Y2=1.205
r37 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.205 $Y=1.29
+ $X2=10.595 $Y2=1.29
r38 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.51 $Y=1.205
+ $X2=10.595 $Y2=1.29
r39 7 9 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.51 $Y=1.205
+ $X2=10.51 $Y2=0.835
r40 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.23
+ $Y=0.625 $X2=11.37 $Y2=0.835
r41 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.37
+ $Y=0.625 $X2=10.51 $Y2=0.835
.ends

