* File: sky130_fd_sc_lp__o2bb2ai_m.pex.spice
* Created: Fri Aug 28 11:13:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2AI_M%A1_N 3 7 9 10 11 12 13 20 21 24
c33 24 0 7.35046e-20 $X=0.255 $Y=1.055
c34 21 0 1.46887e-20 $X=0.27 $Y=1.12
r35 21 24 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=0.255 $Y=1.12
+ $X2=0.255 $Y2=1.055
r36 20 23 87.4515 $w=4.75e-07 $l=5.05e-07 $layer=POLY_cond $X=0.342 $Y=1.12
+ $X2=0.342 $Y2=1.625
r37 20 22 47.6426 $w=4.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.342 $Y=1.12
+ $X2=0.342 $Y2=0.955
r38 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r39 12 13 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r40 11 12 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r41 10 11 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r42 10 21 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.12
r43 9 24 8.04083 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=0.255 $Y=0.925 $X2=0.255
+ $Y2=1.055
r44 7 22 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.505 $Y=0.615
+ $X2=0.505 $Y2=0.955
r45 3 23 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=0.475 $Y=2.885
+ $X2=0.475 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_M%A2_N 3 6 9 10 11 12 13 14 20
c46 20 0 7.35046e-20 $X=0.955 $Y=1.1
c47 10 0 1.12137e-19 $X=0.955 $Y=1.44
r48 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=1.1 $X2=0.955 $Y2=1.1
r49 13 14 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.837 $Y=1.665
+ $X2=0.837 $Y2=2.035
r50 12 13 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.837 $Y=1.295
+ $X2=0.837 $Y2=1.665
r51 12 21 5.5488 $w=4.03e-07 $l=1.95e-07 $layer=LI1_cond $X=0.837 $Y=1.295
+ $X2=0.837 $Y2=1.1
r52 11 21 4.97969 $w=4.03e-07 $l=1.75e-07 $layer=LI1_cond $X=0.837 $Y=0.925
+ $X2=0.837 $Y2=1.1
r53 10 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.955 $Y=1.44
+ $X2=0.955 $Y2=1.1
r54 9 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=0.935
+ $X2=0.955 $Y2=1.1
r55 4 10 58.8488 $w=2.58e-07 $l=3.3908e-07 $layer=POLY_cond $X=0.905 $Y=1.755
+ $X2=0.955 $Y2=1.44
r56 4 6 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=0.905 $Y=1.755
+ $X2=0.905 $Y2=2.885
r57 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.865 $Y=0.615
+ $X2=0.865 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_M%A_110_535# 1 2 11 13 14 15 17 19 20 21 24
+ 26 27 28 35 36
c71 26 0 2.52635e-19 $X=1.27 $Y=2.43
r72 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.355
+ $Y=2.01 $X2=1.355 $Y2=2.01
r73 33 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.355 $Y=2.345
+ $X2=1.355 $Y2=2.01
r74 32 35 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=1.355 $Y=0.66
+ $X2=1.355 $Y2=2.01
r75 28 32 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.27 $Y=0.555
+ $X2=1.355 $Y2=0.66
r76 28 30 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=1.27 $Y=0.555
+ $X2=1.08 $Y2=0.555
r77 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.27 $Y=2.43
+ $X2=1.355 $Y2=2.345
r78 26 27 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.27 $Y=2.43
+ $X2=0.795 $Y2=2.43
r79 22 27 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.7 $Y=2.515
+ $X2=0.795 $Y2=2.43
r80 22 24 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=0.7 $Y=2.515
+ $X2=0.7 $Y2=2.82
r81 20 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.355 $Y=2.35
+ $X2=1.355 $Y2=2.01
r82 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=2.35
+ $X2=1.355 $Y2=2.515
r83 19 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.845
+ $X2=1.355 $Y2=2.01
r84 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.975 $Y=0.92
+ $X2=1.975 $Y2=0.6
r85 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.975 $Y2=0.92
r86 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.52 $Y2=0.995
r87 11 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.445 $Y=2.885
+ $X2=1.445 $Y2=2.515
r88 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.445 $Y=1.07
+ $X2=1.52 $Y2=0.995
r89 7 19 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=1.445 $Y=1.07
+ $X2=1.445 $Y2=1.845
r90 2 24 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.675 $X2=0.69 $Y2=2.82
r91 1 30 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.405 $X2=1.08 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_M%B2 3 7 9 10 11 20
c41 3 0 1.55187e-19 $X=1.875 $Y=2.885
r42 18 20 19.5645 $w=6.7e-07 $l=2.45e-07 $layer=POLY_cond $X=2.16 $Y=1.645
+ $X2=2.405 $Y2=1.645
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.16
+ $Y=1.475 $X2=2.16 $Y2=1.475
r44 15 18 22.7587 $w=6.7e-07 $l=2.85e-07 $layer=POLY_cond $X=1.875 $Y=1.645
+ $X2=2.16 $Y2=1.645
r45 10 11 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=2.035
r46 10 19 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.475
r47 9 19 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.475
r48 5 20 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.405 $Y=1.31
+ $X2=2.405 $Y2=1.645
r49 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.405 $Y=1.31
+ $X2=2.405 $Y2=0.6
r50 1 15 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.875 $Y=1.98
+ $X2=1.875 $Y2=1.645
r51 1 3 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.875 $Y=1.98
+ $X2=1.875 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_M%B1 3 5 6 9 13 14 15 16 17 23
r36 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.925
+ $Y=1.765 $X2=2.925 $Y2=1.765
r37 16 17 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.022 $Y=2.035
+ $X2=3.022 $Y2=2.405
r38 16 24 8.52492 $w=3.63e-07 $l=2.7e-07 $layer=LI1_cond $X=3.022 $Y=2.035
+ $X2=3.022 $Y2=1.765
r39 15 24 3.15738 $w=3.63e-07 $l=1e-07 $layer=LI1_cond $X=3.022 $Y=1.665
+ $X2=3.022 $Y2=1.765
r40 14 15 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.022 $Y=1.295
+ $X2=3.022 $Y2=1.665
r41 13 23 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=2.925 $Y=2.22
+ $X2=2.925 $Y2=1.765
r42 12 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.925 $Y=1.6
+ $X2=2.925 $Y2=1.765
r43 9 12 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=2.835 $Y=0.6 $X2=2.835
+ $Y2=1.6
r44 5 13 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.76 $Y=2.295
+ $X2=2.925 $Y2=2.22
r45 5 6 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.76 $Y=2.295 $X2=2.31
+ $Y2=2.295
r46 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.235 $Y=2.37
+ $X2=2.31 $Y2=2.295
r47 1 3 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.235 $Y=2.37
+ $X2=2.235 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_M%VPWR 1 2 3 10 12 16 20 23 24 25 27 37 38
+ 44
r46 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.14 $Y2=3.33
r52 32 34 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 28 41 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r57 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.14 $Y2=3.33
r59 27 30 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 25 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 23 34 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.45 $Y2=3.33
r64 22 37 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=3.12 $Y2=3.33
r65 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=2.45 $Y2=3.33
r66 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=3.245
+ $X2=2.45 $Y2=3.33
r67 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.45 $Y=3.245
+ $X2=2.45 $Y2=2.95
r68 14 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r69 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.95
r70 10 41 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r71 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r72 3 20 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=2.675 $X2=2.45 $Y2=2.95
r73 2 16 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.675 $X2=1.14 $Y2=2.95
r74 1 12 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.675 $X2=0.26 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_M%Y 1 2 9 12 16 19 20
r44 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=2.405
+ $X2=2.16 $Y2=2.405
r45 18 19 1.74598 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.865 $Y=2.405
+ $X2=1.76 $Y2=2.405
r46 14 16 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.66 $Y=2.82 $X2=1.74
+ $Y2=2.82
r47 12 16 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.74 $Y=2.715
+ $X2=1.74 $Y2=2.82
r48 11 19 4.70473 $w=1.9e-07 $l=9.44722e-08 $layer=LI1_cond $X=1.74 $Y=2.49
+ $X2=1.76 $Y2=2.405
r49 11 12 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.74 $Y=2.49
+ $X2=1.74 $Y2=2.715
r50 7 19 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=2.32 $X2=1.76
+ $Y2=2.405
r51 7 9 87.4069 $w=2.08e-07 $l=1.655e-06 $layer=LI1_cond $X=1.76 $Y=2.32
+ $X2=1.76 $Y2=0.665
r52 2 14 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=2.675 $X2=1.66 $Y2=2.82
r53 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.635
+ $Y=0.39 $X2=1.76 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_M%VGND 1 2 7 9 13 15 17 27 28 34
r36 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r37 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r38 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r39 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 25 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.62
+ $Y2=0
r41 25 27 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=3.12
+ $Y2=0
r42 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r43 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r45 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r46 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 18 31 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r48 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r49 17 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.515 $Y=0 $X2=2.62
+ $Y2=0
r50 17 23 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.515 $Y=0 $X2=2.16
+ $Y2=0
r51 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r52 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r53 11 34 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=0.085
+ $X2=2.62 $Y2=0
r54 11 13 22.71 $w=2.08e-07 $l=4.3e-07 $layer=LI1_cond $X=2.62 $Y=0.085 $X2=2.62
+ $Y2=0.515
r55 7 31 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.227 $Y2=0
r56 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.29 $Y=0.085 $X2=0.29
+ $Y2=0.55
r57 2 13 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.39 $X2=2.62 $Y2=0.515
r58 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.405 $X2=0.29 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_M%A_410_78# 1 2 9 11 12 15
r23 13 15 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=3.05 $Y=0.86
+ $X2=3.05 $Y2=0.665
r24 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.945 $Y=0.945
+ $X2=3.05 $Y2=0.86
r25 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.945 $Y=0.945
+ $X2=2.295 $Y2=0.945
r26 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.19 $Y=0.86
+ $X2=2.295 $Y2=0.945
r27 7 9 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=2.19 $Y=0.86 $X2=2.19
+ $Y2=0.685
r28 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.91
+ $Y=0.39 $X2=3.05 $Y2=0.665
r29 1 9 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.05
+ $Y=0.39 $X2=2.19 $Y2=0.685
.ends

