* File: sky130_fd_sc_lp__dfstp_lp.pxi.spice
* Created: Wed Sep  2 09:44:41 2020
* 
x_PM_SKY130_FD_SC_LP__DFSTP_LP%D N_D_c_270_n N_D_M1022_g N_D_M1005_g N_D_c_271_n
+ N_D_M1010_g N_D_c_272_n D D N_D_c_273_n N_D_c_274_n N_D_c_275_n
+ PM_SKY130_FD_SC_LP__DFSTP_LP%D
x_PM_SKY130_FD_SC_LP__DFSTP_LP%CLK N_CLK_M1029_g N_CLK_c_305_n N_CLK_M1023_g
+ N_CLK_c_306_n N_CLK_c_307_n N_CLK_M1013_g N_CLK_c_308_n CLK N_CLK_c_310_n
+ N_CLK_c_311_n PM_SKY130_FD_SC_LP__DFSTP_LP%CLK
x_PM_SKY130_FD_SC_LP__DFSTP_LP%A_479_409# N_A_479_409#_M1011_d
+ N_A_479_409#_M1018_d N_A_479_409#_M1021_g N_A_479_409#_c_362_n
+ N_A_479_409#_M1017_g N_A_479_409#_M1030_g N_A_479_409#_M1024_g
+ N_A_479_409#_c_376_n N_A_479_409#_c_377_n N_A_479_409#_c_378_n
+ N_A_479_409#_c_379_n N_A_479_409#_c_365_n N_A_479_409#_c_390_p
+ N_A_479_409#_c_391_p N_A_479_409#_c_392_p N_A_479_409#_c_393_p
+ N_A_479_409#_c_394_p N_A_479_409#_c_389_p N_A_479_409#_c_414_p
+ N_A_479_409#_c_401_p N_A_479_409#_c_380_n N_A_479_409#_c_381_n
+ N_A_479_409#_c_366_n N_A_479_409#_c_383_n N_A_479_409#_c_367_n
+ N_A_479_409#_c_368_n N_A_479_409#_c_369_n N_A_479_409#_c_370_n
+ N_A_479_409#_c_371_n N_A_479_409#_c_372_n N_A_479_409#_c_410_p
+ N_A_479_409#_c_373_n PM_SKY130_FD_SC_LP__DFSTP_LP%A_479_409#
x_PM_SKY130_FD_SC_LP__DFSTP_LP%A_943_321# N_A_943_321#_M1019_s
+ N_A_943_321#_M1012_d N_A_943_321#_M1027_g N_A_943_321#_M1008_g
+ N_A_943_321#_c_596_n N_A_943_321#_c_597_n N_A_943_321#_c_598_n
+ N_A_943_321#_c_599_n N_A_943_321#_c_605_n N_A_943_321#_c_620_n
+ N_A_943_321#_c_600_n N_A_943_321#_c_621_n N_A_943_321#_c_601_n
+ PM_SKY130_FD_SC_LP__DFSTP_LP%A_943_321#
x_PM_SKY130_FD_SC_LP__DFSTP_LP%A_709_419# N_A_709_419#_M1028_d
+ N_A_709_419#_M1021_d N_A_709_419#_M1012_g N_A_709_419#_c_685_n
+ N_A_709_419#_c_686_n N_A_709_419#_c_687_n N_A_709_419#_M1019_g
+ N_A_709_419#_M1031_g N_A_709_419#_M1002_g N_A_709_419#_c_689_n
+ N_A_709_419#_c_709_n N_A_709_419#_c_730_n N_A_709_419#_c_710_n
+ N_A_709_419#_c_711_n N_A_709_419#_c_690_n N_A_709_419#_c_691_n
+ N_A_709_419#_c_692_n N_A_709_419#_c_693_n N_A_709_419#_c_694_n
+ N_A_709_419#_c_695_n N_A_709_419#_c_696_n N_A_709_419#_c_697_n
+ N_A_709_419#_c_698_n N_A_709_419#_c_699_n N_A_709_419#_c_700_n
+ N_A_709_419#_c_792_n N_A_709_419#_c_701_n N_A_709_419#_c_702_n
+ N_A_709_419#_c_703_n N_A_709_419#_c_704_n N_A_709_419#_c_705_n
+ PM_SKY130_FD_SC_LP__DFSTP_LP%A_709_419#
x_PM_SKY130_FD_SC_LP__DFSTP_LP%SET_B N_SET_B_M1025_g N_SET_B_M1007_g
+ N_SET_B_c_884_n N_SET_B_M1036_g N_SET_B_c_885_n N_SET_B_c_886_n
+ N_SET_B_M1033_g N_SET_B_c_887_n N_SET_B_c_888_n N_SET_B_c_889_n SET_B
+ N_SET_B_c_891_n N_SET_B_c_892_n N_SET_B_c_893_n N_SET_B_c_894_n
+ PM_SKY130_FD_SC_LP__DFSTP_LP%SET_B
x_PM_SKY130_FD_SC_LP__DFSTP_LP%A_266_409# N_A_266_409#_M1023_s
+ N_A_266_409#_M1029_s N_A_266_409#_M1018_g N_A_266_409#_M1014_g
+ N_A_266_409#_c_1015_n N_A_266_409#_c_1016_n N_A_266_409#_M1011_g
+ N_A_266_409#_c_1018_n N_A_266_409#_c_1019_n N_A_266_409#_M1028_g
+ N_A_266_409#_c_1036_n N_A_266_409#_c_1037_n N_A_266_409#_c_1021_n
+ N_A_266_409#_c_1022_n N_A_266_409#_M1026_g N_A_266_409#_c_1039_n
+ N_A_266_409#_M1009_g N_A_266_409#_c_1040_n N_A_266_409#_c_1041_n
+ N_A_266_409#_c_1023_n N_A_266_409#_M1032_g N_A_266_409#_c_1025_n
+ N_A_266_409#_c_1026_n N_A_266_409#_c_1027_n N_A_266_409#_c_1028_n
+ N_A_266_409#_c_1029_n N_A_266_409#_c_1044_n N_A_266_409#_c_1030_n
+ N_A_266_409#_c_1031_n N_A_266_409#_c_1045_n N_A_266_409#_c_1046_n
+ N_A_266_409#_c_1032_n N_A_266_409#_c_1033_n
+ PM_SKY130_FD_SC_LP__DFSTP_LP%A_266_409#
x_PM_SKY130_FD_SC_LP__DFSTP_LP%A_1731_99# N_A_1731_99#_M1035_s
+ N_A_1731_99#_M1034_s N_A_1731_99#_c_1221_n N_A_1731_99#_M1020_g
+ N_A_1731_99#_c_1222_n N_A_1731_99#_M1000_g N_A_1731_99#_c_1223_n
+ N_A_1731_99#_c_1224_n N_A_1731_99#_c_1225_n N_A_1731_99#_c_1226_n
+ N_A_1731_99#_c_1227_n N_A_1731_99#_c_1228_n N_A_1731_99#_c_1234_n
+ N_A_1731_99#_c_1235_n N_A_1731_99#_c_1229_n N_A_1731_99#_c_1230_n
+ PM_SKY130_FD_SC_LP__DFSTP_LP%A_1731_99#
x_PM_SKY130_FD_SC_LP__DFSTP_LP%A_1526_125# N_A_1526_125#_M1030_d
+ N_A_1526_125#_M1009_d N_A_1526_125#_M1033_d N_A_1526_125#_c_1316_n
+ N_A_1526_125#_M1035_g N_A_1526_125#_c_1317_n N_A_1526_125#_c_1318_n
+ N_A_1526_125#_c_1319_n N_A_1526_125#_M1037_g N_A_1526_125#_M1034_g
+ N_A_1526_125#_c_1321_n N_A_1526_125#_M1001_g N_A_1526_125#_c_1323_n
+ N_A_1526_125#_M1016_g N_A_1526_125#_M1003_g N_A_1526_125#_c_1326_n
+ N_A_1526_125#_c_1327_n N_A_1526_125#_c_1328_n N_A_1526_125#_c_1329_n
+ N_A_1526_125#_c_1379_n N_A_1526_125#_c_1330_n N_A_1526_125#_c_1339_n
+ N_A_1526_125#_c_1340_n N_A_1526_125#_c_1331_n N_A_1526_125#_c_1342_n
+ N_A_1526_125#_c_1343_n N_A_1526_125#_c_1344_n N_A_1526_125#_c_1345_n
+ N_A_1526_125#_c_1332_n N_A_1526_125#_c_1333_n N_A_1526_125#_c_1334_n
+ N_A_1526_125#_c_1335_n N_A_1526_125#_c_1336_n N_A_1526_125#_c_1418_n
+ PM_SKY130_FD_SC_LP__DFSTP_LP%A_1526_125#
x_PM_SKY130_FD_SC_LP__DFSTP_LP%A_2287_74# N_A_2287_74#_M1001_s
+ N_A_2287_74#_M1016_s N_A_2287_74#_M1015_g N_A_2287_74#_M1004_g
+ N_A_2287_74#_M1006_g N_A_2287_74#_c_1498_n N_A_2287_74#_c_1499_n
+ N_A_2287_74#_c_1500_n N_A_2287_74#_c_1508_n N_A_2287_74#_c_1501_n
+ N_A_2287_74#_c_1502_n N_A_2287_74#_c_1503_n N_A_2287_74#_c_1504_n
+ N_A_2287_74#_c_1505_n PM_SKY130_FD_SC_LP__DFSTP_LP%A_2287_74#
x_PM_SKY130_FD_SC_LP__DFSTP_LP%VPWR N_VPWR_M1005_s N_VPWR_M1029_d N_VPWR_M1027_d
+ N_VPWR_M1025_d N_VPWR_M1000_d N_VPWR_M1034_d N_VPWR_M1016_d N_VPWR_c_1569_n
+ N_VPWR_c_1570_n N_VPWR_c_1571_n N_VPWR_c_1572_n N_VPWR_c_1573_n
+ N_VPWR_c_1574_n N_VPWR_c_1575_n N_VPWR_c_1576_n N_VPWR_c_1577_n
+ N_VPWR_c_1578_n VPWR N_VPWR_c_1579_n N_VPWR_c_1580_n N_VPWR_c_1581_n
+ N_VPWR_c_1582_n N_VPWR_c_1583_n N_VPWR_c_1584_n N_VPWR_c_1568_n
+ N_VPWR_c_1586_n N_VPWR_c_1587_n N_VPWR_c_1588_n N_VPWR_c_1589_n
+ N_VPWR_c_1590_n PM_SKY130_FD_SC_LP__DFSTP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DFSTP_LP%A_135_409# N_A_135_409#_M1010_d
+ N_A_135_409#_M1028_s N_A_135_409#_M1005_d N_A_135_409#_M1021_s
+ N_A_135_409#_c_1723_n N_A_135_409#_c_1724_n N_A_135_409#_c_1713_n
+ N_A_135_409#_c_1714_n N_A_135_409#_c_1715_n N_A_135_409#_c_1716_n
+ N_A_135_409#_c_1717_n N_A_135_409#_c_1718_n N_A_135_409#_c_1719_n
+ N_A_135_409#_c_1720_n N_A_135_409#_c_1721_n N_A_135_409#_c_1722_n
+ N_A_135_409#_c_1727_n PM_SKY130_FD_SC_LP__DFSTP_LP%A_135_409#
x_PM_SKY130_FD_SC_LP__DFSTP_LP%Q N_Q_M1006_d N_Q_M1004_d Q Q Q Q Q Q Q
+ N_Q_c_1833_n Q PM_SKY130_FD_SC_LP__DFSTP_LP%Q
x_PM_SKY130_FD_SC_LP__DFSTP_LP%VGND N_VGND_M1022_s N_VGND_M1013_d N_VGND_M1008_d
+ N_VGND_M1007_d N_VGND_M1036_d N_VGND_M1037_d N_VGND_M1003_d N_VGND_c_1851_n
+ N_VGND_c_1852_n N_VGND_c_1853_n N_VGND_c_1854_n N_VGND_c_1855_n
+ N_VGND_c_1856_n N_VGND_c_1857_n N_VGND_c_1858_n N_VGND_c_1859_n
+ N_VGND_c_1860_n N_VGND_c_1861_n N_VGND_c_1862_n N_VGND_c_1863_n
+ N_VGND_c_1864_n VGND N_VGND_c_1865_n N_VGND_c_1866_n N_VGND_c_1867_n
+ N_VGND_c_1868_n N_VGND_c_1869_n N_VGND_c_1870_n N_VGND_c_1871_n
+ N_VGND_c_1872_n PM_SKY130_FD_SC_LP__DFSTP_LP%VGND
cc_1 VNB N_D_c_270_n 0.0175093f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.78
cc_2 VNB N_D_c_271_n 0.0174572f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.78
cc_3 VNB N_D_c_272_n 0.0318739f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.855
cc_4 VNB N_D_c_273_n 0.0603619f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_5 VNB N_D_c_274_n 0.0245402f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_6 VNB N_D_c_275_n 0.018257f $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=1.11
cc_7 VNB N_CLK_c_305_n 0.0161086f $X=-0.19 $Y=-0.245 $X2=0.537 $Y2=1.11
cc_8 VNB N_CLK_c_306_n 0.0197939f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.78
cc_9 VNB N_CLK_c_307_n 0.0134887f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.495
cc_10 VNB N_CLK_c_308_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.537 $Y2=0.855
cc_11 VNB CLK 0.00192922f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.855
cc_12 VNB N_CLK_c_310_n 0.0232962f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_CLK_c_311_n 0.018541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_479_409#_c_362_n 0.0348793f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.495
cc_15 VNB N_A_479_409#_M1017_g 0.0191129f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.855
cc_16 VNB N_A_479_409#_M1030_g 0.0265043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_479_409#_c_365_n 0.0140184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_479_409#_c_366_n 0.0117847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_479_409#_c_367_n 0.00896682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_479_409#_c_368_n 0.0179994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_479_409#_c_369_n 0.00743971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_479_409#_c_370_n 0.00429533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_479_409#_c_371_n 0.00230273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_479_409#_c_372_n 0.0136821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_479_409#_c_373_n 0.0277522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_943_321#_M1008_g 0.0419565f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.855
cc_27 VNB N_A_943_321#_c_596_n 0.00408438f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_28 VNB N_A_943_321#_c_597_n 0.0207263f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_A_943_321#_c_598_n 0.0171159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_943_321#_c_599_n 0.00628966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_943_321#_c_600_n 0.00749004f $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=1.11
cc_32 VNB N_A_943_321#_c_601_n 0.00862753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_709_419#_c_685_n 0.0209773f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.855
cc_34 VNB N_A_709_419#_c_686_n 0.0107917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_709_419#_c_687_n 0.0151731f $X=-0.19 $Y=-0.245 $X2=0.537 $Y2=0.855
cc_36 VNB N_A_709_419#_M1002_g 0.0189946f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_37 VNB N_A_709_419#_c_689_n 0.0197009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_709_419#_c_690_n 0.00596276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_709_419#_c_691_n 0.00650994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_709_419#_c_692_n 0.00730002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_709_419#_c_693_n 0.0126521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_709_419#_c_694_n 0.0250768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_709_419#_c_695_n 0.00348498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_709_419#_c_696_n 0.0040819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_709_419#_c_697_n 0.00864449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_709_419#_c_698_n 0.00577427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_709_419#_c_699_n 0.00533661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_709_419#_c_700_n 0.00466721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_709_419#_c_701_n 0.00368221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_709_419#_c_702_n 0.0100876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_709_419#_c_703_n 0.00570695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_709_419#_c_704_n 0.0146511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_709_419#_c_705_n 0.0212375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_SET_B_M1007_g 0.0377722f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.545
cc_55 VNB N_SET_B_c_884_n 0.0191353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_SET_B_c_885_n 0.0415972f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.495
cc_57 VNB N_SET_B_c_886_n 0.0061284f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.855
cc_58 VNB N_SET_B_c_887_n 0.0122451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_SET_B_c_888_n 0.00133855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_SET_B_c_889_n 5.37117e-19 $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_61 VNB SET_B 3.82464e-19 $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=1.78
cc_62 VNB N_SET_B_c_891_n 0.0190914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_SET_B_c_892_n 0.0134682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_SET_B_c_893_n 0.0169693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_SET_B_c_894_n 0.00270858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_266_409#_M1014_g 0.0169747f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.855
cc_67 VNB N_A_266_409#_c_1015_n 0.0164042f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.855
cc_68 VNB N_A_266_409#_c_1016_n 0.00756955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_266_409#_M1011_g 0.01987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_266_409#_c_1018_n 0.045773f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_71 VNB N_A_266_409#_c_1019_n 0.0223979f $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=1.78
cc_72 VNB N_A_266_409#_M1028_g 0.0358023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_266_409#_c_1021_n 0.336215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_266_409#_c_1022_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_266_409#_c_1023_n 0.0211951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_266_409#_M1032_g 0.0333036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_266_409#_c_1025_n 0.00514703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_266_409#_c_1026_n 0.00787172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_266_409#_c_1027_n 0.00662267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_266_409#_c_1028_n 0.0257208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_266_409#_c_1029_n 0.00899408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_266_409#_c_1030_n 0.0163804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_266_409#_c_1031_n 0.00731112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_266_409#_c_1032_n 0.00466452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_266_409#_c_1033_n 0.0224281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1731_99#_c_1221_n 0.0165417f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.545
cc_87 VNB N_A_1731_99#_c_1222_n 0.015767f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.495
cc_88 VNB N_A_1731_99#_c_1223_n 0.0300288f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_89 VNB N_A_1731_99#_c_1224_n 0.0033103f $X=-0.19 $Y=-0.245 $X2=0.447
+ $Y2=1.275
cc_90 VNB N_A_1731_99#_c_1225_n 0.0244688f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.275
cc_91 VNB N_A_1731_99#_c_1226_n 0.00579723f $X=-0.19 $Y=-0.245 $X2=0.447
+ $Y2=1.11
cc_92 VNB N_A_1731_99#_c_1227_n 0.00608946f $X=-0.19 $Y=-0.245 $X2=0.447
+ $Y2=1.78
cc_93 VNB N_A_1731_99#_c_1228_n 0.0158382f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.295
cc_94 VNB N_A_1731_99#_c_1229_n 0.0223741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1731_99#_c_1230_n 0.00486511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1526_125#_c_1316_n 0.0172366f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.78
cc_97 VNB N_A_1526_125#_c_1317_n 0.011952f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=0.855
cc_98 VNB N_A_1526_125#_c_1318_n 0.0109035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1526_125#_c_1319_n 0.0164171f $X=-0.19 $Y=-0.245 $X2=0.537
+ $Y2=0.855
cc_100 VNB N_A_1526_125#_M1034_g 0.0014858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1526_125#_c_1321_n 0.0432915f $X=-0.19 $Y=-0.245 $X2=0.447
+ $Y2=1.275
cc_102 VNB N_A_1526_125#_M1001_g 0.0416085f $X=-0.19 $Y=-0.245 $X2=0.447
+ $Y2=1.78
cc_103 VNB N_A_1526_125#_c_1323_n 0.00703176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1526_125#_M1016_g 0.0103862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1526_125#_M1003_g 0.0377492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1526_125#_c_1326_n 0.0170703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1526_125#_c_1327_n 0.0158468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1526_125#_c_1328_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1526_125#_c_1329_n 0.00881558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1526_125#_c_1330_n 0.00252615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1526_125#_c_1331_n 0.00541581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1526_125#_c_1332_n 0.00256977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1526_125#_c_1333_n 0.0472192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1526_125#_c_1334_n 0.00138224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1526_125#_c_1335_n 3.0401e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_1526_125#_c_1336_n 0.00605326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2287_74#_M1015_g 0.0202817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2287_74#_M1006_g 0.0250727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2287_74#_c_1498_n 0.0255246f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.275
cc_120 VNB N_A_2287_74#_c_1499_n 0.0118058f $X=-0.19 $Y=-0.245 $X2=0.447
+ $Y2=1.78
cc_121 VNB N_A_2287_74#_c_1500_n 0.00638111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2287_74#_c_1501_n 0.00889996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2287_74#_c_1502_n 0.00121962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2287_74#_c_1503_n 0.0276345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2287_74#_c_1504_n 0.0137821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_2287_74#_c_1505_n 0.00207542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VPWR_c_1568_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_135_409#_c_1713_n 0.0185253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_135_409#_c_1714_n 0.00144245f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.275
cc_130 VNB N_A_135_409#_c_1715_n 0.00195831f $X=-0.19 $Y=-0.245 $X2=0.447
+ $Y2=1.78
cc_131 VNB N_A_135_409#_c_1716_n 0.0177005f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.275
cc_132 VNB N_A_135_409#_c_1717_n 0.00269587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_135_409#_c_1718_n 0.00646754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_135_409#_c_1719_n 0.00955637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_135_409#_c_1720_n 0.0185899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_135_409#_c_1721_n 0.0145896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_135_409#_c_1722_n 0.0207859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB Q 0.0227502f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.545
cc_139 VNB Q 0.0432458f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.545
cc_140 VNB N_VGND_c_1851_n 0.0107448f $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=1.275
cc_141 VNB N_VGND_c_1852_n 0.0265531f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_142 VNB N_VGND_c_1853_n 0.012609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1854_n 0.0121111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1855_n 0.0163391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_1856_n 0.0251415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_1857_n 0.00794941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_1858_n 0.0136149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_1859_n 0.046366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_1860_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_1861_n 0.074349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_1862_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_1863_n 0.0305495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_1864_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_1865_n 0.0650087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_1866_n 0.0355252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_1867_n 0.0287283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_1868_n 0.0282219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_1869_n 0.723146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_1870_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_1871_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_1872_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VPB N_D_M1005_g 0.0458742f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.545
cc_163 VPB N_D_c_273_n 0.018523f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_164 VPB N_D_c_274_n 0.00801329f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_165 VPB N_CLK_M1029_g 0.0365469f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.495
cc_166 VPB CLK 9.8164e-19 $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.855
cc_167 VPB N_CLK_c_310_n 0.0131643f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_168 VPB N_A_479_409#_M1021_g 0.037001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_479_409#_M1024_g 0.0330645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_479_409#_c_376_n 0.00170032f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.275
cc_171 VPB N_A_479_409#_c_377_n 0.00234077f $X=-0.19 $Y=1.655 $X2=0.447 $Y2=1.11
cc_172 VPB N_A_479_409#_c_378_n 0.0109902f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.275
cc_173 VPB N_A_479_409#_c_379_n 0.00268878f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_479_409#_c_380_n 0.0075389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_479_409#_c_381_n 5.89321e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_479_409#_c_366_n 0.0010328f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_479_409#_c_383_n 0.00286389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_479_409#_c_367_n 0.0040347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_479_409#_c_368_n 0.0131355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_479_409#_c_370_n 0.0048662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_479_409#_c_372_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_943_321#_M1027_g 0.0277269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_943_321#_c_596_n 0.00251332f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_184 VPB N_A_943_321#_c_597_n 0.0419454f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_185 VPB N_A_943_321#_c_605_n 0.0106408f $X=-0.19 $Y=1.655 $X2=0.447 $Y2=1.275
cc_186 VPB N_A_709_419#_M1012_g 0.0307296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_709_419#_M1031_g 0.0320945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_709_419#_c_689_n 0.00390768f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_709_419#_c_709_n 0.014958f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.295
cc_190 VPB N_A_709_419#_c_710_n 0.00722063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_709_419#_c_711_n 0.00291473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_709_419#_c_691_n 0.00820953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_709_419#_c_701_n 0.00678818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_709_419#_c_702_n 0.0164834f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_709_419#_c_703_n 7.708e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_SET_B_M1025_g 0.0327074f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.495
cc_197 VPB N_SET_B_M1033_g 0.0399421f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.855
cc_198 VPB N_SET_B_c_887_n 0.00637249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_SET_B_c_889_n 0.00132186f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_200 VPB SET_B 3.834e-19 $X=-0.19 $Y=1.655 $X2=0.447 $Y2=1.78
cc_201 VPB N_SET_B_c_891_n 0.0267627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_SET_B_c_892_n 0.0157164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_SET_B_c_894_n 0.00348378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_266_409#_M1018_g 0.0315132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_266_409#_c_1019_n 0.0127792f $X=-0.19 $Y=1.655 $X2=0.447 $Y2=1.78
cc_206 VPB N_A_266_409#_c_1036_n 0.0252071f $X=-0.19 $Y=1.655 $X2=0.337
+ $Y2=1.665
cc_207 VPB N_A_266_409#_c_1037_n 0.0108515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_266_409#_M1026_g 0.0264815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_266_409#_c_1039_n 0.0211314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_266_409#_c_1040_n 0.0312468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_266_409#_c_1041_n 0.00860929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_266_409#_c_1023_n 0.0117257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_266_409#_c_1029_n 0.00674045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_266_409#_c_1044_n 0.016164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_266_409#_c_1045_n 0.00529045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_266_409#_c_1046_n 0.0106801f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_266_409#_c_1032_n 0.00331644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_266_409#_c_1033_n 0.0261411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1731_99#_M1000_g 0.0330223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_1731_99#_c_1224_n 0.0029014f $X=-0.19 $Y=1.655 $X2=0.447
+ $Y2=1.275
cc_221 VPB N_A_1731_99#_c_1225_n 0.0249915f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.275
cc_222 VPB N_A_1731_99#_c_1234_n 0.00474459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_1731_99#_c_1235_n 0.0115467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_1731_99#_c_1230_n 0.00353855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1526_125#_M1034_g 0.0316198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_1526_125#_M1016_g 0.0316655f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_1526_125#_c_1339_n 0.00213964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_1526_125#_c_1340_n 0.00286131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_1526_125#_c_1331_n 0.00267854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_1526_125#_c_1342_n 0.0161866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_1526_125#_c_1343_n 0.00701759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_1526_125#_c_1344_n 0.0246699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_1526_125#_c_1345_n 2.73935e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_1526_125#_c_1335_n 0.00559419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_2287_74#_M1004_g 0.0327251f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.855
cc_236 VPB N_A_2287_74#_c_1499_n 0.00265205f $X=-0.19 $Y=1.655 $X2=0.447
+ $Y2=1.78
cc_237 VPB N_A_2287_74#_c_1508_n 0.017363f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.665
cc_238 VPB N_A_2287_74#_c_1501_n 0.00280416f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1569_n 0.0115163f $X=-0.19 $Y=1.655 $X2=0.447 $Y2=1.275
cc_240 VPB N_VPWR_c_1570_n 0.04683f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_241 VPB N_VPWR_c_1571_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1572_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1573_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1574_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1575_n 0.030435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1576_n 0.0137031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1577_n 0.0216338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1578_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1579_n 0.0352978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1580_n 0.0636302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1581_n 0.0345797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1582_n 0.0625976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1583_n 0.0462007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1584_n 0.0253236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1568_n 0.103797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1586_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1587_n 0.00510584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1588_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1589_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1590_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_135_409#_c_1723_n 0.00698308f $X=-0.19 $Y=1.655 $X2=0.537
+ $Y2=0.855
cc_262 VPB N_A_135_409#_c_1724_n 0.00979164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_135_409#_c_1718_n 0.0103168f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_135_409#_c_1720_n 0.00795625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_135_409#_c_1727_n 0.0203875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB Q 0.0107174f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.545
cc_267 VPB Q 0.0417159f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.495
cc_268 VPB N_Q_c_1833_n 0.0223739f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 N_D_M1005_g N_A_266_409#_c_1044_n 0.00157815f $X=0.55 $Y=2.545 $X2=0
+ $Y2=0
cc_270 N_D_c_271_n N_A_266_409#_c_1031_n 0.00139213f $X=0.835 $Y=0.78 $X2=0
+ $Y2=0
cc_271 N_D_M1005_g N_A_266_409#_c_1046_n 2.35528e-19 $X=0.55 $Y=2.545 $X2=0
+ $Y2=0
cc_272 N_D_M1005_g N_VPWR_c_1570_n 0.0250417f $X=0.55 $Y=2.545 $X2=0 $Y2=0
cc_273 N_D_c_273_n N_VPWR_c_1570_n 0.00153765f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_274 N_D_c_274_n N_VPWR_c_1570_n 0.0221768f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_275 N_D_M1005_g N_VPWR_c_1579_n 0.00769046f $X=0.55 $Y=2.545 $X2=0 $Y2=0
cc_276 N_D_M1005_g N_VPWR_c_1568_n 0.0143431f $X=0.55 $Y=2.545 $X2=0 $Y2=0
cc_277 N_D_M1005_g N_A_135_409#_c_1723_n 0.00451956f $X=0.55 $Y=2.545 $X2=0
+ $Y2=0
cc_278 N_D_M1005_g N_A_135_409#_c_1724_n 0.015872f $X=0.55 $Y=2.545 $X2=0 $Y2=0
cc_279 N_D_c_271_n N_A_135_409#_c_1720_n 0.00199302f $X=0.835 $Y=0.78 $X2=0
+ $Y2=0
cc_280 N_D_c_272_n N_A_135_409#_c_1720_n 0.0123703f $X=0.835 $Y=0.855 $X2=0
+ $Y2=0
cc_281 N_D_c_274_n N_A_135_409#_c_1720_n 0.0373518f $X=0.385 $Y=1.275 $X2=0
+ $Y2=0
cc_282 N_D_c_275_n N_A_135_409#_c_1720_n 0.0334991f $X=0.447 $Y=1.11 $X2=0 $Y2=0
cc_283 N_D_c_270_n N_A_135_409#_c_1721_n 0.00173006f $X=0.475 $Y=0.78 $X2=0
+ $Y2=0
cc_284 N_D_c_271_n N_A_135_409#_c_1721_n 0.0111648f $X=0.835 $Y=0.78 $X2=0 $Y2=0
cc_285 N_D_c_270_n N_VGND_c_1852_n 0.0136234f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_286 N_D_c_271_n N_VGND_c_1852_n 0.00205702f $X=0.835 $Y=0.78 $X2=0 $Y2=0
cc_287 N_D_c_273_n N_VGND_c_1852_n 0.0012686f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_288 N_D_c_274_n N_VGND_c_1852_n 0.014708f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_289 N_D_c_270_n N_VGND_c_1859_n 0.00445056f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_290 N_D_c_271_n N_VGND_c_1859_n 0.00398426f $X=0.835 $Y=0.78 $X2=0 $Y2=0
cc_291 N_D_c_272_n N_VGND_c_1859_n 5.84996e-19 $X=0.835 $Y=0.855 $X2=0 $Y2=0
cc_292 N_D_c_270_n N_VGND_c_1869_n 0.00796275f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_293 N_D_c_271_n N_VGND_c_1869_n 0.00752426f $X=0.835 $Y=0.78 $X2=0 $Y2=0
cc_294 N_D_c_272_n N_VGND_c_1869_n 7.94744e-19 $X=0.835 $Y=0.855 $X2=0 $Y2=0
cc_295 N_CLK_M1029_g N_A_479_409#_c_377_n 9.40572e-19 $X=1.74 $Y=2.545 $X2=0
+ $Y2=0
cc_296 N_CLK_M1029_g N_A_266_409#_M1018_g 0.0205055f $X=1.74 $Y=2.545 $X2=0
+ $Y2=0
cc_297 N_CLK_c_307_n N_A_266_409#_M1014_g 0.00815124f $X=2.15 $Y=1.04 $X2=0
+ $Y2=0
cc_298 CLK N_A_266_409#_c_1015_n 2.99945e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_299 N_CLK_c_310_n N_A_266_409#_c_1015_n 0.0028093f $X=1.675 $Y=1.615 $X2=0
+ $Y2=0
cc_300 N_CLK_c_306_n N_A_266_409#_c_1025_n 0.00815124f $X=2.075 $Y=1.115 $X2=0
+ $Y2=0
cc_301 N_CLK_c_311_n N_A_266_409#_c_1025_n 0.0028093f $X=1.687 $Y=1.45 $X2=0
+ $Y2=0
cc_302 N_CLK_M1029_g N_A_266_409#_c_1029_n 0.00574945f $X=1.74 $Y=2.545 $X2=0
+ $Y2=0
cc_303 CLK N_A_266_409#_c_1029_n 0.0237562f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_304 N_CLK_c_310_n N_A_266_409#_c_1029_n 0.00746219f $X=1.675 $Y=1.615 $X2=0
+ $Y2=0
cc_305 N_CLK_c_311_n N_A_266_409#_c_1029_n 0.00489306f $X=1.687 $Y=1.45 $X2=0
+ $Y2=0
cc_306 N_CLK_M1029_g N_A_266_409#_c_1044_n 0.0172061f $X=1.74 $Y=2.545 $X2=0
+ $Y2=0
cc_307 N_CLK_c_308_n N_A_266_409#_c_1030_n 0.00368311f $X=1.79 $Y=1.115 $X2=0
+ $Y2=0
cc_308 CLK N_A_266_409#_c_1030_n 0.0164679f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_309 N_CLK_c_310_n N_A_266_409#_c_1030_n 0.0014112f $X=1.675 $Y=1.615 $X2=0
+ $Y2=0
cc_310 N_CLK_c_311_n N_A_266_409#_c_1030_n 0.00302257f $X=1.687 $Y=1.45 $X2=0
+ $Y2=0
cc_311 N_CLK_c_305_n N_A_266_409#_c_1031_n 0.00623428f $X=1.79 $Y=1.04 $X2=0
+ $Y2=0
cc_312 N_CLK_c_307_n N_A_266_409#_c_1031_n 3.41958e-19 $X=2.15 $Y=1.04 $X2=0
+ $Y2=0
cc_313 N_CLK_c_308_n N_A_266_409#_c_1031_n 0.00231817f $X=1.79 $Y=1.115 $X2=0
+ $Y2=0
cc_314 N_CLK_M1029_g N_A_266_409#_c_1045_n 0.0186358f $X=1.74 $Y=2.545 $X2=0
+ $Y2=0
cc_315 CLK N_A_266_409#_c_1045_n 0.0136093f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_316 N_CLK_M1029_g N_A_266_409#_c_1046_n 0.00262049f $X=1.74 $Y=2.545 $X2=0
+ $Y2=0
cc_317 CLK N_A_266_409#_c_1046_n 0.010355f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_318 N_CLK_c_310_n N_A_266_409#_c_1046_n 8.1701e-19 $X=1.675 $Y=1.615 $X2=0
+ $Y2=0
cc_319 N_CLK_c_306_n N_A_266_409#_c_1032_n 8.17524e-19 $X=2.075 $Y=1.115 $X2=0
+ $Y2=0
cc_320 CLK N_A_266_409#_c_1032_n 0.0207103f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_321 N_CLK_c_310_n N_A_266_409#_c_1032_n 0.00606856f $X=1.675 $Y=1.615 $X2=0
+ $Y2=0
cc_322 N_CLK_c_306_n N_A_266_409#_c_1033_n 0.00301619f $X=2.075 $Y=1.115 $X2=0
+ $Y2=0
cc_323 CLK N_A_266_409#_c_1033_n 2.60473e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_324 N_CLK_c_310_n N_A_266_409#_c_1033_n 0.0205055f $X=1.675 $Y=1.615 $X2=0
+ $Y2=0
cc_325 N_CLK_M1029_g N_VPWR_c_1571_n 0.0189165f $X=1.74 $Y=2.545 $X2=0 $Y2=0
cc_326 N_CLK_M1029_g N_VPWR_c_1579_n 0.00769046f $X=1.74 $Y=2.545 $X2=0 $Y2=0
cc_327 N_CLK_M1029_g N_VPWR_c_1568_n 0.0143431f $X=1.74 $Y=2.545 $X2=0 $Y2=0
cc_328 N_CLK_c_305_n N_A_135_409#_c_1713_n 0.00933678f $X=1.79 $Y=1.04 $X2=0
+ $Y2=0
cc_329 N_CLK_c_307_n N_A_135_409#_c_1713_n 8.25938e-19 $X=2.15 $Y=1.04 $X2=0
+ $Y2=0
cc_330 N_CLK_c_305_n N_A_135_409#_c_1714_n 0.00668336f $X=1.79 $Y=1.04 $X2=0
+ $Y2=0
cc_331 N_CLK_c_306_n N_A_135_409#_c_1714_n 0.0034077f $X=2.075 $Y=1.115 $X2=0
+ $Y2=0
cc_332 N_CLK_c_307_n N_A_135_409#_c_1714_n 0.0104574f $X=2.15 $Y=1.04 $X2=0
+ $Y2=0
cc_333 N_CLK_c_307_n N_A_135_409#_c_1715_n 7.17933e-19 $X=2.15 $Y=1.04 $X2=0
+ $Y2=0
cc_334 N_CLK_M1029_g N_A_135_409#_c_1720_n 0.0014722f $X=1.74 $Y=2.545 $X2=0
+ $Y2=0
cc_335 N_CLK_c_305_n N_A_135_409#_c_1721_n 0.00479956f $X=1.79 $Y=1.04 $X2=0
+ $Y2=0
cc_336 N_CLK_c_306_n N_A_135_409#_c_1722_n 0.0125242f $X=2.075 $Y=1.115 $X2=0
+ $Y2=0
cc_337 N_CLK_c_311_n N_A_135_409#_c_1722_n 0.00285323f $X=1.687 $Y=1.45 $X2=0
+ $Y2=0
cc_338 N_CLK_c_307_n N_VGND_c_1853_n 9.45515e-19 $X=2.15 $Y=1.04 $X2=0 $Y2=0
cc_339 N_CLK_c_305_n N_VGND_c_1859_n 6.46133e-19 $X=1.79 $Y=1.04 $X2=0 $Y2=0
cc_340 N_CLK_c_307_n N_VGND_c_1859_n 0.00394144f $X=2.15 $Y=1.04 $X2=0 $Y2=0
cc_341 N_CLK_c_307_n N_VGND_c_1869_n 0.00410091f $X=2.15 $Y=1.04 $X2=0 $Y2=0
cc_342 N_A_479_409#_c_389_p N_A_943_321#_M1012_d 0.00370823f $X=6.335 $Y=2.98
+ $X2=0 $Y2=0
cc_343 N_A_479_409#_c_390_p N_A_943_321#_M1027_g 0.00583866f $X=4.59 $Y=2.98
+ $X2=0 $Y2=0
cc_344 N_A_479_409#_c_391_p N_A_943_321#_M1027_g 0.0118612f $X=4.675 $Y=2.895
+ $X2=0 $Y2=0
cc_345 N_A_479_409#_c_392_p N_A_943_321#_M1027_g 0.0176646f $X=5.45 $Y=2.52
+ $X2=0 $Y2=0
cc_346 N_A_479_409#_c_393_p N_A_943_321#_M1027_g 0.00267646f $X=4.76 $Y=2.52
+ $X2=0 $Y2=0
cc_347 N_A_479_409#_c_394_p N_A_943_321#_M1027_g 0.002879f $X=5.535 $Y=2.895
+ $X2=0 $Y2=0
cc_348 N_A_479_409#_c_362_n N_A_943_321#_M1008_g 0.0124638f $X=4.445 $Y=1.215
+ $X2=0 $Y2=0
cc_349 N_A_479_409#_M1017_g N_A_943_321#_M1008_g 0.0535433f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_350 N_A_479_409#_c_365_n N_A_943_321#_M1008_g 3.75931e-19 $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_351 N_A_479_409#_c_392_p N_A_943_321#_c_597_n 0.00233487f $X=5.45 $Y=2.52
+ $X2=0 $Y2=0
cc_352 N_A_479_409#_c_392_p N_A_943_321#_c_605_n 0.0144976f $X=5.45 $Y=2.52
+ $X2=0 $Y2=0
cc_353 N_A_479_409#_c_389_p N_A_943_321#_c_605_n 0.00458866f $X=6.335 $Y=2.98
+ $X2=0 $Y2=0
cc_354 N_A_479_409#_c_401_p N_A_943_321#_c_605_n 0.00178605f $X=6.42 $Y=2.895
+ $X2=0 $Y2=0
cc_355 N_A_479_409#_c_381_n N_A_943_321#_c_605_n 0.011718f $X=6.505 $Y=2.145
+ $X2=0 $Y2=0
cc_356 N_A_479_409#_c_392_p N_A_943_321#_c_620_n 0.0257246f $X=5.45 $Y=2.52
+ $X2=0 $Y2=0
cc_357 N_A_479_409#_c_392_p N_A_943_321#_c_621_n 0.0116726f $X=5.45 $Y=2.52
+ $X2=0 $Y2=0
cc_358 N_A_479_409#_c_394_p N_A_943_321#_c_621_n 0.00673337f $X=5.535 $Y=2.895
+ $X2=0 $Y2=0
cc_359 N_A_479_409#_c_389_p N_A_943_321#_c_621_n 0.0152912f $X=6.335 $Y=2.98
+ $X2=0 $Y2=0
cc_360 N_A_479_409#_c_401_p N_A_943_321#_c_621_n 0.0313422f $X=6.42 $Y=2.895
+ $X2=0 $Y2=0
cc_361 N_A_479_409#_c_379_n N_A_709_419#_M1021_d 0.0086935f $X=3.585 $Y=2.895
+ $X2=0 $Y2=0
cc_362 N_A_479_409#_c_390_p N_A_709_419#_M1021_d 0.0159428f $X=4.59 $Y=2.98
+ $X2=0 $Y2=0
cc_363 N_A_479_409#_c_410_p N_A_709_419#_M1021_d 6.69812e-19 $X=3.585 $Y=2.98
+ $X2=0 $Y2=0
cc_364 N_A_479_409#_c_392_p N_A_709_419#_M1012_g 0.00660978f $X=5.45 $Y=2.52
+ $X2=0 $Y2=0
cc_365 N_A_479_409#_c_394_p N_A_709_419#_M1012_g 0.008974f $X=5.535 $Y=2.895
+ $X2=0 $Y2=0
cc_366 N_A_479_409#_c_389_p N_A_709_419#_M1012_g 0.0138561f $X=6.335 $Y=2.98
+ $X2=0 $Y2=0
cc_367 N_A_479_409#_c_414_p N_A_709_419#_M1012_g 0.00276664f $X=5.62 $Y=2.98
+ $X2=0 $Y2=0
cc_368 N_A_479_409#_c_401_p N_A_709_419#_M1012_g 9.90402e-19 $X=6.42 $Y=2.895
+ $X2=0 $Y2=0
cc_369 N_A_479_409#_c_401_p N_A_709_419#_M1031_g 0.002845f $X=6.42 $Y=2.895
+ $X2=0 $Y2=0
cc_370 N_A_479_409#_c_380_n N_A_709_419#_M1031_g 0.0228027f $X=7.45 $Y=2.145
+ $X2=0 $Y2=0
cc_371 N_A_479_409#_M1030_g N_A_709_419#_M1002_g 0.0440723f $X=7.555 $Y=0.835
+ $X2=0 $Y2=0
cc_372 N_A_479_409#_c_366_n N_A_709_419#_c_689_n 0.00497692f $X=7.615 $Y=1.84
+ $X2=0 $Y2=0
cc_373 N_A_479_409#_c_380_n N_A_709_419#_c_709_n 5.37369e-19 $X=7.45 $Y=2.145
+ $X2=0 $Y2=0
cc_374 N_A_479_409#_c_383_n N_A_709_419#_c_709_n 0.00489191f $X=7.615 $Y=2.06
+ $X2=0 $Y2=0
cc_375 N_A_479_409#_M1021_g N_A_709_419#_c_730_n 0.00152258f $X=3.42 $Y=2.595
+ $X2=0 $Y2=0
cc_376 N_A_479_409#_c_379_n N_A_709_419#_c_730_n 0.0343853f $X=3.585 $Y=2.895
+ $X2=0 $Y2=0
cc_377 N_A_479_409#_c_390_p N_A_709_419#_c_730_n 0.0194739f $X=4.59 $Y=2.98
+ $X2=0 $Y2=0
cc_378 N_A_479_409#_c_391_p N_A_709_419#_c_730_n 0.00409633f $X=4.675 $Y=2.895
+ $X2=0 $Y2=0
cc_379 N_A_479_409#_c_393_p N_A_709_419#_c_730_n 0.00711662f $X=4.76 $Y=2.52
+ $X2=0 $Y2=0
cc_380 N_A_479_409#_c_362_n N_A_709_419#_c_710_n 0.0026089f $X=4.445 $Y=1.215
+ $X2=0 $Y2=0
cc_381 N_A_479_409#_c_365_n N_A_709_419#_c_710_n 0.00998908f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_382 N_A_479_409#_c_390_p N_A_709_419#_c_710_n 0.00835642f $X=4.59 $Y=2.98
+ $X2=0 $Y2=0
cc_383 N_A_479_409#_c_392_p N_A_709_419#_c_710_n 0.00654666f $X=5.45 $Y=2.52
+ $X2=0 $Y2=0
cc_384 N_A_479_409#_c_393_p N_A_709_419#_c_710_n 0.00852071f $X=4.76 $Y=2.52
+ $X2=0 $Y2=0
cc_385 N_A_479_409#_M1021_g N_A_709_419#_c_711_n 6.20042e-19 $X=3.42 $Y=2.595
+ $X2=0 $Y2=0
cc_386 N_A_479_409#_c_379_n N_A_709_419#_c_711_n 0.0133149f $X=3.585 $Y=2.895
+ $X2=0 $Y2=0
cc_387 N_A_479_409#_c_365_n N_A_709_419#_c_711_n 0.0131581f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_388 N_A_479_409#_c_362_n N_A_709_419#_c_690_n 8.24358e-19 $X=4.445 $Y=1.215
+ $X2=0 $Y2=0
cc_389 N_A_479_409#_M1017_g N_A_709_419#_c_690_n 0.0110194f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_390 N_A_479_409#_c_365_n N_A_709_419#_c_690_n 0.0118253f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_391 N_A_479_409#_c_362_n N_A_709_419#_c_691_n 6.29527e-19 $X=4.445 $Y=1.215
+ $X2=0 $Y2=0
cc_392 N_A_479_409#_M1017_g N_A_709_419#_c_691_n 0.00427294f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_393 N_A_479_409#_c_365_n N_A_709_419#_c_691_n 0.0250967f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_394 N_A_479_409#_c_362_n N_A_709_419#_c_700_n 0.00383599f $X=4.445 $Y=1.215
+ $X2=0 $Y2=0
cc_395 N_A_479_409#_M1017_g N_A_709_419#_c_700_n 0.00243817f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_396 N_A_479_409#_c_365_n N_A_709_419#_c_700_n 0.0197699f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_397 N_A_479_409#_M1030_g N_A_709_419#_c_703_n 6.39263e-19 $X=7.555 $Y=0.835
+ $X2=0 $Y2=0
cc_398 N_A_479_409#_c_380_n N_A_709_419#_c_703_n 0.0214711f $X=7.45 $Y=2.145
+ $X2=0 $Y2=0
cc_399 N_A_479_409#_c_366_n N_A_709_419#_c_703_n 0.0345656f $X=7.615 $Y=1.84
+ $X2=0 $Y2=0
cc_400 N_A_479_409#_c_383_n N_A_709_419#_c_703_n 0.00199128f $X=7.615 $Y=2.06
+ $X2=0 $Y2=0
cc_401 N_A_479_409#_c_373_n N_A_709_419#_c_703_n 3.52355e-19 $X=7.615 $Y=1.465
+ $X2=0 $Y2=0
cc_402 N_A_479_409#_c_373_n N_A_709_419#_c_704_n 0.0210393f $X=7.615 $Y=1.465
+ $X2=0 $Y2=0
cc_403 N_A_479_409#_c_394_p N_SET_B_M1025_g 8.36151e-19 $X=5.535 $Y=2.895 $X2=0
+ $Y2=0
cc_404 N_A_479_409#_c_389_p N_SET_B_M1025_g 0.0183686f $X=6.335 $Y=2.98 $X2=0
+ $Y2=0
cc_405 N_A_479_409#_c_401_p N_SET_B_M1025_g 0.0209102f $X=6.42 $Y=2.895 $X2=0
+ $Y2=0
cc_406 N_A_479_409#_c_381_n N_SET_B_M1025_g 0.00794871f $X=6.505 $Y=2.145 $X2=0
+ $Y2=0
cc_407 N_A_479_409#_c_380_n N_SET_B_c_887_n 0.0185192f $X=7.45 $Y=2.145 $X2=0
+ $Y2=0
cc_408 N_A_479_409#_c_366_n N_SET_B_c_887_n 0.030967f $X=7.615 $Y=1.84 $X2=0
+ $Y2=0
cc_409 N_A_479_409#_c_367_n N_SET_B_c_887_n 0.0489827f $X=8.515 $Y=1.675 $X2=0
+ $Y2=0
cc_410 N_A_479_409#_c_368_n N_SET_B_c_887_n 0.00130212f $X=8.515 $Y=1.675 $X2=0
+ $Y2=0
cc_411 N_A_479_409#_c_380_n N_SET_B_c_888_n 7.05558e-19 $X=7.45 $Y=2.145 $X2=0
+ $Y2=0
cc_412 N_A_479_409#_c_381_n N_SET_B_c_888_n 0.00322165f $X=6.505 $Y=2.145 $X2=0
+ $Y2=0
cc_413 N_A_479_409#_c_380_n N_SET_B_c_889_n 0.01292f $X=7.45 $Y=2.145 $X2=0
+ $Y2=0
cc_414 N_A_479_409#_c_381_n N_SET_B_c_889_n 0.0080962f $X=6.505 $Y=2.145 $X2=0
+ $Y2=0
cc_415 N_A_479_409#_c_380_n N_SET_B_c_891_n 0.00492631f $X=7.45 $Y=2.145 $X2=0
+ $Y2=0
cc_416 N_A_479_409#_c_381_n N_SET_B_c_891_n 0.00254989f $X=6.505 $Y=2.145 $X2=0
+ $Y2=0
cc_417 N_A_479_409#_c_376_n N_A_266_409#_M1018_g 0.00359736f $X=2.495 $Y=2.895
+ $X2=0 $Y2=0
cc_418 N_A_479_409#_c_377_n N_A_266_409#_M1018_g 0.015584f $X=2.535 $Y=2.19
+ $X2=0 $Y2=0
cc_419 N_A_479_409#_c_369_n N_A_266_409#_M1014_g 2.98406e-19 $X=3.155 $Y=0.8
+ $X2=0 $Y2=0
cc_420 N_A_479_409#_c_370_n N_A_266_409#_c_1015_n 2.56181e-19 $X=3.41 $Y=1.41
+ $X2=0 $Y2=0
cc_421 N_A_479_409#_c_372_n N_A_266_409#_c_1015_n 0.00501786f $X=3.38 $Y=1.675
+ $X2=0 $Y2=0
cc_422 N_A_479_409#_c_369_n N_A_266_409#_M1011_g 0.00561945f $X=3.155 $Y=0.8
+ $X2=0 $Y2=0
cc_423 N_A_479_409#_c_371_n N_A_266_409#_M1011_g 0.00295297f $X=3.41 $Y=1.245
+ $X2=0 $Y2=0
cc_424 N_A_479_409#_c_365_n N_A_266_409#_c_1018_n 0.00217123f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_425 N_A_479_409#_c_369_n N_A_266_409#_c_1018_n 0.00176206f $X=3.155 $Y=0.8
+ $X2=0 $Y2=0
cc_426 N_A_479_409#_c_370_n N_A_266_409#_c_1018_n 0.019289f $X=3.41 $Y=1.41
+ $X2=0 $Y2=0
cc_427 N_A_479_409#_c_371_n N_A_266_409#_c_1018_n 0.0130753f $X=3.41 $Y=1.245
+ $X2=0 $Y2=0
cc_428 N_A_479_409#_c_372_n N_A_266_409#_c_1018_n 0.0181333f $X=3.38 $Y=1.675
+ $X2=0 $Y2=0
cc_429 N_A_479_409#_c_362_n N_A_266_409#_c_1019_n 0.0166897f $X=4.445 $Y=1.215
+ $X2=0 $Y2=0
cc_430 N_A_479_409#_c_365_n N_A_266_409#_c_1019_n 0.016368f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_431 N_A_479_409#_c_370_n N_A_266_409#_c_1019_n 0.00658409f $X=3.41 $Y=1.41
+ $X2=0 $Y2=0
cc_432 N_A_479_409#_c_372_n N_A_266_409#_c_1019_n 0.0117901f $X=3.38 $Y=1.675
+ $X2=0 $Y2=0
cc_433 N_A_479_409#_M1017_g N_A_266_409#_M1028_g 0.0193205f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_434 N_A_479_409#_c_369_n N_A_266_409#_M1028_g 8.21615e-19 $X=3.155 $Y=0.8
+ $X2=0 $Y2=0
cc_435 N_A_479_409#_c_371_n N_A_266_409#_M1028_g 0.00132699f $X=3.41 $Y=1.245
+ $X2=0 $Y2=0
cc_436 N_A_479_409#_c_362_n N_A_266_409#_c_1036_n 0.0135108f $X=4.445 $Y=1.215
+ $X2=0 $Y2=0
cc_437 N_A_479_409#_c_365_n N_A_266_409#_c_1036_n 0.00606266f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_438 N_A_479_409#_M1021_g N_A_266_409#_c_1037_n 0.0117901f $X=3.42 $Y=2.595
+ $X2=0 $Y2=0
cc_439 N_A_479_409#_c_379_n N_A_266_409#_c_1037_n 0.00503168f $X=3.585 $Y=2.895
+ $X2=0 $Y2=0
cc_440 N_A_479_409#_M1017_g N_A_266_409#_c_1021_n 0.00866282f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_441 N_A_479_409#_M1030_g N_A_266_409#_c_1021_n 0.00907339f $X=7.555 $Y=0.835
+ $X2=0 $Y2=0
cc_442 N_A_479_409#_M1021_g N_A_266_409#_M1026_g 0.0153622f $X=3.42 $Y=2.595
+ $X2=0 $Y2=0
cc_443 N_A_479_409#_c_379_n N_A_266_409#_M1026_g 0.00581636f $X=3.585 $Y=2.895
+ $X2=0 $Y2=0
cc_444 N_A_479_409#_c_390_p N_A_266_409#_M1026_g 0.0184042f $X=4.59 $Y=2.98
+ $X2=0 $Y2=0
cc_445 N_A_479_409#_c_391_p N_A_266_409#_M1026_g 0.00471947f $X=4.675 $Y=2.895
+ $X2=0 $Y2=0
cc_446 N_A_479_409#_c_393_p N_A_266_409#_M1026_g 0.00178453f $X=4.76 $Y=2.52
+ $X2=0 $Y2=0
cc_447 N_A_479_409#_M1024_g N_A_266_409#_c_1039_n 0.0103926f $X=8.505 $Y=2.595
+ $X2=0 $Y2=0
cc_448 N_A_479_409#_c_380_n N_A_266_409#_c_1039_n 0.02055f $X=7.45 $Y=2.145
+ $X2=0 $Y2=0
cc_449 N_A_479_409#_c_383_n N_A_266_409#_c_1039_n 0.00141113f $X=7.615 $Y=2.06
+ $X2=0 $Y2=0
cc_450 N_A_479_409#_c_383_n N_A_266_409#_c_1040_n 0.00509331f $X=7.615 $Y=2.06
+ $X2=0 $Y2=0
cc_451 N_A_479_409#_c_367_n N_A_266_409#_c_1040_n 0.00903469f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_452 N_A_479_409#_c_383_n N_A_266_409#_c_1041_n 0.00657293f $X=7.615 $Y=2.06
+ $X2=0 $Y2=0
cc_453 N_A_479_409#_c_373_n N_A_266_409#_c_1041_n 0.0165515f $X=7.615 $Y=1.465
+ $X2=0 $Y2=0
cc_454 N_A_479_409#_M1024_g N_A_266_409#_c_1023_n 0.0109311f $X=8.505 $Y=2.595
+ $X2=0 $Y2=0
cc_455 N_A_479_409#_c_366_n N_A_266_409#_c_1023_n 0.00140353f $X=7.615 $Y=1.84
+ $X2=0 $Y2=0
cc_456 N_A_479_409#_c_383_n N_A_266_409#_c_1023_n 0.00103042f $X=7.615 $Y=2.06
+ $X2=0 $Y2=0
cc_457 N_A_479_409#_c_367_n N_A_266_409#_c_1023_n 0.0201216f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_458 N_A_479_409#_c_368_n N_A_266_409#_c_1023_n 0.0213335f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_459 N_A_479_409#_c_373_n N_A_266_409#_c_1023_n 0.0202464f $X=7.615 $Y=1.465
+ $X2=0 $Y2=0
cc_460 N_A_479_409#_M1030_g N_A_266_409#_M1032_g 0.00524107f $X=7.555 $Y=0.835
+ $X2=0 $Y2=0
cc_461 N_A_479_409#_c_362_n N_A_266_409#_c_1027_n 0.00401937f $X=4.445 $Y=1.215
+ $X2=0 $Y2=0
cc_462 N_A_479_409#_c_365_n N_A_266_409#_c_1027_n 0.00788189f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_463 N_A_479_409#_M1030_g N_A_266_409#_c_1028_n 0.00776299f $X=7.555 $Y=0.835
+ $X2=0 $Y2=0
cc_464 N_A_479_409#_c_367_n N_A_266_409#_c_1028_n 0.00528753f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_465 N_A_479_409#_c_368_n N_A_266_409#_c_1028_n 0.00384846f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_466 N_A_479_409#_c_377_n N_A_266_409#_c_1032_n 0.0161772f $X=2.535 $Y=2.19
+ $X2=0 $Y2=0
cc_467 N_A_479_409#_c_377_n N_A_266_409#_c_1033_n 0.00740409f $X=2.535 $Y=2.19
+ $X2=0 $Y2=0
cc_468 N_A_479_409#_M1024_g N_A_1731_99#_M1000_g 0.06193f $X=8.505 $Y=2.595
+ $X2=0 $Y2=0
cc_469 N_A_479_409#_c_368_n N_A_1731_99#_c_1223_n 0.00157977f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_470 N_A_479_409#_c_367_n N_A_1731_99#_c_1225_n 4.22956e-19 $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_471 N_A_479_409#_c_368_n N_A_1731_99#_c_1225_n 0.0181638f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_472 N_A_479_409#_c_367_n N_A_1526_125#_c_1330_n 0.010837f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_473 N_A_479_409#_c_368_n N_A_1526_125#_c_1330_n 0.00532716f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_474 N_A_479_409#_M1024_g N_A_1526_125#_c_1339_n 0.0216713f $X=8.505 $Y=2.595
+ $X2=0 $Y2=0
cc_475 N_A_479_409#_c_367_n N_A_1526_125#_c_1339_n 0.0177198f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_476 N_A_479_409#_c_368_n N_A_1526_125#_c_1339_n 0.0015951f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_477 N_A_479_409#_c_380_n N_A_1526_125#_c_1340_n 0.00544411f $X=7.45 $Y=2.145
+ $X2=0 $Y2=0
cc_478 N_A_479_409#_c_383_n N_A_1526_125#_c_1340_n 0.00256314f $X=7.615 $Y=2.06
+ $X2=0 $Y2=0
cc_479 N_A_479_409#_c_367_n N_A_1526_125#_c_1340_n 0.0248301f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_480 N_A_479_409#_c_368_n N_A_1526_125#_c_1340_n 5.79521e-19 $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_481 N_A_479_409#_M1024_g N_A_1526_125#_c_1331_n 0.00363662f $X=8.505 $Y=2.595
+ $X2=0 $Y2=0
cc_482 N_A_479_409#_c_367_n N_A_1526_125#_c_1331_n 0.0234134f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_483 N_A_479_409#_c_368_n N_A_1526_125#_c_1331_n 0.00179723f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_484 N_A_479_409#_M1030_g N_A_1526_125#_c_1336_n 0.0104575f $X=7.555 $Y=0.835
+ $X2=0 $Y2=0
cc_485 N_A_479_409#_c_367_n N_A_1526_125#_c_1336_n 0.0111354f $X=8.515 $Y=1.675
+ $X2=0 $Y2=0
cc_486 N_A_479_409#_c_392_p N_VPWR_M1027_d 0.0139505f $X=5.45 $Y=2.52 $X2=0
+ $Y2=0
cc_487 N_A_479_409#_c_394_p N_VPWR_M1027_d 0.0037717f $X=5.535 $Y=2.895 $X2=0
+ $Y2=0
cc_488 N_A_479_409#_c_414_p N_VPWR_M1027_d 0.00263335f $X=5.62 $Y=2.98 $X2=0
+ $Y2=0
cc_489 N_A_479_409#_c_389_p N_VPWR_M1025_d 0.00223564f $X=6.335 $Y=2.98 $X2=0
+ $Y2=0
cc_490 N_A_479_409#_c_401_p N_VPWR_M1025_d 0.00738592f $X=6.42 $Y=2.895 $X2=0
+ $Y2=0
cc_491 N_A_479_409#_c_380_n N_VPWR_M1025_d 0.0113004f $X=7.45 $Y=2.145 $X2=0
+ $Y2=0
cc_492 N_A_479_409#_c_376_n N_VPWR_c_1571_n 0.0119061f $X=2.495 $Y=2.895 $X2=0
+ $Y2=0
cc_493 N_A_479_409#_c_377_n N_VPWR_c_1571_n 0.0377117f $X=2.535 $Y=2.19 $X2=0
+ $Y2=0
cc_494 N_A_479_409#_c_390_p N_VPWR_c_1572_n 0.0129587f $X=4.59 $Y=2.98 $X2=0
+ $Y2=0
cc_495 N_A_479_409#_c_391_p N_VPWR_c_1572_n 0.00747108f $X=4.675 $Y=2.895 $X2=0
+ $Y2=0
cc_496 N_A_479_409#_c_392_p N_VPWR_c_1572_n 0.020016f $X=5.45 $Y=2.52 $X2=0
+ $Y2=0
cc_497 N_A_479_409#_c_394_p N_VPWR_c_1572_n 0.00802182f $X=5.535 $Y=2.895 $X2=0
+ $Y2=0
cc_498 N_A_479_409#_c_414_p N_VPWR_c_1572_n 0.0138718f $X=5.62 $Y=2.98 $X2=0
+ $Y2=0
cc_499 N_A_479_409#_c_389_p N_VPWR_c_1573_n 0.0138718f $X=6.335 $Y=2.98 $X2=0
+ $Y2=0
cc_500 N_A_479_409#_c_401_p N_VPWR_c_1573_n 0.0354875f $X=6.42 $Y=2.895 $X2=0
+ $Y2=0
cc_501 N_A_479_409#_c_380_n N_VPWR_c_1573_n 0.0209601f $X=7.45 $Y=2.145 $X2=0
+ $Y2=0
cc_502 N_A_479_409#_M1024_g N_VPWR_c_1574_n 0.00396249f $X=8.505 $Y=2.595 $X2=0
+ $Y2=0
cc_503 N_A_479_409#_M1021_g N_VPWR_c_1580_n 0.00599878f $X=3.42 $Y=2.595 $X2=0
+ $Y2=0
cc_504 N_A_479_409#_c_376_n N_VPWR_c_1580_n 0.0167695f $X=2.495 $Y=2.895 $X2=0
+ $Y2=0
cc_505 N_A_479_409#_c_378_n N_VPWR_c_1580_n 0.0509285f $X=3.5 $Y=2.98 $X2=0
+ $Y2=0
cc_506 N_A_479_409#_c_390_p N_VPWR_c_1580_n 0.0605701f $X=4.59 $Y=2.98 $X2=0
+ $Y2=0
cc_507 N_A_479_409#_c_392_p N_VPWR_c_1580_n 0.00239177f $X=5.45 $Y=2.52 $X2=0
+ $Y2=0
cc_508 N_A_479_409#_c_410_p N_VPWR_c_1580_n 0.0092477f $X=3.585 $Y=2.98 $X2=0
+ $Y2=0
cc_509 N_A_479_409#_c_392_p N_VPWR_c_1581_n 0.00258613f $X=5.45 $Y=2.52 $X2=0
+ $Y2=0
cc_510 N_A_479_409#_c_389_p N_VPWR_c_1581_n 0.0480507f $X=6.335 $Y=2.98 $X2=0
+ $Y2=0
cc_511 N_A_479_409#_c_414_p N_VPWR_c_1581_n 0.0092917f $X=5.62 $Y=2.98 $X2=0
+ $Y2=0
cc_512 N_A_479_409#_M1024_g N_VPWR_c_1582_n 0.00975641f $X=8.505 $Y=2.595 $X2=0
+ $Y2=0
cc_513 N_A_479_409#_M1021_g N_VPWR_c_1568_n 0.0100086f $X=3.42 $Y=2.595 $X2=0
+ $Y2=0
cc_514 N_A_479_409#_M1024_g N_VPWR_c_1568_n 0.0177985f $X=8.505 $Y=2.595 $X2=0
+ $Y2=0
cc_515 N_A_479_409#_c_376_n N_VPWR_c_1568_n 0.00955814f $X=2.495 $Y=2.895 $X2=0
+ $Y2=0
cc_516 N_A_479_409#_c_378_n N_VPWR_c_1568_n 0.0319421f $X=3.5 $Y=2.98 $X2=0
+ $Y2=0
cc_517 N_A_479_409#_c_390_p N_VPWR_c_1568_n 0.0395874f $X=4.59 $Y=2.98 $X2=0
+ $Y2=0
cc_518 N_A_479_409#_c_392_p N_VPWR_c_1568_n 0.0100314f $X=5.45 $Y=2.52 $X2=0
+ $Y2=0
cc_519 N_A_479_409#_c_389_p N_VPWR_c_1568_n 0.0310933f $X=6.335 $Y=2.98 $X2=0
+ $Y2=0
cc_520 N_A_479_409#_c_414_p N_VPWR_c_1568_n 0.00647207f $X=5.62 $Y=2.98 $X2=0
+ $Y2=0
cc_521 N_A_479_409#_c_410_p N_VPWR_c_1568_n 0.00636511f $X=3.585 $Y=2.98 $X2=0
+ $Y2=0
cc_522 N_A_479_409#_c_378_n N_A_135_409#_M1021_s 0.00565337f $X=3.5 $Y=2.98
+ $X2=0 $Y2=0
cc_523 N_A_479_409#_c_369_n N_A_135_409#_c_1715_n 0.0250978f $X=3.155 $Y=0.8
+ $X2=0 $Y2=0
cc_524 N_A_479_409#_c_371_n N_A_135_409#_c_1715_n 0.00519103f $X=3.41 $Y=1.245
+ $X2=0 $Y2=0
cc_525 N_A_479_409#_c_369_n N_A_135_409#_c_1716_n 0.0216701f $X=3.155 $Y=0.8
+ $X2=0 $Y2=0
cc_526 N_A_479_409#_M1021_g N_A_135_409#_c_1718_n 0.00477676f $X=3.42 $Y=2.595
+ $X2=0 $Y2=0
cc_527 N_A_479_409#_c_377_n N_A_135_409#_c_1718_n 0.00368124f $X=2.535 $Y=2.19
+ $X2=0 $Y2=0
cc_528 N_A_479_409#_c_379_n N_A_135_409#_c_1718_n 0.00713479f $X=3.585 $Y=2.895
+ $X2=0 $Y2=0
cc_529 N_A_479_409#_c_370_n N_A_135_409#_c_1718_n 0.0398545f $X=3.41 $Y=1.41
+ $X2=0 $Y2=0
cc_530 N_A_479_409#_c_372_n N_A_135_409#_c_1718_n 0.00109107f $X=3.38 $Y=1.675
+ $X2=0 $Y2=0
cc_531 N_A_479_409#_M1017_g N_A_135_409#_c_1719_n 5.84395e-19 $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_532 N_A_479_409#_c_365_n N_A_135_409#_c_1719_n 0.0135077f $X=4.34 $Y=1.41
+ $X2=0 $Y2=0
cc_533 N_A_479_409#_c_369_n N_A_135_409#_c_1719_n 0.0343215f $X=3.155 $Y=0.8
+ $X2=0 $Y2=0
cc_534 N_A_479_409#_c_370_n N_A_135_409#_c_1719_n 0.013485f $X=3.41 $Y=1.41
+ $X2=0 $Y2=0
cc_535 N_A_479_409#_c_371_n N_A_135_409#_c_1722_n 0.0163999f $X=3.41 $Y=1.245
+ $X2=0 $Y2=0
cc_536 N_A_479_409#_M1021_g N_A_135_409#_c_1727_n 0.0172542f $X=3.42 $Y=2.595
+ $X2=0 $Y2=0
cc_537 N_A_479_409#_c_377_n N_A_135_409#_c_1727_n 0.0510745f $X=2.535 $Y=2.19
+ $X2=0 $Y2=0
cc_538 N_A_479_409#_c_378_n N_A_135_409#_c_1727_n 0.0337547f $X=3.5 $Y=2.98
+ $X2=0 $Y2=0
cc_539 N_A_479_409#_c_379_n N_A_135_409#_c_1727_n 0.0453832f $X=3.585 $Y=2.895
+ $X2=0 $Y2=0
cc_540 N_A_479_409#_c_370_n N_A_135_409#_c_1727_n 0.0118927f $X=3.41 $Y=1.41
+ $X2=0 $Y2=0
cc_541 N_A_479_409#_c_372_n N_A_135_409#_c_1727_n 6.00432e-19 $X=3.38 $Y=1.675
+ $X2=0 $Y2=0
cc_542 N_A_479_409#_c_390_p A_881_419# 0.00453514f $X=4.59 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_543 N_A_479_409#_c_391_p A_881_419# 0.00342086f $X=4.675 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_544 N_A_479_409#_c_393_p A_881_419# 0.00294757f $X=4.76 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_545 N_A_479_409#_c_380_n A_1448_419# 0.0048076f $X=7.45 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_546 N_A_479_409#_M1017_g N_VGND_c_1869_n 9.49986e-19 $X=4.445 $Y=0.835 $X2=0
+ $Y2=0
cc_547 N_A_479_409#_M1030_g N_VGND_c_1869_n 9.49986e-19 $X=7.555 $Y=0.835 $X2=0
+ $Y2=0
cc_548 N_A_943_321#_M1027_g N_A_709_419#_M1012_g 0.0162417f $X=4.84 $Y=2.595
+ $X2=0 $Y2=0
cc_549 N_A_943_321#_c_596_n N_A_709_419#_M1012_g 0.00400351f $X=5.2 $Y=1.77
+ $X2=0 $Y2=0
cc_550 N_A_943_321#_c_597_n N_A_709_419#_M1012_g 0.00185332f $X=5.2 $Y=1.77
+ $X2=0 $Y2=0
cc_551 N_A_943_321#_c_605_n N_A_709_419#_M1012_g 0.0181779f $X=5.825 $Y=2.17
+ $X2=0 $Y2=0
cc_552 N_A_943_321#_c_621_n N_A_709_419#_M1012_g 0.0147646f $X=5.99 $Y=2.4 $X2=0
+ $Y2=0
cc_553 N_A_943_321#_c_598_n N_A_709_419#_c_686_n 0.0022395f $X=5.695 $Y=1.31
+ $X2=0 $Y2=0
cc_554 N_A_943_321#_c_600_n N_A_709_419#_c_686_n 0.00633769f $X=5.78 $Y=1.225
+ $X2=0 $Y2=0
cc_555 N_A_943_321#_c_601_n N_A_709_419#_c_686_n 0.0074733f $X=5.99 $Y=0.815
+ $X2=0 $Y2=0
cc_556 N_A_943_321#_c_600_n N_A_709_419#_c_687_n 0.00196192f $X=5.78 $Y=1.225
+ $X2=0 $Y2=0
cc_557 N_A_943_321#_c_601_n N_A_709_419#_c_687_n 0.00508272f $X=5.99 $Y=0.815
+ $X2=0 $Y2=0
cc_558 N_A_943_321#_M1027_g N_A_709_419#_c_730_n 0.00103959f $X=4.84 $Y=2.595
+ $X2=0 $Y2=0
cc_559 N_A_943_321#_M1027_g N_A_709_419#_c_710_n 0.00795583f $X=4.84 $Y=2.595
+ $X2=0 $Y2=0
cc_560 N_A_943_321#_c_596_n N_A_709_419#_c_710_n 7.63318e-19 $X=5.2 $Y=1.77
+ $X2=0 $Y2=0
cc_561 N_A_943_321#_c_620_n N_A_709_419#_c_710_n 0.0133914f $X=5.365 $Y=2.17
+ $X2=0 $Y2=0
cc_562 N_A_943_321#_M1027_g N_A_709_419#_c_691_n 0.00358566f $X=4.84 $Y=2.595
+ $X2=0 $Y2=0
cc_563 N_A_943_321#_M1008_g N_A_709_419#_c_691_n 0.0161946f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_564 N_A_943_321#_c_596_n N_A_709_419#_c_691_n 0.0476915f $X=5.2 $Y=1.77 $X2=0
+ $Y2=0
cc_565 N_A_943_321#_c_597_n N_A_709_419#_c_691_n 0.0129359f $X=5.2 $Y=1.77 $X2=0
+ $Y2=0
cc_566 N_A_943_321#_c_599_n N_A_709_419#_c_691_n 0.0131397f $X=5.365 $Y=1.31
+ $X2=0 $Y2=0
cc_567 N_A_943_321#_M1008_g N_A_709_419#_c_692_n 0.0058447f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_568 N_A_943_321#_c_597_n N_A_709_419#_c_692_n 0.00451047f $X=5.2 $Y=1.77
+ $X2=0 $Y2=0
cc_569 N_A_943_321#_c_598_n N_A_709_419#_c_692_n 0.0121295f $X=5.695 $Y=1.31
+ $X2=0 $Y2=0
cc_570 N_A_943_321#_c_599_n N_A_709_419#_c_692_n 0.0266477f $X=5.365 $Y=1.31
+ $X2=0 $Y2=0
cc_571 N_A_943_321#_c_600_n N_A_709_419#_c_692_n 0.00202763f $X=5.78 $Y=1.225
+ $X2=0 $Y2=0
cc_572 N_A_943_321#_c_601_n N_A_709_419#_c_692_n 0.0125835f $X=5.99 $Y=0.815
+ $X2=0 $Y2=0
cc_573 N_A_943_321#_M1008_g N_A_709_419#_c_693_n 0.00477288f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_574 N_A_943_321#_c_601_n N_A_709_419#_c_693_n 0.0203077f $X=5.99 $Y=0.815
+ $X2=0 $Y2=0
cc_575 N_A_943_321#_c_601_n N_A_709_419#_c_694_n 0.0331438f $X=5.99 $Y=0.815
+ $X2=0 $Y2=0
cc_576 N_A_943_321#_c_598_n N_A_709_419#_c_696_n 0.00191277f $X=5.695 $Y=1.31
+ $X2=0 $Y2=0
cc_577 N_A_943_321#_c_600_n N_A_709_419#_c_697_n 0.00585263f $X=5.78 $Y=1.225
+ $X2=0 $Y2=0
cc_578 N_A_943_321#_c_601_n N_A_709_419#_c_697_n 0.0155651f $X=5.99 $Y=0.815
+ $X2=0 $Y2=0
cc_579 N_A_943_321#_c_598_n N_A_709_419#_c_699_n 0.0120466f $X=5.695 $Y=1.31
+ $X2=0 $Y2=0
cc_580 N_A_943_321#_c_600_n N_A_709_419#_c_699_n 0.0017133f $X=5.78 $Y=1.225
+ $X2=0 $Y2=0
cc_581 N_A_943_321#_c_601_n N_A_709_419#_c_699_n 0.0055626f $X=5.99 $Y=0.815
+ $X2=0 $Y2=0
cc_582 N_A_943_321#_M1008_g N_A_709_419#_c_792_n 0.00751838f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_583 N_A_943_321#_c_596_n N_A_709_419#_c_701_n 0.0217027f $X=5.2 $Y=1.77 $X2=0
+ $Y2=0
cc_584 N_A_943_321#_c_597_n N_A_709_419#_c_701_n 0.00118806f $X=5.2 $Y=1.77
+ $X2=0 $Y2=0
cc_585 N_A_943_321#_c_598_n N_A_709_419#_c_701_n 0.0213298f $X=5.695 $Y=1.31
+ $X2=0 $Y2=0
cc_586 N_A_943_321#_c_605_n N_A_709_419#_c_701_n 0.0367762f $X=5.825 $Y=2.17
+ $X2=0 $Y2=0
cc_587 N_A_943_321#_c_601_n N_A_709_419#_c_701_n 0.00599133f $X=5.99 $Y=0.815
+ $X2=0 $Y2=0
cc_588 N_A_943_321#_M1008_g N_A_709_419#_c_702_n 2.71876e-19 $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_589 N_A_943_321#_c_596_n N_A_709_419#_c_702_n 5.17216e-19 $X=5.2 $Y=1.77
+ $X2=0 $Y2=0
cc_590 N_A_943_321#_c_597_n N_A_709_419#_c_702_n 0.0198572f $X=5.2 $Y=1.77 $X2=0
+ $Y2=0
cc_591 N_A_943_321#_c_598_n N_A_709_419#_c_702_n 0.00126488f $X=5.695 $Y=1.31
+ $X2=0 $Y2=0
cc_592 N_A_943_321#_c_605_n N_A_709_419#_c_702_n 5.95935e-19 $X=5.825 $Y=2.17
+ $X2=0 $Y2=0
cc_593 N_A_943_321#_c_596_n N_A_709_419#_c_705_n 0.00525934f $X=5.2 $Y=1.77
+ $X2=0 $Y2=0
cc_594 N_A_943_321#_c_598_n N_A_709_419#_c_705_n 0.00660224f $X=5.695 $Y=1.31
+ $X2=0 $Y2=0
cc_595 N_A_943_321#_c_605_n N_SET_B_M1025_g 0.00435166f $X=5.825 $Y=2.17 $X2=0
+ $Y2=0
cc_596 N_A_943_321#_c_621_n N_SET_B_M1025_g 0.00862371f $X=5.99 $Y=2.4 $X2=0
+ $Y2=0
cc_597 N_A_943_321#_c_597_n N_A_266_409#_c_1036_n 0.028257f $X=5.2 $Y=1.77 $X2=0
+ $Y2=0
cc_598 N_A_943_321#_M1008_g N_A_266_409#_c_1021_n 0.00866194f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_599 N_A_943_321#_M1027_g N_A_266_409#_M1026_g 0.028257f $X=4.84 $Y=2.595
+ $X2=0 $Y2=0
cc_600 N_A_943_321#_c_605_n N_VPWR_M1027_d 0.00234485f $X=5.825 $Y=2.17 $X2=0
+ $Y2=0
cc_601 N_A_943_321#_c_620_n N_VPWR_M1027_d 0.00772784f $X=5.365 $Y=2.17 $X2=0
+ $Y2=0
cc_602 N_A_943_321#_M1027_g N_VPWR_c_1572_n 0.0109804f $X=4.84 $Y=2.595 $X2=0
+ $Y2=0
cc_603 N_A_943_321#_M1027_g N_VPWR_c_1580_n 0.00632556f $X=4.84 $Y=2.595 $X2=0
+ $Y2=0
cc_604 N_A_943_321#_M1012_d N_VPWR_c_1568_n 0.00237544f $X=5.85 $Y=2.095 $X2=0
+ $Y2=0
cc_605 N_A_943_321#_M1027_g N_VPWR_c_1568_n 0.00726189f $X=4.84 $Y=2.595 $X2=0
+ $Y2=0
cc_606 N_A_943_321#_M1008_g N_VGND_c_1854_n 0.0065032f $X=4.805 $Y=0.835 $X2=0
+ $Y2=0
cc_607 N_A_943_321#_M1008_g N_VGND_c_1869_n 9.49986e-19 $X=4.805 $Y=0.835 $X2=0
+ $Y2=0
cc_608 N_A_709_419#_M1012_g N_SET_B_M1025_g 0.0421444f $X=5.725 $Y=2.595 $X2=0
+ $Y2=0
cc_609 N_A_709_419#_M1031_g N_SET_B_M1025_g 0.0166646f $X=7.115 $Y=2.595 $X2=0
+ $Y2=0
cc_610 N_A_709_419#_c_702_n N_SET_B_M1025_g 0.00969012f $X=5.74 $Y=1.74 $X2=0
+ $Y2=0
cc_611 N_A_709_419#_c_687_n N_SET_B_M1007_g 0.0347345f $X=6.205 $Y=1.12 $X2=0
+ $Y2=0
cc_612 N_A_709_419#_M1002_g N_SET_B_M1007_g 0.0118375f $X=7.165 $Y=0.835 $X2=0
+ $Y2=0
cc_613 N_A_709_419#_c_696_n N_SET_B_M1007_g 0.00361263f $X=6.13 $Y=1.575 $X2=0
+ $Y2=0
cc_614 N_A_709_419#_c_697_n N_SET_B_M1007_g 0.00639012f $X=6.42 $Y=1.2 $X2=0
+ $Y2=0
cc_615 N_A_709_419#_c_698_n N_SET_B_M1007_g 0.0152587f $X=6.91 $Y=1.285 $X2=0
+ $Y2=0
cc_616 N_A_709_419#_c_703_n N_SET_B_M1007_g 0.00115985f $X=7.075 $Y=1.365 $X2=0
+ $Y2=0
cc_617 N_A_709_419#_c_704_n N_SET_B_M1007_g 0.0188683f $X=7.075 $Y=1.365 $X2=0
+ $Y2=0
cc_618 N_A_709_419#_c_705_n N_SET_B_M1007_g 0.00315923f $X=5.74 $Y=1.575 $X2=0
+ $Y2=0
cc_619 N_A_709_419#_c_689_n N_SET_B_c_887_n 0.00192821f $X=7.075 $Y=1.705 $X2=0
+ $Y2=0
cc_620 N_A_709_419#_c_709_n N_SET_B_c_887_n 6.40922e-19 $X=7.075 $Y=1.87 $X2=0
+ $Y2=0
cc_621 N_A_709_419#_c_698_n N_SET_B_c_887_n 0.00949416f $X=6.91 $Y=1.285 $X2=0
+ $Y2=0
cc_622 N_A_709_419#_c_703_n N_SET_B_c_887_n 0.0254227f $X=7.075 $Y=1.365 $X2=0
+ $Y2=0
cc_623 N_A_709_419#_c_696_n N_SET_B_c_888_n 6.64545e-19 $X=6.13 $Y=1.575 $X2=0
+ $Y2=0
cc_624 N_A_709_419#_c_699_n N_SET_B_c_888_n 0.00795812f $X=6.505 $Y=1.285 $X2=0
+ $Y2=0
cc_625 N_A_709_419#_c_701_n N_SET_B_c_888_n 0.00596941f $X=5.74 $Y=1.74 $X2=0
+ $Y2=0
cc_626 N_A_709_419#_c_703_n N_SET_B_c_888_n 5.35001e-19 $X=7.075 $Y=1.365 $X2=0
+ $Y2=0
cc_627 N_A_709_419#_c_689_n N_SET_B_c_889_n 0.00109386f $X=7.075 $Y=1.705 $X2=0
+ $Y2=0
cc_628 N_A_709_419#_c_696_n N_SET_B_c_889_n 0.0013199f $X=6.13 $Y=1.575 $X2=0
+ $Y2=0
cc_629 N_A_709_419#_c_699_n N_SET_B_c_889_n 0.0180783f $X=6.505 $Y=1.285 $X2=0
+ $Y2=0
cc_630 N_A_709_419#_c_701_n N_SET_B_c_889_n 0.0142964f $X=5.74 $Y=1.74 $X2=0
+ $Y2=0
cc_631 N_A_709_419#_c_702_n N_SET_B_c_889_n 2.94012e-19 $X=5.74 $Y=1.74 $X2=0
+ $Y2=0
cc_632 N_A_709_419#_c_703_n N_SET_B_c_889_n 0.0180089f $X=7.075 $Y=1.365 $X2=0
+ $Y2=0
cc_633 N_A_709_419#_c_685_n N_SET_B_c_891_n 0.00618481f $X=6.13 $Y=1.195 $X2=0
+ $Y2=0
cc_634 N_A_709_419#_M1031_g N_SET_B_c_891_n 4.10212e-19 $X=7.115 $Y=2.595 $X2=0
+ $Y2=0
cc_635 N_A_709_419#_c_689_n N_SET_B_c_891_n 0.0208611f $X=7.075 $Y=1.705 $X2=0
+ $Y2=0
cc_636 N_A_709_419#_c_696_n N_SET_B_c_891_n 0.00114006f $X=6.13 $Y=1.575 $X2=0
+ $Y2=0
cc_637 N_A_709_419#_c_698_n N_SET_B_c_891_n 6.68297e-19 $X=6.91 $Y=1.285 $X2=0
+ $Y2=0
cc_638 N_A_709_419#_c_699_n N_SET_B_c_891_n 0.00785599f $X=6.505 $Y=1.285 $X2=0
+ $Y2=0
cc_639 N_A_709_419#_c_701_n N_SET_B_c_891_n 0.00909892f $X=5.74 $Y=1.74 $X2=0
+ $Y2=0
cc_640 N_A_709_419#_c_703_n N_SET_B_c_891_n 4.99368e-19 $X=7.075 $Y=1.365 $X2=0
+ $Y2=0
cc_641 N_A_709_419#_c_705_n N_SET_B_c_891_n 0.00969012f $X=5.74 $Y=1.575 $X2=0
+ $Y2=0
cc_642 N_A_709_419#_c_700_n N_A_266_409#_M1028_g 0.0040354f $X=4.17 $Y=0.835
+ $X2=0 $Y2=0
cc_643 N_A_709_419#_c_691_n N_A_266_409#_c_1036_n 0.00497102f $X=4.77 $Y=2.075
+ $X2=0 $Y2=0
cc_644 N_A_709_419#_c_711_n N_A_266_409#_c_1037_n 0.00875525f $X=4.18 $Y=2.16
+ $X2=0 $Y2=0
cc_645 N_A_709_419#_c_687_n N_A_266_409#_c_1021_n 0.00737233f $X=6.205 $Y=1.12
+ $X2=0 $Y2=0
cc_646 N_A_709_419#_M1002_g N_A_266_409#_c_1021_n 0.00907339f $X=7.165 $Y=0.835
+ $X2=0 $Y2=0
cc_647 N_A_709_419#_c_690_n N_A_266_409#_c_1021_n 0.00330026f $X=4.685 $Y=0.97
+ $X2=0 $Y2=0
cc_648 N_A_709_419#_c_692_n N_A_266_409#_c_1021_n 0.0046601f $X=5.345 $Y=0.96
+ $X2=0 $Y2=0
cc_649 N_A_709_419#_c_694_n N_A_266_409#_c_1021_n 0.0209179f $X=6.335 $Y=0.35
+ $X2=0 $Y2=0
cc_650 N_A_709_419#_c_695_n N_A_266_409#_c_1021_n 0.00418768f $X=5.515 $Y=0.35
+ $X2=0 $Y2=0
cc_651 N_A_709_419#_c_700_n N_A_266_409#_c_1021_n 0.00478092f $X=4.17 $Y=0.835
+ $X2=0 $Y2=0
cc_652 N_A_709_419#_c_792_n N_A_266_409#_c_1021_n 3.9237e-19 $X=4.77 $Y=0.97
+ $X2=0 $Y2=0
cc_653 N_A_709_419#_c_730_n N_A_266_409#_M1026_g 0.0112713f $X=4.015 $Y=2.395
+ $X2=0 $Y2=0
cc_654 N_A_709_419#_c_710_n N_A_266_409#_M1026_g 0.0160425f $X=4.685 $Y=2.16
+ $X2=0 $Y2=0
cc_655 N_A_709_419#_c_711_n N_A_266_409#_M1026_g 0.00278888f $X=4.18 $Y=2.16
+ $X2=0 $Y2=0
cc_656 N_A_709_419#_M1031_g N_A_266_409#_c_1041_n 0.0787068f $X=7.115 $Y=2.595
+ $X2=0 $Y2=0
cc_657 N_A_709_419#_M1012_g N_VPWR_c_1572_n 0.00341965f $X=5.725 $Y=2.595 $X2=0
+ $Y2=0
cc_658 N_A_709_419#_M1031_g N_VPWR_c_1573_n 0.0193116f $X=7.115 $Y=2.595 $X2=0
+ $Y2=0
cc_659 N_A_709_419#_M1012_g N_VPWR_c_1581_n 0.00599913f $X=5.725 $Y=2.595 $X2=0
+ $Y2=0
cc_660 N_A_709_419#_M1031_g N_VPWR_c_1582_n 0.008763f $X=7.115 $Y=2.595 $X2=0
+ $Y2=0
cc_661 N_A_709_419#_M1021_d N_VPWR_c_1568_n 0.00499582f $X=3.545 $Y=2.095 $X2=0
+ $Y2=0
cc_662 N_A_709_419#_M1012_g N_VPWR_c_1568_n 0.00868967f $X=5.725 $Y=2.595 $X2=0
+ $Y2=0
cc_663 N_A_709_419#_M1031_g N_VPWR_c_1568_n 0.0144563f $X=7.115 $Y=2.595 $X2=0
+ $Y2=0
cc_664 N_A_709_419#_c_700_n N_A_135_409#_c_1719_n 0.0264655f $X=4.17 $Y=0.835
+ $X2=0 $Y2=0
cc_665 N_A_709_419#_c_710_n A_881_419# 0.00341639f $X=4.685 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_666 N_A_709_419#_c_692_n N_VGND_M1008_d 0.00829139f $X=5.345 $Y=0.96 $X2=0
+ $Y2=0
cc_667 N_A_709_419#_c_692_n N_VGND_c_1854_n 0.0176954f $X=5.345 $Y=0.96 $X2=0
+ $Y2=0
cc_668 N_A_709_419#_c_693_n N_VGND_c_1854_n 0.0189538f $X=5.43 $Y=0.875 $X2=0
+ $Y2=0
cc_669 N_A_709_419#_c_695_n N_VGND_c_1854_n 0.0140867f $X=5.515 $Y=0.35 $X2=0
+ $Y2=0
cc_670 N_A_709_419#_c_700_n N_VGND_c_1854_n 6.37013e-19 $X=4.17 $Y=0.835 $X2=0
+ $Y2=0
cc_671 N_A_709_419#_M1002_g N_VGND_c_1855_n 0.0147625f $X=7.165 $Y=0.835 $X2=0
+ $Y2=0
cc_672 N_A_709_419#_c_694_n N_VGND_c_1855_n 0.0144411f $X=6.335 $Y=0.35 $X2=0
+ $Y2=0
cc_673 N_A_709_419#_c_697_n N_VGND_c_1855_n 0.0143489f $X=6.42 $Y=1.2 $X2=0
+ $Y2=0
cc_674 N_A_709_419#_c_698_n N_VGND_c_1855_n 0.0154758f $X=6.91 $Y=1.285 $X2=0
+ $Y2=0
cc_675 N_A_709_419#_c_703_n N_VGND_c_1855_n 0.0084084f $X=7.075 $Y=1.365 $X2=0
+ $Y2=0
cc_676 N_A_709_419#_c_704_n N_VGND_c_1855_n 8.08179e-19 $X=7.075 $Y=1.365 $X2=0
+ $Y2=0
cc_677 N_A_709_419#_c_700_n N_VGND_c_1865_n 0.00518815f $X=4.17 $Y=0.835 $X2=0
+ $Y2=0
cc_678 N_A_709_419#_c_694_n N_VGND_c_1866_n 0.0611043f $X=6.335 $Y=0.35 $X2=0
+ $Y2=0
cc_679 N_A_709_419#_c_695_n N_VGND_c_1866_n 0.0114574f $X=5.515 $Y=0.35 $X2=0
+ $Y2=0
cc_680 N_A_709_419#_M1002_g N_VGND_c_1869_n 9.49986e-19 $X=7.165 $Y=0.835 $X2=0
+ $Y2=0
cc_681 N_A_709_419#_c_694_n N_VGND_c_1869_n 0.0332665f $X=6.335 $Y=0.35 $X2=0
+ $Y2=0
cc_682 N_A_709_419#_c_695_n N_VGND_c_1869_n 0.00589978f $X=5.515 $Y=0.35 $X2=0
+ $Y2=0
cc_683 N_A_709_419#_c_700_n N_VGND_c_1869_n 0.00658035f $X=4.17 $Y=0.835 $X2=0
+ $Y2=0
cc_684 N_A_709_419#_c_690_n A_904_125# 0.00165782f $X=4.685 $Y=0.97 $X2=-0.19
+ $Y2=-0.245
cc_685 N_A_709_419#_c_697_n A_1256_125# 0.00276176f $X=6.42 $Y=1.2 $X2=-0.19
+ $Y2=-0.245
cc_686 N_SET_B_M1007_g N_A_266_409#_c_1021_n 0.00907339f $X=6.595 $Y=0.835 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_884_n N_A_1731_99#_c_1221_n 0.0137654f $X=9.385 $Y=1.12 $X2=0
+ $Y2=0
cc_688 N_SET_B_M1033_g N_A_1731_99#_M1000_g 0.0211122f $X=9.825 $Y=2.595 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_886_n N_A_1731_99#_c_1223_n 0.00842804f $X=9.46 $Y=1.195 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_887_n N_A_1731_99#_c_1223_n 0.00391638f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_691 N_SET_B_c_887_n N_A_1731_99#_c_1224_n 0.0216657f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_692 SET_B N_A_1731_99#_c_1224_n 0.00251515f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_693 N_SET_B_c_892_n N_A_1731_99#_c_1224_n 5.11574e-19 $X=9.865 $Y=1.675 $X2=0
+ $Y2=0
cc_694 N_SET_B_c_893_n N_A_1731_99#_c_1224_n 0.00520801f $X=9.865 $Y=1.51 $X2=0
+ $Y2=0
cc_695 N_SET_B_c_894_n N_A_1731_99#_c_1224_n 0.0179394f $X=9.84 $Y=1.665 $X2=0
+ $Y2=0
cc_696 N_SET_B_c_886_n N_A_1731_99#_c_1225_n 0.00990538f $X=9.46 $Y=1.195 $X2=0
+ $Y2=0
cc_697 N_SET_B_c_887_n N_A_1731_99#_c_1225_n 0.00911931f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_698 SET_B N_A_1731_99#_c_1225_n 0.00136744f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_699 N_SET_B_c_892_n N_A_1731_99#_c_1225_n 0.0220623f $X=9.865 $Y=1.675 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_894_n N_A_1731_99#_c_1225_n 0.00128279f $X=9.84 $Y=1.665 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_885_n N_A_1731_99#_c_1226_n 0.0231371f $X=9.88 $Y=1.195 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_887_n N_A_1731_99#_c_1226_n 0.00843014f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_703 SET_B N_A_1731_99#_c_1226_n 0.00211686f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_704 N_SET_B_c_892_n N_A_1731_99#_c_1226_n 0.00114177f $X=9.865 $Y=1.675 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_893_n N_A_1731_99#_c_1226_n 0.00543754f $X=9.865 $Y=1.51 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_894_n N_A_1731_99#_c_1226_n 0.0213366f $X=9.84 $Y=1.665 $X2=0
+ $Y2=0
cc_707 N_SET_B_c_885_n N_A_1731_99#_c_1227_n 7.70696e-19 $X=9.88 $Y=1.195 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_886_n N_A_1731_99#_c_1227_n 0.0104092f $X=9.46 $Y=1.195 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_884_n N_A_1731_99#_c_1228_n 0.00445383f $X=9.385 $Y=1.12 $X2=0
+ $Y2=0
cc_710 N_SET_B_c_885_n N_A_1731_99#_c_1228_n 0.00146245f $X=9.88 $Y=1.195 $X2=0
+ $Y2=0
cc_711 N_SET_B_M1033_g N_A_1731_99#_c_1235_n 0.00652645f $X=9.825 $Y=2.595 $X2=0
+ $Y2=0
cc_712 SET_B N_A_1731_99#_c_1230_n 0.00142847f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_713 N_SET_B_c_892_n N_A_1731_99#_c_1230_n 0.00188194f $X=9.865 $Y=1.675 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_893_n N_A_1731_99#_c_1230_n 0.00323744f $X=9.865 $Y=1.51 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_894_n N_A_1731_99#_c_1230_n 0.0103099f $X=9.84 $Y=1.665 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_893_n N_A_1526_125#_c_1327_n 0.00190545f $X=9.865 $Y=1.51 $X2=0
+ $Y2=0
cc_717 N_SET_B_c_884_n N_A_1526_125#_c_1330_n 0.00297501f $X=9.385 $Y=1.12 $X2=0
+ $Y2=0
cc_718 N_SET_B_c_887_n N_A_1526_125#_c_1330_n 0.00724916f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_719 N_SET_B_c_887_n N_A_1526_125#_c_1339_n 0.00873876f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_720 N_SET_B_c_887_n N_A_1526_125#_c_1340_n 0.00217478f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_721 N_SET_B_c_884_n N_A_1526_125#_c_1331_n 0.00104439f $X=9.385 $Y=1.12 $X2=0
+ $Y2=0
cc_722 N_SET_B_c_886_n N_A_1526_125#_c_1331_n 3.6489e-19 $X=9.46 $Y=1.195 $X2=0
+ $Y2=0
cc_723 N_SET_B_c_887_n N_A_1526_125#_c_1331_n 0.0204045f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_892_n N_A_1526_125#_c_1331_n 7.79626e-19 $X=9.865 $Y=1.675
+ $X2=0 $Y2=0
cc_725 N_SET_B_M1033_g N_A_1526_125#_c_1342_n 0.0218381f $X=9.825 $Y=2.595 $X2=0
+ $Y2=0
cc_726 N_SET_B_c_887_n N_A_1526_125#_c_1342_n 0.016173f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_727 SET_B N_A_1526_125#_c_1342_n 0.00199884f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_728 N_SET_B_c_892_n N_A_1526_125#_c_1342_n 0.00216661f $X=9.865 $Y=1.675
+ $X2=0 $Y2=0
cc_729 N_SET_B_c_894_n N_A_1526_125#_c_1342_n 0.0219324f $X=9.84 $Y=1.665 $X2=0
+ $Y2=0
cc_730 N_SET_B_M1033_g N_A_1526_125#_c_1343_n 0.0238716f $X=9.825 $Y=2.595 $X2=0
+ $Y2=0
cc_731 N_SET_B_M1033_g N_A_1526_125#_c_1345_n 0.0036057f $X=9.825 $Y=2.595 $X2=0
+ $Y2=0
cc_732 N_SET_B_c_885_n N_A_1526_125#_c_1333_n 0.00190545f $X=9.88 $Y=1.195 $X2=0
+ $Y2=0
cc_733 N_SET_B_c_887_n N_A_1526_125#_c_1336_n 0.00218913f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_734 N_SET_B_M1025_g N_VPWR_c_1573_n 0.00488986f $X=6.27 $Y=2.595 $X2=0 $Y2=0
cc_735 N_SET_B_M1033_g N_VPWR_c_1574_n 0.0108253f $X=9.825 $Y=2.595 $X2=0 $Y2=0
cc_736 N_SET_B_M1025_g N_VPWR_c_1581_n 0.00599858f $X=6.27 $Y=2.595 $X2=0 $Y2=0
cc_737 N_SET_B_M1033_g N_VPWR_c_1583_n 0.00938036f $X=9.825 $Y=2.595 $X2=0 $Y2=0
cc_738 N_SET_B_M1025_g N_VPWR_c_1568_n 0.00863224f $X=6.27 $Y=2.595 $X2=0 $Y2=0
cc_739 N_SET_B_M1033_g N_VPWR_c_1568_n 0.0180473f $X=9.825 $Y=2.595 $X2=0 $Y2=0
cc_740 N_SET_B_M1007_g N_VGND_c_1855_n 0.00141528f $X=6.595 $Y=0.835 $X2=0 $Y2=0
cc_741 N_SET_B_c_887_n N_VGND_c_1855_n 4.14819e-19 $X=9.695 $Y=1.665 $X2=0 $Y2=0
cc_742 N_SET_B_c_884_n N_VGND_c_1856_n 0.0135361f $X=9.385 $Y=1.12 $X2=0 $Y2=0
cc_743 N_SET_B_c_885_n N_VGND_c_1856_n 0.00613749f $X=9.88 $Y=1.195 $X2=0 $Y2=0
cc_744 N_SET_B_c_884_n N_VGND_c_1861_n 0.00345209f $X=9.385 $Y=1.12 $X2=0 $Y2=0
cc_745 N_SET_B_M1007_g N_VGND_c_1869_n 9.49986e-19 $X=6.595 $Y=0.835 $X2=0 $Y2=0
cc_746 N_SET_B_c_884_n N_VGND_c_1869_n 0.00394323f $X=9.385 $Y=1.12 $X2=0 $Y2=0
cc_747 N_A_266_409#_M1032_g N_A_1731_99#_c_1221_n 0.0219774f $X=8.34 $Y=0.835
+ $X2=0 $Y2=0
cc_748 N_A_266_409#_c_1028_n N_A_1731_99#_c_1223_n 0.0219774f $X=8.34 $Y=1.195
+ $X2=0 $Y2=0
cc_749 N_A_266_409#_c_1039_n N_A_1526_125#_c_1379_n 0.0195108f $X=7.605 $Y=2.02
+ $X2=0 $Y2=0
cc_750 N_A_266_409#_M1032_g N_A_1526_125#_c_1330_n 0.0117597f $X=8.34 $Y=0.835
+ $X2=0 $Y2=0
cc_751 N_A_266_409#_c_1039_n N_A_1526_125#_c_1340_n 7.95439e-19 $X=7.605 $Y=2.02
+ $X2=0 $Y2=0
cc_752 N_A_266_409#_c_1040_n N_A_1526_125#_c_1340_n 0.00320378f $X=7.99 $Y=1.945
+ $X2=0 $Y2=0
cc_753 N_A_266_409#_c_1023_n N_A_1526_125#_c_1331_n 0.00478169f $X=8.065 $Y=1.87
+ $X2=0 $Y2=0
cc_754 N_A_266_409#_c_1028_n N_A_1526_125#_c_1331_n 7.49766e-19 $X=8.34 $Y=1.195
+ $X2=0 $Y2=0
cc_755 N_A_266_409#_c_1021_n N_A_1526_125#_c_1336_n 0.00412547f $X=8.265 $Y=0.18
+ $X2=0 $Y2=0
cc_756 N_A_266_409#_M1032_g N_A_1526_125#_c_1336_n 0.00752936f $X=8.34 $Y=0.835
+ $X2=0 $Y2=0
cc_757 N_A_266_409#_c_1028_n N_A_1526_125#_c_1336_n 0.00873582f $X=8.34 $Y=1.195
+ $X2=0 $Y2=0
cc_758 N_A_266_409#_c_1045_n N_VPWR_M1029_d 0.00105617f $X=2.02 $Y=2.045 $X2=0
+ $Y2=0
cc_759 N_A_266_409#_c_1032_n N_VPWR_M1029_d 7.68583e-19 $X=2.31 $Y=1.68 $X2=0
+ $Y2=0
cc_760 N_A_266_409#_M1018_g N_VPWR_c_1571_n 0.0189086f $X=2.27 $Y=2.545 $X2=0
+ $Y2=0
cc_761 N_A_266_409#_c_1044_n N_VPWR_c_1571_n 0.0512146f $X=1.475 $Y=2.19 $X2=0
+ $Y2=0
cc_762 N_A_266_409#_c_1045_n N_VPWR_c_1571_n 0.00931009f $X=2.02 $Y=2.045 $X2=0
+ $Y2=0
cc_763 N_A_266_409#_c_1032_n N_VPWR_c_1571_n 0.00771383f $X=2.31 $Y=1.68 $X2=0
+ $Y2=0
cc_764 N_A_266_409#_M1026_g N_VPWR_c_1572_n 0.00107828f $X=4.28 $Y=2.595 $X2=0
+ $Y2=0
cc_765 N_A_266_409#_c_1039_n N_VPWR_c_1573_n 0.00386701f $X=7.605 $Y=2.02 $X2=0
+ $Y2=0
cc_766 N_A_266_409#_c_1044_n N_VPWR_c_1579_n 0.0321458f $X=1.475 $Y=2.19 $X2=0
+ $Y2=0
cc_767 N_A_266_409#_M1018_g N_VPWR_c_1580_n 0.00767656f $X=2.27 $Y=2.545 $X2=0
+ $Y2=0
cc_768 N_A_266_409#_M1026_g N_VPWR_c_1580_n 0.00599941f $X=4.28 $Y=2.595 $X2=0
+ $Y2=0
cc_769 N_A_266_409#_c_1039_n N_VPWR_c_1582_n 0.00975641f $X=7.605 $Y=2.02 $X2=0
+ $Y2=0
cc_770 N_A_266_409#_M1018_g N_VPWR_c_1568_n 0.014306f $X=2.27 $Y=2.545 $X2=0
+ $Y2=0
cc_771 N_A_266_409#_M1026_g N_VPWR_c_1568_n 0.00869224f $X=4.28 $Y=2.595 $X2=0
+ $Y2=0
cc_772 N_A_266_409#_c_1039_n N_VPWR_c_1568_n 0.017824f $X=7.605 $Y=2.02 $X2=0
+ $Y2=0
cc_773 N_A_266_409#_c_1044_n N_VPWR_c_1568_n 0.0183848f $X=1.475 $Y=2.19 $X2=0
+ $Y2=0
cc_774 N_A_266_409#_c_1044_n N_A_135_409#_c_1723_n 0.0768782f $X=1.475 $Y=2.19
+ $X2=0 $Y2=0
cc_775 N_A_266_409#_c_1030_n N_A_135_409#_c_1713_n 0.00570483f $X=1.575 $Y=1.1
+ $X2=0 $Y2=0
cc_776 N_A_266_409#_c_1031_n N_A_135_409#_c_1713_n 0.0214885f $X=1.575 $Y=0.8
+ $X2=0 $Y2=0
cc_777 N_A_266_409#_M1014_g N_A_135_409#_c_1714_n 6.77551e-19 $X=2.58 $Y=0.755
+ $X2=0 $Y2=0
cc_778 N_A_266_409#_c_1031_n N_A_135_409#_c_1714_n 0.032753f $X=1.575 $Y=0.8
+ $X2=0 $Y2=0
cc_779 N_A_266_409#_M1014_g N_A_135_409#_c_1715_n 0.0118405f $X=2.58 $Y=0.755
+ $X2=0 $Y2=0
cc_780 N_A_266_409#_M1011_g N_A_135_409#_c_1715_n 0.00730035f $X=2.94 $Y=0.755
+ $X2=0 $Y2=0
cc_781 N_A_266_409#_M1011_g N_A_135_409#_c_1716_n 0.00941082f $X=2.94 $Y=0.755
+ $X2=0 $Y2=0
cc_782 N_A_266_409#_c_1018_n N_A_135_409#_c_1716_n 0.00433613f $X=3.785 $Y=1.195
+ $X2=0 $Y2=0
cc_783 N_A_266_409#_M1028_g N_A_135_409#_c_1716_n 0.0123397f $X=3.89 $Y=0.835
+ $X2=0 $Y2=0
cc_784 N_A_266_409#_M1014_g N_A_135_409#_c_1717_n 8.25938e-19 $X=2.58 $Y=0.755
+ $X2=0 $Y2=0
cc_785 N_A_266_409#_M1018_g N_A_135_409#_c_1718_n 0.0035665f $X=2.27 $Y=2.545
+ $X2=0 $Y2=0
cc_786 N_A_266_409#_c_1015_n N_A_135_409#_c_1718_n 0.0103672f $X=2.58 $Y=1.515
+ $X2=0 $Y2=0
cc_787 N_A_266_409#_c_1032_n N_A_135_409#_c_1718_n 0.0207668f $X=2.31 $Y=1.68
+ $X2=0 $Y2=0
cc_788 N_A_266_409#_M1011_g N_A_135_409#_c_1719_n 0.00523599f $X=2.94 $Y=0.755
+ $X2=0 $Y2=0
cc_789 N_A_266_409#_c_1018_n N_A_135_409#_c_1719_n 0.00524184f $X=3.785 $Y=1.195
+ $X2=0 $Y2=0
cc_790 N_A_266_409#_M1028_g N_A_135_409#_c_1719_n 0.0155257f $X=3.89 $Y=0.835
+ $X2=0 $Y2=0
cc_791 N_A_266_409#_c_1029_n N_A_135_409#_c_1720_n 0.0498692f $X=1.245 $Y=1.96
+ $X2=0 $Y2=0
cc_792 N_A_266_409#_c_1030_n N_A_135_409#_c_1720_n 0.0134476f $X=1.575 $Y=1.1
+ $X2=0 $Y2=0
cc_793 N_A_266_409#_c_1031_n N_A_135_409#_c_1720_n 0.0156389f $X=1.575 $Y=0.8
+ $X2=0 $Y2=0
cc_794 N_A_266_409#_c_1046_n N_A_135_409#_c_1720_n 0.0141548f $X=1.4 $Y=2.045
+ $X2=0 $Y2=0
cc_795 N_A_266_409#_c_1030_n N_A_135_409#_c_1721_n 0.00255096f $X=1.575 $Y=1.1
+ $X2=0 $Y2=0
cc_796 N_A_266_409#_c_1031_n N_A_135_409#_c_1721_n 0.00844849f $X=1.575 $Y=0.8
+ $X2=0 $Y2=0
cc_797 N_A_266_409#_M1014_g N_A_135_409#_c_1722_n 0.00408844f $X=2.58 $Y=0.755
+ $X2=0 $Y2=0
cc_798 N_A_266_409#_c_1015_n N_A_135_409#_c_1722_n 0.0102576f $X=2.58 $Y=1.515
+ $X2=0 $Y2=0
cc_799 N_A_266_409#_c_1016_n N_A_135_409#_c_1722_n 0.0101385f $X=2.865 $Y=1.195
+ $X2=0 $Y2=0
cc_800 N_A_266_409#_M1011_g N_A_135_409#_c_1722_n 2.04434e-19 $X=2.94 $Y=0.755
+ $X2=0 $Y2=0
cc_801 N_A_266_409#_c_1025_n N_A_135_409#_c_1722_n 0.00450047f $X=2.58 $Y=1.195
+ $X2=0 $Y2=0
cc_802 N_A_266_409#_c_1026_n N_A_135_409#_c_1722_n 0.0106966f $X=2.94 $Y=1.195
+ $X2=0 $Y2=0
cc_803 N_A_266_409#_c_1030_n N_A_135_409#_c_1722_n 0.0131632f $X=1.575 $Y=1.1
+ $X2=0 $Y2=0
cc_804 N_A_266_409#_c_1032_n N_A_135_409#_c_1722_n 0.0345457f $X=2.31 $Y=1.68
+ $X2=0 $Y2=0
cc_805 N_A_266_409#_c_1033_n N_A_135_409#_c_1722_n 0.00320886f $X=2.58 $Y=1.68
+ $X2=0 $Y2=0
cc_806 N_A_266_409#_M1014_g N_VGND_c_1853_n 9.45515e-19 $X=2.58 $Y=0.755 $X2=0
+ $Y2=0
cc_807 N_A_266_409#_c_1021_n N_VGND_c_1854_n 0.0210961f $X=8.265 $Y=0.18 $X2=0
+ $Y2=0
cc_808 N_A_266_409#_c_1021_n N_VGND_c_1855_n 0.0261591f $X=8.265 $Y=0.18 $X2=0
+ $Y2=0
cc_809 N_A_266_409#_c_1021_n N_VGND_c_1861_n 0.0466671f $X=8.265 $Y=0.18 $X2=0
+ $Y2=0
cc_810 N_A_266_409#_M1014_g N_VGND_c_1865_n 0.00394144f $X=2.58 $Y=0.755 $X2=0
+ $Y2=0
cc_811 N_A_266_409#_M1011_g N_VGND_c_1865_n 6.46133e-19 $X=2.94 $Y=0.755 $X2=0
+ $Y2=0
cc_812 N_A_266_409#_c_1022_n N_VGND_c_1865_n 0.0365811f $X=3.965 $Y=0.18 $X2=0
+ $Y2=0
cc_813 N_A_266_409#_c_1021_n N_VGND_c_1866_n 0.0361813f $X=8.265 $Y=0.18 $X2=0
+ $Y2=0
cc_814 N_A_266_409#_M1014_g N_VGND_c_1869_n 0.00410091f $X=2.58 $Y=0.755 $X2=0
+ $Y2=0
cc_815 N_A_266_409#_c_1021_n N_VGND_c_1869_n 0.145439f $X=8.265 $Y=0.18 $X2=0
+ $Y2=0
cc_816 N_A_266_409#_c_1022_n N_VGND_c_1869_n 0.0106778f $X=3.965 $Y=0.18 $X2=0
+ $Y2=0
cc_817 N_A_1731_99#_c_1228_n N_A_1526_125#_c_1316_n 0.00940165f $X=10.23 $Y=0.47
+ $X2=0 $Y2=0
cc_818 N_A_1731_99#_c_1228_n N_A_1526_125#_c_1318_n 0.00941348f $X=10.23 $Y=0.47
+ $X2=0 $Y2=0
cc_819 N_A_1731_99#_c_1229_n N_A_1526_125#_c_1318_n 0.00949856f $X=10.57
+ $Y=1.245 $X2=0 $Y2=0
cc_820 N_A_1731_99#_c_1228_n N_A_1526_125#_c_1319_n 0.00145561f $X=10.23 $Y=0.47
+ $X2=0 $Y2=0
cc_821 N_A_1731_99#_c_1234_n N_A_1526_125#_M1034_g 9.82477e-19 $X=10.61 $Y=1.8
+ $X2=0 $Y2=0
cc_822 N_A_1731_99#_c_1230_n N_A_1526_125#_M1034_g 0.00414914f $X=10.61 $Y=1.675
+ $X2=0 $Y2=0
cc_823 N_A_1731_99#_c_1221_n N_A_1526_125#_c_1330_n 0.0150848f $X=8.73 $Y=1.12
+ $X2=0 $Y2=0
cc_824 N_A_1731_99#_c_1223_n N_A_1526_125#_c_1330_n 0.0011447f $X=8.995 $Y=1.195
+ $X2=0 $Y2=0
cc_825 N_A_1731_99#_c_1221_n N_A_1526_125#_c_1331_n 0.00148326f $X=8.73 $Y=1.12
+ $X2=0 $Y2=0
cc_826 N_A_1731_99#_c_1222_n N_A_1526_125#_c_1331_n 0.00734563f $X=8.995 $Y=1.51
+ $X2=0 $Y2=0
cc_827 N_A_1731_99#_M1000_g N_A_1526_125#_c_1331_n 0.00586296f $X=9.045 $Y=2.595
+ $X2=0 $Y2=0
cc_828 N_A_1731_99#_c_1223_n N_A_1526_125#_c_1331_n 0.0111124f $X=8.995 $Y=1.195
+ $X2=0 $Y2=0
cc_829 N_A_1731_99#_c_1224_n N_A_1526_125#_c_1331_n 0.0342885f $X=9.325 $Y=1.675
+ $X2=0 $Y2=0
cc_830 N_A_1731_99#_c_1225_n N_A_1526_125#_c_1331_n 0.007852f $X=9.325 $Y=1.675
+ $X2=0 $Y2=0
cc_831 N_A_1731_99#_c_1227_n N_A_1526_125#_c_1331_n 0.0131063f $X=9.49 $Y=1.245
+ $X2=0 $Y2=0
cc_832 N_A_1731_99#_M1000_g N_A_1526_125#_c_1342_n 0.0149933f $X=9.045 $Y=2.595
+ $X2=0 $Y2=0
cc_833 N_A_1731_99#_c_1224_n N_A_1526_125#_c_1342_n 0.0214493f $X=9.325 $Y=1.675
+ $X2=0 $Y2=0
cc_834 N_A_1731_99#_c_1225_n N_A_1526_125#_c_1342_n 0.00270418f $X=9.325
+ $Y=1.675 $X2=0 $Y2=0
cc_835 N_A_1731_99#_c_1235_n N_A_1526_125#_c_1342_n 0.011925f $X=10.65 $Y=1.84
+ $X2=0 $Y2=0
cc_836 N_A_1731_99#_c_1235_n N_A_1526_125#_c_1343_n 0.0346325f $X=10.65 $Y=1.84
+ $X2=0 $Y2=0
cc_837 N_A_1731_99#_c_1235_n N_A_1526_125#_c_1344_n 0.0187378f $X=10.65 $Y=1.84
+ $X2=0 $Y2=0
cc_838 N_A_1731_99#_c_1228_n N_A_1526_125#_c_1332_n 0.012792f $X=10.23 $Y=0.47
+ $X2=0 $Y2=0
cc_839 N_A_1731_99#_c_1229_n N_A_1526_125#_c_1332_n 0.0135689f $X=10.57 $Y=1.245
+ $X2=0 $Y2=0
cc_840 N_A_1731_99#_c_1228_n N_A_1526_125#_c_1333_n 0.00581911f $X=10.23 $Y=0.47
+ $X2=0 $Y2=0
cc_841 N_A_1731_99#_c_1229_n N_A_1526_125#_c_1333_n 0.00248465f $X=10.57
+ $Y=1.245 $X2=0 $Y2=0
cc_842 N_A_1731_99#_c_1230_n N_A_1526_125#_c_1333_n 0.00244423f $X=10.61
+ $Y=1.675 $X2=0 $Y2=0
cc_843 N_A_1731_99#_c_1230_n N_A_1526_125#_c_1334_n 0.0118405f $X=10.61 $Y=1.675
+ $X2=0 $Y2=0
cc_844 N_A_1731_99#_c_1234_n N_A_1526_125#_c_1335_n 0.0351227f $X=10.61 $Y=1.8
+ $X2=0 $Y2=0
cc_845 N_A_1731_99#_c_1230_n N_A_1526_125#_c_1335_n 0.00932725f $X=10.61
+ $Y=1.675 $X2=0 $Y2=0
cc_846 N_A_1731_99#_c_1221_n N_A_1526_125#_c_1336_n 0.00151671f $X=8.73 $Y=1.12
+ $X2=0 $Y2=0
cc_847 N_A_1731_99#_M1000_g N_A_1526_125#_c_1418_n 0.00778061f $X=9.045 $Y=2.595
+ $X2=0 $Y2=0
cc_848 N_A_1731_99#_M1000_g N_VPWR_c_1574_n 0.0209217f $X=9.045 $Y=2.595 $X2=0
+ $Y2=0
cc_849 N_A_1731_99#_M1000_g N_VPWR_c_1582_n 0.008763f $X=9.045 $Y=2.595 $X2=0
+ $Y2=0
cc_850 N_A_1731_99#_M1000_g N_VPWR_c_1568_n 0.0145916f $X=9.045 $Y=2.595 $X2=0
+ $Y2=0
cc_851 N_A_1731_99#_c_1221_n N_VGND_c_1856_n 0.00181462f $X=8.73 $Y=1.12 $X2=0
+ $Y2=0
cc_852 N_A_1731_99#_c_1226_n N_VGND_c_1856_n 0.0189292f $X=10.065 $Y=1.245 $X2=0
+ $Y2=0
cc_853 N_A_1731_99#_c_1227_n N_VGND_c_1856_n 0.00302164f $X=9.49 $Y=1.245 $X2=0
+ $Y2=0
cc_854 N_A_1731_99#_c_1228_n N_VGND_c_1856_n 0.0401567f $X=10.23 $Y=0.47 $X2=0
+ $Y2=0
cc_855 N_A_1731_99#_c_1228_n N_VGND_c_1857_n 0.0127138f $X=10.23 $Y=0.47 $X2=0
+ $Y2=0
cc_856 N_A_1731_99#_c_1221_n N_VGND_c_1861_n 0.00415323f $X=8.73 $Y=1.12 $X2=0
+ $Y2=0
cc_857 N_A_1731_99#_c_1228_n N_VGND_c_1863_n 0.0197885f $X=10.23 $Y=0.47 $X2=0
+ $Y2=0
cc_858 N_A_1731_99#_M1035_s N_VGND_c_1869_n 0.00232985f $X=10.085 $Y=0.235 $X2=0
+ $Y2=0
cc_859 N_A_1731_99#_c_1221_n N_VGND_c_1869_n 0.00469432f $X=8.73 $Y=1.12 $X2=0
+ $Y2=0
cc_860 N_A_1731_99#_c_1228_n N_VGND_c_1869_n 0.0125808f $X=10.23 $Y=0.47 $X2=0
+ $Y2=0
cc_861 N_A_1526_125#_M1003_g N_A_2287_74#_M1015_g 0.0325133f $X=12.155 $Y=0.58
+ $X2=0 $Y2=0
cc_862 N_A_1526_125#_M1016_g N_A_2287_74#_M1004_g 0.0163172f $X=12.175 $Y=2.37
+ $X2=0 $Y2=0
cc_863 N_A_1526_125#_M1016_g N_A_2287_74#_c_1499_n 0.0104943f $X=12.175 $Y=2.37
+ $X2=0 $Y2=0
cc_864 N_A_1526_125#_c_1321_n N_A_2287_74#_c_1500_n 0.00399207f $X=11.72 $Y=1.42
+ $X2=0 $Y2=0
cc_865 N_A_1526_125#_M1001_g N_A_2287_74#_c_1500_n 0.0196967f $X=11.795 $Y=0.58
+ $X2=0 $Y2=0
cc_866 N_A_1526_125#_M1003_g N_A_2287_74#_c_1500_n 0.00261832f $X=12.155 $Y=0.58
+ $X2=0 $Y2=0
cc_867 N_A_1526_125#_c_1326_n N_A_2287_74#_c_1500_n 0.00378827f $X=10.73 $Y=0.73
+ $X2=0 $Y2=0
cc_868 N_A_1526_125#_c_1328_n N_A_2287_74#_c_1500_n 0.00526771f $X=11.795
+ $Y=1.42 $X2=0 $Y2=0
cc_869 N_A_1526_125#_c_1332_n N_A_2287_74#_c_1500_n 0.0206128f $X=11 $Y=0.99
+ $X2=0 $Y2=0
cc_870 N_A_1526_125#_M1034_g N_A_2287_74#_c_1508_n 0.00142202f $X=10.915
+ $Y=2.195 $X2=0 $Y2=0
cc_871 N_A_1526_125#_M1016_g N_A_2287_74#_c_1508_n 0.0264529f $X=12.175 $Y=2.37
+ $X2=0 $Y2=0
cc_872 N_A_1526_125#_c_1335_n N_A_2287_74#_c_1508_n 4.76861e-19 $X=11 $Y=2.895
+ $X2=0 $Y2=0
cc_873 N_A_1526_125#_M1016_g N_A_2287_74#_c_1501_n 0.0140667f $X=12.175 $Y=2.37
+ $X2=0 $Y2=0
cc_874 N_A_1526_125#_c_1329_n N_A_2287_74#_c_1501_n 0.00958004f $X=12.175
+ $Y=1.42 $X2=0 $Y2=0
cc_875 N_A_1526_125#_M1003_g N_A_2287_74#_c_1502_n 0.00142287f $X=12.155 $Y=0.58
+ $X2=0 $Y2=0
cc_876 N_A_1526_125#_c_1329_n N_A_2287_74#_c_1502_n 7.32356e-19 $X=12.175
+ $Y=1.42 $X2=0 $Y2=0
cc_877 N_A_1526_125#_c_1329_n N_A_2287_74#_c_1503_n 0.0104943f $X=12.175 $Y=1.42
+ $X2=0 $Y2=0
cc_878 N_A_1526_125#_c_1319_n N_A_2287_74#_c_1504_n 0.00520156f $X=10.805
+ $Y=0.73 $X2=0 $Y2=0
cc_879 N_A_1526_125#_c_1321_n N_A_2287_74#_c_1504_n 0.00568129f $X=11.72 $Y=1.42
+ $X2=0 $Y2=0
cc_880 N_A_1526_125#_M1001_g N_A_2287_74#_c_1504_n 0.013155f $X=11.795 $Y=0.58
+ $X2=0 $Y2=0
cc_881 N_A_1526_125#_M1003_g N_A_2287_74#_c_1504_n 0.00151759f $X=12.155 $Y=0.58
+ $X2=0 $Y2=0
cc_882 N_A_1526_125#_M1034_g N_A_2287_74#_c_1505_n 9.65953e-19 $X=10.915
+ $Y=2.195 $X2=0 $Y2=0
cc_883 N_A_1526_125#_c_1321_n N_A_2287_74#_c_1505_n 7.3935e-19 $X=11.72 $Y=1.42
+ $X2=0 $Y2=0
cc_884 N_A_1526_125#_c_1323_n N_A_2287_74#_c_1505_n 0.0113571f $X=12.05 $Y=1.42
+ $X2=0 $Y2=0
cc_885 N_A_1526_125#_M1016_g N_A_2287_74#_c_1505_n 0.00381724f $X=12.175 $Y=2.37
+ $X2=0 $Y2=0
cc_886 N_A_1526_125#_c_1328_n N_A_2287_74#_c_1505_n 0.00410084f $X=11.795
+ $Y=1.42 $X2=0 $Y2=0
cc_887 N_A_1526_125#_c_1329_n N_A_2287_74#_c_1505_n 0.00129788f $X=12.175
+ $Y=1.42 $X2=0 $Y2=0
cc_888 N_A_1526_125#_c_1335_n N_A_2287_74#_c_1505_n 0.0056952f $X=11 $Y=2.895
+ $X2=0 $Y2=0
cc_889 N_A_1526_125#_c_1342_n N_VPWR_M1000_d 0.0100222f $X=9.925 $Y=2.105 $X2=0
+ $Y2=0
cc_890 N_A_1526_125#_c_1342_n N_VPWR_c_1574_n 0.0209601f $X=9.925 $Y=2.105 $X2=0
+ $Y2=0
cc_891 N_A_1526_125#_c_1343_n N_VPWR_c_1574_n 0.0191838f $X=10.09 $Y=2.24 $X2=0
+ $Y2=0
cc_892 N_A_1526_125#_c_1345_n N_VPWR_c_1574_n 0.00656934f $X=10.255 $Y=2.98
+ $X2=0 $Y2=0
cc_893 N_A_1526_125#_M1034_g N_VPWR_c_1575_n 0.0073647f $X=10.915 $Y=2.195 $X2=0
+ $Y2=0
cc_894 N_A_1526_125#_c_1321_n N_VPWR_c_1575_n 0.0100853f $X=11.72 $Y=1.42 $X2=0
+ $Y2=0
cc_895 N_A_1526_125#_M1016_g N_VPWR_c_1575_n 0.00488877f $X=12.175 $Y=2.37 $X2=0
+ $Y2=0
cc_896 N_A_1526_125#_c_1344_n N_VPWR_c_1575_n 0.0141601f $X=10.915 $Y=2.98 $X2=0
+ $Y2=0
cc_897 N_A_1526_125#_c_1335_n N_VPWR_c_1575_n 0.0531557f $X=11 $Y=2.895 $X2=0
+ $Y2=0
cc_898 N_A_1526_125#_M1016_g N_VPWR_c_1576_n 0.0257488f $X=12.175 $Y=2.37 $X2=0
+ $Y2=0
cc_899 N_A_1526_125#_M1016_g N_VPWR_c_1577_n 0.00747382f $X=12.175 $Y=2.37 $X2=0
+ $Y2=0
cc_900 N_A_1526_125#_c_1379_n N_VPWR_c_1582_n 0.0200085f $X=8.21 $Y=2.24 $X2=0
+ $Y2=0
cc_901 N_A_1526_125#_M1034_g N_VPWR_c_1583_n 5.77289e-19 $X=10.915 $Y=2.195
+ $X2=0 $Y2=0
cc_902 N_A_1526_125#_c_1344_n N_VPWR_c_1583_n 0.0513924f $X=10.915 $Y=2.98 $X2=0
+ $Y2=0
cc_903 N_A_1526_125#_c_1345_n N_VPWR_c_1583_n 0.0198894f $X=10.255 $Y=2.98 $X2=0
+ $Y2=0
cc_904 N_A_1526_125#_M1009_d N_VPWR_c_1568_n 0.0164864f $X=7.73 $Y=2.095 $X2=0
+ $Y2=0
cc_905 N_A_1526_125#_M1033_d N_VPWR_c_1568_n 0.0023218f $X=9.95 $Y=2.095 $X2=0
+ $Y2=0
cc_906 N_A_1526_125#_M1016_g N_VPWR_c_1568_n 0.00779694f $X=12.175 $Y=2.37 $X2=0
+ $Y2=0
cc_907 N_A_1526_125#_c_1379_n N_VPWR_c_1568_n 0.0126914f $X=8.21 $Y=2.24 $X2=0
+ $Y2=0
cc_908 N_A_1526_125#_c_1344_n N_VPWR_c_1568_n 0.0312303f $X=10.915 $Y=2.98 $X2=0
+ $Y2=0
cc_909 N_A_1526_125#_c_1345_n N_VPWR_c_1568_n 0.0125808f $X=10.255 $Y=2.98 $X2=0
+ $Y2=0
cc_910 N_A_1526_125#_c_1339_n A_1726_419# 0.00560887f $X=8.835 $Y=2.105
+ $X2=-0.19 $Y2=-0.245
cc_911 N_A_1526_125#_c_1418_n A_1726_419# 0.00126309f $X=8.92 $Y=2.105 $X2=-0.19
+ $Y2=-0.245
cc_912 N_A_1526_125#_M1016_g N_Q_c_1833_n 2.75707e-19 $X=12.175 $Y=2.37 $X2=0
+ $Y2=0
cc_913 N_A_1526_125#_c_1316_n N_VGND_c_1856_n 0.00397258f $X=10.445 $Y=0.73
+ $X2=0 $Y2=0
cc_914 N_A_1526_125#_c_1330_n N_VGND_c_1856_n 0.00344199f $X=8.835 $Y=0.98 $X2=0
+ $Y2=0
cc_915 N_A_1526_125#_c_1316_n N_VGND_c_1857_n 0.00231629f $X=10.445 $Y=0.73
+ $X2=0 $Y2=0
cc_916 N_A_1526_125#_c_1319_n N_VGND_c_1857_n 0.0132143f $X=10.805 $Y=0.73 $X2=0
+ $Y2=0
cc_917 N_A_1526_125#_M1001_g N_VGND_c_1857_n 0.00334229f $X=11.795 $Y=0.58 $X2=0
+ $Y2=0
cc_918 N_A_1526_125#_c_1326_n N_VGND_c_1857_n 0.0020268f $X=10.73 $Y=0.73 $X2=0
+ $Y2=0
cc_919 N_A_1526_125#_c_1332_n N_VGND_c_1857_n 0.0224559f $X=11 $Y=0.99 $X2=0
+ $Y2=0
cc_920 N_A_1526_125#_M1001_g N_VGND_c_1858_n 0.00173575f $X=11.795 $Y=0.58 $X2=0
+ $Y2=0
cc_921 N_A_1526_125#_M1003_g N_VGND_c_1858_n 0.0120445f $X=12.155 $Y=0.58 $X2=0
+ $Y2=0
cc_922 N_A_1526_125#_c_1329_n N_VGND_c_1858_n 0.00231283f $X=12.175 $Y=1.42
+ $X2=0 $Y2=0
cc_923 N_A_1526_125#_c_1336_n N_VGND_c_1861_n 0.00681209f $X=8.125 $Y=0.835
+ $X2=0 $Y2=0
cc_924 N_A_1526_125#_c_1316_n N_VGND_c_1863_n 0.00549284f $X=10.445 $Y=0.73
+ $X2=0 $Y2=0
cc_925 N_A_1526_125#_c_1317_n N_VGND_c_1863_n 4.87571e-19 $X=10.73 $Y=0.805
+ $X2=0 $Y2=0
cc_926 N_A_1526_125#_c_1319_n N_VGND_c_1863_n 0.00486043f $X=10.805 $Y=0.73
+ $X2=0 $Y2=0
cc_927 N_A_1526_125#_M1001_g N_VGND_c_1867_n 0.00297309f $X=11.795 $Y=0.58 $X2=0
+ $Y2=0
cc_928 N_A_1526_125#_M1003_g N_VGND_c_1867_n 0.00383152f $X=12.155 $Y=0.58 $X2=0
+ $Y2=0
cc_929 N_A_1526_125#_c_1316_n N_VGND_c_1869_n 0.0112805f $X=10.445 $Y=0.73 $X2=0
+ $Y2=0
cc_930 N_A_1526_125#_c_1317_n N_VGND_c_1869_n 6.51792e-19 $X=10.73 $Y=0.805
+ $X2=0 $Y2=0
cc_931 N_A_1526_125#_c_1319_n N_VGND_c_1869_n 0.00754596f $X=10.805 $Y=0.73
+ $X2=0 $Y2=0
cc_932 N_A_1526_125#_M1001_g N_VGND_c_1869_n 0.0038076f $X=11.795 $Y=0.58 $X2=0
+ $Y2=0
cc_933 N_A_1526_125#_M1003_g N_VGND_c_1869_n 0.00756787f $X=12.155 $Y=0.58 $X2=0
+ $Y2=0
cc_934 N_A_1526_125#_c_1332_n N_VGND_c_1869_n 0.00170501f $X=11 $Y=0.99 $X2=0
+ $Y2=0
cc_935 N_A_1526_125#_c_1336_n N_VGND_c_1869_n 0.00865577f $X=8.125 $Y=0.835
+ $X2=0 $Y2=0
cc_936 N_A_1526_125#_c_1330_n A_1683_125# 0.0048076f $X=8.835 $Y=0.98 $X2=-0.19
+ $Y2=-0.245
cc_937 N_A_1526_125#_c_1330_n A_1761_125# 0.00864867f $X=8.835 $Y=0.98 $X2=-0.19
+ $Y2=-0.245
cc_938 N_A_2287_74#_c_1508_n N_VPWR_c_1575_n 0.096225f $X=11.91 $Y=2.015 $X2=0
+ $Y2=0
cc_939 N_A_2287_74#_M1004_g N_VPWR_c_1576_n 0.0257478f $X=12.705 $Y=2.37 $X2=0
+ $Y2=0
cc_940 N_A_2287_74#_c_1499_n N_VPWR_c_1576_n 5.39992e-19 $X=12.675 $Y=1.66 $X2=0
+ $Y2=0
cc_941 N_A_2287_74#_c_1508_n N_VPWR_c_1576_n 0.0692741f $X=11.91 $Y=2.015 $X2=0
+ $Y2=0
cc_942 N_A_2287_74#_c_1501_n N_VPWR_c_1576_n 0.025615f $X=12.51 $Y=1.575 $X2=0
+ $Y2=0
cc_943 N_A_2287_74#_c_1508_n N_VPWR_c_1577_n 0.0122968f $X=11.91 $Y=2.015 $X2=0
+ $Y2=0
cc_944 N_A_2287_74#_M1004_g N_VPWR_c_1584_n 0.00747382f $X=12.705 $Y=2.37 $X2=0
+ $Y2=0
cc_945 N_A_2287_74#_M1004_g N_VPWR_c_1568_n 0.00779694f $X=12.705 $Y=2.37 $X2=0
+ $Y2=0
cc_946 N_A_2287_74#_c_1508_n N_VPWR_c_1568_n 0.0131561f $X=11.91 $Y=2.015 $X2=0
+ $Y2=0
cc_947 N_A_2287_74#_M1015_g Q 0.00125204f $X=12.585 $Y=0.58 $X2=0 $Y2=0
cc_948 N_A_2287_74#_M1006_g Q 0.0100639f $X=12.945 $Y=0.58 $X2=0 $Y2=0
cc_949 N_A_2287_74#_M1004_g Q 0.00651453f $X=12.705 $Y=2.37 $X2=0 $Y2=0
cc_950 N_A_2287_74#_M1006_g Q 0.0115307f $X=12.945 $Y=0.58 $X2=0 $Y2=0
cc_951 N_A_2287_74#_c_1501_n Q 0.0105477f $X=12.51 $Y=1.575 $X2=0 $Y2=0
cc_952 N_A_2287_74#_c_1502_n Q 0.029316f $X=12.675 $Y=1.155 $X2=0 $Y2=0
cc_953 N_A_2287_74#_c_1503_n Q 0.00865955f $X=12.675 $Y=1.155 $X2=0 $Y2=0
cc_954 N_A_2287_74#_M1004_g Q 0.0139894f $X=12.705 $Y=2.37 $X2=0 $Y2=0
cc_955 N_A_2287_74#_M1004_g N_Q_c_1833_n 0.00522616f $X=12.705 $Y=2.37 $X2=0
+ $Y2=0
cc_956 N_A_2287_74#_c_1501_n N_Q_c_1833_n 0.002673f $X=12.51 $Y=1.575 $X2=0
+ $Y2=0
cc_957 N_A_2287_74#_c_1504_n N_VGND_c_1857_n 0.0203649f $X=11.78 $Y=0.58 $X2=0
+ $Y2=0
cc_958 N_A_2287_74#_M1015_g N_VGND_c_1858_n 0.0121853f $X=12.585 $Y=0.58 $X2=0
+ $Y2=0
cc_959 N_A_2287_74#_M1006_g N_VGND_c_1858_n 0.00182089f $X=12.945 $Y=0.58 $X2=0
+ $Y2=0
cc_960 N_A_2287_74#_c_1502_n N_VGND_c_1858_n 0.00185662f $X=12.675 $Y=1.155
+ $X2=0 $Y2=0
cc_961 N_A_2287_74#_c_1504_n N_VGND_c_1858_n 0.0202525f $X=11.78 $Y=0.58 $X2=0
+ $Y2=0
cc_962 N_A_2287_74#_c_1504_n N_VGND_c_1867_n 0.0190286f $X=11.78 $Y=0.58 $X2=0
+ $Y2=0
cc_963 N_A_2287_74#_M1015_g N_VGND_c_1868_n 0.00383152f $X=12.585 $Y=0.58 $X2=0
+ $Y2=0
cc_964 N_A_2287_74#_M1006_g N_VGND_c_1868_n 0.00434272f $X=12.945 $Y=0.58 $X2=0
+ $Y2=0
cc_965 N_A_2287_74#_M1015_g N_VGND_c_1869_n 0.00756787f $X=12.585 $Y=0.58 $X2=0
+ $Y2=0
cc_966 N_A_2287_74#_M1006_g N_VGND_c_1869_n 0.00824175f $X=12.945 $Y=0.58 $X2=0
+ $Y2=0
cc_967 N_A_2287_74#_c_1504_n N_VGND_c_1869_n 0.0156955f $X=11.78 $Y=0.58 $X2=0
+ $Y2=0
cc_968 N_VPWR_c_1568_n N_A_135_409#_M1021_s 0.00233022f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_969 N_VPWR_c_1570_n N_A_135_409#_c_1723_n 0.0684934f $X=0.285 $Y=2.19 $X2=0
+ $Y2=0
cc_970 N_VPWR_c_1579_n N_A_135_409#_c_1724_n 0.0220321f $X=1.84 $Y=3.33 $X2=0
+ $Y2=0
cc_971 N_VPWR_c_1568_n N_A_135_409#_c_1724_n 0.0125808f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_972 N_VPWR_c_1568_n A_881_419# 0.00249606f $X=13.2 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_973 N_VPWR_c_1568_n A_1448_419# 0.010279f $X=13.2 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_974 N_VPWR_c_1568_n A_1726_419# 0.0124205f $X=13.2 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_975 N_VPWR_c_1584_n Q 0.0168747f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_976 N_VPWR_c_1568_n Q 0.0180375f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_977 N_VPWR_c_1576_n N_Q_c_1833_n 0.0709584f $X=12.44 $Y=2.015 $X2=0 $Y2=0
cc_978 N_A_135_409#_c_1721_n N_VGND_c_1852_n 0.0181655f $X=1.012 $Y=0.35 $X2=0
+ $Y2=0
cc_979 N_A_135_409#_c_1713_n N_VGND_c_1853_n 0.0136958f $X=1.93 $Y=0.35 $X2=0
+ $Y2=0
cc_980 N_A_135_409#_c_1714_n N_VGND_c_1853_n 0.0196067f $X=2.015 $Y=1.1 $X2=0
+ $Y2=0
cc_981 N_A_135_409#_c_1715_n N_VGND_c_1853_n 0.0196067f $X=2.715 $Y=1.1 $X2=0
+ $Y2=0
cc_982 N_A_135_409#_c_1717_n N_VGND_c_1853_n 0.0136958f $X=2.8 $Y=0.35 $X2=0
+ $Y2=0
cc_983 N_A_135_409#_c_1722_n N_VGND_c_1853_n 0.0136087f $X=2.715 $Y=1.217 $X2=0
+ $Y2=0
cc_984 N_A_135_409#_c_1713_n N_VGND_c_1859_n 0.0547886f $X=1.93 $Y=0.35 $X2=0
+ $Y2=0
cc_985 N_A_135_409#_c_1721_n N_VGND_c_1859_n 0.0263762f $X=1.012 $Y=0.35 $X2=0
+ $Y2=0
cc_986 N_A_135_409#_c_1716_n N_VGND_c_1865_n 0.0651594f $X=3.51 $Y=0.35 $X2=0
+ $Y2=0
cc_987 N_A_135_409#_c_1717_n N_VGND_c_1865_n 0.0114622f $X=2.8 $Y=0.35 $X2=0
+ $Y2=0
cc_988 N_A_135_409#_c_1713_n N_VGND_c_1869_n 0.0332955f $X=1.93 $Y=0.35 $X2=0
+ $Y2=0
cc_989 N_A_135_409#_c_1716_n N_VGND_c_1869_n 0.0391802f $X=3.51 $Y=0.35 $X2=0
+ $Y2=0
cc_990 N_A_135_409#_c_1717_n N_VGND_c_1869_n 0.00657784f $X=2.8 $Y=0.35 $X2=0
+ $Y2=0
cc_991 N_A_135_409#_c_1721_n N_VGND_c_1869_n 0.015044f $X=1.012 $Y=0.35 $X2=0
+ $Y2=0
cc_992 N_A_135_409#_c_1714_n A_373_109# 0.00374559f $X=2.015 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_993 N_A_135_409#_c_1715_n A_531_109# 0.00374559f $X=2.715 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_994 Q N_VGND_c_1858_n 0.0153904f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_995 Q N_VGND_c_1868_n 0.0144575f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_996 Q N_VGND_c_1869_n 0.0119563f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_997 N_VGND_c_1869_n A_2104_47# 0.00829524f $X=13.2 $Y=0 $X2=-0.19 $Y2=-0.245
