* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21boi_lp A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_513_47# B1_N a_298_318# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_172_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A1 a_29_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 Y a_298_318# a_336_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND B1_N a_513_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND A2 a_172_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_336_47# a_298_318# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_29_409# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VPWR B1_N a_298_318# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_29_409# a_298_318# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
