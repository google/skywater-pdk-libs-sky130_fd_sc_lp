* File: sky130_fd_sc_lp__nand4bb_4.pex.spice
* Created: Fri Aug 28 10:52:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%A_N 3 6 8 9 13 15
c30 15 0 6.64596e-20 $X=0.53 $Y=1.295
c31 6 0 9.81071e-20 $X=0.58 $Y=2.465
r32 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.46
+ $X2=0.53 $Y2=1.625
r33 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.46
+ $X2=0.53 $Y2=1.295
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.46 $X2=0.53 $Y2=1.46
r35 9 14 5.62502 $w=4.18e-07 $l=2.05e-07 $layer=LI1_cond $X=0.655 $Y=1.665
+ $X2=0.655 $Y2=1.46
r36 8 14 4.52745 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=0.655 $Y=1.295
+ $X2=0.655 $Y2=1.46
r37 6 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.58 $Y=2.465
+ $X2=0.58 $Y2=1.625
r38 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.58 $Y=0.765
+ $X2=0.58 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%B_N 1 3 6 8 9 15
c33 8 0 1.64567e-19 $X=1.2 $Y=1.295
r34 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.46 $X2=1.2 $Y2=1.46
r35 12 15 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.01 $Y=1.46 $X2=1.2
+ $Y2=1.46
r36 9 16 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.16 $Y=1.665
+ $X2=1.16 $Y2=1.46
r37 8 16 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=1.295
+ $X2=1.16 $Y2=1.46
r38 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.625
+ $X2=1.01 $Y2=1.46
r39 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.01 $Y=1.625 $X2=1.01
+ $Y2=2.465
r40 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.295
+ $X2=1.01 $Y2=1.46
r41 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.01 $Y=1.295 $X2=1.01
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%A_44_69# 1 2 9 13 17 21 25 29 33 37 41 46
+ 49 52 53 58 61 63 64 66 75
r117 75 76 4.43558 $w=3.26e-07 $l=3e-08 $layer=POLY_cond $X=3.515 $Y=1.51
+ $X2=3.545 $Y2=1.51
r118 72 73 4.43558 $w=3.26e-07 $l=3e-08 $layer=POLY_cond $X=3.085 $Y=1.51
+ $X2=3.115 $Y2=1.51
r119 71 72 63.5767 $w=3.26e-07 $l=4.3e-07 $layer=POLY_cond $X=2.655 $Y=1.51
+ $X2=3.085 $Y2=1.51
r120 70 71 19.2209 $w=3.26e-07 $l=1.3e-07 $layer=POLY_cond $X=2.525 $Y=1.51
+ $X2=2.655 $Y2=1.51
r121 69 70 44.3558 $w=3.26e-07 $l=3e-07 $layer=POLY_cond $X=2.225 $Y=1.51
+ $X2=2.525 $Y2=1.51
r122 63 64 7.84768 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.267 $Y=2.095
+ $X2=0.267 $Y2=1.93
r123 61 64 51.9522 $w=1.88e-07 $l=8.9e-07 $layer=LI1_cond $X=0.18 $Y=1.04
+ $X2=0.18 $Y2=1.93
r124 59 75 50.2699 $w=3.26e-07 $l=3.4e-07 $layer=POLY_cond $X=3.175 $Y=1.51
+ $X2=3.515 $Y2=1.51
r125 59 73 8.87117 $w=3.26e-07 $l=6e-08 $layer=POLY_cond $X=3.175 $Y=1.51
+ $X2=3.115 $Y2=1.51
r126 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.175
+ $Y=1.51 $X2=3.175 $Y2=1.51
r127 56 69 10.3497 $w=3.26e-07 $l=7e-08 $layer=POLY_cond $X=2.155 $Y=1.51
+ $X2=2.225 $Y2=1.51
r128 56 67 8.87117 $w=3.26e-07 $l=6e-08 $layer=POLY_cond $X=2.155 $Y=1.51
+ $X2=2.095 $Y2=1.51
r129 55 58 53.4314 $w=2.18e-07 $l=1.02e-06 $layer=LI1_cond $X=2.155 $Y=1.495
+ $X2=3.175 $Y2=1.495
r130 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.155
+ $Y=1.51 $X2=2.155 $Y2=1.51
r131 53 55 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=2.02 $Y=1.495
+ $X2=2.155 $Y2=1.495
r132 51 53 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.935 $Y=1.605
+ $X2=2.02 $Y2=1.495
r133 51 52 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.935 $Y=1.605
+ $X2=1.935 $Y2=2.34
r134 50 66 4.19346 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.45 $Y=2.425
+ $X2=0.267 $Y2=2.425
r135 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.85 $Y=2.425
+ $X2=1.935 $Y2=2.34
r136 49 50 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.85 $Y=2.425
+ $X2=0.45 $Y2=2.425
r137 46 66 2.63236 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.267 $Y=2.34
+ $X2=0.267 $Y2=2.425
r138 45 63 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=0.267 $Y=2.112
+ $X2=0.267 $Y2=2.095
r139 45 46 7.19882 $w=3.63e-07 $l=2.28e-07 $layer=LI1_cond $X=0.267 $Y=2.112
+ $X2=0.267 $Y2=2.34
r140 39 61 8.5462 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=0.272 $Y=0.853
+ $X2=0.272 $Y2=1.04
r141 39 41 11.1556 $w=3.73e-07 $l=3.63e-07 $layer=LI1_cond $X=0.272 $Y=0.853
+ $X2=0.272 $Y2=0.49
r142 35 76 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.545 $Y=1.345
+ $X2=3.545 $Y2=1.51
r143 35 37 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.545 $Y=1.345
+ $X2=3.545 $Y2=0.755
r144 31 75 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.515 $Y=1.675
+ $X2=3.515 $Y2=1.51
r145 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.515 $Y=1.675
+ $X2=3.515 $Y2=2.465
r146 27 73 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.345
+ $X2=3.115 $Y2=1.51
r147 27 29 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.115 $Y=1.345
+ $X2=3.115 $Y2=0.755
r148 23 72 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.675
+ $X2=3.085 $Y2=1.51
r149 23 25 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.085 $Y=1.675
+ $X2=3.085 $Y2=2.465
r150 19 71 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.675
+ $X2=2.655 $Y2=1.51
r151 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.655 $Y=1.675
+ $X2=2.655 $Y2=2.465
r152 15 70 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.525 $Y=1.345
+ $X2=2.525 $Y2=1.51
r153 15 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.525 $Y=1.345
+ $X2=2.525 $Y2=0.755
r154 11 69 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.675
+ $X2=2.225 $Y2=1.51
r155 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.225 $Y=1.675
+ $X2=2.225 $Y2=2.465
r156 7 67 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.345
+ $X2=2.095 $Y2=1.51
r157 7 9 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.095 $Y=1.345
+ $X2=2.095 $Y2=0.755
r158 2 66 300 $w=1.7e-07 $l=6.59545e-07 $layer=licon1_PDIFF $count=2 $X=0.24
+ $Y=1.835 $X2=0.365 $Y2=2.435
r159 2 63 600 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.24
+ $Y=1.835 $X2=0.365 $Y2=2.095
r160 1 41 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.22
+ $Y=0.345 $X2=0.345 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%A_217_69# 1 2 9 13 17 21 25 29 33 37 39 45
+ 48 49 50 52 55 56 63
c142 56 0 1.72165e-19 $X=5.735 $Y=1.5
c143 55 0 1.21283e-19 $X=5.735 $Y=1.5
c144 37 0 5.86634e-20 $X=5.425 $Y=0.755
c145 21 0 1.51661e-19 $X=4.565 $Y=0.755
r146 74 75 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=5.235 $Y=1.5
+ $X2=5.425 $Y2=1.5
r147 73 74 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.995 $Y=1.5
+ $X2=5.235 $Y2=1.5
r148 72 73 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.805 $Y=1.5
+ $X2=4.995 $Y2=1.5
r149 71 72 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.565 $Y=1.5
+ $X2=4.805 $Y2=1.5
r150 70 71 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.375 $Y=1.5
+ $X2=4.565 $Y2=1.5
r151 69 70 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.135 $Y=1.5
+ $X2=4.375 $Y2=1.5
r152 63 75 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.5 $Y=1.5
+ $X2=5.425 $Y2=1.5
r153 62 69 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.035 $Y=1.5
+ $X2=4.135 $Y2=1.5
r154 62 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.035 $Y=1.5
+ $X2=3.945 $Y2=1.5
r155 61 62 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=4.035
+ $Y=1.5 $X2=4.035 $Y2=1.5
r156 56 63 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=5.735 $Y=1.5
+ $X2=5.5 $Y2=1.5
r157 55 56 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=5.735
+ $Y=1.5 $X2=5.735 $Y2=1.5
r158 53 61 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=1.51
+ $X2=3.955 $Y2=1.51
r159 53 55 98.9426 $w=1.88e-07 $l=1.695e-06 $layer=LI1_cond $X=4.04 $Y=1.51
+ $X2=5.735 $Y2=1.51
r160 52 61 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.955 $Y=1.415
+ $X2=3.955 $Y2=1.51
r161 51 52 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.955 $Y=0.785
+ $X2=3.955 $Y2=1.415
r162 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.87 $Y=0.7
+ $X2=3.955 $Y2=0.785
r163 49 50 142.877 $w=1.68e-07 $l=2.19e-06 $layer=LI1_cond $X=3.87 $Y=0.7
+ $X2=1.68 $Y2=0.7
r164 47 50 5.69269 $w=2.62e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.59 $Y=0.785
+ $X2=1.68 $Y2=0.7
r165 47 58 16.7634 $w=2.62e-07 $l=3.6e-07 $layer=LI1_cond $X=1.59 $Y=0.785
+ $X2=1.23 $Y2=0.785
r166 47 48 69.9343 $w=1.78e-07 $l=1.135e-06 $layer=LI1_cond $X=1.59 $Y=0.785
+ $X2=1.59 $Y2=1.92
r167 43 58 2.32089 $w=2e-07 $l=1.7e-07 $layer=LI1_cond $X=1.23 $Y=0.615 $X2=1.23
+ $Y2=0.785
r168 43 45 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=1.23 $Y=0.615
+ $X2=1.23 $Y2=0.49
r169 39 48 7.0541 $w=2.5e-07 $l=1.63936e-07 $layer=LI1_cond $X=1.5 $Y=2.045
+ $X2=1.59 $Y2=1.92
r170 39 41 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=1.5 $Y=2.045
+ $X2=1.225 $Y2=2.045
r171 35 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.425 $Y=1.335
+ $X2=5.425 $Y2=1.5
r172 35 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.425 $Y=1.335
+ $X2=5.425 $Y2=0.755
r173 31 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.235 $Y=1.665
+ $X2=5.235 $Y2=1.5
r174 31 33 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.235 $Y=1.665
+ $X2=5.235 $Y2=2.465
r175 27 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.995 $Y=1.335
+ $X2=4.995 $Y2=1.5
r176 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.995 $Y=1.335
+ $X2=4.995 $Y2=0.755
r177 23 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.805 $Y=1.665
+ $X2=4.805 $Y2=1.5
r178 23 25 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.805 $Y=1.665
+ $X2=4.805 $Y2=2.465
r179 19 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.565 $Y=1.335
+ $X2=4.565 $Y2=1.5
r180 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.565 $Y=1.335
+ $X2=4.565 $Y2=0.755
r181 15 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.665
+ $X2=4.375 $Y2=1.5
r182 15 17 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.375 $Y=1.665
+ $X2=4.375 $Y2=2.465
r183 11 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.135 $Y=1.335
+ $X2=4.135 $Y2=1.5
r184 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.135 $Y=1.335
+ $X2=4.135 $Y2=0.755
r185 7 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.665
+ $X2=3.945 $Y2=1.5
r186 7 9 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.945 $Y=1.665
+ $X2=3.945 $Y2=2.465
r187 2 41 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.225 $Y2=2.045
r188 1 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.345 $X2=1.225 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%C 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 51
c79 51 0 1.21283e-19 $X=7.885 $Y=1.35
r80 50 51 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=7.855 $Y=1.35
+ $X2=7.885 $Y2=1.35
r81 48 50 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=7.795 $Y=1.35
+ $X2=7.855 $Y2=1.35
r82 48 49 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=7.795
+ $Y=1.35 $X2=7.795 $Y2=1.35
r83 46 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.455 $Y=1.35
+ $X2=7.795 $Y2=1.35
r84 45 46 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=7.425 $Y=1.35
+ $X2=7.455 $Y2=1.35
r85 44 45 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=7.025 $Y=1.35
+ $X2=7.425 $Y2=1.35
r86 43 44 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.995 $Y=1.35
+ $X2=7.025 $Y2=1.35
r87 42 43 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=6.595 $Y=1.35
+ $X2=6.995 $Y2=1.35
r88 41 42 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.565 $Y=1.35
+ $X2=6.595 $Y2=1.35
r89 38 41 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=6.435 $Y=1.35
+ $X2=6.565 $Y2=1.35
r90 32 49 4.57319 $w=3.13e-07 $l=1.25e-07 $layer=LI1_cond $X=7.92 $Y=1.357
+ $X2=7.795 $Y2=1.357
r91 31 49 12.9878 $w=3.13e-07 $l=3.55e-07 $layer=LI1_cond $X=7.44 $Y=1.357
+ $X2=7.795 $Y2=1.357
r92 30 31 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.357
+ $X2=7.44 $Y2=1.357
r93 29 30 19.2074 $w=3.13e-07 $l=5.25e-07 $layer=LI1_cond $X=6.435 $Y=1.357
+ $X2=6.96 $Y2=1.357
r94 29 38 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.435
+ $Y=1.35 $X2=6.435 $Y2=1.35
r95 26 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.885 $Y=1.185
+ $X2=7.885 $Y2=1.35
r96 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.885 $Y=1.185
+ $X2=7.885 $Y2=0.655
r97 22 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.855 $Y=1.515
+ $X2=7.855 $Y2=1.35
r98 22 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.855 $Y=1.515
+ $X2=7.855 $Y2=2.465
r99 19 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.455 $Y=1.185
+ $X2=7.455 $Y2=1.35
r100 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.455 $Y=1.185
+ $X2=7.455 $Y2=0.655
r101 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.425 $Y=1.515
+ $X2=7.425 $Y2=1.35
r102 15 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.425 $Y=1.515
+ $X2=7.425 $Y2=2.465
r103 12 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.185
+ $X2=7.025 $Y2=1.35
r104 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.025 $Y=1.185
+ $X2=7.025 $Y2=0.655
r105 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.995 $Y=1.515
+ $X2=6.995 $Y2=1.35
r106 8 10 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.995 $Y=1.515
+ $X2=6.995 $Y2=2.465
r107 5 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.185
+ $X2=6.595 $Y2=1.35
r108 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.595 $Y=1.185
+ $X2=6.595 $Y2=0.655
r109 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.565 $Y=1.515
+ $X2=6.565 $Y2=1.35
r110 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.565 $Y=1.515
+ $X2=6.565 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%D 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 50
r70 50 51 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.735
+ $Y=1.35 $X2=9.735 $Y2=1.35
r71 48 50 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=9.605 $Y=1.35
+ $X2=9.735 $Y2=1.35
r72 47 48 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=9.575 $Y=1.35
+ $X2=9.605 $Y2=1.35
r73 46 47 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=9.175 $Y=1.35
+ $X2=9.575 $Y2=1.35
r74 45 46 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=9.145 $Y=1.35
+ $X2=9.175 $Y2=1.35
r75 44 45 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=8.745 $Y=1.35
+ $X2=9.145 $Y2=1.35
r76 43 44 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=8.715 $Y=1.35
+ $X2=8.745 $Y2=1.35
r77 41 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.375 $Y=1.35
+ $X2=8.715 $Y2=1.35
r78 39 41 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.315 $Y=1.35
+ $X2=8.375 $Y2=1.35
r79 37 39 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=8.285 $Y=1.35
+ $X2=8.315 $Y2=1.35
r80 32 51 3.84148 $w=3.13e-07 $l=1.05e-07 $layer=LI1_cond $X=9.84 $Y=1.357
+ $X2=9.735 $Y2=1.357
r81 31 51 13.7196 $w=3.13e-07 $l=3.75e-07 $layer=LI1_cond $X=9.36 $Y=1.357
+ $X2=9.735 $Y2=1.357
r82 30 31 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.357
+ $X2=9.36 $Y2=1.357
r83 29 30 18.4757 $w=3.13e-07 $l=5.05e-07 $layer=LI1_cond $X=8.375 $Y=1.357
+ $X2=8.88 $Y2=1.357
r84 29 41 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.375
+ $Y=1.35 $X2=8.375 $Y2=1.35
r85 26 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.605 $Y=1.185
+ $X2=9.605 $Y2=1.35
r86 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.605 $Y=1.185
+ $X2=9.605 $Y2=0.655
r87 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.575 $Y=1.515
+ $X2=9.575 $Y2=1.35
r88 22 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.575 $Y=1.515
+ $X2=9.575 $Y2=2.465
r89 19 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.175 $Y=1.185
+ $X2=9.175 $Y2=1.35
r90 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.175 $Y=1.185
+ $X2=9.175 $Y2=0.655
r91 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.145 $Y=1.515
+ $X2=9.145 $Y2=1.35
r92 15 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.145 $Y=1.515
+ $X2=9.145 $Y2=2.465
r93 12 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.745 $Y=1.185
+ $X2=8.745 $Y2=1.35
r94 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.745 $Y=1.185
+ $X2=8.745 $Y2=0.655
r95 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.715 $Y=1.515
+ $X2=8.715 $Y2=1.35
r96 8 10 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.715 $Y=1.515
+ $X2=8.715 $Y2=2.465
r97 5 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.315 $Y=1.185
+ $X2=8.315 $Y2=1.35
r98 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.315 $Y=1.185
+ $X2=8.315 $Y2=0.655
r99 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.285 $Y=1.515
+ $X2=8.285 $Y2=1.35
r100 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.285 $Y=1.515
+ $X2=8.285 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49
+ 55 59 63 67 73 77 79 84 85 86 87 88 89 90 92 104 109 118 123 129 132 135 144
+ 147 150 154
r151 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r152 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r153 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r154 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r155 142 144 4.24348 $w=1.035e-06 $l=3.6e-07 $layer=LI1_cond $X=5.88 $Y=2.97
+ $X2=5.88 $Y2=3.33
r156 140 142 6.54203 $w=1.035e-06 $l=5.55e-07 $layer=LI1_cond $X=5.88 $Y=2.415
+ $X2=5.88 $Y2=2.97
r157 138 140 1.47343 $w=1.035e-06 $l=5.28819e-07 $layer=LI1_cond $X=6.35 $Y=2.29
+ $X2=5.88 $Y2=2.415
r158 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r159 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r160 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r161 127 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r162 127 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r163 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r164 124 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.095 $Y=3.33
+ $X2=8.93 $Y2=3.33
r165 124 126 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.095 $Y=3.33
+ $X2=9.36 $Y2=3.33
r166 123 153 4.4394 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=9.655 $Y=3.33
+ $X2=9.867 $Y2=3.33
r167 123 126 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.655 $Y=3.33
+ $X2=9.36 $Y2=3.33
r168 122 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r169 122 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r170 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r171 119 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=8.07 $Y2=3.33
r172 119 121 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=8.4 $Y2=3.33
r173 118 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.765 $Y=3.33
+ $X2=8.93 $Y2=3.33
r174 118 121 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.765 $Y=3.33
+ $X2=8.4 $Y2=3.33
r175 117 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r176 117 145 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6 $Y2=3.33
r177 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r178 114 144 11.9616 $w=1.7e-07 $l=5.95e-07 $layer=LI1_cond $X=6.475 $Y=3.33
+ $X2=5.88 $Y2=3.33
r179 114 116 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.475 $Y=3.33
+ $X2=6.96 $Y2=3.33
r180 110 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=3.33
+ $X2=4.59 $Y2=3.33
r181 110 112 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.755 $Y=3.33
+ $X2=5.04 $Y2=3.33
r182 109 144 11.9616 $w=1.7e-07 $l=5.95e-07 $layer=LI1_cond $X=5.285 $Y=3.33
+ $X2=5.88 $Y2=3.33
r183 109 112 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.285 $Y=3.33
+ $X2=5.04 $Y2=3.33
r184 108 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r185 108 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r186 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r187 105 132 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=3.71 $Y2=3.33
r188 105 107 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=4.08 $Y2=3.33
r189 104 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.59 $Y2=3.33
r190 104 107 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r191 103 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r192 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r193 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r194 100 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r196 97 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=0.795 $Y2=3.33
r197 97 99 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r198 95 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r199 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r200 92 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=3.33
+ $X2=0.795 $Y2=3.33
r201 92 94 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=3.33
+ $X2=0.24 $Y2=3.33
r202 90 145 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r203 90 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r204 90 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r205 88 116 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=6.96 $Y2=3.33
r206 88 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=7.21 $Y2=3.33
r207 86 102 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.64 $Y2=3.33
r208 86 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.87 $Y2=3.33
r209 84 99 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r210 84 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.01 $Y2=3.33
r211 83 102 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.64 $Y2=3.33
r212 83 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.01 $Y2=3.33
r213 79 82 37.2623 $w=2.98e-07 $l=9.7e-07 $layer=LI1_cond $X=9.805 $Y=1.98
+ $X2=9.805 $Y2=2.95
r214 77 153 3.07827 $w=3e-07 $l=1.11781e-07 $layer=LI1_cond $X=9.805 $Y=3.245
+ $X2=9.867 $Y2=3.33
r215 77 82 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=9.805 $Y=3.245
+ $X2=9.805 $Y2=2.95
r216 73 76 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=8.93 $Y=2.2
+ $X2=8.93 $Y2=2.97
r217 71 150 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.93 $Y=3.245
+ $X2=8.93 $Y2=3.33
r218 71 76 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.93 $Y=3.245
+ $X2=8.93 $Y2=2.97
r219 67 70 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=8.07 $Y=2.2
+ $X2=8.07 $Y2=2.97
r220 65 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.07 $Y=3.245
+ $X2=8.07 $Y2=3.33
r221 65 70 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.07 $Y=3.245
+ $X2=8.07 $Y2=2.97
r222 64 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=3.33
+ $X2=7.21 $Y2=3.33
r223 63 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=8.07 $Y2=3.33
r224 63 64 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=7.375 $Y2=3.33
r225 59 62 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=7.21 $Y=2.2
+ $X2=7.21 $Y2=2.97
r226 57 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.21 $Y=3.245
+ $X2=7.21 $Y2=3.33
r227 57 62 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.21 $Y=3.245
+ $X2=7.21 $Y2=2.97
r228 53 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=3.245
+ $X2=4.59 $Y2=3.33
r229 53 55 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=4.59 $Y=3.245
+ $X2=4.59 $Y2=2.375
r230 49 52 34.5733 $w=2.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.71 $Y=2.28
+ $X2=3.71 $Y2=2.97
r231 47 132 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=3.33
r232 47 52 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=2.97
r233 46 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=2.87 $Y2=3.33
r234 45 132 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.71 $Y2=3.33
r235 45 46 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.035 $Y2=3.33
r236 41 44 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.87 $Y=2.2
+ $X2=2.87 $Y2=2.97
r237 39 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=3.245
+ $X2=2.87 $Y2=3.33
r238 39 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.87 $Y=3.245
+ $X2=2.87 $Y2=2.97
r239 35 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=3.245
+ $X2=2.01 $Y2=3.33
r240 35 37 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.01 $Y=3.245 $X2=2.01
+ $Y2=2.845
r241 31 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=3.245
+ $X2=0.795 $Y2=3.33
r242 31 33 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.795 $Y=3.245
+ $X2=0.795 $Y2=2.845
r243 10 82 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.835 $X2=9.79 $Y2=2.95
r244 10 79 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.835 $X2=9.79 $Y2=1.98
r245 9 76 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=8.79
+ $Y=1.835 $X2=8.93 $Y2=2.97
r246 9 73 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=8.79
+ $Y=1.835 $X2=8.93 $Y2=2.2
r247 8 70 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=7.93
+ $Y=1.835 $X2=8.07 $Y2=2.97
r248 8 67 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=7.93
+ $Y=1.835 $X2=8.07 $Y2=2.2
r249 7 62 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=7.07
+ $Y=1.835 $X2=7.21 $Y2=2.97
r250 7 59 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=7.07
+ $Y=1.835 $X2=7.21 $Y2=2.2
r251 6 142 400 $w=1.7e-07 $l=1.57119e-06 $layer=licon1_PDIFF $count=1 $X=5.31
+ $Y=1.835 $X2=6.35 $Y2=2.97
r252 6 140 150 $w=1.7e-07 $l=8.18474e-07 $layer=licon1_PDIFF $count=4 $X=5.31
+ $Y=1.835 $X2=5.885 $Y2=2.415
r253 6 138 400 $w=1.7e-07 $l=1.24692e-06 $layer=licon1_PDIFF $count=1 $X=5.31
+ $Y=1.835 $X2=6.35 $Y2=2.29
r254 5 55 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=4.45
+ $Y=1.835 $X2=4.59 $Y2=2.375
r255 4 52 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.59
+ $Y=1.835 $X2=3.73 $Y2=2.97
r256 4 49 400 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=1 $X=3.59
+ $Y=1.835 $X2=3.73 $Y2=2.28
r257 3 44 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=1.835 $X2=2.87 $Y2=2.97
r258 3 41 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=1.835 $X2=2.87 $Y2=2.2
r259 2 37 600 $w=1.7e-07 $l=1.07068e-06 $layer=licon1_PDIFF $count=1 $X=1.885
+ $Y=1.835 $X2=2.01 $Y2=2.845
r260 1 33 600 $w=1.7e-07 $l=1.07773e-06 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=1.835 $X2=0.795 $Y2=2.845
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%Y 1 2 3 4 5 6 7 8 9 10 31 39 43 44 47 52
+ 53 54 57 61 65 66 69 73 77 81 85 91 92 93 94 95 96 97 105 109 116
c133 66 0 1.72165e-19 $X=6.875 $Y=1.815
r134 97 109 4.52993 $w=3.85e-07 $l=1.2753e-07 $layer=LI1_cond $X=6 $Y=1.922
+ $X2=5.893 $Y2=1.967
r135 96 109 11.1652 $w=3.83e-07 $l=3.73e-07 $layer=LI1_cond $X=5.52 $Y=1.967
+ $X2=5.893 $Y2=1.967
r136 95 105 2.91516 $w=3.65e-07 $l=1.04523e-07 $layer=LI1_cond $X=5.02 $Y=1.967
+ $X2=4.925 $Y2=1.947
r137 95 110 2.91516 $w=3.65e-07 $l=9.5e-08 $layer=LI1_cond $X=5.02 $Y=1.967
+ $X2=5.115 $Y2=1.967
r138 95 96 11.9734 $w=3.83e-07 $l=4e-07 $layer=LI1_cond $X=5.12 $Y=1.967
+ $X2=5.52 $Y2=1.967
r139 95 110 0.149668 $w=3.83e-07 $l=5e-09 $layer=LI1_cond $X=5.12 $Y=1.967
+ $X2=5.115 $Y2=1.967
r140 94 105 12.1925 $w=3.43e-07 $l=3.65e-07 $layer=LI1_cond $X=4.56 $Y=1.947
+ $X2=4.925 $Y2=1.947
r141 94 106 10.1883 $w=3.43e-07 $l=3.05e-07 $layer=LI1_cond $X=4.56 $Y=1.947
+ $X2=4.255 $Y2=1.947
r142 93 106 5.2077 $w=2.57e-07 $l=1.3e-07 $layer=LI1_cond $X=4.125 $Y=1.947
+ $X2=4.255 $Y2=1.947
r143 93 116 10.4982 $w=4.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.125 $Y=2.12
+ $X2=4.125 $Y2=2.445
r144 85 87 49.7646 $w=2.18e-07 $l=9.5e-07 $layer=LI1_cond $X=9.375 $Y=1.96
+ $X2=9.375 $Y2=2.91
r145 83 85 0.785757 $w=2.18e-07 $l=1.5e-08 $layer=LI1_cond $X=9.375 $Y=1.945
+ $X2=9.375 $Y2=1.96
r146 82 92 3.9502 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=8.595 $Y=1.815
+ $X2=8.5 $Y2=1.815
r147 81 83 6.87824 $w=2.6e-07 $l=1.76635e-07 $layer=LI1_cond $X=9.265 $Y=1.815
+ $X2=9.375 $Y2=1.945
r148 81 82 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=9.265 $Y=1.815
+ $X2=8.595 $Y2=1.815
r149 77 79 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=8.5 $Y=1.96 $X2=8.5
+ $Y2=2.91
r150 75 92 2.49283 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=8.5 $Y=1.945 $X2=8.5
+ $Y2=1.815
r151 75 77 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=8.5 $Y=1.945
+ $X2=8.5 $Y2=1.96
r152 74 91 3.9502 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=7.735 $Y=1.815
+ $X2=7.64 $Y2=1.815
r153 73 92 3.9502 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=8.405 $Y=1.815
+ $X2=8.5 $Y2=1.815
r154 73 74 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=8.405 $Y=1.815
+ $X2=7.735 $Y2=1.815
r155 69 71 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=7.64 $Y=1.96
+ $X2=7.64 $Y2=2.91
r156 67 91 2.49283 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=7.64 $Y=1.945
+ $X2=7.64 $Y2=1.815
r157 67 69 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=7.64 $Y=1.945
+ $X2=7.64 $Y2=1.96
r158 65 91 3.9502 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=7.545 $Y=1.815
+ $X2=7.64 $Y2=1.815
r159 65 66 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=7.545 $Y=1.815
+ $X2=6.875 $Y2=1.815
r160 61 63 47.6009 $w=2.28e-07 $l=9.5e-07 $layer=LI1_cond $X=6.76 $Y=1.96
+ $X2=6.76 $Y2=2.91
r161 59 66 5.23507 $w=2.68e-07 $l=1.59781e-07 $layer=LI1_cond $X=6.76 $Y=1.922
+ $X2=6.875 $Y2=1.815
r162 59 97 34.597 $w=2.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.76 $Y=1.922 $X2=6
+ $Y2=1.922
r163 59 61 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.76 $Y=1.945
+ $X2=6.76 $Y2=1.96
r164 55 95 3.76996 $w=1.9e-07 $l=1.93e-07 $layer=LI1_cond $X=5.02 $Y=2.16
+ $X2=5.02 $Y2=1.967
r165 55 57 16.6364 $w=1.88e-07 $l=2.85e-07 $layer=LI1_cond $X=5.02 $Y=2.16
+ $X2=5.02 $Y2=2.445
r166 54 90 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=1.86
+ $X2=3.605 $Y2=1.86
r167 53 93 5.2077 $w=2.57e-07 $l=1.67958e-07 $layer=LI1_cond $X=3.995 $Y=1.86
+ $X2=4.125 $Y2=1.947
r168 53 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.995 $Y=1.86
+ $X2=3.69 $Y2=1.86
r169 52 90 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=1.775
+ $X2=3.605 $Y2=1.86
r170 51 52 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.605 $Y=1.215
+ $X2=3.605 $Y2=1.775
r171 47 49 49.7646 $w=2.18e-07 $l=9.5e-07 $layer=LI1_cond $X=3.315 $Y=1.96
+ $X2=3.315 $Y2=2.91
r172 45 90 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.315 $Y=1.86
+ $X2=3.605 $Y2=1.86
r173 45 47 0.785757 $w=2.18e-07 $l=1.5e-08 $layer=LI1_cond $X=3.315 $Y=1.945
+ $X2=3.315 $Y2=1.96
r174 43 45 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.205 $Y=1.86
+ $X2=3.315 $Y2=1.86
r175 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.205 $Y=1.86
+ $X2=2.535 $Y2=1.86
r176 39 41 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=2.44 $Y=1.96
+ $X2=2.44 $Y2=2.91
r177 37 44 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.44 $Y=1.945
+ $X2=2.535 $Y2=1.86
r178 37 39 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=2.44 $Y=1.945
+ $X2=2.44 $Y2=1.96
r179 33 36 45.2112 $w=2.58e-07 $l=1.02e-06 $layer=LI1_cond $X=2.31 $Y=1.085
+ $X2=3.33 $Y2=1.085
r180 31 51 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.52 $Y=1.085
+ $X2=3.605 $Y2=1.215
r181 31 36 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=3.52 $Y=1.085
+ $X2=3.33 $Y2=1.085
r182 10 87 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.22
+ $Y=1.835 $X2=9.36 $Y2=2.91
r183 10 85 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=9.22
+ $Y=1.835 $X2=9.36 $Y2=1.96
r184 9 79 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.36
+ $Y=1.835 $X2=8.5 $Y2=2.91
r185 9 77 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=8.36
+ $Y=1.835 $X2=8.5 $Y2=1.96
r186 8 71 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.5
+ $Y=1.835 $X2=7.64 $Y2=2.91
r187 8 69 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.5
+ $Y=1.835 $X2=7.64 $Y2=1.96
r188 7 63 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.64
+ $Y=1.835 $X2=6.78 $Y2=2.91
r189 7 61 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=6.64
+ $Y=1.835 $X2=6.78 $Y2=1.96
r190 6 95 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.835 $X2=5.02 $Y2=1.96
r191 6 57 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=4.88
+ $Y=1.835 $X2=5.02 $Y2=2.445
r192 5 93 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.835 $X2=4.16 $Y2=1.96
r193 5 116 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=4.02
+ $Y=1.835 $X2=4.16 $Y2=2.445
r194 4 49 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=1.835 $X2=3.3 $Y2=2.91
r195 4 47 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=1.835 $X2=3.3 $Y2=1.96
r196 3 41 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=1.835 $X2=2.44 $Y2=2.91
r197 3 39 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=1.835 $X2=2.44 $Y2=1.96
r198 2 36 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.335 $X2=3.33 $Y2=1.05
r199 1 33 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=2.17
+ $Y=0.335 $X2=2.31 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%VGND 1 2 3 12 16 20 22 24 29 34 41 42 45
+ 48 51
r101 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r102 48 49 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r103 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r104 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r105 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r106 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.555 $Y=0 $X2=9.39
+ $Y2=0
r107 39 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.555 $Y=0
+ $X2=9.84 $Y2=0
r108 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r109 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r110 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r111 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=0 $X2=8.53
+ $Y2=0
r112 35 37 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.695 $Y=0
+ $X2=8.88 $Y2=0
r113 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.225 $Y=0 $X2=9.39
+ $Y2=0
r114 34 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.225 $Y=0 $X2=8.88
+ $Y2=0
r115 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r116 32 33 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r117 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.795
+ $Y2=0
r118 30 32 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r119 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.365 $Y=0 $X2=8.53
+ $Y2=0
r120 29 32 467.449 $w=1.68e-07 $l=7.165e-06 $layer=LI1_cond $X=8.365 $Y=0
+ $X2=1.2 $Y2=0
r121 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r122 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.795
+ $Y2=0
r124 24 26 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r125 22 49 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=8.4
+ $Y2=0
r126 22 33 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=1.2
+ $Y2=0
r127 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=0.085
+ $X2=9.39 $Y2=0
r128 18 20 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=9.39 $Y=0.085
+ $X2=9.39 $Y2=0.525
r129 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.53 $Y=0.085
+ $X2=8.53 $Y2=0
r130 14 16 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=8.53 $Y=0.085
+ $X2=8.53 $Y2=0.525
r131 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r132 10 12 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.47
r133 3 20 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=9.25
+ $Y=0.235 $X2=9.39 $Y2=0.525
r134 2 16 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=8.39
+ $Y=0.235 $X2=8.53 $Y2=0.525
r135 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.655
+ $Y=0.345 $X2=0.795 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%A_324_45# 1 2 3 4 5 16 26 28 32 34
c57 34 0 5.86634e-20 $X=4.78 $Y=0.35
r58 30 32 8.08732 $w=2.83e-07 $l=2e-07 $layer=LI1_cond $X=5.617 $Y=0.425
+ $X2=5.617 $Y2=0.625
r59 29 34 8.26956 $w=1.8e-07 $l=1.69926e-07 $layer=LI1_cond $X=4.945 $Y=0.34
+ $X2=4.78 $Y2=0.35
r60 28 30 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=5.475 $Y=0.34
+ $X2=5.617 $Y2=0.425
r61 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.475 $Y=0.34
+ $X2=4.945 $Y2=0.34
r62 24 34 0.718145 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.78 $Y=0.445
+ $X2=4.78 $Y2=0.35
r63 24 26 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.78 $Y=0.445
+ $X2=4.78 $Y2=0.46
r64 21 23 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=2.82 $Y=0.35
+ $X2=3.84 $Y2=0.35
r65 18 21 61.5837 $w=1.88e-07 $l=1.055e-06 $layer=LI1_cond $X=1.765 $Y=0.35
+ $X2=2.82 $Y2=0.35
r66 16 34 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.615 $Y=0.35
+ $X2=4.78 $Y2=0.35
r67 16 23 45.2392 $w=1.88e-07 $l=7.75e-07 $layer=LI1_cond $X=4.615 $Y=0.35
+ $X2=3.84 $Y2=0.35
r68 5 32 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=5.5
+ $Y=0.335 $X2=5.64 $Y2=0.625
r69 4 26 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.64
+ $Y=0.335 $X2=4.78 $Y2=0.46
r70 3 23 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=3.62
+ $Y=0.335 $X2=3.84 $Y2=0.35
r71 2 21 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=2.6
+ $Y=0.335 $X2=2.82 $Y2=0.35
r72 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.62
+ $Y=0.225 $X2=1.765 $Y2=0.35
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%A_842_67# 1 2 3 4 15 18 19 20 24 30 31 32
c62 24 0 1.51661e-19 $X=4.35 $Y=1.05
r63 32 35 2.65948 $w=2.58e-07 $l=6e-08 $layer=LI1_cond $X=7.645 $Y=0.415
+ $X2=7.645 $Y2=0.475
r64 29 31 3.64489 $w=3.83e-07 $l=9.5e-08 $layer=LI1_cond $X=5.21 $Y=1.052
+ $X2=5.305 $Y2=1.052
r65 29 30 5.80212 $w=3.83e-07 $l=9.5e-08 $layer=LI1_cond $X=5.21 $Y=1.052
+ $X2=5.115 $Y2=1.052
r66 24 26 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=4.345 $Y=1.05
+ $X2=4.345 $Y2=1.15
r67 20 22 37.4978 $w=2.08e-07 $l=7.1e-07 $layer=LI1_cond $X=6.1 $Y=0.415
+ $X2=6.81 $Y2=0.415
r68 19 32 1.99039 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=7.515 $Y=0.415
+ $X2=7.645 $Y2=0.415
r69 19 22 37.2338 $w=2.08e-07 $l=7.05e-07 $layer=LI1_cond $X=7.515 $Y=0.415
+ $X2=6.81 $Y2=0.415
r70 17 20 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.015 $Y=0.52
+ $X2=6.1 $Y2=0.415
r71 17 18 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.015 $Y=0.52
+ $X2=6.015 $Y2=0.96
r72 15 18 7.39867 $w=2.85e-07 $l=1.79538e-07 $layer=LI1_cond $X=5.93 $Y=1.102
+ $X2=6.015 $Y2=0.96
r73 15 31 25.2729 $w=2.83e-07 $l=6.25e-07 $layer=LI1_cond $X=5.93 $Y=1.102
+ $X2=5.305 $Y2=1.102
r74 14 26 1.02732 $w=1.9e-07 $l=1e-07 $layer=LI1_cond $X=4.445 $Y=1.15 $X2=4.345
+ $Y2=1.15
r75 14 30 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=4.445 $Y=1.15
+ $X2=5.115 $Y2=1.15
r76 4 35 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=7.53
+ $Y=0.235 $X2=7.67 $Y2=0.475
r77 3 22 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.67 $Y=0.235
+ $X2=6.81 $Y2=0.415
r78 2 29 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=5.07
+ $Y=0.335 $X2=5.21 $Y2=1.025
r79 1 24 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=4.21
+ $Y=0.335 $X2=4.35 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_4%A_1251_47# 1 2 3 4 5 16 20 24 26 30 32 36
+ 40 41 42
r46 39 40 6.36683 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.24 $Y=0.865
+ $X2=7.345 $Y2=0.865
r47 34 36 24.4 $w=1.98e-07 $l=4.4e-07 $layer=LI1_cond $X=9.825 $Y=0.86 $X2=9.825
+ $Y2=0.42
r48 33 42 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.045 $Y=0.945
+ $X2=8.955 $Y2=0.945
r49 32 34 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=9.725 $Y=0.945
+ $X2=9.825 $Y2=0.86
r50 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.725 $Y=0.945
+ $X2=9.045 $Y2=0.945
r51 28 42 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=0.86
+ $X2=8.955 $Y2=0.945
r52 28 30 27.1111 $w=1.78e-07 $l=4.4e-07 $layer=LI1_cond $X=8.955 $Y=0.86
+ $X2=8.955 $Y2=0.42
r53 27 41 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=8.195 $Y=0.945
+ $X2=8.095 $Y2=0.945
r54 26 42 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.865 $Y=0.945
+ $X2=8.955 $Y2=0.945
r55 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.865 $Y=0.945
+ $X2=8.195 $Y2=0.945
r56 22 41 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.095 $Y=0.86
+ $X2=8.095 $Y2=0.945
r57 22 24 24.4 $w=1.98e-07 $l=4.4e-07 $layer=LI1_cond $X=8.095 $Y=0.86 $X2=8.095
+ $Y2=0.42
r58 20 41 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.995 $Y=0.945
+ $X2=8.095 $Y2=0.945
r59 20 40 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.995 $Y=0.945
+ $X2=7.345 $Y2=0.945
r60 16 39 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=7.18 $Y=0.865 $X2=7.24
+ $Y2=0.865
r61 16 18 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=7.18 $Y=0.865 $X2=6.38
+ $Y2=0.865
r62 5 36 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.68
+ $Y=0.235 $X2=9.82 $Y2=0.42
r63 4 30 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.82
+ $Y=0.235 $X2=8.96 $Y2=0.42
r64 3 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.96
+ $Y=0.235 $X2=8.1 $Y2=0.42
r65 2 39 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=7.1
+ $Y=0.235 $X2=7.24 $Y2=0.865
r66 1 18 182 $w=1.7e-07 $l=6.89674e-07 $layer=licon1_NDIFF $count=1 $X=6.255
+ $Y=0.235 $X2=6.38 $Y2=0.865
.ends

