* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxbp_lp D GATE VGND VNB VPB VPWR Q Q_N
M1000 a_1597_361# a_969_407# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.6753e+12p ps=1.397e+07u
M1001 VGND a_969_407# a_900_47# VNB nshort w=420000u l=150000u
+  ad=1.0794e+12p pd=1.015e+07u as=1.638e+11p ps=1.62e+06u
M1002 VGND a_969_407# a_1403_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1003 a_1662_131# a_969_407# a_1597_361# VPB phighvt w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=0p ps=0u
M1004 a_1863_367# a_1662_131# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1005 VPWR a_969_407# a_927_519# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 Q_N a_1662_131# a_1863_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.402e+11p pd=3.06e+06u as=0p ps=0u
M1007 a_556_47# a_350_111# a_469_47# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1008 VGND a_350_111# a_556_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_720_47# a_27_111# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1010 VGND D a_114_111# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1011 a_272_111# GATE VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1012 a_567_475# a_350_111# a_469_47# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.76e+11p ps=1.83e+06u
M1013 a_741_475# a_27_111# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1014 a_969_407# a_798_47# a_1152_361# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.465e+11p pd=3.07e+06u as=2.646e+11p ps=2.94e+06u
M1015 VPWR a_350_111# a_567_475# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_969_407# a_1418_361# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1017 a_798_47# a_350_111# a_741_475# VPB phighvt w=640000u l=150000u
+  ad=2.254e+11p pd=2.06e+06u as=0p ps=0u
M1018 a_1418_361# a_969_407# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.465e+11p ps=3.07e+06u
M1019 a_798_47# a_469_47# a_720_47# VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1020 a_900_47# a_350_111# a_798_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_114_111# D a_27_111# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1022 a_969_407# a_798_47# a_1133_47# VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=1.764e+11p ps=2.1e+06u
M1023 a_350_111# GATE a_278_481# VPB phighvt w=640000u l=150000u
+  ad=4.904e+11p pd=3.78e+06u as=1.344e+11p ps=1.7e+06u
M1024 a_1662_131# a_969_407# a_1584_131# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1025 a_278_481# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1152_361# a_798_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1860_53# a_1662_131# VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1028 VPWR D a_112_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1029 a_927_519# a_469_47# a_798_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Q_N a_1662_131# a_1860_53# VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1031 a_1133_47# a_798_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_112_481# D a_27_111# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1033 a_350_111# GATE a_272_111# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1034 a_1403_47# a_969_407# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1035 a_1584_131# a_969_407# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
