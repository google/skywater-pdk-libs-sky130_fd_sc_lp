# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a21bo_m
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a21bo_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 0.765000 2.445000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.975000 0.840000 3.205000 1.750000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 1.025000 1.285000 2.120000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 0.470000 0.365000 0.800000 ;
        RECT 0.155000 0.800000 0.325000 2.685000 ;
        RECT 0.155000 2.685000 0.365000 3.015000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.505000  1.475000 0.675000 2.335000 ;
      RECT 0.505000  2.335000 1.910000 2.505000 ;
      RECT 0.585000  0.085000 0.795000 0.800000 ;
      RECT 0.585000  2.755000 0.795000 3.245000 ;
      RECT 1.015000  0.515000 1.225000 0.675000 ;
      RECT 1.015000  0.675000 1.875000 0.845000 ;
      RECT 1.015000  2.695000 1.735000 3.025000 ;
      RECT 1.530000  0.085000 1.860000 0.485000 ;
      RECT 1.700000  1.625000 2.795000 1.795000 ;
      RECT 1.700000  1.795000 1.910000 2.335000 ;
      RECT 1.705000  0.845000 1.875000 1.435000 ;
      RECT 2.040000  0.285000 2.795000 0.495000 ;
      RECT 2.130000  1.975000 3.200000 2.145000 ;
      RECT 2.130000  2.145000 2.340000 2.505000 ;
      RECT 2.560000  2.325000 2.770000 3.245000 ;
      RECT 2.625000  0.495000 2.795000 1.625000 ;
      RECT 2.975000  0.085000 3.165000 0.545000 ;
      RECT 2.990000  2.145000 3.200000 2.505000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__a21bo_m
