* File: sky130_fd_sc_lp__o32ai_m.pex.spice
* Created: Fri Aug 28 11:18:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32AI_M%B1 2 3 4 5 6 7 9 12 16 17 18 19 20 21 28
r41 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.105 $X2=0.27 $Y2=1.105
r42 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r43 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r44 18 19 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r45 18 29 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.105
r46 17 29 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.105
r47 15 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.445
+ $X2=0.27 $Y2=1.105
r48 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.445
+ $X2=0.27 $Y2=1.61
r49 14 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.09
+ $X2=0.27 $Y2=1.105
r50 10 12 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.82 $Y=2.39
+ $X2=0.82 $Y2=2.885
r51 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.75 $Y=0.94 $X2=0.75
+ $Y2=0.62
r52 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.745 $Y=2.315
+ $X2=0.82 $Y2=2.39
r53 5 6 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.745 $Y=2.315
+ $X2=0.435 $Y2=2.315
r54 4 14 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=1.015
+ $X2=0.27 $Y2=1.09
r55 3 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.675 $Y=1.015
+ $X2=0.75 $Y2=0.94
r56 3 4 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.675 $Y=1.015
+ $X2=0.435 $Y2=1.015
r57 2 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.36 $Y=2.24
+ $X2=0.435 $Y2=2.315
r58 2 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.36 $Y=2.24 $X2=0.36
+ $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_M%B2 3 7 11 12 13 14 15 16 22
c40 3 0 1.00733e-19 $X=1.18 $Y=0.62
r41 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.09
+ $Y=1.495 $X2=1.09 $Y2=1.495
r42 15 16 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.145 $Y=2.035
+ $X2=1.145 $Y2=2.405
r43 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.145 $Y=1.665
+ $X2=1.145 $Y2=2.035
r44 14 23 6.99698 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=1.145 $Y=1.665
+ $X2=1.145 $Y2=1.495
r45 13 23 8.23174 $w=2.78e-07 $l=2e-07 $layer=LI1_cond $X=1.145 $Y=1.295
+ $X2=1.145 $Y2=1.495
r46 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.09 $Y=1.835
+ $X2=1.09 $Y2=1.495
r47 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.835
+ $X2=1.09 $Y2=2
r48 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.33
+ $X2=1.09 $Y2=1.495
r49 7 12 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=1.18 $Y=2.885
+ $X2=1.18 $Y2=2
r50 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.18 $Y=0.62 $X2=1.18
+ $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_M%A3 3 7 11 12 13 14 15 16 22
r40 15 16 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.655 $Y=2.035
+ $X2=1.655 $Y2=2.405
r41 14 15 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.655 $Y=1.665
+ $X2=1.655 $Y2=2.035
r42 13 14 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.655 $Y=1.295
+ $X2=1.655 $Y2=1.665
r43 13 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.375 $X2=1.63 $Y2=1.375
r44 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.63 $Y=1.715
+ $X2=1.63 $Y2=1.375
r45 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.715
+ $X2=1.63 $Y2=1.88
r46 10 22 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.21
+ $X2=1.63 $Y2=1.375
r47 7 12 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.61 $Y=2.885
+ $X2=1.61 $Y2=1.88
r48 3 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.61 $Y=0.62 $X2=1.61
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_M%A2 3 7 11 12 13 14 15 16 22
r42 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.17
+ $Y=1.495 $X2=2.17 $Y2=1.495
r43 15 16 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.165 $Y=2.035
+ $X2=2.165 $Y2=2.405
r44 14 15 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.165 $Y=1.665
+ $X2=2.165 $Y2=2.035
r45 14 23 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=2.165 $Y=1.665
+ $X2=2.165 $Y2=1.495
r46 13 23 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=2.165 $Y=1.295
+ $X2=2.165 $Y2=1.495
r47 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.17 $Y=1.835
+ $X2=2.17 $Y2=1.495
r48 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.835
+ $X2=2.17 $Y2=2
r49 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.33
+ $X2=2.17 $Y2=1.495
r50 7 12 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=2.08 $Y=2.885
+ $X2=2.08 $Y2=2
r51 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.08 $Y=0.62 $X2=2.08
+ $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_M%A1 3 5 7 8 9 10 11 13 16 17 18 19 20 21 28
r40 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.975
+ $Y=1.105 $X2=2.975 $Y2=1.105
r41 20 21 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.047 $Y=2.035
+ $X2=3.047 $Y2=2.405
r42 19 20 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.047 $Y=1.665
+ $X2=3.047 $Y2=2.035
r43 18 19 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.047 $Y=1.295
+ $X2=3.047 $Y2=1.665
r44 18 29 6.95124 $w=3.13e-07 $l=1.9e-07 $layer=LI1_cond $X=3.047 $Y=1.295
+ $X2=3.047 $Y2=1.105
r45 17 29 6.58539 $w=3.13e-07 $l=1.8e-07 $layer=LI1_cond $X=3.047 $Y=0.925
+ $X2=3.047 $Y2=1.105
r46 15 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.975 $Y=1.445
+ $X2=2.975 $Y2=1.105
r47 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.445
+ $X2=2.975 $Y2=1.61
r48 14 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.975 $Y=1.09
+ $X2=2.975 $Y2=1.105
r49 13 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.885 $Y=2.24
+ $X2=2.885 $Y2=1.61
r50 10 14 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.81 $Y=1.015
+ $X2=2.975 $Y2=1.09
r51 10 11 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.81 $Y=1.015
+ $X2=2.585 $Y2=1.015
r52 8 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.81 $Y=2.315
+ $X2=2.885 $Y2=2.24
r53 8 9 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.81 $Y=2.315
+ $X2=2.515 $Y2=2.315
r54 5 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.51 $Y=0.94
+ $X2=2.585 $Y2=1.015
r55 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.51 $Y=0.94 $X2=2.51
+ $Y2=0.62
r56 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.44 $Y=2.39
+ $X2=2.515 $Y2=2.315
r57 1 3 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.44 $Y=2.39 $X2=2.44
+ $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_M%VPWR 1 2 7 9 11 13 15 17 30
r37 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r39 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 23 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 20 23 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 18 26 3.49867 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r45 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 17 29 3.49902 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=3.132 $Y2=3.33
r47 17 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 15 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 11 29 3.34488 $w=1.9e-07 $l=1.69245e-07 $layer=LI1_cond $X=3 $Y=3.245
+ $X2=3.132 $Y2=3.33
r51 11 13 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.95
r52 7 26 3.34522 $w=1.9e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.227 $Y2=3.33
r53 7 9 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.36 $Y2=2.95
r54 2 13 600 $w=1.7e-07 $l=5.96867e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=2.675 $X2=2.99 $Y2=2.95
r55 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=2.675 $X2=0.37 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_M%Y 1 2 7 8 12 13 14 15 16
r46 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.835
+ $X2=2.64 $Y2=2.835
r47 14 15 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.835
+ $X2=2.16 $Y2=2.835
r48 14 26 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.68 $Y=2.835
+ $X2=1.395 $Y2=2.835
r49 13 26 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.2 $Y=2.835
+ $X2=1.395 $Y2=2.835
r50 13 22 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.2 $Y=2.835
+ $X2=0.825 $Y2=2.835
r51 12 22 2.73254 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=0.73 $Y=2.835
+ $X2=0.825 $Y2=2.835
r52 8 12 5.03363 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=0.74 $Y=2.67
+ $X2=0.73 $Y2=2.835
r53 7 11 8.52485 $w=3.22e-07 $l=3.07409e-07 $layer=LI1_cond $X=0.74 $Y=1.01
+ $X2=0.965 $Y2=0.815
r54 7 8 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=0.74 $Y=1.01 $X2=0.74
+ $Y2=2.67
r55 2 26 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=1.255
+ $Y=2.675 $X2=1.395 $Y2=2.835
r56 1 11 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=0.825
+ $Y=0.41 $X2=0.965 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_M%A_66_82# 1 2 3 10 16 17 20 22
r33 22 25 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.455 $Y=0.355
+ $X2=0.455 $Y2=0.555
r34 18 20 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=2.285 $Y=0.82
+ $X2=2.285 $Y2=0.685
r35 16 18 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.19 $Y=0.905
+ $X2=2.285 $Y2=0.82
r36 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.19 $Y=0.905 $X2=1.5
+ $Y2=0.905
r37 13 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.405 $Y=0.82
+ $X2=1.5 $Y2=0.905
r38 13 15 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=1.405 $Y=0.82
+ $X2=1.405 $Y2=0.555
r39 12 15 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=1.405 $Y=0.44
+ $X2=1.405 $Y2=0.555
r40 11 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=0.355
+ $X2=0.455 $Y2=0.355
r41 10 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.31 $Y=0.355
+ $X2=1.405 $Y2=0.44
r42 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.31 $Y=0.355
+ $X2=0.62 $Y2=0.355
r43 3 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.41 $X2=2.295 $Y2=0.685
r44 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.255
+ $Y=0.41 $X2=1.395 $Y2=0.555
r45 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.33
+ $Y=0.41 $X2=0.455 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_M%VGND 1 2 9 11 15 17 19 26 27 30 33
c34 9 0 1.00733e-19 $X=1.845 $Y=0.555
r35 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r36 27 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r37 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r38 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.725
+ $Y2=0
r39 24 26 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.12
+ $Y2=0
r40 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r41 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.845
+ $Y2=0
r42 19 21 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r43 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r44 17 22 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r45 17 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r46 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0
r47 13 15 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0.555
r48 12 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.845
+ $Y2=0
r49 11 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.725
+ $Y2=0
r50 11 12 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.01
+ $Y2=0
r51 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=0.085
+ $X2=1.845 $Y2=0
r52 7 9 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.845 $Y=0.085
+ $X2=1.845 $Y2=0.555
r53 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.41 $X2=2.725 $Y2=0.555
r54 1 9 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.41 $X2=1.845 $Y2=0.555
.ends

