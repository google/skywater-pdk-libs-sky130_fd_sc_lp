* File: sky130_fd_sc_lp__and3b_4.pxi.spice
* Created: Fri Aug 28 10:06:52 2020
* 
x_PM_SKY130_FD_SC_LP__AND3B_4%A_N N_A_N_M1015_g N_A_N_M1009_g A_N A_N A_N A_N
+ A_N N_A_N_c_86_n N_A_N_c_87_n PM_SKY130_FD_SC_LP__AND3B_4%A_N
x_PM_SKY130_FD_SC_LP__AND3B_4%A_242_23# N_A_242_23#_M1010_d N_A_242_23#_M1001_d
+ N_A_242_23#_M1007_d N_A_242_23#_M1002_g N_A_242_23#_M1000_g
+ N_A_242_23#_M1003_g N_A_242_23#_M1006_g N_A_242_23#_M1008_g
+ N_A_242_23#_M1013_g N_A_242_23#_M1012_g N_A_242_23#_M1014_g
+ N_A_242_23#_c_204_p N_A_242_23#_c_117_n N_A_242_23#_c_118_n
+ N_A_242_23#_c_212_p N_A_242_23#_c_173_p N_A_242_23#_c_141_p
+ N_A_242_23#_c_119_n N_A_242_23#_c_120_n N_A_242_23#_c_130_n
+ N_A_242_23#_c_121_n N_A_242_23#_c_122_n N_A_242_23#_c_131_n
+ N_A_242_23#_c_123_n N_A_242_23#_c_124_n PM_SKY130_FD_SC_LP__AND3B_4%A_242_23#
x_PM_SKY130_FD_SC_LP__AND3B_4%C N_C_M1001_g N_C_M1011_g C N_C_c_250_n
+ N_C_c_251_n PM_SKY130_FD_SC_LP__AND3B_4%C
x_PM_SKY130_FD_SC_LP__AND3B_4%B N_B_M1004_g N_B_M1005_g B N_B_c_290_n
+ N_B_c_291_n PM_SKY130_FD_SC_LP__AND3B_4%B
x_PM_SKY130_FD_SC_LP__AND3B_4%A_49_133# N_A_49_133#_M1015_s N_A_49_133#_M1009_s
+ N_A_49_133#_M1010_g N_A_49_133#_c_322_n N_A_49_133#_M1007_g
+ N_A_49_133#_c_323_n N_A_49_133#_c_329_n N_A_49_133#_c_330_n
+ N_A_49_133#_c_346_n N_A_49_133#_c_324_n N_A_49_133#_c_375_p
+ N_A_49_133#_c_325_n PM_SKY130_FD_SC_LP__AND3B_4%A_49_133#
x_PM_SKY130_FD_SC_LP__AND3B_4%VPWR N_VPWR_M1009_d N_VPWR_M1006_s N_VPWR_M1014_s
+ N_VPWR_M1005_d N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n N_VPWR_c_401_n
+ N_VPWR_c_402_n N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n
+ N_VPWR_c_407_n VPWR N_VPWR_c_408_n N_VPWR_c_397_n N_VPWR_c_410_n
+ N_VPWR_c_411_n PM_SKY130_FD_SC_LP__AND3B_4%VPWR
x_PM_SKY130_FD_SC_LP__AND3B_4%X N_X_M1002_d N_X_M1008_d N_X_M1000_d N_X_M1013_d
+ N_X_c_467_n N_X_c_468_n N_X_c_469_n N_X_c_513_p N_X_c_470_n N_X_c_514_p
+ N_X_c_471_n X X X X N_X_c_473_n PM_SKY130_FD_SC_LP__AND3B_4%X
x_PM_SKY130_FD_SC_LP__AND3B_4%VGND N_VGND_M1015_d N_VGND_M1003_s N_VGND_M1012_s
+ N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n
+ N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n N_VGND_c_527_n VGND
+ N_VGND_c_528_n N_VGND_c_529_n PM_SKY130_FD_SC_LP__AND3B_4%VGND
cc_1 VNB N_A_N_M1009_g 0.00750648f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.045
cc_2 VNB A_N 0.00710732f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_3 VNB N_A_N_c_86_n 0.0424024f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_4 VNB N_A_N_c_87_n 0.0218059f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.195
cc_5 VNB N_A_242_23#_M1002_g 0.0262975f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_6 VNB N_A_242_23#_M1003_g 0.022241f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_7 VNB N_A_242_23#_M1008_g 0.0222554f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.295
cc_8 VNB N_A_242_23#_M1012_g 0.0246709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_242_23#_c_117_n 0.00233717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_242_23#_c_118_n 3.45182e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_242_23#_c_119_n 0.057808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_242_23#_c_120_n 0.00636685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_242_23#_c_121_n 0.0010166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_242_23#_c_122_n 0.00779277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_242_23#_c_123_n 0.0237994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_242_23#_c_124_n 0.067061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_M1011_g 0.0245715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C_c_250_n 0.0239669f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_19 VNB N_C_c_251_n 0.00319189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_M1004_g 0.0242252f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.875
cc_21 VNB N_B_c_290_n 0.0241877f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_22 VNB N_B_c_291_n 0.00302401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_49_133#_M1010_g 0.0303761f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_24 VNB N_A_49_133#_c_322_n 0.0307783f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_25 VNB N_A_49_133#_c_323_n 0.043909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_49_133#_c_324_n 4.36972e-19 $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.925
cc_27 VNB N_A_49_133#_c_325_n 0.00824297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_397_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_467_n 0.00732741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_468_n 7.4031e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_469_n 0.00130814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_470_n 0.00577414f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.195
cc_33 VNB N_X_c_471_n 0.00185325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_519_n 0.00466354f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_35 VNB N_VGND_c_520_n 5.00391e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_521_n 0.00534544f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_37 VNB N_VGND_c_522_n 0.0311014f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.555
cc_38 VNB N_VGND_c_523_n 0.00423165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_524_n 0.014949f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.925
cc_40 VNB N_VGND_c_525_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_526_n 0.01628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_527_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.665
cc_43 VNB N_VGND_c_528_n 0.0455532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_529_n 0.270875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A_N_M1009_g 0.0231652f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.045
cc_46 VPB A_N 0.00124334f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_47 VPB N_A_242_23#_M1000_g 0.0216446f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_242_23#_M1006_g 0.0183243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_242_23#_M1013_g 0.0183375f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.035
cc_50 VPB N_A_242_23#_M1014_g 0.0186863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_242_23#_c_118_n 0.00141617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_242_23#_c_130_n 0.0515828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_242_23#_c_131_n 0.0154772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_242_23#_c_123_n 0.00798114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_242_23#_c_124_n 0.0120167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_C_M1001_g 0.0193048f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.875
cc_57 VPB N_C_c_250_n 0.00616042f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_58 VPB N_C_c_251_n 0.00237922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_B_M1005_g 0.0196909f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_B_c_290_n 0.00800268f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_61 VPB N_B_c_291_n 0.00560319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_49_133#_c_322_n 0.00695615f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_63 VPB N_A_49_133#_M1007_g 0.0234048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_49_133#_c_323_n 0.0278744f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_49_133#_c_329_n 0.0172364f $X=-0.19 $Y=1.655 $X2=0.707 $Y2=1.195
cc_66 VPB N_A_49_133#_c_330_n 0.0129205f $X=-0.19 $Y=1.655 $X2=0.707 $Y2=1.525
cc_67 VPB N_A_49_133#_c_324_n 0.00148424f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.925
cc_68 VPB N_VPWR_c_398_n 0.019911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_399_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.36
cc_70 VPB N_VPWR_c_400_n 0.0133553f $X=-0.19 $Y=1.655 $X2=0.707 $Y2=1.195
cc_71 VPB N_VPWR_c_401_n 0.00213954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_402_n 0.0158804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_403_n 0.00276847f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_404_n 0.0309422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_405_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_406_n 0.0147084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_407_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_408_n 0.0260163f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_397_n 0.0615123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_410_n 0.00510611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_411_n 0.00510611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_X_c_467_n 0.00291334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_X_c_473_n 0.00777464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 A_N N_A_242_23#_M1002_g 0.00226073f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_85 N_A_N_c_86_n N_A_242_23#_M1002_g 0.0108689f $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_86 N_A_N_c_87_n N_A_242_23#_M1002_g 0.0078602f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_87 A_N N_A_242_23#_M1000_g 0.0011393f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_88 N_A_N_M1009_g N_A_242_23#_c_124_n 0.0163658f $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_89 A_N N_A_49_133#_c_323_n 0.104179f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_90 N_A_N_c_87_n N_A_49_133#_c_323_n 0.0252067f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_91 N_A_N_M1009_g N_A_49_133#_c_329_n 0.0111117f $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_92 A_N N_A_49_133#_c_329_n 0.0106526f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_93 A_N N_VPWR_M1009_d 0.00345784f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_94 N_A_N_M1009_g N_X_c_467_n 0.00217229f $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_95 A_N N_X_c_467_n 0.0641855f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_96 N_A_N_c_86_n N_X_c_467_n 0.0022345f $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_97 A_N N_X_c_469_n 0.0136165f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_98 N_A_N_c_86_n N_X_c_469_n 4.51926e-19 $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_99 N_A_N_c_87_n N_X_c_469_n 4.23027e-19 $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_100 A_N N_VGND_M1015_d 0.00490698f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_101 A_N N_VGND_c_519_n 0.0326166f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_102 N_A_N_c_87_n N_VGND_c_519_n 0.00107846f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_103 A_N N_VGND_c_522_n 0.00533686f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_104 N_A_N_c_87_n N_VGND_c_522_n 0.00275448f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_105 A_N N_VGND_c_529_n 0.00608074f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_106 N_A_N_c_87_n N_VGND_c_529_n 0.00293451f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_107 N_A_242_23#_M1014_g N_C_M1001_g 0.04509f $X=2.575 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_242_23#_c_118_n N_C_M1001_g 0.00388767f $X=2.71 $Y=1.93 $X2=0 $Y2=0
cc_109 N_A_242_23#_c_141_p N_C_M1001_g 0.013472f $X=3.295 $Y=2.095 $X2=0 $Y2=0
cc_110 N_A_242_23#_M1012_g N_C_M1011_g 0.0276701f $X=2.575 $Y=0.665 $X2=0 $Y2=0
cc_111 N_A_242_23#_c_117_n N_C_M1011_g 0.0034595f $X=2.71 $Y=1.425 $X2=0 $Y2=0
cc_112 N_A_242_23#_c_120_n N_C_M1011_g 0.00993576f $X=3.785 $Y=0.71 $X2=0 $Y2=0
cc_113 N_A_242_23#_c_122_n N_C_M1011_g 0.015296f $X=3.33 $Y=0.71 $X2=0 $Y2=0
cc_114 N_A_242_23#_c_117_n N_C_c_250_n 4.83438e-19 $X=2.71 $Y=1.425 $X2=0 $Y2=0
cc_115 N_A_242_23#_c_118_n N_C_c_250_n 4.83438e-19 $X=2.71 $Y=1.93 $X2=0 $Y2=0
cc_116 N_A_242_23#_c_141_p N_C_c_250_n 0.00257775f $X=3.295 $Y=2.095 $X2=0 $Y2=0
cc_117 N_A_242_23#_c_121_n N_C_c_250_n 0.00120117f $X=2.71 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A_242_23#_c_122_n N_C_c_250_n 0.00339108f $X=3.33 $Y=0.71 $X2=0 $Y2=0
cc_119 N_A_242_23#_c_124_n N_C_c_250_n 0.0205364f $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_120 N_A_242_23#_c_117_n N_C_c_251_n 0.00591553f $X=2.71 $Y=1.425 $X2=0 $Y2=0
cc_121 N_A_242_23#_c_118_n N_C_c_251_n 0.0118001f $X=2.71 $Y=1.93 $X2=0 $Y2=0
cc_122 N_A_242_23#_c_141_p N_C_c_251_n 0.0182805f $X=3.295 $Y=2.095 $X2=0 $Y2=0
cc_123 N_A_242_23#_c_121_n N_C_c_251_n 0.0142096f $X=2.71 $Y=1.51 $X2=0 $Y2=0
cc_124 N_A_242_23#_c_122_n N_C_c_251_n 0.0207162f $X=3.33 $Y=0.71 $X2=0 $Y2=0
cc_125 N_A_242_23#_c_124_n N_C_c_251_n 2.99608e-19 $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_126 N_A_242_23#_c_120_n N_B_M1004_g 0.0348067f $X=3.785 $Y=0.71 $X2=0 $Y2=0
cc_127 N_A_242_23#_c_120_n N_B_c_290_n 0.00397376f $X=3.785 $Y=0.71 $X2=0 $Y2=0
cc_128 N_A_242_23#_c_120_n N_B_c_291_n 0.0213194f $X=3.785 $Y=0.71 $X2=0 $Y2=0
cc_129 N_A_242_23#_c_119_n N_A_49_133#_M1010_g 0.0346367f $X=4.52 $Y=0.71 $X2=0
+ $Y2=0
cc_130 N_A_242_23#_c_123_n N_A_49_133#_M1010_g 0.00463554f $X=4.447 $Y=1.815
+ $X2=0 $Y2=0
cc_131 N_A_242_23#_c_119_n N_A_49_133#_c_322_n 0.00165323f $X=4.52 $Y=0.71 $X2=0
+ $Y2=0
cc_132 N_A_242_23#_c_131_n N_A_49_133#_c_322_n 0.00323663f $X=4.3 $Y=1.98 $X2=0
+ $Y2=0
cc_133 N_A_242_23#_c_123_n N_A_49_133#_c_322_n 0.00287983f $X=4.447 $Y=1.815
+ $X2=0 $Y2=0
cc_134 N_A_242_23#_c_131_n N_A_49_133#_M1007_g 0.00336104f $X=4.3 $Y=1.98 $X2=0
+ $Y2=0
cc_135 N_A_242_23#_c_123_n N_A_49_133#_M1007_g 0.002463f $X=4.447 $Y=1.815 $X2=0
+ $Y2=0
cc_136 N_A_242_23#_M1000_g N_A_49_133#_c_329_n 0.0134403f $X=1.285 $Y=2.465
+ $X2=0 $Y2=0
cc_137 N_A_242_23#_M1006_g N_A_49_133#_c_329_n 0.0117636f $X=1.715 $Y=2.465
+ $X2=0 $Y2=0
cc_138 N_A_242_23#_M1013_g N_A_49_133#_c_329_n 0.0105439f $X=2.145 $Y=2.465
+ $X2=0 $Y2=0
cc_139 N_A_242_23#_M1001_d N_A_49_133#_c_346_n 0.00494544f $X=3.155 $Y=1.835
+ $X2=0 $Y2=0
cc_140 N_A_242_23#_M1014_g N_A_49_133#_c_346_n 0.0151726f $X=2.575 $Y=2.465
+ $X2=0 $Y2=0
cc_141 N_A_242_23#_c_173_p N_A_49_133#_c_346_n 0.0090121f $X=2.795 $Y=2.095
+ $X2=0 $Y2=0
cc_142 N_A_242_23#_c_141_p N_A_49_133#_c_346_n 0.0351575f $X=3.295 $Y=2.095
+ $X2=0 $Y2=0
cc_143 N_A_242_23#_c_131_n N_A_49_133#_c_324_n 0.0216464f $X=4.3 $Y=1.98 $X2=0
+ $Y2=0
cc_144 N_A_242_23#_c_123_n N_A_49_133#_c_324_n 0.00551246f $X=4.447 $Y=1.815
+ $X2=0 $Y2=0
cc_145 N_A_242_23#_c_119_n N_A_49_133#_c_325_n 0.0403625f $X=4.52 $Y=0.71 $X2=0
+ $Y2=0
cc_146 N_A_242_23#_c_131_n N_A_49_133#_c_325_n 0.011252f $X=4.3 $Y=1.98 $X2=0
+ $Y2=0
cc_147 N_A_242_23#_c_123_n N_A_49_133#_c_325_n 0.0229477f $X=4.447 $Y=1.815
+ $X2=0 $Y2=0
cc_148 N_A_242_23#_c_118_n N_VPWR_M1014_s 0.00112177f $X=2.71 $Y=1.93 $X2=0
+ $Y2=0
cc_149 N_A_242_23#_c_173_p N_VPWR_M1014_s 9.65132e-19 $X=2.795 $Y=2.095 $X2=0
+ $Y2=0
cc_150 N_A_242_23#_c_141_p N_VPWR_M1014_s 0.00645603f $X=3.295 $Y=2.095 $X2=0
+ $Y2=0
cc_151 N_A_242_23#_M1000_g N_VPWR_c_398_n 0.0148577f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_242_23#_M1006_g N_VPWR_c_398_n 0.00172252f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A_242_23#_M1000_g N_VPWR_c_399_n 0.00172252f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_154 N_A_242_23#_M1006_g N_VPWR_c_399_n 0.0129203f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_242_23#_M1013_g N_VPWR_c_399_n 0.013023f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_242_23#_M1014_g N_VPWR_c_399_n 0.00196407f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_242_23#_M1013_g N_VPWR_c_400_n 0.00486043f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A_242_23#_M1014_g N_VPWR_c_400_n 0.0036352f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A_242_23#_M1013_g N_VPWR_c_401_n 0.00135454f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_242_23#_M1014_g N_VPWR_c_401_n 0.00948316f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_242_23#_M1000_g N_VPWR_c_406_n 0.00486043f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_242_23#_M1006_g N_VPWR_c_406_n 0.00486043f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_242_23#_c_130_n N_VPWR_c_408_n 0.0339406f $X=4.3 $Y=2.91 $X2=0 $Y2=0
cc_164 N_A_242_23#_M1001_d N_VPWR_c_397_n 0.00360572f $X=3.155 $Y=1.835 $X2=0
+ $Y2=0
cc_165 N_A_242_23#_M1007_d N_VPWR_c_397_n 0.00371702f $X=4.16 $Y=1.835 $X2=0
+ $Y2=0
cc_166 N_A_242_23#_M1000_g N_VPWR_c_397_n 0.00462979f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_242_23#_M1006_g N_VPWR_c_397_n 0.00462979f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_242_23#_M1013_g N_VPWR_c_397_n 0.00462979f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_242_23#_M1014_g N_VPWR_c_397_n 0.00436741f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_242_23#_c_130_n N_VPWR_c_397_n 0.0187779f $X=4.3 $Y=2.91 $X2=0 $Y2=0
cc_171 N_A_242_23#_M1002_g N_X_c_467_n 0.0125982f $X=1.285 $Y=0.665 $X2=0 $Y2=0
cc_172 N_A_242_23#_c_204_p N_X_c_467_n 0.0128525f $X=2.625 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A_242_23#_M1002_g N_X_c_468_n 0.0165573f $X=1.285 $Y=0.665 $X2=0 $Y2=0
cc_174 N_A_242_23#_c_204_p N_X_c_468_n 0.00192511f $X=2.625 $Y=1.51 $X2=0 $Y2=0
cc_175 N_A_242_23#_M1003_g N_X_c_470_n 0.0141561f $X=1.715 $Y=0.665 $X2=0 $Y2=0
cc_176 N_A_242_23#_M1008_g N_X_c_470_n 0.0138236f $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_177 N_A_242_23#_M1012_g N_X_c_470_n 0.00131418f $X=2.575 $Y=0.665 $X2=0 $Y2=0
cc_178 N_A_242_23#_c_204_p N_X_c_470_n 0.0593934f $X=2.625 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A_242_23#_c_117_n N_X_c_470_n 0.00641961f $X=2.71 $Y=1.425 $X2=0 $Y2=0
cc_180 N_A_242_23#_c_212_p N_X_c_470_n 0.00750776f $X=2.795 $Y=1.08 $X2=0 $Y2=0
cc_181 N_A_242_23#_c_124_n N_X_c_470_n 0.00500423f $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A_242_23#_c_204_p N_X_c_471_n 0.0177796f $X=2.625 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A_242_23#_c_124_n N_X_c_471_n 0.00255521f $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_184 N_A_242_23#_M1000_g N_X_c_473_n 0.0150311f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_242_23#_M1006_g N_X_c_473_n 0.0131615f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_242_23#_M1013_g N_X_c_473_n 0.0132057f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A_242_23#_c_204_p N_X_c_473_n 0.0678136f $X=2.625 $Y=1.51 $X2=0 $Y2=0
cc_188 N_A_242_23#_c_118_n N_X_c_473_n 0.00448013f $X=2.71 $Y=1.93 $X2=0 $Y2=0
cc_189 N_A_242_23#_c_124_n N_X_c_473_n 0.00729892f $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A_242_23#_c_212_p N_VGND_M1012_s 9.73829e-19 $X=2.795 $Y=1.08 $X2=0
+ $Y2=0
cc_191 N_A_242_23#_c_122_n N_VGND_M1012_s 0.0026801f $X=3.33 $Y=0.71 $X2=0 $Y2=0
cc_192 N_A_242_23#_M1002_g N_VGND_c_519_n 0.00328513f $X=1.285 $Y=0.665 $X2=0
+ $Y2=0
cc_193 N_A_242_23#_M1002_g N_VGND_c_520_n 6.28047e-19 $X=1.285 $Y=0.665 $X2=0
+ $Y2=0
cc_194 N_A_242_23#_M1003_g N_VGND_c_520_n 0.0108141f $X=1.715 $Y=0.665 $X2=0
+ $Y2=0
cc_195 N_A_242_23#_M1008_g N_VGND_c_520_n 0.010876f $X=2.145 $Y=0.665 $X2=0
+ $Y2=0
cc_196 N_A_242_23#_M1012_g N_VGND_c_520_n 6.39121e-19 $X=2.575 $Y=0.665 $X2=0
+ $Y2=0
cc_197 N_A_242_23#_M1012_g N_VGND_c_521_n 0.00524422f $X=2.575 $Y=0.665 $X2=0
+ $Y2=0
cc_198 N_A_242_23#_c_212_p N_VGND_c_521_n 0.00793424f $X=2.795 $Y=1.08 $X2=0
+ $Y2=0
cc_199 N_A_242_23#_c_122_n N_VGND_c_521_n 0.0181065f $X=3.33 $Y=0.71 $X2=0 $Y2=0
cc_200 N_A_242_23#_M1002_g N_VGND_c_524_n 0.00575161f $X=1.285 $Y=0.665 $X2=0
+ $Y2=0
cc_201 N_A_242_23#_M1003_g N_VGND_c_524_n 0.00477554f $X=1.715 $Y=0.665 $X2=0
+ $Y2=0
cc_202 N_A_242_23#_M1008_g N_VGND_c_526_n 0.00477554f $X=2.145 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_242_23#_M1012_g N_VGND_c_526_n 0.00575161f $X=2.575 $Y=0.665 $X2=0
+ $Y2=0
cc_204 N_A_242_23#_c_119_n N_VGND_c_528_n 0.0121867f $X=4.52 $Y=0.71 $X2=0 $Y2=0
cc_205 N_A_242_23#_c_120_n N_VGND_c_528_n 0.0746856f $X=3.785 $Y=0.71 $X2=0
+ $Y2=0
cc_206 N_A_242_23#_M1010_d N_VGND_c_529_n 0.00212318f $X=4.125 $Y=0.245 $X2=0
+ $Y2=0
cc_207 N_A_242_23#_M1002_g N_VGND_c_529_n 0.0118487f $X=1.285 $Y=0.665 $X2=0
+ $Y2=0
cc_208 N_A_242_23#_M1003_g N_VGND_c_529_n 0.00825815f $X=1.715 $Y=0.665 $X2=0
+ $Y2=0
cc_209 N_A_242_23#_M1008_g N_VGND_c_529_n 0.00825815f $X=2.145 $Y=0.665 $X2=0
+ $Y2=0
cc_210 N_A_242_23#_M1012_g N_VGND_c_529_n 0.0110121f $X=2.575 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_242_23#_c_119_n N_VGND_c_529_n 0.00660921f $X=4.52 $Y=0.71 $X2=0
+ $Y2=0
cc_212 N_A_242_23#_c_120_n N_VGND_c_529_n 0.0447855f $X=3.785 $Y=0.71 $X2=0
+ $Y2=0
cc_213 N_A_242_23#_c_120_n A_645_49# 0.00889726f $X=3.785 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_214 N_A_242_23#_c_122_n A_645_49# 0.00179331f $X=3.33 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A_242_23#_c_119_n A_717_49# 0.00170656f $X=4.52 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A_242_23#_c_120_n A_717_49# 0.0023191f $X=3.785 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_217 N_C_M1011_g N_B_M1004_g 0.0483068f $X=3.15 $Y=0.665 $X2=0 $Y2=0
cc_218 N_C_M1001_g N_B_M1005_g 0.0539248f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_219 N_C_c_250_n N_B_c_290_n 0.0483068f $X=3.06 $Y=1.51 $X2=0 $Y2=0
cc_220 N_C_c_251_n N_B_c_290_n 0.00128896f $X=3.06 $Y=1.51 $X2=0 $Y2=0
cc_221 N_C_M1001_g N_B_c_291_n 2.0072e-19 $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_222 N_C_c_250_n N_B_c_291_n 9.75099e-19 $X=3.06 $Y=1.51 $X2=0 $Y2=0
cc_223 N_C_c_251_n N_B_c_291_n 0.0328813f $X=3.06 $Y=1.51 $X2=0 $Y2=0
cc_224 N_C_M1001_g N_A_49_133#_c_346_n 0.0129331f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_225 N_C_M1001_g N_VPWR_c_401_n 0.00325225f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_226 N_C_M1001_g N_VPWR_c_402_n 0.00437171f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_227 N_C_M1001_g N_VPWR_c_403_n 0.00141133f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_228 N_C_M1001_g N_VPWR_c_397_n 0.00633763f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_229 N_C_M1011_g N_VGND_c_521_n 0.00657275f $X=3.15 $Y=0.665 $X2=0 $Y2=0
cc_230 N_C_M1011_g N_VGND_c_528_n 0.00575161f $X=3.15 $Y=0.665 $X2=0 $Y2=0
cc_231 N_C_M1011_g N_VGND_c_529_n 0.010916f $X=3.15 $Y=0.665 $X2=0 $Y2=0
cc_232 N_B_M1004_g N_A_49_133#_M1010_g 0.0376659f $X=3.51 $Y=0.665 $X2=0 $Y2=0
cc_233 N_B_c_290_n N_A_49_133#_c_322_n 0.0184515f $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_234 N_B_c_291_n N_A_49_133#_c_322_n 2.91848e-19 $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_235 N_B_M1005_g N_A_49_133#_M1007_g 0.032992f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_236 N_B_c_291_n N_A_49_133#_M1007_g 2.01271e-19 $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_237 N_B_M1005_g N_A_49_133#_c_346_n 0.0175798f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B_M1005_g N_A_49_133#_c_324_n 0.00969841f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B_c_291_n N_A_49_133#_c_324_n 0.00807248f $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_240 N_B_M1004_g N_A_49_133#_c_325_n 2.05149e-19 $X=3.51 $Y=0.665 $X2=0 $Y2=0
cc_241 N_B_c_290_n N_A_49_133#_c_325_n 0.00209704f $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_242 N_B_c_291_n N_A_49_133#_c_325_n 0.0241398f $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_243 N_B_M1005_g N_VPWR_c_402_n 0.0036352f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B_M1005_g N_VPWR_c_403_n 0.0101666f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B_M1005_g N_VPWR_c_397_n 0.00439469f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B_M1004_g N_VGND_c_528_n 0.00351226f $X=3.51 $Y=0.665 $X2=0 $Y2=0
cc_247 N_B_M1004_g N_VGND_c_529_n 0.00542362f $X=3.51 $Y=0.665 $X2=0 $Y2=0
cc_248 N_A_49_133#_c_329_n N_VPWR_M1009_d 0.00628441f $X=2.265 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_249 N_A_49_133#_c_329_n N_VPWR_M1006_s 0.00342847f $X=2.265 $Y=2.4 $X2=0
+ $Y2=0
cc_250 N_A_49_133#_c_346_n N_VPWR_M1014_s 0.00506052f $X=3.865 $Y=2.52 $X2=0
+ $Y2=0
cc_251 N_A_49_133#_c_346_n N_VPWR_M1005_d 0.012983f $X=3.865 $Y=2.52 $X2=0 $Y2=0
cc_252 N_A_49_133#_c_324_n N_VPWR_M1005_d 0.00774256f $X=3.95 $Y=2.43 $X2=0
+ $Y2=0
cc_253 N_A_49_133#_c_329_n N_VPWR_c_398_n 0.021529f $X=2.265 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A_49_133#_c_329_n N_VPWR_c_399_n 0.016709f $X=2.265 $Y=2.4 $X2=0 $Y2=0
cc_255 N_A_49_133#_c_346_n N_VPWR_c_400_n 0.00204011f $X=3.865 $Y=2.52 $X2=0
+ $Y2=0
cc_256 N_A_49_133#_c_375_p N_VPWR_c_400_n 0.00269838f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_257 N_A_49_133#_c_346_n N_VPWR_c_401_n 0.0206179f $X=3.865 $Y=2.52 $X2=0
+ $Y2=0
cc_258 N_A_49_133#_c_346_n N_VPWR_c_402_n 0.00743264f $X=3.865 $Y=2.52 $X2=0
+ $Y2=0
cc_259 N_A_49_133#_M1007_g N_VPWR_c_403_n 0.0061506f $X=4.085 $Y=2.465 $X2=0
+ $Y2=0
cc_260 N_A_49_133#_c_346_n N_VPWR_c_403_n 0.0212022f $X=3.865 $Y=2.52 $X2=0
+ $Y2=0
cc_261 N_A_49_133#_M1007_g N_VPWR_c_408_n 0.0056066f $X=4.085 $Y=2.465 $X2=0
+ $Y2=0
cc_262 N_A_49_133#_c_346_n N_VPWR_c_408_n 0.00182519f $X=3.865 $Y=2.52 $X2=0
+ $Y2=0
cc_263 N_A_49_133#_M1007_g N_VPWR_c_397_n 0.0115363f $X=4.085 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A_49_133#_c_329_n N_VPWR_c_397_n 0.0390492f $X=2.265 $Y=2.4 $X2=0 $Y2=0
cc_265 N_A_49_133#_c_330_n N_VPWR_c_397_n 0.00977402f $X=0.455 $Y=2.4 $X2=0
+ $Y2=0
cc_266 N_A_49_133#_c_346_n N_VPWR_c_397_n 0.0254104f $X=3.865 $Y=2.52 $X2=0
+ $Y2=0
cc_267 N_A_49_133#_c_375_p N_VPWR_c_397_n 0.00515293f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_268 N_A_49_133#_c_329_n N_X_M1000_d 0.00503872f $X=2.265 $Y=2.4 $X2=0 $Y2=0
cc_269 N_A_49_133#_c_375_p N_X_M1013_d 0.00493947f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_270 N_A_49_133#_c_323_n N_X_c_467_n 8.91818e-19 $X=0.37 $Y=0.875 $X2=0 $Y2=0
cc_271 N_A_49_133#_c_329_n N_X_c_467_n 0.0136682f $X=2.265 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A_49_133#_c_329_n N_X_c_473_n 0.0573951f $X=2.265 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A_49_133#_c_375_p N_X_c_473_n 0.0132692f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_274 N_A_49_133#_c_323_n N_VGND_c_522_n 0.00421272f $X=0.37 $Y=0.875 $X2=0
+ $Y2=0
cc_275 N_A_49_133#_M1010_g N_VGND_c_528_n 0.00351226f $X=4.05 $Y=0.665 $X2=0
+ $Y2=0
cc_276 N_A_49_133#_M1010_g N_VGND_c_529_n 0.0066798f $X=4.05 $Y=0.665 $X2=0
+ $Y2=0
cc_277 N_A_49_133#_c_323_n N_VGND_c_529_n 0.00717262f $X=0.37 $Y=0.875 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_397_n N_X_M1000_d 0.00412982f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_279 N_VPWR_c_397_n N_X_M1013_d 0.00366139f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_280 N_VPWR_M1009_d N_X_c_467_n 0.00568373f $X=0.68 $Y=1.835 $X2=0 $Y2=0
cc_281 N_VPWR_M1006_s N_X_c_473_n 0.00180541f $X=1.79 $Y=1.835 $X2=0 $Y2=0
cc_282 N_X_c_469_n N_VGND_M1015_d 0.00197782f $X=1.155 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_283 N_X_c_470_n N_VGND_M1003_s 0.00180746f $X=2.265 $Y=1.16 $X2=0 $Y2=0
cc_284 N_X_c_469_n N_VGND_c_519_n 0.0151472f $X=1.155 $Y=1.16 $X2=0 $Y2=0
cc_285 N_X_c_470_n N_VGND_c_520_n 0.0163515f $X=2.265 $Y=1.16 $X2=0 $Y2=0
cc_286 N_X_c_513_p N_VGND_c_524_n 0.0138717f $X=1.5 $Y=0.42 $X2=0 $Y2=0
cc_287 N_X_c_514_p N_VGND_c_526_n 0.0124525f $X=2.36 $Y=0.42 $X2=0 $Y2=0
cc_288 N_X_M1002_d N_VGND_c_529_n 0.00397496f $X=1.36 $Y=0.245 $X2=0 $Y2=0
cc_289 N_X_M1008_d N_VGND_c_529_n 0.00536646f $X=2.22 $Y=0.245 $X2=0 $Y2=0
cc_290 N_X_c_513_p N_VGND_c_529_n 0.00886411f $X=1.5 $Y=0.42 $X2=0 $Y2=0
cc_291 N_X_c_514_p N_VGND_c_529_n 0.00730901f $X=2.36 $Y=0.42 $X2=0 $Y2=0
cc_292 N_VGND_c_529_n A_645_49# 0.00534151f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
cc_293 N_VGND_c_529_n A_717_49# 0.00313651f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
