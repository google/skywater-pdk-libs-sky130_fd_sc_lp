* File: sky130_fd_sc_lp__a211o_2.pex.spice
* Created: Fri Aug 28 09:47:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211O_2%A_80_21# 1 2 3 12 16 20 24 27 28 29 30 34 36
+ 40 46 49 50 52
c107 50 0 1.55843e-19 $X=1.105 $Y=1.51
r108 53 55 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.51
+ $X2=0.905 $Y2=1.51
r109 50 55 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.105 $Y=1.51
+ $X2=0.905 $Y2=1.51
r110 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=1.51 $X2=1.105 $Y2=1.51
r111 44 46 19.2813 $w=2.58e-07 $l=4.35e-07 $layer=LI1_cond $X=3.545 $Y=0.855
+ $X2=3.545 $Y2=0.42
r112 40 42 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=3.51 $Y=1.98
+ $X2=3.51 $Y2=2.95
r113 38 40 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.51 $Y=1.875
+ $X2=3.51 $Y2=1.98
r114 37 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0.94
+ $X2=2.53 $Y2=0.94
r115 36 44 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.415 $Y=0.94
+ $X2=3.545 $Y2=0.855
r116 36 37 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.415 $Y=0.94
+ $X2=2.695 $Y2=0.94
r117 32 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=0.855
+ $X2=2.53 $Y2=0.94
r118 32 34 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.53 $Y=0.855
+ $X2=2.53 $Y2=0.42
r119 31 49 10.4193 $w=3.22e-07 $l=3.64452e-07 $layer=LI1_cond $X=1.415 $Y=1.785
+ $X2=1.207 $Y2=1.51
r120 30 38 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.345 $Y=1.785
+ $X2=3.51 $Y2=1.875
r121 30 31 118.919 $w=1.78e-07 $l=1.93e-06 $layer=LI1_cond $X=3.345 $Y=1.785
+ $X2=1.415 $Y2=1.785
r122 28 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0.94
+ $X2=2.53 $Y2=0.94
r123 28 29 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.365 $Y=0.94
+ $X2=1.415 $Y2=0.94
r124 27 49 8.95589 $w=3.22e-07 $l=2.17991e-07 $layer=LI1_cond $X=1.33 $Y=1.345
+ $X2=1.207 $Y2=1.51
r125 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.33 $Y=1.025
+ $X2=1.415 $Y2=0.94
r126 26 27 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.33 $Y=1.025
+ $X2=1.33 $Y2=1.345
r127 22 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.905 $Y2=1.51
r128 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.905 $Y2=2.465
r129 18 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=1.51
r130 18 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=0.655
r131 14 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.675
+ $X2=0.475 $Y2=1.51
r132 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=1.675
+ $X2=0.475 $Y2=2.465
r133 10 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=1.51
r134 10 12 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=0.655
r135 3 42 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=1.835 $X2=3.51 $Y2=2.95
r136 3 40 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=1.835 $X2=3.51 $Y2=1.98
r137 2 46 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.37
+ $Y=0.235 $X2=3.51 $Y2=0.42
r138 1 34 91 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.235 $X2=2.53 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_2%A2 1 3 6 8 14
c37 8 0 2.03038e-19 $X=1.68 $Y=1.295
r38 11 14 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.68 $Y=1.36
+ $X2=1.855 $Y2=1.36
r39 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.36 $X2=1.68 $Y2=1.36
r40 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.525
+ $X2=1.855 $Y2=1.36
r41 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.855 $Y=1.525 $X2=1.855
+ $Y2=2.465
r42 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.195
+ $X2=1.855 $Y2=1.36
r43 1 3 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.855 $Y=1.195
+ $X2=1.855 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_2%A1 3 6 8 11 12 13
c37 6 0 4.71948e-20 $X=2.395 $Y=2.465
r38 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.35
+ $X2=2.305 $Y2=1.515
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.35
+ $X2=2.305 $Y2=1.185
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.305
+ $Y=1.35 $X2=2.305 $Y2=1.35
r41 8 12 5.22201 $w=3.18e-07 $l=1.45e-07 $layer=LI1_cond $X=2.16 $Y=1.355
+ $X2=2.305 $Y2=1.355
r42 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.395 $Y=2.465
+ $X2=2.395 $Y2=1.515
r43 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.215 $Y=0.655
+ $X2=2.215 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_2%B1 3 6 8 11 13
r32 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.35
+ $X2=2.845 $Y2=1.515
r33 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.35
+ $X2=2.845 $Y2=1.185
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.35 $X2=2.845 $Y2=1.35
r35 8 12 9.90381 $w=3.18e-07 $l=2.75e-07 $layer=LI1_cond $X=3.12 $Y=1.355
+ $X2=2.845 $Y2=1.355
r36 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.875 $Y=2.465
+ $X2=2.875 $Y2=1.515
r37 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.865 $Y=0.655
+ $X2=2.865 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_2%C1 1 3 6 8 13
r23 10 13 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=3.295 $Y=1.35
+ $X2=3.55 $Y2=1.35
r24 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.35 $X2=3.55 $Y2=1.35
r25 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.515
+ $X2=3.295 $Y2=1.35
r26 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.295 $Y=1.515
+ $X2=3.295 $Y2=2.465
r27 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.185
+ $X2=3.295 $Y2=1.35
r28 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.295 $Y=1.185
+ $X2=3.295 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_2%VPWR 1 2 3 10 12 18 24 26 28 33 43 44 50 53
r50 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r54 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r55 41 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 40 43 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 38 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=2.125 $Y2=3.33
r59 38 40 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 34 50 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.142 $Y2=3.33
r63 34 36 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 33 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.96 $Y=3.33
+ $X2=2.125 $Y2=3.33
r65 33 36 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 32 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r67 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r68 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 29 47 4.40339 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.192 $Y2=3.33
r70 29 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 28 50 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=1.142
+ $Y2=3.33
r72 28 31 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r73 26 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 26 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 22 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=3.33
r76 22 24 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=2.505
r77 18 21 29.9231 $w=2.83e-07 $l=7.4e-07 $layer=LI1_cond $X=1.142 $Y=2.21
+ $X2=1.142 $Y2=2.95
r78 16 50 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.142 $Y=3.245
+ $X2=1.142 $Y2=3.33
r79 16 21 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=1.142 $Y=3.245
+ $X2=1.142 $Y2=2.95
r80 12 15 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=0.24 $Y=1.98
+ $X2=0.24 $Y2=2.95
r81 10 47 3.03446 $w=2.9e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.192 $Y2=3.33
r82 10 15 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.95
r83 3 24 300 $w=1.7e-07 $l=7.61282e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.835 $X2=2.125 $Y2=2.505
r84 2 21 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.95
r85 2 18 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.21
r86 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r87 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_2%X 1 2 7 8 9 10 11 12 13 22
r17 13 40 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.69 $Y=2.775
+ $X2=0.69 $Y2=2.91
r18 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=2.405
+ $X2=0.69 $Y2=2.775
r19 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.69 $Y=1.98
+ $X2=0.69 $Y2=2.405
r20 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=1.665
+ $X2=0.69 $Y2=1.98
r21 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=1.295
+ $X2=0.69 $Y2=1.665
r22 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=0.925 $X2=0.69
+ $Y2=1.295
r23 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=0.555 $X2=0.69
+ $Y2=0.925
r24 7 22 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.69 $Y=0.555
+ $X2=0.69 $Y2=0.42
r25 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.91
r26 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=1.98
r27 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_2%A_303_367# 1 2 7 9 11 13 15
r25 13 20 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.625 $Y=2.225
+ $X2=2.625 $Y2=2.135
r26 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.625 $Y=2.225
+ $X2=2.625 $Y2=2.9
r27 12 18 4.77666 $w=1.8e-07 $l=1.58e-07 $layer=LI1_cond $X=1.79 $Y=2.135
+ $X2=1.632 $Y2=2.135
r28 11 20 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=2.135
+ $X2=2.625 $Y2=2.135
r29 11 12 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.46 $Y=2.135
+ $X2=1.79 $Y2=2.135
r30 7 18 2.72088 $w=3.15e-07 $l=9e-08 $layer=LI1_cond $X=1.632 $Y=2.225
+ $X2=1.632 $Y2=2.135
r31 7 9 25.0611 $w=3.13e-07 $l=6.85e-07 $layer=LI1_cond $X=1.632 $Y=2.225
+ $X2=1.632 $Y2=2.91
r32 2 20 400 $w=1.7e-07 $l=3.64349e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.835 $X2=2.625 $Y2=2.13
r33 2 15 400 $w=1.7e-07 $l=1.13987e-06 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.835 $X2=2.625 $Y2=2.9
r34 1 18 400 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.835 $X2=1.64 $Y2=2.13
r35 1 9 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.835 $X2=1.64 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_2%VGND 1 2 3 10 12 16 18 25 32 33 41 47 49
r53 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r54 45 47 10.6269 $w=7.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.68 $Y=0.3
+ $X2=1.805 $Y2=0.3
r55 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 43 45 0.621339 $w=7.68e-07 $l=4e-08 $layer=LI1_cond $X=1.64 $Y=0.3 $X2=1.68
+ $Y2=0.3
r57 40 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r58 39 43 6.83473 $w=7.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.2 $Y=0.3 $X2=1.64
+ $Y2=0.3
r59 39 41 11.8696 $w=7.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.2 $Y=0.3
+ $X2=0.995 $Y2=0.3
r60 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r61 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r62 33 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r63 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r64 30 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.08
+ $Y2=0
r65 30 32 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.6
+ $Y2=0
r66 29 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r67 28 47 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=1.805
+ $Y2=0
r68 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r69 25 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.08
+ $Y2=0
r70 25 28 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r71 24 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r72 24 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r73 23 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.995
+ $Y2=0
r74 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r75 21 36 4.40339 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.192
+ $Y2=0
r76 21 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.72
+ $Y2=0
r77 18 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r78 18 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r79 14 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0
r80 14 16 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.56
r81 10 36 3.03446 $w=2.9e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.192 $Y2=0
r82 10 12 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.38
r83 3 16 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.56
r84 2 43 91 $w=1.7e-07 $l=8.1037e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.235 $X2=1.64 $Y2=0.57
r85 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

