* File: sky130_fd_sc_lp__nand4bb_2.pxi.spice
* Created: Fri Aug 28 10:52:27 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4BB_2%B_N N_B_N_M1000_g N_B_N_M1015_g N_B_N_c_115_n
+ N_B_N_c_116_n N_B_N_c_117_n B_N B_N N_B_N_c_119_n
+ PM_SKY130_FD_SC_LP__NAND4BB_2%B_N
x_PM_SKY130_FD_SC_LP__NAND4BB_2%A_N N_A_N_M1016_g N_A_N_M1006_g N_A_N_c_148_n
+ N_A_N_c_149_n N_A_N_c_150_n A_N A_N N_A_N_c_152_n
+ PM_SKY130_FD_SC_LP__NAND4BB_2%A_N
x_PM_SKY130_FD_SC_LP__NAND4BB_2%A_223_49# N_A_223_49#_M1016_d
+ N_A_223_49#_M1006_d N_A_223_49#_M1008_g N_A_223_49#_M1003_g
+ N_A_223_49#_M1013_g N_A_223_49#_M1018_g N_A_223_49#_c_187_n
+ N_A_223_49#_c_188_n N_A_223_49#_c_189_n N_A_223_49#_c_197_n
+ N_A_223_49#_c_190_n N_A_223_49#_c_191_n N_A_223_49#_c_192_n
+ PM_SKY130_FD_SC_LP__NAND4BB_2%A_223_49#
x_PM_SKY130_FD_SC_LP__NAND4BB_2%A_27_373# N_A_27_373#_M1015_s
+ N_A_27_373#_M1000_s N_A_27_373#_M1005_g N_A_27_373#_M1001_g
+ N_A_27_373#_M1009_g N_A_27_373#_M1012_g N_A_27_373#_c_262_n
+ N_A_27_373#_c_270_n N_A_27_373#_c_263_n N_A_27_373#_c_272_n
+ N_A_27_373#_c_273_n N_A_27_373#_c_274_n N_A_27_373#_c_275_n
+ N_A_27_373#_c_307_n N_A_27_373#_c_264_n N_A_27_373#_c_265_n
+ N_A_27_373#_c_266_n N_A_27_373#_c_267_n
+ PM_SKY130_FD_SC_LP__NAND4BB_2%A_27_373#
x_PM_SKY130_FD_SC_LP__NAND4BB_2%C N_C_M1004_g N_C_M1019_g N_C_c_365_n
+ N_C_M1007_g N_C_c_366_n N_C_c_367_n N_C_c_368_n N_C_M1017_g C C
+ PM_SKY130_FD_SC_LP__NAND4BB_2%C
x_PM_SKY130_FD_SC_LP__NAND4BB_2%D N_D_c_423_n N_D_M1011_g N_D_c_417_n
+ N_D_c_418_n N_D_M1002_g N_D_c_426_n N_D_M1014_g N_D_M1010_g D D N_D_c_422_n
+ PM_SKY130_FD_SC_LP__NAND4BB_2%D
x_PM_SKY130_FD_SC_LP__NAND4BB_2%VPWR N_VPWR_M1000_d N_VPWR_M1003_s
+ N_VPWR_M1018_s N_VPWR_M1012_s N_VPWR_M1019_s N_VPWR_M1014_s N_VPWR_c_464_n
+ N_VPWR_c_465_n N_VPWR_c_466_n N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_469_n
+ N_VPWR_c_470_n N_VPWR_c_471_n N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n
+ N_VPWR_c_475_n VPWR N_VPWR_c_476_n N_VPWR_c_477_n N_VPWR_c_478_n
+ N_VPWR_c_479_n N_VPWR_c_480_n N_VPWR_c_481_n N_VPWR_c_463_n
+ PM_SKY130_FD_SC_LP__NAND4BB_2%VPWR
x_PM_SKY130_FD_SC_LP__NAND4BB_2%Y N_Y_M1008_d N_Y_M1003_d N_Y_M1001_d
+ N_Y_M1004_d N_Y_M1011_d N_Y_c_629_p N_Y_c_609_n N_Y_c_545_n N_Y_c_546_n
+ N_Y_c_551_n N_Y_c_552_n N_Y_c_613_n N_Y_c_615_n N_Y_c_547_n N_Y_c_554_n
+ N_Y_c_618_n N_Y_c_548_n N_Y_c_549_n Y Y PM_SKY130_FD_SC_LP__NAND4BB_2%Y
x_PM_SKY130_FD_SC_LP__NAND4BB_2%VGND N_VGND_M1015_d N_VGND_M1002_d
+ N_VGND_c_637_n N_VGND_c_638_n VGND N_VGND_c_639_n N_VGND_c_640_n
+ N_VGND_c_641_n N_VGND_c_642_n N_VGND_c_643_n
+ PM_SKY130_FD_SC_LP__NAND4BB_2%VGND
x_PM_SKY130_FD_SC_LP__NAND4BB_2%A_357_47# N_A_357_47#_M1008_s
+ N_A_357_47#_M1013_s N_A_357_47#_M1009_d N_A_357_47#_c_707_n
+ N_A_357_47#_c_713_n N_A_357_47#_c_715_n N_A_357_47#_c_708_n
+ N_A_357_47#_c_716_n PM_SKY130_FD_SC_LP__NAND4BB_2%A_357_47#
x_PM_SKY130_FD_SC_LP__NAND4BB_2%A_614_47# N_A_614_47#_M1005_s
+ N_A_614_47#_M1007_d N_A_614_47#_c_746_n
+ PM_SKY130_FD_SC_LP__NAND4BB_2%A_614_47#
x_PM_SKY130_FD_SC_LP__NAND4BB_2%A_821_47# N_A_821_47#_M1007_s
+ N_A_821_47#_M1017_s N_A_821_47#_M1010_s N_A_821_47#_c_765_n
+ N_A_821_47#_c_786_n N_A_821_47#_c_766_n N_A_821_47#_c_767_n
+ N_A_821_47#_c_768_n PM_SKY130_FD_SC_LP__NAND4BB_2%A_821_47#
cc_1 VNB N_B_N_M1000_g 0.0136599f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.075
cc_2 VNB N_B_N_c_115_n 0.0194856f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.775
cc_3 VNB N_B_N_c_116_n 0.0236573f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.28
cc_4 VNB N_B_N_c_117_n 0.0166738f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.445
cc_5 VNB B_N 0.00941401f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_B_N_c_119_n 0.0165169f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.94
cc_7 VNB N_A_N_M1006_g 0.0129556f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.455
cc_8 VNB N_A_N_c_148_n 0.0197192f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.775
cc_9 VNB N_A_N_c_149_n 0.0275044f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.28
cc_10 VNB N_A_N_c_150_n 0.0164114f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.445
cc_11 VNB A_N 0.0109774f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_12 VNB N_A_N_c_152_n 0.0185639f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.94
cc_13 VNB N_A_223_49#_M1008_g 0.0280382f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.775
cc_14 VNB N_A_223_49#_M1013_g 0.0226194f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.94
cc_15 VNB N_A_223_49#_c_187_n 0.0369125f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.295
cc_16 VNB N_A_223_49#_c_188_n 0.031985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_223_49#_c_189_n 0.0114809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_223_49#_c_190_n 0.00164208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_223_49#_c_191_n 0.00816022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_223_49#_c_192_n 0.0149334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_373#_M1005_g 0.0233277f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.775
cc_22 VNB N_A_27_373#_M1009_g 0.0267955f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.94
cc_23 VNB N_A_27_373#_c_262_n 0.0502498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_373#_c_263_n 0.00766971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_373#_c_264_n 0.00386753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_373#_c_265_n 0.0166914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_373#_c_266_n 0.00515346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_373#_c_267_n 0.0396819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_C_M1004_g 0.00677274f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.075
cc_30 VNB N_C_M1019_g 0.00844382f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.455
cc_31 VNB N_C_c_365_n 0.0204041f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.775
cc_32 VNB N_C_c_366_n 0.0215078f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_33 VNB N_C_c_367_n 0.0545104f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_34 VNB N_C_c_368_n 0.0164056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB C 0.00264221f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.94
cc_36 VNB N_D_c_417_n 0.0103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_D_c_418_n 0.00530688f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.775
cc_38 VNB N_D_M1002_g 0.0231295f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.94
cc_39 VNB N_D_M1010_g 0.0311025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB D 0.0120055f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.94
cc_41 VNB N_D_c_422_n 0.0474804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_463_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_545_n 0.00813267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_546_n 0.00327323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_547_n 0.00240309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_548_n 0.00648585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_549_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB Y 0.0031126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_637_n 7.46595e-19 $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.445
cc_50 VNB N_VGND_c_638_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_639_n 0.100854f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.925
cc_52 VNB N_VGND_c_640_n 0.0163305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_641_n 0.321849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_642_n 0.0229928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_643_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_357_47#_c_707_n 0.00263155f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_57 VNB N_A_357_47#_c_708_n 0.00253352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_614_47#_c_746_n 0.00807993f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.445
cc_59 VNB N_A_821_47#_c_765_n 0.00253352f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.28
cc_60 VNB N_A_821_47#_c_766_n 0.015414f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.94
cc_61 VNB N_A_821_47#_c_767_n 0.00361594f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.94
cc_62 VNB N_A_821_47#_c_768_n 0.0307328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VPB N_B_N_M1000_g 0.0336124f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.075
cc_64 VPB N_A_N_M1006_g 0.0264728f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.455
cc_65 VPB N_A_223_49#_M1003_g 0.0234845f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_66 VPB N_A_223_49#_M1018_g 0.0188922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_223_49#_c_187_n 0.0156811f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.295
cc_68 VPB N_A_223_49#_c_188_n 0.00476146f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_223_49#_c_197_n 0.0152012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_223_49#_c_190_n 0.00285119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_27_373#_M1001_g 0.0189206f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_72 VPB N_A_27_373#_M1012_g 0.0180918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_27_373#_c_270_n 0.0199438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_27_373#_c_263_n 0.00964028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_27_373#_c_272_n 0.00106573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_27_373#_c_273_n 0.0216253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_27_373#_c_274_n 0.00482359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_27_373#_c_275_n 0.00165358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_27_373#_c_266_n 0.00640089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_C_M1004_g 0.0180918f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.075
cc_81 VPB N_C_M1019_g 0.0186849f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.455
cc_82 VPB N_D_c_423_n 0.0182173f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.445
cc_83 VPB N_D_c_417_n 0.00819946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_D_c_418_n 0.00204547f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.775
cc_85 VPB N_D_c_426_n 0.0233104f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.28
cc_86 VPB D 0.0131726f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=0.94
cc_87 VPB N_D_c_422_n 0.0186876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_464_n 0.0596488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_465_n 0.0187497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_466_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_467_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_468_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_469_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_470_n 0.0157625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_471_n 0.0484537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_472_n 0.032713f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_473_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_474_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_475_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_476_n 0.0199636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_477_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_478_n 0.0214572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_479_n 0.00449427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_480_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_481_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_463_n 0.0896102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_Y_c_551_n 0.00314908f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_Y_c_552_n 0.00214217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_Y_c_547_n 0.00256721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_Y_c_554_n 0.0016492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_Y_c_549_n 5.05803e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB Y 0.00339666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 N_B_N_M1000_g N_A_N_M1006_g 0.0145182f $X=0.475 $Y=2.075 $X2=0 $Y2=0
cc_114 N_B_N_c_115_n N_A_N_c_148_n 0.012977f $X=0.56 $Y=0.775 $X2=0 $Y2=0
cc_115 N_B_N_c_116_n N_A_N_c_149_n 0.0116433f $X=0.56 $Y=1.28 $X2=0 $Y2=0
cc_116 N_B_N_c_117_n N_A_N_c_150_n 0.0116433f $X=0.56 $Y=1.445 $X2=0 $Y2=0
cc_117 B_N A_N 0.0530546f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_118 N_B_N_c_119_n A_N 6.26206e-19 $X=0.56 $Y=0.94 $X2=0 $Y2=0
cc_119 B_N N_A_N_c_152_n 0.00452408f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_120 N_B_N_c_119_n N_A_N_c_152_n 0.0116433f $X=0.56 $Y=0.94 $X2=0 $Y2=0
cc_121 N_B_N_M1000_g N_A_27_373#_c_262_n 0.00674303f $X=0.475 $Y=2.075 $X2=0
+ $Y2=0
cc_122 N_B_N_c_115_n N_A_27_373#_c_262_n 0.00504932f $X=0.56 $Y=0.775 $X2=0
+ $Y2=0
cc_123 B_N N_A_27_373#_c_262_n 0.0516451f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_124 N_B_N_c_119_n N_A_27_373#_c_262_n 0.0163583f $X=0.56 $Y=0.94 $X2=0 $Y2=0
cc_125 N_B_N_M1000_g N_A_27_373#_c_270_n 0.00237971f $X=0.475 $Y=2.075 $X2=0
+ $Y2=0
cc_126 N_B_N_M1000_g N_A_27_373#_c_263_n 0.0193889f $X=0.475 $Y=2.075 $X2=0
+ $Y2=0
cc_127 N_B_N_c_117_n N_A_27_373#_c_263_n 0.00140616f $X=0.56 $Y=1.445 $X2=0
+ $Y2=0
cc_128 B_N N_A_27_373#_c_263_n 0.0291167f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_129 N_B_N_M1000_g N_A_27_373#_c_272_n 0.00175577f $X=0.475 $Y=2.075 $X2=0
+ $Y2=0
cc_130 B_N N_A_27_373#_c_265_n 0.00142887f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_131 N_B_N_c_119_n N_A_27_373#_c_265_n 0.00329303f $X=0.56 $Y=0.94 $X2=0 $Y2=0
cc_132 N_B_N_M1000_g N_VPWR_c_464_n 0.00392114f $X=0.475 $Y=2.075 $X2=0 $Y2=0
cc_133 N_B_N_c_115_n N_VGND_c_637_n 0.00943603f $X=0.56 $Y=0.775 $X2=0 $Y2=0
cc_134 B_N N_VGND_c_637_n 0.0105781f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_135 N_B_N_c_115_n N_VGND_c_641_n 0.00545225f $X=0.56 $Y=0.775 $X2=0 $Y2=0
cc_136 B_N N_VGND_c_641_n 0.00678029f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_137 N_B_N_c_115_n N_VGND_c_642_n 0.00477554f $X=0.56 $Y=0.775 $X2=0 $Y2=0
cc_138 N_B_N_c_119_n N_VGND_c_642_n 3.32067e-19 $X=0.56 $Y=0.94 $X2=0 $Y2=0
cc_139 N_A_N_M1006_g N_A_223_49#_c_187_n 0.00848125f $X=1.175 $Y=2.075 $X2=0
+ $Y2=0
cc_140 N_A_N_c_150_n N_A_223_49#_c_187_n 0.00662704f $X=1.13 $Y=1.445 $X2=0
+ $Y2=0
cc_141 A_N N_A_223_49#_c_187_n 3.4245e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_142 A_N N_A_223_49#_c_189_n 0.0110282f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_143 N_A_N_c_152_n N_A_223_49#_c_189_n 9.57425e-19 $X=1.13 $Y=0.94 $X2=0 $Y2=0
cc_144 N_A_N_M1006_g N_A_223_49#_c_197_n 4.51053e-19 $X=1.175 $Y=2.075 $X2=0
+ $Y2=0
cc_145 N_A_N_M1006_g N_A_223_49#_c_191_n 0.00803905f $X=1.175 $Y=2.075 $X2=0
+ $Y2=0
cc_146 N_A_N_c_149_n N_A_223_49#_c_191_n 0.00207953f $X=1.13 $Y=1.28 $X2=0 $Y2=0
cc_147 N_A_N_c_148_n N_A_223_49#_c_192_n 0.00432812f $X=1.13 $Y=0.775 $X2=0
+ $Y2=0
cc_148 A_N N_A_223_49#_c_192_n 0.0530324f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_149 N_A_N_c_152_n N_A_223_49#_c_192_n 0.00207953f $X=1.13 $Y=0.94 $X2=0 $Y2=0
cc_150 N_A_N_M1006_g N_A_27_373#_c_263_n 0.0063289f $X=1.175 $Y=2.075 $X2=0
+ $Y2=0
cc_151 N_A_N_c_150_n N_A_27_373#_c_263_n 0.00309338f $X=1.13 $Y=1.445 $X2=0
+ $Y2=0
cc_152 A_N N_A_27_373#_c_263_n 0.00998813f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_153 N_A_N_M1006_g N_A_27_373#_c_272_n 0.018013f $X=1.175 $Y=2.075 $X2=0 $Y2=0
cc_154 N_A_N_M1006_g N_A_27_373#_c_273_n 0.00929412f $X=1.175 $Y=2.075 $X2=0
+ $Y2=0
cc_155 N_A_N_M1006_g N_A_27_373#_c_274_n 0.00163211f $X=1.175 $Y=2.075 $X2=0
+ $Y2=0
cc_156 N_A_N_M1006_g N_VPWR_c_464_n 0.00131163f $X=1.175 $Y=2.075 $X2=0 $Y2=0
cc_157 N_A_N_c_148_n N_VGND_c_637_n 0.0102414f $X=1.13 $Y=0.775 $X2=0 $Y2=0
cc_158 N_A_N_c_148_n N_VGND_c_639_n 0.00477554f $X=1.13 $Y=0.775 $X2=0 $Y2=0
cc_159 N_A_N_c_152_n N_VGND_c_639_n 3.89791e-19 $X=1.13 $Y=0.94 $X2=0 $Y2=0
cc_160 N_A_N_c_148_n N_VGND_c_641_n 0.00654451f $X=1.13 $Y=0.775 $X2=0 $Y2=0
cc_161 A_N N_VGND_c_641_n 0.00526159f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_162 N_A_223_49#_M1013_g N_A_27_373#_M1005_g 0.0239765f $X=2.555 $Y=0.655
+ $X2=0 $Y2=0
cc_163 N_A_223_49#_c_188_n N_A_27_373#_M1001_g 0.0249914f $X=2.635 $Y=1.49 $X2=0
+ $Y2=0
cc_164 N_A_223_49#_c_190_n N_A_27_373#_c_263_n 0.00850128f $X=1.56 $Y=1.845
+ $X2=0 $Y2=0
cc_165 N_A_223_49#_c_197_n N_A_27_373#_c_272_n 0.012028f $X=1.39 $Y=2.01 $X2=0
+ $Y2=0
cc_166 N_A_223_49#_c_190_n N_A_27_373#_c_272_n 0.00221907f $X=1.56 $Y=1.845
+ $X2=0 $Y2=0
cc_167 N_A_223_49#_M1003_g N_A_27_373#_c_273_n 0.00618257f $X=2.205 $Y=2.465
+ $X2=0 $Y2=0
cc_168 N_A_223_49#_c_187_n N_A_27_373#_c_273_n 0.00446267f $X=2.05 $Y=1.49 $X2=0
+ $Y2=0
cc_169 N_A_223_49#_c_197_n N_A_27_373#_c_273_n 0.0417242f $X=1.39 $Y=2.01 $X2=0
+ $Y2=0
cc_170 N_A_223_49#_M1003_g N_A_27_373#_c_275_n 0.0194386f $X=2.205 $Y=2.465
+ $X2=0 $Y2=0
cc_171 N_A_223_49#_M1018_g N_A_27_373#_c_275_n 5.09517e-19 $X=2.635 $Y=2.465
+ $X2=0 $Y2=0
cc_172 N_A_223_49#_c_187_n N_A_27_373#_c_275_n 0.00319862f $X=2.05 $Y=1.49 $X2=0
+ $Y2=0
cc_173 N_A_223_49#_c_188_n N_A_27_373#_c_275_n 0.00637555f $X=2.635 $Y=1.49
+ $X2=0 $Y2=0
cc_174 N_A_223_49#_c_190_n N_A_27_373#_c_275_n 0.0477508f $X=1.56 $Y=1.845 $X2=0
+ $Y2=0
cc_175 N_A_223_49#_c_187_n N_A_27_373#_c_307_n 0.00577524f $X=2.05 $Y=1.49 $X2=0
+ $Y2=0
cc_176 N_A_223_49#_c_188_n N_A_27_373#_c_307_n 0.00737912f $X=2.635 $Y=1.49
+ $X2=0 $Y2=0
cc_177 N_A_223_49#_c_191_n N_A_27_373#_c_307_n 0.0155616f $X=1.7 $Y=1.49 $X2=0
+ $Y2=0
cc_178 N_A_223_49#_c_188_n N_A_27_373#_c_264_n 0.0320692f $X=2.635 $Y=1.49 $X2=0
+ $Y2=0
cc_179 N_A_223_49#_c_188_n N_A_27_373#_c_267_n 0.0235692f $X=2.635 $Y=1.49 $X2=0
+ $Y2=0
cc_180 N_A_223_49#_M1003_g N_VPWR_c_465_n 0.0109623f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_223_49#_M1018_g N_VPWR_c_465_n 5.60256e-19 $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_223_49#_M1003_g N_VPWR_c_466_n 7.24342e-19 $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_223_49#_M1018_g N_VPWR_c_466_n 0.0140971f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_223_49#_M1003_g N_VPWR_c_474_n 0.00486043f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A_223_49#_M1018_g N_VPWR_c_474_n 0.00486043f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A_223_49#_M1003_g N_VPWR_c_463_n 0.00824727f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_223_49#_M1018_g N_VPWR_c_463_n 0.00824727f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_223_49#_M1013_g N_Y_c_545_n 0.0119156f $X=2.555 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A_223_49#_c_188_n N_Y_c_545_n 0.00223526f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_190 N_A_223_49#_M1008_g N_Y_c_546_n 0.00218057f $X=2.125 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A_223_49#_c_188_n N_Y_c_546_n 0.00279547f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_192 N_A_223_49#_c_192_n N_Y_c_546_n 0.0039884f $X=1.645 $Y=1.325 $X2=0 $Y2=0
cc_193 N_A_223_49#_M1018_g N_Y_c_551_n 0.0134118f $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A_223_49#_M1003_g N_Y_c_552_n 7.79693e-19 $X=2.205 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A_223_49#_c_188_n N_Y_c_552_n 0.00292959f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_196 N_A_223_49#_M1008_g N_VGND_c_639_n 0.00357877f $X=2.125 $Y=0.655 $X2=0
+ $Y2=0
cc_197 N_A_223_49#_M1013_g N_VGND_c_639_n 0.00357842f $X=2.555 $Y=0.655 $X2=0
+ $Y2=0
cc_198 N_A_223_49#_c_189_n N_VGND_c_639_n 0.0285099f $X=1.56 $Y=0.44 $X2=0 $Y2=0
cc_199 N_A_223_49#_M1016_d N_VGND_c_641_n 0.00237724f $X=1.115 $Y=0.245 $X2=0
+ $Y2=0
cc_200 N_A_223_49#_M1008_g N_VGND_c_641_n 0.00681251f $X=2.125 $Y=0.655 $X2=0
+ $Y2=0
cc_201 N_A_223_49#_M1013_g N_VGND_c_641_n 0.00540059f $X=2.555 $Y=0.655 $X2=0
+ $Y2=0
cc_202 N_A_223_49#_c_189_n N_VGND_c_641_n 0.018304f $X=1.56 $Y=0.44 $X2=0 $Y2=0
cc_203 N_A_223_49#_M1008_g N_A_357_47#_c_707_n 0.00241433f $X=2.125 $Y=0.655
+ $X2=0 $Y2=0
cc_204 N_A_223_49#_c_187_n N_A_357_47#_c_707_n 0.00771551f $X=2.05 $Y=1.49 $X2=0
+ $Y2=0
cc_205 N_A_223_49#_c_189_n N_A_357_47#_c_707_n 0.0145897f $X=1.56 $Y=0.44 $X2=0
+ $Y2=0
cc_206 N_A_223_49#_c_192_n N_A_357_47#_c_707_n 0.0367095f $X=1.645 $Y=1.325
+ $X2=0 $Y2=0
cc_207 N_A_223_49#_M1008_g N_A_357_47#_c_713_n 0.012237f $X=2.125 $Y=0.655 $X2=0
+ $Y2=0
cc_208 N_A_223_49#_M1013_g N_A_357_47#_c_713_n 0.008403f $X=2.555 $Y=0.655 $X2=0
+ $Y2=0
cc_209 N_A_223_49#_c_189_n N_A_357_47#_c_715_n 0.0133514f $X=1.56 $Y=0.44 $X2=0
+ $Y2=0
cc_210 N_A_223_49#_M1008_g N_A_357_47#_c_716_n 3.91551e-19 $X=2.125 $Y=0.655
+ $X2=0 $Y2=0
cc_211 N_A_223_49#_M1013_g N_A_357_47#_c_716_n 0.00638661f $X=2.555 $Y=0.655
+ $X2=0 $Y2=0
cc_212 N_A_27_373#_c_267_n N_C_M1004_g 0.0209293f $X=3.495 $Y=1.485 $X2=0 $Y2=0
cc_213 N_A_27_373#_M1009_g N_C_c_367_n 0.0209293f $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A_27_373#_M1009_g C 2.28598e-19 $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_215 N_A_27_373#_c_272_n N_VPWR_M1000_d 0.00440581f $X=1.05 $Y=2.345 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A_27_373#_c_273_n N_VPWR_M1003_s 0.00512367f $X=1.985 $Y=2.43 $X2=0
+ $Y2=0
cc_217 N_A_27_373#_c_275_n N_VPWR_M1003_s 0.0100714f $X=2.07 $Y=2.345 $X2=0
+ $Y2=0
cc_218 N_A_27_373#_c_263_n N_VPWR_c_464_n 0.0172021f $X=0.965 $Y=1.71 $X2=0
+ $Y2=0
cc_219 N_A_27_373#_c_272_n N_VPWR_c_464_n 0.028414f $X=1.05 $Y=2.345 $X2=0 $Y2=0
cc_220 N_A_27_373#_c_274_n N_VPWR_c_464_n 0.0146817f $X=1.135 $Y=2.43 $X2=0
+ $Y2=0
cc_221 N_A_27_373#_c_273_n N_VPWR_c_465_n 0.0223246f $X=1.985 $Y=2.43 $X2=0
+ $Y2=0
cc_222 N_A_27_373#_M1001_g N_VPWR_c_466_n 0.0140971f $X=3.065 $Y=2.465 $X2=0
+ $Y2=0
cc_223 N_A_27_373#_M1012_g N_VPWR_c_466_n 7.24342e-19 $X=3.495 $Y=2.465 $X2=0
+ $Y2=0
cc_224 N_A_27_373#_M1001_g N_VPWR_c_467_n 0.00486043f $X=3.065 $Y=2.465 $X2=0
+ $Y2=0
cc_225 N_A_27_373#_M1012_g N_VPWR_c_467_n 0.00486043f $X=3.495 $Y=2.465 $X2=0
+ $Y2=0
cc_226 N_A_27_373#_M1001_g N_VPWR_c_468_n 7.28586e-19 $X=3.065 $Y=2.465 $X2=0
+ $Y2=0
cc_227 N_A_27_373#_M1012_g N_VPWR_c_468_n 0.0144091f $X=3.495 $Y=2.465 $X2=0
+ $Y2=0
cc_228 N_A_27_373#_M1001_g N_VPWR_c_463_n 0.00824727f $X=3.065 $Y=2.465 $X2=0
+ $Y2=0
cc_229 N_A_27_373#_M1012_g N_VPWR_c_463_n 0.00824727f $X=3.495 $Y=2.465 $X2=0
+ $Y2=0
cc_230 N_A_27_373#_c_273_n N_VPWR_c_463_n 0.0255484f $X=1.985 $Y=2.43 $X2=0
+ $Y2=0
cc_231 N_A_27_373#_c_274_n N_VPWR_c_463_n 0.00685203f $X=1.135 $Y=2.43 $X2=0
+ $Y2=0
cc_232 N_A_27_373#_M1005_g N_Y_c_545_n 0.0125841f $X=2.995 $Y=0.655 $X2=0 $Y2=0
cc_233 N_A_27_373#_M1009_g N_Y_c_545_n 0.00962275f $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_234 N_A_27_373#_c_264_n N_Y_c_545_n 0.05853f $X=3.085 $Y=1.485 $X2=0 $Y2=0
cc_235 N_A_27_373#_c_267_n N_Y_c_545_n 0.00469285f $X=3.495 $Y=1.485 $X2=0 $Y2=0
cc_236 N_A_27_373#_c_264_n N_Y_c_546_n 0.0181507f $X=3.085 $Y=1.485 $X2=0 $Y2=0
cc_237 N_A_27_373#_M1001_g N_Y_c_551_n 0.0136606f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A_27_373#_c_264_n N_Y_c_551_n 0.0482269f $X=3.085 $Y=1.485 $X2=0 $Y2=0
cc_239 N_A_27_373#_c_267_n N_Y_c_551_n 0.00202857f $X=3.495 $Y=1.485 $X2=0 $Y2=0
cc_240 N_A_27_373#_c_275_n N_Y_c_552_n 0.0105115f $X=2.07 $Y=2.345 $X2=0 $Y2=0
cc_241 N_A_27_373#_c_264_n N_Y_c_552_n 0.0154688f $X=3.085 $Y=1.485 $X2=0 $Y2=0
cc_242 N_A_27_373#_M1005_g Y 6.77067e-19 $X=2.995 $Y=0.655 $X2=0 $Y2=0
cc_243 N_A_27_373#_M1009_g Y 0.00393422f $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_244 N_A_27_373#_c_264_n Y 0.0151657f $X=3.085 $Y=1.485 $X2=0 $Y2=0
cc_245 N_A_27_373#_c_267_n Y 0.0125076f $X=3.495 $Y=1.485 $X2=0 $Y2=0
cc_246 N_A_27_373#_M1001_g Y 5.52814e-19 $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_247 N_A_27_373#_M1012_g Y 0.0152767f $X=3.495 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A_27_373#_c_264_n Y 0.00529238f $X=3.085 $Y=1.485 $X2=0 $Y2=0
cc_249 N_A_27_373#_c_267_n Y 0.00642554f $X=3.495 $Y=1.485 $X2=0 $Y2=0
cc_250 N_A_27_373#_M1005_g N_VGND_c_639_n 0.00357856f $X=2.995 $Y=0.655 $X2=0
+ $Y2=0
cc_251 N_A_27_373#_M1009_g N_VGND_c_639_n 0.00357877f $X=3.495 $Y=0.655 $X2=0
+ $Y2=0
cc_252 N_A_27_373#_M1015_s N_VGND_c_641_n 0.00237724f $X=0.27 $Y=0.245 $X2=0
+ $Y2=0
cc_253 N_A_27_373#_M1005_g N_VGND_c_641_n 0.00558488f $X=2.995 $Y=0.655 $X2=0
+ $Y2=0
cc_254 N_A_27_373#_M1009_g N_VGND_c_641_n 0.00683518f $X=3.495 $Y=0.655 $X2=0
+ $Y2=0
cc_255 N_A_27_373#_c_265_n N_VGND_c_641_n 0.0152848f $X=0.395 $Y=0.44 $X2=0
+ $Y2=0
cc_256 N_A_27_373#_c_265_n N_VGND_c_642_n 0.0237112f $X=0.395 $Y=0.44 $X2=0
+ $Y2=0
cc_257 N_A_27_373#_c_307_n N_A_357_47#_c_707_n 0.00177712f $X=2.155 $Y=1.472
+ $X2=0 $Y2=0
cc_258 N_A_27_373#_M1005_g N_A_357_47#_c_708_n 0.0103448f $X=2.995 $Y=0.655
+ $X2=0 $Y2=0
cc_259 N_A_27_373#_M1009_g N_A_357_47#_c_708_n 0.00923113f $X=3.495 $Y=0.655
+ $X2=0 $Y2=0
cc_260 N_A_27_373#_M1005_g N_A_357_47#_c_716_n 0.00559453f $X=2.995 $Y=0.655
+ $X2=0 $Y2=0
cc_261 N_A_27_373#_M1009_g N_A_357_47#_c_716_n 5.59125e-19 $X=3.495 $Y=0.655
+ $X2=0 $Y2=0
cc_262 N_A_27_373#_M1009_g N_A_614_47#_c_746_n 0.012794f $X=3.495 $Y=0.655 $X2=0
+ $Y2=0
cc_263 N_C_M1019_g N_D_c_418_n 0.0240783f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_264 N_C_c_366_n N_D_c_418_n 0.0158972f $X=4.8 $Y=1.26 $X2=0 $Y2=0
cc_265 N_C_c_368_n N_D_M1002_g 0.0216905f $X=4.875 $Y=1.185 $X2=0 $Y2=0
cc_266 C N_D_M1002_g 5.59438e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_267 N_C_c_367_n N_D_c_422_n 0.00367671f $X=4.525 $Y=1.26 $X2=0 $Y2=0
cc_268 C N_D_c_422_n 0.00196364f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_269 N_C_M1004_g N_VPWR_c_468_n 0.0143521f $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_270 N_C_M1019_g N_VPWR_c_468_n 7.28586e-19 $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_271 N_C_M1004_g N_VPWR_c_469_n 7.69607e-19 $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_272 N_C_M1019_g N_VPWR_c_469_n 0.0173454f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_273 N_C_M1004_g N_VPWR_c_477_n 0.00486043f $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_274 N_C_M1019_g N_VPWR_c_477_n 0.00486043f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_275 N_C_M1004_g N_VPWR_c_463_n 0.00824727f $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_276 N_C_M1019_g N_VPWR_c_463_n 0.00824727f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_277 N_C_c_365_n N_Y_c_545_n 0.00361972f $X=4.445 $Y=1.185 $X2=0 $Y2=0
cc_278 N_C_c_367_n N_Y_c_545_n 5.83137e-19 $X=4.525 $Y=1.26 $X2=0 $Y2=0
cc_279 N_C_M1019_g N_Y_c_547_n 0.0140763f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_280 N_C_c_366_n N_Y_c_547_n 0.00402152f $X=4.8 $Y=1.26 $X2=0 $Y2=0
cc_281 N_C_c_367_n N_Y_c_547_n 0.0027281f $X=4.525 $Y=1.26 $X2=0 $Y2=0
cc_282 C N_Y_c_547_n 0.0302352f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_283 N_C_c_366_n N_Y_c_554_n 3.15974e-19 $X=4.8 $Y=1.26 $X2=0 $Y2=0
cc_284 N_C_M1004_g N_Y_c_548_n 0.0191633f $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_285 C N_Y_c_548_n 0.0139439f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_286 N_C_M1019_g N_Y_c_549_n 9.97365e-19 $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_287 N_C_c_367_n N_Y_c_549_n 0.00256759f $X=4.525 $Y=1.26 $X2=0 $Y2=0
cc_288 C N_Y_c_549_n 0.0156157f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_289 N_C_c_367_n Y 0.00570538f $X=4.525 $Y=1.26 $X2=0 $Y2=0
cc_290 C Y 0.0184086f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_291 N_C_c_368_n N_VGND_c_638_n 0.00109252f $X=4.875 $Y=1.185 $X2=0 $Y2=0
cc_292 N_C_c_365_n N_VGND_c_639_n 0.00357877f $X=4.445 $Y=1.185 $X2=0 $Y2=0
cc_293 N_C_c_368_n N_VGND_c_639_n 0.00357877f $X=4.875 $Y=1.185 $X2=0 $Y2=0
cc_294 N_C_c_365_n N_VGND_c_641_n 0.00665089f $X=4.445 $Y=1.185 $X2=0 $Y2=0
cc_295 N_C_c_368_n N_VGND_c_641_n 0.00537654f $X=4.875 $Y=1.185 $X2=0 $Y2=0
cc_296 N_C_c_365_n N_A_614_47#_c_746_n 0.0136938f $X=4.445 $Y=1.185 $X2=0 $Y2=0
cc_297 N_C_c_366_n N_A_614_47#_c_746_n 0.0025871f $X=4.8 $Y=1.26 $X2=0 $Y2=0
cc_298 N_C_c_367_n N_A_614_47#_c_746_n 0.0119892f $X=4.525 $Y=1.26 $X2=0 $Y2=0
cc_299 N_C_c_368_n N_A_614_47#_c_746_n 0.00367457f $X=4.875 $Y=1.185 $X2=0 $Y2=0
cc_300 C N_A_614_47#_c_746_n 0.0310938f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_301 N_C_c_365_n N_A_821_47#_c_765_n 0.0086866f $X=4.445 $Y=1.185 $X2=0 $Y2=0
cc_302 N_C_c_368_n N_A_821_47#_c_765_n 0.0126515f $X=4.875 $Y=1.185 $X2=0 $Y2=0
cc_303 N_C_c_368_n N_A_821_47#_c_767_n 0.00470011f $X=4.875 $Y=1.185 $X2=0 $Y2=0
cc_304 C N_A_821_47#_c_767_n 0.00124306f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_305 N_D_c_423_n N_VPWR_c_469_n 0.0193907f $X=4.785 $Y=1.725 $X2=0 $Y2=0
cc_306 N_D_c_426_n N_VPWR_c_471_n 0.0224661f $X=5.595 $Y=1.725 $X2=0 $Y2=0
cc_307 D N_VPWR_c_471_n 0.0257069f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_308 N_D_c_422_n N_VPWR_c_471_n 0.00101486f $X=5.685 $Y=1.51 $X2=0 $Y2=0
cc_309 N_D_c_423_n N_VPWR_c_478_n 0.00486043f $X=4.785 $Y=1.725 $X2=0 $Y2=0
cc_310 N_D_c_426_n N_VPWR_c_478_n 0.00486043f $X=5.595 $Y=1.725 $X2=0 $Y2=0
cc_311 N_D_c_423_n N_VPWR_c_463_n 0.00895189f $X=4.785 $Y=1.725 $X2=0 $Y2=0
cc_312 N_D_c_426_n N_VPWR_c_463_n 0.00895189f $X=5.595 $Y=1.725 $X2=0 $Y2=0
cc_313 N_D_c_423_n N_Y_c_547_n 0.0077773f $X=4.785 $Y=1.725 $X2=0 $Y2=0
cc_314 N_D_c_417_n N_Y_c_547_n 0.00113014f $X=5.16 $Y=1.65 $X2=0 $Y2=0
cc_315 N_D_c_418_n N_Y_c_547_n 0.00503429f $X=4.86 $Y=1.65 $X2=0 $Y2=0
cc_316 N_D_c_423_n N_Y_c_554_n 0.00141051f $X=4.785 $Y=1.725 $X2=0 $Y2=0
cc_317 N_D_c_417_n N_Y_c_554_n 0.0123188f $X=5.16 $Y=1.65 $X2=0 $Y2=0
cc_318 N_D_c_426_n N_Y_c_554_n 0.00423318f $X=5.595 $Y=1.725 $X2=0 $Y2=0
cc_319 D N_Y_c_554_n 0.0152894f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_320 N_D_c_422_n N_Y_c_554_n 0.0152323f $X=5.685 $Y=1.51 $X2=0 $Y2=0
cc_321 N_D_M1002_g N_VGND_c_638_n 0.0124368f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_322 N_D_M1010_g N_VGND_c_638_n 0.0130588f $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_323 N_D_M1002_g N_VGND_c_639_n 0.00486043f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_324 N_D_M1010_g N_VGND_c_640_n 0.00486043f $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_325 N_D_M1002_g N_VGND_c_641_n 0.0082726f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_326 N_D_M1010_g N_VGND_c_641_n 0.00920706f $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_327 N_D_M1002_g N_A_821_47#_c_766_n 0.0172265f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_328 N_D_M1010_g N_A_821_47#_c_766_n 0.0155556f $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_329 D N_A_821_47#_c_766_n 0.0472013f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_330 N_D_c_422_n N_A_821_47#_c_766_n 0.00504716f $X=5.685 $Y=1.51 $X2=0 $Y2=0
cc_331 N_D_c_417_n N_A_821_47#_c_767_n 0.00305093f $X=5.16 $Y=1.65 $X2=0 $Y2=0
cc_332 N_D_c_422_n N_A_821_47#_c_767_n 7.29777e-19 $X=5.685 $Y=1.51 $X2=0 $Y2=0
cc_333 N_VPWR_c_463_n N_Y_M1003_d 0.00536646f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_334 N_VPWR_c_463_n N_Y_M1001_d 0.00536646f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_335 N_VPWR_c_463_n N_Y_M1004_d 0.00536646f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_336 N_VPWR_c_463_n N_Y_M1011_d 0.00852317f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_337 N_VPWR_c_474_n N_Y_c_609_n 0.0124525f $X=2.685 $Y=3.33 $X2=0 $Y2=0
cc_338 N_VPWR_c_463_n N_Y_c_609_n 0.00730901f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_339 N_VPWR_M1018_s N_Y_c_551_n 0.00183199f $X=2.71 $Y=1.835 $X2=0 $Y2=0
cc_340 N_VPWR_c_466_n N_Y_c_551_n 0.0160778f $X=2.85 $Y=2.27 $X2=0 $Y2=0
cc_341 N_VPWR_c_467_n N_Y_c_613_n 0.0124525f $X=3.545 $Y=3.33 $X2=0 $Y2=0
cc_342 N_VPWR_c_463_n N_Y_c_613_n 0.00730901f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_343 N_VPWR_c_477_n N_Y_c_615_n 0.0124525f $X=4.405 $Y=3.33 $X2=0 $Y2=0
cc_344 N_VPWR_c_463_n N_Y_c_615_n 0.00730901f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_345 N_VPWR_c_469_n N_Y_c_547_n 0.0216087f $X=4.57 $Y=2.03 $X2=0 $Y2=0
cc_346 N_VPWR_c_478_n N_Y_c_618_n 0.0391712f $X=5.645 $Y=3.33 $X2=0 $Y2=0
cc_347 N_VPWR_c_463_n N_Y_c_618_n 0.0220825f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_348 N_VPWR_M1012_s N_Y_c_548_n 0.00115923f $X=3.57 $Y=1.835 $X2=0 $Y2=0
cc_349 N_VPWR_c_468_n N_Y_c_548_n 0.0109948f $X=3.71 $Y=2.175 $X2=0 $Y2=0
cc_350 N_VPWR_M1012_s Y 6.41842e-19 $X=3.57 $Y=1.835 $X2=0 $Y2=0
cc_351 N_VPWR_c_468_n Y 0.00721868f $X=3.71 $Y=2.175 $X2=0 $Y2=0
cc_352 N_Y_M1008_d N_VGND_c_641_n 0.00225186f $X=2.2 $Y=0.235 $X2=0 $Y2=0
cc_353 N_Y_c_545_n N_A_357_47#_M1013_s 0.00205023f $X=3.42 $Y=1.12 $X2=0 $Y2=0
cc_354 N_Y_c_545_n N_A_357_47#_M1009_d 0.0014901f $X=3.42 $Y=1.12 $X2=0 $Y2=0
cc_355 N_Y_c_546_n N_A_357_47#_c_707_n 0.00147129f $X=2.435 $Y=1.12 $X2=0 $Y2=0
cc_356 N_Y_M1008_d N_A_357_47#_c_713_n 0.00332344f $X=2.2 $Y=0.235 $X2=0 $Y2=0
cc_357 N_Y_c_629_p N_A_357_47#_c_713_n 0.0125296f $X=2.34 $Y=0.76 $X2=0 $Y2=0
cc_358 N_Y_c_545_n N_A_357_47#_c_713_n 0.00292867f $X=3.42 $Y=1.12 $X2=0 $Y2=0
cc_359 N_Y_c_545_n N_A_357_47#_c_708_n 0.00342201f $X=3.42 $Y=1.12 $X2=0 $Y2=0
cc_360 N_Y_c_545_n N_A_357_47#_c_716_n 0.0143984f $X=3.42 $Y=1.12 $X2=0 $Y2=0
cc_361 N_Y_c_545_n N_A_614_47#_M1005_s 0.00251484f $X=3.42 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_362 N_Y_c_545_n N_A_614_47#_c_746_n 0.033989f $X=3.42 $Y=1.12 $X2=0 $Y2=0
cc_363 N_Y_c_554_n N_A_821_47#_c_766_n 0.00340169f $X=5.19 $Y=2.205 $X2=0 $Y2=0
cc_364 N_Y_c_554_n N_A_821_47#_c_767_n 0.00942952f $X=5.19 $Y=2.205 $X2=0 $Y2=0
cc_365 N_VGND_c_641_n N_A_357_47#_M1008_s 0.00319523f $X=6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_366 N_VGND_c_641_n N_A_357_47#_M1013_s 0.00231601f $X=6 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_641_n N_A_357_47#_M1009_d 0.00215176f $X=6 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_639_n N_A_357_47#_c_713_n 0.0326395f $X=5.355 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_641_n N_A_357_47#_c_713_n 0.0208532f $X=6 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_639_n N_A_357_47#_c_715_n 0.0132962f $X=5.355 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_641_n N_A_357_47#_c_715_n 0.00777554f $X=6 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_639_n N_A_357_47#_c_708_n 0.0549136f $X=5.355 $Y=0 $X2=0 $Y2=0
cc_373 N_VGND_c_641_n N_A_357_47#_c_708_n 0.0341296f $X=6 $Y=0 $X2=0 $Y2=0
cc_374 N_VGND_c_639_n N_A_357_47#_c_716_n 0.0188918f $X=5.355 $Y=0 $X2=0 $Y2=0
cc_375 N_VGND_c_641_n N_A_357_47#_c_716_n 0.0124426f $X=6 $Y=0 $X2=0 $Y2=0
cc_376 N_VGND_c_641_n N_A_614_47#_M1005_s 0.00281482f $X=6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_377 N_VGND_c_641_n N_A_614_47#_M1007_d 0.00225186f $X=6 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_639_n N_A_614_47#_c_746_n 0.00353981f $X=5.355 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_641_n N_A_614_47#_c_746_n 0.00852678f $X=6 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_641_n N_A_821_47#_M1007_s 0.00215176f $X=6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_381 N_VGND_c_641_n N_A_821_47#_M1017_s 0.00376627f $X=6 $Y=0 $X2=0 $Y2=0
cc_382 N_VGND_c_641_n N_A_821_47#_M1010_s 0.00371702f $X=6 $Y=0 $X2=0 $Y2=0
cc_383 N_VGND_c_639_n N_A_821_47#_c_765_n 0.0529361f $X=5.355 $Y=0 $X2=0 $Y2=0
cc_384 N_VGND_c_641_n N_A_821_47#_c_765_n 0.033612f $X=6 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_c_639_n N_A_821_47#_c_786_n 0.0125234f $X=5.355 $Y=0 $X2=0 $Y2=0
cc_386 N_VGND_c_641_n N_A_821_47#_c_786_n 0.00738676f $X=6 $Y=0 $X2=0 $Y2=0
cc_387 N_VGND_M1002_d N_A_821_47#_c_766_n 0.00176461f $X=5.38 $Y=0.235 $X2=0
+ $Y2=0
cc_388 N_VGND_c_638_n N_A_821_47#_c_766_n 0.0170777f $X=5.52 $Y=0.38 $X2=0 $Y2=0
cc_389 N_VGND_c_640_n N_A_821_47#_c_768_n 0.0178111f $X=6 $Y=0 $X2=0 $Y2=0
cc_390 N_VGND_c_641_n N_A_821_47#_c_768_n 0.0100304f $X=6 $Y=0 $X2=0 $Y2=0
cc_391 N_A_357_47#_c_708_n N_A_614_47#_M1005_s 0.00476194f $X=3.71 $Y=0.38
+ $X2=-0.19 $Y2=-0.245
cc_392 N_A_357_47#_M1009_d N_A_614_47#_c_746_n 0.00978161f $X=3.57 $Y=0.235
+ $X2=0 $Y2=0
cc_393 N_A_357_47#_c_708_n N_A_614_47#_c_746_n 0.0446918f $X=3.71 $Y=0.38 $X2=0
+ $Y2=0
cc_394 N_A_357_47#_c_708_n N_A_821_47#_c_765_n 0.0180051f $X=3.71 $Y=0.38 $X2=0
+ $Y2=0
cc_395 N_A_614_47#_c_746_n N_A_821_47#_M1007_s 0.00572927f $X=4.66 $Y=0.75
+ $X2=-0.19 $Y2=-0.245
cc_396 N_A_614_47#_M1007_d N_A_821_47#_c_765_n 0.0033495f $X=4.52 $Y=0.235 $X2=0
+ $Y2=0
cc_397 N_A_614_47#_c_746_n N_A_821_47#_c_765_n 0.0413226f $X=4.66 $Y=0.75 $X2=0
+ $Y2=0
