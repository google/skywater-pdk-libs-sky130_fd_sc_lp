* File: sky130_fd_sc_lp__dlrtn_2.spice
* Created: Wed Sep  2 09:46:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrtn_2.pex.spice"
.subckt sky130_fd_sc_lp__dlrtn_2  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_D_M1003_g N_A_31_464#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_221_70#_M1004_d N_GATE_N_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_221_70#_M1018_g N_A_372_397#_M1018_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1019 A_554_125# N_A_31_464#_M1019_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1015 N_A_626_125#_M1015_d N_A_221_70#_M1015_g A_554_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.0735 AS=0.0441 PD=0.77 PS=0.63 NRD=19.992 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1016 A_726_125# N_A_372_397#_M1016_g N_A_626_125#_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0525 AS=0.0735 PD=0.67 PS=0.77 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_776_99#_M1021_g A_726_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0525 PD=1.37 PS=0.67 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 A_996_47# N_A_626_125#_M1017_g N_A_776_99#_M1017_s VNB NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_RESET_B_M1011_g A_996_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.0882 PD=1.23 PS=1.05 NRD=5.712 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1001 N_Q_M1001_d N_A_776_99#_M1001_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1638 PD=1.12 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1006 N_Q_M1001_d N_A_776_99#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_D_M1013_g N_A_31_464#_M1013_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1712 AS=0.1696 PD=1.175 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1005 N_A_221_70#_M1005_d N_GATE_N_M1005_g N_VPWR_M1013_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1792 AS=0.1712 PD=1.84 PS=1.175 NRD=4.6098 NRS=78.4848 M=1
+ R=4.26667 SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_221_70#_M1000_g N_A_372_397#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1248 AS=0.3254 PD=1.03 PS=2.76 NRD=16.9223 NRS=139.555 M=1
+ R=4.26667 SA=75000.3 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1007 A_582_473# N_A_31_464#_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1248 PD=0.85 PS=1.03 NRD=15.3857 NRS=16.9223 M=1 R=4.26667
+ SA=75000.8 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1009 N_A_626_125#_M1009_d N_A_372_397#_M1009_g A_582_473# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.138023 AS=0.0672 PD=1.24981 PS=0.85 NRD=6.1464 NRS=15.3857 M=1
+ R=4.26667 SA=75001.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1012 A_763_473# N_A_221_70#_M1012_g N_A_626_125#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0905774 PD=0.63 PS=0.820189 NRD=23.443 NRS=45.7237 M=1
+ R=2.8 SA=75001.7 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_776_99#_M1014_g A_763_473# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.124425 AS=0.0441 PD=0.9575 PS=0.63 NRD=113.157 NRS=23.443 M=1 R=2.8
+ SA=75002.1 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1002 N_A_776_99#_M1002_d N_A_626_125#_M1002_g N_VPWR_M1014_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.373275 PD=1.54 PS=2.8725 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_RESET_B_M1010_g N_A_776_99#_M1002_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_Q_M1008_d N_A_776_99#_M1008_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75002
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1020 N_Q_M1008_d N_A_776_99#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX22_noxref VNB VPB NWDIODE A=13.2415 P=17.93
c_148 VPB 0 1.48338e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlrtn_2.pxi.spice"
*
.ends
*
*
