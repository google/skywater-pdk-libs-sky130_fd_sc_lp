* File: sky130_fd_sc_lp__or4b_4.spice
* Created: Wed Sep  2 10:32:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4b_4.pex.spice"
.subckt sky130_fd_sc_lp__or4b_4  VNB VPB A B C D_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D_N	D_N
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_X_M1000_d N_A_83_21#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75004
+ A=0.126 P=1.98 MULT=1
MM1007 N_X_M1000_d N_A_83_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1008_d N_A_83_21#_M1008_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1012 N_X_M1008_d N_A_83_21#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.856 M=1 R=5.6 SA=75001.5
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1006 N_A_83_21#_M1006_d N_A_M1006_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.856 M=1 R=5.6 SA=75001.9
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_B_M1013_g N_A_83_21#_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1003 N_A_83_21#_M1003_d N_C_M1003_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2604 PD=1.12 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75003.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_737_315#_M1009_g N_A_83_21#_M1003_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2758 AS=0.1176 PD=2.08 PS=1.12 NRD=20.952 NRS=0 M=1 R=5.6
+ SA=75003.6 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_A_737_315#_M1017_d N_D_N_M1017_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1379 PD=1.37 PS=1.04 NRD=0 NRS=63.564 M=1 R=2.8
+ SA=75004.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_83_21#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_83_21#_M1005_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6 SB=75003
+ A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1005_d N_A_83_21#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A_83_21#_M1014_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.1764 PD=1.65 PS=1.54 NRD=8.5892 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1015 A_479_367# N_A_M1015_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.2457 PD=1.47 PS=1.65 NRD=7.8012 NRS=8.5892 M=1 R=8.4 SA=75002 SB=75001.6
+ A=0.189 P=2.82 MULT=1
MM1016 A_551_367# N_B_M1016_g A_479_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75002.4
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1004 A_659_367# N_C_M1004_g A_551_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.2457 PD=1.65 PS=1.65 NRD=21.8867 NRS=21.8867 M=1 R=8.4 SA=75002.9
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1010 N_A_83_21#_M1010_d N_A_737_315#_M1010_g A_659_367# VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4
+ SA=75003.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_A_737_315#_M1002_d N_D_N_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX18_noxref VNB VPB NWDIODE A=10.5559 P=15.05
c_54 VNB 0 1.31108e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__or4b_4.pxi.spice"
*
.ends
*
*
