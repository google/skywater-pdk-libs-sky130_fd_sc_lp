* File: sky130_fd_sc_lp__and3b_4.pex.spice
* Created: Fri Aug 28 10:06:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3B_4%A_N 3 6 8 9 10 11 12 19 21
r29 19 22 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.707 $Y=1.36
+ $X2=0.707 $Y2=1.525
r30 19 21 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.707 $Y=1.36
+ $X2=0.707 $Y2=1.195
r31 11 12 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=1.665
+ $X2=0.715 $Y2=2.035
r32 10 11 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=1.295
+ $X2=0.715 $Y2=1.665
r33 10 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.36 $X2=0.72 $Y2=1.36
r34 9 10 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.925
+ $X2=0.715 $Y2=1.295
r35 8 9 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.555
+ $X2=0.715 $Y2=0.925
r36 6 22 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.605 $Y=2.045
+ $X2=0.605 $Y2=1.525
r37 3 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.605 $Y=0.875
+ $X2=0.605 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_4%A_242_23# 1 2 3 12 16 20 24 28 32 36 40 42
+ 51 53 55 56 58 60 61 66 70 71 73 74 81
c136 40 0 3.47797e-19 $X=2.575 $Y=2.465
r137 78 79 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.715 $Y=1.51
+ $X2=2.145 $Y2=1.51
r138 73 74 9.42615 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=4.447 $Y=1.98
+ $X2=4.447 $Y2=1.815
r139 68 74 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.605 $Y=1.165
+ $X2=4.605 $Y2=1.815
r140 64 73 1.89893 $w=4.83e-07 $l=7.7e-08 $layer=LI1_cond $X=4.447 $Y=2.057
+ $X2=4.447 $Y2=1.98
r141 64 66 21.0362 $w=4.83e-07 $l=8.53e-07 $layer=LI1_cond $X=4.447 $Y=2.057
+ $X2=4.447 $Y2=2.91
r142 61 71 16.2203 $w=9.08e-07 $l=4.55e-07 $layer=LI1_cond $X=3.785 $Y=0.71
+ $X2=3.33 $Y2=0.71
r143 61 63 6.43516 $w=9.08e-07 $l=4.8e-07 $layer=LI1_cond $X=3.785 $Y=0.71
+ $X2=4.265 $Y2=0.71
r144 60 68 12.2187 $w=9.1e-07 $l=4.95681e-07 $layer=LI1_cond $X=4.52 $Y=0.71
+ $X2=4.605 $Y2=1.165
r145 60 63 3.41868 $w=9.08e-07 $l=2.55e-07 $layer=LI1_cond $X=4.52 $Y=0.71
+ $X2=4.265 $Y2=0.71
r146 56 58 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.795 $Y=2.095
+ $X2=3.295 $Y2=2.095
r147 55 71 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.795 $Y=1.08
+ $X2=3.33 $Y2=1.08
r148 53 56 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.71 $Y=1.93
+ $X2=2.795 $Y2=2.095
r149 52 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=1.595
+ $X2=2.71 $Y2=1.51
r150 52 53 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.71 $Y=1.595
+ $X2=2.71 $Y2=1.93
r151 51 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=1.425
+ $X2=2.71 $Y2=1.51
r152 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.71 $Y=1.165
+ $X2=2.795 $Y2=1.08
r153 50 51 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.71 $Y=1.165
+ $X2=2.71 $Y2=1.425
r154 49 81 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.52 $Y=1.51
+ $X2=2.575 $Y2=1.51
r155 49 79 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=2.52 $Y=1.51
+ $X2=2.145 $Y2=1.51
r156 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.51 $X2=2.52 $Y2=1.51
r157 45 78 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.5 $Y=1.51
+ $X2=1.715 $Y2=1.51
r158 45 75 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.5 $Y=1.51
+ $X2=1.285 $Y2=1.51
r159 44 48 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.5 $Y=1.51
+ $X2=2.52 $Y2=1.51
r160 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.5
+ $Y=1.51 $X2=1.5 $Y2=1.51
r161 42 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=1.51
+ $X2=2.71 $Y2=1.51
r162 42 48 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.625 $Y=1.51
+ $X2=2.52 $Y2=1.51
r163 38 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.675
+ $X2=2.575 $Y2=1.51
r164 38 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.575 $Y=1.675
+ $X2=2.575 $Y2=2.465
r165 34 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.345
+ $X2=2.575 $Y2=1.51
r166 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.575 $Y=1.345
+ $X2=2.575 $Y2=0.665
r167 30 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.145 $Y=1.675
+ $X2=2.145 $Y2=1.51
r168 30 32 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.145 $Y=1.675
+ $X2=2.145 $Y2=2.465
r169 26 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.145 $Y=1.345
+ $X2=2.145 $Y2=1.51
r170 26 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.145 $Y=1.345
+ $X2=2.145 $Y2=0.665
r171 22 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.675
+ $X2=1.715 $Y2=1.51
r172 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.715 $Y=1.675
+ $X2=1.715 $Y2=2.465
r173 18 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.345
+ $X2=1.715 $Y2=1.51
r174 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.715 $Y=1.345
+ $X2=1.715 $Y2=0.665
r175 14 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.675
+ $X2=1.285 $Y2=1.51
r176 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.285 $Y=1.675
+ $X2=1.285 $Y2=2.465
r177 10 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.345
+ $X2=1.285 $Y2=1.51
r178 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.285 $Y=1.345
+ $X2=1.285 $Y2=0.665
r179 3 73 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=1.835 $X2=4.3 $Y2=1.98
r180 3 66 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=1.835 $X2=4.3 $Y2=2.91
r181 2 58 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=1.835 $X2=3.295 $Y2=2.095
r182 1 63 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=4.125
+ $Y=0.245 $X2=4.265 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_4%C 3 7 9 12 13
c40 13 0 1.94442e-19 $X=3.06 $Y=1.51
r41 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.51
+ $X2=3.06 $Y2=1.675
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.51
+ $X2=3.06 $Y2=1.345
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=1.51 $X2=3.06 $Y2=1.51
r44 9 13 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=3.11 $Y=1.665
+ $X2=3.11 $Y2=1.51
r45 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.15 $Y=0.665
+ $X2=3.15 $Y2=1.345
r46 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.08 $Y=2.465
+ $X2=3.08 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_4%B 3 7 9 12 13
c32 12 0 1.98204e-19 $X=3.6 $Y=1.51
r33 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=1.51 $X2=3.6
+ $Y2=1.675
r34 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=1.51 $X2=3.6
+ $Y2=1.345
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.6
+ $Y=1.51 $X2=3.6 $Y2=1.51
r36 9 13 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.56 $Y=1.665
+ $X2=3.56 $Y2=1.51
r37 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.51 $Y=2.465
+ $X2=3.51 $Y2=1.675
r38 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.51 $Y=0.665
+ $X2=3.51 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_4%A_49_133# 1 2 9 11 13 17 21 22 23 26 27 34
c76 26 0 1.98204e-19 $X=3.95 $Y=2.43
r77 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.175
+ $Y=1.51 $X2=4.175 $Y2=1.51
r78 31 34 8.36451 $w=3.08e-07 $l=2.25e-07 $layer=LI1_cond $X=3.95 $Y=1.49
+ $X2=4.175 $Y2=1.49
r79 27 29 7.00478 $w=1.88e-07 $l=1.2e-07 $layer=LI1_cond $X=2.36 $Y=2.4 $X2=2.36
+ $Y2=2.52
r80 25 31 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.95 $Y=1.645
+ $X2=3.95 $Y2=1.49
r81 25 26 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.95 $Y=1.645
+ $X2=3.95 $Y2=2.43
r82 24 29 1.04402 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.455 $Y=2.52
+ $X2=2.36 $Y2=2.52
r83 23 26 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.865 $Y=2.52
+ $X2=3.95 $Y2=2.43
r84 23 24 86.8788 $w=1.78e-07 $l=1.41e-06 $layer=LI1_cond $X=3.865 $Y=2.52
+ $X2=2.455 $Y2=2.52
r85 21 27 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.265 $Y=2.4 $X2=2.36
+ $Y2=2.4
r86 21 22 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=2.265 $Y=2.4
+ $X2=0.455 $Y2=2.4
r87 17 20 53.9343 $w=2.48e-07 $l=1.17e-06 $layer=LI1_cond $X=0.33 $Y=0.875
+ $X2=0.33 $Y2=2.045
r88 15 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.33 $Y=2.315
+ $X2=0.455 $Y2=2.4
r89 15 20 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=0.33 $Y=2.315
+ $X2=0.33 $Y2=2.045
r90 11 35 38.7288 $w=3.45e-07 $l=1.9775e-07 $layer=POLY_cond $X=4.085 $Y=1.675
+ $X2=4.157 $Y2=1.51
r91 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.085 $Y=1.675
+ $X2=4.085 $Y2=2.465
r92 7 35 38.7288 $w=3.45e-07 $l=2.11849e-07 $layer=POLY_cond $X=4.05 $Y=1.345
+ $X2=4.157 $Y2=1.51
r93 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.05 $Y=1.345 $X2=4.05
+ $Y2=0.665
r94 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.045
r95 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.665 $X2=0.37 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_4%VPWR 1 2 3 4 15 19 21 25 27 31 34 35 36 37
+ 38 49 50 53 56
r70 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r71 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r72 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r73 50 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r74 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 47 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=3.33
+ $X2=3.725 $Y2=3.33
r76 47 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.89 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r78 42 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 38 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 38 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r82 36 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.93 $Y2=3.33
r84 34 41 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.07 $Y2=3.33
r86 33 45 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.235 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=3.33
+ $X2=1.07 $Y2=3.33
r88 29 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=3.245
+ $X2=3.725 $Y2=3.33
r89 29 31 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.725 $Y=3.245
+ $X2=3.725 $Y2=2.905
r90 28 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=3.33
+ $X2=2.79 $Y2=3.33
r91 27 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=3.33
+ $X2=3.725 $Y2=3.33
r92 27 28 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.56 $Y=3.33
+ $X2=2.955 $Y2=3.33
r93 23 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=3.33
r94 23 25 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=2.905
r95 22 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=1.93 $Y2=3.33
r96 21 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.79 $Y2=3.33
r97 21 22 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.095 $Y2=3.33
r98 17 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r99 17 19 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.795
r100 13 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=3.33
r101 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.795
r102 4 31 600 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.835 $X2=3.725 $Y2=2.905
r103 3 25 600 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.835 $X2=2.79 $Y2=2.905
r104 2 19 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.835 $X2=1.93 $Y2=2.795
r105 1 15 600 $w=1.7e-07 $l=1.13842e-06 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.835 $X2=1.07 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_4%X 1 2 3 4 14 15 16 19 21 25 27 28 29 30 37
+ 46
c52 46 0 1.53355e-19 $X=2.36 $Y=1.98
r53 35 37 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.155 $Y=1.98
+ $X2=1.2 $Y2=1.98
r54 30 46 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.16 $Y=1.98 $X2=2.36
+ $Y2=1.98
r55 29 30 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.98
+ $X2=2.16 $Y2=1.98
r56 29 40 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=1.98 $X2=1.5
+ $Y2=1.98
r57 28 35 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=1.98 $X2=1.155
+ $Y2=1.98
r58 28 40 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.22 $Y=1.98 $X2=1.5
+ $Y2=1.98
r59 28 37 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=1.22 $Y=1.98 $X2=1.2
+ $Y2=1.98
r60 23 25 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=2.36 $Y=1.075
+ $X2=2.36 $Y2=0.42
r61 22 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.48 $Y2=1.16
r62 21 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.265 $Y=1.16
+ $X2=2.36 $Y2=1.075
r63 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.265 $Y=1.16
+ $X2=1.595 $Y2=1.16
r64 17 27 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=1.075
+ $X2=1.48 $Y2=1.16
r65 17 19 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.48 $Y=1.075
+ $X2=1.48 $Y2=0.42
r66 15 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.365 $Y=1.16
+ $X2=1.48 $Y2=1.16
r67 15 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.365 $Y=1.16
+ $X2=1.155 $Y2=1.16
r68 14 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=1.815
+ $X2=1.07 $Y2=1.98
r69 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.07 $Y=1.245
+ $X2=1.155 $Y2=1.16
r70 13 14 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.07 $Y=1.245
+ $X2=1.07 $Y2=1.815
r71 4 46 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.835 $X2=2.36 $Y2=1.98
r72 3 40 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=1.98
r73 2 25 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.22
+ $Y=0.245 $X2=2.36 $Y2=0.42
r74 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.36
+ $Y=0.245 $X2=1.5 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_4%VGND 1 2 3 12 16 20 23 24 26 27 29 30 31 47
+ 48
r62 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r63 45 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r64 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r65 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r66 42 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r67 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 35 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r70 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r71 31 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r72 31 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r73 29 41 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.64
+ $Y2=0
r74 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.86
+ $Y2=0
r75 28 44 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.025 $Y=0 $X2=3.12
+ $Y2=0
r76 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=2.86
+ $Y2=0
r77 26 38 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r78 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.93
+ $Y2=0
r79 25 41 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.64
+ $Y2=0
r80 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=1.93
+ $Y2=0
r81 23 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r82 23 24 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.085
+ $Y2=0
r83 22 38 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.68
+ $Y2=0
r84 22 24 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.085
+ $Y2=0
r85 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0
r86 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0.37
r87 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0
r88 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0.39
r89 10 24 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=0.085
+ $X2=1.085 $Y2=0
r90 10 12 15.9771 $w=2.18e-07 $l=3.05e-07 $layer=LI1_cond $X=1.085 $Y=0.085
+ $X2=1.085 $Y2=0.39
r91 3 20 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=2.65
+ $Y=0.245 $X2=2.86 $Y2=0.37
r92 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.79
+ $Y=0.245 $X2=1.93 $Y2=0.39
r93 1 12 91 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=2 $X=0.68
+ $Y=0.665 $X2=1.07 $Y2=0.39
.ends

