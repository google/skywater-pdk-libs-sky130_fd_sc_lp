* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
X0 VPWR GATE_N a_219_135# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VGND GATE_N a_219_135# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_363_483# a_219_135# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_1069_161# a_806_385# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_1069_161# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_626_47# a_219_135# a_764_483# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_764_483# a_806_385# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_626_47# a_806_385# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_1069_161# a_806_385# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VPWR a_34_407# a_584_483# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_584_483# a_363_483# a_626_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_626_47# a_363_483# a_734_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_1069_161# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_734_47# a_806_385# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND a_806_385# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR a_806_385# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_363_483# a_219_135# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_34_407# a_554_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_626_47# a_806_385# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_34_407# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_34_407# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_554_47# a_219_135# a_626_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
