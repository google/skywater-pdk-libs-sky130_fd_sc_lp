* File: sky130_fd_sc_lp__nor3b_1.pex.spice
* Created: Wed Sep  2 10:09:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3B_1%C_N 1 3 4 6 7 8
c25 4 0 1.10796e-20 $X=0.75 $Y=1.725
r26 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.375 $X2=0.63 $Y2=1.375
r27 8 13 8.68074 $w=3.83e-07 $l=2.9e-07 $layer=LI1_cond $X=0.667 $Y=1.665
+ $X2=0.667 $Y2=1.375
r28 7 13 2.39469 $w=3.83e-07 $l=8e-08 $layer=LI1_cond $X=0.667 $Y=1.295
+ $X2=0.667 $Y2=1.375
r29 4 12 69.9537 $w=2.85e-07 $l=3.99061e-07 $layer=POLY_cond $X=0.75 $Y=1.725
+ $X2=0.645 $Y2=1.375
r30 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.75 $Y=1.725 $X2=0.75
+ $Y2=2.045
r31 1 12 42.8941 $w=2.85e-07 $l=2.36749e-07 $layer=POLY_cond $X=0.75 $Y=1.185
+ $X2=0.645 $Y2=1.375
r32 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.75 $Y=1.185 $X2=0.75
+ $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_1%A 3 7 9 10 14
c35 14 0 2.33147e-20 $X=1.2 $Y=1.375
c36 10 0 2.71618e-19 $X=1.2 $Y=1.665
r37 14 17 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.205 $Y=1.375
+ $X2=1.205 $Y2=1.54
r38 14 16 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.205 $Y=1.375
+ $X2=1.205 $Y2=1.21
r39 9 10 14.6084 $w=3.09e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.665
r40 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.375 $X2=1.2 $Y2=1.375
r41 7 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.3 $Y=2.465 $X2=1.3
+ $Y2=1.54
r42 3 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.3 $Y=0.655 $X2=1.3
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_1%B 3 7 9 12 13
c37 12 0 3.10063e-20 $X=1.75 $Y=1.51
c38 3 0 1.94574e-20 $X=1.66 $Y=2.465
r39 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.51
+ $X2=1.75 $Y2=1.675
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.51
+ $X2=1.75 $Y2=1.345
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.51 $X2=1.75 $Y2=1.51
r42 9 13 5.85668 $w=3.03e-07 $l=1.55e-07 $layer=LI1_cond $X=1.682 $Y=1.665
+ $X2=1.682 $Y2=1.51
r43 7 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.765 $Y=0.655
+ $X2=1.765 $Y2=1.345
r44 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.66 $Y=2.465
+ $X2=1.66 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_1%A_82_131# 1 2 9 13 16 17 18 22 26 31 32
c61 31 0 1.40129e-19 $X=2.29 $Y=1.505
c62 22 0 1.66352e-19 $X=2.09 $Y=1.93
r63 32 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.505
+ $X2=2.29 $Y2=1.67
r64 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.505
+ $X2=2.29 $Y2=1.34
r65 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.505 $X2=2.29 $Y2=1.505
r66 28 31 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.09 $Y=1.505 $X2=2.29
+ $Y2=1.505
r67 23 26 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.195 $Y=0.865
+ $X2=0.535 $Y2=0.865
r68 21 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=1.67
+ $X2=2.09 $Y2=1.505
r69 21 22 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.09 $Y=1.67
+ $X2=2.09 $Y2=1.93
r70 18 20 12.1472 $w=2.08e-07 $l=2.3e-07 $layer=LI1_cond $X=0.305 $Y=2.035
+ $X2=0.535 $Y2=2.035
r71 17 22 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.005 $Y=2.035
+ $X2=2.09 $Y2=1.93
r72 17 20 77.6364 $w=2.08e-07 $l=1.47e-06 $layer=LI1_cond $X=2.005 $Y=2.035
+ $X2=0.535 $Y2=2.035
r73 16 18 6.82129 $w=2.1e-07 $l=1.53786e-07 $layer=LI1_cond $X=0.195 $Y=1.93
+ $X2=0.305 $Y2=2.035
r74 15 23 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.195 $Y=1.03
+ $X2=0.195 $Y2=0.865
r75 15 16 47.1454 $w=2.18e-07 $l=9e-07 $layer=LI1_cond $X=0.195 $Y=1.03
+ $X2=0.195 $Y2=1.93
r76 13 36 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.2 $Y=2.465
+ $X2=2.2 $Y2=1.67
r77 9 35 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.2 $Y=0.655 $X2=2.2
+ $Y2=1.34
r78 2 20 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.41
+ $Y=1.835 $X2=0.535 $Y2=2.035
r79 1 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.41
+ $Y=0.655 $X2=0.535 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_1%VPWR 1 6 8 10 17 18 21
r22 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r23 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r24 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.085 $Y2=3.33
r25 15 17 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=2.64 $Y2=3.33
r26 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r27 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=3.33
+ $X2=1.085 $Y2=3.33
r29 10 12 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.92 $Y=3.33 $X2=0.72
+ $Y2=3.33
r30 8 18 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r32 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=3.245
+ $X2=1.085 $Y2=3.33
r33 4 6 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.085 $Y=3.245
+ $X2=1.085 $Y2=2.415
r34 1 6 300 $w=1.7e-07 $l=6.97997e-07 $layer=licon1_PDIFF $count=2 $X=0.825
+ $Y=1.835 $X2=1.085 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_1%Y 1 2 3 12 14 15 16 17 18 19 20 21 22 34 40
+ 58 62
r43 58 59 6.97512 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=2.005
+ $X2=2.57 $Y2=1.84
r44 47 62 0.797386 $w=4.48e-07 $l=3e-08 $layer=LI1_cond $X=2.57 $Y=2.065
+ $X2=2.57 $Y2=2.035
r45 32 40 1.86887 $w=4.78e-07 $l=7.5e-08 $layer=LI1_cond $X=2.555 $Y=1 $X2=2.555
+ $Y2=0.925
r46 22 54 3.58824 $w=4.48e-07 $l=1.35e-07 $layer=LI1_cond $X=2.57 $Y=2.775
+ $X2=2.57 $Y2=2.91
r47 21 22 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.57 $Y=2.405
+ $X2=2.57 $Y2=2.775
r48 20 62 0.744227 $w=4.48e-07 $l=2.8e-08 $layer=LI1_cond $X=2.57 $Y=2.007
+ $X2=2.57 $Y2=2.035
r49 20 58 0.053159 $w=4.48e-07 $l=2e-09 $layer=LI1_cond $X=2.57 $Y=2.007
+ $X2=2.57 $Y2=2.005
r50 20 21 8.31939 $w=4.48e-07 $l=3.13e-07 $layer=LI1_cond $X=2.57 $Y=2.092
+ $X2=2.57 $Y2=2.405
r51 20 47 0.717647 $w=4.48e-07 $l=2.7e-08 $layer=LI1_cond $X=2.57 $Y=2.092
+ $X2=2.57 $Y2=2.065
r52 19 59 8.40323 $w=2.38e-07 $l=1.75e-07 $layer=LI1_cond $X=2.675 $Y=1.665
+ $X2=2.675 $Y2=1.84
r53 18 19 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.675 $Y=1.295
+ $X2=2.675 $Y2=1.665
r54 18 41 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=2.675 $Y=1.295
+ $X2=2.675 $Y2=1.17
r55 17 32 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=1.085
+ $X2=2.555 $Y2=1
r56 17 41 2.66603 $w=3.6e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.555 $Y=1.085
+ $X2=2.675 $Y2=1.17
r57 17 40 0.124591 $w=4.78e-07 $l=5e-09 $layer=LI1_cond $X=2.555 $Y=0.92
+ $X2=2.555 $Y2=0.925
r58 16 17 9.09518 $w=4.78e-07 $l=3.65e-07 $layer=LI1_cond $X=2.555 $Y=0.555
+ $X2=2.555 $Y2=0.92
r59 16 34 3.36397 $w=4.78e-07 $l=1.35e-07 $layer=LI1_cond $X=2.555 $Y=0.555
+ $X2=2.555 $Y2=0.42
r60 14 17 4.14084 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=2.315 $Y=1.085
+ $X2=2.555 $Y2=1.085
r61 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.315 $Y=1.085
+ $X2=1.645 $Y2=1.085
r62 10 15 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.55 $Y=1
+ $X2=1.645 $Y2=1.085
r63 10 12 33.8565 $w=1.88e-07 $l=5.8e-07 $layer=LI1_cond $X=1.55 $Y=1 $X2=1.55
+ $Y2=0.42
r64 3 58 400 $w=1.7e-07 $l=2.35053e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.835 $X2=2.43 $Y2=2.005
r65 3 54 400 $w=1.7e-07 $l=1.14989e-06 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.835 $X2=2.43 $Y2=2.91
r66 2 34 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.275
+ $Y=0.235 $X2=2.415 $Y2=0.42
r67 1 12 91 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_NDIFF $count=2 $X=1.375
+ $Y=0.235 $X2=1.55 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_1%VGND 1 2 9 15 18 19 21 22 23 33 34
c37 9 0 1.10796e-20 $X=1.085 $Y=0.38
r38 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r40 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r41 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 23 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r43 23 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r44 21 30 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.68
+ $Y2=0
r45 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.98
+ $Y2=0
r46 20 33 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.64
+ $Y2=0
r47 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=1.98
+ $Y2=0
r48 18 26 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.8 $Y=0 $X2=0.72
+ $Y2=0
r49 18 19 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.8 $Y=0 $X2=1.025
+ $Y2=0
r50 17 30 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.68
+ $Y2=0
r51 17 19 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.025
+ $Y2=0
r52 13 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r53 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.36
r54 9 11 13.1569 $w=4.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.025 $Y=0.38
+ $X2=1.025 $Y2=0.875
r55 7 19 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.025 $Y=0.085
+ $X2=1.025 $Y2=0
r56 7 9 7.84096 $w=4.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.025 $Y=0.085
+ $X2=1.025 $Y2=0.38
r57 2 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.36
r58 1 11 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=0.825
+ $Y=0.655 $X2=0.965 $Y2=0.875
r59 1 9 182 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_NDIFF $count=1 $X=0.825
+ $Y=0.655 $X2=1.085 $Y2=0.38
.ends

