* File: sky130_fd_sc_lp__a22oi_0.pxi.spice
* Created: Fri Aug 28 09:54:45 2020
* 
x_PM_SKY130_FD_SC_LP__A22OI_0%B2 N_B2_M1006_g N_B2_M1004_g N_B2_c_54_n
+ N_B2_c_59_n B2 B2 B2 N_B2_c_56_n PM_SKY130_FD_SC_LP__A22OI_0%B2
x_PM_SKY130_FD_SC_LP__A22OI_0%B1 N_B1_M1003_g N_B1_M1005_g N_B1_c_89_n
+ N_B1_c_90_n B1 B1 N_B1_c_92_n PM_SKY130_FD_SC_LP__A22OI_0%B1
x_PM_SKY130_FD_SC_LP__A22OI_0%A1 N_A1_M1007_g N_A1_M1002_g A1 A1 A1 N_A1_c_126_n
+ PM_SKY130_FD_SC_LP__A22OI_0%A1
x_PM_SKY130_FD_SC_LP__A22OI_0%A2 N_A2_c_161_n N_A2_M1001_g N_A2_M1000_g
+ N_A2_c_162_n N_A2_c_163_n N_A2_c_169_n N_A2_c_164_n A2 A2 N_A2_c_166_n
+ PM_SKY130_FD_SC_LP__A22OI_0%A2
x_PM_SKY130_FD_SC_LP__A22OI_0%A_45_405# N_A_45_405#_M1004_s N_A_45_405#_M1005_d
+ N_A_45_405#_M1000_d N_A_45_405#_c_199_n N_A_45_405#_c_200_n
+ N_A_45_405#_c_201_n N_A_45_405#_c_202_n N_A_45_405#_c_203_n
+ N_A_45_405#_c_204_n N_A_45_405#_c_205_n PM_SKY130_FD_SC_LP__A22OI_0%A_45_405#
x_PM_SKY130_FD_SC_LP__A22OI_0%Y N_Y_M1003_d N_Y_M1004_d N_Y_c_243_n N_Y_c_252_n
+ N_Y_c_240_n N_Y_c_241_n Y Y PM_SKY130_FD_SC_LP__A22OI_0%Y
x_PM_SKY130_FD_SC_LP__A22OI_0%VPWR N_VPWR_M1002_d N_VPWR_c_277_n VPWR
+ N_VPWR_c_278_n N_VPWR_c_279_n N_VPWR_c_276_n N_VPWR_c_281_n
+ PM_SKY130_FD_SC_LP__A22OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A22OI_0%VGND N_VGND_M1006_s N_VGND_M1001_d N_VGND_c_298_n
+ N_VGND_c_299_n N_VGND_c_300_n N_VGND_c_301_n VGND N_VGND_c_302_n
+ N_VGND_c_303_n PM_SKY130_FD_SC_LP__A22OI_0%VGND
cc_1 VNB N_B2_M1006_g 0.0254253f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.445
cc_2 VNB N_B2_c_54_n 0.00817002f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.725
cc_3 VNB B2 0.0355661f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_4 VNB N_B2_c_56_n 0.0808125f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.005
cc_5 VNB N_B1_M1003_g 0.0196413f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.84
cc_6 VNB N_B1_M1005_g 0.00954729f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.875
cc_7 VNB N_B1_c_89_n 0.0213485f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.725
cc_8 VNB N_B1_c_90_n 0.0153782f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.875
cc_9 VNB B1 0.0101857f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_10 VNB N_B1_c_92_n 0.0155588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_M1007_g 0.035627f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.84
cc_12 VNB N_A1_M1002_g 0.00999475f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.875
cc_13 VNB A1 0.00576459f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.345
cc_14 VNB N_A1_c_126_n 0.0315331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_161_n 0.0209394f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.51
cc_16 VNB N_A2_c_162_n 0.0147148f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.345
cc_17 VNB N_A2_c_163_n 0.0358094f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_18 VNB N_A2_c_164_n 0.0175467f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.005
cc_19 VNB A2 0.0378618f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.005
cc_20 VNB N_A2_c_166_n 0.0318729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_240_n 0.00702037f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_VPWR_c_276_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.005
cc_23 VNB N_VGND_c_298_n 0.0109711f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.875
cc_24 VNB N_VGND_c_299_n 0.0186631f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.345
cc_25 VNB N_VGND_c_300_n 0.0123757f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.725
cc_26 VNB N_VGND_c_301_n 0.0203983f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_27 VNB N_VGND_c_302_n 0.0407636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_303_n 0.147626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_B2_M1004_g 0.0217905f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.345
cc_30 VPB N_B2_c_54_n 0.00389882f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.725
cc_31 VPB N_B2_c_59_n 0.0170801f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.875
cc_32 VPB B2 0.01499f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_33 VPB N_B1_M1005_g 0.0307266f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.875
cc_34 VPB N_A1_M1002_g 0.0300746f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.875
cc_35 VPB N_A2_M1000_g 0.0232788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A2_c_162_n 0.00457782f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.345
cc_37 VPB N_A2_c_169_n 0.0195286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_45_405#_c_199_n 0.0383046f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.875
cc_39 VPB N_A_45_405#_c_200_n 0.0223771f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_40 VPB N_A_45_405#_c_201_n 0.0107624f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_41 VPB N_A_45_405#_c_202_n 0.00825887f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.005
cc_42 VPB N_A_45_405#_c_203_n 0.0194365f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.005
cc_43 VPB N_A_45_405#_c_204_n 0.00627443f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.005
cc_44 VPB N_A_45_405#_c_205_n 0.0373787f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=0.925
cc_45 VPB N_Y_c_241_n 0.00684097f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_46 VPB Y 0.0041639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_277_n 0.0290777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_278_n 0.040999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_279_n 0.0196102f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.005
cc_50 VPB N_VPWR_c_276_n 0.0692884f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.005
cc_51 VPB N_VPWR_c_281_n 0.00516749f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=0.925
cc_52 N_B2_M1006_g N_B1_M1003_g 0.0432461f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_53 N_B2_c_59_n N_B1_M1005_g 0.0173461f $X=0.55 $Y=1.875 $X2=0 $Y2=0
cc_54 N_B2_c_56_n N_B1_M1005_g 0.00718662f $X=0.28 $Y=1.005 $X2=0 $Y2=0
cc_55 N_B2_c_56_n N_B1_c_89_n 0.0432461f $X=0.28 $Y=1.005 $X2=0 $Y2=0
cc_56 N_B2_M1006_g B1 6.38981e-19 $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_57 N_B2_M1004_g N_A_45_405#_c_199_n 0.00589996f $X=0.6 $Y=2.345 $X2=0 $Y2=0
cc_58 N_B2_c_59_n N_A_45_405#_c_199_n 0.00146537f $X=0.55 $Y=1.875 $X2=0 $Y2=0
cc_59 B2 N_A_45_405#_c_199_n 0.017615f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_60 N_B2_c_56_n N_A_45_405#_c_199_n 0.00247799f $X=0.28 $Y=1.005 $X2=0 $Y2=0
cc_61 N_B2_M1004_g N_A_45_405#_c_200_n 0.00619529f $X=0.6 $Y=2.345 $X2=0 $Y2=0
cc_62 N_B2_M1006_g N_Y_c_243_n 0.00781888f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_63 N_B2_M1006_g N_Y_c_240_n 0.0104441f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_64 N_B2_c_54_n N_Y_c_240_n 0.0033337f $X=0.55 $Y=1.725 $X2=0 $Y2=0
cc_65 B2 N_Y_c_240_n 0.0752834f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_66 N_B2_c_56_n N_Y_c_240_n 0.0160547f $X=0.28 $Y=1.005 $X2=0 $Y2=0
cc_67 N_B2_c_54_n N_Y_c_241_n 0.00156016f $X=0.55 $Y=1.725 $X2=0 $Y2=0
cc_68 N_B2_c_59_n N_Y_c_241_n 0.00920403f $X=0.55 $Y=1.875 $X2=0 $Y2=0
cc_69 N_B2_M1004_g Y 0.0162866f $X=0.6 $Y=2.345 $X2=0 $Y2=0
cc_70 N_B2_c_59_n Y 0.00220168f $X=0.55 $Y=1.875 $X2=0 $Y2=0
cc_71 N_B2_M1006_g N_VGND_c_299_n 0.00576179f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_72 B2 N_VGND_c_299_n 0.0190277f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_73 N_B2_c_56_n N_VGND_c_299_n 0.00171268f $X=0.28 $Y=1.005 $X2=0 $Y2=0
cc_74 N_B2_M1006_g N_VGND_c_302_n 0.00495133f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_75 N_B2_M1006_g N_VGND_c_303_n 0.00941123f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_76 B2 N_VGND_c_303_n 0.00268635f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_77 N_B2_c_56_n N_VGND_c_303_n 0.00204523f $X=0.28 $Y=1.005 $X2=0 $Y2=0
cc_78 N_B1_M1003_g N_A1_M1007_g 0.0128757f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_79 B1 N_A1_M1007_g 0.00504593f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_80 N_B1_c_92_n N_A1_M1007_g 0.0169469f $X=0.98 $Y=0.98 $X2=0 $Y2=0
cc_81 N_B1_M1005_g N_A1_M1002_g 0.0264829f $X=1.03 $Y=2.345 $X2=0 $Y2=0
cc_82 N_B1_M1003_g A1 7.9655e-19 $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_83 B1 A1 0.0575638f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_84 N_B1_c_92_n A1 5.70429e-19 $X=0.98 $Y=0.98 $X2=0 $Y2=0
cc_85 N_B1_c_89_n N_A1_c_126_n 0.0169469f $X=0.98 $Y=1.32 $X2=0 $Y2=0
cc_86 N_B1_M1005_g N_A_45_405#_c_200_n 0.00701919f $X=1.03 $Y=2.345 $X2=0 $Y2=0
cc_87 N_B1_M1005_g N_A_45_405#_c_202_n 0.00332444f $X=1.03 $Y=2.345 $X2=0 $Y2=0
cc_88 N_B1_M1005_g N_A_45_405#_c_204_n 0.00151072f $X=1.03 $Y=2.345 $X2=0 $Y2=0
cc_89 N_B1_c_90_n N_A_45_405#_c_204_n 2.33186e-19 $X=0.98 $Y=1.485 $X2=0 $Y2=0
cc_90 B1 N_A_45_405#_c_204_n 0.0160323f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_91 N_B1_M1003_g N_Y_c_252_n 0.0137141f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_92 B1 N_Y_c_252_n 0.0307363f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_93 N_B1_c_92_n N_Y_c_252_n 0.00101885f $X=0.98 $Y=0.98 $X2=0 $Y2=0
cc_94 N_B1_M1003_g N_Y_c_240_n 0.00809798f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_95 N_B1_M1005_g N_Y_c_240_n 0.0035162f $X=1.03 $Y=2.345 $X2=0 $Y2=0
cc_96 B1 N_Y_c_240_n 0.0524857f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_97 N_B1_M1005_g N_Y_c_241_n 0.00317904f $X=1.03 $Y=2.345 $X2=0 $Y2=0
cc_98 N_B1_c_90_n N_Y_c_241_n 0.00424983f $X=0.98 $Y=1.485 $X2=0 $Y2=0
cc_99 B1 N_Y_c_241_n 0.00411436f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_100 N_B1_M1003_g N_VGND_c_302_n 0.00359964f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_101 N_B1_M1003_g N_VGND_c_303_n 0.00551049f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A1_M1007_g N_A2_c_161_n 0.0520681f $X=1.46 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_103 A1 N_A2_c_161_n 0.0133974f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_104 N_A1_M1002_g N_A2_c_162_n 0.00783362f $X=1.46 $Y=2.345 $X2=0 $Y2=0
cc_105 A1 N_A2_c_163_n 0.00455699f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_106 N_A1_M1002_g N_A2_c_169_n 0.017264f $X=1.46 $Y=2.345 $X2=0 $Y2=0
cc_107 N_A1_M1007_g A2 6.47847e-19 $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_108 A1 A2 0.0589432f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_109 N_A1_c_126_n A2 9.87809e-19 $X=1.55 $Y=1.32 $X2=0 $Y2=0
cc_110 N_A1_M1007_g N_A2_c_166_n 0.00615982f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_111 A1 N_A2_c_166_n 0.00198555f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_112 N_A1_c_126_n N_A2_c_166_n 0.0181238f $X=1.55 $Y=1.32 $X2=0 $Y2=0
cc_113 N_A1_M1002_g N_A_45_405#_c_202_n 0.0036065f $X=1.46 $Y=2.345 $X2=0 $Y2=0
cc_114 N_A1_M1002_g N_A_45_405#_c_203_n 0.0174277f $X=1.46 $Y=2.345 $X2=0 $Y2=0
cc_115 A1 N_A_45_405#_c_203_n 0.0235772f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_116 N_A1_c_126_n N_A_45_405#_c_203_n 0.00125321f $X=1.55 $Y=1.32 $X2=0 $Y2=0
cc_117 N_A1_M1007_g N_Y_c_252_n 0.00395186f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_118 A1 N_Y_c_252_n 0.0167729f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_119 N_A1_M1002_g N_VPWR_c_277_n 0.00121054f $X=1.46 $Y=2.345 $X2=0 $Y2=0
cc_120 N_A1_M1002_g N_VPWR_c_278_n 0.00394852f $X=1.46 $Y=2.345 $X2=0 $Y2=0
cc_121 N_A1_M1002_g N_VPWR_c_276_n 0.00458517f $X=1.46 $Y=2.345 $X2=0 $Y2=0
cc_122 N_A1_M1007_g N_VGND_c_302_n 0.00492889f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_123 A1 N_VGND_c_302_n 0.00933827f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_124 N_A1_M1007_g N_VGND_c_303_n 0.0086545f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_125 A1 N_VGND_c_303_n 0.0106165f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_126 A1 A_307_47# 0.00122477f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_127 N_A2_c_162_n N_A_45_405#_c_203_n 0.00498368f $X=2.03 $Y=1.725 $X2=0 $Y2=0
cc_128 N_A2_c_169_n N_A_45_405#_c_203_n 0.0154955f $X=2.03 $Y=1.8 $X2=0 $Y2=0
cc_129 N_A2_c_164_n N_A_45_405#_c_203_n 0.00128115f $X=2.12 $Y=1.485 $X2=0 $Y2=0
cc_130 A2 N_A_45_405#_c_203_n 0.0268171f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_131 N_A2_M1000_g N_A_45_405#_c_205_n 0.00482091f $X=1.89 $Y=2.345 $X2=0 $Y2=0
cc_132 N_A2_c_169_n N_A_45_405#_c_205_n 0.00494594f $X=2.03 $Y=1.8 $X2=0 $Y2=0
cc_133 N_A2_M1000_g N_VPWR_c_277_n 0.00337384f $X=1.89 $Y=2.345 $X2=0 $Y2=0
cc_134 N_A2_M1000_g N_VPWR_c_279_n 0.00394852f $X=1.89 $Y=2.345 $X2=0 $Y2=0
cc_135 N_A2_M1000_g N_VPWR_c_276_n 0.00458517f $X=1.89 $Y=2.345 $X2=0 $Y2=0
cc_136 A2 N_VGND_c_300_n 5.97714e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_137 N_A2_c_161_n N_VGND_c_301_n 0.00462277f $X=1.82 $Y=0.765 $X2=0 $Y2=0
cc_138 N_A2_c_163_n N_VGND_c_301_n 0.00253595f $X=2.12 $Y=0.915 $X2=0 $Y2=0
cc_139 A2 N_VGND_c_301_n 0.0277706f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_140 N_A2_c_161_n N_VGND_c_302_n 0.0054651f $X=1.82 $Y=0.765 $X2=0 $Y2=0
cc_141 N_A2_c_163_n N_VGND_c_302_n 7.72001e-19 $X=2.12 $Y=0.915 $X2=0 $Y2=0
cc_142 N_A2_c_161_n N_VGND_c_303_n 0.0105349f $X=1.82 $Y=0.765 $X2=0 $Y2=0
cc_143 N_A2_c_163_n N_VGND_c_303_n 0.00104801f $X=2.12 $Y=0.915 $X2=0 $Y2=0
cc_144 A2 N_VGND_c_303_n 0.00232495f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_145 N_A_45_405#_c_204_n N_Y_c_241_n 0.015237f $X=1.37 $Y=1.75 $X2=0 $Y2=0
cc_146 N_A_45_405#_c_199_n Y 0.0519175f $X=0.35 $Y=2.17 $X2=0 $Y2=0
cc_147 N_A_45_405#_c_200_n Y 0.025184f $X=1.115 $Y=2.94 $X2=0 $Y2=0
cc_148 N_A_45_405#_c_202_n Y 0.0168544f $X=1.245 $Y=2.17 $X2=0 $Y2=0
cc_149 N_A_45_405#_c_200_n N_VPWR_c_277_n 0.0148258f $X=1.115 $Y=2.94 $X2=0
+ $Y2=0
cc_150 N_A_45_405#_c_202_n N_VPWR_c_277_n 0.0166806f $X=1.245 $Y=2.17 $X2=0
+ $Y2=0
cc_151 N_A_45_405#_c_203_n N_VPWR_c_277_n 0.0226353f $X=1.98 $Y=1.75 $X2=0 $Y2=0
cc_152 N_A_45_405#_c_205_n N_VPWR_c_277_n 0.00308399f $X=2.105 $Y=2.17 $X2=0
+ $Y2=0
cc_153 N_A_45_405#_c_200_n N_VPWR_c_278_n 0.0462126f $X=1.115 $Y=2.94 $X2=0
+ $Y2=0
cc_154 N_A_45_405#_c_201_n N_VPWR_c_278_n 0.0146885f $X=0.455 $Y=2.94 $X2=0
+ $Y2=0
cc_155 N_A_45_405#_c_205_n N_VPWR_c_279_n 0.00571379f $X=2.105 $Y=2.17 $X2=0
+ $Y2=0
cc_156 N_A_45_405#_c_200_n N_VPWR_c_276_n 0.033709f $X=1.115 $Y=2.94 $X2=0 $Y2=0
cc_157 N_A_45_405#_c_201_n N_VPWR_c_276_n 0.0102333f $X=0.455 $Y=2.94 $X2=0
+ $Y2=0
cc_158 N_A_45_405#_c_205_n N_VPWR_c_276_n 0.00867559f $X=2.105 $Y=2.17 $X2=0
+ $Y2=0
cc_159 N_Y_c_243_n N_VGND_c_299_n 0.0266531f $X=0.715 $Y=0.43 $X2=0 $Y2=0
cc_160 N_Y_c_243_n N_VGND_c_302_n 0.00924872f $X=0.715 $Y=0.43 $X2=0 $Y2=0
cc_161 N_Y_c_252_n N_VGND_c_302_n 0.0325038f $X=1.13 $Y=0.43 $X2=0 $Y2=0
cc_162 N_Y_M1003_d N_VGND_c_303_n 0.00651597f $X=0.965 $Y=0.235 $X2=0 $Y2=0
cc_163 N_Y_c_243_n N_VGND_c_303_n 0.00630147f $X=0.715 $Y=0.43 $X2=0 $Y2=0
cc_164 N_Y_c_252_n N_VGND_c_303_n 0.0212465f $X=1.13 $Y=0.43 $X2=0 $Y2=0
cc_165 N_Y_c_243_n A_121_47# 5.29851e-19 $X=0.715 $Y=0.43 $X2=-0.19 $Y2=-0.245
cc_166 N_Y_c_252_n A_121_47# 0.00214773f $X=1.13 $Y=0.43 $X2=-0.19 $Y2=-0.245
cc_167 N_Y_c_240_n A_121_47# 6.58248e-19 $X=0.745 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_168 N_VGND_c_303_n A_121_47# 0.00169085f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
cc_169 N_VGND_c_303_n A_307_47# 0.00181925f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
