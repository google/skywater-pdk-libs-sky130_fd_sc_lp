# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfstp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfstp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.84000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.460000 2.300000 1.790000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.205000 1.850000 15.725000 2.890000 ;
        RECT 15.395000 0.265000 15.725000 0.725000 ;
        RECT 15.485000 0.725000 15.725000 1.850000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.160000 3.685000 1.830000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.750000 0.855000 2.275000 1.110000 ;
        RECT 0.750000 1.110000 2.835000 1.185000 ;
        RECT 1.565000 0.810000 2.275000 0.855000 ;
        RECT 1.565000 1.185000 2.835000 1.280000 ;
        RECT 2.510000 1.280000 2.835000 1.790000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  8.735000 1.920000  9.025000 1.965000 ;
        RECT  8.735000 1.965000 12.385000 2.105000 ;
        RECT  8.735000 2.105000  9.025000 2.150000 ;
        RECT 12.095000 1.920000 12.385000 1.965000 ;
        RECT 12.095000 2.105000 12.385000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.215000 1.510000 4.645000 1.840000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.840000 0.085000 ;
      RECT  0.000000  3.245000 15.840000 3.415000 ;
      RECT  0.115000  0.265000  0.595000 0.675000 ;
      RECT  0.115000  0.675000  0.445000 1.460000 ;
      RECT  0.115000  1.460000  1.385000 1.790000 ;
      RECT  0.115000  1.790000  0.445000 3.065000 ;
      RECT  0.645000  2.025000  0.975000 3.245000 ;
      RECT  1.055000  0.085000  1.385000 0.675000 ;
      RECT  1.205000  2.010000  1.535000 2.895000 ;
      RECT  1.205000  2.895000  2.415000 3.065000 ;
      RECT  1.735000  1.970000  3.185000 2.140000 ;
      RECT  1.735000  2.140000  2.065000 2.715000 ;
      RECT  2.205000  0.265000  2.625000 0.630000 ;
      RECT  2.245000  2.320000  3.615000 2.490000 ;
      RECT  2.245000  2.490000  2.415000 2.895000 ;
      RECT  2.455000  0.630000  2.625000 0.760000 ;
      RECT  2.455000  0.760000  3.625000 0.930000 ;
      RECT  2.755000  2.670000  3.085000 3.245000 ;
      RECT  3.015000  0.930000  3.185000 1.970000 ;
      RECT  3.025000  0.085000  3.275000 0.580000 ;
      RECT  3.365000  2.010000  3.615000 2.320000 ;
      RECT  3.365000  2.490000  3.615000 3.050000 ;
      RECT  3.455000  0.265000  4.410000 0.435000 ;
      RECT  3.455000  0.435000  3.625000 0.760000 ;
      RECT  3.810000  0.615000  4.060000 0.980000 ;
      RECT  3.845000  2.020000  5.100000 2.190000 ;
      RECT  3.845000  2.190000  4.175000 3.065000 ;
      RECT  3.865000  0.980000  4.035000 2.020000 ;
      RECT  4.240000  0.435000  4.410000 1.160000 ;
      RECT  4.240000  1.160000  5.450000 1.330000 ;
      RECT  4.375000  2.370000  4.705000 3.245000 ;
      RECT  4.630000  0.085000  4.800000 0.980000 ;
      RECT  4.825000  1.555000  5.100000 2.020000 ;
      RECT  4.905000  2.370000  5.235000 2.895000 ;
      RECT  4.905000  2.895000  6.980000 3.065000 ;
      RECT  4.990000  0.265000  6.150000 0.435000 ;
      RECT  4.990000  0.435000  5.160000 1.160000 ;
      RECT  5.280000  1.330000  5.450000 2.020000 ;
      RECT  5.280000  2.020000  5.770000 2.190000 ;
      RECT  5.340000  0.615000  5.800000 0.980000 ;
      RECT  5.440000  2.190000  5.770000 2.715000 ;
      RECT  5.630000  0.980000  5.800000 1.300000 ;
      RECT  5.630000  1.300000  6.895000 1.630000 ;
      RECT  5.630000  1.630000  6.120000 1.840000 ;
      RECT  5.950000  1.840000  6.120000 2.895000 ;
      RECT  5.980000  0.435000  6.150000 1.065000 ;
      RECT  6.300000  2.075000  7.245000 2.245000 ;
      RECT  6.300000  2.245000  6.630000 2.715000 ;
      RECT  6.395000  0.605000  6.725000 0.865000 ;
      RECT  6.395000  0.865000  7.915000 1.035000 ;
      RECT  6.395000  1.035000  7.245000 1.065000 ;
      RECT  6.810000  2.505000 10.020000 2.675000 ;
      RECT  6.810000  2.675000  6.980000 2.895000 ;
      RECT  7.075000  1.065000  7.245000 2.075000 ;
      RECT  7.315000  0.085000  7.565000 0.685000 ;
      RECT  7.425000  1.215000  8.265000 1.385000 ;
      RECT  7.425000  1.385000  7.755000 2.075000 ;
      RECT  7.425000  2.075000  8.590000 2.325000 ;
      RECT  7.440000  2.855000  7.770000 3.245000 ;
      RECT  7.745000  0.265000  8.905000 0.435000 ;
      RECT  7.745000  0.435000  7.915000 0.865000 ;
      RECT  7.995000  1.565000  8.615000 1.895000 ;
      RECT  8.095000  0.615000  8.555000 1.065000 ;
      RECT  8.095000  1.065000  8.265000 1.215000 ;
      RECT  8.445000  1.245000  9.640000 1.415000 ;
      RECT  8.445000  1.415000  8.615000 1.565000 ;
      RECT  8.735000  0.435000  8.905000 1.245000 ;
      RECT  8.790000  2.855000  9.120000 3.245000 ;
      RECT  8.795000  1.605000  9.100000 2.150000 ;
      RECT  9.085000  0.085000  9.415000 1.065000 ;
      RECT  9.310000  1.415000  9.640000 1.915000 ;
      RECT  9.850000  1.300000 10.180000 1.460000 ;
      RECT  9.850000  1.460000 11.055000 1.630000 ;
      RECT  9.850000  1.630000 10.020000 2.505000 ;
      RECT 10.085000  0.310000 10.530000 0.915000 ;
      RECT 10.085000  0.915000 11.405000 1.085000 ;
      RECT 10.240000  2.075000 10.570000 2.330000 ;
      RECT 10.240000  2.330000 12.655000 2.500000 ;
      RECT 10.240000  2.500000 10.570000 3.065000 ;
      RECT 10.750000  1.630000 11.055000 1.935000 ;
      RECT 11.235000  1.085000 11.405000 2.330000 ;
      RECT 11.375000  0.085000 11.705000 0.735000 ;
      RECT 11.545000  2.680000 11.875000 3.245000 ;
      RECT 11.585000  0.915000 13.135000 1.085000 ;
      RECT 11.585000  1.085000 11.890000 1.885000 ;
      RECT 12.100000  1.265000 12.430000 2.150000 ;
      RECT 12.325000  2.500000 12.655000 2.895000 ;
      RECT 12.325000  2.895000 13.485000 3.065000 ;
      RECT 12.465000  0.265000 12.795000 0.915000 ;
      RECT 12.885000  1.085000 13.135000 2.715000 ;
      RECT 13.255000  0.085000 13.585000 0.725000 ;
      RECT 13.315000  0.905000 13.645000 1.575000 ;
      RECT 13.315000  1.575000 13.485000 2.895000 ;
      RECT 13.665000  1.755000 13.915000 3.245000 ;
      RECT 13.815000  0.265000 14.265000 0.725000 ;
      RECT 14.095000  0.725000 14.265000 0.990000 ;
      RECT 14.095000  0.990000 15.240000 1.160000 ;
      RECT 14.095000  1.160000 14.475000 2.890000 ;
      RECT 14.605000  0.085000 14.935000 0.725000 ;
      RECT 14.675000  1.850000 15.005000 3.245000 ;
      RECT 14.910000  1.160000 15.240000 1.660000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.950000  8.965000 2.120000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  1.950000 12.325000 2.120000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfstp_lp
