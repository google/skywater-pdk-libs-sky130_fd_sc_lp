* File: sky130_fd_sc_lp__o21ai_4.pex.spice
* Created: Fri Aug 28 11:04:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21AI_4%A1 1 3 6 8 10 13 15 17 20 24 28 29 31 35 37
+ 38 39 40 54 57 69 71
c111 54 0 4.30413e-20 $X=1.36 $Y=1.35
c112 31 0 7.69757e-20 $X=3.57 $Y=1.16
r113 53 69 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=1.31 $Y=1.362
+ $X2=1.42 $Y2=1.362
r114 52 54 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.31 $Y=1.35 $X2=1.36
+ $Y2=1.35
r115 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.31
+ $Y=1.35 $X2=1.31 $Y2=1.35
r116 50 52 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=0.93 $Y=1.35
+ $X2=1.31 $Y2=1.35
r117 49 50 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.5 $Y=1.35
+ $X2=0.93 $Y2=1.35
r118 46 49 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.29 $Y=1.35
+ $X2=0.5 $Y2=1.35
r119 40 71 8.31148 $w=4.38e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=1.295
+ $X2=1.825 $Y2=1.295
r120 40 69 7.90579 $w=4.38e-07 $l=2.6e-07 $layer=LI1_cond $X=1.68 $Y=1.295
+ $X2=1.42 $Y2=1.295
r121 39 53 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=1.2 $Y=1.362
+ $X2=1.31 $Y2=1.362
r122 38 39 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.362
+ $X2=1.2 $Y2=1.362
r123 37 38 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.362
+ $X2=0.72 $Y2=1.362
r124 37 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=1.35 $X2=0.29 $Y2=1.35
r125 35 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.35
+ $X2=3.53 $Y2=1.515
r126 35 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.35
+ $X2=3.53 $Y2=1.185
r127 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.53
+ $Y=1.35 $X2=3.53 $Y2=1.35
r128 31 34 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=3.57 $Y=1.16
+ $X2=3.57 $Y2=1.35
r129 29 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.445 $Y=1.16
+ $X2=3.57 $Y2=1.16
r130 29 71 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=3.445 $Y=1.16
+ $X2=1.825 $Y2=1.16
r131 28 57 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.55 $Y=0.655
+ $X2=3.55 $Y2=1.185
r132 24 58 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.51 $Y=2.465
+ $X2=3.51 $Y2=1.515
r133 18 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.515
+ $X2=1.36 $Y2=1.35
r134 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.36 $Y=1.515
+ $X2=1.36 $Y2=2.465
r135 15 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.36 $Y2=1.35
r136 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.36 $Y2=0.655
r137 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.515
+ $X2=0.93 $Y2=1.35
r138 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.93 $Y=1.515
+ $X2=0.93 $Y2=2.465
r139 8 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=1.35
r140 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=0.655
r141 4 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.515
+ $X2=0.5 $Y2=1.35
r142 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.5 $Y=1.515 $X2=0.5
+ $Y2=2.465
r143 1 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.185
+ $X2=0.5 $Y2=1.35
r144 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.5 $Y=1.185 $X2=0.5
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_4%A2 3 7 11 15 19 23 27 31 33 34 35 52
c86 52 0 7.69757e-20 $X=3.08 $Y=1.51
c87 35 0 4.30413e-20 $X=3.12 $Y=1.665
r88 50 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.99 $Y=1.51 $X2=3.08
+ $Y2=1.51
r89 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.51 $X2=2.99 $Y2=1.51
r90 48 50 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.65 $Y=1.51
+ $X2=2.99 $Y2=1.51
r91 46 48 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.59 $Y=1.51 $X2=2.65
+ $Y2=1.51
r92 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.51 $X2=2.59 $Y2=1.51
r93 44 46 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=2.22 $Y=1.51
+ $X2=2.59 $Y2=1.51
r94 42 44 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.16 $Y=1.51 $X2=2.22
+ $Y2=1.51
r95 39 42 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=1.79 $Y=1.51
+ $X2=2.16 $Y2=1.51
r96 35 51 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.592
+ $X2=2.99 $Y2=1.592
r97 34 51 12.0404 $w=3.33e-07 $l=3.5e-07 $layer=LI1_cond $X=2.64 $Y=1.592
+ $X2=2.99 $Y2=1.592
r98 34 47 1.72006 $w=3.33e-07 $l=5e-08 $layer=LI1_cond $X=2.64 $Y=1.592 $X2=2.59
+ $Y2=1.592
r99 33 47 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=2.59 $Y2=1.592
r100 33 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.51 $X2=2.16 $Y2=1.51
r101 29 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=1.675
+ $X2=3.08 $Y2=1.51
r102 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.08 $Y=1.675
+ $X2=3.08 $Y2=2.465
r103 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=1.345
+ $X2=3.08 $Y2=1.51
r104 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.08 $Y=1.345
+ $X2=3.08 $Y2=0.655
r105 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.675
+ $X2=2.65 $Y2=1.51
r106 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.65 $Y=1.675
+ $X2=2.65 $Y2=2.465
r107 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.345
+ $X2=2.65 $Y2=1.51
r108 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.65 $Y=1.345
+ $X2=2.65 $Y2=0.655
r109 13 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.675
+ $X2=2.22 $Y2=1.51
r110 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.22 $Y=1.675
+ $X2=2.22 $Y2=2.465
r111 9 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.345
+ $X2=2.22 $Y2=1.51
r112 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.22 $Y=1.345
+ $X2=2.22 $Y2=0.655
r113 5 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.675
+ $X2=1.79 $Y2=1.51
r114 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.79 $Y=1.675
+ $X2=1.79 $Y2=2.465
r115 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.345
+ $X2=1.79 $Y2=1.51
r116 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.79 $Y=1.345
+ $X2=1.79 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 45
r69 43 45 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.09 $Y=1.35 $X2=5.27
+ $Y2=1.35
r70 41 43 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=4.84 $Y=1.35
+ $X2=5.09 $Y2=1.35
r71 40 41 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.41 $Y=1.35
+ $X2=4.84 $Y2=1.35
r72 38 40 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.07 $Y=1.35
+ $X2=4.41 $Y2=1.35
r73 35 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.98 $Y=1.35 $X2=4.07
+ $Y2=1.35
r74 31 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.09
+ $Y=1.35 $X2=5.09 $Y2=1.35
r75 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.322
+ $X2=5.04 $Y2=1.322
r76 29 30 25.0976 $w=2.23e-07 $l=4.9e-07 $layer=LI1_cond $X=4.07 $Y=1.322
+ $X2=4.56 $Y2=1.322
r77 29 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.07
+ $Y=1.35 $X2=4.07 $Y2=1.35
r78 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.27 $Y=1.515
+ $X2=5.27 $Y2=1.35
r79 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.27 $Y=1.515
+ $X2=5.27 $Y2=2.465
r80 22 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.27 $Y=1.185
+ $X2=5.27 $Y2=1.35
r81 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.27 $Y=1.185
+ $X2=5.27 $Y2=0.655
r82 18 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.84 $Y=1.515
+ $X2=4.84 $Y2=1.35
r83 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.84 $Y=1.515
+ $X2=4.84 $Y2=2.465
r84 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.84 $Y=1.185
+ $X2=4.84 $Y2=1.35
r85 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.84 $Y=1.185
+ $X2=4.84 $Y2=0.655
r86 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=1.515
+ $X2=4.41 $Y2=1.35
r87 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.41 $Y=1.515
+ $X2=4.41 $Y2=2.465
r88 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=1.185
+ $X2=4.41 $Y2=1.35
r89 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.41 $Y=1.185
+ $X2=4.41 $Y2=0.655
r90 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=1.515
+ $X2=3.98 $Y2=1.35
r91 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.98 $Y=1.515 $X2=3.98
+ $Y2=2.465
r92 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=1.185
+ $X2=3.98 $Y2=1.35
r93 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.98 $Y=1.185 $X2=3.98
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_4%VPWR 1 2 3 4 5 16 18 24 30 34 38 40 44 46 51
+ 56 61 70 73 76 80
r88 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r89 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r91 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r92 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r93 65 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r94 65 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r95 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r96 62 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.79 $Y=3.33
+ $X2=4.625 $Y2=3.33
r97 62 64 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.79 $Y=3.33
+ $X2=5.04 $Y2=3.33
r98 61 79 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=5.32 $Y=3.33 $X2=5.54
+ $Y2=3.33
r99 61 64 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.32 $Y=3.33
+ $X2=5.04 $Y2=3.33
r100 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r101 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r102 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r103 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=3.33
+ $X2=3.745 $Y2=3.33
r104 57 59 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.91 $Y=3.33
+ $X2=4.08 $Y2=3.33
r105 56 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.625 $Y2=3.33
r106 56 59 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 55 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r108 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 52 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=3.33
+ $X2=1.145 $Y2=3.33
r110 52 54 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.31 $Y=3.33
+ $X2=1.68 $Y2=3.33
r111 51 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=3.33
+ $X2=3.745 $Y2=3.33
r112 51 54 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=3.58 $Y=3.33
+ $X2=1.68 $Y2=3.33
r113 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r114 50 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r115 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 47 67 4.31589 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.202 $Y2=3.33
r117 47 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 46 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.145 $Y2=3.33
r119 46 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 44 74 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r121 44 55 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.68 $Y2=3.33
r122 40 43 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.485 $Y=2.19
+ $X2=5.485 $Y2=2.95
r123 38 79 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=5.485 $Y=3.245
+ $X2=5.54 $Y2=3.33
r124 38 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.485 $Y=3.245
+ $X2=5.485 $Y2=2.95
r125 34 37 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=4.625 $Y=2.19
+ $X2=4.625 $Y2=2.95
r126 32 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=3.33
r127 32 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=2.95
r128 28 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.745 $Y=3.245
+ $X2=3.745 $Y2=3.33
r129 28 30 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=3.745 $Y=3.245
+ $X2=3.745 $Y2=2.4
r130 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.145 $Y=2.18
+ $X2=1.145 $Y2=2.95
r131 22 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=3.33
r132 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=2.95
r133 18 21 39.2235 $w=2.83e-07 $l=9.7e-07 $layer=LI1_cond $X=0.262 $Y=1.98
+ $X2=0.262 $Y2=2.95
r134 16 67 3.08278 $w=2.85e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.262 $Y=3.245
+ $X2=0.202 $Y2=3.33
r135 16 21 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.262 $Y=3.245
+ $X2=0.262 $Y2=2.95
r136 5 43 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.345
+ $Y=1.835 $X2=5.485 $Y2=2.95
r137 5 40 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=5.345
+ $Y=1.835 $X2=5.485 $Y2=2.19
r138 4 37 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.835 $X2=4.625 $Y2=2.95
r139 4 34 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.835 $X2=4.625 $Y2=2.19
r140 3 30 300 $w=1.7e-07 $l=6.4002e-07 $layer=licon1_PDIFF $count=2 $X=3.585
+ $Y=1.835 $X2=3.745 $Y2=2.4
r141 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.835 $X2=1.145 $Y2=2.95
r142 2 24 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.835 $X2=1.145 $Y2=2.18
r143 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=2.95
r144 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_4%A_115_367# 1 2 3 4 15 19 20 22 25 29 31 35
+ 39
r40 33 35 24.8225 $w=2.08e-07 $l=4.7e-07 $layer=LI1_cond $X=3.305 $Y=2.905
+ $X2=3.305 $Y2=2.435
r41 32 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.53 $Y=2.99
+ $X2=2.435 $Y2=2.99
r42 31 33 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.2 $Y=2.99
+ $X2=3.305 $Y2=2.905
r43 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.2 $Y=2.99 $X2=2.53
+ $Y2=2.99
r44 27 39 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=2.905
+ $X2=2.435 $Y2=2.99
r45 27 29 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=2.435 $Y=2.905
+ $X2=2.435 $Y2=2.435
r46 26 38 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.67 $Y=2.99
+ $X2=1.575 $Y2=2.99
r47 25 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.34 $Y=2.99
+ $X2=2.435 $Y2=2.99
r48 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.34 $Y=2.99
+ $X2=1.67 $Y2=2.99
r49 22 38 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=2.905
+ $X2=1.575 $Y2=2.99
r50 22 24 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=1.575 $Y=2.905
+ $X2=1.575 $Y2=1.98
r51 21 24 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.575 $Y=1.925
+ $X2=1.575 $Y2=1.98
r52 19 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.48 $Y=1.84
+ $X2=1.575 $Y2=1.925
r53 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.48 $Y=1.84
+ $X2=0.81 $Y2=1.84
r54 15 17 45.6073 $w=2.33e-07 $l=9.3e-07 $layer=LI1_cond $X=0.692 $Y=1.98
+ $X2=0.692 $Y2=2.91
r55 13 20 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.692 $Y=1.925
+ $X2=0.81 $Y2=1.84
r56 13 15 2.69721 $w=2.33e-07 $l=5.5e-08 $layer=LI1_cond $X=0.692 $Y=1.925
+ $X2=0.692 $Y2=1.98
r57 4 35 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=3.155
+ $Y=1.835 $X2=3.295 $Y2=2.435
r58 3 29 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=2.295
+ $Y=1.835 $X2=2.435 $Y2=2.435
r59 2 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.835 $X2=1.575 $Y2=2.91
r60 2 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.835 $X2=1.575 $Y2=1.98
r61 1 17 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.715 $Y2=2.91
r62 1 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.715 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_4%Y 1 2 3 4 5 6 21 25 29 31 37 38 41 46 48 53
+ 57
r79 56 57 12.4652 $w=2.43e-07 $l=2.65e-07 $layer=LI1_cond $X=5.547 $Y=1.03
+ $X2=5.547 $Y2=1.295
r80 54 57 14.5819 $w=2.43e-07 $l=3.1e-07 $layer=LI1_cond $X=5.547 $Y=1.605
+ $X2=5.547 $Y2=1.295
r81 53 54 2.32264 $w=2.45e-07 $l=1.6e-07 $layer=LI1_cond $X=5.547 $Y=1.765
+ $X2=5.547 $Y2=1.605
r82 52 53 17.7188 $w=3.18e-07 $l=4.92e-07 $layer=LI1_cond $X=5.055 $Y=1.765
+ $X2=5.547 $Y2=1.765
r83 49 51 0.290476 $w=4.2e-07 $l=1e-08 $layer=LI1_cond $X=4.185 $Y=1.852
+ $X2=4.195 $Y2=1.852
r84 41 43 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=5.055 $Y=1.98
+ $X2=5.055 $Y2=2.91
r85 39 52 3.78705 $w=1.9e-07 $l=1.6e-07 $layer=LI1_cond $X=5.055 $Y=1.925
+ $X2=5.055 $Y2=1.765
r86 39 41 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=5.055 $Y=1.925
+ $X2=5.055 $Y2=1.98
r87 38 51 3.48098 $w=4.2e-07 $l=1.31491e-07 $layer=LI1_cond $X=4.29 $Y=1.765
+ $X2=4.195 $Y2=1.852
r88 37 52 3.42132 $w=3.18e-07 $l=9.5e-08 $layer=LI1_cond $X=4.96 $Y=1.765
+ $X2=5.055 $Y2=1.765
r89 37 38 24.1293 $w=3.18e-07 $l=6.7e-07 $layer=LI1_cond $X=4.96 $Y=1.765
+ $X2=4.29 $Y2=1.765
r90 33 36 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.195 $Y=0.865
+ $X2=5.055 $Y2=0.865
r91 31 56 7.01204 $w=3.3e-07 $l=2.17612e-07 $layer=LI1_cond $X=5.425 $Y=0.865
+ $X2=5.547 $Y2=1.03
r92 31 36 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.425 $Y=0.865
+ $X2=5.055 $Y2=0.865
r93 27 49 4.80115 $w=2.1e-07 $l=2.48e-07 $layer=LI1_cond $X=4.185 $Y=2.1
+ $X2=4.185 $Y2=1.852
r94 27 29 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=4.185 $Y=2.1
+ $X2=4.185 $Y2=2.435
r95 26 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=2.015
+ $X2=2.865 $Y2=2.015
r96 25 49 25.9511 $w=4.2e-07 $l=8.17447e-07 $layer=LI1_cond $X=3.445 $Y=2.015
+ $X2=4.185 $Y2=1.852
r97 25 26 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.445 $Y=2.015
+ $X2=3.03 $Y2=2.015
r98 22 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=2.015
+ $X2=2.005 $Y2=2.015
r99 21 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=2.015
+ $X2=2.865 $Y2=2.015
r100 21 22 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.7 $Y=2.015
+ $X2=2.17 $Y2=2.015
r101 6 43 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.915
+ $Y=1.835 $X2=5.055 $Y2=2.91
r102 6 41 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.915
+ $Y=1.835 $X2=5.055 $Y2=1.98
r103 5 51 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.835 $X2=4.195 $Y2=1.98
r104 5 29 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=4.055
+ $Y=1.835 $X2=4.195 $Y2=2.435
r105 4 48 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=2.725
+ $Y=1.835 $X2=2.865 $Y2=2.085
r106 3 46 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=1.865
+ $Y=1.835 $X2=2.005 $Y2=2.085
r107 2 36 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=4.915
+ $Y=0.235 $X2=5.055 $Y2=0.865
r108 1 33 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=4.055
+ $Y=0.235 $X2=4.195 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_4%A_32_47# 1 2 3 4 5 6 7 24 26 27 30 32 36 38
+ 42 44 46 47 52 54 59 61
r79 54 56 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=1.15 $Y=0.82
+ $X2=1.15 $Y2=0.955
r80 54 55 4.75232 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.82
+ $X2=1.15 $Y2=0.735
r81 50 52 36.04 $w=2.73e-07 $l=8.6e-07 $layer=LI1_cond $X=4.625 $Y=0.392
+ $X2=5.485 $Y2=0.392
r82 48 63 3.55899 $w=2.75e-07 $l=1.5e-07 $layer=LI1_cond $X=3.93 $Y=0.392
+ $X2=3.78 $Y2=0.392
r83 48 50 29.1254 $w=2.73e-07 $l=6.95e-07 $layer=LI1_cond $X=3.93 $Y=0.392
+ $X2=4.625 $Y2=0.392
r84 47 65 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=0.735 $X2=3.78
+ $Y2=0.82
r85 46 63 3.27427 $w=3e-07 $l=1.38e-07 $layer=LI1_cond $X=3.78 $Y=0.53 $X2=3.78
+ $Y2=0.392
r86 46 47 7.87503 $w=2.98e-07 $l=2.05e-07 $layer=LI1_cond $X=3.78 $Y=0.53
+ $X2=3.78 $Y2=0.735
r87 45 61 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.96 $Y=0.82
+ $X2=2.865 $Y2=0.82
r88 44 65 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.63 $Y=0.82 $X2=3.78
+ $Y2=0.82
r89 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.63 $Y=0.82
+ $X2=2.96 $Y2=0.82
r90 40 61 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0.735
+ $X2=2.865 $Y2=0.82
r91 40 42 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=2.865 $Y=0.735
+ $X2=2.865 $Y2=0.42
r92 39 59 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.1 $Y=0.82 $X2=2.005
+ $Y2=0.82
r93 38 61 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.77 $Y=0.82
+ $X2=2.865 $Y2=0.82
r94 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.77 $Y=0.82 $X2=2.1
+ $Y2=0.82
r95 34 59 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=0.735
+ $X2=2.005 $Y2=0.82
r96 34 36 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=2.005 $Y=0.735
+ $X2=2.005 $Y2=0.42
r97 33 54 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.25 $Y=0.82 $X2=1.15
+ $Y2=0.82
r98 32 59 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.91 $Y=0.82
+ $X2=2.005 $Y2=0.82
r99 32 33 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.91 $Y=0.82
+ $X2=1.25 $Y2=0.82
r100 30 55 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.145 $Y=0.43
+ $X2=1.145 $Y2=0.735
r101 26 56 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.05 $Y=0.955 $X2=1.15
+ $Y2=0.955
r102 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.05 $Y=0.955
+ $X2=0.38 $Y2=0.955
r103 22 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.25 $Y=0.87
+ $X2=0.38 $Y2=0.955
r104 22 24 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=0.25 $Y=0.87
+ $X2=0.25 $Y2=0.42
r105 7 52 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.235 $X2=5.485 $Y2=0.435
r106 6 50 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.485
+ $Y=0.235 $X2=4.625 $Y2=0.415
r107 5 65 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=3.625
+ $Y=0.235 $X2=3.765 $Y2=0.82
r108 5 63 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.625
+ $Y=0.235 $X2=3.765 $Y2=0.42
r109 4 61 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=2.725
+ $Y=0.235 $X2=2.865 $Y2=0.82
r110 4 42 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.725
+ $Y=0.235 $X2=2.865 $Y2=0.42
r111 3 59 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.235 $X2=2.005 $Y2=0.82
r112 3 36 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.235 $X2=2.005 $Y2=0.42
r113 2 30 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.235 $X2=1.145 $Y2=0.43
r114 1 24 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 40 59 60 63
r94 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r95 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r96 57 60 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=5.52
+ $Y2=0
r97 56 59 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.52
+ $Y2=0
r98 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r99 54 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r100 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r101 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r102 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r103 48 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r104 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r105 45 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.715
+ $Y2=0
r106 45 47 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.2
+ $Y2=0
r107 43 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r108 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r109 40 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.715
+ $Y2=0
r110 40 42 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r111 38 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r112 38 51 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r113 36 53 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.13 $Y=0 $X2=3.12
+ $Y2=0
r114 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=3.295
+ $Y2=0
r115 35 56 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.46 $Y=0 $X2=3.6
+ $Y2=0
r116 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=0 $X2=3.295
+ $Y2=0
r117 33 50 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.16
+ $Y2=0
r118 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.435
+ $Y2=0
r119 32 53 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.6 $Y=0 $X2=3.12
+ $Y2=0
r120 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=0 $X2=2.435
+ $Y2=0
r121 30 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.2
+ $Y2=0
r122 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.575
+ $Y2=0
r123 29 50 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=2.16
+ $Y2=0
r124 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.575
+ $Y2=0
r125 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=0.085
+ $X2=3.295 $Y2=0
r126 25 27 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.295 $Y=0.085
+ $X2=3.295 $Y2=0.44
r127 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0.085
+ $X2=2.435 $Y2=0
r128 21 23 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.435 $Y=0.085
+ $X2=2.435 $Y2=0.44
r129 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0
r130 17 19 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0.44
r131 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r132 13 15 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.555
r133 4 27 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.235 $X2=3.295 $Y2=0.44
r134 3 23 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.235 $X2=2.435 $Y2=0.44
r135 2 19 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.235 $X2=1.575 $Y2=0.44
r136 1 15 182 $w=1.7e-07 $l=3.83667e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.555
.ends

