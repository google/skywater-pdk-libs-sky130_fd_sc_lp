* File: sky130_fd_sc_lp__o32a_4.spice
* Created: Fri Aug 28 11:17:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32a_4.pex.spice"
.subckt sky130_fd_sc_lp__o32a_4  VNB VPB A2 A1 A3 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A3	A3
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A2_M1012_g N_A_44_65#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.2226 PD=1.46 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75005
+ A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1012_d N_A1_M1006_g N_A_44_65#_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=48.564 NRS=0 M=1 R=5.6 SA=75001
+ SB=75004.3 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1019_d N_A1_M1019_g N_A_44_65#_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75003.8 A=0.126 P=1.98 MULT=1
MM1018 N_VGND_M1019_d N_A2_M1018_g N_A_44_65#_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=4.284 M=1 R=5.6 SA=75001.8
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1017_d N_A3_M1017_g N_A_44_65#_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.1344 PD=1.14 PS=1.16 NRD=2.856 NRS=1.428 M=1 R=5.6 SA=75002.3
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1017_d N_A3_M1022_g N_A_44_65#_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.3003 PD=1.14 PS=1.555 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.7
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1003 N_A_44_65#_M1022_s N_B2_M1003_g N_A_547_367#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.3003 AS=0.147 PD=1.555 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1008 N_A_547_367#_M1003_s N_B1_M1008_g N_A_44_65#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75004.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1021 N_A_547_367#_M1021_d N_B1_M1021_g N_A_44_65#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1197 AS=0.1176 PD=1.125 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.5
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1023 N_A_44_65#_M1023_d N_B2_M1023_g N_A_547_367#_M1021_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2856 AS=0.1197 PD=2.36 PS=1.125 NRD=10.704 NRS=0.708 M=1 R=5.6
+ SA=75005 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1000 N_X_M1000_d N_A_547_367#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1000_d N_A_547_367#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1009 N_X_M1009_d N_A_547_367#_M1009_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1020 N_X_M1009_d N_A_547_367#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_A_195_367#_M1013_d N_A2_M1013_g N_A_112_367#_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_195_367#_M1013_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002 A=0.189 P=2.82 MULT=1
MM1024 N_VPWR_M1002_d N_A1_M1024_g N_A_195_367#_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=6.2449 M=1 R=8.4
+ SA=75001.1 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1015 N_A_195_367#_M1024_s N_A2_M1015_g N_A_112_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_A_547_367#_M1005_d N_A3_M1005_g N_A_112_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_A_547_367#_M1005_d N_A3_M1025_g N_A_112_367#_M1025_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1014 N_A_547_367#_M1014_d N_B2_M1014_g N_A_823_367#_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.17955 PD=3.05 PS=1.545 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1001 N_A_823_367#_M1014_s N_B1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.17955 AS=0.1764 PD=1.545 PS=1.54 NRD=0.7683 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1010 N_A_823_367#_M1010_d N_B1_M1010_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1026 N_A_547_367#_M1026_d N_B2_M1026_g N_A_823_367#_M1010_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A_547_367#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_547_367#_M1011_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1011_d N_A_547_367#_M1016_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_VPWR_M1027_d N_A_547_367#_M1027_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.9271 P=20.81
*
.include "sky130_fd_sc_lp__o32a_4.pxi.spice"
*
.ends
*
*
