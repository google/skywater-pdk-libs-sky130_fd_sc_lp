* File: sky130_fd_sc_lp__or4b_1.spice
* Created: Fri Aug 28 11:25:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4b_1.pex.spice"
.subckt sky130_fd_sc_lp__or4b_1  VNB VPB D_N C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_D_N_M1006_g N_A_64_131#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1002 N_A_220_367#_M1002_d N_A_64_131#_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.7
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_C_M1010_g N_A_220_367#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0588 PD=0.98 PS=0.7 NRD=4.284 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 N_A_220_367#_M1011_d N_B_M1011_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1176 PD=0.7 PS=0.98 NRD=0 NRS=75.708 M=1 R=2.8 SA=75001.8
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_220_367#_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.098 AS=0.0588 PD=0.85 PS=0.7 NRD=27.132 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_X_M1008_d N_A_220_367#_M1008_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.196 PD=2.21 PS=1.7 NRD=0 NRS=4.284 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_D_N_M1005_g N_A_64_131#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_303_367# N_A_64_131#_M1009_g N_A_220_367#_M1009_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=49.25 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1007 A_397_367# N_C_M1007_g A_303_367# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0672 PD=0.7 PS=0.74 NRD=39.8531 NRS=49.25 M=1 R=2.8 SA=75000.7 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1003 A_483_367# N_B_M1003_g A_397_367# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=39.8531 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_483_367# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0441 PD=0.8175 PS=0.63 NRD=44.5417 NRS=23.443 M=1 R=2.8
+ SA=75001.4 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_220_367#_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__or4b_1.pxi.spice"
*
.ends
*
*
