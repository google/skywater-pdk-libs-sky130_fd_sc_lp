* File: sky130_fd_sc_lp__o21ai_1.pex.spice
* Created: Wed Sep  2 10:15:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21AI_1%A1 3 7 9 10 17
r26 14 17 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.295 $Y=1.375
+ $X2=0.485 $Y2=1.375
r27 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.665
r28 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.295
+ $Y=1.375 $X2=0.295 $Y2=1.375
r29 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.54
+ $X2=0.485 $Y2=1.375
r30 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.485 $Y=1.54
+ $X2=0.485 $Y2=2.465
r31 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.21
+ $X2=0.485 $Y2=1.375
r32 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.485 $Y=1.21
+ $X2=0.485 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_1%A2 3 7 9 12 13
r33 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.51
+ $X2=0.935 $Y2=1.675
r34 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.51
+ $X2=0.935 $Y2=1.345
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.935
+ $Y=1.51 $X2=0.935 $Y2=1.51
r36 9 13 6.11791 $w=4.03e-07 $l=2.15e-07 $layer=LI1_cond $X=0.72 $Y=1.547
+ $X2=0.935 $Y2=1.547
r37 7 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.015 $Y=0.655
+ $X2=1.015 $Y2=1.345
r38 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.845 $Y=2.465
+ $X2=0.845 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_1%B1 3 7 9 14 15
r23 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.48 $X2=1.65 $Y2=1.48
r24 11 14 33.7982 $w=3.5e-07 $l=2.05e-07 $layer=POLY_cond $X=1.445 $Y=1.47
+ $X2=1.65 $Y2=1.47
r25 9 15 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=1.682 $Y=1.665
+ $X2=1.682 $Y2=1.48
r26 5 11 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.445 $Y=1.645
+ $X2=1.445 $Y2=1.47
r27 5 7 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.445 $Y=1.645
+ $X2=1.445 $Y2=2.465
r28 1 11 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.445 $Y=1.295
+ $X2=1.445 $Y2=1.47
r29 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.445 $Y=1.295
+ $X2=1.445 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_1%VPWR 1 2 7 9 13 15 19 21 31
r24 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r25 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r26 25 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r28 22 27 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r29 22 24 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=1.2 $Y2=3.33
r30 21 30 4.44548 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.53 $Y=3.33
+ $X2=1.725 $Y2=3.33
r31 21 24 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.53 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 19 25 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 19 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 15 18 33.792 $w=2.93e-07 $l=8.65e-07 $layer=LI1_cond $X=1.677 $Y=2.085
+ $X2=1.677 $Y2=2.95
r35 13 30 3.03205 $w=2.95e-07 $l=1.06325e-07 $layer=LI1_cond $X=1.677 $Y=3.245
+ $X2=1.725 $Y2=3.33
r36 13 18 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=1.677 $Y=3.245
+ $X2=1.677 $Y2=2.95
r37 9 12 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.27 $Y=2.005
+ $X2=0.27 $Y2=2.95
r38 7 27 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r39 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.95
r40 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.835 $X2=1.66 $Y2=2.95
r41 2 15 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.835 $X2=1.66 $Y2=2.085
r42 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.95
r43 1 9 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_1%Y 1 2 9 10 13 15 16 17 30
r26 17 27 4.80185 $w=4.18e-07 $l=1.75e-07 $layer=LI1_cond $X=1.15 $Y=2.775
+ $X2=1.15 $Y2=2.95
r27 16 17 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=2.405
+ $X2=1.15 $Y2=2.775
r28 16 21 7.54576 $w=4.18e-07 $l=2.75e-07 $layer=LI1_cond $X=1.15 $Y=2.405
+ $X2=1.15 $Y2=2.13
r29 15 21 2.60672 $w=4.18e-07 $l=9.5e-08 $layer=LI1_cond $X=1.15 $Y=2.035
+ $X2=1.15 $Y2=2.13
r30 15 30 7.36464 $w=4.18e-07 $l=1.15e-07 $layer=LI1_cond $X=1.15 $Y=2.035
+ $X2=1.15 $Y2=1.92
r31 11 13 24.6002 $w=2.58e-07 $l=5.55e-07 $layer=LI1_cond $X=1.695 $Y=0.975
+ $X2=1.695 $Y2=0.42
r32 9 11 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.565 $Y=1.06
+ $X2=1.695 $Y2=0.975
r33 9 10 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.565 $Y=1.06
+ $X2=1.36 $Y2=1.06
r34 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.275 $Y=1.145
+ $X2=1.36 $Y2=1.06
r35 7 30 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.275 $Y=1.145
+ $X2=1.275 $Y2=1.92
r36 2 15 400 $w=1.7e-07 $l=3.55106e-07 $layer=licon1_PDIFF $count=1 $X=0.92
+ $Y=1.835 $X2=1.145 $Y2=2.095
r37 2 27 400 $w=1.7e-07 $l=1.22233e-06 $layer=licon1_PDIFF $count=1 $X=0.92
+ $Y=1.835 $X2=1.145 $Y2=2.95
r38 1 13 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.52
+ $Y=0.235 $X2=1.66 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_1%A_29_47# 1 2 7 9 11 15
r27 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.23 $Y=0.635
+ $X2=1.23 $Y2=0.36
r28 12 18 2.87515 $w=4.05e-07 $l=1.35e-07 $layer=LI1_cond $X=0.375 $Y=0.837
+ $X2=0.24 $Y2=0.837
r29 11 13 14.1419 $w=4.05e-07 $l=4.27701e-07 $layer=LI1_cond $X=0.818 $Y=0.837
+ $X2=1.23 $Y2=0.805
r30 11 12 12.6057 $w=4.03e-07 $l=4.43e-07 $layer=LI1_cond $X=0.818 $Y=0.837
+ $X2=0.375 $Y2=0.837
r31 7 18 4.30208 $w=2.7e-07 $l=2.02e-07 $layer=LI1_cond $X=0.24 $Y=0.635
+ $X2=0.24 $Y2=0.837
r32 7 9 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.24 $Y=0.635
+ $X2=0.24 $Y2=0.43
r33 2 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.36
r34 1 18 182 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.93
r35 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_1%VGND 1 6 8 10 17 18 21
r27 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r28 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r29 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.73
+ $Y2=0
r30 15 17 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.68
+ $Y2=0
r31 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r32 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.73
+ $Y2=0
r34 10 12 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.24
+ $Y2=0
r35 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r36 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r37 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085 $X2=0.73
+ $Y2=0
r38 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r39 1 6 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

