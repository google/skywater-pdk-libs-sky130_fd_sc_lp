* File: sky130_fd_sc_lp__a221oi_0.pxi.spice
* Created: Fri Aug 28 09:53:02 2020
* 
x_PM_SKY130_FD_SC_LP__A221OI_0%C1 N_C1_M1009_g N_C1_c_75_n N_C1_M1007_g
+ N_C1_c_80_n C1 C1 C1 N_C1_c_77_n PM_SKY130_FD_SC_LP__A221OI_0%C1
x_PM_SKY130_FD_SC_LP__A221OI_0%B2 N_B2_M1000_g N_B2_M1002_g N_B2_c_116_n
+ N_B2_c_122_n B2 B2 N_B2_c_118_n N_B2_c_119_n B2
+ PM_SKY130_FD_SC_LP__A221OI_0%B2
x_PM_SKY130_FD_SC_LP__A221OI_0%B1 N_B1_M1001_g N_B1_c_177_n N_B1_M1008_g
+ N_B1_c_178_n N_B1_c_179_n N_B1_c_180_n N_B1_c_171_n N_B1_c_172_n N_B1_c_173_n
+ B1 B1 B1 B1 N_B1_c_174_n N_B1_c_175_n N_B1_c_176_n
+ PM_SKY130_FD_SC_LP__A221OI_0%B1
x_PM_SKY130_FD_SC_LP__A221OI_0%A1 N_A1_M1003_g N_A1_M1006_g N_A1_c_230_n
+ N_A1_c_234_n A1 A1 N_A1_c_232_n PM_SKY130_FD_SC_LP__A221OI_0%A1
x_PM_SKY130_FD_SC_LP__A221OI_0%A2 N_A2_M1004_g N_A2_c_279_n N_A2_M1005_g A2 A2
+ N_A2_c_285_n N_A2_c_282_n PM_SKY130_FD_SC_LP__A221OI_0%A2
x_PM_SKY130_FD_SC_LP__A221OI_0%Y N_Y_M1009_s N_Y_M1001_d N_Y_M1007_s N_Y_c_322_n
+ N_Y_c_323_n N_Y_c_342_n N_Y_c_343_n N_Y_c_324_n Y Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__A221OI_0%Y
x_PM_SKY130_FD_SC_LP__A221OI_0%A_156_487# N_A_156_487#_M1007_d
+ N_A_156_487#_M1008_d N_A_156_487#_c_372_n N_A_156_487#_c_373_n
+ N_A_156_487#_c_374_n N_A_156_487#_c_375_n
+ PM_SKY130_FD_SC_LP__A221OI_0%A_156_487#
x_PM_SKY130_FD_SC_LP__A221OI_0%A_242_487# N_A_242_487#_M1002_d
+ N_A_242_487#_M1004_d N_A_242_487#_c_412_n N_A_242_487#_c_408_n
+ N_A_242_487#_c_409_n PM_SKY130_FD_SC_LP__A221OI_0%A_242_487#
x_PM_SKY130_FD_SC_LP__A221OI_0%VPWR N_VPWR_M1003_d N_VPWR_c_430_n N_VPWR_c_431_n
+ N_VPWR_c_432_n VPWR N_VPWR_c_433_n N_VPWR_c_429_n
+ PM_SKY130_FD_SC_LP__A221OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A221OI_0%VGND N_VGND_M1009_d N_VGND_M1005_d N_VGND_c_463_n
+ N_VGND_c_464_n VGND N_VGND_c_465_n N_VGND_c_466_n N_VGND_c_467_n
+ N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n PM_SKY130_FD_SC_LP__A221OI_0%VGND
cc_1 VNB N_C1_M1009_g 0.0479066f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_2 VNB N_C1_c_75_n 0.0189931f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.703
cc_3 VNB C1 0.00516937f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C1_c_77_n 0.0184417f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.375
cc_5 VNB N_B2_M1000_g 0.0484625f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_6 VNB N_B2_c_116_n 0.00976743f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.88
cc_7 VNB B2 0.00170357f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_B2_c_118_n 0.0153219f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.375
cc_9 VNB N_B2_c_119_n 0.00596961f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.21
cc_10 VNB N_B1_c_171_n 0.0223196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_c_172_n 0.0325984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_173_n 0.0320015f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.375
cc_13 VNB N_B1_c_174_n 0.0362271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_175_n 0.016978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_c_176_n 0.0224795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_M1006_g 0.0470746f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.88
cc_17 VNB N_A1_c_230_n 0.024459f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.88
cc_18 VNB A1 0.00580421f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_19 VNB N_A1_c_232_n 0.0116307f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.375
cc_20 VNB N_A2_c_279_n 0.0166295f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.387
cc_21 VNB N_A2_M1005_g 0.0529883f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.755
cc_22 VNB A2 0.00747704f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.88
cc_23 VNB N_A2_c_282_n 0.0104297f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.21
cc_24 VNB N_Y_c_322_n 0.0193082f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_25 VNB N_Y_c_323_n 0.00121229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_324_n 0.0168177f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.375
cc_27 VNB Y 0.0113548f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.21
cc_28 VNB Y 0.0309246f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.905
cc_29 VNB N_VPWR_c_429_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_463_n 0.00496638f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.755
cc_31 VNB N_VGND_c_464_n 0.017485f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_32 VNB N_VGND_c_465_n 0.0194672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_466_n 0.0409141f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.905
cc_34 VNB N_VGND_c_467_n 0.022032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_468_n 0.198888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_469_n 0.00420624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_470_n 0.00510915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_C1_c_75_n 0.00334336f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.703
cc_39 VPB N_C1_M1007_g 0.0454431f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.755
cc_40 VPB N_C1_c_80_n 0.0190133f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.88
cc_41 VPB C1 0.00173234f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_42 VPB C1 0.00675862f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_43 VPB N_B2_M1002_g 0.0339093f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=1.88
cc_44 VPB N_B2_c_116_n 0.0116702f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.88
cc_45 VPB N_B2_c_122_n 0.0153125f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_46 VPB B2 0.0024136f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_47 VPB N_B1_c_177_n 0.0188087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_B1_c_178_n 0.0130969f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.755
cc_49 VPB N_B1_c_179_n 0.0228069f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.88
cc_50 VPB N_B1_c_180_n 0.0208555f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_51 VPB N_B1_c_172_n 0.0166077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_B1_c_173_n 0.0154843f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.375
cc_53 VPB N_A1_M1003_g 0.0361241f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_54 VPB N_A1_c_234_n 0.0154101f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_55 VPB A1 0.00211554f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_56 VPB N_A1_c_232_n 0.0119748f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.375
cc_57 VPB N_A2_M1004_g 0.0366673f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_58 VPB A2 0.00240545f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.88
cc_59 VPB N_A2_c_285_n 0.0344043f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.375
cc_60 VPB N_A2_c_282_n 0.00264128f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.21
cc_61 VPB Y 0.0379718f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.905
cc_62 VPB Y 0.039243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_156_487#_c_372_n 0.0100886f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=1.88
cc_64 VPB N_A_156_487#_c_373_n 0.00120843f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.755
cc_65 VPB N_A_156_487#_c_374_n 0.0412865f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.88
cc_66 VPB N_A_156_487#_c_375_n 0.0327779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_242_487#_c_408_n 0.00179423f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_68 VPB N_A_242_487#_c_409_n 0.00171433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_430_n 0.00336216f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.703
cc_70 VPB N_VPWR_c_431_n 0.0480325f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.755
cc_71 VPB N_VPWR_c_432_n 0.00525195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_433_n 0.0328868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_429_n 0.0725323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 N_C1_M1009_g N_B2_M1000_g 0.0241793f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_75 C1 N_B2_M1000_g 6.52403e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_C1_c_77_n N_B2_M1000_g 0.0124625f $X=0.615 $Y=1.375 $X2=0 $Y2=0
cc_77 N_C1_M1007_g N_B2_M1002_g 0.0241299f $X=0.705 $Y=2.755 $X2=0 $Y2=0
cc_78 C1 N_B2_M1002_g 0.0023895f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_79 N_C1_c_80_n N_B2_c_116_n 0.0124625f $X=0.602 $Y=1.88 $X2=0 $Y2=0
cc_80 N_C1_M1007_g N_B2_c_122_n 0.0124625f $X=0.705 $Y=2.755 $X2=0 $Y2=0
cc_81 C1 N_B2_c_122_n 0.00124354f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_82 C1 B2 0.0416769f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 C1 B2 0.00477749f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_84 N_C1_c_77_n B2 6.75702e-19 $X=0.615 $Y=1.375 $X2=0 $Y2=0
cc_85 N_C1_c_75_n N_B2_c_118_n 0.0124625f $X=0.602 $Y=1.703 $X2=0 $Y2=0
cc_86 C1 N_B2_c_118_n 0.00292718f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 C1 N_B2_c_119_n 0.0156393f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_C1_M1009_g N_Y_c_322_n 0.00387498f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_89 N_C1_M1009_g N_Y_c_323_n 5.58244e-19 $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_90 N_C1_M1009_g N_Y_c_324_n 0.0201739f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_91 C1 N_Y_c_324_n 0.024462f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_92 N_C1_c_77_n N_Y_c_324_n 0.00134056f $X=0.615 $Y=1.375 $X2=0 $Y2=0
cc_93 N_C1_M1009_g Y 0.024593f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_94 N_C1_M1007_g Y 0.00756296f $X=0.705 $Y=2.755 $X2=0 $Y2=0
cc_95 C1 Y 0.0546862f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_96 C1 Y 0.0171628f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_97 N_C1_M1007_g Y 0.00774782f $X=0.705 $Y=2.755 $X2=0 $Y2=0
cc_98 N_C1_c_80_n Y 0.00391531f $X=0.602 $Y=1.88 $X2=0 $Y2=0
cc_99 C1 Y 0.00765419f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_100 N_C1_M1007_g N_A_156_487#_c_372_n 0.00353962f $X=0.705 $Y=2.755 $X2=0
+ $Y2=0
cc_101 N_C1_M1007_g N_VPWR_c_431_n 0.00529818f $X=0.705 $Y=2.755 $X2=0 $Y2=0
cc_102 N_C1_M1007_g N_VPWR_c_429_n 0.0109004f $X=0.705 $Y=2.755 $X2=0 $Y2=0
cc_103 N_C1_M1009_g N_VGND_c_463_n 0.00318338f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_104 N_C1_M1009_g N_VGND_c_465_n 0.00585385f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_105 N_C1_M1009_g N_VGND_c_468_n 0.00757798f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_106 N_B2_M1000_g N_B1_c_174_n 0.0217466f $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_107 N_B2_c_119_n N_B1_c_174_n 6.41898e-19 $X=1.182 $Y=1.377 $X2=0 $Y2=0
cc_108 N_B2_M1000_g N_B1_c_175_n 0.0360084f $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_109 N_B2_M1000_g N_B1_c_176_n 2.70847e-19 $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_110 N_B2_c_119_n N_B1_c_176_n 0.0020603f $X=1.182 $Y=1.377 $X2=0 $Y2=0
cc_111 N_B2_M1002_g N_A1_M1003_g 0.0240542f $X=1.135 $Y=2.755 $X2=0 $Y2=0
cc_112 N_B2_c_119_n N_A1_M1006_g 6.67896e-19 $X=1.182 $Y=1.377 $X2=0 $Y2=0
cc_113 B2 N_A1_c_230_n 0.00195285f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B2_c_118_n N_A1_c_230_n 0.0120899f $X=1.155 $Y=1.5 $X2=0 $Y2=0
cc_115 N_B2_c_122_n N_A1_c_234_n 0.0120899f $X=1.155 $Y=2.005 $X2=0 $Y2=0
cc_116 N_B2_M1000_g A1 6.60754e-19 $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_117 B2 A1 0.0496996f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B2_c_118_n A1 0.00189762f $X=1.155 $Y=1.5 $X2=0 $Y2=0
cc_119 N_B2_c_119_n A1 0.0163205f $X=1.182 $Y=1.377 $X2=0 $Y2=0
cc_120 N_B2_c_116_n N_A1_c_232_n 0.0120899f $X=1.155 $Y=1.84 $X2=0 $Y2=0
cc_121 N_B2_M1000_g N_Y_c_323_n 0.00500806f $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_122 N_B2_M1000_g N_Y_c_342_n 0.0106317f $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B2_c_119_n N_Y_c_343_n 0.00566233f $X=1.182 $Y=1.377 $X2=0 $Y2=0
cc_124 N_B2_M1000_g N_Y_c_324_n 0.00964608f $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_125 N_B2_c_119_n N_Y_c_324_n 0.0154042f $X=1.182 $Y=1.377 $X2=0 $Y2=0
cc_126 N_B2_M1002_g N_A_156_487#_c_372_n 0.00870222f $X=1.135 $Y=2.755 $X2=0
+ $Y2=0
cc_127 N_B2_c_122_n N_A_156_487#_c_372_n 0.00202048f $X=1.155 $Y=2.005 $X2=0
+ $Y2=0
cc_128 B2 N_A_156_487#_c_372_n 0.0133466f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B2_M1002_g N_A_156_487#_c_373_n 0.00947124f $X=1.135 $Y=2.755 $X2=0
+ $Y2=0
cc_130 N_B2_M1002_g N_A_156_487#_c_374_n 0.00732984f $X=1.135 $Y=2.755 $X2=0
+ $Y2=0
cc_131 N_B2_c_122_n N_A_156_487#_c_374_n 0.00299108f $X=1.155 $Y=2.005 $X2=0
+ $Y2=0
cc_132 B2 N_A_156_487#_c_374_n 0.0182685f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_133 N_B2_M1002_g N_A_242_487#_c_408_n 0.00501863f $X=1.135 $Y=2.755 $X2=0
+ $Y2=0
cc_134 N_B2_M1002_g N_VPWR_c_431_n 0.00441574f $X=1.135 $Y=2.755 $X2=0 $Y2=0
cc_135 N_B2_M1002_g N_VPWR_c_429_n 0.00795405f $X=1.135 $Y=2.755 $X2=0 $Y2=0
cc_136 N_B2_M1000_g N_VGND_c_463_n 0.00572707f $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_137 N_B2_M1000_g N_VGND_c_466_n 0.00377689f $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_138 N_B2_M1000_g N_VGND_c_468_n 0.00575065f $X=1.065 $Y=0.445 $X2=0 $Y2=0
cc_139 N_B1_c_174_n N_A1_M1006_g 0.0218601f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_140 N_B1_c_175_n N_A1_M1006_g 0.0105532f $X=1.515 $Y=0.765 $X2=0 $Y2=0
cc_141 N_B1_c_176_n N_A1_M1006_g 0.0173028f $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_142 N_B1_c_174_n N_A1_c_230_n 0.00601589f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_143 N_B1_c_176_n N_A1_c_230_n 0.00113544f $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_144 N_B1_c_174_n A1 0.00137108f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_145 N_B1_c_176_n A1 0.0294907f $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_146 N_B1_c_179_n N_A2_M1004_g 0.0224188f $X=2.865 $Y=2.275 $X2=0 $Y2=0
cc_147 N_B1_c_180_n N_A2_M1004_g 0.00541244f $X=2.965 $Y=2.035 $X2=0 $Y2=0
cc_148 N_B1_c_172_n N_A2_c_279_n 0.00458493f $X=2.975 $Y=1.53 $X2=0 $Y2=0
cc_149 N_B1_c_173_n N_A2_c_279_n 0.0198796f $X=2.975 $Y=1.53 $X2=0 $Y2=0
cc_150 N_B1_c_176_n N_A2_c_279_n 9.09231e-19 $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_151 N_B1_c_172_n N_A2_M1005_g 0.00630051f $X=2.975 $Y=1.53 $X2=0 $Y2=0
cc_152 N_B1_c_176_n N_A2_M1005_g 0.0165755f $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_153 N_B1_c_172_n A2 0.0659157f $X=2.975 $Y=1.53 $X2=0 $Y2=0
cc_154 N_B1_c_173_n A2 6.86429e-19 $X=2.975 $Y=1.53 $X2=0 $Y2=0
cc_155 N_B1_c_176_n A2 0.0430369f $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_156 N_B1_c_176_n N_A2_c_285_n 3.4028e-19 $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_157 N_B1_c_180_n N_A2_c_282_n 0.0198796f $X=2.965 $Y=2.035 $X2=0 $Y2=0
cc_158 N_B1_c_174_n N_Y_c_323_n 2.85435e-19 $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_159 N_B1_c_175_n N_Y_c_323_n 0.00222435f $X=1.515 $Y=0.765 $X2=0 $Y2=0
cc_160 N_B1_c_174_n N_Y_c_343_n 0.00332855f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_161 N_B1_c_175_n N_Y_c_343_n 0.0114914f $X=1.515 $Y=0.765 $X2=0 $Y2=0
cc_162 N_B1_c_176_n N_Y_c_343_n 0.0352933f $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_163 N_B1_c_174_n N_Y_c_324_n 8.80896e-19 $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_164 N_B1_c_176_n N_Y_c_324_n 0.0195481f $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_165 N_B1_c_178_n N_A_156_487#_c_374_n 0.00534368f $X=2.865 $Y=2.2 $X2=0 $Y2=0
cc_166 N_B1_c_179_n N_A_156_487#_c_374_n 0.0166565f $X=2.865 $Y=2.275 $X2=0
+ $Y2=0
cc_167 N_B1_c_180_n N_A_156_487#_c_374_n 0.00583474f $X=2.965 $Y=2.035 $X2=0
+ $Y2=0
cc_168 N_B1_c_172_n N_A_156_487#_c_374_n 0.0340429f $X=2.975 $Y=1.53 $X2=0 $Y2=0
cc_169 N_B1_c_177_n N_A_156_487#_c_375_n 0.0159666f $X=2.695 $Y=2.35 $X2=0 $Y2=0
cc_170 N_B1_c_179_n N_A_156_487#_c_375_n 0.0052604f $X=2.865 $Y=2.275 $X2=0
+ $Y2=0
cc_171 N_B1_c_177_n N_A_242_487#_c_409_n 0.00690653f $X=2.695 $Y=2.35 $X2=0
+ $Y2=0
cc_172 N_B1_c_177_n N_VPWR_c_430_n 8.8746e-19 $X=2.695 $Y=2.35 $X2=0 $Y2=0
cc_173 N_B1_c_177_n N_VPWR_c_433_n 0.00529818f $X=2.695 $Y=2.35 $X2=0 $Y2=0
cc_174 N_B1_c_177_n N_VPWR_c_429_n 0.0110293f $X=2.695 $Y=2.35 $X2=0 $Y2=0
cc_175 N_B1_c_176_n N_VGND_c_464_n 0.0243027f $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_176 N_B1_c_175_n N_VGND_c_466_n 0.00363059f $X=1.515 $Y=0.765 $X2=0 $Y2=0
cc_177 N_B1_c_171_n N_VGND_c_468_n 0.0189186f $X=2.977 $Y=1.015 $X2=0 $Y2=0
cc_178 N_B1_c_175_n N_VGND_c_468_n 0.00556891f $X=1.515 $Y=0.765 $X2=0 $Y2=0
cc_179 N_B1_c_176_n N_VGND_c_468_n 0.0194231f $X=2.75 $Y=0.897 $X2=0 $Y2=0
cc_180 N_A1_M1003_g N_A2_M1004_g 0.0359062f $X=1.695 $Y=2.755 $X2=0 $Y2=0
cc_181 N_A1_c_234_n N_A2_M1004_g 0.00910131f $X=1.73 $Y=2.005 $X2=0 $Y2=0
cc_182 N_A1_c_230_n N_A2_c_279_n 0.00949617f $X=1.802 $Y=1.485 $X2=0 $Y2=0
cc_183 A1 N_A2_c_279_n 3.07037e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A1_c_232_n N_A2_c_279_n 0.00646312f $X=1.73 $Y=1.5 $X2=0 $Y2=0
cc_185 N_A1_M1006_g N_A2_M1005_g 0.0662288f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A1_M1006_g A2 0.00240519f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_187 A1 A2 0.0641339f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A1_c_232_n A2 0.00327073f $X=1.73 $Y=1.5 $X2=0 $Y2=0
cc_189 A1 N_A2_c_285_n 3.029e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A1_c_232_n N_A2_c_285_n 0.00910131f $X=1.73 $Y=1.5 $X2=0 $Y2=0
cc_191 N_A1_M1006_g N_Y_c_343_n 0.00557832f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A1_M1003_g N_A_156_487#_c_372_n 7.33361e-19 $X=1.695 $Y=2.755 $X2=0
+ $Y2=0
cc_193 N_A1_M1003_g N_A_156_487#_c_374_n 0.0114246f $X=1.695 $Y=2.755 $X2=0
+ $Y2=0
cc_194 N_A1_c_230_n N_A_156_487#_c_374_n 0.0036662f $X=1.802 $Y=1.485 $X2=0
+ $Y2=0
cc_195 N_A1_c_234_n N_A_156_487#_c_374_n 0.00491229f $X=1.73 $Y=2.005 $X2=0
+ $Y2=0
cc_196 A1 N_A_156_487#_c_374_n 0.0273353f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A1_M1003_g N_A_242_487#_c_412_n 0.0092159f $X=1.695 $Y=2.755 $X2=0
+ $Y2=0
cc_198 N_A1_M1003_g N_A_242_487#_c_408_n 0.00685497f $X=1.695 $Y=2.755 $X2=0
+ $Y2=0
cc_199 N_A1_M1003_g N_VPWR_c_430_n 0.00432115f $X=1.695 $Y=2.755 $X2=0 $Y2=0
cc_200 N_A1_M1003_g N_VPWR_c_431_n 0.00404007f $X=1.695 $Y=2.755 $X2=0 $Y2=0
cc_201 N_A1_M1003_g N_VPWR_c_429_n 0.00608234f $X=1.695 $Y=2.755 $X2=0 $Y2=0
cc_202 N_A1_M1006_g N_VGND_c_464_n 0.00225331f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_203 N_A1_M1006_g N_VGND_c_466_n 0.00563152f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_204 N_A1_M1006_g N_VGND_c_468_n 0.00642886f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A2_M1005_g N_Y_c_343_n 9.10137e-19 $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_206 N_A2_M1004_g N_A_156_487#_c_374_n 0.0114096f $X=2.195 $Y=2.755 $X2=0
+ $Y2=0
cc_207 A2 N_A_156_487#_c_374_n 0.0406804f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_208 N_A2_c_285_n N_A_156_487#_c_374_n 0.00835797f $X=2.415 $Y=1.825 $X2=0
+ $Y2=0
cc_209 N_A2_M1004_g N_A_242_487#_c_412_n 0.0128361f $X=2.195 $Y=2.755 $X2=0
+ $Y2=0
cc_210 N_A2_M1004_g N_A_242_487#_c_408_n 3.10406e-19 $X=2.195 $Y=2.755 $X2=0
+ $Y2=0
cc_211 N_A2_M1004_g N_VPWR_c_430_n 0.00765971f $X=2.195 $Y=2.755 $X2=0 $Y2=0
cc_212 N_A2_M1004_g N_VPWR_c_433_n 0.0034441f $X=2.195 $Y=2.755 $X2=0 $Y2=0
cc_213 N_A2_M1004_g N_VPWR_c_429_n 0.0043427f $X=2.195 $Y=2.755 $X2=0 $Y2=0
cc_214 N_A2_M1005_g N_VGND_c_464_n 0.0128416f $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A2_M1005_g N_VGND_c_466_n 0.00486043f $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_216 N_A2_M1005_g N_VGND_c_468_n 0.00441216f $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_217 Y N_A_156_487#_c_372_n 0.0102253f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_218 Y N_A_156_487#_c_372_n 0.00279957f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_219 Y N_VPWR_c_431_n 0.0331972f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_220 Y N_VPWR_c_429_n 0.0192324f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_221 N_Y_c_342_n N_VGND_c_463_n 0.0264119f $X=1.17 $Y=0.445 $X2=0 $Y2=0
cc_222 N_Y_c_324_n N_VGND_c_463_n 0.016971f $X=1 $Y=0.895 $X2=0 $Y2=0
cc_223 N_Y_c_343_n N_VGND_c_464_n 0.0108275f $X=1.715 $Y=0.445 $X2=0 $Y2=0
cc_224 N_Y_c_322_n N_VGND_c_465_n 0.0134923f $X=0.285 $Y=0.445 $X2=0 $Y2=0
cc_225 N_Y_c_342_n N_VGND_c_466_n 0.00911951f $X=1.17 $Y=0.445 $X2=0 $Y2=0
cc_226 N_Y_c_343_n N_VGND_c_466_n 0.0364511f $X=1.715 $Y=0.445 $X2=0 $Y2=0
cc_227 N_Y_M1009_s N_VGND_c_468_n 0.00236029f $X=0.16 $Y=0.235 $X2=0 $Y2=0
cc_228 N_Y_M1001_d N_VGND_c_468_n 0.00290843f $X=1.53 $Y=0.235 $X2=0 $Y2=0
cc_229 N_Y_c_322_n N_VGND_c_468_n 0.00894849f $X=0.285 $Y=0.445 $X2=0 $Y2=0
cc_230 N_Y_c_342_n N_VGND_c_468_n 0.00587796f $X=1.17 $Y=0.445 $X2=0 $Y2=0
cc_231 N_Y_c_343_n N_VGND_c_468_n 0.0268715f $X=1.715 $Y=0.445 $X2=0 $Y2=0
cc_232 N_Y_c_324_n N_VGND_c_468_n 0.0142087f $X=1 $Y=0.895 $X2=0 $Y2=0
cc_233 N_Y_c_343_n A_228_47# 0.00377228f $X=1.715 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_234 N_A_156_487#_c_374_n N_A_242_487#_c_412_n 0.0422043f $X=2.815 $Y=2.22
+ $X2=0 $Y2=0
cc_235 N_A_156_487#_c_373_n N_A_242_487#_c_408_n 0.0473207f $X=0.92 $Y=2.56
+ $X2=0 $Y2=0
cc_236 N_A_156_487#_c_374_n N_A_242_487#_c_408_n 0.0243022f $X=2.815 $Y=2.22
+ $X2=0 $Y2=0
cc_237 N_A_156_487#_c_374_n N_A_242_487#_c_409_n 0.0237727f $X=2.815 $Y=2.22
+ $X2=0 $Y2=0
cc_238 N_A_156_487#_c_373_n N_VPWR_c_431_n 0.0197784f $X=0.92 $Y=2.56 $X2=0
+ $Y2=0
cc_239 N_A_156_487#_c_375_n N_VPWR_c_433_n 0.022733f $X=2.98 $Y=2.58 $X2=0 $Y2=0
cc_240 N_A_156_487#_c_373_n N_VPWR_c_429_n 0.0119688f $X=0.92 $Y=2.56 $X2=0
+ $Y2=0
cc_241 N_A_156_487#_c_375_n N_VPWR_c_429_n 0.0127519f $X=2.98 $Y=2.58 $X2=0
+ $Y2=0
cc_242 N_A_242_487#_c_412_n N_VPWR_M1003_d 0.00485551f $X=2.315 $Y=2.565
+ $X2=-0.19 $Y2=1.655
cc_243 N_A_242_487#_c_412_n N_VPWR_c_430_n 0.0199771f $X=2.315 $Y=2.565 $X2=0
+ $Y2=0
cc_244 N_A_242_487#_c_412_n N_VPWR_c_431_n 0.00225191f $X=2.315 $Y=2.565 $X2=0
+ $Y2=0
cc_245 N_A_242_487#_c_408_n N_VPWR_c_431_n 0.0208206f $X=1.48 $Y=2.59 $X2=0
+ $Y2=0
cc_246 N_A_242_487#_c_412_n N_VPWR_c_433_n 0.00225806f $X=2.315 $Y=2.565 $X2=0
+ $Y2=0
cc_247 N_A_242_487#_c_409_n N_VPWR_c_433_n 0.0204446f $X=2.48 $Y=2.59 $X2=0
+ $Y2=0
cc_248 N_A_242_487#_c_412_n N_VPWR_c_429_n 0.00961527f $X=2.315 $Y=2.565 $X2=0
+ $Y2=0
cc_249 N_A_242_487#_c_408_n N_VPWR_c_429_n 0.0125907f $X=1.48 $Y=2.59 $X2=0
+ $Y2=0
cc_250 N_A_242_487#_c_409_n N_VPWR_c_429_n 0.0125907f $X=2.48 $Y=2.59 $X2=0
+ $Y2=0
cc_251 N_VGND_c_468_n A_228_47# 0.00193888f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_252 N_VGND_c_468_n A_408_47# 0.00330611f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
