# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__inv_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.395000 3.815000 1.585000 ;
        RECT 2.060000 1.160000 2.365000 1.385000 ;
        RECT 2.060000 1.385000 3.815000 1.395000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.045000 1.890000 1.215000 ;
        RECT 0.085000 1.215000 0.255000 1.755000 ;
        RECT 0.085000 1.755000 4.225000 1.925000 ;
        RECT 0.815000 0.255000 1.075000 1.045000 ;
        RECT 0.815000 1.925000 1.075000 3.075000 ;
        RECT 1.675000 0.255000 1.935000 0.820000 ;
        RECT 1.675000 0.820000 2.795000 0.990000 ;
        RECT 1.675000 0.990000 1.890000 1.045000 ;
        RECT 1.675000 1.925000 1.935000 3.075000 ;
        RECT 2.535000 0.255000 2.795000 0.820000 ;
        RECT 2.535000 0.990000 2.795000 1.045000 ;
        RECT 2.535000 1.045000 4.225000 1.215000 ;
        RECT 2.535000 1.925000 2.795000 3.075000 ;
        RECT 3.395000 0.255000 3.655000 1.045000 ;
        RECT 3.395000 1.925000 3.655000 3.075000 ;
        RECT 3.985000 1.215000 4.225000 1.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.350000  0.085000 0.645000 0.875000 ;
      RECT 0.350000  2.105000 0.645000 3.245000 ;
      RECT 1.245000  0.085000 1.505000 0.875000 ;
      RECT 1.245000  2.095000 1.505000 3.245000 ;
      RECT 2.105000  0.085000 2.365000 0.650000 ;
      RECT 2.105000  2.095000 2.365000 3.245000 ;
      RECT 2.965000  0.085000 3.225000 0.875000 ;
      RECT 2.965000  2.095000 3.225000 3.245000 ;
      RECT 3.825000  0.085000 4.120000 0.875000 ;
      RECT 3.825000  2.095000 4.120000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__inv_8
