* NGSPICE file created from sky130_fd_sc_lp__or4b_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or4b_m A B C D_N VGND VNB VPB VPWR X
M1000 a_338_397# a_38_125# a_215_125# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1001 X a_215_125# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.751e+11p ps=2.99e+06u
M1002 a_215_125# B VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=5.943e+11p ps=5.35e+06u
M1003 VGND D_N a_38_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 VPWR D_N a_38_125# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 a_215_125# a_38_125# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C a_215_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_215_125# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 a_410_397# C a_338_397# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 a_482_397# B a_410_397# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 VPWR A a_482_397# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A a_215_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

