* File: sky130_fd_sc_lp__o32ai_m.spice
* Created: Wed Sep  2 10:27:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32ai_m.pex.spice"
.subckt sky130_fd_sc_lp__o32ai_m  VNB VPB B1 B2 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_66_82#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1449 PD=0.7 PS=1.53 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.3
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1009 N_A_66_82#_M1009_d N_B2_M1009_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.7 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A3_M1006_g N_A_66_82#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_A_66_82#_M1003_d N_A2_M1003_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_66_82#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 A_179_535# N_B1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.21 PD=0.63 PS=1.84 NRD=23.443 NRS=110.222 M=1 R=2.8 SA=75000.4
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g A_179_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.8 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1008 A_337_535# N_A3_M1008_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0672
+ AS=0.0588 PD=0.74 PS=0.7 NRD=49.25 NRS=0 M=1 R=2.8 SA=75001.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1005 A_431_535# N_A2_M1005_g A_337_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0672 PD=0.63 PS=0.74 NRD=23.443 NRS=49.25 M=1 R=2.8 SA=75001.7 SB=75000.9
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g A_431_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.252
+ AS=0.0441 PD=2.04 PS=0.63 NRD=157.127 NRS=23.443 M=1 R=2.8 SA=75002 SB=75000.5
+ A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o32ai_m.pxi.spice"
*
.ends
*
*
