* File: sky130_fd_sc_lp__o21ba_1.pxi.spice
* Created: Wed Sep  2 10:16:42 2020
* 
x_PM_SKY130_FD_SC_LP__O21BA_1%A_84_28# N_A_84_28#_M1002_s N_A_84_28#_M1001_d
+ N_A_84_28#_c_67_n N_A_84_28#_M1005_g N_A_84_28#_M1008_g N_A_84_28#_c_69_n
+ N_A_84_28#_c_81_p N_A_84_28#_c_135_p N_A_84_28#_c_70_n N_A_84_28#_c_71_n
+ N_A_84_28#_c_72_n N_A_84_28#_c_73_n N_A_84_28#_c_95_p N_A_84_28#_c_102_p
+ N_A_84_28#_c_105_p N_A_84_28#_c_106_p N_A_84_28#_c_74_n N_A_84_28#_c_75_n
+ PM_SKY130_FD_SC_LP__O21BA_1%A_84_28#
x_PM_SKY130_FD_SC_LP__O21BA_1%B1_N N_B1_N_M1006_g N_B1_N_M1000_g B1_N B1_N
+ N_B1_N_c_152_n N_B1_N_c_153_n PM_SKY130_FD_SC_LP__O21BA_1%B1_N
x_PM_SKY130_FD_SC_LP__O21BA_1%A_281_138# N_A_281_138#_M1006_d
+ N_A_281_138#_M1000_d N_A_281_138#_c_183_n N_A_281_138#_M1002_g
+ N_A_281_138#_M1001_g N_A_281_138#_c_185_n N_A_281_138#_c_186_n
+ N_A_281_138#_c_187_n N_A_281_138#_c_191_n N_A_281_138#_c_188_n
+ N_A_281_138#_c_189_n PM_SKY130_FD_SC_LP__O21BA_1%A_281_138#
x_PM_SKY130_FD_SC_LP__O21BA_1%A2 N_A2_M1007_g N_A2_M1003_g A2 A2 N_A2_c_222_n
+ PM_SKY130_FD_SC_LP__O21BA_1%A2
x_PM_SKY130_FD_SC_LP__O21BA_1%A1 N_A1_M1009_g N_A1_M1004_g A1 N_A1_c_257_n
+ N_A1_c_258_n PM_SKY130_FD_SC_LP__O21BA_1%A1
x_PM_SKY130_FD_SC_LP__O21BA_1%X N_X_M1005_s N_X_M1008_s X X X X X X X
+ N_X_c_281_n N_X_c_284_n X PM_SKY130_FD_SC_LP__O21BA_1%X
x_PM_SKY130_FD_SC_LP__O21BA_1%VPWR N_VPWR_M1008_d N_VPWR_M1001_s N_VPWR_M1004_d
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n
+ N_VPWR_c_304_n VPWR N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n
+ N_VPWR_c_298_n PM_SKY130_FD_SC_LP__O21BA_1%VPWR
x_PM_SKY130_FD_SC_LP__O21BA_1%VGND N_VGND_M1005_d N_VGND_M1007_d N_VGND_c_343_n
+ N_VGND_c_344_n VGND N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n
+ N_VGND_c_348_n N_VGND_c_349_n N_VGND_c_350_n PM_SKY130_FD_SC_LP__O21BA_1%VGND
x_PM_SKY130_FD_SC_LP__O21BA_1%A_494_51# N_A_494_51#_M1002_d N_A_494_51#_M1009_d
+ N_A_494_51#_c_386_n N_A_494_51#_c_387_n N_A_494_51#_c_388_n
+ N_A_494_51#_c_389_n PM_SKY130_FD_SC_LP__O21BA_1%A_494_51#
cc_1 VNB N_A_84_28#_c_67_n 0.0223582f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A_84_28#_M1008_g 0.00673391f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_3 VNB N_A_84_28#_c_69_n 0.0022826f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.22
cc_4 VNB N_A_84_28#_c_70_n 0.00672468f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.87
cc_5 VNB N_A_84_28#_c_71_n 0.0254109f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=0.34
cc_6 VNB N_A_84_28#_c_72_n 0.00342101f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=0.34
cc_7 VNB N_A_84_28#_c_73_n 0.00336246f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=0.43
cc_8 VNB N_A_84_28#_c_74_n 0.00382633f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.385
cc_9 VNB N_A_84_28#_c_75_n 0.0408775f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_10 VNB N_B1_N_M1000_g 0.00594297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB B1_N 0.00264399f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_12 VNB N_B1_N_c_152_n 0.0351097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_N_c_153_n 0.0204534f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.22
cc_14 VNB N_A_281_138#_c_183_n 0.0204825f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_15 VNB N_A_281_138#_M1001_g 0.00565738f $X=-0.19 $Y=-0.245 $X2=0.695
+ $Y2=2.465
cc_16 VNB N_A_281_138#_c_185_n 0.0738337f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.04
cc_17 VNB N_A_281_138#_c_186_n 0.0114969f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.22
cc_18 VNB N_A_281_138#_c_187_n 0.00666233f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.425
cc_19 VNB N_A_281_138#_c_188_n 0.00157838f $X=-0.19 $Y=-0.245 $X2=2.192 $Y2=0.43
cc_20 VNB N_A_281_138#_c_189_n 0.00734155f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=2.012
cc_21 VNB N_A2_M1007_g 0.024424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A2 0.00717506f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.55
cc_23 VNB N_A2_c_222_n 0.0233959f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.04
cc_24 VNB N_A1_M1009_g 0.0283095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_M1004_g 0.00179511f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_26 VNB N_A1_c_257_n 0.0475599f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.04
cc_27 VNB N_A1_c_258_n 0.0114877f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.22
cc_28 VNB N_X_c_281_n 0.0654263f $X=-0.19 $Y=-0.245 $X2=2.192 $Y2=0.43
cc_29 VNB N_VPWR_c_298_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_343_n 0.00889273f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_31 VNB N_VGND_c_344_n 0.00626815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_345_n 0.0161846f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.955
cc_33 VNB N_VGND_c_346_n 0.0499757f $X=-0.19 $Y=-0.245 $X2=2.192 $Y2=0.425
cc_34 VNB N_VGND_c_347_n 0.0181857f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.385
cc_35 VNB N_VGND_c_348_n 0.238462f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.385
cc_36 VNB N_VGND_c_349_n 0.00602297f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.385
cc_37 VNB N_VGND_c_350_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=2.63 $Y2=2.01
cc_38 VNB N_A_494_51#_c_386_n 0.00120843f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_39 VNB N_A_494_51#_c_387_n 0.0145535f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_40 VNB N_A_494_51#_c_388_n 0.00337303f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_41 VNB N_A_494_51#_c_389_n 0.031954f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.22
cc_42 VPB N_A_84_28#_M1008_g 0.0267444f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_43 VPB N_A_84_28#_c_73_n 0.00343976f $X=-0.19 $Y=1.655 $X2=2.18 $Y2=0.43
cc_44 VPB N_B1_N_M1000_g 0.0285919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB B1_N 0.00246236f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.69
cc_46 VPB N_A_281_138#_M1001_g 0.0227747f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_47 VPB N_A_281_138#_c_191_n 0.00421112f $X=-0.19 $Y=1.655 $X2=2.192 $Y2=1.925
cc_48 VPB N_A_281_138#_c_188_n 0.00499911f $X=-0.19 $Y=1.655 $X2=2.192 $Y2=0.43
cc_49 VPB N_A2_M1003_g 0.0196172f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.22
cc_50 VPB A2 0.0149439f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.55
cc_51 VPB N_A2_c_222_n 0.00630939f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.04
cc_52 VPB N_A1_M1004_g 0.0263066f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.22
cc_53 VPB N_A1_c_258_n 0.00716831f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.22
cc_54 VPB X 0.0517099f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_55 VPB N_X_c_281_n 0.00932789f $X=-0.19 $Y=1.655 $X2=2.192 $Y2=0.43
cc_56 VPB N_X_c_284_n 0.0156412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_299_n 0.0396224f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_58 VPB N_VPWR_c_300_n 0.0336019f $X=-0.19 $Y=1.655 $X2=1.22 $Y2=0.425
cc_59 VPB N_VPWR_c_301_n 0.0106587f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=0.34
cc_60 VPB N_VPWR_c_302_n 0.0483963f $X=-0.19 $Y=1.655 $X2=2.192 $Y2=0.425
cc_61 VPB N_VPWR_c_303_n 0.0202129f $X=-0.19 $Y=1.655 $X2=2.31 $Y2=2.012
cc_62 VPB N_VPWR_c_304_n 0.00857067f $X=-0.19 $Y=1.655 $X2=2.66 $Y2=2.1
cc_63 VPB N_VPWR_c_305_n 0.0241211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_306_n 0.0289253f $X=-0.19 $Y=1.655 $X2=2.63 $Y2=2.01
cc_65 VPB N_VPWR_c_307_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_298_n 0.0774902f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 N_A_84_28#_M1008_g N_B1_N_M1000_g 0.015974f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A_84_28#_M1008_g B1_N 0.00380985f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_69 N_A_84_28#_c_69_n B1_N 7.62376e-19 $X=0.85 $Y=1.22 $X2=0 $Y2=0
cc_70 N_A_84_28#_c_81_p B1_N 0.0146298f $X=1.135 $Y=0.955 $X2=0 $Y2=0
cc_71 N_A_84_28#_c_74_n B1_N 0.0254078f $X=0.85 $Y=1.385 $X2=0 $Y2=0
cc_72 N_A_84_28#_c_75_n B1_N 3.07192e-19 $X=0.695 $Y=1.385 $X2=0 $Y2=0
cc_73 N_A_84_28#_c_81_p N_B1_N_c_152_n 0.00284256f $X=1.135 $Y=0.955 $X2=0 $Y2=0
cc_74 N_A_84_28#_c_74_n N_B1_N_c_152_n 0.00223028f $X=0.85 $Y=1.385 $X2=0 $Y2=0
cc_75 N_A_84_28#_c_75_n N_B1_N_c_152_n 0.0173669f $X=0.695 $Y=1.385 $X2=0 $Y2=0
cc_76 N_A_84_28#_c_67_n N_B1_N_c_153_n 0.00551887f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_77 N_A_84_28#_c_69_n N_B1_N_c_153_n 0.00172067f $X=0.85 $Y=1.22 $X2=0 $Y2=0
cc_78 N_A_84_28#_c_81_p N_B1_N_c_153_n 0.00606715f $X=1.135 $Y=0.955 $X2=0 $Y2=0
cc_79 N_A_84_28#_c_70_n N_B1_N_c_153_n 0.0178739f $X=1.22 $Y=0.87 $X2=0 $Y2=0
cc_80 N_A_84_28#_c_71_n N_B1_N_c_153_n 0.00429306f $X=2.075 $Y=0.34 $X2=0 $Y2=0
cc_81 N_A_84_28#_c_73_n N_B1_N_c_153_n 0.00672527f $X=2.18 $Y=0.43 $X2=0 $Y2=0
cc_82 N_A_84_28#_c_73_n N_A_281_138#_c_183_n 0.00580465f $X=2.18 $Y=0.43 $X2=0
+ $Y2=0
cc_83 N_A_84_28#_c_73_n N_A_281_138#_M1001_g 0.0100736f $X=2.18 $Y=0.43 $X2=0
+ $Y2=0
cc_84 N_A_84_28#_c_95_p N_A_281_138#_M1001_g 0.0182393f $X=2.525 $Y=2.012 $X2=0
+ $Y2=0
cc_85 N_A_84_28#_c_73_n N_A_281_138#_c_185_n 0.0271433f $X=2.18 $Y=0.43 $X2=0
+ $Y2=0
cc_86 N_A_84_28#_c_69_n N_A_281_138#_c_187_n 0.00589331f $X=0.85 $Y=1.22 $X2=0
+ $Y2=0
cc_87 N_A_84_28#_c_81_p N_A_281_138#_c_187_n 0.0140373f $X=1.135 $Y=0.955 $X2=0
+ $Y2=0
cc_88 N_A_84_28#_c_70_n N_A_281_138#_c_187_n 7.22177e-19 $X=1.22 $Y=0.87 $X2=0
+ $Y2=0
cc_89 N_A_84_28#_c_71_n N_A_281_138#_c_187_n 0.0153464f $X=2.075 $Y=0.34 $X2=0
+ $Y2=0
cc_90 N_A_84_28#_c_73_n N_A_281_138#_c_187_n 0.0541114f $X=2.18 $Y=0.43 $X2=0
+ $Y2=0
cc_91 N_A_84_28#_c_102_p N_A_281_138#_c_191_n 0.00967746f $X=2.31 $Y=2.012 $X2=0
+ $Y2=0
cc_92 N_A_84_28#_c_73_n N_A_281_138#_c_188_n 0.0191801f $X=2.18 $Y=0.43 $X2=0
+ $Y2=0
cc_93 N_A_84_28#_c_73_n N_A2_M1007_g 5.72261e-19 $X=2.18 $Y=0.43 $X2=0 $Y2=0
cc_94 N_A_84_28#_c_105_p N_A2_M1003_g 0.00371196f $X=2.66 $Y=2.1 $X2=0 $Y2=0
cc_95 N_A_84_28#_c_106_p N_A2_M1003_g 0.0200396f $X=2.63 $Y=2.435 $X2=0 $Y2=0
cc_96 N_A_84_28#_c_73_n A2 0.0273928f $X=2.18 $Y=0.43 $X2=0 $Y2=0
cc_97 N_A_84_28#_c_105_p A2 0.0200863f $X=2.66 $Y=2.1 $X2=0 $Y2=0
cc_98 N_A_84_28#_c_73_n N_A2_c_222_n 4.91707e-19 $X=2.18 $Y=0.43 $X2=0 $Y2=0
cc_99 N_A_84_28#_c_105_p N_A2_c_222_n 2.3741e-19 $X=2.66 $Y=2.1 $X2=0 $Y2=0
cc_100 N_A_84_28#_c_105_p N_A1_M1004_g 5.37969e-19 $X=2.66 $Y=2.1 $X2=0 $Y2=0
cc_101 N_A_84_28#_c_106_p N_A1_M1004_g 0.00300918f $X=2.63 $Y=2.435 $X2=0 $Y2=0
cc_102 N_A_84_28#_c_67_n N_X_c_281_n 0.015677f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_103 N_A_84_28#_M1008_g N_X_c_281_n 0.00902497f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A_84_28#_c_69_n N_X_c_281_n 0.00630628f $X=0.85 $Y=1.22 $X2=0 $Y2=0
cc_105 N_A_84_28#_c_74_n N_X_c_281_n 0.0249965f $X=0.85 $Y=1.385 $X2=0 $Y2=0
cc_106 N_A_84_28#_M1008_g N_X_c_284_n 0.00377403f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_84_28#_c_74_n N_X_c_284_n 5.45223e-19 $X=0.85 $Y=1.385 $X2=0 $Y2=0
cc_108 N_A_84_28#_c_75_n N_X_c_284_n 0.00655331f $X=0.695 $Y=1.385 $X2=0 $Y2=0
cc_109 N_A_84_28#_c_73_n N_VPWR_M1001_s 0.00148947f $X=2.18 $Y=0.43 $X2=0 $Y2=0
cc_110 N_A_84_28#_c_102_p N_VPWR_M1001_s 0.00508878f $X=2.31 $Y=2.012 $X2=0
+ $Y2=0
cc_111 N_A_84_28#_M1008_g N_VPWR_c_299_n 0.02728f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_84_28#_c_74_n N_VPWR_c_299_n 0.00750783f $X=0.85 $Y=1.385 $X2=0 $Y2=0
cc_113 N_A_84_28#_c_95_p N_VPWR_c_300_n 0.00178974f $X=2.525 $Y=2.012 $X2=0
+ $Y2=0
cc_114 N_A_84_28#_c_102_p N_VPWR_c_300_n 0.0169053f $X=2.31 $Y=2.012 $X2=0 $Y2=0
cc_115 N_A_84_28#_c_105_p N_VPWR_c_302_n 0.00485263f $X=2.66 $Y=2.1 $X2=0 $Y2=0
cc_116 N_A_84_28#_c_106_p N_VPWR_c_302_n 0.0249852f $X=2.63 $Y=2.435 $X2=0 $Y2=0
cc_117 N_A_84_28#_M1008_g N_VPWR_c_303_n 0.00486043f $X=0.695 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_84_28#_c_106_p N_VPWR_c_306_n 0.0167395f $X=2.63 $Y=2.435 $X2=0 $Y2=0
cc_119 N_A_84_28#_M1001_d N_VPWR_c_298_n 0.00430974f $X=2.47 $Y=1.835 $X2=0
+ $Y2=0
cc_120 N_A_84_28#_M1008_g N_VPWR_c_298_n 0.00933203f $X=0.695 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_A_84_28#_c_106_p N_VPWR_c_298_n 0.0102309f $X=2.63 $Y=2.435 $X2=0 $Y2=0
cc_122 N_A_84_28#_c_69_n N_VGND_M1005_d 0.0018166f $X=0.85 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_84_28#_c_81_p N_VGND_M1005_d 0.0147588f $X=1.135 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_84_28#_c_135_p N_VGND_M1005_d 0.00611744f $X=0.935 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_84_28#_c_70_n N_VGND_M1005_d 0.00286001f $X=1.22 $Y=0.87 $X2=-0.19
+ $Y2=-0.245
cc_126 N_A_84_28#_c_67_n N_VGND_c_343_n 0.0126696f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_127 N_A_84_28#_c_135_p N_VGND_c_343_n 0.0128082f $X=0.935 $Y=0.955 $X2=0
+ $Y2=0
cc_128 N_A_84_28#_c_70_n N_VGND_c_343_n 0.0182686f $X=1.22 $Y=0.87 $X2=0 $Y2=0
cc_129 N_A_84_28#_c_72_n N_VGND_c_343_n 0.0126224f $X=1.305 $Y=0.34 $X2=0 $Y2=0
cc_130 N_A_84_28#_c_74_n N_VGND_c_343_n 0.00578976f $X=0.85 $Y=1.385 $X2=0 $Y2=0
cc_131 N_A_84_28#_c_75_n N_VGND_c_343_n 0.00394744f $X=0.695 $Y=1.385 $X2=0
+ $Y2=0
cc_132 N_A_84_28#_c_67_n N_VGND_c_345_n 0.00493667f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A_84_28#_c_71_n N_VGND_c_346_n 0.0644106f $X=2.075 $Y=0.34 $X2=0 $Y2=0
cc_134 N_A_84_28#_c_72_n N_VGND_c_346_n 0.0121867f $X=1.305 $Y=0.34 $X2=0 $Y2=0
cc_135 N_A_84_28#_c_67_n N_VGND_c_348_n 0.00956483f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_136 N_A_84_28#_c_71_n N_VGND_c_348_n 0.0380785f $X=2.075 $Y=0.34 $X2=0 $Y2=0
cc_137 N_A_84_28#_c_72_n N_VGND_c_348_n 0.00660921f $X=1.305 $Y=0.34 $X2=0 $Y2=0
cc_138 N_A_84_28#_c_73_n N_A_494_51#_c_388_n 0.00940701f $X=2.18 $Y=0.43 $X2=0
+ $Y2=0
cc_139 B1_N N_A_281_138#_c_185_n 2.6616e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B1_N_c_152_n N_A_281_138#_c_185_n 0.017311f $X=1.22 $Y=1.385 $X2=0
+ $Y2=0
cc_141 B1_N N_A_281_138#_c_187_n 0.0414514f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_142 N_B1_N_c_153_n N_A_281_138#_c_187_n 0.00715166f $X=1.23 $Y=1.22 $X2=0
+ $Y2=0
cc_143 N_B1_N_M1000_g N_A_281_138#_c_188_n 0.00715166f $X=1.33 $Y=2.045 $X2=0
+ $Y2=0
cc_144 N_B1_N_c_152_n N_A_281_138#_c_189_n 0.00715166f $X=1.22 $Y=1.385 $X2=0
+ $Y2=0
cc_145 N_B1_N_M1000_g N_VPWR_c_299_n 0.00690562f $X=1.33 $Y=2.045 $X2=0 $Y2=0
cc_146 B1_N N_VPWR_c_299_n 0.0106179f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_147 N_B1_N_c_152_n N_VPWR_c_299_n 0.00244497f $X=1.22 $Y=1.385 $X2=0 $Y2=0
cc_148 N_B1_N_M1000_g N_VPWR_c_300_n 0.00270314f $X=1.33 $Y=2.045 $X2=0 $Y2=0
cc_149 N_B1_N_c_153_n N_VGND_c_343_n 4.98627e-19 $X=1.23 $Y=1.22 $X2=0 $Y2=0
cc_150 N_B1_N_c_153_n N_VGND_c_346_n 2.50133e-19 $X=1.23 $Y=1.22 $X2=0 $Y2=0
cc_151 N_A_281_138#_c_183_n N_A2_M1007_g 0.0226504f $X=2.395 $Y=1.22 $X2=0 $Y2=0
cc_152 N_A_281_138#_M1001_g N_A2_M1003_g 0.016785f $X=2.395 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_281_138#_c_186_n A2 0.00295634f $X=2.395 $Y=1.385 $X2=0 $Y2=0
cc_154 N_A_281_138#_c_186_n N_A2_c_222_n 0.0181687f $X=2.395 $Y=1.385 $X2=0
+ $Y2=0
cc_155 N_A_281_138#_M1001_g N_VPWR_c_300_n 0.0185741f $X=2.395 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_281_138#_M1001_g N_VPWR_c_306_n 0.00486043f $X=2.395 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_281_138#_M1001_g N_VPWR_c_298_n 0.0083203f $X=2.395 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A_281_138#_c_183_n N_VGND_c_346_n 0.00565115f $X=2.395 $Y=1.22 $X2=0
+ $Y2=0
cc_159 N_A_281_138#_c_183_n N_VGND_c_348_n 0.0119838f $X=2.395 $Y=1.22 $X2=0
+ $Y2=0
cc_160 N_A_281_138#_c_183_n N_A_494_51#_c_388_n 9.73274e-19 $X=2.395 $Y=1.22
+ $X2=0 $Y2=0
cc_161 N_A2_M1007_g N_A1_M1009_g 0.0251886f $X=2.825 $Y=0.675 $X2=0 $Y2=0
cc_162 N_A2_M1003_g N_A1_M1004_g 0.0493825f $X=2.845 $Y=2.465 $X2=0 $Y2=0
cc_163 A2 N_A1_c_257_n 0.0026909f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A2_c_222_n N_A1_c_257_n 0.018139f $X=2.875 $Y=1.51 $X2=0 $Y2=0
cc_165 A2 N_A1_c_258_n 0.0274126f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_166 N_A2_c_222_n N_A1_c_258_n 4.79693e-19 $X=2.875 $Y=1.51 $X2=0 $Y2=0
cc_167 N_A2_M1003_g N_VPWR_c_300_n 0.00132953f $X=2.845 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A2_M1003_g N_VPWR_c_302_n 0.00458595f $X=2.845 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A2_M1003_g N_VPWR_c_306_n 0.0054895f $X=2.845 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A2_M1003_g N_VPWR_c_298_n 0.0103157f $X=2.845 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A2_M1007_g N_VGND_c_344_n 0.00330325f $X=2.825 $Y=0.675 $X2=0 $Y2=0
cc_172 N_A2_M1007_g N_VGND_c_346_n 0.00565115f $X=2.825 $Y=0.675 $X2=0 $Y2=0
cc_173 N_A2_M1007_g N_VGND_c_348_n 0.0107556f $X=2.825 $Y=0.675 $X2=0 $Y2=0
cc_174 N_A2_M1007_g N_A_494_51#_c_387_n 0.014861f $X=2.825 $Y=0.675 $X2=0 $Y2=0
cc_175 A2 N_A_494_51#_c_387_n 0.0310725f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A2_c_222_n N_A_494_51#_c_387_n 0.00425107f $X=2.875 $Y=1.51 $X2=0 $Y2=0
cc_177 A2 N_A_494_51#_c_388_n 0.0173f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A2_M1007_g N_A_494_51#_c_389_n 6.59263e-19 $X=2.825 $Y=0.675 $X2=0
+ $Y2=0
cc_179 N_A1_M1004_g N_VPWR_c_302_n 0.0320364f $X=3.355 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A1_c_257_n N_VPWR_c_302_n 0.00152318f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_181 N_A1_c_258_n N_VPWR_c_302_n 0.0261279f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_182 N_A1_M1004_g N_VPWR_c_306_n 0.00486043f $X=3.355 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A1_M1004_g N_VPWR_c_298_n 0.0085771f $X=3.355 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A1_M1009_g N_VGND_c_344_n 0.00646956f $X=3.355 $Y=0.675 $X2=0 $Y2=0
cc_185 N_A1_M1009_g N_VGND_c_347_n 0.00529818f $X=3.355 $Y=0.675 $X2=0 $Y2=0
cc_186 N_A1_M1009_g N_VGND_c_348_n 0.0108215f $X=3.355 $Y=0.675 $X2=0 $Y2=0
cc_187 N_A1_M1009_g N_A_494_51#_c_387_n 0.0178197f $X=3.355 $Y=0.675 $X2=0 $Y2=0
cc_188 N_A1_c_257_n N_A_494_51#_c_387_n 0.00731208f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_189 N_A1_c_258_n N_A_494_51#_c_387_n 0.0295243f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_190 N_A1_M1009_g N_A_494_51#_c_389_n 0.013029f $X=3.355 $Y=0.675 $X2=0 $Y2=0
cc_191 X N_VPWR_c_303_n 0.034299f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_192 N_X_M1008_s N_VPWR_c_298_n 0.00371702f $X=0.355 $Y=1.835 $X2=0 $Y2=0
cc_193 X N_VPWR_c_298_n 0.0189723f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_194 N_X_c_281_n N_VGND_c_343_n 0.0174954f $X=0.28 $Y=0.42 $X2=0 $Y2=0
cc_195 N_X_c_281_n N_VGND_c_345_n 0.0213627f $X=0.28 $Y=0.42 $X2=0 $Y2=0
cc_196 N_X_c_281_n N_VGND_c_348_n 0.0115856f $X=0.28 $Y=0.42 $X2=0 $Y2=0
cc_197 N_VPWR_c_298_n A_584_367# 0.0154185f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_198 N_VGND_c_346_n N_A_494_51#_c_386_n 0.0140491f $X=2.905 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_348_n N_A_494_51#_c_386_n 0.0090585f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_200 N_VGND_M1007_d N_A_494_51#_c_387_n 0.00289294f $X=2.9 $Y=0.255 $X2=0
+ $Y2=0
cc_201 N_VGND_c_344_n N_A_494_51#_c_387_n 0.0216414f $X=3.07 $Y=0.4 $X2=0 $Y2=0
cc_202 N_VGND_c_347_n N_A_494_51#_c_389_n 0.0210467f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_c_348_n N_A_494_51#_c_389_n 0.0126321f $X=3.6 $Y=0 $X2=0 $Y2=0
