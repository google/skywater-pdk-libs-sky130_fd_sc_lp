* File: sky130_fd_sc_lp__dlxbn_2.spice
* Created: Fri Aug 28 10:27:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxbn_2.pex.spice"
.subckt sky130_fd_sc_lp__dlxbn_2  VNB VPB D GATE_N VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_D_M1014_g N_A_45_136#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1013 N_A_214_136#_M1013_d N_GATE_N_M1013_g N_VGND_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_214_136#_M1010_g N_A_354_47#_M1010_s VNB NSHORT L=0.15
+ W=0.42 AD=0.08775 AS=0.1113 PD=0.85 PS=1.37 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1001 A_547_47# N_A_45_136#_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.08775 PD=0.63 PS=0.85 NRD=14.28 NRS=17.136 M=1 R=2.8 SA=75000.7
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1022 N_A_619_47#_M1022_d N_A_214_136#_M1022_g A_547_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.09385 AS=0.0441 PD=0.87 PS=0.63 NRD=22.848 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1002 A_737_47# N_A_354_47#_M1002_g N_A_619_47#_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0714 AS=0.09385 PD=0.76 PS=0.87 NRD=32.856 NRS=22.848 M=1 R=2.8
+ SA=75001.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_805_21#_M1017_g A_737_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.138033 AS=0.0714 PD=0.973333 PS=0.76 NRD=32.856 NRS=32.856 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1012 N_A_805_21#_M1012_d N_A_619_47#_M1012_g N_VGND_M1017_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.276067 PD=2.25 PS=1.94667 NRD=0 NRS=16.776 M=1 R=5.6
+ SA=75001.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1018 N_VGND_M1018_d N_A_805_21#_M1018_g N_A_1138_153#_M1018_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.138733 AS=0.1197 PD=0.976667 PS=1.41 NRD=78.66 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1018_d N_A_1138_153#_M1007_g N_Q_N_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.277467 AS=0.1176 PD=1.95333 PS=1.12 NRD=17.136 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1024_d N_A_1138_153#_M1024_g N_Q_N_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.20075 AS=0.1176 PD=1.39 PS=1.12 NRD=12.132 NRS=0 M=1 R=5.6
+ SA=75001 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1008 N_Q_M1008_d N_A_805_21#_M1008_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6 SA=75001.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1025 N_Q_M1008_d N_A_805_21#_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1011 N_VPWR_M1011_d N_D_M1011_g N_A_45_136#_M1011_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.2048 PD=0.92 PS=1.92 NRD=0 NRS=16.9223 M=1 R=4.26667 SA=75000.2
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1019 N_A_214_136#_M1019_d N_GATE_N_M1019_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.3459 AS=0.0896 PD=2.7 PS=0.92 NRD=149.424 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_214_136#_M1000_g N_A_354_47#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1696 PD=1.21 PS=1.81 NRD=43.0839 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1023 A_589_491# N_A_45_136#_M1023_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.21 NRD=15.3857 NRS=46.1571 M=1 R=4.26667
+ SA=75000.9 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_619_47#_M1020_d N_A_354_47#_M1020_g A_589_491# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.134098 AS=0.0672 PD=1.24377 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.3 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1006 A_769_491# N_A_214_136#_M1006_g N_A_619_47#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0880019 PD=0.63 PS=0.816226 NRD=23.443 NRS=52.7566 M=1
+ R=2.8 SA=75001.8 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_805_21#_M1005_g A_769_491# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.120025 AS=0.0441 PD=0.9325 PS=0.63 NRD=77.3816 NRS=23.443 M=1 R=2.8
+ SA=75002.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1016 N_A_805_21#_M1016_d N_A_619_47#_M1016_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.360075 PD=3.05 PS=2.7975 NRD=0 NRS=16.9223 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_805_21#_M1009_g N_A_1138_153#_M1009_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.17472 AS=0.1696 PD=1.19579 PS=1.81 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1009_d N_A_1138_153#_M1003_g N_Q_N_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.34398 AS=0.1764 PD=2.35421 PS=1.54 NRD=18.3604 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1015 N_VPWR_M1015_d N_A_1138_153#_M1015_g N_Q_N_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75001 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_Q_M1004_d N_A_805_21#_M1004_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2268 PD=1.54 PS=1.62 NRD=0 NRS=1.5563 M=1 R=8.4 SA=75001.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1021 N_Q_M1004_d N_A_805_21#_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=17.0653 P=21.91
*
.include "sky130_fd_sc_lp__dlxbn_2.pxi.spice"
*
.ends
*
*
