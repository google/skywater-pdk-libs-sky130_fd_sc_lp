* NGSPICE file created from sky130_fd_sc_lp__dfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
M1000 a_423_191# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.7428e+12p ps=1.451e+07u
M1001 VPWR a_1440_304# a_1398_472# VPB phighvt w=420000u l=150000u
+  ad=1.8202e+12p pd=1.66e+07u as=8.82e+10p ps=1.26e+06u
M1002 a_1398_472# a_197_108# a_1245_128# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.43e+06u
M1003 a_603_191# a_28_108# a_304_463# VNB nshort w=420000u l=150000u
+  ad=2.709e+11p pd=2.13e+06u as=1.638e+11p ps=1.62e+06u
M1004 VPWR a_1796_139# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1005 a_1420_128# a_28_108# a_1245_128# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=4.398e+11p ps=2.73e+06u
M1006 VPWR a_1245_128# a_1440_304# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1007 Q a_1796_139# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1008 Q_N a_1245_128# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1009 VPWR a_804_328# a_789_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 a_848_191# a_804_328# a_762_191# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=1.176e+11p ps=1.4e+06u
M1011 a_789_463# a_28_108# a_603_191# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.289e+11p ps=2.77e+06u
M1012 VPWR CLK a_28_108# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1013 a_304_463# D VPWR VPB phighvt w=420000u l=150000u
+  ad=3.465e+11p pd=4.17e+06u as=0p ps=0u
M1014 a_197_108# a_28_108# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1015 a_603_191# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1440_304# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1578_128# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1018 a_603_191# a_197_108# a_304_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_762_191# a_197_108# a_603_191# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_804_328# a_603_191# VGND VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1021 a_1245_128# a_197_108# a_804_328# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_304_463# D a_423_191# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q_N a_1245_128# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1024 a_1440_304# a_1245_128# a_1578_128# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1025 VPWR RESET_B a_304_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND RESET_B a_848_191# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND CLK a_28_108# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1028 a_197_108# a_28_108# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1029 a_1245_128# a_28_108# a_804_328# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=4.6965e+11p ps=3.03e+06u
M1030 VPWR a_1245_128# a_1796_139# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1031 VGND a_1245_128# a_1796_139# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.883e+11p ps=1.78e+06u
M1032 a_804_328# a_603_191# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_1440_304# a_1420_128# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

