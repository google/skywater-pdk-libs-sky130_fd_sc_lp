* File: sky130_fd_sc_lp__or4_4.pxi.spice
* Created: Fri Aug 28 11:25:10 2020
* 
x_PM_SKY130_FD_SC_LP__OR4_4%D N_D_c_87_n N_D_M1004_g N_D_M1000_g N_D_c_89_n
+ N_D_c_90_n D D PM_SKY130_FD_SC_LP__OR4_4%D
x_PM_SKY130_FD_SC_LP__OR4_4%C N_C_M1012_g N_C_M1009_g C C N_C_c_117_n
+ PM_SKY130_FD_SC_LP__OR4_4%C
x_PM_SKY130_FD_SC_LP__OR4_4%B N_B_M1002_g N_B_M1007_g B N_B_c_154_n N_B_c_155_n
+ PM_SKY130_FD_SC_LP__OR4_4%B
x_PM_SKY130_FD_SC_LP__OR4_4%A N_A_M1013_g N_A_M1008_g A N_A_c_188_n N_A_c_189_n
+ PM_SKY130_FD_SC_LP__OR4_4%A
x_PM_SKY130_FD_SC_LP__OR4_4%A_58_367# N_A_58_367#_M1004_d N_A_58_367#_M1007_d
+ N_A_58_367#_M1000_s N_A_58_367#_M1005_g N_A_58_367#_M1001_g
+ N_A_58_367#_M1011_g N_A_58_367#_M1003_g N_A_58_367#_M1014_g
+ N_A_58_367#_M1006_g N_A_58_367#_M1015_g N_A_58_367#_M1010_g
+ N_A_58_367#_c_244_n N_A_58_367#_c_245_n N_A_58_367#_c_252_n
+ N_A_58_367#_c_258_n N_A_58_367#_c_231_n N_A_58_367#_c_232_n
+ N_A_58_367#_c_265_n N_A_58_367#_c_233_n N_A_58_367#_c_234_n
+ N_A_58_367#_c_235_n N_A_58_367#_c_236_n N_A_58_367#_c_237_n
+ N_A_58_367#_c_238_n N_A_58_367#_c_239_n PM_SKY130_FD_SC_LP__OR4_4%A_58_367#
x_PM_SKY130_FD_SC_LP__OR4_4%VPWR N_VPWR_M1008_d N_VPWR_M1003_d N_VPWR_M1010_d
+ N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_390_n
+ N_VPWR_c_391_n N_VPWR_c_392_n VPWR N_VPWR_c_393_n N_VPWR_c_394_n
+ N_VPWR_c_385_n N_VPWR_c_396_n PM_SKY130_FD_SC_LP__OR4_4%VPWR
x_PM_SKY130_FD_SC_LP__OR4_4%X N_X_M1005_s N_X_M1014_s N_X_M1001_s N_X_M1006_s
+ N_X_c_498_p N_X_c_486_n N_X_c_440_n N_X_c_441_n N_X_c_447_n N_X_c_448_n
+ N_X_c_495_p N_X_c_490_n N_X_c_449_n N_X_c_442_n N_X_c_443_n N_X_c_450_n X X X
+ X X PM_SKY130_FD_SC_LP__OR4_4%X
x_PM_SKY130_FD_SC_LP__OR4_4%VGND N_VGND_M1004_s N_VGND_M1009_d N_VGND_M1013_d
+ N_VGND_M1011_d N_VGND_M1015_d N_VGND_c_505_n N_VGND_c_506_n N_VGND_c_507_n
+ N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n N_VGND_c_511_n N_VGND_c_512_n
+ N_VGND_c_513_n N_VGND_c_514_n N_VGND_c_515_n N_VGND_c_516_n VGND
+ N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n
+ PM_SKY130_FD_SC_LP__OR4_4%VGND
cc_1 VNB N_D_c_87_n 0.022658f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.21
cc_2 VNB N_D_M1000_g 0.00543551f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.465
cc_3 VNB N_D_c_89_n 0.0411225f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.375
cc_4 VNB N_D_c_90_n 0.010462f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.375
cc_5 VNB D 0.0259435f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_C_M1009_g 0.0258602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB C 0.00572903f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_C_c_117_n 0.0227321f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_9 VNB N_B_M1007_g 0.0258648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_154_n 0.0242072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_155_n 0.00361559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_M1013_g 0.0257061f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.665
cc_13 VNB N_A_c_188_n 0.0264005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_c_189_n 0.00103489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_58_367#_M1005_g 0.0246677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_58_367#_M1011_g 0.0221884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_58_367#_M1014_g 0.022195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_58_367#_M1015_g 0.02842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_58_367#_c_231_n 0.0071123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_58_367#_c_232_n 0.00329865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_58_367#_c_233_n 0.00494517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_58_367#_c_234_n 0.00233717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_58_367#_c_235_n 3.45182e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_58_367#_c_236_n 0.0015776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_58_367#_c_237_n 0.0805522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_58_367#_c_238_n 0.00761983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_58_367#_c_239_n 0.0010166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_385_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_440_n 0.0086357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_441_n 0.00270104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_442_n 0.0131919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_443_n 0.00177012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB X 0.0355993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.00973053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB X 0.0222482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_505_n 0.0153857f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_37 VNB N_VGND_c_506_n 0.0340321f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_38 VNB N_VGND_c_507_n 0.0158122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_508_n 0.00474659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_509_n 0.00473997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_510_n 5.00305e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_511_n 0.0148369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_512_n 0.0175141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_513_n 0.017949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_514_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_515_n 0.0164391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_516_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_517_n 0.0169395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_518_n 0.262847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_519_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_520_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_D_M1000_g 0.023939f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_53 VPB D 0.0135036f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_54 VPB N_C_M1012_g 0.0187037f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.665
cc_55 VPB C 0.00499702f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_56 VPB N_C_c_117_n 0.00624994f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.375
cc_57 VPB N_B_M1002_g 0.0211328f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.665
cc_58 VPB N_B_c_154_n 0.00637553f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_B_c_155_n 0.00272262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_M1008_g 0.0213955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_c_188_n 0.00632004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_c_189_n 0.00157004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_58_367#_M1001_g 0.0195477f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.375
cc_64 VPB N_A_58_367#_M1003_g 0.0179231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_58_367#_M1006_g 0.0179297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_58_367#_M1010_g 0.0217531f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_58_367#_c_244_n 0.00745115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_58_367#_c_245_n 0.0379885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_58_367#_c_235_n 0.00144307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_58_367#_c_237_n 0.0171528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_386_n 0.00501995f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_387_n 3.22457e-19 $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.375
cc_73 VPB N_VPWR_c_388_n 0.0412021f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.665
cc_74 VPB N_VPWR_c_389_n 0.0684612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_390_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_391_n 0.0165323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_392_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_393_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_394_n 0.017577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_385_n 0.0670347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_396_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_X_c_447_n 0.00304538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_X_c_448_n 0.00195054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_X_c_449_n 0.0296689f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_X_c_450_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB X 0.00642948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 N_D_M1000_g N_C_M1012_g 0.059852f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_88 N_D_c_87_n N_C_M1009_g 0.0241685f $X=0.63 $Y=1.21 $X2=0 $Y2=0
cc_89 D N_C_M1009_g 5.24962e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_90 N_D_M1000_g C 0.00623353f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_91 N_D_c_90_n C 0.00738079f $X=0.63 $Y=1.375 $X2=0 $Y2=0
cc_92 D C 0.0277311f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_93 N_D_c_90_n N_C_c_117_n 0.059852f $X=0.63 $Y=1.375 $X2=0 $Y2=0
cc_94 D N_C_c_117_n 4.04893e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_95 N_D_M1000_g N_A_58_367#_c_244_n 0.00163016f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_96 N_D_c_89_n N_A_58_367#_c_244_n 0.00342614f $X=0.555 $Y=1.375 $X2=0 $Y2=0
cc_97 D N_A_58_367#_c_244_n 0.0185242f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_98 N_D_M1000_g N_A_58_367#_c_245_n 0.0197753f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_99 N_D_M1000_g N_A_58_367#_c_252_n 0.0119921f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_100 N_D_c_87_n N_A_58_367#_c_232_n 0.00253514f $X=0.63 $Y=1.21 $X2=0 $Y2=0
cc_101 N_D_M1000_g N_VPWR_c_389_n 0.0054895f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_102 N_D_M1000_g N_VPWR_c_385_n 0.0109026f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_103 N_D_c_87_n N_VGND_c_506_n 0.0172566f $X=0.63 $Y=1.21 $X2=0 $Y2=0
cc_104 N_D_c_89_n N_VGND_c_506_n 0.00469603f $X=0.555 $Y=1.375 $X2=0 $Y2=0
cc_105 D N_VGND_c_506_n 0.0175384f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_106 N_D_c_87_n N_VGND_c_507_n 0.00477554f $X=0.63 $Y=1.21 $X2=0 $Y2=0
cc_107 N_D_c_87_n N_VGND_c_518_n 0.00828349f $X=0.63 $Y=1.21 $X2=0 $Y2=0
cc_108 N_C_M1012_g N_B_M1002_g 0.0553412f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_109 N_C_M1009_g N_B_M1007_g 0.0291164f $X=1.06 $Y=0.665 $X2=0 $Y2=0
cc_110 C N_B_c_154_n 0.00232612f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_C_c_117_n N_B_c_154_n 0.0209912f $X=1.08 $Y=1.51 $X2=0 $Y2=0
cc_112 C N_B_c_155_n 0.0281403f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_113 N_C_c_117_n N_B_c_155_n 7.72092e-19 $X=1.08 $Y=1.51 $X2=0 $Y2=0
cc_114 N_C_M1012_g N_A_58_367#_c_245_n 0.0048871f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_115 N_C_M1012_g N_A_58_367#_c_252_n 0.0150921f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_116 C N_A_58_367#_c_252_n 0.0469164f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_117 N_C_c_117_n N_A_58_367#_c_252_n 9.05333e-19 $X=1.08 $Y=1.51 $X2=0 $Y2=0
cc_118 N_C_M1009_g N_A_58_367#_c_258_n 0.0108095f $X=1.06 $Y=0.665 $X2=0 $Y2=0
cc_119 N_C_M1009_g N_A_58_367#_c_231_n 0.0122728f $X=1.06 $Y=0.665 $X2=0 $Y2=0
cc_120 C N_A_58_367#_c_231_n 0.0170899f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_121 N_C_c_117_n N_A_58_367#_c_231_n 0.00254934f $X=1.08 $Y=1.51 $X2=0 $Y2=0
cc_122 N_C_M1009_g N_A_58_367#_c_232_n 0.00157969f $X=1.06 $Y=0.665 $X2=0 $Y2=0
cc_123 C N_A_58_367#_c_232_n 0.0165798f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_124 N_C_c_117_n N_A_58_367#_c_232_n 0.00198375f $X=1.08 $Y=1.51 $X2=0 $Y2=0
cc_125 N_C_M1009_g N_A_58_367#_c_265_n 8.80337e-19 $X=1.06 $Y=0.665 $X2=0 $Y2=0
cc_126 N_C_M1012_g N_VPWR_c_389_n 0.00585385f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_127 N_C_M1012_g N_VPWR_c_385_n 0.011101f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_128 N_C_M1009_g N_VGND_c_506_n 7.42749e-19 $X=1.06 $Y=0.665 $X2=0 $Y2=0
cc_129 N_C_M1009_g N_VGND_c_507_n 0.00539298f $X=1.06 $Y=0.665 $X2=0 $Y2=0
cc_130 N_C_M1009_g N_VGND_c_508_n 0.00518195f $X=1.06 $Y=0.665 $X2=0 $Y2=0
cc_131 N_C_M1009_g N_VGND_c_518_n 0.0102217f $X=1.06 $Y=0.665 $X2=0 $Y2=0
cc_132 N_B_M1007_g N_A_M1013_g 0.02734f $X=1.64 $Y=0.665 $X2=0 $Y2=0
cc_133 N_B_M1002_g N_A_M1008_g 0.0515392f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B_c_154_n N_A_c_188_n 0.0206141f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_135 N_B_c_155_n N_A_c_188_n 0.00247975f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_136 N_B_c_154_n N_A_c_189_n 3.74634e-19 $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_137 N_B_c_155_n N_A_c_189_n 0.0322427f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_138 N_B_M1002_g N_A_58_367#_c_252_n 0.0172852f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_139 N_B_c_154_n N_A_58_367#_c_252_n 9.01154e-19 $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_140 N_B_c_155_n N_A_58_367#_c_252_n 0.0237646f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_141 N_B_M1007_g N_A_58_367#_c_258_n 8.89265e-19 $X=1.64 $Y=0.665 $X2=0 $Y2=0
cc_142 N_B_M1007_g N_A_58_367#_c_231_n 0.0118846f $X=1.64 $Y=0.665 $X2=0 $Y2=0
cc_143 N_B_c_154_n N_A_58_367#_c_231_n 0.0021576f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_144 N_B_c_155_n N_A_58_367#_c_231_n 0.0137749f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_145 N_B_M1007_g N_A_58_367#_c_265_n 0.0116603f $X=1.64 $Y=0.665 $X2=0 $Y2=0
cc_146 N_B_M1007_g N_A_58_367#_c_238_n 0.00168563f $X=1.64 $Y=0.665 $X2=0 $Y2=0
cc_147 N_B_c_154_n N_A_58_367#_c_238_n 5.49911e-19 $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_148 N_B_c_155_n N_A_58_367#_c_238_n 0.0115342f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_149 N_B_M1002_g N_VPWR_c_389_n 0.00585385f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_150 N_B_M1002_g N_VPWR_c_385_n 0.011557f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_151 N_B_M1007_g N_VGND_c_508_n 0.00536995f $X=1.64 $Y=0.665 $X2=0 $Y2=0
cc_152 N_B_M1007_g N_VGND_c_513_n 0.00539298f $X=1.64 $Y=0.665 $X2=0 $Y2=0
cc_153 N_B_M1007_g N_VGND_c_518_n 0.0101944f $X=1.64 $Y=0.665 $X2=0 $Y2=0
cc_154 N_A_M1013_g N_A_58_367#_M1005_g 0.0275237f $X=2.07 $Y=0.665 $X2=0 $Y2=0
cc_155 N_A_M1008_g N_A_58_367#_M1001_g 0.0349795f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A_c_189_n N_A_58_367#_M1001_g 2.26172e-19 $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A_M1008_g N_A_58_367#_c_252_n 0.0163762f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_c_188_n N_A_58_367#_c_252_n 0.0029438f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A_c_189_n N_A_58_367#_c_252_n 0.0171481f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A_M1013_g N_A_58_367#_c_265_n 0.0116441f $X=2.07 $Y=0.665 $X2=0 $Y2=0
cc_161 N_A_M1013_g N_A_58_367#_c_233_n 0.0118485f $X=2.07 $Y=0.665 $X2=0 $Y2=0
cc_162 N_A_c_188_n N_A_58_367#_c_233_n 0.00339745f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_163 N_A_c_189_n N_A_58_367#_c_233_n 0.016719f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A_M1013_g N_A_58_367#_c_234_n 0.0034595f $X=2.07 $Y=0.665 $X2=0 $Y2=0
cc_165 N_A_c_188_n N_A_58_367#_c_234_n 5.26016e-19 $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_166 N_A_c_189_n N_A_58_367#_c_234_n 0.00585807f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_167 N_A_M1008_g N_A_58_367#_c_235_n 0.00350021f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A_c_188_n N_A_58_367#_c_235_n 5.26016e-19 $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A_c_189_n N_A_58_367#_c_235_n 0.0124608f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A_c_188_n N_A_58_367#_c_237_n 0.0168326f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_171 N_A_c_189_n N_A_58_367#_c_237_n 2.91526e-19 $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_172 N_A_M1013_g N_A_58_367#_c_238_n 0.00190778f $X=2.07 $Y=0.665 $X2=0 $Y2=0
cc_173 N_A_c_189_n N_A_58_367#_c_238_n 0.00147988f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_174 N_A_c_188_n N_A_58_367#_c_239_n 0.00129183f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_175 N_A_c_189_n N_A_58_367#_c_239_n 0.014087f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A_M1008_g N_VPWR_c_386_n 0.00830791f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A_M1008_g N_VPWR_c_389_n 0.00585385f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_M1008_g N_VPWR_c_385_n 0.0114683f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A_M1013_g N_VGND_c_509_n 0.00532898f $X=2.07 $Y=0.665 $X2=0 $Y2=0
cc_180 N_A_M1013_g N_VGND_c_513_n 0.00539298f $X=2.07 $Y=0.665 $X2=0 $Y2=0
cc_181 N_A_M1013_g N_VGND_c_518_n 0.0101851f $X=2.07 $Y=0.665 $X2=0 $Y2=0
cc_182 N_A_58_367#_c_252_n A_141_367# 0.00468592f $X=2.425 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_58_367#_c_252_n A_213_367# 0.0155103f $X=2.425 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_58_367#_c_252_n A_321_367# 0.0164968f $X=2.425 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_58_367#_c_252_n N_VPWR_M1008_d 0.00903103f $X=2.425 $Y=2.015
+ $X2=-0.19 $Y2=-0.245
cc_186 N_A_58_367#_c_235_n N_VPWR_M1008_d 0.00118786f $X=2.51 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_58_367#_M1001_g N_VPWR_c_386_n 0.00664393f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_58_367#_c_252_n N_VPWR_c_386_n 0.0259956f $X=2.425 $Y=2.015 $X2=0
+ $Y2=0
cc_189 N_A_58_367#_M1001_g N_VPWR_c_387_n 7.56381e-19 $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A_58_367#_M1003_g N_VPWR_c_387_n 0.0143579f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A_58_367#_M1006_g N_VPWR_c_387_n 0.0141781f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_192 N_A_58_367#_M1010_g N_VPWR_c_387_n 7.24342e-19 $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_A_58_367#_M1006_g N_VPWR_c_388_n 7.24342e-19 $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_A_58_367#_M1010_g N_VPWR_c_388_n 0.0152828f $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_58_367#_c_245_n N_VPWR_c_389_n 0.0210467f $X=0.415 $Y=2.95 $X2=0
+ $Y2=0
cc_196 N_A_58_367#_M1001_g N_VPWR_c_391_n 0.00585385f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_A_58_367#_M1003_g N_VPWR_c_391_n 0.00486043f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A_58_367#_M1006_g N_VPWR_c_393_n 0.00486043f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A_58_367#_M1010_g N_VPWR_c_393_n 0.00486043f $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_200 N_A_58_367#_M1000_s N_VPWR_c_385_n 0.00215158f $X=0.29 $Y=1.835 $X2=0
+ $Y2=0
cc_201 N_A_58_367#_M1001_g N_VPWR_c_385_n 0.0111134f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_202 N_A_58_367#_M1003_g N_VPWR_c_385_n 0.00824727f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_203 N_A_58_367#_M1006_g N_VPWR_c_385_n 0.00824727f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_A_58_367#_M1010_g N_VPWR_c_385_n 0.00824727f $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_205 N_A_58_367#_c_245_n N_VPWR_c_385_n 0.0125689f $X=0.415 $Y=2.95 $X2=0
+ $Y2=0
cc_206 N_A_58_367#_M1011_g N_X_c_440_n 0.0138902f $X=3.075 $Y=0.665 $X2=0 $Y2=0
cc_207 N_A_58_367#_M1014_g N_X_c_440_n 0.0142932f $X=3.505 $Y=0.665 $X2=0 $Y2=0
cc_208 N_A_58_367#_c_236_n N_X_c_440_n 0.0467265f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_209 N_A_58_367#_c_237_n N_X_c_440_n 0.00246472f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_210 N_A_58_367#_M1005_g N_X_c_441_n 0.00139667f $X=2.645 $Y=0.665 $X2=0 $Y2=0
cc_211 N_A_58_367#_c_233_n N_X_c_441_n 0.00708451f $X=2.425 $Y=1.08 $X2=0 $Y2=0
cc_212 N_A_58_367#_c_234_n N_X_c_441_n 0.00722632f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_213 N_A_58_367#_c_236_n N_X_c_441_n 0.0153308f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_214 N_A_58_367#_c_237_n N_X_c_441_n 0.00256759f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_215 N_A_58_367#_M1003_g N_X_c_447_n 0.0129099f $X=3.075 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A_58_367#_M1006_g N_X_c_447_n 0.0130453f $X=3.505 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_58_367#_c_236_n N_X_c_447_n 0.0467265f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_218 N_A_58_367#_c_237_n N_X_c_447_n 0.00246472f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_219 N_A_58_367#_M1001_g N_X_c_448_n 5.73473e-19 $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A_58_367#_c_235_n N_X_c_448_n 0.00880114f $X=2.51 $Y=1.93 $X2=0 $Y2=0
cc_221 N_A_58_367#_c_236_n N_X_c_448_n 0.0153308f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_222 N_A_58_367#_c_237_n N_X_c_448_n 0.00256759f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_223 N_A_58_367#_M1010_g N_X_c_449_n 0.0150864f $X=3.935 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_58_367#_c_236_n N_X_c_449_n 0.0312279f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_225 N_A_58_367#_c_237_n N_X_c_449_n 0.0061618f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_226 N_A_58_367#_M1015_g N_X_c_442_n 0.0170683f $X=3.935 $Y=0.665 $X2=0 $Y2=0
cc_227 N_A_58_367#_c_236_n N_X_c_442_n 0.028724f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A_58_367#_c_237_n N_X_c_442_n 0.0061618f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_229 N_A_58_367#_c_236_n N_X_c_443_n 0.0181554f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_230 N_A_58_367#_c_237_n N_X_c_443_n 0.00256759f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_231 N_A_58_367#_c_236_n N_X_c_450_n 0.0153308f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_232 N_A_58_367#_c_237_n N_X_c_450_n 0.00256759f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_233 N_A_58_367#_M1015_g X 0.00317266f $X=3.935 $Y=0.665 $X2=0 $Y2=0
cc_234 N_A_58_367#_M1015_g X 0.00248935f $X=3.935 $Y=0.665 $X2=0 $Y2=0
cc_235 N_A_58_367#_M1010_g X 0.00248935f $X=3.935 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A_58_367#_c_236_n X 0.0139437f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_237 N_A_58_367#_c_237_n X 0.00829366f $X=4.095 $Y=1.51 $X2=0 $Y2=0
cc_238 N_A_58_367#_c_231_n N_VGND_M1009_d 0.00370397f $X=1.69 $Y=1.08 $X2=0
+ $Y2=0
cc_239 N_A_58_367#_c_233_n N_VGND_M1013_d 0.00365393f $X=2.425 $Y=1.08 $X2=0
+ $Y2=0
cc_240 N_A_58_367#_c_258_n N_VGND_c_507_n 0.015688f $X=0.845 $Y=0.42 $X2=0 $Y2=0
cc_241 N_A_58_367#_c_231_n N_VGND_c_508_n 0.0257093f $X=1.69 $Y=1.08 $X2=0 $Y2=0
cc_242 N_A_58_367#_M1005_g N_VGND_c_509_n 0.00519269f $X=2.645 $Y=0.665 $X2=0
+ $Y2=0
cc_243 N_A_58_367#_c_233_n N_VGND_c_509_n 0.0260407f $X=2.425 $Y=1.08 $X2=0
+ $Y2=0
cc_244 N_A_58_367#_M1005_g N_VGND_c_510_n 6.46604e-19 $X=2.645 $Y=0.665 $X2=0
+ $Y2=0
cc_245 N_A_58_367#_M1011_g N_VGND_c_510_n 0.0116199f $X=3.075 $Y=0.665 $X2=0
+ $Y2=0
cc_246 N_A_58_367#_M1014_g N_VGND_c_510_n 0.0115373f $X=3.505 $Y=0.665 $X2=0
+ $Y2=0
cc_247 N_A_58_367#_M1015_g N_VGND_c_510_n 6.31838e-19 $X=3.935 $Y=0.665 $X2=0
+ $Y2=0
cc_248 N_A_58_367#_M1014_g N_VGND_c_511_n 0.00477554f $X=3.505 $Y=0.665 $X2=0
+ $Y2=0
cc_249 N_A_58_367#_M1015_g N_VGND_c_511_n 0.00575161f $X=3.935 $Y=0.665 $X2=0
+ $Y2=0
cc_250 N_A_58_367#_M1015_g N_VGND_c_512_n 0.00333511f $X=3.935 $Y=0.665 $X2=0
+ $Y2=0
cc_251 N_A_58_367#_c_265_n N_VGND_c_513_n 0.0189236f $X=1.855 $Y=0.37 $X2=0
+ $Y2=0
cc_252 N_A_58_367#_M1005_g N_VGND_c_515_n 0.00575161f $X=2.645 $Y=0.665 $X2=0
+ $Y2=0
cc_253 N_A_58_367#_M1011_g N_VGND_c_515_n 0.00477554f $X=3.075 $Y=0.665 $X2=0
+ $Y2=0
cc_254 N_A_58_367#_M1004_d N_VGND_c_518_n 0.00380103f $X=0.705 $Y=0.245 $X2=0
+ $Y2=0
cc_255 N_A_58_367#_M1007_d N_VGND_c_518_n 0.00223559f $X=1.715 $Y=0.245 $X2=0
+ $Y2=0
cc_256 N_A_58_367#_M1005_g N_VGND_c_518_n 0.0110258f $X=2.645 $Y=0.665 $X2=0
+ $Y2=0
cc_257 N_A_58_367#_M1011_g N_VGND_c_518_n 0.00825815f $X=3.075 $Y=0.665 $X2=0
+ $Y2=0
cc_258 N_A_58_367#_M1014_g N_VGND_c_518_n 0.00825815f $X=3.505 $Y=0.665 $X2=0
+ $Y2=0
cc_259 N_A_58_367#_M1015_g N_VGND_c_518_n 0.0118351f $X=3.935 $Y=0.665 $X2=0
+ $Y2=0
cc_260 N_A_58_367#_c_258_n N_VGND_c_518_n 0.00984745f $X=0.845 $Y=0.42 $X2=0
+ $Y2=0
cc_261 N_A_58_367#_c_265_n N_VGND_c_518_n 0.0123859f $X=1.855 $Y=0.37 $X2=0
+ $Y2=0
cc_262 A_141_367# N_VPWR_c_385_n 0.00899413f $X=0.705 $Y=1.835 $X2=0 $Y2=0
cc_263 A_213_367# N_VPWR_c_385_n 0.0167135f $X=1.065 $Y=1.835 $X2=0 $Y2=0
cc_264 A_321_367# N_VPWR_c_385_n 0.0167135f $X=1.605 $Y=1.835 $X2=0 $Y2=0
cc_265 N_VPWR_c_385_n N_X_M1001_s 0.00536646f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_266 N_VPWR_c_385_n N_X_M1006_s 0.00536646f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_267 N_VPWR_c_391_n N_X_c_486_n 0.0124525f $X=3.125 $Y=3.33 $X2=0 $Y2=0
cc_268 N_VPWR_c_385_n N_X_c_486_n 0.00730901f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_M1003_d N_X_c_447_n 0.00176461f $X=3.15 $Y=1.835 $X2=0 $Y2=0
cc_270 N_VPWR_c_387_n N_X_c_447_n 0.0170777f $X=3.29 $Y=2.19 $X2=0 $Y2=0
cc_271 N_VPWR_c_393_n N_X_c_490_n 0.0124525f $X=3.985 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_c_385_n N_X_c_490_n 0.00730901f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_273 N_VPWR_M1010_d N_X_c_449_n 0.00267685f $X=4.01 $Y=1.835 $X2=0 $Y2=0
cc_274 N_VPWR_c_388_n N_X_c_449_n 0.0220026f $X=4.15 $Y=2.19 $X2=0 $Y2=0
cc_275 N_X_c_440_n N_VGND_c_510_n 0.0216087f $X=3.625 $Y=1.17 $X2=0 $Y2=0
cc_276 N_X_c_495_p N_VGND_c_511_n 0.0136943f $X=3.72 $Y=0.42 $X2=0 $Y2=0
cc_277 N_X_c_442_n N_VGND_c_512_n 0.0196987f $X=4.43 $Y=1.17 $X2=0 $Y2=0
cc_278 X N_VGND_c_512_n 0.0357926f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_279 N_X_c_498_p N_VGND_c_515_n 0.0124525f $X=2.86 $Y=0.42 $X2=0 $Y2=0
cc_280 X N_VGND_c_517_n 0.00773544f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_281 N_X_M1005_s N_VGND_c_518_n 0.00536646f $X=2.72 $Y=0.245 $X2=0 $Y2=0
cc_282 N_X_M1014_s N_VGND_c_518_n 0.0041489f $X=3.58 $Y=0.245 $X2=0 $Y2=0
cc_283 N_X_c_498_p N_VGND_c_518_n 0.00730901f $X=2.86 $Y=0.42 $X2=0 $Y2=0
cc_284 N_X_c_495_p N_VGND_c_518_n 0.00866972f $X=3.72 $Y=0.42 $X2=0 $Y2=0
cc_285 X N_VGND_c_518_n 0.00881366f $X=4.475 $Y=0.47 $X2=0 $Y2=0
