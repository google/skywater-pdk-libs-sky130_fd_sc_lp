* File: sky130_fd_sc_lp__or3_4.pex.spice
* Created: Wed Sep  2 10:30:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3_4%C 3 7 9 10 14
r28 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=1.46
+ $X2=0.635 $Y2=1.625
r29 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=1.46
+ $X2=0.635 $Y2=1.295
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=1.46 $X2=0.635 $Y2=1.46
r31 10 15 2.6122 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.562
+ $X2=0.635 $Y2=1.562
r32 9 15 12.1391 $w=3.73e-07 $l=3.95e-07 $layer=LI1_cond $X=0.24 $Y=1.562
+ $X2=0.635 $Y2=1.562
r33 7 17 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.725 $Y=2.465
+ $X2=0.725 $Y2=1.625
r34 3 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.725 $Y=0.665
+ $X2=0.725 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_4%B 3 7 9 12 13
c33 3 0 1.78332e-19 $X=1.085 $Y=2.465
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.51
+ $X2=1.175 $Y2=1.675
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.51
+ $X2=1.175 $Y2=1.345
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.175
+ $Y=1.51 $X2=1.175 $Y2=1.51
r37 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.19 $Y=1.665
+ $X2=1.19 $Y2=1.51
r38 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.235 $Y=0.665
+ $X2=1.235 $Y2=1.345
r39 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.085 $Y=2.465
+ $X2=1.085 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_4%A 3 7 9 12 13
c41 13 0 1.78332e-19 $X=1.715 $Y=1.51
r42 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.51
+ $X2=1.715 $Y2=1.675
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.51
+ $X2=1.715 $Y2=1.345
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.715
+ $Y=1.51 $X2=1.715 $Y2=1.51
r45 9 13 6.26767 $w=2.83e-07 $l=1.55e-07 $layer=LI1_cond $X=1.667 $Y=1.665
+ $X2=1.667 $Y2=1.51
r46 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.665 $Y=0.665
+ $X2=1.665 $Y2=1.345
r47 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.625 $Y=2.465
+ $X2=1.625 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_4%A_77_49# 1 2 3 12 16 20 24 28 32 36 40 44 46
+ 48 50 51 52 56 58 61 63 69 70 74 75
r146 80 81 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.06 $Y=1.51
+ $X2=3.49 $Y2=1.51
r147 79 80 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.63 $Y=1.51
+ $X2=3.06 $Y2=1.51
r148 70 81 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.65 $Y=1.51
+ $X2=3.49 $Y2=1.51
r149 69 70 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.65
+ $Y=1.51 $X2=3.65 $Y2=1.51
r150 67 79 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.29 $Y=1.51
+ $X2=2.63 $Y2=1.51
r151 67 76 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.29 $Y=1.51 $X2=2.2
+ $Y2=1.51
r152 66 69 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.29 $Y=1.51
+ $X2=3.65 $Y2=1.51
r153 66 67 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.51 $X2=2.29 $Y2=1.51
r154 64 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=1.51
+ $X2=2.065 $Y2=1.51
r155 64 66 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.15 $Y=1.51
+ $X2=2.29 $Y2=1.51
r156 62 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=1.595
+ $X2=2.065 $Y2=1.51
r157 62 63 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.065 $Y=1.595
+ $X2=2.065 $Y2=1.92
r158 61 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=1.425
+ $X2=2.065 $Y2=1.51
r159 60 61 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.065 $Y=1.165
+ $X2=2.065 $Y2=1.425
r160 59 74 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.595 $Y=1.08
+ $X2=1.452 $Y2=1.08
r161 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.98 $Y=1.08
+ $X2=2.065 $Y2=1.165
r162 58 59 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.98 $Y=1.08
+ $X2=1.595 $Y2=1.08
r163 54 74 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.452 $Y=0.995
+ $X2=1.452 $Y2=1.08
r164 54 56 23.251 $w=2.83e-07 $l=5.75e-07 $layer=LI1_cond $X=1.452 $Y=0.995
+ $X2=1.452 $Y2=0.42
r165 53 73 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.675 $Y=2.01
+ $X2=0.51 $Y2=2.01
r166 52 63 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.98 $Y=2.01
+ $X2=2.065 $Y2=1.92
r167 52 53 80.4091 $w=1.78e-07 $l=1.305e-06 $layer=LI1_cond $X=1.98 $Y=2.01
+ $X2=0.675 $Y2=2.01
r168 50 74 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.31 $Y=1.08
+ $X2=1.452 $Y2=1.08
r169 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.31 $Y=1.08
+ $X2=0.64 $Y2=1.08
r170 46 73 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.51 $Y=2.1 $X2=0.51
+ $Y2=2.01
r171 46 48 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.51 $Y=2.1
+ $X2=0.51 $Y2=2.95
r172 42 51 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=0.492 $Y=0.995
+ $X2=0.64 $Y2=1.08
r173 42 44 22.4629 $w=2.93e-07 $l=5.75e-07 $layer=LI1_cond $X=0.492 $Y=0.995
+ $X2=0.492 $Y2=0.42
r174 38 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=1.675
+ $X2=3.49 $Y2=1.51
r175 38 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.49 $Y=1.675
+ $X2=3.49 $Y2=2.465
r176 34 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=1.345
+ $X2=3.49 $Y2=1.51
r177 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.49 $Y=1.345
+ $X2=3.49 $Y2=0.665
r178 30 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.675
+ $X2=3.06 $Y2=1.51
r179 30 32 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.06 $Y=1.675
+ $X2=3.06 $Y2=2.465
r180 26 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.345
+ $X2=3.06 $Y2=1.51
r181 26 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.06 $Y=1.345
+ $X2=3.06 $Y2=0.665
r182 22 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.63 $Y=1.675
+ $X2=2.63 $Y2=1.51
r183 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.63 $Y=1.675
+ $X2=2.63 $Y2=2.465
r184 18 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.63 $Y=1.345
+ $X2=2.63 $Y2=1.51
r185 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.63 $Y=1.345
+ $X2=2.63 $Y2=0.665
r186 14 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.675
+ $X2=2.2 $Y2=1.51
r187 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.2 $Y=1.675
+ $X2=2.2 $Y2=2.465
r188 10 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.345
+ $X2=2.2 $Y2=1.51
r189 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.2 $Y=1.345
+ $X2=2.2 $Y2=0.665
r190 3 73 400 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.385
+ $Y=1.835 $X2=0.51 $Y2=2.045
r191 3 48 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.385
+ $Y=1.835 $X2=0.51 $Y2=2.95
r192 2 56 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.31
+ $Y=0.245 $X2=1.45 $Y2=0.42
r193 1 44 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=0.385
+ $Y=0.245 $X2=0.51 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_4%VPWR 1 2 3 12 16 20 24 29 30 31 32 33 47 48 51
r52 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 48 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 45 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.87 $Y=3.33
+ $X2=3.705 $Y2=3.33
r56 45 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.87 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 44 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 37 41 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 36 40 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 33 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 31 43 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r66 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=3.33
+ $X2=2.845 $Y2=3.33
r67 29 40 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.745 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 29 30 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.745 $Y=3.33
+ $X2=1.922 $Y2=3.33
r69 28 43 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.1 $Y=3.33 $X2=2.64
+ $Y2=3.33
r70 28 30 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=2.1 $Y=3.33
+ $X2=1.922 $Y2=3.33
r71 24 27 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=3.705 $Y=2.2
+ $X2=3.705 $Y2=2.95
r72 22 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=3.245
+ $X2=3.705 $Y2=3.33
r73 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.705 $Y=3.245
+ $X2=3.705 $Y2=2.95
r74 21 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=3.33
+ $X2=2.845 $Y2=3.33
r75 20 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=3.33
+ $X2=3.705 $Y2=3.33
r76 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.54 $Y=3.33
+ $X2=3.01 $Y2=3.33
r77 16 19 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.845 $Y=2.2
+ $X2=2.845 $Y2=2.97
r78 14 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=3.245
+ $X2=2.845 $Y2=3.33
r79 14 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.845 $Y=3.245
+ $X2=2.845 $Y2=2.97
r80 10 30 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.922 $Y=3.245
+ $X2=1.922 $Y2=3.33
r81 10 12 27.1068 $w=3.53e-07 $l=8.35e-07 $layer=LI1_cond $X=1.922 $Y=3.245
+ $X2=1.922 $Y2=2.41
r82 3 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.835 $X2=3.705 $Y2=2.95
r83 3 24 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.835 $X2=3.705 $Y2=2.2
r84 2 19 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.835 $X2=2.845 $Y2=2.97
r85 2 16 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.835 $X2=2.845 $Y2=2.2
r86 1 12 300 $w=1.7e-07 $l=6.71844e-07 $layer=licon1_PDIFF $count=2 $X=1.7
+ $Y=1.835 $X2=1.91 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41 42
+ 44 45 46 47 61
r67 59 61 3.08081 $w=1.78e-07 $l=5e-08 $layer=LI1_cond $X=4.075 $Y=1.245
+ $X2=4.075 $Y2=1.295
r68 46 53 4.86787 $w=1.82e-07 $l=8.5e-08 $layer=LI1_cond $X=4.072 $Y=1.16
+ $X2=4.072 $Y2=1.075
r69 46 59 4.86787 $w=1.82e-07 $l=8.6487e-08 $layer=LI1_cond $X=4.072 $Y=1.16
+ $X2=4.075 $Y2=1.245
r70 46 47 21.7505 $w=1.78e-07 $l=3.53e-07 $layer=LI1_cond $X=4.075 $Y=1.312
+ $X2=4.075 $Y2=1.665
r71 46 61 1.04747 $w=1.78e-07 $l=1.7e-08 $layer=LI1_cond $X=4.075 $Y=1.312
+ $X2=4.075 $Y2=1.295
r72 45 53 8.99263 $w=1.83e-07 $l=1.5e-07 $layer=LI1_cond $X=4.072 $Y=0.925
+ $X2=4.072 $Y2=1.075
r73 44 45 22.1818 $w=1.83e-07 $l=3.7e-07 $layer=LI1_cond $X=4.072 $Y=0.555
+ $X2=4.072 $Y2=0.925
r74 43 47 6.77778 $w=1.78e-07 $l=1.1e-07 $layer=LI1_cond $X=4.075 $Y=1.775
+ $X2=4.075 $Y2=1.665
r75 40 41 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.405 $Y=1.16
+ $X2=3.292 $Y2=1.16
r76 39 46 1.59926 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=3.98 $Y=1.16
+ $X2=4.072 $Y2=1.16
r77 39 40 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.98 $Y=1.16
+ $X2=3.405 $Y2=1.16
r78 38 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.37 $Y=1.86
+ $X2=3.275 $Y2=1.86
r79 37 43 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.985 $Y=1.86
+ $X2=4.075 $Y2=1.775
r80 37 38 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.985 $Y=1.86
+ $X2=3.37 $Y2=1.86
r81 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.275 $Y=1.98
+ $X2=3.275 $Y2=2.91
r82 31 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=1.945
+ $X2=3.275 $Y2=1.86
r83 31 33 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=3.275 $Y=1.945
+ $X2=3.275 $Y2=1.98
r84 27 41 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.292 $Y=1.075
+ $X2=3.292 $Y2=1.16
r85 27 29 33.5489 $w=2.23e-07 $l=6.55e-07 $layer=LI1_cond $X=3.292 $Y=1.075
+ $X2=3.292 $Y2=0.42
r86 25 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.18 $Y=1.86
+ $X2=3.275 $Y2=1.86
r87 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.18 $Y=1.86
+ $X2=2.51 $Y2=1.86
r88 23 41 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.18 $Y=1.16
+ $X2=3.292 $Y2=1.16
r89 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.18 $Y=1.16
+ $X2=2.51 $Y2=1.16
r90 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.415 $Y=1.98
+ $X2=2.415 $Y2=2.91
r91 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.415 $Y=1.945
+ $X2=2.51 $Y2=1.86
r92 17 19 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=2.415 $Y=1.945
+ $X2=2.415 $Y2=1.98
r93 13 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.415 $Y=1.075
+ $X2=2.51 $Y2=1.16
r94 13 15 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=2.415 $Y=1.075
+ $X2=2.415 $Y2=0.42
r95 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.135
+ $Y=1.835 $X2=3.275 $Y2=2.91
r96 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.135
+ $Y=1.835 $X2=3.275 $Y2=1.98
r97 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.835 $X2=2.415 $Y2=2.91
r98 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.835 $X2=2.415 $Y2=1.98
r99 2 29 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.135
+ $Y=0.245 $X2=3.275 $Y2=0.42
r100 1 15 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.275
+ $Y=0.245 $X2=2.415 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_4%VGND 1 2 3 4 15 19 23 25 29 32 33 35 36 37 38
+ 39 53 54 57
r61 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r62 54 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r63 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r64 51 57 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.692
+ $Y2=0
r65 51 53 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=4.08
+ $Y2=0
r66 50 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r67 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 43 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r70 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r71 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r72 39 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r73 37 49 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.64
+ $Y2=0
r74 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.845
+ $Y2=0
r75 35 46 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r76 35 36 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.947
+ $Y2=0
r77 34 49 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=2.64
+ $Y2=0
r78 34 36 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=1.947
+ $Y2=0
r79 32 42 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.72
+ $Y2=0
r80 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.975
+ $Y2=0
r81 31 46 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.14 $Y=0 $X2=1.68
+ $Y2=0
r82 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=0 $X2=0.975
+ $Y2=0
r83 27 57 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.692 $Y=0.085
+ $X2=3.692 $Y2=0
r84 27 29 14.9572 $w=2.33e-07 $l=3.05e-07 $layer=LI1_cond $X=3.692 $Y=0.085
+ $X2=3.692 $Y2=0.39
r85 26 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=0 $X2=2.845
+ $Y2=0
r86 25 57 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=3.575 $Y=0 $X2=3.692
+ $Y2=0
r87 25 26 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.575 $Y=0 $X2=3.01
+ $Y2=0
r88 21 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0
r89 21 23 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0.39
r90 17 36 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.947 $Y=0.085
+ $X2=1.947 $Y2=0
r91 17 19 8.99853 $w=3.63e-07 $l=2.85e-07 $layer=LI1_cond $X=1.947 $Y=0.085
+ $X2=1.947 $Y2=0.37
r92 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0
r93 13 15 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0.37
r94 4 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.565
+ $Y=0.245 $X2=3.705 $Y2=0.39
r95 3 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.705
+ $Y=0.245 $X2=2.845 $Y2=0.39
r96 2 19 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=1.74
+ $Y=0.245 $X2=1.93 $Y2=0.37
r97 1 15 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=0.8
+ $Y=0.245 $X2=0.975 $Y2=0.37
.ends

