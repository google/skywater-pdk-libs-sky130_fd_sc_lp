# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xnor2_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__xnor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.415000 1.570000 1.750000 ;
        RECT 1.285000 1.750000 1.570000 1.930000 ;
        RECT 1.285000 1.930000 6.475000 1.935000 ;
        RECT 1.285000 1.935000 3.670000 2.100000 ;
        RECT 3.500000 1.415000 3.830000 1.765000 ;
        RECT 3.500000 1.765000 6.475000 1.930000 ;
        RECT 6.305000 1.425000 7.960000 1.595000 ;
        RECT 6.305000 1.595000 6.475000 1.765000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.810000 1.415000 3.160000 1.595000 ;
        RECT 2.075000 1.595000 3.160000 1.750000 ;
        RECT 8.240000 1.425000 9.590000 1.750000 ;
      LAYER mcon ;
        RECT 2.075000 1.580000 2.245000 1.750000 ;
        RECT 8.315000 1.580000 8.485000 1.750000 ;
      LAYER met1 ;
        RECT 2.015000 1.550000 2.305000 1.595000 ;
        RECT 2.015000 1.595000 8.545000 1.735000 ;
        RECT 2.015000 1.735000 2.305000 1.780000 ;
        RECT 8.255000 1.550000 8.545000 1.595000 ;
        RECT 8.255000 1.735000 8.545000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.940400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.075000 5.435000 1.245000 ;
        RECT 0.095000 1.245000 0.275000 1.920000 ;
        RECT 0.095000 1.920000 1.115000 2.090000 ;
        RECT 0.945000 2.090000 1.115000 2.270000 ;
        RECT 0.945000 2.270000 6.080000 2.275000 ;
        RECT 0.945000 2.275000 4.645000 2.450000 ;
        RECT 4.165000 2.105000 6.080000 2.270000 ;
        RECT 4.215000 2.450000 4.645000 3.075000 ;
        RECT 4.235000 0.605000 4.435000 1.075000 ;
        RECT 5.105000 0.595000 5.435000 1.075000 ;
        RECT 5.820000 2.275000 6.080000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
        RECT 0.635000  0.085000  0.965000 0.565000 ;
        RECT 1.505000  0.085000  1.835000 0.565000 ;
        RECT 2.365000  0.085000  2.695000 0.565000 ;
        RECT 3.225000  0.085000  3.555000 0.565000 ;
        RECT 6.635000  0.085000  6.965000 0.575000 ;
        RECT 7.505000  0.085000  7.835000 0.575000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
        RECT 9.755000 -0.085000 9.925000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.080000 3.415000 ;
        RECT 0.095000 2.260000  0.425000 3.245000 ;
        RECT 1.035000 2.960000  1.365000 3.245000 ;
        RECT 3.715000 2.620000  4.045000 3.245000 ;
        RECT 4.815000 2.445000  5.650000 3.245000 ;
        RECT 6.250000 2.125000  6.470000 3.245000 ;
        RECT 7.040000 2.125000  7.370000 3.245000 ;
        RECT 7.900000 2.260000  8.230000 3.245000 ;
        RECT 8.760000 2.260000  9.090000 3.245000 ;
        RECT 9.620000 2.260000  9.950000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
        RECT 9.755000 3.245000 9.925000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.135000 0.295000 0.465000 0.735000 ;
      RECT 0.135000 0.735000 4.065000 0.905000 ;
      RECT 0.595000 2.620000 3.545000 2.790000 ;
      RECT 0.595000 2.790000 0.865000 2.950000 ;
      RECT 1.155000 0.285000 1.335000 0.735000 ;
      RECT 1.535000 2.790000 3.545000 2.960000 ;
      RECT 2.005000 0.285000 2.195000 0.735000 ;
      RECT 2.865000 0.285000 3.055000 0.735000 ;
      RECT 3.735000 0.255000 5.935000 0.425000 ;
      RECT 3.735000 0.425000 4.935000 0.435000 ;
      RECT 3.735000 0.435000 4.065000 0.735000 ;
      RECT 4.040000 1.415000 6.135000 1.585000 ;
      RECT 4.605000 0.435000 4.935000 0.905000 ;
      RECT 5.605000 0.425000 5.935000 0.915000 ;
      RECT 5.625000 1.085000 9.990000 1.255000 ;
      RECT 5.625000 1.255000 6.135000 1.415000 ;
      RECT 6.135000 0.305000 6.465000 0.745000 ;
      RECT 6.135000 0.745000 8.195000 0.915000 ;
      RECT 6.645000 1.775000 7.800000 1.920000 ;
      RECT 6.645000 1.920000 9.990000 1.945000 ;
      RECT 6.645000 1.945000 6.870000 3.075000 ;
      RECT 7.135000 0.285000 7.335000 0.745000 ;
      RECT 7.540000 1.945000 9.990000 2.090000 ;
      RECT 7.540000 2.090000 7.730000 3.075000 ;
      RECT 8.005000 0.255000 9.985000 0.425000 ;
      RECT 8.005000 0.425000 9.055000 0.435000 ;
      RECT 8.005000 0.435000 8.195000 0.745000 ;
      RECT 8.365000 0.615000 8.695000 1.065000 ;
      RECT 8.365000 1.065000 9.990000 1.085000 ;
      RECT 8.400000 2.090000 8.590000 3.075000 ;
      RECT 8.865000 0.435000 9.055000 0.895000 ;
      RECT 9.225000 0.615000 9.555000 1.065000 ;
      RECT 9.260000 2.090000 9.450000 3.075000 ;
      RECT 9.725000 0.425000 9.985000 0.895000 ;
      RECT 9.770000 1.255000 9.990000 1.920000 ;
  END
END sky130_fd_sc_lp__xnor2_4
