* File: sky130_fd_sc_lp__mux2_1.pex.spice
* Created: Fri Aug 28 10:43:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2_1%A_105_22# 1 2 9 12 16 17 19 20 23 26 29
c65 19 0 1.30219e-19 $X=1.775 $Y=1.075
r66 21 26 8.31818 $w=3.52e-07 $l=3.35142e-07 $layer=LI1_cond $X=2.18 $Y=1.16
+ $X2=1.94 $Y2=0.932
r67 21 23 63.6463 $w=2.18e-07 $l=1.215e-06 $layer=LI1_cond $X=2.18 $Y=1.16
+ $X2=2.18 $Y2=2.375
r68 19 26 8.99038 $w=3.52e-07 $l=2.25433e-07 $layer=LI1_cond $X=1.775 $Y=1.075
+ $X2=1.94 $Y2=0.932
r69 19 20 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.775 $Y=1.075
+ $X2=0.9 $Y2=1.075
r70 17 30 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.712 $Y=1.355
+ $X2=0.712 $Y2=1.52
r71 17 29 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.712 $Y=1.355
+ $X2=0.712 $Y2=1.19
r72 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.735
+ $Y=1.355 $X2=0.735 $Y2=1.355
r73 14 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.77 $Y=1.16
+ $X2=0.9 $Y2=1.075
r74 14 16 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=0.77 $Y=1.16
+ $X2=0.77 $Y2=1.355
r75 12 30 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=0.6 $Y=2.465
+ $X2=0.6 $Y2=1.52
r76 9 29 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.6 $Y=0.66 $X2=0.6
+ $Y2=1.19
r77 2 23 600 $w=1.7e-07 $l=4.76603e-07 $layer=licon1_PDIFF $count=1 $X=1.8
+ $Y=2.17 $X2=2.185 $Y2=2.375
r78 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.8
+ $Y=0.66 $X2=1.94 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_1%S 3 7 11 15 19 20 23 24 26 27 28 29 30 35 36
+ 41
r95 39 41 1.26488 $w=4.08e-07 $l=4.5e-08 $layer=LI1_cond $X=3.075 $Y=1.925
+ $X2=3.12 $Y2=1.925
r96 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=1.845
+ $X2=3.685 $Y2=2.01
r97 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=1.845
+ $X2=3.685 $Y2=1.68
r98 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=1.845 $X2=3.685 $Y2=1.845
r99 30 39 2.47908 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=1.925
+ $X2=3.075 $Y2=1.925
r100 30 36 15.3191 $w=4.08e-07 $l=5.45e-07 $layer=LI1_cond $X=3.14 $Y=1.925
+ $X2=3.685 $Y2=1.925
r101 30 41 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=3.14 $Y=1.925
+ $X2=3.12 $Y2=1.925
r102 28 30 5.97895 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.99 $Y=2.13
+ $X2=2.99 $Y2=1.925
r103 28 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.99 $Y=2.13
+ $X2=2.99 $Y2=2.885
r104 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=2.97
+ $X2=2.99 $Y2=2.885
r105 26 27 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=2.905 $Y=2.97
+ $X2=1.36 $Y2=2.97
r106 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.275
+ $Y=1.505 $X2=1.275 $Y2=1.505
r107 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.275 $Y=2.885
+ $X2=1.36 $Y2=2.97
r108 21 23 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.275 $Y=2.885
+ $X2=1.275 $Y2=1.505
r109 19 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.275 $Y=1.845
+ $X2=1.275 $Y2=1.505
r110 19 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.275 $Y=1.845
+ $X2=1.275 $Y2=2.01
r111 18 24 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.275 $Y=1.34
+ $X2=1.275 $Y2=1.505
r112 15 38 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.595 $Y=2.38
+ $X2=3.595 $Y2=2.01
r113 11 37 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.595 $Y=0.87
+ $X2=3.595 $Y2=1.68
r114 7 20 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.365 $Y=2.38
+ $X2=1.365 $Y2=2.01
r115 3 18 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.255 $Y=0.87 $X2=1.255
+ $Y2=1.34
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_1%A1 3 6 8 11 13 14 15 16 17 18 28 30 34 36
r62 34 36 0.83814 $w=2.73e-07 $l=2e-08 $layer=LI1_cond $X=2.597 $Y=0.535
+ $X2=2.597 $Y2=0.555
r63 30 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.605 $Y=1.845
+ $X2=2.605 $Y2=2.01
r64 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.605
+ $Y=1.845 $X2=2.605 $Y2=1.845
r65 17 18 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.597 $Y=2.035
+ $X2=2.597 $Y2=2.405
r66 17 31 7.96233 $w=2.73e-07 $l=1.9e-07 $layer=LI1_cond $X=2.597 $Y=2.035
+ $X2=2.597 $Y2=1.845
r67 16 31 7.54326 $w=2.73e-07 $l=1.8e-07 $layer=LI1_cond $X=2.597 $Y=1.665
+ $X2=2.597 $Y2=1.845
r68 15 16 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.597 $Y=1.295
+ $X2=2.597 $Y2=1.665
r69 14 15 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.597 $Y=0.925
+ $X2=2.597 $Y2=1.295
r70 13 34 3.44552 $w=2.75e-07 $l=1.4e-07 $layer=LI1_cond $X=2.597 $Y=0.395
+ $X2=2.597 $Y2=0.535
r71 13 14 14.1646 $w=2.73e-07 $l=3.38e-07 $layer=LI1_cond $X=2.597 $Y=0.587
+ $X2=2.597 $Y2=0.925
r72 13 36 1.34102 $w=2.73e-07 $l=3.2e-08 $layer=LI1_cond $X=2.597 $Y=0.587
+ $X2=2.597 $Y2=0.555
r73 11 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=0.385
+ $X2=1.705 $Y2=0.55
r74 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.705
+ $Y=0.385 $X2=1.705 $Y2=0.385
r75 8 13 3.37169 $w=2.8e-07 $l=1.37e-07 $layer=LI1_cond $X=2.46 $Y=0.395
+ $X2=2.597 $Y2=0.395
r76 8 10 31.0748 $w=2.78e-07 $l=7.55e-07 $layer=LI1_cond $X=2.46 $Y=0.395
+ $X2=1.705 $Y2=0.395
r77 6 33 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.515 $Y=2.38
+ $X2=2.515 $Y2=2.01
r78 3 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.725 $Y=0.87
+ $X2=1.725 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_1%A0 3 7 9 10 11 20
c39 20 0 1.30219e-19 $X=2.155 $Y=1.745
r40 18 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.815 $Y=1.745
+ $X2=2.155 $Y2=1.745
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.815
+ $Y=1.745 $X2=1.815 $Y2=1.745
r42 15 18 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.725 $Y=1.745
+ $X2=1.815 $Y2=1.745
r43 10 11 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.715 $Y=2.035
+ $X2=1.715 $Y2=2.405
r44 10 19 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.715 $Y=2.035
+ $X2=1.715 $Y2=1.745
r45 9 19 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=1.715 $Y=1.665
+ $X2=1.715 $Y2=1.745
r46 5 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.58
+ $X2=2.155 $Y2=1.745
r47 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.155 $Y=1.58
+ $X2=2.155 $Y2=0.87
r48 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.91
+ $X2=1.725 $Y2=1.745
r49 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.725 $Y=1.91 $X2=1.725
+ $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_1%A_488_106# 1 2 9 11 12 15 17 22 28 31 32 33
r58 30 32 5.86749 $w=2.82e-07 $l=5.92453e-07 $layer=LI1_cond $X=4.115 $Y=1.55
+ $X2=3.665 $Y2=1.22
r59 30 31 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.115 $Y=1.55
+ $X2=4.115 $Y2=2.3
r60 26 32 5.86749 $w=2.82e-07 $l=1.97e-07 $layer=LI1_cond $X=3.862 $Y=1.22
+ $X2=3.665 $Y2=1.22
r61 26 28 10.2115 $w=3.93e-07 $l=3.5e-07 $layer=LI1_cond $X=3.862 $Y=1.22
+ $X2=3.862 $Y2=0.87
r62 22 31 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.03 $Y=2.435
+ $X2=4.115 $Y2=2.3
r63 22 24 9.39028 $w=2.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.03 $Y=2.435
+ $X2=3.81 $Y2=2.435
r64 20 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.385
+ $X2=3.145 $Y2=1.55
r65 20 33 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.145 $Y=1.385
+ $X2=3.145 $Y2=1.295
r66 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.145
+ $Y=1.385 $X2=3.145 $Y2=1.385
r67 17 32 0.789365 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=1.385
+ $X2=3.665 $Y2=1.22
r68 17 19 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.665 $Y=1.385
+ $X2=3.145 $Y2=1.385
r69 15 36 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.055 $Y=2.38
+ $X2=3.055 $Y2=1.55
r70 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.98 $Y=1.295
+ $X2=3.145 $Y2=1.295
r71 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.98 $Y=1.295
+ $X2=2.59 $Y2=1.295
r72 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.515 $Y=1.22
+ $X2=2.59 $Y2=1.295
r73 7 9 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.515 $Y=1.22
+ $X2=2.515 $Y2=0.87
r74 2 24 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=2.17 $X2=3.81 $Y2=2.405
r75 1 28 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.66 $X2=3.83 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_1%X 1 2 7 8 9 10 11 12 13 22
r12 13 41 4.04103 $w=3.83e-07 $l=1.35e-07 $layer=LI1_cond $X=0.277 $Y=2.775
+ $X2=0.277 $Y2=2.91
r13 12 13 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=2.405
+ $X2=0.277 $Y2=2.775
r14 11 12 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=2.035
+ $X2=0.277 $Y2=2.405
r15 11 33 1.64635 $w=3.83e-07 $l=5.5e-08 $layer=LI1_cond $X=0.277 $Y=2.035
+ $X2=0.277 $Y2=1.98
r16 10 33 9.42908 $w=3.83e-07 $l=3.15e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.98
r17 9 10 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.665
r18 8 9 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=0.925
+ $X2=0.277 $Y2=1.295
r19 7 8 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=0.555
+ $X2=0.277 $Y2=0.925
r20 7 22 4.04103 $w=3.83e-07 $l=1.35e-07 $layer=LI1_cond $X=0.277 $Y=0.555
+ $X2=0.277 $Y2=0.42
r21 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.835 $X2=0.385 $Y2=2.91
r22 2 33 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.835 $X2=0.385 $Y2=1.98
r23 1 22 91 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=2 $X=0.26
+ $Y=0.24 $X2=0.385 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_1%VPWR 1 2 11 19 22 23 24 34 35 38
r39 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r41 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r42 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 29 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 28 31 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 26 38 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.02 $Y=3.33
+ $X2=0.865 $Y2=3.33
r47 26 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.02 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 24 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 24 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 22 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 22 23 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.36 $Y2=3.33
r52 21 34 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.475 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 21 23 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.475 $Y=3.33
+ $X2=3.36 $Y2=3.33
r54 17 23 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=3.245
+ $X2=3.36 $Y2=3.33
r55 17 19 39.0829 $w=2.28e-07 $l=7.8e-07 $layer=LI1_cond $X=3.36 $Y=3.245
+ $X2=3.36 $Y2=2.465
r56 14 16 18.9595 $w=3.08e-07 $l=5.1e-07 $layer=LI1_cond $X=0.865 $Y=2.44
+ $X2=0.865 $Y2=2.95
r57 11 14 17.1008 $w=3.08e-07 $l=4.6e-07 $layer=LI1_cond $X=0.865 $Y=1.98
+ $X2=0.865 $Y2=2.44
r58 9 38 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=3.33
r59 9 16 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=2.95
r60 2 19 600 $w=1.7e-07 $l=3.89776e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.17 $X2=3.35 $Y2=2.465
r61 1 16 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=1.835 $X2=0.815 $Y2=2.95
r62 1 14 600 $w=1.7e-07 $l=7.23412e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=1.835 $X2=0.935 $Y2=2.44
r63 1 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=1.835 $X2=0.815 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_1%VGND 1 2 11 15 17 19 29 30 33 36
r42 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r45 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r46 27 36 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.2
+ $Y2=0
r47 27 29 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.495 $Y=0 $X2=4.08
+ $Y2=0
r48 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r49 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r50 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r52 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r54 20 22 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r55 19 36 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.2
+ $Y2=0
r56 19 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.64
+ $Y2=0
r57 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r58 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r59 13 36 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0.085 $X2=3.2
+ $Y2=0
r60 13 15 15.9139 $w=5.88e-07 $l=7.85e-07 $layer=LI1_cond $X=3.2 $Y=0.085
+ $X2=3.2 $Y2=0.87
r61 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r62 9 11 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.385
r63 2 15 91 $w=1.7e-07 $l=8.88819e-07 $layer=licon1_NDIFF $count=2 $X=2.59
+ $Y=0.66 $X2=3.38 $Y2=0.87
r64 1 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.675
+ $Y=0.24 $X2=0.815 $Y2=0.385
.ends

