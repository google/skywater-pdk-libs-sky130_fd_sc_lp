* File: sky130_fd_sc_lp__a2111o_m.pxi.spice
* Created: Wed Sep  2 09:16:37 2020
* 
x_PM_SKY130_FD_SC_LP__A2111O_M%A_85_21# N_A_85_21#_M1001_d N_A_85_21#_M1009_d
+ N_A_85_21#_M1011_s N_A_85_21#_M1010_g N_A_85_21#_M1007_g N_A_85_21#_c_85_n
+ N_A_85_21#_c_95_n N_A_85_21#_c_86_n N_A_85_21#_c_87_n N_A_85_21#_c_96_n
+ N_A_85_21#_c_97_n N_A_85_21#_c_88_n N_A_85_21#_c_89_n N_A_85_21#_c_90_n
+ N_A_85_21#_c_91_n N_A_85_21#_c_92_n PM_SKY130_FD_SC_LP__A2111O_M%A_85_21#
x_PM_SKY130_FD_SC_LP__A2111O_M%D1 N_D1_M1001_g N_D1_M1011_g N_D1_c_174_n
+ N_D1_c_175_n D1 D1 N_D1_c_176_n N_D1_c_179_n PM_SKY130_FD_SC_LP__A2111O_M%D1
x_PM_SKY130_FD_SC_LP__A2111O_M%C1 N_C1_M1006_g N_C1_M1003_g N_C1_c_220_n
+ N_C1_c_222_n C1 C1 PM_SKY130_FD_SC_LP__A2111O_M%C1
x_PM_SKY130_FD_SC_LP__A2111O_M%B1 N_B1_M1008_g N_B1_M1009_g N_B1_c_266_n B1 B1
+ N_B1_c_270_n N_B1_c_271_n N_B1_c_272_n PM_SKY130_FD_SC_LP__A2111O_M%B1
x_PM_SKY130_FD_SC_LP__A2111O_M%A1 N_A1_M1005_g N_A1_M1000_g N_A1_c_320_n
+ N_A1_c_318_n N_A1_c_321_n A1 A1 PM_SKY130_FD_SC_LP__A2111O_M%A1
x_PM_SKY130_FD_SC_LP__A2111O_M%A2 N_A2_M1002_g N_A2_M1004_g N_A2_c_366_n
+ N_A2_c_367_n N_A2_c_368_n A2 A2 N_A2_c_370_n PM_SKY130_FD_SC_LP__A2111O_M%A2
x_PM_SKY130_FD_SC_LP__A2111O_M%X N_X_M1010_s N_X_M1007_s X X X X X X X
+ PM_SKY130_FD_SC_LP__A2111O_M%X
x_PM_SKY130_FD_SC_LP__A2111O_M%VPWR N_VPWR_M1007_d N_VPWR_M1005_d N_VPWR_c_412_n
+ N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n
+ VPWR N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_411_n N_VPWR_c_421_n
+ PM_SKY130_FD_SC_LP__A2111O_M%VPWR
x_PM_SKY130_FD_SC_LP__A2111O_M%A_411_369# N_A_411_369#_M1008_d
+ N_A_411_369#_M1004_d N_A_411_369#_c_473_n N_A_411_369#_c_470_n
+ N_A_411_369#_c_471_n N_A_411_369#_c_472_n
+ PM_SKY130_FD_SC_LP__A2111O_M%A_411_369#
x_PM_SKY130_FD_SC_LP__A2111O_M%VGND N_VGND_M1010_d N_VGND_M1006_d N_VGND_M1002_d
+ N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n N_VGND_c_503_n N_VGND_c_504_n
+ N_VGND_c_505_n VGND N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n
+ N_VGND_c_509_n PM_SKY130_FD_SC_LP__A2111O_M%VGND
cc_1 VNB N_A_85_21#_M1010_g 0.0644046f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_2 VNB N_A_85_21#_c_85_n 0.00142488f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.975
cc_3 VNB N_A_85_21#_c_86_n 0.00402475f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.635
cc_4 VNB N_A_85_21#_c_87_n 0.019644f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.635
cc_5 VNB N_A_85_21#_c_88_n 0.00195279f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.51
cc_6 VNB N_A_85_21#_c_89_n 0.00550631f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=1.93
cc_7 VNB N_A_85_21#_c_90_n 0.022777f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=0.81
cc_8 VNB N_A_85_21#_c_91_n 0.00899387f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=0.81
cc_9 VNB N_A_85_21#_c_92_n 0.00136805f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.51
cc_10 VNB N_D1_M1001_g 0.0336543f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.845
cc_11 VNB N_D1_c_174_n 0.0264859f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_12 VNB N_D1_c_175_n 0.0101622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D1_c_176_n 0.0212449f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.47
cc_14 VNB N_C1_M1006_g 0.0334079f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.845
cc_15 VNB N_C1_M1003_g 0.0160544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C1_c_220_n 0.00945474f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.47
cc_17 VNB N_B1_M1009_g 0.0582153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_266_n 0.00485514f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.47
cc_19 VNB N_A1_M1005_g 8.1542e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_M1000_g 0.0529932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_318_n 0.010695f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_22 VNB N_A2_M1004_g 0.0168968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_c_366_n 0.0207539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_367_n 0.0249397f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.47
cc_25 VNB N_A2_c_368_n 0.0184894f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_26 VNB A2 0.0359616f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.14
cc_27 VNB N_A2_c_370_n 0.0194195f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.14
cc_28 VNB X 0.0145804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB X 0.0482264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_411_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.51
cc_31 VNB N_A_411_369#_c_470_n 0.00479367f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_32 VNB N_A_411_369#_c_471_n 0.00875383f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_33 VNB N_A_411_369#_c_472_n 0.00642375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_500_n 0.00295613f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_35 VNB N_VGND_c_501_n 0.00494119f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.745
cc_36 VNB N_VGND_c_502_n 0.0130452f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.635
cc_37 VNB N_VGND_c_503_n 0.0127707f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.975
cc_38 VNB N_VGND_c_504_n 0.0226052f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.635
cc_39 VNB N_VGND_c_505_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.635
cc_40 VNB N_VGND_c_506_n 0.0173969f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.035
cc_41 VNB N_VGND_c_507_n 0.0266536f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=1.93
cc_42 VNB N_VGND_c_508_n 0.00522083f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.51
cc_43 VNB N_VGND_c_509_n 0.192829f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=0.81
cc_44 VPB N_A_85_21#_M1007_g 0.0420156f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.745
cc_45 VPB N_A_85_21#_c_85_n 0.0260204f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.975
cc_46 VPB N_A_85_21#_c_95_n 0.0181495f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.14
cc_47 VPB N_A_85_21#_c_96_n 0.0103143f $X=-0.19 $Y=1.655 $X2=1.475 $Y2=2.035
cc_48 VPB N_A_85_21#_c_97_n 0.002407f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.035
cc_49 VPB N_A_85_21#_c_89_n 0.00146799f $X=-0.19 $Y=1.655 $X2=1.56 $Y2=1.93
cc_50 VPB N_D1_M1011_g 0.0178536f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_D1_c_175_n 0.00842792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_D1_c_179_n 0.00257727f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.975
cc_53 VPB N_C1_M1003_g 0.0265188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_C1_c_222_n 0.0684991f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_55 VPB C1 0.00950841f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_56 VPB N_B1_M1008_g 0.0302934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_B1_c_266_n 0.00591829f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.47
cc_58 VPB B1 0.00974708f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_59 VPB N_B1_c_270_n 0.0386395f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.635
cc_60 VPB N_B1_c_271_n 0.0061991f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.47
cc_61 VPB N_B1_c_272_n 0.00598815f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.93
cc_62 VPB N_A1_M1005_g 0.0147111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A1_c_320_n 0.0611492f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.47
cc_64 VPB N_A1_c_321_n 0.0172504f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.745
cc_65 VPB A1 0.0189919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB A1 0.0166222f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.635
cc_67 VPB N_A2_M1004_g 0.0235671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB X 0.0420159f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB X 0.0142745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_412_n 0.0117912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_413_n 0.0145601f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_72 VPB N_VPWR_c_414_n 0.00111297f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.745
cc_73 VPB N_VPWR_c_415_n 0.00308345f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.47
cc_74 VPB N_VPWR_c_416_n 0.0396439f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.93
cc_75 VPB N_VPWR_c_417_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.635
cc_76 VPB N_VPWR_c_418_n 0.0201169f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_419_n 0.024496f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=0.725
cc_78 VPB N_VPWR_c_411_n 0.0850672f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=0.51
cc_79 VPB N_VPWR_c_421_n 0.00401341f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=0.81
cc_80 VPB N_A_411_369#_c_473_n 0.00128085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_411_369#_c_470_n 0.00647715f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_82 VPB N_A_411_369#_c_471_n 0.00128625f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_83 VPB N_A_411_369#_c_472_n 0.0191565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 N_A_85_21#_M1010_g N_D1_M1001_g 0.0170758f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_85_21#_c_88_n N_D1_M1001_g 0.0017629f $X=1.365 $Y=0.51 $X2=0 $Y2=0
cc_86 N_A_85_21#_c_89_n N_D1_M1001_g 0.00225047f $X=1.56 $Y=1.93 $X2=0 $Y2=0
cc_87 N_A_85_21#_c_91_n N_D1_M1001_g 0.00544896f $X=1.645 $Y=0.81 $X2=0 $Y2=0
cc_88 N_A_85_21#_M1007_g N_D1_M1011_g 0.00431797f $X=0.5 $Y=2.745 $X2=0 $Y2=0
cc_89 N_A_85_21#_c_85_n N_D1_M1011_g 0.00874466f $X=0.59 $Y=1.975 $X2=0 $Y2=0
cc_90 N_A_85_21#_c_86_n N_D1_M1011_g 7.15973e-19 $X=0.59 $Y=1.635 $X2=0 $Y2=0
cc_91 N_A_85_21#_c_96_n N_D1_M1011_g 0.0100231f $X=1.475 $Y=2.035 $X2=0 $Y2=0
cc_92 N_A_85_21#_c_86_n N_D1_c_174_n 6.73349e-19 $X=0.59 $Y=1.635 $X2=0 $Y2=0
cc_93 N_A_85_21#_c_87_n N_D1_c_174_n 0.00665769f $X=0.59 $Y=1.635 $X2=0 $Y2=0
cc_94 N_A_85_21#_c_85_n N_D1_c_175_n 0.00665769f $X=0.59 $Y=1.975 $X2=0 $Y2=0
cc_95 N_A_85_21#_c_96_n N_D1_c_175_n 0.00117387f $X=1.475 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_85_21#_c_89_n N_D1_c_175_n 0.00490404f $X=1.56 $Y=1.93 $X2=0 $Y2=0
cc_97 N_A_85_21#_c_91_n N_D1_c_175_n 0.00102134f $X=1.645 $Y=0.81 $X2=0 $Y2=0
cc_98 N_A_85_21#_M1010_g N_D1_c_176_n 0.0137032f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_85_21#_c_89_n N_D1_c_176_n 0.00405827f $X=1.56 $Y=1.93 $X2=0 $Y2=0
cc_100 N_A_85_21#_c_91_n N_D1_c_176_n 0.0010066f $X=1.645 $Y=0.81 $X2=0 $Y2=0
cc_101 N_A_85_21#_M1010_g N_D1_c_179_n 0.00147247f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A_85_21#_c_85_n N_D1_c_179_n 5.9921e-19 $X=0.59 $Y=1.975 $X2=0 $Y2=0
cc_103 N_A_85_21#_c_86_n N_D1_c_179_n 0.0132744f $X=0.59 $Y=1.635 $X2=0 $Y2=0
cc_104 N_A_85_21#_c_87_n N_D1_c_179_n 7.91268e-19 $X=0.59 $Y=1.635 $X2=0 $Y2=0
cc_105 N_A_85_21#_c_96_n N_D1_c_179_n 0.0235874f $X=1.475 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_85_21#_c_89_n N_D1_c_179_n 0.0470439f $X=1.56 $Y=1.93 $X2=0 $Y2=0
cc_107 N_A_85_21#_c_91_n N_D1_c_179_n 0.00239462f $X=1.645 $Y=0.81 $X2=0 $Y2=0
cc_108 N_A_85_21#_c_88_n N_C1_M1006_g 9.56501e-19 $X=1.365 $Y=0.51 $X2=0 $Y2=0
cc_109 N_A_85_21#_c_89_n N_C1_M1006_g 0.00764879f $X=1.56 $Y=1.93 $X2=0 $Y2=0
cc_110 N_A_85_21#_c_90_n N_C1_M1006_g 0.00272839f $X=2.12 $Y=0.81 $X2=0 $Y2=0
cc_111 N_A_85_21#_c_91_n N_C1_M1006_g 0.00778708f $X=1.645 $Y=0.81 $X2=0 $Y2=0
cc_112 N_A_85_21#_c_96_n N_C1_M1003_g 0.00773951f $X=1.475 $Y=2.035 $X2=0 $Y2=0
cc_113 N_A_85_21#_c_89_n N_C1_M1003_g 0.0160367f $X=1.56 $Y=1.93 $X2=0 $Y2=0
cc_114 N_A_85_21#_c_89_n N_C1_c_220_n 0.0052523f $X=1.56 $Y=1.93 $X2=0 $Y2=0
cc_115 N_A_85_21#_c_90_n N_C1_c_220_n 0.00152366f $X=2.12 $Y=0.81 $X2=0 $Y2=0
cc_116 N_A_85_21#_M1007_g N_C1_c_222_n 0.00419977f $X=0.5 $Y=2.745 $X2=0 $Y2=0
cc_117 N_A_85_21#_c_96_n N_C1_c_222_n 0.00435106f $X=1.475 $Y=2.035 $X2=0 $Y2=0
cc_118 N_A_85_21#_M1007_g C1 0.0047909f $X=0.5 $Y=2.745 $X2=0 $Y2=0
cc_119 N_A_85_21#_c_96_n C1 0.0233089f $X=1.475 $Y=2.035 $X2=0 $Y2=0
cc_120 N_A_85_21#_c_96_n N_B1_M1008_g 6.80947e-19 $X=1.475 $Y=2.035 $X2=0 $Y2=0
cc_121 N_A_85_21#_c_89_n N_B1_M1009_g 0.00410951f $X=1.56 $Y=1.93 $X2=0 $Y2=0
cc_122 N_A_85_21#_c_90_n N_B1_M1009_g 0.0163548f $X=2.12 $Y=0.81 $X2=0 $Y2=0
cc_123 N_A_85_21#_c_92_n N_B1_M1009_g 9.4709e-19 $X=2.225 $Y=0.51 $X2=0 $Y2=0
cc_124 N_A_85_21#_c_89_n N_B1_c_266_n 0.00117316f $X=1.56 $Y=1.93 $X2=0 $Y2=0
cc_125 N_A_85_21#_c_90_n N_B1_c_266_n 7.29492e-19 $X=2.12 $Y=0.81 $X2=0 $Y2=0
cc_126 N_A_85_21#_c_96_n B1 0.0100199f $X=1.475 $Y=2.035 $X2=0 $Y2=0
cc_127 N_A_85_21#_c_90_n N_A1_M1000_g 0.0042793f $X=2.12 $Y=0.81 $X2=0 $Y2=0
cc_128 N_A_85_21#_c_92_n N_A1_M1000_g 0.0017418f $X=2.225 $Y=0.51 $X2=0 $Y2=0
cc_129 N_A_85_21#_c_90_n A2 0.00413071f $X=2.12 $Y=0.81 $X2=0 $Y2=0
cc_130 N_A_85_21#_M1010_g X 8.03018e-19 $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_85_21#_M1010_g X 0.0537766f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A_85_21#_c_86_n X 0.0314501f $X=0.59 $Y=1.635 $X2=0 $Y2=0
cc_133 N_A_85_21#_c_97_n X 0.0160262f $X=0.675 $Y=2.035 $X2=0 $Y2=0
cc_134 N_A_85_21#_M1007_g N_VPWR_c_412_n 0.00513407f $X=0.5 $Y=2.745 $X2=0 $Y2=0
cc_135 N_A_85_21#_c_95_n N_VPWR_c_412_n 0.00202498f $X=0.59 $Y=2.14 $X2=0 $Y2=0
cc_136 N_A_85_21#_c_96_n N_VPWR_c_412_n 0.0051887f $X=1.475 $Y=2.035 $X2=0 $Y2=0
cc_137 N_A_85_21#_c_97_n N_VPWR_c_412_n 0.00196512f $X=0.675 $Y=2.035 $X2=0
+ $Y2=0
cc_138 N_A_85_21#_M1007_g N_VPWR_c_418_n 0.00457417f $X=0.5 $Y=2.745 $X2=0 $Y2=0
cc_139 N_A_85_21#_M1007_g N_VPWR_c_411_n 0.00544287f $X=0.5 $Y=2.745 $X2=0 $Y2=0
cc_140 N_A_85_21#_c_96_n A_267_369# 0.00471742f $X=1.475 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A_85_21#_c_89_n A_267_369# 9.56317e-19 $X=1.56 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_85_21#_c_89_n N_A_411_369#_c_473_n 0.00374237f $X=1.56 $Y=1.93 $X2=0
+ $Y2=0
cc_143 N_A_85_21#_c_89_n N_A_411_369#_c_471_n 0.00668349f $X=1.56 $Y=1.93 $X2=0
+ $Y2=0
cc_144 N_A_85_21#_M1010_g N_VGND_c_500_n 0.0102261f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_145 N_A_85_21#_c_90_n N_VGND_c_501_n 0.0139569f $X=2.12 $Y=0.81 $X2=0 $Y2=0
cc_146 N_A_85_21#_c_88_n N_VGND_c_504_n 0.00805099f $X=1.365 $Y=0.51 $X2=0 $Y2=0
cc_147 N_A_85_21#_c_91_n N_VGND_c_504_n 0.00308568f $X=1.645 $Y=0.81 $X2=0 $Y2=0
cc_148 N_A_85_21#_M1010_g N_VGND_c_506_n 0.00564095f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_85_21#_c_90_n N_VGND_c_507_n 0.00305343f $X=2.12 $Y=0.81 $X2=0 $Y2=0
cc_150 N_A_85_21#_c_92_n N_VGND_c_507_n 0.008231f $X=2.225 $Y=0.51 $X2=0 $Y2=0
cc_151 N_A_85_21#_M1001_d N_VGND_c_509_n 0.00370075f $X=1.225 $Y=0.235 $X2=0
+ $Y2=0
cc_152 N_A_85_21#_M1009_d N_VGND_c_509_n 0.00373063f $X=2.085 $Y=0.235 $X2=0
+ $Y2=0
cc_153 N_A_85_21#_M1010_g N_VGND_c_509_n 0.0106196f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_154 N_A_85_21#_c_88_n N_VGND_c_509_n 0.00756149f $X=1.365 $Y=0.51 $X2=0 $Y2=0
cc_155 N_A_85_21#_c_90_n N_VGND_c_509_n 0.00588128f $X=2.12 $Y=0.81 $X2=0 $Y2=0
cc_156 N_A_85_21#_c_91_n N_VGND_c_509_n 0.00512145f $X=1.645 $Y=0.81 $X2=0 $Y2=0
cc_157 N_A_85_21#_c_92_n N_VGND_c_509_n 0.00765087f $X=2.225 $Y=0.51 $X2=0 $Y2=0
cc_158 N_D1_M1001_g N_C1_M1006_g 0.0242176f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_159 N_D1_c_176_n N_C1_M1006_g 0.00870327f $X=1.13 $Y=1.18 $X2=0 $Y2=0
cc_160 N_D1_c_179_n N_C1_M1006_g 2.37143e-19 $X=1.13 $Y=1.18 $X2=0 $Y2=0
cc_161 N_D1_c_174_n N_C1_M1003_g 0.0119149f $X=1.15 $Y=1.535 $X2=0 $Y2=0
cc_162 N_D1_c_175_n N_C1_M1003_g 0.0535184f $X=1.15 $Y=1.685 $X2=0 $Y2=0
cc_163 N_D1_c_179_n N_C1_M1003_g 4.91642e-19 $X=1.13 $Y=1.18 $X2=0 $Y2=0
cc_164 N_D1_c_174_n N_C1_c_220_n 0.00870327f $X=1.15 $Y=1.535 $X2=0 $Y2=0
cc_165 N_D1_M1011_g N_C1_c_222_n 0.00834678f $X=1.26 $Y=2.055 $X2=0 $Y2=0
cc_166 N_D1_M1011_g C1 0.00603083f $X=1.26 $Y=2.055 $X2=0 $Y2=0
cc_167 N_D1_M1011_g B1 3.78935e-19 $X=1.26 $Y=2.055 $X2=0 $Y2=0
cc_168 N_D1_c_179_n X 0.0101548f $X=1.13 $Y=1.18 $X2=0 $Y2=0
cc_169 N_D1_M1001_g N_VGND_c_500_n 0.00666961f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_170 N_D1_M1001_g N_VGND_c_504_n 0.00585385f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_171 N_D1_M1001_g N_VGND_c_509_n 0.0115097f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_172 N_C1_c_222_n N_B1_M1008_g 0.0413373f $X=1.545 $Y=2.8 $X2=0 $Y2=0
cc_173 N_C1_M1006_g N_B1_M1009_g 0.0315403f $X=1.58 $Y=0.445 $X2=0 $Y2=0
cc_174 N_C1_c_220_n N_B1_M1009_g 0.0232826f $X=1.6 $Y=1.295 $X2=0 $Y2=0
cc_175 N_C1_M1003_g N_B1_c_266_n 0.0413373f $X=1.62 $Y=2.055 $X2=0 $Y2=0
cc_176 N_C1_M1003_g B1 0.0133299f $X=1.62 $Y=2.055 $X2=0 $Y2=0
cc_177 N_C1_c_222_n B1 0.00439543f $X=1.545 $Y=2.8 $X2=0 $Y2=0
cc_178 C1 B1 0.0328329f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_179 N_C1_c_222_n N_B1_c_272_n 0.0127802f $X=1.545 $Y=2.8 $X2=0 $Y2=0
cc_180 C1 N_B1_c_272_n 0.018338f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_181 C1 X 0.00626066f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_182 C1 X 0.00198529f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_183 N_C1_c_222_n N_VPWR_c_412_n 0.00290028f $X=1.545 $Y=2.8 $X2=0 $Y2=0
cc_184 C1 N_VPWR_c_412_n 0.022979f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_185 N_C1_c_222_n N_VPWR_c_416_n 0.00777516f $X=1.545 $Y=2.8 $X2=0 $Y2=0
cc_186 C1 N_VPWR_c_416_n 0.0128005f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_187 N_C1_c_222_n N_VPWR_c_411_n 0.00515305f $X=1.545 $Y=2.8 $X2=0 $Y2=0
cc_188 C1 N_VPWR_c_411_n 0.0117057f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_189 N_C1_M1006_g N_VGND_c_501_n 0.00288714f $X=1.58 $Y=0.445 $X2=0 $Y2=0
cc_190 N_C1_M1006_g N_VGND_c_504_n 0.00437852f $X=1.58 $Y=0.445 $X2=0 $Y2=0
cc_191 N_C1_M1006_g N_VGND_c_509_n 0.00604796f $X=1.58 $Y=0.445 $X2=0 $Y2=0
cc_192 N_B1_M1008_g N_A1_M1005_g 0.0197742f $X=1.98 $Y=2.055 $X2=0 $Y2=0
cc_193 N_B1_c_266_n N_A1_M1005_g 0.00630693f $X=1.995 $Y=1.735 $X2=0 $Y2=0
cc_194 N_B1_M1009_g N_A1_M1000_g 0.0472357f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_195 N_B1_M1008_g N_A1_c_320_n 0.00548026f $X=1.98 $Y=2.055 $X2=0 $Y2=0
cc_196 N_B1_c_270_n N_A1_c_320_n 0.00943165f $X=2.07 $Y=2.9 $X2=0 $Y2=0
cc_197 N_B1_M1009_g N_A1_c_318_n 0.00630693f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_198 N_B1_M1008_g N_VPWR_c_413_n 0.00197548f $X=1.98 $Y=2.055 $X2=0 $Y2=0
cc_199 B1 N_VPWR_c_413_n 0.00788678f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_200 N_B1_c_270_n N_VPWR_c_413_n 0.00375554f $X=2.07 $Y=2.9 $X2=0 $Y2=0
cc_201 N_B1_c_271_n N_VPWR_c_413_n 0.0263906f $X=2.07 $Y=2.9 $X2=0 $Y2=0
cc_202 N_B1_M1008_g N_VPWR_c_415_n 7.58114e-19 $X=1.98 $Y=2.055 $X2=0 $Y2=0
cc_203 B1 N_VPWR_c_415_n 0.00539659f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_204 N_B1_c_270_n N_VPWR_c_416_n 0.00852872f $X=2.07 $Y=2.9 $X2=0 $Y2=0
cc_205 N_B1_c_271_n N_VPWR_c_416_n 0.024867f $X=2.07 $Y=2.9 $X2=0 $Y2=0
cc_206 N_B1_c_272_n N_VPWR_c_416_n 0.0178675f $X=1.632 $Y=2.735 $X2=0 $Y2=0
cc_207 N_B1_c_270_n N_VPWR_c_411_n 0.0111008f $X=2.07 $Y=2.9 $X2=0 $Y2=0
cc_208 N_B1_c_271_n N_VPWR_c_411_n 0.0152046f $X=2.07 $Y=2.9 $X2=0 $Y2=0
cc_209 N_B1_c_272_n N_VPWR_c_411_n 0.0102537f $X=1.632 $Y=2.735 $X2=0 $Y2=0
cc_210 N_B1_M1008_g N_A_411_369#_c_473_n 7.84892e-19 $X=1.98 $Y=2.055 $X2=0
+ $Y2=0
cc_211 N_B1_c_270_n N_A_411_369#_c_473_n 0.00304132f $X=2.07 $Y=2.9 $X2=0 $Y2=0
cc_212 N_B1_c_271_n N_A_411_369#_c_473_n 0.00202022f $X=2.07 $Y=2.9 $X2=0 $Y2=0
cc_213 N_B1_M1008_g N_A_411_369#_c_471_n 5.4461e-19 $X=1.98 $Y=2.055 $X2=0 $Y2=0
cc_214 N_B1_c_266_n N_A_411_369#_c_471_n 0.00186347f $X=1.995 $Y=1.735 $X2=0
+ $Y2=0
cc_215 N_B1_M1009_g N_VGND_c_501_n 0.00288714f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_216 N_B1_M1009_g N_VGND_c_507_n 0.00437852f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_217 N_B1_M1009_g N_VGND_c_509_n 0.00604796f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_218 N_A1_M1005_g N_A2_M1004_g 0.0140324f $X=2.41 $Y=2.055 $X2=0 $Y2=0
cc_219 N_A1_M1000_g N_A2_M1004_g 0.00969976f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A1_c_320_n N_A2_M1004_g 0.00752517f $X=2.52 $Y=2.665 $X2=0 $Y2=0
cc_221 N_A1_c_321_n N_A2_M1004_g 0.00117059f $X=2.52 $Y=2.45 $X2=0 $Y2=0
cc_222 A1 N_A2_M1004_g 0.00464826f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_223 A1 N_A2_M1004_g 6.97298e-19 $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_224 N_A1_M1000_g N_A2_c_366_n 0.0813918f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A1_M1000_g A2 0.0152643f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_226 N_A1_c_320_n N_VPWR_c_413_n 0.0116238f $X=2.52 $Y=2.665 $X2=0 $Y2=0
cc_227 N_A1_c_321_n N_VPWR_c_413_n 0.00446653f $X=2.52 $Y=2.45 $X2=0 $Y2=0
cc_228 A1 N_VPWR_c_413_n 0.00734934f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_229 A1 N_VPWR_c_413_n 0.025245f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_230 N_A1_M1005_g N_VPWR_c_414_n 0.0010012f $X=2.41 $Y=2.055 $X2=0 $Y2=0
cc_231 N_A1_c_321_n N_VPWR_c_414_n 5.78451e-19 $X=2.52 $Y=2.45 $X2=0 $Y2=0
cc_232 N_A1_M1005_g N_VPWR_c_415_n 0.00620255f $X=2.41 $Y=2.055 $X2=0 $Y2=0
cc_233 N_A1_c_320_n N_VPWR_c_415_n 0.00413331f $X=2.52 $Y=2.665 $X2=0 $Y2=0
cc_234 N_A1_c_321_n N_VPWR_c_415_n 0.00983465f $X=2.52 $Y=2.45 $X2=0 $Y2=0
cc_235 A1 N_VPWR_c_415_n 0.0137383f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_236 A1 N_VPWR_c_415_n 7.38584e-19 $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_237 N_A1_c_320_n N_VPWR_c_419_n 0.00972723f $X=2.52 $Y=2.665 $X2=0 $Y2=0
cc_238 A1 N_VPWR_c_419_n 0.0219703f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_239 N_A1_c_320_n N_VPWR_c_411_n 0.0125687f $X=2.52 $Y=2.665 $X2=0 $Y2=0
cc_240 A1 N_VPWR_c_411_n 0.0181915f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_241 N_A1_M1005_g N_A_411_369#_c_473_n 9.32559e-19 $X=2.41 $Y=2.055 $X2=0
+ $Y2=0
cc_242 N_A1_M1005_g N_A_411_369#_c_470_n 0.00890337f $X=2.41 $Y=2.055 $X2=0
+ $Y2=0
cc_243 N_A1_c_318_n N_A_411_369#_c_470_n 0.00938333f $X=2.425 $Y=1.635 $X2=0
+ $Y2=0
cc_244 N_A1_c_321_n N_A_411_369#_c_470_n 2.4916e-19 $X=2.52 $Y=2.45 $X2=0 $Y2=0
cc_245 A1 N_A_411_369#_c_470_n 0.00107699f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_246 N_A1_M1005_g N_A_411_369#_c_472_n 6.02135e-19 $X=2.41 $Y=2.055 $X2=0
+ $Y2=0
cc_247 A1 N_A_411_369#_c_472_n 0.0167974f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_248 N_A1_M1000_g N_VGND_c_503_n 0.00207709f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_249 N_A1_M1000_g N_VGND_c_507_n 0.00585385f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_250 N_A1_M1000_g N_VGND_c_509_n 0.0108402f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_251 N_A2_M1004_g N_VPWR_c_414_n 0.00469177f $X=2.88 $Y=2.055 $X2=0 $Y2=0
cc_252 N_A2_M1004_g N_VPWR_c_415_n 9.18177e-19 $X=2.88 $Y=2.055 $X2=0 $Y2=0
cc_253 N_A2_M1004_g N_A_411_369#_c_470_n 0.0113212f $X=2.88 $Y=2.055 $X2=0 $Y2=0
cc_254 N_A2_c_368_n N_A_411_369#_c_470_n 0.00216013f $X=2.89 $Y=1.435 $X2=0
+ $Y2=0
cc_255 A2 N_A_411_369#_c_470_n 0.0240185f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_256 N_A2_M1004_g N_A_411_369#_c_472_n 0.0114726f $X=2.88 $Y=2.055 $X2=0 $Y2=0
cc_257 N_A2_c_368_n N_A_411_369#_c_472_n 0.00274105f $X=2.89 $Y=1.435 $X2=0
+ $Y2=0
cc_258 A2 N_A_411_369#_c_472_n 0.0194534f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_259 N_A2_c_366_n N_VGND_c_503_n 0.0106506f $X=2.89 $Y=0.765 $X2=0 $Y2=0
cc_260 A2 N_VGND_c_503_n 0.0129339f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_261 N_A2_c_370_n N_VGND_c_503_n 0.00439657f $X=2.89 $Y=0.93 $X2=0 $Y2=0
cc_262 N_A2_c_366_n N_VGND_c_507_n 0.00486043f $X=2.89 $Y=0.765 $X2=0 $Y2=0
cc_263 N_A2_c_366_n N_VGND_c_509_n 0.00445138f $X=2.89 $Y=0.765 $X2=0 $Y2=0
cc_264 A2 N_VGND_c_509_n 0.0130291f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_265 X N_VPWR_c_418_n 0.00640351f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_266 X N_VPWR_c_411_n 0.00789919f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_267 X N_VGND_c_506_n 0.00980051f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_268 N_X_M1010_s N_VGND_c_509_n 0.0034811f $X=0.16 $Y=0.235 $X2=0 $Y2=0
cc_269 X N_VGND_c_509_n 0.00857705f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_270 N_VPWR_c_414_n N_A_411_369#_c_470_n 0.0133334f $X=2.625 $Y=2.12 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_415_n N_A_411_369#_c_470_n 0.00518537f $X=2.615 $Y=2.4 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_414_n N_A_411_369#_c_472_n 0.00854666f $X=2.625 $Y=2.12 $X2=0
+ $Y2=0
cc_273 N_VGND_c_509_n A_503_47# 0.00420785f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
