* File: sky130_fd_sc_lp__o32a_0.spice
* Created: Fri Aug 28 11:17:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32a_0.pex.spice"
.subckt sky130_fd_sc_lp__o32a_0  VNB VPB A1 A2 A3 B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_97_309#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.1113 PD=0.84 PS=1.37 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1005 N_A_271_85#_M1005_d N_A1_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.8
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_271_85#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.105 AS=0.0588 PD=0.92 PS=0.7 NRD=31.428 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 N_A_271_85#_M1001_d N_A3_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.105 PD=0.7 PS=0.92 NRD=0 NRS=31.428 M=1 R=2.8 SA=75001.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_A_97_309#_M1007_d N_B2_M1007_g N_A_271_85#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_A_271_85#_M1006_d N_B1_M1006_g N_A_97_309#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1218 AS=0.0735 PD=1.42 PS=0.77 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_97_309#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1728 AS=0.1696 PD=1.18 PS=1.81 NRD=40.0107 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1003 A_301_481# N_A1_M1003_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1728 PD=0.88 PS=1.18 NRD=19.9955 NRS=40.0107 M=1 R=4.26667
+ SA=75000.9 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1009 A_379_481# N_A2_M1009_g A_301_481# VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0768 PD=0.88 PS=0.88 NRD=19.9955 NRS=19.9955 M=1 R=4.26667 SA=75001.3
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1002 N_A_97_309#_M1002_d N_A3_M1002_g A_379_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1152 AS=0.0768 PD=1 PS=0.88 NRD=12.2928 NRS=19.9955 M=1 R=4.26667
+ SA=75001.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 A_559_481# N_B2_M1004_g N_A_97_309#_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1152 PD=0.88 PS=1 NRD=19.9955 NRS=12.2928 M=1 R=4.26667
+ SA=75002.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_B1_M1008_g A_559_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75002.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o32a_0.pxi.spice"
*
.ends
*
*
