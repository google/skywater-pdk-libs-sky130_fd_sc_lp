/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_LP__ISO0P_TB_V
`define SKY130_FD_SC_LP__ISO0P_TB_V

/**
 * iso0p: ????.
 *
 * Autogenerated test bench.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

`include "sky130_fd_sc_lp__iso0p.v"

module top();

    // Inputs are registered
    reg A;
    reg SLEEP;
    reg KAPWR;
    reg VGND;
    reg VPB;
    reg VNB;

    // Outputs are wires
    wire X;

    initial
    begin
        // Initial state is x for all inputs.
        A     = 1'bX;
        KAPWR = 1'bX;
        SLEEP = 1'bX;
        VGND  = 1'bX;
        VNB   = 1'bX;
        VPB   = 1'bX;

        #20   A     = 1'b0;
        #40   KAPWR = 1'b0;
        #60   SLEEP = 1'b0;
        #80   VGND  = 1'b0;
        #100  VNB   = 1'b0;
        #120  VPB   = 1'b0;
        #140  A     = 1'b1;
        #160  KAPWR = 1'b1;
        #180  SLEEP = 1'b1;
        #200  VGND  = 1'b1;
        #220  VNB   = 1'b1;
        #240  VPB   = 1'b1;
        #260  A     = 1'b0;
        #280  KAPWR = 1'b0;
        #300  SLEEP = 1'b0;
        #320  VGND  = 1'b0;
        #340  VNB   = 1'b0;
        #360  VPB   = 1'b0;
        #380  VPB   = 1'b1;
        #400  VNB   = 1'b1;
        #420  VGND  = 1'b1;
        #440  SLEEP = 1'b1;
        #460  KAPWR = 1'b1;
        #480  A     = 1'b1;
        #500  VPB   = 1'bx;
        #520  VNB   = 1'bx;
        #540  VGND  = 1'bx;
        #560  SLEEP = 1'bx;
        #580  KAPWR = 1'bx;
        #600  A     = 1'bx;
    end

    sky130_fd_sc_lp__iso0p dut (.A(A), .SLEEP(SLEEP), .KAPWR(KAPWR), .VGND(VGND), .VPB(VPB), .VNB(VNB), .X(X));

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_LP__ISO0P_TB_V
