* NGSPICE file created from sky130_fd_sc_lp__srsdfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__srsdfxtp_1 CLK D SCD SCE SLEEP_B KAPWR VGND VNB VPB VPWR
+ Q
M1000 a_204_477# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.52888e+12p ps=1.147e+07u
M1001 a_1858_419# a_570_47# a_1319_69# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=5.244e+11p ps=4.82e+06u
M1002 a_2321_178# SLEEP_B a_2243_178# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.008e+11p ps=1.32e+06u
M1003 a_282_477# D a_210_47# VNB nshort w=420000u l=150000u
+  ad=2.835e+11p pd=3.03e+06u as=1.008e+11p ps=1.32e+06u
M1004 a_368_477# a_31_477# a_282_477# VPB phighvt w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=3.283e+11p ps=3.39e+06u
M1005 a_786_139# a_540_21# a_282_477# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1006 VGND a_1493_21# a_1523_113# VNB nshort w=420000u l=150000u
+  ad=1.3371e+12p pd=1.18e+07u as=8.82e+10p ps=1.26e+06u
M1007 a_1493_21# a_1319_69# a_1704_125# VNB nshort w=420000u l=150000u
+  ad=1.738e+11p pd=1.68e+06u as=8.82e+10p ps=1.26e+06u
M1008 a_872_139# a_570_47# a_786_139# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 a_1372_379# a_540_21# a_914_245# VPB phighvt w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=3.346e+11p ps=2.86e+06u
M1010 a_540_21# SLEEP_B KAPWR VPB phighvt w=640000u l=150000u
+  ad=3.52e+11p pd=2.38e+06u as=7.108e+11p ps=5.58e+06u
M1011 VPWR a_1319_69# a_2504_57# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1012 a_1319_69# a_570_47# a_1247_69# VNB nshort w=640000u l=150000u
+  ad=3.099e+11p pd=2.3e+06u as=1.344e+11p ps=1.7e+06u
M1013 a_2243_178# CLK a_540_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.68e+11p ps=1.64e+06u
M1014 a_1319_69# a_540_21# a_1372_379# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 KAPWR CLK a_540_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND SCD a_396_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1017 KAPWR a_1493_21# a_1858_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_396_47# SCE a_282_477# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1523_113# a_1493_21# a_1451_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1020 a_1704_125# a_1319_69# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_282_477# D a_204_477# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1010_530# a_540_21# a_786_139# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.176e+11p ps=1.4e+06u
M1023 a_914_245# a_786_139# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Q a_2504_57# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1025 a_570_47# a_540_21# VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1026 a_1451_113# a_540_21# a_1319_69# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_570_47# a_540_21# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1028 a_1247_69# a_570_47# a_914_245# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.392e+11p ps=2.34e+06u
M1029 a_1493_21# a_1319_69# KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=4.35e+11p pd=2.87e+06u as=0p ps=0u
M1030 VPWR SCE a_31_477# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1031 Q a_2504_57# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1032 VGND a_1319_69# a_2504_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1033 VGND SLEEP_B a_2321_178# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_914_245# a_872_139# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_786_139# a_570_47# a_282_477# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_914_245# a_1010_530# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_210_47# a_31_477# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_914_245# a_786_139# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR SCD a_368_477# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND SCE a_31_477# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends

