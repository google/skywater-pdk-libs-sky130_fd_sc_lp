* File: sky130_fd_sc_lp__o41ai_m.spice
* Created: Fri Aug 28 11:20:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41ai_m.pex.spice"
.subckt sky130_fd_sc_lp__o41ai_m  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_A_175_47#_M1006_d N_B1_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.2058 PD=0.755 PS=1.82 NRD=15.708 NRS=64.284 M=1 R=2.8
+ SA=75000.4 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A4_M1004_g N_A_175_47#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07875 AS=0.07035 PD=0.795 PS=0.755 NRD=0 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_175_47#_M1007_d N_A3_M1007_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.07875 PD=0.7 PS=0.795 NRD=0 NRS=27.132 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_175_47#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.0588 PD=0.72 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_175_47#_M1002_d N_A1_M1002_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.063 PD=1.37 PS=0.72 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09555 AS=0.1113 PD=0.875 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1005 A_247_371# N_A4_M1005_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.09555 PD=0.81 PS=0.875 NRD=65.6601 NRS=82.0702 M=1 R=2.8 SA=75000.8
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 A_355_371# N_A3_M1008_g A_247_371# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0819 PD=0.81 PS=0.81 NRD=65.6601 NRS=65.6601 M=1 R=2.8 SA=75001.3
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_463_371# N_A2_M1001_g A_355_371# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=65.6601 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g A_463_371# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_43 VNB 0 2.89541e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o41ai_m.pxi.spice"
*
.ends
*
*
