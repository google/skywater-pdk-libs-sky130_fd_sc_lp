* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
M1000 X a_79_47# a_283_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=6.174e+11p pd=3.5e+06u as=2.646e+11p ps=2.94e+06u
M1001 VGND a_79_47# X VNB nshort w=840000u l=150000u
+  ad=5.334e+11p pd=4.8e+06u as=2.352e+11p ps=2.24e+06u
M1002 VGND A a_79_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 VPWR A a_79_47# VPB phighvt w=420000u l=150000u
+  ad=3.864e+11p pd=3.3e+06u as=1.113e+11p ps=1.37e+06u
M1004 X SLEEP VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_283_367# SLEEP VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
