* File: sky130_fd_sc_lp__a21bo_1.pxi.spice
* Created: Fri Aug 28 09:49:09 2020
* 
x_PM_SKY130_FD_SC_LP__A21BO_1%A_80_43# N_A_80_43#_M1007_d N_A_80_43#_M1001_s
+ N_A_80_43#_M1005_g N_A_80_43#_M1009_g N_A_80_43#_c_76_n N_A_80_43#_c_70_n
+ N_A_80_43#_c_140_p N_A_80_43#_c_77_n N_A_80_43#_c_128_p N_A_80_43#_c_81_p
+ N_A_80_43#_c_96_p N_A_80_43#_c_71_n N_A_80_43#_c_72_n N_A_80_43#_c_73_n
+ N_A_80_43#_c_78_n N_A_80_43#_c_97_p N_A_80_43#_c_74_n
+ PM_SKY130_FD_SC_LP__A21BO_1%A_80_43#
x_PM_SKY130_FD_SC_LP__A21BO_1%B1_N N_B1_N_M1006_g N_B1_N_M1002_g B1_N
+ N_B1_N_c_158_n N_B1_N_c_159_n PM_SKY130_FD_SC_LP__A21BO_1%B1_N
x_PM_SKY130_FD_SC_LP__A21BO_1%A_237_367# N_A_237_367#_M1002_d
+ N_A_237_367#_M1006_d N_A_237_367#_M1007_g N_A_237_367#_M1001_g
+ N_A_237_367#_c_194_n N_A_237_367#_c_195_n N_A_237_367#_c_202_n
+ N_A_237_367#_c_196_n N_A_237_367#_c_197_n N_A_237_367#_c_203_n
+ N_A_237_367#_c_198_n PM_SKY130_FD_SC_LP__A21BO_1%A_237_367#
x_PM_SKY130_FD_SC_LP__A21BO_1%A1 N_A1_M1004_g N_A1_M1003_g A1 A1 N_A1_c_260_n
+ N_A1_c_261_n PM_SKY130_FD_SC_LP__A21BO_1%A1
x_PM_SKY130_FD_SC_LP__A21BO_1%A2 N_A2_M1008_g N_A2_M1000_g A2 A2 N_A2_c_295_n
+ N_A2_c_296_n PM_SKY130_FD_SC_LP__A21BO_1%A2
x_PM_SKY130_FD_SC_LP__A21BO_1%X N_X_M1005_s N_X_M1009_s X X X X X X X
+ PM_SKY130_FD_SC_LP__A21BO_1%X
x_PM_SKY130_FD_SC_LP__A21BO_1%VPWR N_VPWR_M1009_d N_VPWR_M1004_d N_VPWR_c_335_n
+ N_VPWR_c_336_n VPWR N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n
+ N_VPWR_c_334_n N_VPWR_c_341_n N_VPWR_c_342_n PM_SKY130_FD_SC_LP__A21BO_1%VPWR
x_PM_SKY130_FD_SC_LP__A21BO_1%A_436_367# N_A_436_367#_M1001_d
+ N_A_436_367#_M1000_d N_A_436_367#_c_376_n N_A_436_367#_c_374_n
+ N_A_436_367#_c_375_n N_A_436_367#_c_379_n
+ PM_SKY130_FD_SC_LP__A21BO_1%A_436_367#
x_PM_SKY130_FD_SC_LP__A21BO_1%VGND N_VGND_M1005_d N_VGND_M1007_s N_VGND_M1008_d
+ N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n
+ VGND N_VGND_c_406_n N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n
+ N_VGND_c_410_n PM_SKY130_FD_SC_LP__A21BO_1%VGND
cc_1 VNB N_A_80_43#_M1009_g 0.00158724f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_2 VNB N_A_80_43#_c_70_n 0.0132213f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=0.72
cc_3 VNB N_A_80_43#_c_71_n 0.00618095f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.46
cc_4 VNB N_A_80_43#_c_72_n 0.0403779f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.46
cc_5 VNB N_A_80_43#_c_73_n 0.001861f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.295
cc_6 VNB N_A_80_43#_c_74_n 0.0223851f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.295
cc_7 VNB N_B1_N_M1002_g 0.0235217f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.295
cc_8 VNB N_B1_N_c_158_n 0.0253515f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_9 VNB N_B1_N_c_159_n 0.00347984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_237_367#_M1007_g 0.0295216f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_11 VNB N_A_237_367#_c_194_n 0.0288276f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_12 VNB N_A_237_367#_c_195_n 0.0102703f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.625
cc_13 VNB N_A_237_367#_c_196_n 0.00475267f $X=-0.19 $Y=-0.245 $X2=0.825
+ $Y2=2.405
cc_14 VNB N_A_237_367#_c_197_n 0.00380131f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=2.01
cc_15 VNB N_A_237_367#_c_198_n 0.00251304f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.46
cc_16 VNB N_A1_M1004_g 0.00775904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A1 0.00862464f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_18 VNB N_A1_c_260_n 0.0309452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_261_n 0.0173739f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_20 VNB N_A2_M1000_g 0.0113394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A2 0.0370818f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_22 VNB N_A2_c_295_n 0.0393572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_c_296_n 0.0207587f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_24 VNB X 0.0603078f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.295
cc_25 VNB N_VPWR_c_334_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.46
cc_26 VNB N_A_436_367#_c_374_n 0.0104065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_436_367#_c_375_n 0.00265307f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=0.805
cc_28 VNB N_VGND_c_401_n 0.0152316f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=0.805
cc_29 VNB N_VGND_c_402_n 0.0118704f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=0.72
cc_30 VNB N_VGND_c_403_n 0.0341176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_404_n 0.0206164f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=2.01
cc_32 VNB N_VGND_c_405_n 0.00510127f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=2.01
cc_33 VNB N_VGND_c_406_n 0.0276359f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.46
cc_34 VNB N_VGND_c_407_n 0.014713f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=0.72
cc_35 VNB N_VGND_c_408_n 0.235404f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=0.93
cc_36 VNB N_VGND_c_409_n 0.0265431f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.46
cc_37 VNB N_VGND_c_410_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_80_43#_M1009_g 0.0249101f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_39 VPB N_A_80_43#_c_76_n 0.00143034f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.32
cc_40 VPB N_A_80_43#_c_77_n 0.0240029f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=2.405
cc_41 VPB N_A_80_43#_c_78_n 0.0234191f $X=-0.19 $Y=1.655 $X2=1.89 $Y2=2.455
cc_42 VPB N_B1_N_M1006_g 0.0225045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_B1_N_c_158_n 0.00629975f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_44 VPB N_B1_N_c_159_n 0.00274851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_237_367#_M1001_g 0.0230427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_237_367#_c_194_n 0.0119686f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.295
cc_47 VPB N_A_237_367#_c_195_n 7.08598e-19 $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.625
cc_48 VPB N_A_237_367#_c_202_n 0.00508434f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.32
cc_49 VPB N_A_237_367#_c_203_n 0.00564892f $X=-0.19 $Y=1.655 $X2=2.41 $Y2=0.635
cc_50 VPB N_A_237_367#_c_198_n 7.78427e-19 $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.46
cc_51 VPB N_A1_M1004_g 0.0199258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A2_M1000_g 0.0248037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB X 0.00853703f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.295
cc_54 VPB X 0.010762f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_55 VPB X 0.0479783f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.46
cc_56 VPB N_VPWR_c_335_n 0.0198075f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_57 VPB N_VPWR_c_336_n 0.00561552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_337_n 0.0177474f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=0.72
cc_59 VPB N_VPWR_c_338_n 0.0478356f $X=-0.19 $Y=1.655 $X2=1.915 $Y2=2.32
cc_60 VPB N_VPWR_c_339_n 0.0277357f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_334_n 0.0701076f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.46
cc_62 VPB N_VPWR_c_341_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.295
cc_63 VPB N_VPWR_c_342_n 0.00632158f $X=-0.19 $Y=1.655 $X2=1.89 $Y2=2.455
cc_64 VPB N_A_436_367#_c_376_n 7.12009e-19 $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_65 VPB N_A_436_367#_c_374_n 0.0124832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_436_367#_c_375_n 0.0017297f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=0.805
cc_67 VPB N_A_436_367#_c_379_n 0.0465699f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.32
cc_68 N_A_80_43#_c_76_n N_B1_N_M1006_g 0.00784919f $X=0.74 $Y=2.32 $X2=0 $Y2=0
cc_69 N_A_80_43#_c_77_n N_B1_N_M1006_g 0.00950315f $X=1.725 $Y=2.405 $X2=0 $Y2=0
cc_70 N_A_80_43#_c_81_p N_B1_N_M1006_g 0.00302177f $X=1.89 $Y=2.01 $X2=0 $Y2=0
cc_71 N_A_80_43#_c_70_n N_B1_N_M1002_g 0.0147368f $X=2.245 $Y=0.72 $X2=0 $Y2=0
cc_72 N_A_80_43#_c_72_n N_B1_N_M1002_g 0.00220127f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_73 N_A_80_43#_c_73_n N_B1_N_M1002_g 0.00715125f $X=0.68 $Y=1.295 $X2=0 $Y2=0
cc_74 N_A_80_43#_c_74_n N_B1_N_M1002_g 0.00993804f $X=0.597 $Y=1.295 $X2=0 $Y2=0
cc_75 N_A_80_43#_M1009_g N_B1_N_c_158_n 0.0212911f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_76 N_A_80_43#_c_71_n N_B1_N_c_158_n 6.37069e-19 $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_77 N_A_80_43#_c_72_n N_B1_N_c_158_n 0.0154153f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_78 N_A_80_43#_M1009_g N_B1_N_c_159_n 3.18639e-19 $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_79 N_A_80_43#_c_70_n N_B1_N_c_159_n 0.00446217f $X=2.245 $Y=0.72 $X2=0 $Y2=0
cc_80 N_A_80_43#_c_77_n N_B1_N_c_159_n 0.00436934f $X=1.725 $Y=2.405 $X2=0 $Y2=0
cc_81 N_A_80_43#_c_71_n N_B1_N_c_159_n 0.031253f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_82 N_A_80_43#_c_72_n N_B1_N_c_159_n 8.69838e-19 $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_83 N_A_80_43#_c_70_n N_A_237_367#_M1002_d 0.00253998f $X=2.245 $Y=0.72
+ $X2=-0.19 $Y2=-0.245
cc_84 N_A_80_43#_c_70_n N_A_237_367#_M1007_g 0.0153202f $X=2.245 $Y=0.72 $X2=0
+ $Y2=0
cc_85 N_A_80_43#_c_96_p N_A_237_367#_M1007_g 0.00693908f $X=2.41 $Y=0.38 $X2=0
+ $Y2=0
cc_86 N_A_80_43#_c_97_p N_A_237_367#_M1007_g 0.00639508f $X=2.41 $Y=0.72 $X2=0
+ $Y2=0
cc_87 N_A_80_43#_c_70_n N_A_237_367#_c_194_n 0.00698832f $X=2.245 $Y=0.72 $X2=0
+ $Y2=0
cc_88 N_A_80_43#_c_77_n N_A_237_367#_c_194_n 0.00123673f $X=1.725 $Y=2.405 $X2=0
+ $Y2=0
cc_89 N_A_80_43#_c_81_p N_A_237_367#_c_194_n 0.00657241f $X=1.89 $Y=2.01 $X2=0
+ $Y2=0
cc_90 N_A_80_43#_c_78_n N_A_237_367#_c_194_n 0.00133906f $X=1.89 $Y=2.455 $X2=0
+ $Y2=0
cc_91 N_A_80_43#_c_76_n N_A_237_367#_c_202_n 0.00940273f $X=0.74 $Y=2.32 $X2=0
+ $Y2=0
cc_92 N_A_80_43#_c_77_n N_A_237_367#_c_202_n 0.033103f $X=1.725 $Y=2.405 $X2=0
+ $Y2=0
cc_93 N_A_80_43#_c_81_p N_A_237_367#_c_202_n 0.0172488f $X=1.89 $Y=2.01 $X2=0
+ $Y2=0
cc_94 N_A_80_43#_c_70_n N_A_237_367#_c_196_n 0.0297886f $X=2.245 $Y=0.72 $X2=0
+ $Y2=0
cc_95 N_A_80_43#_c_73_n N_A_237_367#_c_196_n 0.00842652f $X=0.68 $Y=1.295 $X2=0
+ $Y2=0
cc_96 N_A_80_43#_c_97_p N_A_237_367#_c_196_n 0.00215878f $X=2.41 $Y=0.72 $X2=0
+ $Y2=0
cc_97 N_A_80_43#_c_73_n N_A_237_367#_c_197_n 0.00503082f $X=0.68 $Y=1.295 $X2=0
+ $Y2=0
cc_98 N_A_80_43#_c_76_n N_A_237_367#_c_203_n 0.00517087f $X=0.74 $Y=2.32 $X2=0
+ $Y2=0
cc_99 N_A_80_43#_c_81_p N_A_237_367#_c_203_n 0.00637099f $X=1.89 $Y=2.01 $X2=0
+ $Y2=0
cc_100 N_A_80_43#_c_70_n N_A_237_367#_c_198_n 0.00805574f $X=2.245 $Y=0.72 $X2=0
+ $Y2=0
cc_101 N_A_80_43#_c_77_n N_A_237_367#_c_198_n 0.00250742f $X=1.725 $Y=2.405
+ $X2=0 $Y2=0
cc_102 N_A_80_43#_c_81_p N_A_237_367#_c_198_n 0.00734967f $X=1.89 $Y=2.01 $X2=0
+ $Y2=0
cc_103 N_A_80_43#_c_78_n N_A_237_367#_c_198_n 0.00238105f $X=1.89 $Y=2.455 $X2=0
+ $Y2=0
cc_104 N_A_80_43#_c_70_n A1 0.00522081f $X=2.245 $Y=0.72 $X2=0 $Y2=0
cc_105 N_A_80_43#_c_97_p A1 0.0273342f $X=2.41 $Y=0.72 $X2=0 $Y2=0
cc_106 N_A_80_43#_c_97_p N_A1_c_260_n 0.00343578f $X=2.41 $Y=0.72 $X2=0 $Y2=0
cc_107 N_A_80_43#_M1009_g X 0.0040734f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_80_43#_c_76_n X 0.00946825f $X=0.74 $Y=2.32 $X2=0 $Y2=0
cc_109 N_A_80_43#_c_71_n X 0.0255321f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_110 N_A_80_43#_c_73_n X 0.015163f $X=0.68 $Y=1.295 $X2=0 $Y2=0
cc_111 N_A_80_43#_c_74_n X 0.0154581f $X=0.597 $Y=1.295 $X2=0 $Y2=0
cc_112 N_A_80_43#_M1009_g X 0.00336422f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_80_43#_c_76_n X 0.0163712f $X=0.74 $Y=2.32 $X2=0 $Y2=0
cc_114 N_A_80_43#_c_72_n X 0.00303057f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_115 N_A_80_43#_c_76_n N_VPWR_M1009_d 0.00588397f $X=0.74 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A_80_43#_c_77_n N_VPWR_M1009_d 0.00495501f $X=1.725 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_80_43#_c_128_p N_VPWR_M1009_d 0.00116801f $X=0.825 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_80_43#_M1009_g N_VPWR_c_335_n 0.0142495f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_A_80_43#_c_77_n N_VPWR_c_335_n 0.0111448f $X=1.725 $Y=2.405 $X2=0 $Y2=0
cc_120 N_A_80_43#_c_128_p N_VPWR_c_335_n 0.00983065f $X=0.825 $Y=2.405 $X2=0
+ $Y2=0
cc_121 N_A_80_43#_M1009_g N_VPWR_c_337_n 0.00486043f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_A_80_43#_c_78_n N_VPWR_c_338_n 0.0192303f $X=1.89 $Y=2.455 $X2=0 $Y2=0
cc_123 N_A_80_43#_M1001_s N_VPWR_c_334_n 0.00232552f $X=1.765 $Y=1.835 $X2=0
+ $Y2=0
cc_124 N_A_80_43#_M1009_g N_VPWR_c_334_n 0.00926856f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_80_43#_c_77_n N_VPWR_c_334_n 0.0267261f $X=1.725 $Y=2.405 $X2=0 $Y2=0
cc_126 N_A_80_43#_c_128_p N_VPWR_c_334_n 6.15123e-19 $X=0.825 $Y=2.405 $X2=0
+ $Y2=0
cc_127 N_A_80_43#_c_78_n N_VPWR_c_334_n 0.0115856f $X=1.89 $Y=2.455 $X2=0 $Y2=0
cc_128 N_A_80_43#_c_70_n N_VGND_M1005_d 0.0085226f $X=2.245 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_80_43#_c_140_p N_VGND_M1005_d 0.00521432f $X=0.825 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_130 N_A_80_43#_c_73_n N_VGND_M1005_d 0.011267f $X=0.68 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_80_43#_c_70_n N_VGND_M1007_s 0.00624226f $X=2.245 $Y=0.72 $X2=0 $Y2=0
cc_132 N_A_80_43#_c_70_n N_VGND_c_401_n 0.0110001f $X=2.245 $Y=0.72 $X2=0 $Y2=0
cc_133 N_A_80_43#_c_140_p N_VGND_c_401_n 0.0143137f $X=0.825 $Y=0.72 $X2=0 $Y2=0
cc_134 N_A_80_43#_c_74_n N_VGND_c_401_n 0.00744387f $X=0.597 $Y=1.295 $X2=0
+ $Y2=0
cc_135 N_A_80_43#_c_70_n N_VGND_c_402_n 0.0206145f $X=2.245 $Y=0.72 $X2=0 $Y2=0
cc_136 N_A_80_43#_c_96_p N_VGND_c_402_n 0.0149618f $X=2.41 $Y=0.38 $X2=0 $Y2=0
cc_137 N_A_80_43#_c_70_n N_VGND_c_404_n 0.0134614f $X=2.245 $Y=0.72 $X2=0 $Y2=0
cc_138 N_A_80_43#_c_70_n N_VGND_c_406_n 0.00272902f $X=2.245 $Y=0.72 $X2=0 $Y2=0
cc_139 N_A_80_43#_c_96_p N_VGND_c_406_n 0.0230277f $X=2.41 $Y=0.38 $X2=0 $Y2=0
cc_140 N_A_80_43#_M1007_d N_VGND_c_408_n 0.00582224f $X=2.18 $Y=0.235 $X2=0
+ $Y2=0
cc_141 N_A_80_43#_c_70_n N_VGND_c_408_n 0.028435f $X=2.245 $Y=0.72 $X2=0 $Y2=0
cc_142 N_A_80_43#_c_140_p N_VGND_c_408_n 8.64211e-19 $X=0.825 $Y=0.72 $X2=0
+ $Y2=0
cc_143 N_A_80_43#_c_96_p N_VGND_c_408_n 0.0127466f $X=2.41 $Y=0.38 $X2=0 $Y2=0
cc_144 N_A_80_43#_c_74_n N_VGND_c_408_n 0.0100483f $X=0.597 $Y=1.295 $X2=0 $Y2=0
cc_145 N_A_80_43#_c_74_n N_VGND_c_409_n 0.00482246f $X=0.597 $Y=1.295 $X2=0
+ $Y2=0
cc_146 N_B1_N_c_158_n N_A_237_367#_c_194_n 0.014118f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_147 N_B1_N_c_159_n N_A_237_367#_c_194_n 2.74127e-19 $X=1.2 $Y=1.51 $X2=0
+ $Y2=0
cc_148 N_B1_N_M1006_g N_A_237_367#_c_202_n 0.0036177f $X=1.11 $Y=2.045 $X2=0
+ $Y2=0
cc_149 N_B1_N_c_158_n N_A_237_367#_c_202_n 0.00330087f $X=1.2 $Y=1.51 $X2=0
+ $Y2=0
cc_150 N_B1_N_c_159_n N_A_237_367#_c_202_n 0.00735337f $X=1.2 $Y=1.51 $X2=0
+ $Y2=0
cc_151 N_B1_N_M1002_g N_A_237_367#_c_196_n 0.00362675f $X=1.135 $Y=0.975 $X2=0
+ $Y2=0
cc_152 N_B1_N_c_158_n N_A_237_367#_c_196_n 0.00349522f $X=1.2 $Y=1.51 $X2=0
+ $Y2=0
cc_153 N_B1_N_c_159_n N_A_237_367#_c_196_n 0.00532736f $X=1.2 $Y=1.51 $X2=0
+ $Y2=0
cc_154 N_B1_N_M1002_g N_A_237_367#_c_197_n 0.00344926f $X=1.135 $Y=0.975 $X2=0
+ $Y2=0
cc_155 N_B1_N_M1006_g N_A_237_367#_c_203_n 0.00277072f $X=1.11 $Y=2.045 $X2=0
+ $Y2=0
cc_156 N_B1_N_c_159_n N_A_237_367#_c_203_n 0.00563737f $X=1.2 $Y=1.51 $X2=0
+ $Y2=0
cc_157 N_B1_N_c_158_n N_A_237_367#_c_198_n 0.00258991f $X=1.2 $Y=1.51 $X2=0
+ $Y2=0
cc_158 N_B1_N_c_159_n N_A_237_367#_c_198_n 0.0252213f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_159 N_B1_N_M1002_g N_VGND_c_404_n 0.00272283f $X=1.135 $Y=0.975 $X2=0 $Y2=0
cc_160 N_B1_N_M1002_g N_VGND_c_408_n 0.00432409f $X=1.135 $Y=0.975 $X2=0 $Y2=0
cc_161 N_A_237_367#_c_195_n N_A1_M1004_g 0.0259227f $X=2.105 $Y=1.51 $X2=0 $Y2=0
cc_162 N_A_237_367#_c_198_n N_A1_M1004_g 4.5018e-19 $X=1.81 $Y=1.51 $X2=0 $Y2=0
cc_163 N_A_237_367#_M1007_g A1 0.00691125f $X=2.105 $Y=0.655 $X2=0 $Y2=0
cc_164 N_A_237_367#_c_195_n A1 0.00898093f $X=2.105 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A_237_367#_c_197_n A1 0.00520396f $X=1.55 $Y=1.345 $X2=0 $Y2=0
cc_166 N_A_237_367#_c_198_n A1 0.00882436f $X=1.81 $Y=1.51 $X2=0 $Y2=0
cc_167 N_A_237_367#_M1007_g N_A1_c_260_n 0.0164024f $X=2.105 $Y=0.655 $X2=0
+ $Y2=0
cc_168 N_A_237_367#_c_198_n N_A1_c_260_n 2.80625e-19 $X=1.81 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A_237_367#_M1007_g N_A1_c_261_n 0.0229759f $X=2.105 $Y=0.655 $X2=0
+ $Y2=0
cc_170 N_A_237_367#_M1001_g N_VPWR_c_338_n 0.00585385f $X=2.105 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_237_367#_M1001_g N_VPWR_c_334_n 0.0120903f $X=2.105 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_237_367#_M1001_g N_A_436_367#_c_376_n 0.00115015f $X=2.105 $Y=2.465
+ $X2=0 $Y2=0
cc_173 N_A_237_367#_c_203_n N_A_436_367#_c_376_n 0.00131014f $X=1.55 $Y=1.93
+ $X2=0 $Y2=0
cc_174 N_A_237_367#_c_195_n N_A_436_367#_c_375_n 0.00263367f $X=2.105 $Y=1.51
+ $X2=0 $Y2=0
cc_175 N_A_237_367#_c_203_n N_A_436_367#_c_375_n 0.00456198f $X=1.55 $Y=1.93
+ $X2=0 $Y2=0
cc_176 N_A_237_367#_c_198_n N_A_436_367#_c_375_n 0.00247948f $X=1.81 $Y=1.51
+ $X2=0 $Y2=0
cc_177 N_A_237_367#_M1007_g N_VGND_c_402_n 0.00886947f $X=2.105 $Y=0.655 $X2=0
+ $Y2=0
cc_178 N_A_237_367#_M1007_g N_VGND_c_406_n 0.00353537f $X=2.105 $Y=0.655 $X2=0
+ $Y2=0
cc_179 N_A_237_367#_M1007_g N_VGND_c_408_n 0.00460168f $X=2.105 $Y=0.655 $X2=0
+ $Y2=0
cc_180 N_A1_M1004_g N_A2_M1000_g 0.0183877f $X=2.535 $Y=2.465 $X2=0 $Y2=0
cc_181 A1 A2 0.0188435f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A1_c_260_n A2 2.78241e-19 $X=2.615 $Y=1.35 $X2=0 $Y2=0
cc_183 A1 N_A2_c_295_n 0.00166163f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A1_c_260_n N_A2_c_295_n 0.0433148f $X=2.615 $Y=1.35 $X2=0 $Y2=0
cc_185 N_A1_c_261_n N_A2_c_296_n 0.0433148f $X=2.615 $Y=1.185 $X2=0 $Y2=0
cc_186 N_A1_M1004_g N_VPWR_c_336_n 0.00390609f $X=2.535 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A1_M1004_g N_VPWR_c_338_n 0.00585385f $X=2.535 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A1_M1004_g N_VPWR_c_334_n 0.0108362f $X=2.535 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A1_M1004_g N_A_436_367#_c_376_n 0.00162073f $X=2.535 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A1_M1004_g N_A_436_367#_c_374_n 0.0151914f $X=2.535 $Y=2.465 $X2=0
+ $Y2=0
cc_191 A1 N_A_436_367#_c_374_n 0.0256449f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A1_c_260_n N_A_436_367#_c_374_n 0.00481139f $X=2.615 $Y=1.35 $X2=0
+ $Y2=0
cc_193 A1 N_A_436_367#_c_375_n 0.0225326f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A1_c_261_n N_VGND_c_402_n 9.43385e-19 $X=2.615 $Y=1.185 $X2=0 $Y2=0
cc_195 N_A1_c_261_n N_VGND_c_403_n 0.00346344f $X=2.615 $Y=1.185 $X2=0 $Y2=0
cc_196 N_A1_c_261_n N_VGND_c_406_n 0.00585385f $X=2.615 $Y=1.185 $X2=0 $Y2=0
cc_197 N_A1_c_261_n N_VGND_c_408_n 0.0112227f $X=2.615 $Y=1.185 $X2=0 $Y2=0
cc_198 N_A2_M1000_g N_VPWR_c_336_n 0.00390609f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A2_M1000_g N_VPWR_c_339_n 0.00585385f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A2_M1000_g N_VPWR_c_334_n 0.01193f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_201 N_A2_M1000_g N_A_436_367#_c_374_n 0.0177726f $X=3.065 $Y=2.465 $X2=0
+ $Y2=0
cc_202 A2 N_A_436_367#_c_374_n 0.0310404f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A2_c_295_n N_A_436_367#_c_374_n 0.00519237f $X=3.185 $Y=1.35 $X2=0
+ $Y2=0
cc_204 N_A2_M1000_g N_A_436_367#_c_379_n 0.00434064f $X=3.065 $Y=2.465 $X2=0
+ $Y2=0
cc_205 A2 N_VGND_c_403_n 0.0243461f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_206 N_A2_c_295_n N_VGND_c_403_n 0.00485909f $X=3.185 $Y=1.35 $X2=0 $Y2=0
cc_207 N_A2_c_296_n N_VGND_c_403_n 0.0233404f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_208 N_A2_c_296_n N_VGND_c_406_n 0.00486043f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_209 N_A2_c_296_n N_VGND_c_408_n 0.00818711f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_210 X N_VPWR_c_337_n 0.0264135f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_211 N_X_M1009_s N_VPWR_c_334_n 0.00371702f $X=0.245 $Y=1.835 $X2=0 $Y2=0
cc_212 X N_VPWR_c_334_n 0.0146958f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_213 X N_VGND_c_401_n 0.00452266f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_214 X N_VGND_c_408_n 0.0104192f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_215 X N_VGND_c_409_n 0.0137839f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_216 N_VPWR_c_334_n N_A_436_367#_M1001_d 0.00293134f $X=3.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_217 N_VPWR_c_334_n N_A_436_367#_M1000_d 0.00336915f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_338_n N_A_436_367#_c_376_n 0.0149362f $X=2.635 $Y=3.33 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_334_n N_A_436_367#_c_376_n 0.0100304f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_220 N_VPWR_c_336_n N_A_436_367#_c_374_n 0.0243395f $X=2.8 $Y=2.055 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_339_n N_A_436_367#_c_379_n 0.0160153f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_334_n N_A_436_367#_c_379_n 0.00925289f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_223 N_VGND_c_408_n A_556_47# 0.00899413f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
