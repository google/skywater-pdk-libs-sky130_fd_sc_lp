* File: sky130_fd_sc_lp__o21bai_4.spice
* Created: Wed Sep  2 10:17:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21bai_4.pex.spice"
.subckt sky130_fd_sc_lp__o21bai_4  VNB VPB B1_N A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_B1_N_M1009_g N_A_27_49#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_A_218_49#_M1006_d N_A_27_49#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75005 A=0.126 P=1.98 MULT=1
MM1008 N_A_218_49#_M1008_d N_A_27_49#_M1008_g N_Y_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.5 A=0.126 P=1.98 MULT=1
MM1015 N_A_218_49#_M1008_d N_A_27_49#_M1015_g N_Y_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1018 N_A_218_49#_M1018_d N_A_27_49#_M1018_g N_Y_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1407 AS=0.1176 PD=1.175 PS=1.12 NRD=7.848 NRS=0 M=1 R=5.6
+ SA=75001.5 SB=75003.7 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A1_M1002_g N_A_218_49#_M1018_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1407 PD=1.12 PS=1.175 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75003.2
+ A=0.126 P=1.98 MULT=1
MM1000 N_A_218_49#_M1000_d N_A2_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1010 N_A_218_49#_M1000_d N_A2_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1012 N_A_218_49#_M1012_d N_A2_M1012_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1016 N_A_218_49#_M1012_d N_A2_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.7
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1016_s N_A1_M1005_g N_A_218_49#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1020 N_VGND_M1020_d N_A1_M1020_g N_A_218_49#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1020_d N_A1_M1022_g N_A_218_49#_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75005 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1024 N_VPWR_M1024_d N_B1_N_M1024_g N_A_27_49#_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.4725 AS=0.3339 PD=2.01 PS=3.05 NRD=73.481 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75005.9 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1024_d N_A_27_49#_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4725 AS=0.1764 PD=2.01 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1 SB=75005
+ A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A_27_49#_M1003_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1003_d N_A_27_49#_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75004.1
+ A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1021_d N_A_27_49#_M1021_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1004 N_A_653_367#_M1004_d N_A1_M1004_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75002.8 SB=75003.2 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1007_d N_A2_M1007_g N_A_653_367#_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.3
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1014 N_Y_M1007_d N_A2_M1014_g N_A_653_367#_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1017 N_Y_M1017_d N_A2_M1017_g N_A_653_367#_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1025 N_Y_M1017_d N_A2_M1025_g N_A_653_367#_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1013 N_A_653_367#_M1025_s N_A1_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1019 N_A_653_367#_M1019_d N_A1_M1019_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1023 N_A_653_367#_M1019_d N_A1_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75005.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=13.2415 P=17.93
*
.include "sky130_fd_sc_lp__o21bai_4.pxi.spice"
*
.ends
*
*
