* File: sky130_fd_sc_lp__a2bb2oi_m.spice
* Created: Wed Sep  2 09:24:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2oi_m.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2oi_m  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1005 N_A_202_47#_M1005_d N_A1_N_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A2_N_M1000_g N_A_202_47#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.06615 AS=0.0588 PD=0.735 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_202_47#_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.06615 PD=0.7 PS=0.735 NRD=0 NRS=9.996 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 A_467_47# N_B2_M1008_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0672
+ AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.7 A=0.063
+ P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g A_467_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75002 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1007 A_132_517# N_A1_N_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1449 PD=0.63 PS=1.53 NRD=23.443 NRS=37.5088 M=1 R=2.8
+ SA=75000.3 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_202_47#_M1002_d N_A2_N_M1002_g A_132_517# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_403_387#_M1006_d N_A_202_47#_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_B2_M1003_g N_A_403_387#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_403_387#_M1009_d N_B1_M1009_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_75 VPB 0 1.44327e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a2bb2oi_m.pxi.spice"
*
.ends
*
*
