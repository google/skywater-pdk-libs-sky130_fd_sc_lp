* File: sky130_fd_sc_lp__a311oi_4.pxi.spice
* Created: Fri Aug 28 09:58:36 2020
* 
x_PM_SKY130_FD_SC_LP__A311OI_4%A3 N_A3_c_151_n N_A3_M1012_g N_A3_M1008_g
+ N_A3_c_153_n N_A3_M1022_g N_A3_M1023_g N_A3_c_155_n N_A3_M1024_g N_A3_M1026_g
+ N_A3_c_157_n N_A3_M1039_g N_A3_M1034_g A3 A3 A3 A3 N_A3_c_160_n
+ PM_SKY130_FD_SC_LP__A311OI_4%A3
x_PM_SKY130_FD_SC_LP__A311OI_4%A2 N_A2_c_231_n N_A2_M1009_g N_A2_M1004_g
+ N_A2_c_233_n N_A2_M1018_g N_A2_M1014_g N_A2_c_235_n N_A2_M1032_g N_A2_M1020_g
+ N_A2_c_237_n N_A2_M1033_g N_A2_M1035_g A2 A2 A2 A2 N_A2_c_240_n
+ PM_SKY130_FD_SC_LP__A311OI_4%A2
x_PM_SKY130_FD_SC_LP__A311OI_4%A1 N_A1_M1002_g N_A1_c_318_n N_A1_c_319_n
+ N_A1_c_320_n N_A1_M1000_g N_A1_M1006_g N_A1_c_321_n N_A1_M1021_g N_A1_M1010_g
+ N_A1_c_322_n N_A1_M1028_g N_A1_M1017_g N_A1_c_323_n N_A1_M1037_g A1 A1 A1
+ N_A1_c_325_n PM_SKY130_FD_SC_LP__A311OI_4%A1
x_PM_SKY130_FD_SC_LP__A311OI_4%B1 N_B1_c_404_n N_B1_M1001_g N_B1_M1007_g
+ N_B1_c_406_n N_B1_M1013_g N_B1_M1025_g N_B1_c_408_n N_B1_M1015_g N_B1_M1029_g
+ N_B1_c_410_n N_B1_M1019_g N_B1_M1036_g B1 B1 B1 B1 N_B1_c_412_n N_B1_c_413_n
+ PM_SKY130_FD_SC_LP__A311OI_4%B1
x_PM_SKY130_FD_SC_LP__A311OI_4%C1 N_C1_c_493_n N_C1_M1005_g N_C1_M1003_g
+ N_C1_c_495_n N_C1_M1016_g N_C1_M1011_g N_C1_c_497_n N_C1_M1030_g N_C1_M1027_g
+ N_C1_c_499_n N_C1_M1031_g N_C1_M1038_g C1 C1 C1 C1 N_C1_c_502_n N_C1_c_503_n
+ PM_SKY130_FD_SC_LP__A311OI_4%C1
x_PM_SKY130_FD_SC_LP__A311OI_4%VPWR N_VPWR_M1008_d N_VPWR_M1023_d N_VPWR_M1034_d
+ N_VPWR_M1014_s N_VPWR_M1035_s N_VPWR_M1006_s N_VPWR_M1017_s N_VPWR_c_577_n
+ N_VPWR_c_578_n N_VPWR_c_579_n N_VPWR_c_580_n N_VPWR_c_581_n N_VPWR_c_582_n
+ N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n N_VPWR_c_587_n
+ N_VPWR_c_588_n N_VPWR_c_589_n N_VPWR_c_590_n N_VPWR_c_591_n N_VPWR_c_592_n
+ VPWR N_VPWR_c_593_n N_VPWR_c_594_n N_VPWR_c_595_n N_VPWR_c_576_n
+ N_VPWR_c_597_n N_VPWR_c_598_n PM_SKY130_FD_SC_LP__A311OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A311OI_4%A_124_367# N_A_124_367#_M1008_s
+ N_A_124_367#_M1026_s N_A_124_367#_M1004_d N_A_124_367#_M1020_d
+ N_A_124_367#_M1002_d N_A_124_367#_M1010_d N_A_124_367#_M1007_d
+ N_A_124_367#_M1029_d N_A_124_367#_c_727_n N_A_124_367#_c_721_n
+ N_A_124_367#_c_722_n N_A_124_367#_c_730_n N_A_124_367#_c_723_n
+ N_A_124_367#_c_732_n N_A_124_367#_c_724_n N_A_124_367#_c_734_n
+ N_A_124_367#_c_763_n N_A_124_367#_c_764_n N_A_124_367#_c_767_n
+ N_A_124_367#_c_775_n N_A_124_367#_c_811_n N_A_124_367#_c_735_n
+ N_A_124_367#_c_819_p N_A_124_367#_c_783_n N_A_124_367#_c_725_n
+ N_A_124_367#_c_726_n N_A_124_367#_c_770_n N_A_124_367#_c_779_n
+ N_A_124_367#_c_781_n N_A_124_367#_c_828_p N_A_124_367#_c_822_p
+ PM_SKY130_FD_SC_LP__A311OI_4%A_124_367#
x_PM_SKY130_FD_SC_LP__A311OI_4%A_1199_367# N_A_1199_367#_M1007_s
+ N_A_1199_367#_M1025_s N_A_1199_367#_M1036_s N_A_1199_367#_M1011_s
+ N_A_1199_367#_M1038_s N_A_1199_367#_c_834_n N_A_1199_367#_c_841_n
+ N_A_1199_367#_c_835_n N_A_1199_367#_c_844_n N_A_1199_367#_c_848_n
+ N_A_1199_367#_c_850_n N_A_1199_367#_c_857_n N_A_1199_367#_c_859_n
+ N_A_1199_367#_c_863_n N_A_1199_367#_c_836_n N_A_1199_367#_c_837_n
+ N_A_1199_367#_c_852_n N_A_1199_367#_c_854_n N_A_1199_367#_c_869_n
+ PM_SKY130_FD_SC_LP__A311OI_4%A_1199_367#
x_PM_SKY130_FD_SC_LP__A311OI_4%Y N_Y_M1000_d N_Y_M1021_d N_Y_M1037_d N_Y_M1013_s
+ N_Y_M1019_s N_Y_M1016_d N_Y_M1031_d N_Y_M1003_d N_Y_M1027_d N_Y_c_911_n
+ N_Y_c_912_n N_Y_c_937_n N_Y_c_941_n N_Y_c_1029_p N_Y_c_960_n N_Y_c_1030_p
+ N_Y_c_964_n N_Y_c_968_n N_Y_c_980_n N_Y_c_921_n N_Y_c_913_n N_Y_c_1032_p
+ N_Y_c_914_n N_Y_c_923_n N_Y_c_915_n N_Y_c_916_n N_Y_c_947_n N_Y_c_970_n
+ N_Y_c_972_n N_Y_c_974_n N_Y_c_917_n N_Y_c_999_n Y
+ PM_SKY130_FD_SC_LP__A311OI_4%Y
x_PM_SKY130_FD_SC_LP__A311OI_4%A_27_47# N_A_27_47#_M1012_s N_A_27_47#_M1022_s
+ N_A_27_47#_M1039_s N_A_27_47#_M1018_d N_A_27_47#_M1033_d N_A_27_47#_c_1055_n
+ N_A_27_47#_c_1057_n N_A_27_47#_c_1056_n N_A_27_47#_c_1092_p
+ N_A_27_47#_c_1063_n N_A_27_47#_c_1090_p N_A_27_47#_c_1070_n
+ N_A_27_47#_c_1074_n N_A_27_47#_c_1067_n N_A_27_47#_c_1069_n
+ N_A_27_47#_c_1079_n N_A_27_47#_c_1081_n PM_SKY130_FD_SC_LP__A311OI_4%A_27_47#
x_PM_SKY130_FD_SC_LP__A311OI_4%VGND N_VGND_M1012_d N_VGND_M1024_d N_VGND_M1001_d
+ N_VGND_M1015_d N_VGND_M1005_s N_VGND_M1030_s N_VGND_c_1111_n N_VGND_c_1112_n
+ N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n N_VGND_c_1116_n
+ N_VGND_c_1117_n N_VGND_c_1118_n N_VGND_c_1119_n N_VGND_c_1120_n
+ N_VGND_c_1121_n N_VGND_c_1122_n N_VGND_c_1123_n N_VGND_c_1124_n VGND
+ N_VGND_c_1125_n N_VGND_c_1126_n N_VGND_c_1127_n N_VGND_c_1128_n
+ N_VGND_c_1129_n N_VGND_c_1130_n PM_SKY130_FD_SC_LP__A311OI_4%VGND
x_PM_SKY130_FD_SC_LP__A311OI_4%A_454_47# N_A_454_47#_M1009_s N_A_454_47#_M1032_s
+ N_A_454_47#_M1000_s N_A_454_47#_M1028_s N_A_454_47#_c_1244_n
+ N_A_454_47#_c_1243_n N_A_454_47#_c_1248_n N_A_454_47#_c_1268_n
+ PM_SKY130_FD_SC_LP__A311OI_4%A_454_47#
cc_1 VNB N_A3_c_151_n 0.0218823f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_A3_M1008_g 0.0111699f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_3 VNB N_A3_c_153_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.185
cc_4 VNB N_A3_M1023_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_5 VNB N_A3_c_155_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.185
cc_6 VNB N_A3_M1026_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_7 VNB N_A3_c_157_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.185
cc_8 VNB N_A3_M1034_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_9 VNB A3 0.0132546f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_10 VNB N_A3_c_160_n 0.10964f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.35
cc_11 VNB N_A2_c_231_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_12 VNB N_A2_M1004_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_13 VNB N_A2_c_233_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.185
cc_14 VNB N_A2_M1014_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_15 VNB N_A2_c_235_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.185
cc_16 VNB N_A2_M1020_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_17 VNB N_A2_c_237_n 0.0198856f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.185
cc_18 VNB N_A2_M1035_g 0.00760942f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_19 VNB A2 0.00509024f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_20 VNB N_A2_c_240_n 0.0995122f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=1.35
cc_21 VNB N_A1_c_318_n 0.00770059f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_22 VNB N_A1_c_319_n 0.00890299f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_23 VNB N_A1_c_320_n 0.0194007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_321_n 0.0162036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_c_322_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A1_c_323_n 0.0165366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A1 0.00231539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_c_325_n 0.101875f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.35
cc_29 VNB N_B1_c_404_n 0.0163375f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_30 VNB N_B1_M1007_g 0.0100771f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_31 VNB N_B1_c_406_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.185
cc_32 VNB N_B1_M1025_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_33 VNB N_B1_c_408_n 0.0171175f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.185
cc_34 VNB N_B1_M1029_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_35 VNB N_B1_c_410_n 0.0173559f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.185
cc_36 VNB N_B1_M1036_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_37 VNB N_B1_c_412_n 0.00550454f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.35
cc_38 VNB N_B1_c_413_n 0.0958134f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.322
cc_39 VNB N_C1_c_493_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_40 VNB N_C1_M1003_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_41 VNB N_C1_c_495_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.185
cc_42 VNB N_C1_M1011_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_43 VNB N_C1_c_497_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.185
cc_44 VNB N_C1_M1027_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_45 VNB N_C1_c_499_n 0.0218823f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.185
cc_46 VNB N_C1_M1038_g 0.0111696f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_47 VNB C1 0.0144832f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_48 VNB N_C1_c_502_n 0.0755077f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.35
cc_49 VNB N_C1_c_503_n 0.0699596f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.35
cc_50 VNB N_VPWR_c_576_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_124_367#_c_721_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_52 VNB N_A_124_367#_c_722_n 0.00205518f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_53 VNB N_A_124_367#_c_723_n 0.00376651f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.35
cc_54 VNB N_A_124_367#_c_724_n 0.00486347f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.35
cc_55 VNB N_A_124_367#_c_725_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_124_367#_c_726_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Y_c_911_n 0.0170086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Y_c_912_n 5.04753e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_59 VNB N_Y_c_913_n 0.00554103f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.322
cc_60 VNB N_Y_c_914_n 0.00740486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_Y_c_915_n 0.0233935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_Y_c_916_n 0.00522433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_Y_c_917_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB Y 0.0106911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_27_47#_c_1055_n 0.0233935f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.515
cc_66 VNB N_A_27_47#_c_1056_n 0.00753748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1111_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1112_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=1.515
cc_69 VNB N_VGND_c_1113_n 4.06898e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_70 VNB N_VGND_c_1114_n 0.00430308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1115_n 3.18512e-19 $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.35
cc_72 VNB N_VGND_c_1116_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.35
cc_73 VNB N_VGND_c_1117_n 0.104372f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.35
cc_74 VNB N_VGND_c_1118_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.35
cc_75 VNB N_VGND_c_1119_n 0.0149824f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.35
cc_76 VNB N_VGND_c_1120_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.35
cc_77 VNB N_VGND_c_1121_n 0.0151002f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=1.35
cc_78 VNB N_VGND_c_1122_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.322
cc_79 VNB N_VGND_c_1123_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1124_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.322
cc_81 VNB N_VGND_c_1125_n 0.0153759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1126_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1127_n 0.0258771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1128_n 0.484337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1129_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1130_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_454_47#_c_1243_n 0.0111849f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.185
cc_88 VPB N_A3_M1008_g 0.0264709f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_89 VPB N_A3_M1023_g 0.0185652f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_90 VPB N_A3_M1026_g 0.0185652f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.465
cc_91 VPB N_A3_M1034_g 0.0186849f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_92 VPB N_A2_M1004_g 0.0186849f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_93 VPB N_A2_M1014_g 0.0185652f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_94 VPB N_A2_M1020_g 0.0185652f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.465
cc_95 VPB N_A2_M1035_g 0.0205851f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_96 VPB N_A1_M1002_g 0.0196795f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_97 VPB N_A1_c_318_n 0.0025893f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_98 VPB N_A1_c_319_n 3.31384e-19 $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_99 VPB N_A1_M1006_g 0.0181546f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_100 VPB N_A1_M1010_g 0.0181546f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.465
cc_101 VPB N_A1_M1017_g 0.0235997f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_102 VPB N_A1_c_325_n 0.00760551f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.35
cc_103 VPB N_B1_M1007_g 0.0251023f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_104 VPB N_B1_M1025_g 0.0188212f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_105 VPB N_B1_M1029_g 0.0188212f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.465
cc_106 VPB N_B1_M1036_g 0.0189644f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_107 VPB N_C1_M1003_g 0.0189499f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_108 VPB N_C1_M1011_g 0.0187643f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_109 VPB N_C1_M1027_g 0.0187643f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.465
cc_110 VPB N_C1_M1038_g 0.0272177f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_111 VPB N_VPWR_c_577_n 0.0125726f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.185
cc_112 VPB N_VPWR_c_578_n 0.0547871f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.655
cc_113 VPB N_VPWR_c_579_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_114 VPB N_VPWR_c_580_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_581_n 3.18512e-19 $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.35
cc_116 VPB N_VPWR_c_582_n 0.00427239f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.35
cc_117 VPB N_VPWR_c_583_n 3.18512e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_584_n 0.010471f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.322
cc_119 VPB N_VPWR_c_585_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_586_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_587_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_588_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_589_n 0.0151002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_590_n 0.00631492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_591_n 0.0149978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_592_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_593_n 0.012927f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_594_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_595_n 0.102893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_576_n 0.0669799f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_597_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_598_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_124_367#_c_727_n 0.00106657f $X=-0.19 $Y=1.655 $X2=1.835
+ $Y2=2.465
cc_134 VPB N_A_124_367#_c_721_n 0.00559032f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_135 VPB N_A_124_367#_c_722_n 0.00149292f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_136 VPB N_A_124_367#_c_730_n 9.96097e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_124_367#_c_723_n 0.00559032f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=1.35
cc_138 VPB N_A_124_367#_c_732_n 9.96097e-19 $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.35
cc_139 VPB N_A_124_367#_c_724_n 0.00559032f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.35
cc_140 VPB N_A_124_367#_c_734_n 4.98048e-19 $X=-0.19 $Y=1.655 $X2=1.835 $Y2=1.35
cc_141 VPB N_A_124_367#_c_735_n 0.011345f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_1199_367#_c_834_n 0.00589404f $X=-0.19 $Y=1.655 $X2=1.405
+ $Y2=1.515
cc_143 VPB N_A_1199_367#_c_835_n 0.001829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_1199_367#_c_836_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=1.35
cc_145 VPB N_A_1199_367#_c_837_n 0.044334f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.35
cc_146 VPB N_Y_c_911_n 0.0298611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_Y_c_912_n 0.00149303f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_148 VPB N_Y_c_921_n 0.00103081f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.322
cc_149 VPB N_Y_c_913_n 0.0072948f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.322
cc_150 VPB N_Y_c_923_n 0.00117631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 N_A3_c_157_n N_A2_c_231_n 0.0116592f $X=1.765 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A3_M1034_g N_A2_M1004_g 0.0268449f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_153 A3 A2 0.0198809f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A3_c_160_n A2 0.00114658f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_155 A3 N_A2_c_240_n 2.19457e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A3_c_160_n N_A2_c_240_n 0.0229793f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_157 N_A3_M1008_g N_VPWR_c_578_n 0.0225598f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A3_M1023_g N_VPWR_c_578_n 8.06385e-19 $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_159 A3 N_VPWR_c_578_n 0.014722f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A3_c_160_n N_VPWR_c_578_n 0.00709291f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A3_M1008_g N_VPWR_c_579_n 7.69607e-19 $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A3_M1023_g N_VPWR_c_579_n 0.01742f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A3_M1026_g N_VPWR_c_579_n 0.01742f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A3_M1034_g N_VPWR_c_579_n 7.69607e-19 $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A3_M1026_g N_VPWR_c_580_n 7.69607e-19 $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A3_M1034_g N_VPWR_c_580_n 0.0173454f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A3_M1026_g N_VPWR_c_585_n 0.00486043f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A3_M1034_g N_VPWR_c_585_n 0.00486043f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A3_M1008_g N_VPWR_c_593_n 0.00486043f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A3_M1023_g N_VPWR_c_593_n 0.00486043f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A3_M1008_g N_VPWR_c_576_n 0.00824727f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A3_M1023_g N_VPWR_c_576_n 0.00824727f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A3_M1026_g N_VPWR_c_576_n 0.00824727f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A3_M1034_g N_VPWR_c_576_n 0.00824727f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A3_M1008_g N_A_124_367#_c_727_n 0.00175293f $X=0.545 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A3_M1023_g N_A_124_367#_c_727_n 0.0014373f $X=0.975 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A3_M1023_g N_A_124_367#_c_721_n 0.0138902f $X=0.975 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A3_M1026_g N_A_124_367#_c_721_n 0.0142932f $X=1.405 $Y=2.465 $X2=0
+ $Y2=0
cc_179 A3 N_A_124_367#_c_721_n 0.0477264f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A3_c_160_n N_A_124_367#_c_721_n 0.00276559f $X=1.765 $Y=1.35 $X2=0
+ $Y2=0
cc_181 N_A3_M1008_g N_A_124_367#_c_722_n 0.00544609f $X=0.545 $Y=2.465 $X2=0
+ $Y2=0
cc_182 A3 N_A_124_367#_c_722_n 0.0156157f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A3_c_160_n N_A_124_367#_c_722_n 0.00286879f $X=1.765 $Y=1.35 $X2=0
+ $Y2=0
cc_184 N_A3_M1026_g N_A_124_367#_c_730_n 0.0014373f $X=1.405 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A3_M1034_g N_A_124_367#_c_730_n 0.0014373f $X=1.835 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A3_M1034_g N_A_124_367#_c_723_n 0.0147682f $X=1.835 $Y=2.465 $X2=0
+ $Y2=0
cc_187 A3 N_A_124_367#_c_723_n 0.00879067f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_188 A3 N_A_124_367#_c_725_n 0.0156157f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A3_c_160_n N_A_124_367#_c_725_n 0.00286879f $X=1.765 $Y=1.35 $X2=0
+ $Y2=0
cc_190 N_A3_c_151_n N_A_27_47#_c_1057_n 0.0122595f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_191 N_A3_c_153_n N_A_27_47#_c_1057_n 0.0122458f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_192 A3 N_A_27_47#_c_1057_n 0.039834f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_193 N_A3_c_160_n N_A_27_47#_c_1057_n 0.0025922f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_194 A3 N_A_27_47#_c_1056_n 0.0206589f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_195 N_A3_c_160_n N_A_27_47#_c_1056_n 0.00488323f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_196 N_A3_c_155_n N_A_27_47#_c_1063_n 0.0122595f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_197 N_A3_c_157_n N_A_27_47#_c_1063_n 0.0122458f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_198 A3 N_A_27_47#_c_1063_n 0.0382418f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_199 N_A3_c_160_n N_A_27_47#_c_1063_n 0.0025922f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_200 A3 N_A_27_47#_c_1067_n 0.0142048f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_201 N_A3_c_160_n N_A_27_47#_c_1067_n 0.00268449f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_202 N_A3_c_160_n N_A_27_47#_c_1069_n 5.98225e-19 $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_203 N_A3_c_151_n N_VGND_c_1111_n 0.0122575f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_204 N_A3_c_153_n N_VGND_c_1111_n 0.0105703f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_205 N_A3_c_155_n N_VGND_c_1111_n 5.75816e-19 $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_206 N_A3_c_153_n N_VGND_c_1112_n 5.75816e-19 $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_207 N_A3_c_155_n N_VGND_c_1112_n 0.0105703f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_208 N_A3_c_157_n N_VGND_c_1112_n 0.011763f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_209 N_A3_c_157_n N_VGND_c_1117_n 0.00486043f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_210 N_A3_c_151_n N_VGND_c_1125_n 0.00486043f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_211 N_A3_c_153_n N_VGND_c_1126_n 0.00486043f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_212 N_A3_c_155_n N_VGND_c_1126_n 0.00486043f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_213 N_A3_c_151_n N_VGND_c_1128_n 0.00917987f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_214 N_A3_c_153_n N_VGND_c_1128_n 0.00824727f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_215 N_A3_c_155_n N_VGND_c_1128_n 0.00824727f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_216 N_A3_c_157_n N_VGND_c_1128_n 0.0082726f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_217 N_A2_M1035_g N_A1_c_319_n 0.0277253f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A2_c_240_n N_A1_c_325_n 0.0056812f $X=3.645 $Y=1.35 $X2=0 $Y2=0
cc_219 N_A2_M1004_g N_VPWR_c_580_n 0.0173454f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A2_M1014_g N_VPWR_c_580_n 7.69607e-19 $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A2_M1004_g N_VPWR_c_581_n 7.69607e-19 $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A2_M1014_g N_VPWR_c_581_n 0.01742f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A2_M1020_g N_VPWR_c_581_n 0.0175335f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A2_M1035_g N_VPWR_c_581_n 8.59659e-19 $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A2_M1035_g N_VPWR_c_582_n 0.00272685f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A2_M1004_g N_VPWR_c_587_n 0.00486043f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_227 N_A2_M1014_g N_VPWR_c_587_n 0.00486043f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A2_M1020_g N_VPWR_c_589_n 0.00486043f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A2_M1035_g N_VPWR_c_589_n 0.00571722f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A2_M1004_g N_VPWR_c_576_n 0.00824727f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A2_M1014_g N_VPWR_c_576_n 0.00824727f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A2_M1020_g N_VPWR_c_576_n 0.00824727f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A2_M1035_g N_VPWR_c_576_n 0.0105481f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A2_M1004_g N_A_124_367#_c_723_n 0.0142932f $X=2.265 $Y=2.465 $X2=0
+ $Y2=0
cc_235 A2 N_A_124_367#_c_723_n 0.0272137f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_236 N_A2_c_240_n N_A_124_367#_c_723_n 0.00202617f $X=3.645 $Y=1.35 $X2=0
+ $Y2=0
cc_237 N_A2_M1004_g N_A_124_367#_c_732_n 0.0014373f $X=2.265 $Y=2.465 $X2=0
+ $Y2=0
cc_238 N_A2_M1014_g N_A_124_367#_c_732_n 0.0014373f $X=2.695 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A2_M1014_g N_A_124_367#_c_724_n 0.0143261f $X=2.695 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_A2_M1020_g N_A_124_367#_c_724_n 0.0143398f $X=3.125 $Y=2.465 $X2=0
+ $Y2=0
cc_241 N_A2_M1035_g N_A_124_367#_c_724_n 0.00534248f $X=3.555 $Y=2.465 $X2=0
+ $Y2=0
cc_242 A2 N_A_124_367#_c_724_n 0.0689561f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_243 N_A2_c_240_n N_A_124_367#_c_724_n 0.00563437f $X=3.645 $Y=1.35 $X2=0
+ $Y2=0
cc_244 N_A2_M1020_g N_A_124_367#_c_734_n 8.32811e-19 $X=3.125 $Y=2.465 $X2=0
+ $Y2=0
cc_245 N_A2_M1035_g N_A_124_367#_c_734_n 0.00380374f $X=3.555 $Y=2.465 $X2=0
+ $Y2=0
cc_246 N_A2_M1035_g N_A_124_367#_c_763_n 0.0120133f $X=3.555 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_A2_M1035_g N_A_124_367#_c_764_n 0.0130767f $X=3.555 $Y=2.465 $X2=0
+ $Y2=0
cc_248 A2 N_A_124_367#_c_764_n 0.00809206f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_249 N_A2_c_240_n N_A_124_367#_c_764_n 0.00321206f $X=3.645 $Y=1.35 $X2=0
+ $Y2=0
cc_250 N_A2_M1035_g N_A_124_367#_c_767_n 4.71645e-19 $X=3.555 $Y=2.465 $X2=0
+ $Y2=0
cc_251 A2 N_A_124_367#_c_726_n 0.0156157f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_252 N_A2_c_240_n N_A_124_367#_c_726_n 0.00286879f $X=3.645 $Y=1.35 $X2=0
+ $Y2=0
cc_253 N_A2_M1035_g N_A_124_367#_c_770_n 0.00113767f $X=3.555 $Y=2.465 $X2=0
+ $Y2=0
cc_254 N_A2_M1035_g N_Y_c_912_n 0.00145643f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_255 N_A2_c_237_n Y 0.00376583f $X=3.485 $Y=1.185 $X2=0 $Y2=0
cc_256 N_A2_M1035_g Y 0.00154884f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_257 A2 Y 0.0167812f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_258 N_A2_c_240_n Y 0.00357481f $X=3.645 $Y=1.35 $X2=0 $Y2=0
cc_259 N_A2_c_231_n N_A_27_47#_c_1070_n 0.0129469f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_260 N_A2_c_233_n N_A_27_47#_c_1070_n 0.00983632f $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_261 A2 N_A_27_47#_c_1070_n 0.0372338f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_262 N_A2_c_240_n N_A_27_47#_c_1070_n 0.0025922f $X=3.645 $Y=1.35 $X2=0 $Y2=0
cc_263 N_A2_c_235_n N_A_27_47#_c_1074_n 0.00979232f $X=3.055 $Y=1.185 $X2=0
+ $Y2=0
cc_264 N_A2_c_237_n N_A_27_47#_c_1074_n 0.00975958f $X=3.485 $Y=1.185 $X2=0
+ $Y2=0
cc_265 A2 N_A_27_47#_c_1074_n 0.0376019f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_266 N_A2_c_240_n N_A_27_47#_c_1074_n 0.0025922f $X=3.645 $Y=1.35 $X2=0 $Y2=0
cc_267 A2 N_A_27_47#_c_1069_n 0.00652125f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_268 A2 N_A_27_47#_c_1079_n 0.015815f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_269 N_A2_c_240_n N_A_27_47#_c_1079_n 0.00264019f $X=3.645 $Y=1.35 $X2=0 $Y2=0
cc_270 A2 N_A_27_47#_c_1081_n 0.0164266f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_271 N_A2_c_240_n N_A_27_47#_c_1081_n 0.00574416f $X=3.645 $Y=1.35 $X2=0 $Y2=0
cc_272 N_A2_c_231_n N_VGND_c_1112_n 0.00121814f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_273 N_A2_c_231_n N_VGND_c_1117_n 0.00585385f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_274 N_A2_c_233_n N_VGND_c_1117_n 0.00357877f $X=2.625 $Y=1.185 $X2=0 $Y2=0
cc_275 N_A2_c_235_n N_VGND_c_1117_n 0.00357877f $X=3.055 $Y=1.185 $X2=0 $Y2=0
cc_276 N_A2_c_237_n N_VGND_c_1117_n 0.00357877f $X=3.485 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A2_c_231_n N_VGND_c_1128_n 0.0108984f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_278 N_A2_c_233_n N_VGND_c_1128_n 0.00542194f $X=2.625 $Y=1.185 $X2=0 $Y2=0
cc_279 N_A2_c_235_n N_VGND_c_1128_n 0.00542194f $X=3.055 $Y=1.185 $X2=0 $Y2=0
cc_280 N_A2_c_237_n N_VGND_c_1128_n 0.0068216f $X=3.485 $Y=1.185 $X2=0 $Y2=0
cc_281 N_A2_c_233_n N_A_454_47#_c_1244_n 0.00978832f $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_282 N_A2_c_235_n N_A_454_47#_c_1244_n 0.00977268f $X=3.055 $Y=1.185 $X2=0
+ $Y2=0
cc_283 N_A2_c_237_n N_A_454_47#_c_1243_n 0.0134939f $X=3.485 $Y=1.185 $X2=0
+ $Y2=0
cc_284 N_A1_c_323_n N_B1_c_404_n 0.0140578f $X=5.725 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_285 A1 N_B1_c_412_n 0.01988f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_286 N_A1_c_325_n N_B1_c_412_n 0.00143623f $X=5.53 $Y=1.35 $X2=0 $Y2=0
cc_287 N_A1_c_325_n N_B1_c_413_n 0.0189016f $X=5.53 $Y=1.35 $X2=0 $Y2=0
cc_288 N_A1_M1002_g N_VPWR_c_582_n 0.00272685f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_289 N_A1_M1002_g N_VPWR_c_583_n 7.13785e-19 $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_290 N_A1_M1006_g N_VPWR_c_583_n 0.0144708f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A1_M1010_g N_VPWR_c_583_n 0.0143455f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A1_M1017_g N_VPWR_c_583_n 6.73419e-19 $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A1_M1010_g N_VPWR_c_584_n 6.73419e-19 $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A1_M1017_g N_VPWR_c_584_n 0.0168105f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_295 N_A1_M1002_g N_VPWR_c_591_n 0.00571722f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_296 N_A1_M1006_g N_VPWR_c_591_n 0.00486043f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A1_M1010_g N_VPWR_c_594_n 0.00486043f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A1_M1017_g N_VPWR_c_594_n 0.00486043f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A1_M1002_g N_VPWR_c_576_n 0.0105481f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A1_M1006_g N_VPWR_c_576_n 0.00824727f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A1_M1010_g N_VPWR_c_576_n 0.00824727f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A1_M1017_g N_VPWR_c_576_n 0.00824727f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A1_M1002_g N_A_124_367#_c_734_n 7.85616e-19 $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_304 N_A1_M1002_g N_A_124_367#_c_763_n 4.71645e-19 $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_A1_M1002_g N_A_124_367#_c_764_n 0.0127704f $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_306 N_A1_M1002_g N_A_124_367#_c_767_n 0.0115461f $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A1_M1006_g N_A_124_367#_c_775_n 0.0122595f $X=4.525 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A1_M1010_g N_A_124_367#_c_775_n 0.0122595f $X=4.955 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A1_c_325_n N_A_124_367#_c_775_n 5.26522e-19 $X=5.53 $Y=1.35 $X2=0 $Y2=0
cc_310 N_A1_M1017_g N_A_124_367#_c_735_n 0.0143f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_311 N_A1_M1002_g N_A_124_367#_c_779_n 2.7414e-19 $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_312 N_A1_c_318_n N_A_124_367#_c_779_n 6.04715e-19 $X=4.345 $Y=1.59 $X2=0
+ $Y2=0
cc_313 N_A1_c_325_n N_A_124_367#_c_781_n 5.96266e-19 $X=5.53 $Y=1.35 $X2=0 $Y2=0
cc_314 N_A1_M1017_g N_A_1199_367#_c_834_n 0.00136133f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_315 N_A1_c_318_n N_Y_c_911_n 0.00520284f $X=4.345 $Y=1.59 $X2=0 $Y2=0
cc_316 N_A1_M1006_g N_Y_c_911_n 0.00612865f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_317 N_A1_M1010_g N_Y_c_911_n 0.00615859f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A1_M1017_g N_Y_c_911_n 0.00747036f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_319 A1 N_Y_c_911_n 0.0943964f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_320 N_A1_c_325_n N_Y_c_911_n 0.0356479f $X=5.53 $Y=1.35 $X2=0 $Y2=0
cc_321 N_A1_M1002_g N_Y_c_912_n 0.00567237f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A1_c_319_n N_Y_c_912_n 0.00120909f $X=4.17 $Y=1.59 $X2=0 $Y2=0
cc_323 N_A1_c_320_n N_Y_c_937_n 0.01007f $X=4.435 $Y=1.185 $X2=0 $Y2=0
cc_324 N_A1_c_321_n N_Y_c_937_n 0.0096875f $X=4.865 $Y=1.185 $X2=0 $Y2=0
cc_325 A1 N_Y_c_937_n 0.0376019f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_326 N_A1_c_325_n N_Y_c_937_n 0.0026917f $X=5.53 $Y=1.35 $X2=0 $Y2=0
cc_327 N_A1_c_322_n N_Y_c_941_n 0.0096875f $X=5.295 $Y=1.185 $X2=0 $Y2=0
cc_328 N_A1_c_323_n N_Y_c_941_n 0.0137508f $X=5.725 $Y=1.185 $X2=0 $Y2=0
cc_329 A1 N_Y_c_941_n 0.0297976f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_330 N_A1_c_325_n N_Y_c_941_n 0.00230884f $X=5.53 $Y=1.35 $X2=0 $Y2=0
cc_331 N_A1_c_318_n N_Y_c_916_n 0.00311869f $X=4.345 $Y=1.59 $X2=0 $Y2=0
cc_332 N_A1_c_319_n N_Y_c_916_n 3.58832e-19 $X=4.17 $Y=1.59 $X2=0 $Y2=0
cc_333 A1 N_Y_c_947_n 0.0160195f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_334 N_A1_c_325_n N_Y_c_947_n 0.00274146f $X=5.53 $Y=1.35 $X2=0 $Y2=0
cc_335 N_A1_c_318_n Y 0.00398774f $X=4.345 $Y=1.59 $X2=0 $Y2=0
cc_336 N_A1_c_319_n Y 0.0051342f $X=4.17 $Y=1.59 $X2=0 $Y2=0
cc_337 N_A1_c_320_n Y 0.00490083f $X=4.435 $Y=1.185 $X2=0 $Y2=0
cc_338 A1 Y 0.0178948f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_339 N_A1_c_325_n Y 0.00362672f $X=5.53 $Y=1.35 $X2=0 $Y2=0
cc_340 N_A1_c_320_n N_A_27_47#_c_1081_n 2.58648e-19 $X=4.435 $Y=1.185 $X2=0
+ $Y2=0
cc_341 N_A1_c_323_n N_VGND_c_1113_n 0.00120001f $X=5.725 $Y=1.185 $X2=0 $Y2=0
cc_342 N_A1_c_320_n N_VGND_c_1117_n 0.00357877f $X=4.435 $Y=1.185 $X2=0 $Y2=0
cc_343 N_A1_c_321_n N_VGND_c_1117_n 0.00357877f $X=4.865 $Y=1.185 $X2=0 $Y2=0
cc_344 N_A1_c_322_n N_VGND_c_1117_n 0.00357877f $X=5.295 $Y=1.185 $X2=0 $Y2=0
cc_345 N_A1_c_323_n N_VGND_c_1117_n 0.00585385f $X=5.725 $Y=1.185 $X2=0 $Y2=0
cc_346 N_A1_c_320_n N_VGND_c_1128_n 0.0068216f $X=4.435 $Y=1.185 $X2=0 $Y2=0
cc_347 N_A1_c_321_n N_VGND_c_1128_n 0.00542194f $X=4.865 $Y=1.185 $X2=0 $Y2=0
cc_348 N_A1_c_322_n N_VGND_c_1128_n 0.00542194f $X=5.295 $Y=1.185 $X2=0 $Y2=0
cc_349 N_A1_c_323_n N_VGND_c_1128_n 0.0109224f $X=5.725 $Y=1.185 $X2=0 $Y2=0
cc_350 N_A1_c_320_n N_A_454_47#_c_1243_n 0.0135093f $X=4.435 $Y=1.185 $X2=0
+ $Y2=0
cc_351 N_A1_c_321_n N_A_454_47#_c_1248_n 0.0106614f $X=4.865 $Y=1.185 $X2=0
+ $Y2=0
cc_352 N_A1_c_322_n N_A_454_47#_c_1248_n 0.0106614f $X=5.295 $Y=1.185 $X2=0
+ $Y2=0
cc_353 N_B1_c_410_n N_C1_c_493_n 0.0149306f $X=7.555 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_354 N_B1_M1036_g N_C1_M1003_g 0.0278063f $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_355 N_B1_c_412_n C1 0.0159115f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_356 N_B1_c_413_n C1 2.76649e-19 $X=7.625 $Y=1.35 $X2=0 $Y2=0
cc_357 N_B1_c_412_n N_C1_c_502_n 2.76649e-19 $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_358 N_B1_c_413_n N_C1_c_502_n 0.0235325f $X=7.625 $Y=1.35 $X2=0 $Y2=0
cc_359 N_B1_M1007_g N_VPWR_c_584_n 0.00392606f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_360 N_B1_M1007_g N_VPWR_c_595_n 0.00357842f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_361 N_B1_M1025_g N_VPWR_c_595_n 0.00357842f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_362 N_B1_M1029_g N_VPWR_c_595_n 0.00357842f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_363 N_B1_M1036_g N_VPWR_c_595_n 0.00357842f $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_364 N_B1_M1007_g N_VPWR_c_576_n 0.00665087f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_365 N_B1_M1025_g N_VPWR_c_576_n 0.00535118f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_366 N_B1_M1029_g N_VPWR_c_576_n 0.00535118f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_367 N_B1_M1036_g N_VPWR_c_576_n 0.00537652f $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_368 N_B1_M1007_g N_A_124_367#_c_735_n 0.0143f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_369 N_B1_M1025_g N_A_124_367#_c_783_n 0.0122129f $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_370 N_B1_M1029_g N_A_124_367#_c_783_n 0.0122595f $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_371 N_B1_M1007_g N_A_1199_367#_c_834_n 0.0112773f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_372 N_B1_M1025_g N_A_1199_367#_c_834_n 5.62159e-19 $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_373 N_B1_M1007_g N_A_1199_367#_c_841_n 0.0105205f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_374 N_B1_M1025_g N_A_1199_367#_c_841_n 0.0105205f $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_375 N_B1_M1007_g N_A_1199_367#_c_835_n 5.89773e-19 $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_376 N_B1_M1007_g N_A_1199_367#_c_844_n 5.62159e-19 $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_377 N_B1_M1025_g N_A_1199_367#_c_844_n 0.00987577f $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_378 N_B1_M1029_g N_A_1199_367#_c_844_n 0.00987577f $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_379 N_B1_M1036_g N_A_1199_367#_c_844_n 5.62159e-19 $X=7.625 $Y=2.465 $X2=0
+ $Y2=0
cc_380 N_B1_M1029_g N_A_1199_367#_c_848_n 0.0105205f $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_381 N_B1_M1036_g N_A_1199_367#_c_848_n 0.0105205f $X=7.625 $Y=2.465 $X2=0
+ $Y2=0
cc_382 N_B1_M1029_g N_A_1199_367#_c_850_n 6.10534e-19 $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_383 N_B1_M1036_g N_A_1199_367#_c_850_n 0.0128917f $X=7.625 $Y=2.465 $X2=0
+ $Y2=0
cc_384 N_B1_M1025_g N_A_1199_367#_c_852_n 5.89773e-19 $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_385 N_B1_M1029_g N_A_1199_367#_c_852_n 5.89773e-19 $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_386 N_B1_M1036_g N_A_1199_367#_c_854_n 5.89773e-19 $X=7.625 $Y=2.465 $X2=0
+ $Y2=0
cc_387 N_B1_M1007_g N_Y_c_911_n 0.0125331f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_388 N_B1_M1025_g N_Y_c_911_n 0.0104926f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_389 N_B1_M1029_g N_Y_c_911_n 0.0104926f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_390 N_B1_M1036_g N_Y_c_911_n 0.0142932f $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_391 N_B1_c_412_n N_Y_c_911_n 0.132313f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_392 N_B1_c_413_n N_Y_c_911_n 0.0154471f $X=7.625 $Y=1.35 $X2=0 $Y2=0
cc_393 N_B1_c_404_n N_Y_c_960_n 0.0122595f $X=6.165 $Y=1.185 $X2=0 $Y2=0
cc_394 N_B1_c_406_n N_Y_c_960_n 0.0122595f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_395 N_B1_c_412_n N_Y_c_960_n 0.039834f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_396 N_B1_c_413_n N_Y_c_960_n 0.00271364f $X=7.625 $Y=1.35 $X2=0 $Y2=0
cc_397 N_B1_c_408_n N_Y_c_964_n 0.0135339f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_398 N_B1_c_410_n N_Y_c_964_n 0.0127965f $X=7.555 $Y=1.185 $X2=0 $Y2=0
cc_399 N_B1_c_412_n N_Y_c_964_n 0.0431266f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_400 N_B1_c_413_n N_Y_c_964_n 0.00530584f $X=7.625 $Y=1.35 $X2=0 $Y2=0
cc_401 N_B1_c_408_n N_Y_c_968_n 4.50559e-19 $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_402 N_B1_c_410_n N_Y_c_968_n 0.00801502f $X=7.555 $Y=1.185 $X2=0 $Y2=0
cc_403 N_B1_c_412_n N_Y_c_970_n 0.014505f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_404 N_B1_c_413_n N_Y_c_970_n 8.01838e-19 $X=7.625 $Y=1.35 $X2=0 $Y2=0
cc_405 N_B1_c_412_n N_Y_c_972_n 0.0158046f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_406 N_B1_c_413_n N_Y_c_972_n 0.00280606f $X=7.625 $Y=1.35 $X2=0 $Y2=0
cc_407 N_B1_c_410_n N_Y_c_974_n 2.74535e-19 $X=7.555 $Y=1.185 $X2=0 $Y2=0
cc_408 N_B1_c_412_n N_Y_c_974_n 0.00380661f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_409 N_B1_c_413_n N_Y_c_974_n 0.00178162f $X=7.625 $Y=1.35 $X2=0 $Y2=0
cc_410 N_B1_c_404_n N_VGND_c_1113_n 0.0117721f $X=6.165 $Y=1.185 $X2=0 $Y2=0
cc_411 N_B1_c_406_n N_VGND_c_1113_n 0.0106734f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_412 N_B1_c_408_n N_VGND_c_1113_n 5.94039e-19 $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_413 N_B1_c_408_n N_VGND_c_1114_n 0.00258937f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_414 N_B1_c_410_n N_VGND_c_1114_n 0.00253973f $X=7.555 $Y=1.185 $X2=0 $Y2=0
cc_415 N_B1_c_410_n N_VGND_c_1115_n 6.27534e-19 $X=7.555 $Y=1.185 $X2=0 $Y2=0
cc_416 N_B1_c_404_n N_VGND_c_1117_n 0.00486043f $X=6.165 $Y=1.185 $X2=0 $Y2=0
cc_417 N_B1_c_406_n N_VGND_c_1119_n 0.00486043f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_418 N_B1_c_408_n N_VGND_c_1119_n 0.00585385f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_419 N_B1_c_410_n N_VGND_c_1121_n 0.00571722f $X=7.555 $Y=1.185 $X2=0 $Y2=0
cc_420 N_B1_c_404_n N_VGND_c_1128_n 0.00829667f $X=6.165 $Y=1.185 $X2=0 $Y2=0
cc_421 N_B1_c_406_n N_VGND_c_1128_n 0.00824727f $X=6.595 $Y=1.185 $X2=0 $Y2=0
cc_422 N_B1_c_408_n N_VGND_c_1128_n 0.0109131f $X=7.025 $Y=1.185 $X2=0 $Y2=0
cc_423 N_B1_c_410_n N_VGND_c_1128_n 0.0106693f $X=7.555 $Y=1.185 $X2=0 $Y2=0
cc_424 N_C1_M1003_g N_VPWR_c_595_n 0.00357842f $X=8.055 $Y=2.465 $X2=0 $Y2=0
cc_425 N_C1_M1011_g N_VPWR_c_595_n 0.00357842f $X=8.485 $Y=2.465 $X2=0 $Y2=0
cc_426 N_C1_M1027_g N_VPWR_c_595_n 0.00357842f $X=8.915 $Y=2.465 $X2=0 $Y2=0
cc_427 N_C1_M1038_g N_VPWR_c_595_n 0.00357877f $X=9.345 $Y=2.465 $X2=0 $Y2=0
cc_428 N_C1_M1003_g N_VPWR_c_576_n 0.00537652f $X=8.055 $Y=2.465 $X2=0 $Y2=0
cc_429 N_C1_M1011_g N_VPWR_c_576_n 0.00535118f $X=8.485 $Y=2.465 $X2=0 $Y2=0
cc_430 N_C1_M1027_g N_VPWR_c_576_n 0.00535118f $X=8.915 $Y=2.465 $X2=0 $Y2=0
cc_431 N_C1_M1038_g N_VPWR_c_576_n 0.00645423f $X=9.345 $Y=2.465 $X2=0 $Y2=0
cc_432 N_C1_M1003_g N_A_1199_367#_c_850_n 0.0129114f $X=8.055 $Y=2.465 $X2=0
+ $Y2=0
cc_433 N_C1_M1011_g N_A_1199_367#_c_850_n 6.58347e-19 $X=8.485 $Y=2.465 $X2=0
+ $Y2=0
cc_434 N_C1_M1003_g N_A_1199_367#_c_857_n 0.0105205f $X=8.055 $Y=2.465 $X2=0
+ $Y2=0
cc_435 N_C1_M1011_g N_A_1199_367#_c_857_n 0.0105205f $X=8.485 $Y=2.465 $X2=0
+ $Y2=0
cc_436 N_C1_M1003_g N_A_1199_367#_c_859_n 6.58347e-19 $X=8.055 $Y=2.465 $X2=0
+ $Y2=0
cc_437 N_C1_M1011_g N_A_1199_367#_c_859_n 0.0129502f $X=8.485 $Y=2.465 $X2=0
+ $Y2=0
cc_438 N_C1_M1027_g N_A_1199_367#_c_859_n 0.0130588f $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_439 N_C1_M1038_g N_A_1199_367#_c_859_n 6.66596e-19 $X=9.345 $Y=2.465 $X2=0
+ $Y2=0
cc_440 N_C1_M1027_g N_A_1199_367#_c_863_n 0.0105205f $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_441 N_C1_M1038_g N_A_1199_367#_c_863_n 0.012237f $X=9.345 $Y=2.465 $X2=0
+ $Y2=0
cc_442 N_C1_M1038_g N_A_1199_367#_c_837_n 0.00346841f $X=9.345 $Y=2.465 $X2=0
+ $Y2=0
cc_443 C1 N_A_1199_367#_c_837_n 0.0130246f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_444 N_C1_c_503_n N_A_1199_367#_c_837_n 0.00649196f $X=9.775 $Y=1.35 $X2=0
+ $Y2=0
cc_445 N_C1_M1003_g N_A_1199_367#_c_854_n 5.89773e-19 $X=8.055 $Y=2.465 $X2=0
+ $Y2=0
cc_446 N_C1_M1011_g N_A_1199_367#_c_869_n 5.89773e-19 $X=8.485 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_C1_M1027_g N_A_1199_367#_c_869_n 5.89773e-19 $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_448 N_C1_M1003_g N_Y_c_911_n 0.0142932f $X=8.055 $Y=2.465 $X2=0 $Y2=0
cc_449 C1 N_Y_c_911_n 0.0187504f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_450 N_C1_c_502_n N_Y_c_911_n 0.00202617f $X=9.42 $Y=1.35 $X2=0 $Y2=0
cc_451 N_C1_c_493_n N_Y_c_980_n 0.0122595f $X=7.985 $Y=1.185 $X2=0 $Y2=0
cc_452 N_C1_c_495_n N_Y_c_980_n 0.0122458f $X=8.415 $Y=1.185 $X2=0 $Y2=0
cc_453 C1 N_Y_c_980_n 0.0382418f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_454 N_C1_c_502_n N_Y_c_980_n 0.0025922f $X=9.42 $Y=1.35 $X2=0 $Y2=0
cc_455 N_C1_M1003_g N_Y_c_921_n 0.00229987f $X=8.055 $Y=2.465 $X2=0 $Y2=0
cc_456 N_C1_M1011_g N_Y_c_921_n 0.00165214f $X=8.485 $Y=2.465 $X2=0 $Y2=0
cc_457 N_C1_M1011_g N_Y_c_913_n 0.0142932f $X=8.485 $Y=2.465 $X2=0 $Y2=0
cc_458 N_C1_M1027_g N_Y_c_913_n 0.0140113f $X=8.915 $Y=2.465 $X2=0 $Y2=0
cc_459 N_C1_M1038_g N_Y_c_913_n 0.00572358f $X=9.345 $Y=2.465 $X2=0 $Y2=0
cc_460 C1 N_Y_c_913_n 0.0666303f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_461 N_C1_c_502_n N_Y_c_913_n 0.00563437f $X=9.42 $Y=1.35 $X2=0 $Y2=0
cc_462 N_C1_c_497_n N_Y_c_914_n 0.0122595f $X=8.845 $Y=1.185 $X2=0 $Y2=0
cc_463 N_C1_c_499_n N_Y_c_914_n 0.0122595f $X=9.275 $Y=1.185 $X2=0 $Y2=0
cc_464 C1 N_Y_c_914_n 0.0602418f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_465 N_C1_c_502_n N_Y_c_914_n 0.00887638f $X=9.42 $Y=1.35 $X2=0 $Y2=0
cc_466 N_C1_M1027_g N_Y_c_923_n 0.00167621f $X=8.915 $Y=2.465 $X2=0 $Y2=0
cc_467 N_C1_M1038_g N_Y_c_923_n 0.00214694f $X=9.345 $Y=2.465 $X2=0 $Y2=0
cc_468 C1 N_Y_c_917_n 0.0156157f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_469 N_C1_c_502_n N_Y_c_917_n 0.00286879f $X=9.42 $Y=1.35 $X2=0 $Y2=0
cc_470 C1 N_Y_c_999_n 0.0142048f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_471 N_C1_c_502_n N_Y_c_999_n 0.00268449f $X=9.42 $Y=1.35 $X2=0 $Y2=0
cc_472 N_C1_c_493_n N_VGND_c_1115_n 0.0106956f $X=7.985 $Y=1.185 $X2=0 $Y2=0
cc_473 N_C1_c_495_n N_VGND_c_1115_n 0.0105703f $X=8.415 $Y=1.185 $X2=0 $Y2=0
cc_474 N_C1_c_497_n N_VGND_c_1115_n 5.75816e-19 $X=8.845 $Y=1.185 $X2=0 $Y2=0
cc_475 N_C1_c_495_n N_VGND_c_1116_n 5.75816e-19 $X=8.415 $Y=1.185 $X2=0 $Y2=0
cc_476 N_C1_c_497_n N_VGND_c_1116_n 0.0105703f $X=8.845 $Y=1.185 $X2=0 $Y2=0
cc_477 N_C1_c_499_n N_VGND_c_1116_n 0.0122575f $X=9.275 $Y=1.185 $X2=0 $Y2=0
cc_478 N_C1_c_493_n N_VGND_c_1121_n 0.00486043f $X=7.985 $Y=1.185 $X2=0 $Y2=0
cc_479 N_C1_c_495_n N_VGND_c_1123_n 0.00486043f $X=8.415 $Y=1.185 $X2=0 $Y2=0
cc_480 N_C1_c_497_n N_VGND_c_1123_n 0.00486043f $X=8.845 $Y=1.185 $X2=0 $Y2=0
cc_481 N_C1_c_499_n N_VGND_c_1127_n 0.00486043f $X=9.275 $Y=1.185 $X2=0 $Y2=0
cc_482 N_C1_c_493_n N_VGND_c_1128_n 0.0082726f $X=7.985 $Y=1.185 $X2=0 $Y2=0
cc_483 N_C1_c_495_n N_VGND_c_1128_n 0.00824727f $X=8.415 $Y=1.185 $X2=0 $Y2=0
cc_484 N_C1_c_497_n N_VGND_c_1128_n 0.00824727f $X=8.845 $Y=1.185 $X2=0 $Y2=0
cc_485 N_C1_c_499_n N_VGND_c_1128_n 0.00954696f $X=9.275 $Y=1.185 $X2=0 $Y2=0
cc_486 N_VPWR_c_576_n N_A_124_367#_M1008_s 0.00536646f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_487 N_VPWR_c_576_n N_A_124_367#_M1026_s 0.00536646f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_576_n N_A_124_367#_M1004_d 0.00536646f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_576_n N_A_124_367#_M1020_d 0.00380103f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_576_n N_A_124_367#_M1002_d 0.00380103f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_576_n N_A_124_367#_M1010_d 0.00536646f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_576_n N_A_124_367#_M1007_d 0.00225186f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_576_n N_A_124_367#_M1029_d 0.00225186f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_578_n N_A_124_367#_c_727_n 0.0480052f $X=0.33 $Y=1.98 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_593_n N_A_124_367#_c_727_n 0.0124525f $X=1.025 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_576_n N_A_124_367#_c_727_n 0.00730901f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_579_n N_A_124_367#_c_721_n 0.0216087f $X=1.19 $Y=2.03 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_585_n N_A_124_367#_c_730_n 0.0124525f $X=1.885 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_576_n N_A_124_367#_c_730_n 0.00730901f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_580_n N_A_124_367#_c_723_n 0.0216087f $X=2.05 $Y=2.03 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_587_n N_A_124_367#_c_732_n 0.0124525f $X=2.745 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_576_n N_A_124_367#_c_732_n 0.00730901f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_581_n N_A_124_367#_c_724_n 0.0216087f $X=2.91 $Y=2.03 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_589_n N_A_124_367#_c_763_n 0.0146655f $X=3.66 $Y=3.33 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_576_n N_A_124_367#_c_763_n 0.00933292f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_506 N_VPWR_M1035_s N_A_124_367#_c_764_n 0.0108868f $X=3.63 $Y=1.835 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_582_n N_A_124_367#_c_764_n 0.022455f $X=3.825 $Y=2.39 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_591_n N_A_124_367#_c_767_n 0.0146655f $X=4.575 $Y=3.33 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_576_n N_A_124_367#_c_767_n 0.00933292f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_510 N_VPWR_M1006_s N_A_124_367#_c_775_n 0.00334047f $X=4.6 $Y=1.835 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_583_n N_A_124_367#_c_775_n 0.0170777f $X=4.74 $Y=2.39 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_594_n N_A_124_367#_c_811_n 0.0124525f $X=5.435 $Y=3.33 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_576_n N_A_124_367#_c_811_n 0.00730901f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_514 N_VPWR_M1017_s N_A_124_367#_c_735_n 0.0049409f $X=5.46 $Y=1.835 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_584_n N_A_124_367#_c_735_n 0.0220026f $X=5.6 $Y=2.39 $X2=0 $Y2=0
cc_516 N_VPWR_c_576_n N_A_1199_367#_M1007_s 0.00215158f $X=9.84 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_517 N_VPWR_c_576_n N_A_1199_367#_M1025_s 0.00223559f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_576_n N_A_1199_367#_M1036_s 0.00223559f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_576_n N_A_1199_367#_M1011_s 0.00223559f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_576_n N_A_1199_367#_M1038_s 0.00215159f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_584_n N_A_1199_367#_c_834_n 0.047703f $X=5.6 $Y=2.39 $X2=0 $Y2=0
cc_522 N_VPWR_c_595_n N_A_1199_367#_c_841_n 0.0298674f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_576_n N_A_1199_367#_c_841_n 0.0187823f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_584_n N_A_1199_367#_c_835_n 0.0139f $X=5.6 $Y=2.39 $X2=0 $Y2=0
cc_525 N_VPWR_c_595_n N_A_1199_367#_c_835_n 0.0211865f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_576_n N_A_1199_367#_c_835_n 0.0126421f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_595_n N_A_1199_367#_c_848_n 0.0298674f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_576_n N_A_1199_367#_c_848_n 0.0187823f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_595_n N_A_1199_367#_c_857_n 0.0298674f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_576_n N_A_1199_367#_c_857_n 0.0187823f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_595_n N_A_1199_367#_c_863_n 0.0319341f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_576_n N_A_1199_367#_c_863_n 0.0201012f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_595_n N_A_1199_367#_c_836_n 0.0189827f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_576_n N_A_1199_367#_c_836_n 0.0112692f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_595_n N_A_1199_367#_c_852_n 0.01906f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_536 N_VPWR_c_576_n N_A_1199_367#_c_852_n 0.0124545f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_595_n N_A_1199_367#_c_854_n 0.01906f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_538 N_VPWR_c_576_n N_A_1199_367#_c_854_n 0.0124545f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_595_n N_A_1199_367#_c_869_n 0.01906f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_540 N_VPWR_c_576_n N_A_1199_367#_c_869_n 0.0124545f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_576_n N_Y_M1003_d 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_542 N_VPWR_c_576_n N_Y_M1027_d 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_543 N_A_124_367#_c_735_n N_A_1199_367#_M1007_s 0.00494644f $X=6.455 $Y=2.03
+ $X2=-0.19 $Y2=-0.245
cc_544 N_A_124_367#_c_783_n N_A_1199_367#_M1025_s 0.00339285f $X=7.315 $Y=2.03
+ $X2=0 $Y2=0
cc_545 N_A_124_367#_c_735_n N_A_1199_367#_c_834_n 0.0220026f $X=6.455 $Y=2.03
+ $X2=0 $Y2=0
cc_546 N_A_124_367#_M1007_d N_A_1199_367#_c_841_n 0.00332344f $X=6.41 $Y=1.835
+ $X2=0 $Y2=0
cc_547 N_A_124_367#_c_819_p N_A_1199_367#_c_841_n 0.0126348f $X=6.55 $Y=2.57
+ $X2=0 $Y2=0
cc_548 N_A_124_367#_c_783_n N_A_1199_367#_c_844_n 0.0170777f $X=7.315 $Y=2.03
+ $X2=0 $Y2=0
cc_549 N_A_124_367#_M1029_d N_A_1199_367#_c_848_n 0.00332344f $X=7.27 $Y=1.835
+ $X2=0 $Y2=0
cc_550 N_A_124_367#_c_822_p N_A_1199_367#_c_848_n 0.0126348f $X=7.41 $Y=2.11
+ $X2=0 $Y2=0
cc_551 N_A_124_367#_c_775_n N_Y_c_911_n 0.0402255f $X=5.075 $Y=2.03 $X2=0 $Y2=0
cc_552 N_A_124_367#_c_735_n N_Y_c_911_n 0.0790486f $X=6.455 $Y=2.03 $X2=0 $Y2=0
cc_553 N_A_124_367#_c_783_n N_Y_c_911_n 0.0402256f $X=7.315 $Y=2.03 $X2=0 $Y2=0
cc_554 N_A_124_367#_c_779_n N_Y_c_911_n 0.0161083f $X=4.31 $Y=2.03 $X2=0 $Y2=0
cc_555 N_A_124_367#_c_781_n N_Y_c_911_n 0.0146338f $X=5.17 $Y=2.03 $X2=0 $Y2=0
cc_556 N_A_124_367#_c_828_p N_Y_c_911_n 0.0146339f $X=6.55 $Y=2.03 $X2=0 $Y2=0
cc_557 N_A_124_367#_c_822_p N_Y_c_911_n 0.0146339f $X=7.41 $Y=2.11 $X2=0 $Y2=0
cc_558 N_A_124_367#_c_724_n N_Y_c_912_n 0.00682007f $X=3.245 $Y=1.69 $X2=0 $Y2=0
cc_559 N_A_124_367#_c_764_n N_Y_c_912_n 0.0117968f $X=4.16 $Y=2.03 $X2=0 $Y2=0
cc_560 N_A_124_367#_c_779_n N_Y_c_912_n 0.00103843f $X=4.31 $Y=2.03 $X2=0 $Y2=0
cc_561 N_A_124_367#_c_723_n N_A_27_47#_c_1069_n 0.00402068f $X=2.385 $Y=1.69
+ $X2=0 $Y2=0
cc_562 N_A_1199_367#_c_857_n N_Y_M1003_d 0.00332344f $X=8.535 $Y=2.99 $X2=0
+ $Y2=0
cc_563 N_A_1199_367#_c_863_n N_Y_M1027_d 0.00332344f $X=9.435 $Y=2.99 $X2=0
+ $Y2=0
cc_564 N_A_1199_367#_c_850_n N_Y_c_911_n 0.0216087f $X=7.84 $Y=2.03 $X2=0 $Y2=0
cc_565 N_A_1199_367#_c_857_n N_Y_c_921_n 0.0126348f $X=8.535 $Y=2.99 $X2=0 $Y2=0
cc_566 N_A_1199_367#_c_859_n N_Y_c_913_n 0.0216087f $X=8.7 $Y=2.03 $X2=0 $Y2=0
cc_567 N_A_1199_367#_c_863_n N_Y_c_923_n 0.0126348f $X=9.435 $Y=2.99 $X2=0 $Y2=0
cc_568 N_A_1199_367#_c_837_n N_Y_c_923_n 0.00152359f $X=9.56 $Y=1.98 $X2=0 $Y2=0
cc_569 N_Y_c_916_n N_A_27_47#_c_1081_n 0.0310717f $X=4.355 $Y=0.847 $X2=0 $Y2=0
cc_570 N_Y_c_960_n N_VGND_M1001_d 0.00329816f $X=6.715 $Y=0.955 $X2=0 $Y2=0
cc_571 N_Y_c_964_n N_VGND_M1015_d 0.00536854f $X=7.62 $Y=0.955 $X2=0 $Y2=0
cc_572 N_Y_c_980_n N_VGND_M1005_s 0.00329816f $X=8.535 $Y=0.955 $X2=0 $Y2=0
cc_573 N_Y_c_914_n N_VGND_M1030_s 0.00329816f $X=9.395 $Y=0.955 $X2=0 $Y2=0
cc_574 N_Y_c_960_n N_VGND_c_1113_n 0.0170777f $X=6.715 $Y=0.955 $X2=0 $Y2=0
cc_575 N_Y_c_964_n N_VGND_c_1114_n 0.0216414f $X=7.62 $Y=0.955 $X2=0 $Y2=0
cc_576 N_Y_c_980_n N_VGND_c_1115_n 0.0170777f $X=8.535 $Y=0.955 $X2=0 $Y2=0
cc_577 N_Y_c_914_n N_VGND_c_1116_n 0.0170777f $X=9.395 $Y=0.955 $X2=0 $Y2=0
cc_578 N_Y_c_1029_p N_VGND_c_1117_n 0.0145748f $X=5.94 $Y=0.42 $X2=0 $Y2=0
cc_579 N_Y_c_1030_p N_VGND_c_1119_n 0.0140491f $X=6.81 $Y=0.42 $X2=0 $Y2=0
cc_580 N_Y_c_968_n N_VGND_c_1121_n 0.0146655f $X=7.77 $Y=0.42 $X2=0 $Y2=0
cc_581 N_Y_c_1032_p N_VGND_c_1123_n 0.0124525f $X=8.63 $Y=0.42 $X2=0 $Y2=0
cc_582 N_Y_c_915_n N_VGND_c_1127_n 0.0178111f $X=9.49 $Y=0.42 $X2=0 $Y2=0
cc_583 N_Y_M1000_d N_VGND_c_1128_n 0.0021598f $X=4.095 $Y=0.235 $X2=0 $Y2=0
cc_584 N_Y_M1021_d N_VGND_c_1128_n 0.00225186f $X=4.94 $Y=0.235 $X2=0 $Y2=0
cc_585 N_Y_M1037_d N_VGND_c_1128_n 0.00405538f $X=5.8 $Y=0.235 $X2=0 $Y2=0
cc_586 N_Y_M1013_s N_VGND_c_1128_n 0.00380103f $X=6.67 $Y=0.235 $X2=0 $Y2=0
cc_587 N_Y_M1019_s N_VGND_c_1128_n 0.00380103f $X=7.63 $Y=0.235 $X2=0 $Y2=0
cc_588 N_Y_M1016_d N_VGND_c_1128_n 0.00536646f $X=8.49 $Y=0.235 $X2=0 $Y2=0
cc_589 N_Y_M1031_d N_VGND_c_1128_n 0.00371702f $X=9.35 $Y=0.235 $X2=0 $Y2=0
cc_590 N_Y_c_1029_p N_VGND_c_1128_n 0.00925289f $X=5.94 $Y=0.42 $X2=0 $Y2=0
cc_591 N_Y_c_1030_p N_VGND_c_1128_n 0.0090585f $X=6.81 $Y=0.42 $X2=0 $Y2=0
cc_592 N_Y_c_968_n N_VGND_c_1128_n 0.00933292f $X=7.77 $Y=0.42 $X2=0 $Y2=0
cc_593 N_Y_c_1032_p N_VGND_c_1128_n 0.00730901f $X=8.63 $Y=0.42 $X2=0 $Y2=0
cc_594 N_Y_c_915_n N_VGND_c_1128_n 0.0100304f $X=9.49 $Y=0.42 $X2=0 $Y2=0
cc_595 N_Y_c_937_n N_A_454_47#_M1000_s 0.00329816f $X=4.95 $Y=0.955 $X2=0 $Y2=0
cc_596 N_Y_c_941_n N_A_454_47#_M1028_s 0.00329816f $X=5.805 $Y=0.955 $X2=0 $Y2=0
cc_597 N_Y_M1000_d N_A_454_47#_c_1243_n 0.00528143f $X=4.095 $Y=0.235 $X2=0
+ $Y2=0
cc_598 N_Y_c_937_n N_A_454_47#_c_1243_n 0.018408f $X=4.95 $Y=0.955 $X2=0 $Y2=0
cc_599 N_Y_c_916_n N_A_454_47#_c_1243_n 0.0234019f $X=4.355 $Y=0.847 $X2=0 $Y2=0
cc_600 N_Y_M1021_d N_A_454_47#_c_1248_n 0.00335455f $X=4.94 $Y=0.235 $X2=0 $Y2=0
cc_601 N_Y_c_937_n N_A_454_47#_c_1248_n 0.00535657f $X=4.95 $Y=0.955 $X2=0 $Y2=0
cc_602 N_Y_c_941_n N_A_454_47#_c_1248_n 0.018408f $X=5.805 $Y=0.955 $X2=0 $Y2=0
cc_603 N_Y_c_947_n N_A_454_47#_c_1248_n 0.0125258f $X=5.08 $Y=0.82 $X2=0 $Y2=0
cc_604 N_A_27_47#_c_1057_n N_VGND_M1012_d 0.00329816f $X=1.025 $Y=0.955
+ $X2=-0.19 $Y2=-0.245
cc_605 N_A_27_47#_c_1063_n N_VGND_M1024_d 0.00329816f $X=1.885 $Y=0.955 $X2=0
+ $Y2=0
cc_606 N_A_27_47#_c_1057_n N_VGND_c_1111_n 0.0170777f $X=1.025 $Y=0.955 $X2=0
+ $Y2=0
cc_607 N_A_27_47#_c_1063_n N_VGND_c_1112_n 0.0170777f $X=1.885 $Y=0.955 $X2=0
+ $Y2=0
cc_608 N_A_27_47#_c_1090_p N_VGND_c_1117_n 0.0138717f $X=1.98 $Y=0.42 $X2=0
+ $Y2=0
cc_609 N_A_27_47#_c_1055_n N_VGND_c_1125_n 0.0178111f $X=0.26 $Y=0.42 $X2=0
+ $Y2=0
cc_610 N_A_27_47#_c_1092_p N_VGND_c_1126_n 0.0124525f $X=1.12 $Y=0.42 $X2=0
+ $Y2=0
cc_611 N_A_27_47#_M1012_s N_VGND_c_1128_n 0.00371702f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_612 N_A_27_47#_M1022_s N_VGND_c_1128_n 0.00536646f $X=0.98 $Y=0.235 $X2=0
+ $Y2=0
cc_613 N_A_27_47#_M1039_s N_VGND_c_1128_n 0.00397496f $X=1.84 $Y=0.235 $X2=0
+ $Y2=0
cc_614 N_A_27_47#_M1018_d N_VGND_c_1128_n 0.00225186f $X=2.7 $Y=0.235 $X2=0
+ $Y2=0
cc_615 N_A_27_47#_M1033_d N_VGND_c_1128_n 0.00215176f $X=3.56 $Y=0.235 $X2=0
+ $Y2=0
cc_616 N_A_27_47#_c_1055_n N_VGND_c_1128_n 0.0100304f $X=0.26 $Y=0.42 $X2=0
+ $Y2=0
cc_617 N_A_27_47#_c_1092_p N_VGND_c_1128_n 0.00730901f $X=1.12 $Y=0.42 $X2=0
+ $Y2=0
cc_618 N_A_27_47#_c_1090_p N_VGND_c_1128_n 0.00886411f $X=1.98 $Y=0.42 $X2=0
+ $Y2=0
cc_619 N_A_27_47#_c_1070_n N_A_454_47#_M1009_s 0.00329816f $X=2.71 $Y=0.955
+ $X2=-0.19 $Y2=-0.245
cc_620 N_A_27_47#_c_1074_n N_A_454_47#_M1032_s 0.00329816f $X=3.57 $Y=0.955
+ $X2=0 $Y2=0
cc_621 N_A_27_47#_M1018_d N_A_454_47#_c_1244_n 0.00354618f $X=2.7 $Y=0.235 $X2=0
+ $Y2=0
cc_622 N_A_27_47#_c_1070_n N_A_454_47#_c_1244_n 0.00485898f $X=2.71 $Y=0.955
+ $X2=0 $Y2=0
cc_623 N_A_27_47#_c_1074_n N_A_454_47#_c_1244_n 0.0179104f $X=3.57 $Y=0.955
+ $X2=0 $Y2=0
cc_624 N_A_27_47#_c_1079_n N_A_454_47#_c_1244_n 0.00981998f $X=2.84 $Y=0.83
+ $X2=0 $Y2=0
cc_625 N_A_27_47#_M1033_d N_A_454_47#_c_1243_n 0.00531926f $X=3.56 $Y=0.235
+ $X2=0 $Y2=0
cc_626 N_A_27_47#_c_1074_n N_A_454_47#_c_1243_n 0.00535657f $X=3.57 $Y=0.955
+ $X2=0 $Y2=0
cc_627 N_A_27_47#_c_1081_n N_A_454_47#_c_1243_n 0.014857f $X=3.7 $Y=0.83 $X2=0
+ $Y2=0
cc_628 N_A_27_47#_c_1070_n N_A_454_47#_c_1268_n 0.0130514f $X=2.71 $Y=0.955
+ $X2=0 $Y2=0
cc_629 N_VGND_c_1128_n N_A_454_47#_M1009_s 0.00280024f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_630 N_VGND_c_1128_n N_A_454_47#_M1032_s 0.0022356f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_631 N_VGND_c_1128_n N_A_454_47#_M1000_s 0.00223561f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_632 N_VGND_c_1128_n N_A_454_47#_M1028_s 0.00280024f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_633 N_VGND_c_1117_n N_A_454_47#_c_1244_n 0.0484998f $X=6.215 $Y=0 $X2=0 $Y2=0
cc_634 N_VGND_c_1128_n N_A_454_47#_c_1244_n 0.0311725f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_635 N_VGND_c_1117_n N_A_454_47#_c_1243_n 0.0828087f $X=6.215 $Y=0 $X2=0 $Y2=0
cc_636 N_VGND_c_1128_n N_A_454_47#_c_1243_n 0.050938f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_637 N_VGND_c_1117_n N_A_454_47#_c_1248_n 0.0486976f $X=6.215 $Y=0 $X2=0 $Y2=0
cc_638 N_VGND_c_1128_n N_A_454_47#_c_1248_n 0.0310694f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_639 N_VGND_c_1117_n N_A_454_47#_c_1268_n 0.0144063f $X=6.215 $Y=0 $X2=0 $Y2=0
cc_640 N_VGND_c_1128_n N_A_454_47#_c_1268_n 0.00973027f $X=9.84 $Y=0 $X2=0 $Y2=0
