* File: sky130_fd_sc_lp__o2111a_1.pxi.spice
* Created: Fri Aug 28 10:59:54 2020
* 
x_PM_SKY130_FD_SC_LP__O2111A_1%A_80_21# N_A_80_21#_M1005_s N_A_80_21#_M1010_d
+ N_A_80_21#_M1001_d N_A_80_21#_M1003_g N_A_80_21#_M1011_g N_A_80_21#_c_66_n
+ N_A_80_21#_c_67_n N_A_80_21#_c_68_n N_A_80_21#_c_75_p N_A_80_21#_c_104_p
+ N_A_80_21#_c_69_n N_A_80_21#_c_117_p N_A_80_21#_c_86_p N_A_80_21#_c_96_p
+ N_A_80_21#_c_118_p N_A_80_21#_c_70_n N_A_80_21#_c_81_p N_A_80_21#_c_71_n
+ PM_SKY130_FD_SC_LP__O2111A_1%A_80_21#
x_PM_SKY130_FD_SC_LP__O2111A_1%D1 N_D1_M1010_g N_D1_M1005_g D1 N_D1_c_135_n
+ PM_SKY130_FD_SC_LP__O2111A_1%D1
x_PM_SKY130_FD_SC_LP__O2111A_1%C1 N_C1_M1002_g N_C1_M1006_g C1 C1 C1 C1
+ N_C1_c_169_n N_C1_c_170_n PM_SKY130_FD_SC_LP__O2111A_1%C1
x_PM_SKY130_FD_SC_LP__O2111A_1%B1 N_B1_M1004_g N_B1_M1001_g B1 N_B1_c_209_n
+ N_B1_c_210_n PM_SKY130_FD_SC_LP__O2111A_1%B1
x_PM_SKY130_FD_SC_LP__O2111A_1%A2 N_A2_M1000_g N_A2_M1007_g A2 A2 N_A2_c_242_n
+ PM_SKY130_FD_SC_LP__O2111A_1%A2
x_PM_SKY130_FD_SC_LP__O2111A_1%A1 N_A1_M1009_g N_A1_M1008_g A1 N_A1_c_275_n
+ N_A1_c_276_n PM_SKY130_FD_SC_LP__O2111A_1%A1
x_PM_SKY130_FD_SC_LP__O2111A_1%X N_X_M1003_s N_X_M1011_s X X X X X X X
+ N_X_c_296_n PM_SKY130_FD_SC_LP__O2111A_1%X
x_PM_SKY130_FD_SC_LP__O2111A_1%VPWR N_VPWR_M1011_d N_VPWR_M1006_d N_VPWR_M1008_d
+ N_VPWR_c_310_n N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n
+ N_VPWR_c_332_n VPWR N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n
+ N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_309_n PM_SKY130_FD_SC_LP__O2111A_1%VPWR
x_PM_SKY130_FD_SC_LP__O2111A_1%VGND N_VGND_M1003_d N_VGND_M1000_d N_VGND_c_371_n
+ N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n VGND N_VGND_c_375_n
+ N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n PM_SKY130_FD_SC_LP__O2111A_1%VGND
x_PM_SKY130_FD_SC_LP__O2111A_1%A_517_49# N_A_517_49#_M1004_d N_A_517_49#_M1009_d
+ N_A_517_49#_c_422_n N_A_517_49#_c_419_n N_A_517_49#_c_420_n
+ N_A_517_49#_c_421_n PM_SKY130_FD_SC_LP__O2111A_1%A_517_49#
cc_1 VNB N_A_80_21#_M1011_g 0.00887657f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB N_A_80_21#_c_66_n 0.0115278f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.35
cc_3 VNB N_A_80_21#_c_67_n 0.0420003f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.35
cc_4 VNB N_A_80_21#_c_68_n 0.00326276f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.93
cc_5 VNB N_A_80_21#_c_69_n 0.0104472f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=0.42
cc_6 VNB N_A_80_21#_c_70_n 0.0259107f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.245
cc_7 VNB N_A_80_21#_c_71_n 0.0221055f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.185
cc_8 VNB N_D1_M1005_g 0.0284411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB D1 0.00798137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_D1_c_135_n 0.0284882f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_11 VNB N_C1_M1006_g 0.00636982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB C1 0.00422379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C1_c_169_n 0.0307041f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.35
cc_14 VNB N_C1_c_170_n 0.0162639f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.35
cc_15 VNB N_B1_M1004_g 0.0286697f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.835
cc_16 VNB N_B1_c_209_n 0.0020279f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_17 VNB N_B1_c_210_n 0.0343807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_M1000_g 0.027414f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.835
cc_19 VNB A2 0.00675347f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_20 VNB N_A2_c_242_n 0.0223079f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_21 VNB N_A1_M1009_g 0.0283203f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.835
cc_22 VNB N_A1_M1008_g 0.00137845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_275_n 0.0579531f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_24 VNB N_A1_c_276_n 0.0137708f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_25 VNB N_X_c_296_n 0.0621369f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.515
cc_26 VNB N_VPWR_c_309_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_371_n 0.0113576f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_28 VNB N_VGND_c_372_n 7.46595e-19 $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.515
cc_29 VNB N_VGND_c_373_n 0.0663794f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.35
cc_30 VNB N_VGND_c_374_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.35
cc_31 VNB N_VGND_c_375_n 0.0156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_376_n 0.0197377f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=2.015
cc_33 VNB N_VGND_c_377_n 0.250498f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=2.015
cc_34 VNB N_VGND_c_378_n 0.00500114f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=2.5
cc_35 VNB N_A_517_49#_c_419_n 0.0121597f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_36 VNB N_A_517_49#_c_420_n 0.00813124f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_37 VNB N_A_517_49#_c_421_n 0.0280982f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_38 VPB N_A_80_21#_M1011_g 0.0266493f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_39 VPB N_A_80_21#_c_68_n 0.00453994f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.93
cc_40 VPB N_D1_M1010_g 0.0218483f $X=-0.19 $Y=1.655 $X2=2.885 $Y2=1.835
cc_41 VPB D1 0.00467255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_D1_c_135_n 0.0075394f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_43 VPB N_C1_M1006_g 0.0227878f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB C1 0.0032835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_B1_M1001_g 0.0228528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_B1_c_209_n 0.0029989f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_47 VPB N_B1_c_210_n 0.0102865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_M1007_g 0.0187037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB A2 0.0119697f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_50 VPB N_A2_c_242_n 0.00624994f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_51 VPB N_A1_M1008_g 0.0228896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A1_c_276_n 0.012231f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_53 VPB N_X_c_296_n 0.0570269f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.515
cc_54 VPB N_VPWR_c_310_n 0.00227117f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_55 VPB N_VPWR_c_311_n 0.00345916f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.35
cc_56 VPB N_VPWR_c_312_n 0.00221918f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.35
cc_57 VPB N_VPWR_c_313_n 0.0150456f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.515
cc_58 VPB N_VPWR_c_314_n 0.0484195f $X=-0.19 $Y=1.655 $X2=1.66 $Y2=2.015
cc_59 VPB N_VPWR_c_315_n 0.0156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_316_n 0.0129398f $X=-0.19 $Y=1.655 $X2=3.095 $Y2=2.5
cc_61 VPB N_VPWR_c_317_n 0.0256244f $X=-0.19 $Y=1.655 $X2=1.755 $Y2=2.015
cc_62 VPB N_VPWR_c_318_n 0.0159762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_319_n 0.0117815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_309_n 0.0498577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_68_n N_D1_M1010_g 0.00539353f $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_75_p N_D1_M1010_g 0.0140214f $X=1.66 $Y=2.015 $X2=0 $Y2=0
cc_67 N_A_80_21#_c_69_n N_D1_M1005_g 0.0154988f $X=1.395 $Y=0.42 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_70_n N_D1_M1005_g 0.00984861f $X=1.06 $Y=1.245 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_68_n D1 0.0184943f $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_75_p D1 0.0214851f $X=1.66 $Y=2.015 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_70_n D1 0.0279374f $X=1.06 $Y=1.245 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_81_p D1 0.0120725f $X=1.755 $Y=2.015 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_67_n N_D1_c_135_n 0.0029114f $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_68_n N_D1_c_135_n 0.00111007f $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_75_p N_D1_c_135_n 6.84596e-19 $X=1.66 $Y=2.015 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_70_n N_D1_c_135_n 0.00820784f $X=1.06 $Y=1.245 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_86_p N_C1_M1006_g 0.0161441f $X=2.93 $Y=2.015 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_69_n C1 0.0249927f $X=1.395 $Y=0.42 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_86_p C1 0.0247074f $X=2.93 $Y=2.015 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_70_n C1 0.0065154f $X=1.06 $Y=1.245 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_86_p N_C1_c_169_n 6.61061e-19 $X=2.93 $Y=2.015 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_69_n N_C1_c_170_n 0.00249217f $X=1.395 $Y=0.42 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_70_n N_C1_c_170_n 4.65879e-19 $X=1.06 $Y=1.245 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_86_p N_B1_M1001_g 0.0185594f $X=2.93 $Y=2.015 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_86_p N_B1_c_209_n 0.0232666f $X=2.93 $Y=2.015 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_86_p N_B1_c_210_n 0.00289997f $X=2.93 $Y=2.015 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_96_p A2 0.0237279f $X=3.095 $Y=2.1 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_96_p N_A2_c_242_n 9.40088e-19 $X=3.095 $Y=2.1 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_66_n N_X_c_296_n 0.0269244f $X=0.975 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_68_n N_X_c_296_n 0.00950755f $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_70_n N_X_c_296_n 0.0038303f $X=1.06 $Y=1.245 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_71_n N_X_c_296_n 0.0267759f $X=0.597 $Y=1.185 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_68_n N_VPWR_M1011_d 0.00297253f $X=1.06 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_80_21#_c_75_p N_VPWR_M1011_d 0.0116245f $X=1.66 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A_80_21#_c_104_p N_VPWR_M1011_d 0.00509242f $X=1.145 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_96 N_A_80_21#_c_86_p N_VPWR_M1006_d 0.0184029f $X=2.93 $Y=2.015 $X2=0 $Y2=0
cc_97 N_A_80_21#_M1011_g N_VPWR_c_310_n 0.00517001f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_98 N_A_80_21#_c_66_n N_VPWR_c_310_n 0.0147857f $X=0.975 $Y=1.35 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_67_n N_VPWR_c_310_n 0.0052955f $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_68_n N_VPWR_c_310_n 0.00867205f $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_104_p N_VPWR_c_310_n 0.0142757f $X=1.145 $Y=2.015 $X2=0
+ $Y2=0
cc_102 N_A_80_21#_M1011_g N_VPWR_c_311_n 0.0101615f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_103 N_A_80_21#_c_86_p N_VPWR_c_312_n 0.0504347f $X=2.93 $Y=2.015 $X2=0 $Y2=0
cc_104 N_A_80_21#_M1011_g N_VPWR_c_332_n 0.00951683f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_105 N_A_80_21#_c_75_p N_VPWR_c_332_n 0.0231469f $X=1.66 $Y=2.015 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_104_p N_VPWR_c_332_n 0.0152373f $X=1.145 $Y=2.015 $X2=0
+ $Y2=0
cc_107 N_A_80_21#_M1011_g N_VPWR_c_315_n 0.00525069f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_A_80_21#_c_117_p N_VPWR_c_316_n 0.0124525f $X=1.755 $Y=2.47 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_118_p N_VPWR_c_317_n 0.0212513f $X=3.095 $Y=2.5 $X2=0 $Y2=0
cc_110 N_A_80_21#_M1010_d N_VPWR_c_309_n 0.00536646f $X=1.615 $Y=1.835 $X2=0
+ $Y2=0
cc_111 N_A_80_21#_M1001_d N_VPWR_c_309_n 0.00526034f $X=2.885 $Y=1.835 $X2=0
+ $Y2=0
cc_112 N_A_80_21#_M1011_g N_VPWR_c_309_n 0.00979769f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_80_21#_c_117_p N_VPWR_c_309_n 0.00730901f $X=1.755 $Y=2.47 $X2=0
+ $Y2=0
cc_114 N_A_80_21#_c_118_p N_VPWR_c_309_n 0.0127519f $X=3.095 $Y=2.5 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_66_n N_VGND_c_371_n 0.0227575f $X=0.975 $Y=1.35 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_67_n N_VGND_c_371_n 0.00553375f $X=0.63 $Y=1.35 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_69_n N_VGND_c_371_n 0.0358726f $X=1.395 $Y=0.42 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_71_n N_VGND_c_371_n 0.0155752f $X=0.597 $Y=1.185 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_69_n N_VGND_c_373_n 0.0210467f $X=1.395 $Y=0.42 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_71_n N_VGND_c_375_n 0.00525069f $X=0.597 $Y=1.185 $X2=0
+ $Y2=0
cc_121 N_A_80_21#_M1005_s N_VGND_c_377_n 0.00212301f $X=1.27 $Y=0.245 $X2=0
+ $Y2=0
cc_122 N_A_80_21#_c_69_n N_VGND_c_377_n 0.0125689f $X=1.395 $Y=0.42 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_71_n N_VGND_c_377_n 0.00979769f $X=0.597 $Y=1.185 $X2=0
+ $Y2=0
cc_124 N_D1_M1010_g N_C1_M1006_g 0.0177628f $X=1.54 $Y=2.465 $X2=0 $Y2=0
cc_125 N_D1_M1005_g C1 0.00347396f $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_126 D1 C1 0.0280694f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_127 N_D1_c_135_n C1 2.2502e-19 $X=1.49 $Y=1.51 $X2=0 $Y2=0
cc_128 D1 N_C1_c_169_n 0.00229792f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_129 N_D1_c_135_n N_C1_c_169_n 0.0464846f $X=1.49 $Y=1.51 $X2=0 $Y2=0
cc_130 N_D1_M1005_g N_C1_c_170_n 0.0464846f $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_131 N_D1_M1010_g N_VPWR_c_310_n 0.00318793f $X=1.54 $Y=2.465 $X2=0 $Y2=0
cc_132 N_D1_M1010_g N_VPWR_c_311_n 0.00902321f $X=1.54 $Y=2.465 $X2=0 $Y2=0
cc_133 N_D1_M1010_g N_VPWR_c_312_n 6.92059e-19 $X=1.54 $Y=2.465 $X2=0 $Y2=0
cc_134 N_D1_M1010_g N_VPWR_c_332_n 0.00991769f $X=1.54 $Y=2.465 $X2=0 $Y2=0
cc_135 N_D1_M1010_g N_VPWR_c_316_n 0.00486043f $X=1.54 $Y=2.465 $X2=0 $Y2=0
cc_136 N_D1_M1010_g N_VPWR_c_309_n 0.0082726f $X=1.54 $Y=2.465 $X2=0 $Y2=0
cc_137 N_D1_M1005_g N_VGND_c_371_n 0.00287921f $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_138 N_D1_M1005_g N_VGND_c_373_n 0.00539298f $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_139 N_D1_M1005_g N_VGND_c_377_n 0.0111162f $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_140 C1 N_B1_M1004_g 0.0135705f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_141 N_C1_c_169_n N_B1_M1004_g 0.0202453f $X=2.06 $Y=1.36 $X2=0 $Y2=0
cc_142 N_C1_c_170_n N_B1_M1004_g 0.0295795f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_143 N_C1_M1006_g N_B1_M1001_g 0.0112614f $X=1.97 $Y=2.465 $X2=0 $Y2=0
cc_144 C1 N_B1_M1001_g 2.11299e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_145 N_C1_M1006_g N_B1_c_209_n 3.36806e-19 $X=1.97 $Y=2.465 $X2=0 $Y2=0
cc_146 C1 N_B1_c_209_n 0.0331551f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_147 N_C1_M1006_g N_B1_c_210_n 0.00407215f $X=1.97 $Y=2.465 $X2=0 $Y2=0
cc_148 C1 A2 3.02628e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_149 N_C1_M1006_g N_VPWR_c_312_n 0.0172736f $X=1.97 $Y=2.465 $X2=0 $Y2=0
cc_150 N_C1_M1006_g N_VPWR_c_332_n 6.91782e-19 $X=1.97 $Y=2.465 $X2=0 $Y2=0
cc_151 N_C1_M1006_g N_VPWR_c_316_n 0.00486043f $X=1.97 $Y=2.465 $X2=0 $Y2=0
cc_152 N_C1_M1006_g N_VPWR_c_309_n 0.0082726f $X=1.97 $Y=2.465 $X2=0 $Y2=0
cc_153 C1 N_VGND_c_373_n 0.0111245f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_154 N_C1_c_170_n N_VGND_c_373_n 0.0048399f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_155 C1 N_VGND_c_377_n 0.0114793f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_156 N_C1_c_170_n N_VGND_c_377_n 0.00847353f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_157 C1 A_409_49# 0.0122009f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_158 C1 N_A_517_49#_c_422_n 0.0359541f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_159 N_C1_c_170_n N_A_517_49#_c_422_n 0.00108733f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_160 C1 N_A_517_49#_c_420_n 0.0103705f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_161 N_B1_M1004_g N_A2_M1000_g 0.00914214f $X=2.51 $Y=0.665 $X2=0 $Y2=0
cc_162 N_B1_M1001_g N_A2_M1007_g 0.0260551f $X=2.81 $Y=2.465 $X2=0 $Y2=0
cc_163 N_B1_c_209_n A2 0.0348358f $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_164 N_B1_c_210_n A2 0.00323651f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_165 N_B1_c_209_n N_A2_c_242_n 2.83062e-19 $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_166 N_B1_c_210_n N_A2_c_242_n 0.0208818f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_167 N_B1_M1001_g N_VPWR_c_312_n 0.0186379f $X=2.81 $Y=2.465 $X2=0 $Y2=0
cc_168 N_B1_M1001_g N_VPWR_c_317_n 0.00486043f $X=2.81 $Y=2.465 $X2=0 $Y2=0
cc_169 N_B1_M1001_g N_VPWR_c_309_n 0.00864313f $X=2.81 $Y=2.465 $X2=0 $Y2=0
cc_170 N_B1_M1004_g N_VGND_c_373_n 0.00539298f $X=2.51 $Y=0.665 $X2=0 $Y2=0
cc_171 N_B1_M1004_g N_VGND_c_377_n 0.0108811f $X=2.51 $Y=0.665 $X2=0 $Y2=0
cc_172 N_B1_M1004_g N_A_517_49#_c_422_n 0.0129702f $X=2.51 $Y=0.665 $X2=0 $Y2=0
cc_173 N_B1_M1004_g N_A_517_49#_c_420_n 0.00402623f $X=2.51 $Y=0.665 $X2=0 $Y2=0
cc_174 N_B1_c_209_n N_A_517_49#_c_420_n 0.0195889f $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_175 N_B1_c_210_n N_A_517_49#_c_420_n 0.00579177f $X=2.81 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A2_M1000_g N_A1_M1009_g 0.0252978f $X=3.28 $Y=0.665 $X2=0 $Y2=0
cc_177 N_A2_M1007_g N_A1_M1008_g 0.0566514f $X=3.35 $Y=2.465 $X2=0 $Y2=0
cc_178 A2 N_A1_M1008_g 0.00589031f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_179 A2 N_A1_c_275_n 0.00934403f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A2_c_242_n N_A1_c_275_n 0.0566514f $X=3.26 $Y=1.51 $X2=0 $Y2=0
cc_181 A2 N_A1_c_276_n 0.0345608f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_182 N_A2_M1007_g N_VPWR_c_312_n 0.00116001f $X=3.35 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A2_M1007_g N_VPWR_c_314_n 0.00466081f $X=3.35 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A2_M1007_g N_VPWR_c_317_n 0.00585385f $X=3.35 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A2_M1007_g N_VPWR_c_309_n 0.0109726f $X=3.35 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A2_M1000_g N_VGND_c_372_n 0.011586f $X=3.28 $Y=0.665 $X2=0 $Y2=0
cc_187 N_A2_M1000_g N_VGND_c_373_n 0.00477554f $X=3.28 $Y=0.665 $X2=0 $Y2=0
cc_188 N_A2_M1000_g N_VGND_c_377_n 0.00889934f $X=3.28 $Y=0.665 $X2=0 $Y2=0
cc_189 N_A2_M1000_g N_A_517_49#_c_419_n 0.0137639f $X=3.28 $Y=0.665 $X2=0 $Y2=0
cc_190 A2 N_A_517_49#_c_419_n 0.0415635f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A2_c_242_n N_A_517_49#_c_419_n 7.80086e-19 $X=3.26 $Y=1.51 $X2=0 $Y2=0
cc_192 A2 N_A_517_49#_c_420_n 0.0171162f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A2_c_242_n N_A_517_49#_c_420_n 5.01112e-19 $X=3.26 $Y=1.51 $X2=0 $Y2=0
cc_194 N_A1_M1008_g N_VPWR_c_314_n 0.0337522f $X=3.71 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A1_c_275_n N_VPWR_c_314_n 0.00319295f $X=4.03 $Y=1.46 $X2=0 $Y2=0
cc_196 N_A1_c_276_n N_VPWR_c_314_n 0.0198561f $X=4.03 $Y=1.46 $X2=0 $Y2=0
cc_197 N_A1_M1008_g N_VPWR_c_317_n 0.00368966f $X=3.71 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A1_M1008_g N_VPWR_c_309_n 0.00634462f $X=3.71 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A1_M1009_g N_VGND_c_372_n 0.011586f $X=3.71 $Y=0.665 $X2=0 $Y2=0
cc_200 N_A1_M1009_g N_VGND_c_376_n 0.00477554f $X=3.71 $Y=0.665 $X2=0 $Y2=0
cc_201 N_A1_M1009_g N_VGND_c_377_n 0.00929579f $X=3.71 $Y=0.665 $X2=0 $Y2=0
cc_202 N_A1_M1009_g N_A_517_49#_c_419_n 0.0165586f $X=3.71 $Y=0.665 $X2=0 $Y2=0
cc_203 N_A1_c_275_n N_A_517_49#_c_419_n 0.00889063f $X=4.03 $Y=1.46 $X2=0 $Y2=0
cc_204 N_A1_c_276_n N_A_517_49#_c_419_n 0.0193151f $X=4.03 $Y=1.46 $X2=0 $Y2=0
cc_205 N_X_c_296_n N_VPWR_c_310_n 0.050994f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_206 N_X_c_296_n N_VPWR_c_315_n 0.0181659f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_207 N_X_M1011_s N_VPWR_c_309_n 0.00336915f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_208 N_X_c_296_n N_VPWR_c_309_n 0.0104192f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_209 N_X_c_296_n N_VGND_c_375_n 0.0181659f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_210 N_X_M1003_s N_VGND_c_377_n 0.00336915f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_211 N_X_c_296_n N_VGND_c_377_n 0.0104192f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_212 N_VPWR_c_309_n A_685_367# 0.00900287f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_213 N_VGND_c_377_n A_337_49# 0.00899413f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_214 N_VGND_c_377_n A_409_49# 0.00785437f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_215 N_VGND_c_377_n N_A_517_49#_M1004_d 0.0065352f $X=4.08 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_216 N_VGND_c_377_n N_A_517_49#_M1009_d 0.00368844f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_373_n N_A_517_49#_c_422_n 0.0395943f $X=3.33 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_377_n N_A_517_49#_c_422_n 0.0230659f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_M1000_d N_A_517_49#_c_419_n 0.00176461f $X=3.355 $Y=0.245 $X2=0
+ $Y2=0
cc_220 N_VGND_c_372_n N_A_517_49#_c_419_n 0.0170777f $X=3.495 $Y=0.37 $X2=0
+ $Y2=0
cc_221 N_VGND_c_376_n N_A_517_49#_c_421_n 0.0178111f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_377_n N_A_517_49#_c_421_n 0.0100304f $X=4.08 $Y=0 $X2=0 $Y2=0
