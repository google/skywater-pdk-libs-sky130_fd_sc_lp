* File: sky130_fd_sc_lp__a221o_1.spice
* Created: Wed Sep  2 09:21:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a221o_1.pex.spice"
.subckt sky130_fd_sc_lp__a221o_1  VNB VPB A2 A1 B1 B2 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_80_21#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.2226 PD=1.46 PS=2.21 NRD=12.852 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1007 A_264_47# N_A2_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84 AD=0.1197
+ AS=0.2604 PD=1.125 PS=1.46 NRD=12.492 NRS=35.712 M=1 R=5.6 SA=75001 SB=75002.5
+ A=0.126 P=1.98 MULT=1
MM1009 N_A_80_21#_M1009_d N_A1_M1009_g A_264_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.336 AS=0.1197 PD=1.64 PS=1.125 NRD=17.856 NRS=12.492 M=1 R=5.6 SA=75001.4
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1010 A_541_47# N_B1_M1010_g N_A_80_21#_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.336 PD=1.05 PS=1.64 NRD=7.14 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_B2_M1004_g A_541_47# VNB NSHORT L=0.15 W=0.84 AD=0.189
+ AS=0.0882 PD=1.29 PS=1.05 NRD=12.852 NRS=7.14 M=1 R=5.6 SA=75002.7 SB=75000.8
+ A=0.126 P=1.98 MULT=1
MM1003 N_A_80_21#_M1003_d N_C1_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.189 PD=2.21 PS=1.29 NRD=0 NRS=11.424 M=1 R=5.6 SA=75003.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_VPWR_M1011_d N_A_80_21#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.3339 PD=1.88 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1008 N_A_264_367#_M1008_d N_A2_M1008_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.17955 AS=0.3906 PD=1.545 PS=1.88 NRD=0.7683 NRS=0 M=1 R=8.4
+ SA=75001 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_264_367#_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.17955 PD=3.05 PS=1.545 NRD=0 NRS=0 M=1 R=8.4 SA=75001.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_A_264_367#_M1005_d N_B1_M1005_g N_A_458_367#_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.3339 PD=1.62 PS=3.05 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_A_458_367#_M1006_d N_B2_M1006_g N_A_264_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.189 AS=0.2268 PD=1.56 PS=1.62 NRD=0.7683 NRS=1.5563 M=1 R=8.4
+ SA=75000.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_A_80_21#_M1000_d N_C1_M1000_g N_A_458_367#_M1006_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.189 PD=3.05 PS=1.56 NRD=0 NRS=2.3443 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
c_65 VPB 0 1.10918e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a221o_1.pxi.spice"
*
.ends
*
*
