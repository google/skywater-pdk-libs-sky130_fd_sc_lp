* File: sky130_fd_sc_lp__and2b_1.spice
* Created: Wed Sep  2 09:30:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and2b_1.pex.spice"
.subckt sky130_fd_sc_lp__and2b_1  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_N_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_300_131# N_A_27_47#_M1006_g N_A_217_131#_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g A_300_131# VNB NSHORT L=0.15 W=0.42 AD=0.098
+ AS=0.0441 PD=0.85 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_217_131#_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.196 PD=2.21 PS=1.7 NRD=0 NRS=11.064 M=1 R=5.6 SA=75000.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_A_N_M1007_g N_A_27_47#_M1007_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09345 AS=0.1113 PD=0.865 PS=1.37 NRD=37.5088 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1000 N_A_217_131#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.08505 AS=0.09345 PD=0.825 PS=0.865 NRD=39.8531 NRS=39.8531 M=1
+ R=2.8 SA=75000.8 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_A_217_131#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0987 AS=0.08505 PD=0.835 PS=0.825 NRD=0 NRS=18.7544 M=1 R=2.8 SA=75001.3
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_217_131#_M1002_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2961 PD=3.05 PS=2.505 NRD=0 NRS=6.7571 M=1 R=8.4 SA=75000.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__and2b_1.pxi.spice"
*
.ends
*
*
