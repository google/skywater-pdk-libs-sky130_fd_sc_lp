* File: sky130_fd_sc_lp__dfstp_2.pex.spice
* Created: Fri Aug 28 10:23:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFSTP_2%CLK 2 3 5 8 12 14 15 19
c43 8 0 6.03026e-20 $X=0.505 $Y=0.58
r44 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.09 $X2=0.525 $Y2=1.09
r45 19 21 3.69349 $w=2.61e-07 $l=2e-08 $layer=POLY_cond $X=0.505 $Y=1.09
+ $X2=0.525 $Y2=1.09
r46 15 22 6.14496 $w=4.07e-07 $l=2.05e-07 $layer=LI1_cond $X=0.642 $Y=1.295
+ $X2=0.642 $Y2=1.09
r47 14 22 4.94595 $w=4.07e-07 $l=1.65e-07 $layer=LI1_cond $X=0.642 $Y=0.925
+ $X2=0.642 $Y2=1.09
r48 10 12 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=0.23 $Y=2.14
+ $X2=0.475 $Y2=2.14
r49 6 19 15.717 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=0.925
+ $X2=0.505 $Y2=1.09
r50 6 8 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.505 $Y=0.925
+ $X2=0.505 $Y2=0.58
r51 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.215
+ $X2=0.475 $Y2=2.14
r52 3 5 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=2.215
+ $X2=0.475 $Y2=2.645
r53 2 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.23 $Y=2.065
+ $X2=0.23 $Y2=2.14
r54 1 19 50.7854 $w=2.61e-07 $l=3.47851e-07 $layer=POLY_cond $X=0.23 $Y=1.255
+ $X2=0.505 $Y2=1.09
r55 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.23 $Y=1.255 $X2=0.23
+ $Y2=2.065
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%D 1 2 3 4 5 7 8 10 13 16
c56 16 0 3.54564e-20 $X=1.49 $Y=1.97
c57 13 0 1.75573e-20 $X=1.68 $Y=2.035
c58 5 0 1.22143e-19 $X=1.925 $Y=1.125
c59 3 0 2.05317e-19 $X=1.85 $Y=2.13
r60 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.97 $X2=1.49 $Y2=1.97
r61 13 17 5.68738 $w=3.83e-07 $l=1.9e-07 $layer=LI1_cond $X=1.68 $Y=1.997
+ $X2=1.49 $Y2=1.997
r62 12 16 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.49 $Y=2.055
+ $X2=1.49 $Y2=1.97
r63 11 16 121.529 $w=3.3e-07 $l=6.95e-07 $layer=POLY_cond $X=1.49 $Y=1.275
+ $X2=1.49 $Y2=1.97
r64 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.925 $Y=2.205
+ $X2=1.925 $Y2=2.525
r65 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.925 $Y=1.125
+ $X2=1.925 $Y2=0.805
r66 4 12 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.655 $Y=2.13
+ $X2=1.49 $Y2=2.055
r67 3 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.85 $Y=2.13
+ $X2=1.925 $Y2=2.205
r68 3 4 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.85 $Y=2.13
+ $X2=1.655 $Y2=2.13
r69 2 11 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.655 $Y=1.2
+ $X2=1.49 $Y2=1.275
r70 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.85 $Y=1.2
+ $X2=1.925 $Y2=1.125
r71 1 2 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.85 $Y=1.2 $X2=1.655
+ $Y2=1.2
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_196_465# 1 2 9 11 13 15 19 23 25 26 30 32
+ 36 38 40 43 44 45 51 52 55 58 59 66
c181 58 0 1.12351e-19 $X=5.52 $Y=1.295
c182 44 0 1.77925e-19 $X=1.13 $Y=2.315
c183 40 0 6.03026e-20 $X=1.19 $Y=1.005
c184 26 0 1.96081e-19 $X=2.355 $Y=1.68
c185 25 0 3.43944e-20 $X=2.28 $Y=1.68
c186 11 0 8.73851e-20 $X=2.67 $Y=1.59
r187 64 66 23.9349 $w=2.92e-07 $l=1.45e-07 $layer=POLY_cond $X=5.57 $Y=1.51
+ $X2=5.715 $Y2=1.51
r188 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.57
+ $Y=1.51 $X2=5.57 $Y2=1.51
r189 59 65 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=5.57 $Y=1.295
+ $X2=5.57 $Y2=1.51
r190 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r191 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.295
+ $X2=1.2 $Y2=1.295
r192 52 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.295
+ $X2=1.2 $Y2=1.295
r193 51 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=5.52 $Y2=1.295
r194 51 52 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=1.345 $Y2=1.295
r195 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.68 $X2=2.03 $Y2=1.68
r196 45 48 8.31818 $w=1.78e-07 $l=1.35e-07 $layer=LI1_cond $X=2.035 $Y=1.545
+ $X2=2.035 $Y2=1.68
r197 42 55 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.19 $Y=1.455
+ $X2=1.19 $Y2=1.295
r198 42 43 3.89906 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=1.19 $Y=1.455 $X2=1.19
+ $Y2=1.545
r199 40 55 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.19 $Y=1.005
+ $X2=1.19 $Y2=1.295
r200 40 41 6.05995 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=1.005
+ $X2=1.19 $Y2=0.84
r201 39 43 2.54814 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.545
+ $X2=1.19 $Y2=1.545
r202 38 45 0.716491 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=1.945 $Y=1.545
+ $X2=2.035 $Y2=1.545
r203 38 39 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=1.945 $Y=1.545
+ $X2=1.355 $Y2=1.545
r204 36 41 10.7013 $w=2.78e-07 $l=2.6e-07 $layer=LI1_cond $X=1.215 $Y=0.58
+ $X2=1.215 $Y2=0.84
r205 30 44 5.98033 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=1.13 $Y=2.42
+ $X2=1.13 $Y2=2.315
r206 30 32 3.16883 $w=2.08e-07 $l=6e-08 $layer=LI1_cond $X=1.13 $Y=2.42 $X2=1.13
+ $Y2=2.48
r207 28 43 3.89906 $w=2.5e-07 $l=1.23693e-07 $layer=LI1_cond $X=1.11 $Y=1.635
+ $X2=1.19 $Y2=1.545
r208 28 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.11 $Y=1.635
+ $X2=1.11 $Y2=2.315
r209 25 49 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.28 $Y=1.68
+ $X2=2.03 $Y2=1.68
r210 25 26 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=2.28 $Y=1.68
+ $X2=2.355 $Y2=1.68
r211 21 66 16.5068 $w=2.92e-07 $l=2.09105e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.715 $Y2=1.51
r212 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.815 $Y2=2.335
r213 17 66 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.345
+ $X2=5.715 $Y2=1.51
r214 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.715 $Y=1.345
+ $X2=5.715 $Y2=0.555
r215 13 27 43.6381 $w=1.76e-07 $l=1.64697e-07 $layer=POLY_cond $X=2.785 $Y=1.435
+ $X2=2.765 $Y2=1.59
r216 13 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.785 $Y=1.435
+ $X2=2.785 $Y2=0.805
r217 12 26 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.43 $Y=1.59
+ $X2=2.355 $Y2=1.68
r218 11 27 6.61437 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=2.67 $Y=1.59
+ $X2=2.765 $Y2=1.59
r219 11 12 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.67 $Y=1.59
+ $X2=2.43 $Y2=1.59
r220 7 26 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.845
+ $X2=2.355 $Y2=1.68
r221 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.355 $Y=1.845
+ $X2=2.355 $Y2=2.525
r222 2 32 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.325 $X2=1.13 $Y2=2.48
r223 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.37 $X2=1.19 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_614_93# 1 2 9 14 16 19 21 24 26 27 31 36
+ 41 44 47
c84 36 0 1.09601e-19 $X=3.9 $Y=2.525
r85 45 47 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.145 $Y=1.455
+ $X2=3.145 $Y2=1.825
r86 38 41 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.87 $Y=0.445
+ $X2=3.995 $Y2=0.445
r87 33 36 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.72 $Y=2.525
+ $X2=3.9 $Y2=2.525
r88 31 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=1.29
+ $X2=3.235 $Y2=1.455
r89 31 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=1.29
+ $X2=3.235 $Y2=1.125
r90 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.235
+ $Y=1.29 $X2=3.235 $Y2=1.29
r91 27 30 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.235 $Y=1.1
+ $X2=3.235 $Y2=1.29
r92 25 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.87 $Y=0.61
+ $X2=3.87 $Y2=0.445
r93 25 26 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.87 $Y=0.61
+ $X2=3.87 $Y2=1.015
r94 24 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.72 $Y=2.36
+ $X2=3.72 $Y2=2.525
r95 23 24 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.72 $Y=2.155
+ $X2=3.72 $Y2=2.36
r96 22 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=1.1 $X2=3.235
+ $Y2=1.1
r97 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.785 $Y=1.1
+ $X2=3.87 $Y2=1.015
r98 21 22 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.785 $Y=1.1
+ $X2=3.4 $Y2=1.1
r99 19 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=1.99
+ $X2=3.235 $Y2=2.155
r100 19 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=1.99
+ $X2=3.235 $Y2=1.825
r101 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.235
+ $Y=1.99 $X2=3.235 $Y2=1.99
r102 16 23 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.635 $Y=2.025
+ $X2=3.72 $Y2=2.155
r103 16 18 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=3.635 $Y=2.025
+ $X2=3.235 $Y2=2.025
r104 14 48 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.145 $Y=2.525
+ $X2=3.145 $Y2=2.155
r105 9 44 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.145 $Y=0.805
+ $X2=3.145 $Y2=1.125
r106 2 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.76
+ $Y=2.315 $X2=3.9 $Y2=2.525
r107 1 41 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.87
+ $Y=0.235 $X2=3.995 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%SET_B 3 7 9 11 12 13 16 21 23 24 26 27 31 34
+ 35 36 37 38 64
c122 38 0 1.59619e-19 $X=7.44 $Y=1.665
c123 34 0 1.09601e-19 $X=4.14 $Y=1.99
c124 9 0 2.38286e-19 $X=6.98 $Y=0.985
r125 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.285
+ $Y=1.41 $X2=7.285 $Y2=1.41
r126 38 46 2.76705 $w=6.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.44 $Y=1.58
+ $X2=7.285 $Y2=1.58
r127 37 46 5.80187 $w=6.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.96 $Y=1.58
+ $X2=7.285 $Y2=1.58
r128 36 37 8.56892 $w=6.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.58
+ $X2=6.96 $Y2=1.58
r129 35 64 9.52743 $w=6.88e-07 $l=9.5e-08 $layer=LI1_cond $X=6 $Y=1.59 $X2=5.905
+ $Y2=1.59
r130 35 36 6.14854 $w=8.38e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=1.58
+ $X2=6.48 $Y2=1.58
r131 34 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.99
+ $X2=4.14 $Y2=2.155
r132 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.14
+ $Y=1.99 $X2=4.14 $Y2=1.99
r133 31 33 6.18841 $w=2.76e-07 $l=1.4e-07 $layer=LI1_cond $X=4.14 $Y=1.85
+ $X2=4.14 $Y2=1.99
r134 30 31 3.57235 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=1.85
+ $X2=4.14 $Y2=1.85
r135 30 64 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=4.305 $Y=1.85
+ $X2=5.905 $Y2=1.85
r136 27 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.66 $Y=1.07
+ $X2=4.66 $Y2=0.905
r137 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.66
+ $Y=1.07 $X2=4.66 $Y2=1.07
r138 24 26 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=4.305 $Y=1.11
+ $X2=4.66 $Y2=1.11
r139 23 31 5.54508 $w=2.76e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.22 $Y=1.765
+ $X2=4.14 $Y2=1.85
r140 22 24 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.22 $Y=1.235
+ $X2=4.305 $Y2=1.11
r141 22 23 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.22 $Y=1.235
+ $X2=4.22 $Y2=1.765
r142 21 45 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=7.285 $Y=1.765
+ $X2=7.285 $Y2=1.41
r143 14 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.865 $Y=1.915
+ $X2=7.865 $Y2=2.525
r144 13 21 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.45 $Y=1.84
+ $X2=7.285 $Y2=1.765
r145 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.79 $Y=1.84
+ $X2=7.865 $Y2=1.915
r146 12 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.79 $Y=1.84
+ $X2=7.45 $Y2=1.84
r147 9 45 63.9174 $w=2.3e-07 $l=5.57001e-07 $layer=POLY_cond $X=6.98 $Y=0.985
+ $X2=7.285 $Y2=1.41
r148 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.98 $Y=0.985
+ $X2=6.98 $Y2=0.665
r149 7 51 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.57 $Y=0.445
+ $X2=4.57 $Y2=0.905
r150 3 49 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.115 $Y=2.525
+ $X2=4.115 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_486_119# 1 2 9 13 15 19 22 23 25 26 27 28
+ 30 34 37 39 40 45 52 54
c148 39 0 1.40946e-20 $X=2.73 $Y=2.435
c149 37 0 1.22143e-19 $X=2.73 $Y=1.555
r150 54 57 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.78 $Y=1.45
+ $X2=3.78 $Y2=1.64
r151 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.45 $X2=3.78 $Y2=1.45
r152 43 45 8.3814 $w=2.18e-07 $l=1.6e-07 $layer=LI1_cond $X=2.57 $Y=0.725
+ $X2=2.73 $Y2=0.725
r153 41 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=1.64
+ $X2=2.73 $Y2=1.64
r154 40 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=1.64
+ $X2=3.78 $Y2=1.64
r155 40 41 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.615 $Y=1.64
+ $X2=2.815 $Y2=1.64
r156 39 48 6.70512 $w=2.73e-07 $l=1.6e-07 $layer=LI1_cond $X=2.73 $Y=2.572
+ $X2=2.57 $Y2=2.572
r157 38 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=1.725
+ $X2=2.73 $Y2=1.64
r158 38 39 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.73 $Y=1.725
+ $X2=2.73 $Y2=2.435
r159 37 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=1.555
+ $X2=2.73 $Y2=1.64
r160 36 45 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.73 $Y=0.835
+ $X2=2.73 $Y2=0.725
r161 36 37 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.73 $Y=0.835
+ $X2=2.73 $Y2=1.555
r162 32 34 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=5.11 $Y=1.06
+ $X2=5.355 $Y2=1.06
r163 29 30 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=4.865 $Y=1.54
+ $X2=5.11 $Y2=1.54
r164 27 55 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.135 $Y=1.45
+ $X2=3.78 $Y2=1.45
r165 27 28 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.135 $Y=1.45
+ $X2=4.21 $Y2=1.45
r166 26 55 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.76 $Y=1.45 $X2=3.78
+ $Y2=1.45
r167 23 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.355 $Y=0.985
+ $X2=5.355 $Y2=1.06
r168 23 25 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.355 $Y=0.985
+ $X2=5.355 $Y2=0.555
r169 22 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.11 $Y=1.465
+ $X2=5.11 $Y2=1.54
r170 21 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.11 $Y=1.135
+ $X2=5.11 $Y2=1.06
r171 21 22 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.11 $Y=1.135
+ $X2=5.11 $Y2=1.465
r172 17 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.865 $Y=1.615
+ $X2=4.865 $Y2=1.54
r173 17 19 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.865 $Y=1.615
+ $X2=4.865 $Y2=2.315
r174 16 28 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.285 $Y=1.54
+ $X2=4.21 $Y2=1.45
r175 15 29 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.79 $Y=1.54
+ $X2=4.865 $Y2=1.54
r176 15 16 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.79 $Y=1.54
+ $X2=4.285 $Y2=1.54
r177 11 28 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.285
+ $X2=4.21 $Y2=1.45
r178 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.21 $Y=1.285
+ $X2=4.21 $Y2=0.445
r179 7 26 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.685 $Y=1.615
+ $X2=3.76 $Y2=1.45
r180 7 9 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3.685 $Y=1.615
+ $X2=3.685 $Y2=2.525
r181 2 48 600 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=2.315 $X2=2.57 $Y2=2.545
r182 1 43 182 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.595 $X2=2.57 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_27_465# 1 2 10 14 15 16 17 18 21 25 27 31
+ 36 37 40 43 46 50 56 58 62
c143 62 0 1.75573e-20 $X=0.975 $Y=1.66
c144 50 0 3.54564e-20 $X=0.68 $Y=1.66
c145 31 0 1.12351e-19 $X=6.26 $Y=0.665
r146 61 62 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.905 $Y=1.66
+ $X2=0.975 $Y2=1.66
r147 53 56 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.175 $Y=0.575
+ $X2=0.27 $Y2=0.575
r148 51 61 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.68 $Y=1.66
+ $X2=0.905 $Y2=1.66
r149 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.68
+ $Y=1.66 $X2=0.68 $Y2=1.66
r150 48 58 0.926478 $w=2.5e-07 $l=1.38e-07 $layer=LI1_cond $X=0.365 $Y=1.7
+ $X2=0.227 $Y2=1.7
r151 48 50 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.365 $Y=1.7
+ $X2=0.68 $Y2=1.7
r152 44 58 5.68576 $w=2.22e-07 $l=1.25e-07 $layer=LI1_cond $X=0.227 $Y=1.825
+ $X2=0.227 $Y2=1.7
r153 44 46 27.03 $w=2.73e-07 $l=6.45e-07 $layer=LI1_cond $X=0.227 $Y=1.825
+ $X2=0.227 $Y2=2.47
r154 43 58 5.68576 $w=2.22e-07 $l=1.48745e-07 $layer=LI1_cond $X=0.175 $Y=1.575
+ $X2=0.227 $Y2=1.7
r155 42 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.175 $Y=0.74
+ $X2=0.175 $Y2=0.575
r156 42 43 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=0.175 $Y=0.74
+ $X2=0.175 $Y2=1.575
r157 38 40 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=6.26 $Y=1.94 $X2=6.36
+ $Y2=1.94
r158 34 36 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.36 $Y=3.075
+ $X2=6.36 $Y2=2.545
r159 33 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.36 $Y=2.015
+ $X2=6.36 $Y2=1.94
r160 33 36 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.36 $Y=2.015
+ $X2=6.36 $Y2=2.545
r161 29 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.26 $Y=1.865
+ $X2=6.26 $Y2=1.94
r162 29 31 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=6.26 $Y=1.865
+ $X2=6.26 $Y2=0.665
r163 28 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.86 $Y=3.15
+ $X2=2.785 $Y2=3.15
r164 27 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.285 $Y=3.15
+ $X2=6.36 $Y2=3.075
r165 27 28 1756.22 $w=1.5e-07 $l=3.425e-06 $layer=POLY_cond $X=6.285 $Y=3.15
+ $X2=2.86 $Y2=3.15
r166 23 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.785 $Y=3.075
+ $X2=2.785 $Y2=3.15
r167 23 25 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.785 $Y=3.075
+ $X2=2.785 $Y2=2.525
r168 19 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.355 $Y=0.255
+ $X2=2.355 $Y2=0.805
r169 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.28 $Y=0.18
+ $X2=2.355 $Y2=0.255
r170 17 18 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=2.28 $Y=0.18
+ $X2=1.05 $Y2=0.18
r171 15 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.71 $Y=3.15
+ $X2=2.785 $Y2=3.15
r172 15 16 887.085 $w=1.5e-07 $l=1.73e-06 $layer=POLY_cond $X=2.71 $Y=3.15
+ $X2=0.98 $Y2=3.15
r173 12 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.495
+ $X2=0.975 $Y2=1.66
r174 12 14 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=0.975 $Y=1.495
+ $X2=0.975 $Y2=0.58
r175 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.975 $Y=0.255
+ $X2=1.05 $Y2=0.18
r176 11 14 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.975 $Y=0.255
+ $X2=0.975 $Y2=0.58
r177 8 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=3.075
+ $X2=0.98 $Y2=3.15
r178 8 10 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.905 $Y=3.075
+ $X2=0.905 $Y2=2.645
r179 7 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.825
+ $X2=0.905 $Y2=1.66
r180 7 10 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.905 $Y=1.825
+ $X2=0.905 $Y2=2.645
r181 2 46 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.325 $X2=0.26 $Y2=2.47
r182 1 56 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.37 $X2=0.27 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_1309_65# 1 2 9 12 14 15 16 19 21 25 29 31
+ 33 37 40 45
c94 45 0 6.50956e-20 $X=7.955 $Y=0.57
c95 25 0 1.7319e-19 $X=6.835 $Y=1.55
c96 19 0 1.59619e-19 $X=7.435 $Y=2.525
c97 14 0 1.85795e-19 $X=6.945 $Y=3.075
r98 43 45 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.79 $Y=0.57
+ $X2=7.955 $Y2=0.57
r99 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.9 $Y=2.6
+ $X2=8.9 $Y2=2.6
r100 37 39 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=8.9 $Y=1.835
+ $X2=8.9 $Y2=2.6
r101 35 37 42.6055 $w=3.28e-07 $l=1.22e-06 $layer=LI1_cond $X=8.9 $Y=0.615
+ $X2=8.9 $Y2=1.835
r102 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.735 $Y=0.53
+ $X2=8.9 $Y2=0.615
r103 33 45 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=8.735 $Y=0.53
+ $X2=7.955 $Y2=0.53
r104 32 40 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=8.9 $Y=3.075
+ $X2=8.9 $Y2=2.6
r105 27 29 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=6.835 $Y=2.23
+ $X2=6.945 $Y2=2.23
r106 23 25 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=6.62 $Y=1.55
+ $X2=6.835 $Y2=1.55
r107 22 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.51 $Y=3.15
+ $X2=7.435 $Y2=3.15
r108 21 32 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.735 $Y=3.15
+ $X2=8.9 $Y2=3.075
r109 21 22 628.138 $w=1.5e-07 $l=1.225e-06 $layer=POLY_cond $X=8.735 $Y=3.15
+ $X2=7.51 $Y2=3.15
r110 17 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.435 $Y=3.075
+ $X2=7.435 $Y2=3.15
r111 17 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.435 $Y=3.075
+ $X2=7.435 $Y2=2.525
r112 15 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.36 $Y=3.15
+ $X2=7.435 $Y2=3.15
r113 15 16 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.36 $Y=3.15
+ $X2=7.02 $Y2=3.15
r114 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.945 $Y=3.075
+ $X2=7.02 $Y2=3.15
r115 13 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.945 $Y=2.305
+ $X2=6.945 $Y2=2.23
r116 13 14 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=6.945 $Y=2.305
+ $X2=6.945 $Y2=3.075
r117 12 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.835 $Y=2.155
+ $X2=6.835 $Y2=2.23
r118 11 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.835 $Y=1.625
+ $X2=6.835 $Y2=1.55
r119 11 12 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.835 $Y=1.625
+ $X2=6.835 $Y2=2.155
r120 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.62 $Y=1.475
+ $X2=6.62 $Y2=1.55
r121 7 9 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.62 $Y=1.475 $X2=6.62
+ $Y2=0.665
r122 2 37 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.74
+ $Y=1.625 $X2=8.88 $Y2=1.835
r123 1 43 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=7.63
+ $Y=0.455 $X2=7.79 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_1158_47# 1 2 3 10 12 13 14 17 19 22 24 25
+ 26 27 28 31 33 35 38 39 42 50 51 52 56 58 59 60 61 62 66
c142 61 0 1.85795e-19 $X=6.35 $Y=2.22
r143 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.45
+ $Y=0.96 $X2=8.45 $Y2=0.96
r144 63 65 0.231499 $w=5.27e-07 $l=1e-08 $layer=LI1_cond $X=8.255 $Y=0.95
+ $X2=8.255 $Y2=0.96
r145 60 61 5.55755 $w=2.38e-07 $l=9.5e-08 $layer=LI1_cond $X=6.255 $Y=2.22
+ $X2=6.35 $Y2=2.22
r146 59 62 3.98977 $w=2.3e-07 $l=8.9861e-08 $layer=LI1_cond $X=8.085 $Y=2.095
+ $X2=8.075 $Y2=2.18
r147 58 65 15.9347 $w=5.27e-07 $l=5.83845e-07 $layer=LI1_cond $X=8.085 $Y=1.465
+ $X2=8.255 $Y2=0.96
r148 58 59 33.0018 $w=2.18e-07 $l=6.3e-07 $layer=LI1_cond $X=8.085 $Y=1.465
+ $X2=8.085 $Y2=2.095
r149 54 62 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.075 $Y=2.265
+ $X2=8.075 $Y2=2.18
r150 54 56 12.4848 $w=2.38e-07 $l=2.6e-07 $layer=LI1_cond $X=8.075 $Y=2.265
+ $X2=8.075 $Y2=2.525
r151 52 62 2.45049 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.955 $Y=2.18
+ $X2=8.075 $Y2=2.18
r152 52 61 104.711 $w=1.68e-07 $l=1.605e-06 $layer=LI1_cond $X=7.955 $Y=2.18
+ $X2=6.35 $Y2=2.18
r153 50 63 7.48814 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=7.975 $Y=0.95
+ $X2=8.255 $Y2=0.95
r154 50 51 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=7.975 $Y=0.95
+ $X2=6.115 $Y2=0.95
r155 48 60 7.92305 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=6.09 $Y=2.225
+ $X2=6.255 $Y2=2.225
r156 42 45 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.95 $Y=0.39
+ $X2=5.95 $Y2=0.73
r157 40 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.95 $Y=0.865
+ $X2=6.115 $Y2=0.95
r158 40 45 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.95 $Y=0.865
+ $X2=5.95 $Y2=0.73
r159 37 66 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=8.45 $Y=1.315
+ $X2=8.45 $Y2=0.96
r160 37 38 13.5877 $w=2.4e-07 $l=1.01366e-07 $layer=POLY_cond $X=8.45 $Y=1.315
+ $X2=8.512 $Y2=1.39
r161 36 66 107.54 $w=3.3e-07 $l=6.15e-07 $layer=POLY_cond $X=8.45 $Y=0.345
+ $X2=8.45 $Y2=0.96
r162 33 35 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.615 $Y=1.875
+ $X2=9.615 $Y2=2.305
r163 29 31 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.615 $Y=0.795
+ $X2=9.615 $Y2=0.445
r164 27 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.54 $Y=1.8
+ $X2=9.615 $Y2=1.875
r165 27 28 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=9.54 $Y=1.8
+ $X2=9.23 $Y2=1.8
r166 25 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.54 $Y=0.87
+ $X2=9.615 $Y2=0.795
r167 25 26 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=9.54 $Y=0.87
+ $X2=9.23 $Y2=0.87
r168 24 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.155 $Y=1.725
+ $X2=9.23 $Y2=1.8
r169 23 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.155 $Y=1.465
+ $X2=9.155 $Y2=1.39
r170 23 24 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=9.155 $Y=1.465
+ $X2=9.155 $Y2=1.725
r171 22 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.155 $Y=1.315
+ $X2=9.155 $Y2=1.39
r172 21 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.155 $Y=0.945
+ $X2=9.23 $Y2=0.87
r173 21 22 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.155 $Y=0.945
+ $X2=9.155 $Y2=1.315
r174 20 38 12.1617 $w=1.5e-07 $l=2.28e-07 $layer=POLY_cond $X=8.74 $Y=1.39
+ $X2=8.512 $Y2=1.39
r175 19 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.08 $Y=1.39
+ $X2=9.155 $Y2=1.39
r176 19 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=9.08 $Y=1.39
+ $X2=8.74 $Y2=1.39
r177 15 38 13.5877 $w=2.4e-07 $l=1.86773e-07 $layer=POLY_cond $X=8.665 $Y=1.465
+ $X2=8.512 $Y2=1.39
r178 15 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.665 $Y=1.465
+ $X2=8.665 $Y2=1.835
r179 13 36 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.285 $Y=0.27
+ $X2=8.45 $Y2=0.345
r180 13 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=8.285 $Y=0.27
+ $X2=7.63 $Y2=0.27
r181 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.555 $Y=0.345
+ $X2=7.63 $Y2=0.27
r182 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.555 $Y=0.345
+ $X2=7.555 $Y2=0.665
r183 3 56 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.94
+ $Y=2.315 $X2=8.08 $Y2=2.525
r184 2 48 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=2.125 $X2=6.09 $Y2=2.25
r185 1 45 182 $w=1.7e-07 $l=5.69408e-07 $layer=licon1_NDIFF $count=1 $X=5.79
+ $Y=0.235 $X2=5.95 $Y2=0.73
r186 1 42 182 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_NDIFF $count=1 $X=5.79
+ $Y=0.235 $X2=5.95 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_1855_47# 1 2 9 12 14 16 18 21 23 26 30 34
+ 37 38 39
r68 38 39 32.8921 $w=3.95e-07 $l=7.5e-08 $layer=POLY_cond $X=10.002 $Y=1.26
+ $X2=10.002 $Y2=1.185
r69 35 41 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=10.002 $Y=1.35
+ $X2=10.002 $Y2=1.515
r70 35 38 12.6719 $w=3.95e-07 $l=9e-08 $layer=POLY_cond $X=10.002 $Y=1.35
+ $X2=10.002 $Y2=1.26
r71 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.97
+ $Y=1.35 $X2=9.97 $Y2=1.35
r72 32 37 0.695019 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=9.515 $Y=1.35
+ $X2=9.375 $Y2=1.35
r73 32 34 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=9.515 $Y=1.35
+ $X2=9.97 $Y2=1.35
r74 28 37 5.99569 $w=2.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=9.37 $Y=1.515
+ $X2=9.375 $Y2=1.35
r75 28 30 26.2501 $w=2.68e-07 $l=6.15e-07 $layer=LI1_cond $X=9.37 $Y=1.515
+ $X2=9.37 $Y2=2.13
r76 24 37 5.99569 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=9.375 $Y=1.185
+ $X2=9.375 $Y2=1.35
r77 24 26 31.4864 $w=2.78e-07 $l=7.65e-07 $layer=LI1_cond $X=9.375 $Y=1.185
+ $X2=9.375 $Y2=0.42
r78 19 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.555 $Y=1.335
+ $X2=10.555 $Y2=1.26
r79 19 21 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=10.555 $Y=1.335
+ $X2=10.555 $Y2=2.465
r80 16 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.555 $Y=1.185
+ $X2=10.555 $Y2=1.26
r81 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.555 $Y=1.185
+ $X2=10.555 $Y2=0.655
r82 15 38 25.5547 $w=1.5e-07 $l=1.98e-07 $layer=POLY_cond $X=10.2 $Y=1.26
+ $X2=10.002 $Y2=1.26
r83 14 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.48 $Y=1.26
+ $X2=10.555 $Y2=1.26
r84 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.48 $Y=1.26
+ $X2=10.2 $Y2=1.26
r85 12 41 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=10.125 $Y=2.465
+ $X2=10.125 $Y2=1.515
r86 9 39 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.125 $Y=0.655
+ $X2=10.125 $Y2=1.185
r87 2 30 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=9.275
+ $Y=1.985 $X2=9.4 $Y2=2.13
r88 1 26 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=9.275
+ $Y=0.235 $X2=9.4 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%VPWR 1 2 3 4 5 6 7 8 27 31 35 37 38 41 43 47
+ 51 53 55 60 61 63 64 67 68 69 75 86 97 102 108 111 114 117 121
c139 31 0 3.43944e-20 $X=1.71 $Y=2.525
r140 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r141 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r142 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r143 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r144 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r145 106 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r146 106 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r147 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r148 103 117 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=9.935 $Y=3.33
+ $X2=9.83 $Y2=3.33
r149 103 105 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.935 $Y=3.33
+ $X2=10.32 $Y2=3.33
r150 102 120 4.47956 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=10.635 $Y=3.33
+ $X2=10.837 $Y2=3.33
r151 102 105 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.635 $Y=3.33
+ $X2=10.32 $Y2=3.33
r152 101 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r153 101 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.4 $Y2=3.33
r154 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r155 98 114 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=8.565 $Y=3.33
+ $X2=8.465 $Y2=3.33
r156 98 100 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=8.565 $Y=3.33
+ $X2=9.36 $Y2=3.33
r157 97 117 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=9.725 $Y=3.33
+ $X2=9.83 $Y2=3.33
r158 97 100 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.725 $Y=3.33
+ $X2=9.36 $Y2=3.33
r159 96 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r160 95 96 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r161 93 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r162 92 95 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r163 92 93 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r164 90 111 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=4.455 $Y2=3.33
r165 90 92 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=5.04 $Y2=3.33
r166 89 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r167 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r168 86 111 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=4.165 $Y=3.33
+ $X2=4.455 $Y2=3.33
r169 86 88 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=3.33
+ $X2=4.08 $Y2=3.33
r170 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r171 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r172 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r173 82 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r174 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r175 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r176 79 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.71 $Y2=3.33
r177 79 81 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=2.16 $Y2=3.33
r178 78 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r179 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r180 75 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.71 $Y2=3.33
r181 75 77 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r182 73 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r183 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r184 69 96 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=7.44 $Y2=3.33
r185 69 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r186 67 95 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.555 $Y=3.33
+ $X2=7.44 $Y2=3.33
r187 67 68 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.555 $Y=3.33
+ $X2=7.67 $Y2=3.33
r188 63 84 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.12 $Y2=3.33
r189 63 64 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.33 $Y2=3.33
r190 62 88 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=4.08 $Y2=3.33
r191 62 64 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.33 $Y2=3.33
r192 60 72 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.24 $Y2=3.33
r193 60 61 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.69 $Y2=3.33
r194 59 77 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=1.2 $Y2=3.33
r195 59 61 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.69 $Y2=3.33
r196 55 58 37.2623 $w=2.98e-07 $l=9.7e-07 $layer=LI1_cond $X=10.785 $Y=1.98
+ $X2=10.785 $Y2=2.95
r197 53 120 3.03811 $w=3e-07 $l=1.07912e-07 $layer=LI1_cond $X=10.785 $Y=3.245
+ $X2=10.837 $Y2=3.33
r198 53 58 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=10.785 $Y=3.245
+ $X2=10.785 $Y2=2.95
r199 49 117 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=9.83 $Y=3.245
+ $X2=9.83 $Y2=3.33
r200 49 51 58.3593 $w=2.08e-07 $l=1.105e-06 $layer=LI1_cond $X=9.83 $Y=3.245
+ $X2=9.83 $Y2=2.14
r201 45 114 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=3.245
+ $X2=8.465 $Y2=3.33
r202 45 47 78.1909 $w=1.98e-07 $l=1.41e-06 $layer=LI1_cond $X=8.465 $Y=3.245
+ $X2=8.465 $Y2=1.835
r203 44 68 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.785 $Y=3.33
+ $X2=7.67 $Y2=3.33
r204 43 114 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=8.465 $Y2=3.33
r205 43 44 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=7.785 $Y2=3.33
r206 39 68 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=3.245
+ $X2=7.67 $Y2=3.33
r207 39 41 32.3185 $w=2.28e-07 $l=6.45e-07 $layer=LI1_cond $X=7.67 $Y=3.245
+ $X2=7.67 $Y2=2.6
r208 38 111 2.44113 $w=5.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=3.245
+ $X2=4.455 $Y2=3.33
r209 37 66 8.83446 $w=5.8e-07 $l=4.6744e-07 $layer=LI1_cond $X=4.455 $Y=2.65
+ $X2=4.65 $Y2=2.27
r210 37 38 12.2701 $w=5.78e-07 $l=5.95e-07 $layer=LI1_cond $X=4.455 $Y=2.65
+ $X2=4.455 $Y2=3.245
r211 33 64 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=3.245
+ $X2=3.33 $Y2=3.33
r212 33 35 30.7318 $w=2.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.33 $Y=3.245
+ $X2=3.33 $Y2=2.525
r213 29 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=3.33
r214 29 31 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=2.525
r215 25 61 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r216 25 27 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.48
r217 8 58 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.835 $X2=10.77 $Y2=2.95
r218 8 55 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.835 $X2=10.77 $Y2=1.98
r219 7 51 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=9.69
+ $Y=1.985 $X2=9.83 $Y2=2.14
r220 6 47 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=8.325
+ $Y=1.625 $X2=8.45 $Y2=1.835
r221 5 41 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=7.51
+ $Y=2.315 $X2=7.65 $Y2=2.6
r222 4 66 300 $w=1.7e-07 $l=4.81975e-07 $layer=licon1_PDIFF $count=2 $X=4.19
+ $Y=2.315 $X2=4.65 $Y2=2.27
r223 3 35 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=3.22
+ $Y=2.315 $X2=3.37 $Y2=2.525
r224 2 31 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=2.315 $X2=1.71 $Y2=2.525
r225 1 27 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.325 $X2=0.69 $Y2=2.48
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_400_119# 1 2 9 13 16 19 23
c45 23 0 8.73851e-20 $X=2.38 $Y=2.18
c46 19 0 1.96081e-19 $X=2.38 $Y=1.09
c47 16 0 1.91223e-19 $X=2.38 $Y=2.095
r48 21 23 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.14 $Y=2.18
+ $X2=2.38 $Y2=2.18
r49 16 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=2.095
+ $X2=2.38 $Y2=2.18
r50 15 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=1.175
+ $X2=2.38 $Y2=1.09
r51 15 16 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.38 $Y=1.175
+ $X2=2.38 $Y2=2.095
r52 11 21 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.265
+ $X2=2.14 $Y2=2.18
r53 11 13 15.177 $w=1.88e-07 $l=2.6e-07 $layer=LI1_cond $X=2.14 $Y=2.265
+ $X2=2.14 $Y2=2.525
r54 7 19 16.8321 $w=1.68e-07 $l=2.58e-07 $layer=LI1_cond $X=2.122 $Y=1.09
+ $X2=2.38 $Y2=1.09
r55 7 9 10.2439 $w=2.23e-07 $l=2e-07 $layer=LI1_cond $X=2.122 $Y=1.005 $X2=2.122
+ $Y2=0.805
r56 2 13 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=2.315 $X2=2.14 $Y2=2.525
r57 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.595
+ $X2=2.14 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_988_379# 1 2 9 11 13
r27 11 13 79.0227 $w=1.98e-07 $l=1.425e-06 $layer=LI1_cond $X=5.245 $Y=2.955
+ $X2=6.67 $Y2=2.955
r28 7 11 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=5.08 $Y=2.855
+ $X2=5.245 $Y2=2.955
r29 7 9 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=5.08 $Y=2.855
+ $X2=5.08 $Y2=2.19
r30 2 13 600 $w=1.7e-07 $l=9.35147e-07 $layer=licon1_PDIFF $count=1 $X=6.435
+ $Y=2.125 $X2=6.67 $Y2=2.95
r31 1 9 300 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=2 $X=4.94
+ $Y=1.895 $X2=5.08 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%A_1095_425# 1 2 9 12 14 15
r25 14 15 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.22 $Y=2.56
+ $X2=7.055 $Y2=2.56
r26 12 15 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.71 $Y=2.6
+ $X2=7.055 $Y2=2.6
r27 7 12 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=5.572 $Y=2.515
+ $X2=5.71 $Y2=2.6
r28 7 9 7.54326 $w=2.73e-07 $l=1.8e-07 $layer=LI1_cond $X=5.572 $Y=2.515
+ $X2=5.572 $Y2=2.335
r29 2 14 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=7.095
+ $Y=2.315 $X2=7.22 $Y2=2.54
r30 1 9 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=5.475
+ $Y=2.125 $X2=5.6 $Y2=2.335
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%Q 1 2 7 8 9 10 11 12 13 22
r16 13 40 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=10.345 $Y=2.775
+ $X2=10.345 $Y2=2.91
r17 12 13 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=2.405
+ $X2=10.345 $Y2=2.775
r18 11 12 18.7272 $w=2.38e-07 $l=3.9e-07 $layer=LI1_cond $X=10.345 $Y=2.015
+ $X2=10.345 $Y2=2.405
r19 10 11 16.8065 $w=2.38e-07 $l=3.5e-07 $layer=LI1_cond $X=10.345 $Y=1.665
+ $X2=10.345 $Y2=2.015
r20 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=1.295
+ $X2=10.345 $Y2=1.665
r21 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=0.925
+ $X2=10.345 $Y2=1.295
r22 7 8 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=0.555
+ $X2=10.345 $Y2=0.925
r23 7 22 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=10.345 $Y=0.555
+ $X2=10.345 $Y2=0.42
r24 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.2
+ $Y=1.835 $X2=10.34 $Y2=2.91
r25 2 11 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=10.2 $Y=1.835
+ $X2=10.34 $Y2=2.015
r26 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=10.2
+ $Y=0.235 $X2=10.34 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 43 46 48
+ 50 53 54 56 57 59 61 63 68 80 94 101 107 110 113 116 120
r135 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r136 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r137 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r138 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r139 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r140 105 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r141 105 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r142 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r143 102 116 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=10.055 $Y=0
+ $X2=9.87 $Y2=0
r144 102 104 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=10.055 $Y=0
+ $X2=10.32 $Y2=0
r145 101 119 4.47956 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.837 $Y2=0
r146 101 104 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.32 $Y2=0
r147 100 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r148 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r149 97 100 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=9.36 $Y2=0
r150 96 99 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.44 $Y=0 $X2=9.36
+ $Y2=0
r151 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r152 94 116 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=9.685 $Y=0
+ $X2=9.87 $Y2=0
r153 94 99 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.685 $Y=0
+ $X2=9.36 $Y2=0
r154 93 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r155 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r156 89 92 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=6.96
+ $Y2=0
r157 87 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0
+ $X2=5.06 $Y2=0
r158 87 89 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.52
+ $Y2=0
r159 86 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r160 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r161 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r162 82 85 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r163 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r164 80 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=5.06 $Y2=0
r165 80 85 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=4.56 $Y2=0
r166 79 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r167 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r168 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r169 76 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r170 75 78 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r171 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r172 73 110 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.84 $Y=0
+ $X2=1.692 $Y2=0
r173 73 75 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=2.16
+ $Y2=0
r174 72 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r175 72 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r176 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r177 69 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.74 $Y2=0
r178 69 71 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.2
+ $Y2=0
r179 68 110 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=1.545 $Y=0
+ $X2=1.692 $Y2=0
r180 68 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r181 66 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r182 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r183 63 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0
+ $X2=0.74 $Y2=0
r184 63 65 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0
+ $X2=0.24 $Y2=0
r185 61 93 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.96 $Y2=0
r186 61 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r187 61 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r188 59 60 5.47614 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.87 $Y=0.38
+ $X2=9.87 $Y2=0.545
r189 56 92 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=7.03 $Y=0 $X2=6.96
+ $Y2=0
r190 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.03 $Y=0 $X2=7.195
+ $Y2=0
r191 55 96 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.36 $Y=0 $X2=7.44
+ $Y2=0
r192 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.36 $Y=0 $X2=7.195
+ $Y2=0
r193 53 78 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.195 $Y=0 $X2=3.12
+ $Y2=0
r194 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=0 $X2=3.36
+ $Y2=0
r195 52 82 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.525 $Y=0 $X2=3.6
+ $Y2=0
r196 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=0 $X2=3.36
+ $Y2=0
r197 48 119 3.03811 $w=3e-07 $l=1.07912e-07 $layer=LI1_cond $X=10.785 $Y=0.085
+ $X2=10.837 $Y2=0
r198 48 50 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=10.785 $Y=0.085
+ $X2=10.785 $Y2=0.38
r199 46 60 11.3386 $w=3.08e-07 $l=3.05e-07 $layer=LI1_cond $X=9.9 $Y=0.85
+ $X2=9.9 $Y2=0.545
r200 43 59 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=9.87 $Y=0.36
+ $X2=9.87 $Y2=0.38
r201 42 116 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.87 $Y=0.085
+ $X2=9.87 $Y2=0
r202 42 43 8.56545 $w=3.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.87 $Y=0.085
+ $X2=9.87 $Y2=0.36
r203 38 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.195 $Y=0.085
+ $X2=7.195 $Y2=0
r204 38 40 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=7.195 $Y=0.085
+ $X2=7.195 $Y2=0.58
r205 34 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0
r206 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0.38
r207 30 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=0.085
+ $X2=3.36 $Y2=0
r208 30 32 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.36 $Y=0.085
+ $X2=3.36 $Y2=0.74
r209 26 110 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.692 $Y=0.085
+ $X2=1.692 $Y2=0
r210 26 28 28.1274 $w=2.93e-07 $l=7.2e-07 $layer=LI1_cond $X=1.692 $Y=0.085
+ $X2=1.692 $Y2=0.805
r211 22 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r212 22 24 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.545
r213 7 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.63
+ $Y=0.235 $X2=10.77 $Y2=0.38
r214 6 59 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=9.69
+ $Y=0.235 $X2=9.85 $Y2=0.38
r215 6 46 182 $w=1.7e-07 $l=7.16607e-07 $layer=licon1_NDIFF $count=1 $X=9.69
+ $Y=0.235 $X2=9.91 $Y2=0.85
r216 5 40 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=7.055
+ $Y=0.455 $X2=7.195 $Y2=0.58
r217 4 36 91 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_NDIFF $count=2 $X=4.645
+ $Y=0.235 $X2=5.06 $Y2=0.38
r218 3 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.595 $X2=3.36 $Y2=0.74
r219 2 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.595 $X2=1.71 $Y2=0.805
r220 1 24 182 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.37 $X2=0.74 $Y2=0.545
.ends

