* File: sky130_fd_sc_lp__einvn_0.pxi.spice
* Created: Fri Aug 28 10:32:33 2020
* 
x_PM_SKY130_FD_SC_LP__EINVN_0%A_28_141# N_A_28_141#_M1004_s N_A_28_141#_M1001_s
+ N_A_28_141#_c_35_n N_A_28_141#_M1005_g N_A_28_141#_c_36_n N_A_28_141#_c_37_n
+ N_A_28_141#_c_38_n N_A_28_141#_c_39_n PM_SKY130_FD_SC_LP__EINVN_0%A_28_141#
x_PM_SKY130_FD_SC_LP__EINVN_0%TE_B N_TE_B_M1004_g N_TE_B_c_73_n N_TE_B_M1001_g
+ N_TE_B_M1003_g N_TE_B_c_76_n TE_B TE_B TE_B N_TE_B_c_72_n
+ PM_SKY130_FD_SC_LP__EINVN_0%TE_B
x_PM_SKY130_FD_SC_LP__EINVN_0%A N_A_M1002_g N_A_M1000_g A A A A A N_A_c_116_n
+ PM_SKY130_FD_SC_LP__EINVN_0%A
x_PM_SKY130_FD_SC_LP__EINVN_0%VPWR N_VPWR_M1001_d N_VPWR_c_152_n VPWR
+ N_VPWR_c_153_n N_VPWR_c_154_n N_VPWR_c_151_n N_VPWR_c_156_n
+ PM_SKY130_FD_SC_LP__EINVN_0%VPWR
x_PM_SKY130_FD_SC_LP__EINVN_0%Z N_Z_M1002_d N_Z_M1000_d Z Z Z Z Z Z
+ PM_SKY130_FD_SC_LP__EINVN_0%Z
x_PM_SKY130_FD_SC_LP__EINVN_0%VGND N_VGND_M1004_d N_VGND_c_192_n N_VGND_c_187_n
+ VGND N_VGND_c_188_n N_VGND_c_189_n N_VGND_c_190_n N_VGND_c_191_n
+ PM_SKY130_FD_SC_LP__EINVN_0%VGND
cc_1 VNB N_A_28_141#_c_35_n 0.021204f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.595
cc_2 VNB N_A_28_141#_c_36_n 0.0430039f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.915
cc_3 VNB N_A_28_141#_c_37_n 0.0183964f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=0.43
cc_4 VNB N_A_28_141#_c_38_n 0.0064136f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.43
cc_5 VNB N_A_28_141#_c_39_n 0.0429677f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.43
cc_6 VNB N_TE_B_M1004_g 0.04092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB TE_B 0.00836194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_TE_B_c_72_n 0.0209459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_M1002_g 0.0365041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A 0.00537642f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.915
cc_11 VNB N_A_c_116_n 0.0197192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_151_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.43
cc_13 VNB Z 0.0497685f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.595
cc_14 VNB N_VGND_c_187_n 0.0209654f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.915
cc_15 VNB N_VGND_c_188_n 0.0317396f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.915
cc_16 VNB N_VGND_c_189_n 0.0186439f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.43
cc_17 VNB N_VGND_c_190_n 0.145051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_191_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.43
cc_19 VPB N_A_28_141#_c_36_n 0.0487039f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=0.915
cc_20 VPB N_TE_B_c_73_n 0.0292671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_21 VPB N_TE_B_M1001_g 0.0260994f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=0.915
cc_22 VPB N_TE_B_M1003_g 0.0220286f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=2.615
cc_23 VPB N_TE_B_c_76_n 0.0375161f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.43
cc_24 VPB TE_B 0.00177129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 VPB N_TE_B_c_72_n 0.0120584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_A_M1000_g 0.0438148f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=0.595
cc_27 VPB A 0.00281675f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=0.915
cc_28 VPB N_A_c_116_n 0.0199951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_152_n 0.0184055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_153_n 0.019457f $X=-0.19 $Y=1.655 $X2=0.265 $Y2=0.595
cc_31 VPB N_VPWR_c_154_n 0.0288092f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.43
cc_32 VPB N_VPWR_c_151_n 0.057094f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.43
cc_33 VPB N_VPWR_c_156_n 0.00641775f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.43
cc_34 VPB Z 0.0672407f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=0.595
cc_35 N_A_28_141#_c_35_n N_TE_B_M1004_g 0.0167815f $X=1.045 $Y=0.595 $X2=0 $Y2=0
cc_36 N_A_28_141#_c_36_n N_TE_B_M1004_g 0.0246734f $X=0.265 $Y=0.915 $X2=0 $Y2=0
cc_37 N_A_28_141#_c_37_n N_TE_B_M1004_g 9.58137e-19 $X=0.43 $Y=0.43 $X2=0 $Y2=0
cc_38 N_A_28_141#_c_38_n N_TE_B_M1004_g 0.00882631f $X=0.93 $Y=0.43 $X2=0 $Y2=0
cc_39 N_A_28_141#_c_39_n N_TE_B_M1004_g 0.00129679f $X=1.045 $Y=0.43 $X2=0 $Y2=0
cc_40 N_A_28_141#_c_36_n N_TE_B_c_73_n 0.0103255f $X=0.265 $Y=0.915 $X2=0 $Y2=0
cc_41 N_A_28_141#_c_36_n N_TE_B_M1001_g 0.00604718f $X=0.265 $Y=0.915 $X2=0
+ $Y2=0
cc_42 N_A_28_141#_c_36_n N_TE_B_c_76_n 0.00603347f $X=0.265 $Y=0.915 $X2=0 $Y2=0
cc_43 N_A_28_141#_c_35_n TE_B 4.13922e-19 $X=1.045 $Y=0.595 $X2=0 $Y2=0
cc_44 N_A_28_141#_c_36_n TE_B 0.0755304f $X=0.265 $Y=0.915 $X2=0 $Y2=0
cc_45 N_A_28_141#_c_36_n N_TE_B_c_72_n 0.00850854f $X=0.265 $Y=0.915 $X2=0 $Y2=0
cc_46 N_A_28_141#_c_39_n N_A_M1002_g 0.0359447f $X=1.045 $Y=0.43 $X2=0 $Y2=0
cc_47 N_A_28_141#_c_35_n A 0.00144136f $X=1.045 $Y=0.595 $X2=0 $Y2=0
cc_48 N_A_28_141#_c_36_n A 0.00457839f $X=0.265 $Y=0.915 $X2=0 $Y2=0
cc_49 N_A_28_141#_c_35_n N_A_c_116_n 2.76127e-19 $X=1.045 $Y=0.595 $X2=0 $Y2=0
cc_50 N_A_28_141#_c_36_n N_VPWR_c_152_n 0.00158275f $X=0.265 $Y=0.915 $X2=0
+ $Y2=0
cc_51 N_A_28_141#_c_36_n N_VPWR_c_153_n 0.00728859f $X=0.265 $Y=0.915 $X2=0
+ $Y2=0
cc_52 N_A_28_141#_c_36_n N_VPWR_c_151_n 0.01059f $X=0.265 $Y=0.915 $X2=0 $Y2=0
cc_53 N_A_28_141#_c_35_n N_VGND_c_192_n 0.0189365f $X=1.045 $Y=0.595 $X2=0 $Y2=0
cc_54 N_A_28_141#_c_38_n N_VGND_c_192_n 0.0273732f $X=0.93 $Y=0.43 $X2=0 $Y2=0
cc_55 N_A_28_141#_c_39_n N_VGND_c_192_n 0.00447359f $X=1.045 $Y=0.43 $X2=0 $Y2=0
cc_56 N_A_28_141#_c_38_n N_VGND_c_187_n 0.0250935f $X=0.93 $Y=0.43 $X2=0 $Y2=0
cc_57 N_A_28_141#_c_39_n N_VGND_c_187_n 0.0121828f $X=1.045 $Y=0.43 $X2=0 $Y2=0
cc_58 N_A_28_141#_c_37_n N_VGND_c_188_n 0.0222501f $X=0.43 $Y=0.43 $X2=0 $Y2=0
cc_59 N_A_28_141#_c_38_n N_VGND_c_188_n 0.0363486f $X=0.93 $Y=0.43 $X2=0 $Y2=0
cc_60 N_A_28_141#_c_39_n N_VGND_c_188_n 0.00953864f $X=1.045 $Y=0.43 $X2=0 $Y2=0
cc_61 N_A_28_141#_c_37_n N_VGND_c_190_n 0.0127687f $X=0.43 $Y=0.43 $X2=0 $Y2=0
cc_62 N_A_28_141#_c_38_n N_VGND_c_190_n 0.0220451f $X=0.93 $Y=0.43 $X2=0 $Y2=0
cc_63 N_A_28_141#_c_39_n N_VGND_c_190_n 0.0118956f $X=1.045 $Y=0.43 $X2=0 $Y2=0
cc_64 TE_B N_A_M1002_g 0.00101972f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_TE_B_c_73_n N_A_M1000_g 0.00474576f $X=0.64 $Y=2.065 $X2=0 $Y2=0
cc_66 N_TE_B_c_76_n N_A_M1000_g 0.0606473f $X=1.045 $Y=2.14 $X2=0 $Y2=0
cc_67 TE_B N_A_M1000_g 3.11508e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_68 N_TE_B_M1001_g A 6.46404e-19 $X=0.52 $Y=2.615 $X2=0 $Y2=0
cc_69 N_TE_B_M1003_g A 0.0169155f $X=1.045 $Y=2.725 $X2=0 $Y2=0
cc_70 N_TE_B_c_76_n A 0.00450006f $X=1.045 $Y=2.14 $X2=0 $Y2=0
cc_71 TE_B A 0.0621757f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_TE_B_c_72_n A 0.00391181f $X=0.71 $Y=1.71 $X2=0 $Y2=0
cc_73 N_TE_B_M1004_g N_A_c_116_n 6.83675e-19 $X=0.48 $Y=0.915 $X2=0 $Y2=0
cc_74 N_TE_B_c_76_n N_A_c_116_n 2.76127e-19 $X=1.045 $Y=2.14 $X2=0 $Y2=0
cc_75 TE_B N_A_c_116_n 5.58633e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_TE_B_c_72_n N_A_c_116_n 0.0153015f $X=0.71 $Y=1.71 $X2=0 $Y2=0
cc_77 N_TE_B_M1001_g N_VPWR_c_152_n 0.00461133f $X=0.52 $Y=2.615 $X2=0 $Y2=0
cc_78 N_TE_B_M1003_g N_VPWR_c_152_n 0.00667803f $X=1.045 $Y=2.725 $X2=0 $Y2=0
cc_79 N_TE_B_c_76_n N_VPWR_c_152_n 0.00173319f $X=1.045 $Y=2.14 $X2=0 $Y2=0
cc_80 TE_B N_VPWR_c_152_n 0.0243408f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_81 N_TE_B_M1001_g N_VPWR_c_153_n 0.00484506f $X=0.52 $Y=2.615 $X2=0 $Y2=0
cc_82 N_TE_B_M1003_g N_VPWR_c_154_n 0.0051803f $X=1.045 $Y=2.725 $X2=0 $Y2=0
cc_83 N_TE_B_M1001_g N_VPWR_c_151_n 0.00503886f $X=0.52 $Y=2.615 $X2=0 $Y2=0
cc_84 N_TE_B_M1003_g N_VPWR_c_151_n 0.0105874f $X=1.045 $Y=2.725 $X2=0 $Y2=0
cc_85 TE_B N_VGND_c_192_n 0.0229499f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_86 N_TE_B_c_72_n N_VGND_c_192_n 9.46865e-19 $X=0.71 $Y=1.71 $X2=0 $Y2=0
cc_87 N_TE_B_M1004_g N_VGND_c_188_n 4.76376e-19 $X=0.48 $Y=0.915 $X2=0 $Y2=0
cc_88 A N_VPWR_c_152_n 0.0222602f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A_M1000_g N_VPWR_c_154_n 0.0051803f $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_90 A N_VPWR_c_154_n 0.00906797f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A_M1000_g N_VPWR_c_151_n 0.0105147f $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_92 A N_VPWR_c_151_n 0.00973298f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_93 A A_224_481# 0.00150892f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_94 N_A_M1002_g Z 0.0337745f $X=1.435 $Y=0.915 $X2=0 $Y2=0
cc_95 A Z 0.112863f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A_M1002_g N_VGND_c_192_n 0.00525871f $X=1.435 $Y=0.915 $X2=0 $Y2=0
cc_97 A N_VGND_c_192_n 0.0181964f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_98 N_A_c_116_n N_VGND_c_192_n 8.1119e-19 $X=1.28 $Y=1.66 $X2=0 $Y2=0
cc_99 N_A_M1002_g N_VGND_c_187_n 0.0064653f $X=1.435 $Y=0.915 $X2=0 $Y2=0
cc_100 N_A_M1002_g N_VGND_c_189_n 0.00362253f $X=1.435 $Y=0.915 $X2=0 $Y2=0
cc_101 N_A_M1002_g N_VGND_c_190_n 0.00435931f $X=1.435 $Y=0.915 $X2=0 $Y2=0
cc_102 N_VPWR_c_152_n Z 3.00164e-19 $X=0.765 $Y=2.545 $X2=0 $Y2=0
cc_103 N_VPWR_c_154_n Z 0.0183256f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_104 N_VPWR_c_151_n Z 0.0110888f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_105 Z N_VGND_c_187_n 0.0036256f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_106 Z N_VGND_c_189_n 0.00527604f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_107 Z N_VGND_c_190_n 0.00842268f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_108 N_VGND_c_192_n A_224_141# 0.00153763f $X=1.195 $Y=0.907 $X2=-0.19
+ $Y2=-0.245
cc_109 N_VGND_c_187_n A_224_141# 7.62448e-19 $X=1.28 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
