* File: sky130_fd_sc_lp__or3_1.pex.spice
* Created: Fri Aug 28 11:23:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3_1%C 2 5 9 11 12 13 14 19
c40 5 0 1.40402e-19 $X=0.575 $Y=0.445
r41 19 21 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.005
+ $X2=0.605 $Y2=0.84
r42 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.005 $X2=0.59 $Y2=1.005
r43 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.67 $Y=1.295
+ $X2=0.67 $Y2=1.665
r44 13 20 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=0.67 $Y=1.295
+ $X2=0.67 $Y2=1.005
r45 12 20 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=0.67 $Y=0.925 $X2=0.67
+ $Y2=1.005
r46 9 11 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.71 $Y=2.52
+ $X2=0.71 $Y2=1.51
r47 5 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.575 $Y=0.445
+ $X2=0.575 $Y2=0.84
r48 2 11 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.605 $Y=1.33
+ $X2=0.605 $Y2=1.51
r49 1 19 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=0.605 $Y=1.02
+ $X2=0.605 $Y2=1.005
r50 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=0.605 $Y=1.02
+ $X2=0.605 $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_1%B 3 7 9 10 12 13 14 15 20
c48 13 0 1.40402e-19 $X=1.2 $Y=0.925
c49 12 0 3.36215e-20 $X=1.16 $Y=1.435
r50 15 29 9.0969 $w=3.08e-07 $l=2.4e-07 $layer=LI1_cond $X=1.175 $Y=1.665
+ $X2=1.175 $Y2=1.425
r51 14 29 5.44791 $w=2.73e-07 $l=1.3e-07 $layer=LI1_cond $X=1.157 $Y=1.295
+ $X2=1.157 $Y2=1.425
r52 13 14 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.157 $Y=0.925
+ $X2=1.157 $Y2=1.295
r53 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=0.93 $X2=1.16 $Y2=0.93
r54 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.16 $Y=1.27
+ $X2=1.16 $Y2=0.93
r55 11 12 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.27
+ $X2=1.16 $Y2=1.435
r56 10 20 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.16 $Y=0.915
+ $X2=1.16 $Y2=0.93
r57 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.212 $Y=0.765
+ $X2=1.212 $Y2=0.915
r58 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.355 $Y=0.445
+ $X2=1.355 $Y2=0.765
r59 3 12 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=1.15 $Y=2.52
+ $X2=1.15 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_1%A 3 7 9 12 13
c43 13 0 3.36215e-20 $X=1.73 $Y=1.51
r44 12 15 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.51
+ $X2=1.715 $Y2=1.675
r45 12 14 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.51
+ $X2=1.715 $Y2=1.345
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.51 $X2=1.73 $Y2=1.51
r47 9 13 4.52224 $w=3.93e-07 $l=1.55e-07 $layer=LI1_cond $X=1.697 $Y=1.665
+ $X2=1.697 $Y2=1.51
r48 7 14 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.785 $Y=0.445
+ $X2=1.785 $Y2=1.345
r49 3 15 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=1.61 $Y=2.52
+ $X2=1.61 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_1%A_47_47# 1 2 3 12 15 18 21 23 27 29 30 34 35
+ 39 41 43
r83 36 39 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=0.205 $Y=0.445
+ $X2=0.36 $Y2=0.445
r84 35 44 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.292 $Y=1.35
+ $X2=2.292 $Y2=1.515
r85 35 43 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.292 $Y=1.35
+ $X2=2.292 $Y2=1.185
r86 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.27
+ $Y=1.35 $X2=2.27 $Y2=1.35
r87 32 34 27.3705 $w=2.38e-07 $l=5.7e-07 $layer=LI1_cond $X=2.235 $Y=1.92
+ $X2=2.235 $Y2=1.35
r88 31 34 4.56175 $w=2.38e-07 $l=9.5e-08 $layer=LI1_cond $X=2.235 $Y=1.255
+ $X2=2.235 $Y2=1.35
r89 29 31 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.115 $Y=1.17
+ $X2=2.235 $Y2=1.255
r90 29 30 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.115 $Y=1.17
+ $X2=1.715 $Y2=1.17
r91 25 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.59 $Y=1.085
+ $X2=1.715 $Y2=1.17
r92 25 27 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=1.59 $Y=1.085
+ $X2=1.59 $Y2=0.445
r93 24 41 3.63156 $w=2.2e-07 $l=2.88e-07 $layer=LI1_cond $X=0.66 $Y=2.03
+ $X2=0.372 $Y2=2.03
r94 23 32 6.83327 $w=2.2e-07 $l=1.66132e-07 $layer=LI1_cond $X=2.115 $Y=2.03
+ $X2=2.235 $Y2=1.92
r95 23 24 76.2184 $w=2.18e-07 $l=1.455e-06 $layer=LI1_cond $X=2.115 $Y=2.03
+ $X2=0.66 $Y2=2.03
r96 19 41 3.01362 $w=4.07e-07 $l=1.1e-07 $layer=LI1_cond $X=0.372 $Y=2.14
+ $X2=0.372 $Y2=2.03
r97 19 21 7.90452 $w=5.73e-07 $l=3.8e-07 $layer=LI1_cond $X=0.372 $Y=2.14
+ $X2=0.372 $Y2=2.52
r98 18 41 3.01362 $w=4.07e-07 $l=2.15079e-07 $layer=LI1_cond $X=0.205 $Y=1.92
+ $X2=0.372 $Y2=2.03
r99 17 36 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.205 $Y=0.61
+ $X2=0.205 $Y2=0.445
r100 17 18 62.9042 $w=2.38e-07 $l=1.31e-06 $layer=LI1_cond $X=0.205 $Y=0.61
+ $X2=0.205 $Y2=1.92
r101 15 44 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.405 $Y=2.465
+ $X2=2.405 $Y2=1.515
r102 12 43 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.33 $Y=0.655
+ $X2=2.33 $Y2=1.185
r103 3 21 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.37
+ $Y=2.31 $X2=0.495 $Y2=2.52
r104 2 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.445
r105 1 39 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.235 $X2=0.36 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_1%VPWR 1 6 10 12 19 20 23
r25 24 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 23 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 20 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 17 23 13.6095 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.007 $Y2=3.33
r31 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 12 23 13.6095 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=1.66 $Y=3.33
+ $X2=2.007 $Y2=3.33
r34 12 14 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=1.66 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 10 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 10 15 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 6 9 9.12117 $w=6.93e-07 $l=5.3e-07 $layer=LI1_cond $X=2.007 $Y=2.42
+ $X2=2.007 $Y2=2.95
r38 4 23 2.84707 $w=6.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.007 $Y=3.245
+ $X2=2.007 $Y2=3.33
r39 4 9 5.07688 $w=6.93e-07 $l=2.95e-07 $layer=LI1_cond $X=2.007 $Y=3.245
+ $X2=2.007 $Y2=2.95
r40 1 9 600 $w=1.7e-07 $l=8.56037e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=2.31 $X2=2.19 $Y2=2.95
r41 1 6 300 $w=1.7e-07 $l=5.57293e-07 $layer=licon1_PDIFF $count=2 $X=1.685
+ $Y=2.31 $X2=2.19 $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_1%X 1 2 7 8 9 10 11 12 13 24 30
r17 30 47 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=2.655 $Y=0.925
+ $X2=2.655 $Y2=0.905
r18 13 44 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=2.655 $Y=2.775
+ $X2=2.655 $Y2=2.91
r19 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.655 $Y=2.405
+ $X2=2.655 $Y2=2.775
r20 11 12 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=2.655 $Y=1.98
+ $X2=2.655 $Y2=2.405
r21 10 11 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.655 $Y=1.665
+ $X2=2.655 $Y2=1.98
r22 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.655 $Y=1.295
+ $X2=2.655 $Y2=1.665
r23 8 47 2.41196 $w=4.03e-07 $l=3.3e-08 $layer=LI1_cond $X=2.582 $Y=0.872
+ $X2=2.582 $Y2=0.905
r24 8 22 4.80896 $w=4.03e-07 $l=1.69e-07 $layer=LI1_cond $X=2.582 $Y=0.872
+ $X2=2.582 $Y2=0.703
r25 8 9 14.9818 $w=2.58e-07 $l=3.38e-07 $layer=LI1_cond $X=2.655 $Y=0.957
+ $X2=2.655 $Y2=1.295
r26 8 30 1.41839 $w=2.58e-07 $l=3.2e-08 $layer=LI1_cond $X=2.655 $Y=0.957
+ $X2=2.655 $Y2=0.925
r27 7 22 4.2114 $w=4.03e-07 $l=1.48e-07 $layer=LI1_cond $X=2.582 $Y=0.555
+ $X2=2.582 $Y2=0.703
r28 7 24 3.84148 $w=4.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.582 $Y=0.555
+ $X2=2.582 $Y2=0.42
r29 2 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2.91
r30 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=1.98
r31 1 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.405
+ $Y=0.235 $X2=2.545 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_1%VGND 1 2 11 14 15 16 23 24 27 35
r39 33 35 9.44511 $w=6.78e-07 $l=9.5e-08 $layer=LI1_cond $X=1.2 $Y=0.255
+ $X2=1.295 $Y2=0.255
r40 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 31 33 1.05536 $w=6.78e-07 $l=6e-08 $layer=LI1_cond $X=1.14 $Y=0.255 $X2=1.2
+ $Y2=0.255
r42 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r43 27 31 7.38754 $w=6.78e-07 $l=4.2e-07 $layer=LI1_cond $X=0.72 $Y=0.255
+ $X2=1.14 $Y2=0.255
r44 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 21 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r47 20 35 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.295
+ $Y2=0
r48 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r49 16 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r50 16 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r51 14 20 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=1.68
+ $Y2=0
r52 14 15 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=2.047
+ $Y2=0
r53 13 23 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.64
+ $Y2=0
r54 13 15 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.047
+ $Y2=0
r55 9 15 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.047 $Y=0.085
+ $X2=2.047 $Y2=0
r56 9 11 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=2.047 $Y=0.085
+ $X2=2.047 $Y2=0.38
r57 2 11 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=1.86
+ $Y=0.235 $X2=2.05 $Y2=0.38
r58 1 31 91 $w=1.7e-07 $l=5.79353e-07 $layer=licon1_NDIFF $count=2 $X=0.65
+ $Y=0.235 $X2=1.14 $Y2=0.43
.ends

