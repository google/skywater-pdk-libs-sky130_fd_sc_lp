# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__sdfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.24000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 0.810000 1.795000 1.795000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.365000 0.265000 17.695000 3.065000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.410000 0.265000 15.765000 1.125000 ;
        RECT 15.485000 1.815000 15.765000 3.065000 ;
        RECT 15.595000 1.125000 15.765000 1.815000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.525000 1.345000 14.920000 1.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.215000 0.550000 1.885000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895000 1.215000 1.315000 1.885000 ;
    END
  END SCE
  PIN SET_B
    ANTENNADIFFAREA  2.773000 ;
    ANTENNAPARTIALMETALSIDEAREA  3.451000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.605000 1.180000 12.950000 1.780000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.870000 1.110000 4.200000 1.780000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 18.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 18.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.240000 0.085000 ;
      RECT  0.000000  3.245000 18.240000 3.415000 ;
      RECT  0.165000  0.085000  0.495000 1.035000 ;
      RECT  0.260000  2.065000  1.470000 2.235000 ;
      RECT  0.260000  2.235000  0.590000 3.065000 ;
      RECT  0.770000  2.415000  1.100000 3.245000 ;
      RECT  0.985000  0.460000  2.145000 0.630000 ;
      RECT  0.985000  0.630000  1.315000 1.035000 ;
      RECT  1.300000  2.235000  1.470000 2.895000 ;
      RECT  1.300000  2.895000  2.490000 3.065000 ;
      RECT  1.650000  2.035000  4.245000 2.205000 ;
      RECT  1.650000  2.205000  1.980000 2.715000 ;
      RECT  1.975000  0.630000  2.145000 2.035000 ;
      RECT  2.160000  2.385000  2.490000 2.895000 ;
      RECT  2.325000  0.085000  2.655000 1.005000 ;
      RECT  2.325000  1.185000  2.580000 1.515000 ;
      RECT  2.325000  1.515000  3.445000 1.855000 ;
      RECT  2.720000  2.425000  3.050000 3.245000 ;
      RECT  2.945000  0.575000  3.445000 1.515000 ;
      RECT  3.645000  2.385000  3.895000 3.245000 ;
      RECT  3.665000  0.085000  3.995000 0.915000 ;
      RECT  4.075000  2.205000  4.245000 2.895000 ;
      RECT  4.075000  2.895000  5.180000 3.065000 ;
      RECT  4.175000  0.455000  4.595000 0.915000 ;
      RECT  4.425000  0.915000  4.595000 1.005000 ;
      RECT  4.425000  1.005000  4.770000 2.715000 ;
      RECT  4.870000  0.315000  5.200000 0.775000 ;
      RECT  4.950000  0.775000  5.200000 1.815000 ;
      RECT  4.950000  1.815000  5.890000 1.985000 ;
      RECT  4.950000  1.985000  5.200000 2.145000 ;
      RECT  5.010000  2.325000  6.240000 2.495000 ;
      RECT  5.010000  2.495000  5.180000 2.895000 ;
      RECT  5.360000  2.675000  5.690000 3.245000 ;
      RECT  5.380000  0.085000  5.710000 0.775000 ;
      RECT  5.615000  1.315000  5.890000 1.815000 ;
      RECT  5.910000  0.665000  6.240000 1.125000 ;
      RECT  5.910000  2.295000  6.240000 2.325000 ;
      RECT  5.910000  2.495000  6.240000 2.755000 ;
      RECT  6.070000  1.125000  6.240000 2.295000 ;
      RECT  6.420000  0.665000  6.590000 2.075000 ;
      RECT  6.420000  2.075000  7.295000 2.245000 ;
      RECT  6.420000  2.245000  6.750000 2.755000 ;
      RECT  6.770000  0.830000  8.145000 1.000000 ;
      RECT  6.770000  1.000000  6.945000 1.545000 ;
      RECT  7.125000  1.475000  8.005000 1.645000 ;
      RECT  7.125000  1.645000  7.295000 2.075000 ;
      RECT  7.465000  0.085000  7.795000 0.650000 ;
      RECT  7.475000  1.825000  7.655000 2.075000 ;
      RECT  7.475000  2.075000  9.330000 2.245000 ;
      RECT  7.835000  1.645000  8.005000 1.725000 ;
      RECT  7.835000  1.725000  8.980000 1.895000 ;
      RECT  7.955000  2.425000  8.285000 3.245000 ;
      RECT  7.975000  0.265000 10.025000 0.435000 ;
      RECT  7.975000  0.435000  8.145000 0.830000 ;
      RECT  8.185000  1.180000  8.515000 1.545000 ;
      RECT  8.325000  0.615000  9.675000 0.785000 ;
      RECT  8.325000  0.785000  8.655000 1.000000 ;
      RECT  8.525000  2.245000  9.330000 2.755000 ;
      RECT  8.705000  1.405000  8.980000 1.725000 ;
      RECT  8.835000  0.965000  9.165000 1.055000 ;
      RECT  8.835000  1.055000  9.330000 1.225000 ;
      RECT  9.160000  1.225000  9.330000 1.445000 ;
      RECT  9.160000  1.445000 10.500000 1.615000 ;
      RECT  9.160000  1.615000  9.330000 2.075000 ;
      RECT  9.345000  0.785000  9.675000 0.875000 ;
      RECT  9.510000  1.875000  9.840000 3.245000 ;
      RECT  9.855000  0.435000 10.025000 1.095000 ;
      RECT  9.855000  1.095000 11.120000 1.265000 ;
      RECT 10.170000  1.615000 10.500000 1.705000 ;
      RECT 10.205000  0.085000 10.455000 0.915000 ;
      RECT 10.680000  1.265000 11.120000 1.675000 ;
      RECT 10.680000  1.675000 10.850000 2.895000 ;
      RECT 10.680000  2.895000 12.020000 3.065000 ;
      RECT 11.030000  2.120000 11.470000 2.715000 ;
      RECT 11.300000  0.575000 11.630000 0.830000 ;
      RECT 11.300000  0.830000 13.300000 1.000000 ;
      RECT 11.300000  1.000000 11.630000 1.255000 ;
      RECT 11.300000  1.255000 11.470000 2.120000 ;
      RECT 11.690000  1.700000 12.020000 2.895000 ;
      RECT 12.230000  1.960000 12.560000 2.120000 ;
      RECT 12.230000  2.120000 13.445000 2.290000 ;
      RECT 12.335000  0.085000 12.665000 0.650000 ;
      RECT 12.685000  2.470000 12.935000 3.245000 ;
      RECT 12.925000  0.265000 14.240000 0.435000 ;
      RECT 12.925000  0.435000 13.255000 0.650000 ;
      RECT 13.115000  2.290000 13.445000 2.390000 ;
      RECT 13.115000  2.390000 15.305000 2.560000 ;
      RECT 13.115000  2.560000 13.445000 3.065000 ;
      RECT 13.130000  1.000000 13.300000 1.460000 ;
      RECT 13.130000  1.460000 13.485000 1.790000 ;
      RECT 13.480000  0.615000 13.810000 0.995000 ;
      RECT 13.480000  0.995000 13.835000 1.165000 ;
      RECT 13.665000  1.165000 13.835000 2.390000 ;
      RECT 13.935000  2.740000 14.265000 3.245000 ;
      RECT 13.990000  0.435000 14.240000 0.815000 ;
      RECT 14.015000  0.995000 14.800000 1.165000 ;
      RECT 14.015000  1.165000 14.340000 1.960000 ;
      RECT 14.015000  1.960000 14.795000 2.210000 ;
      RECT 14.470000  0.665000 14.800000 0.995000 ;
      RECT 14.975000  2.740000 15.305000 3.245000 ;
      RECT 14.980000  0.085000 15.230000 1.125000 ;
      RECT 15.135000  1.305000 15.415000 1.635000 ;
      RECT 15.135000  1.635000 15.305000 2.390000 ;
      RECT 15.945000  0.085000 16.195000 1.125000 ;
      RECT 15.945000  1.815000 16.195000 3.245000 ;
      RECT 16.425000  0.295000 16.755000 1.185000 ;
      RECT 16.425000  1.185000 17.185000 1.515000 ;
      RECT 16.425000  1.515000 16.755000 2.640000 ;
      RECT 16.935000  0.085000 17.185000 1.005000 ;
      RECT 16.935000  1.815000 17.185000 3.245000 ;
      RECT 17.875000  0.085000 18.125000 1.095000 ;
      RECT 17.875000  1.815000 18.125000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.210000  8.485000 1.380000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  1.210000 12.805000 1.380000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.245000 18.085000 3.415000 ;
    LAYER met1 ;
      RECT  8.255000 1.180000  8.545000 1.225000 ;
      RECT  8.255000 1.225000 12.865000 1.365000 ;
      RECT  8.255000 1.365000  8.545000 1.410000 ;
      RECT 12.575000 1.180000 12.865000 1.225000 ;
      RECT 12.575000 1.365000 12.865000 1.410000 ;
  END
END sky130_fd_sc_lp__sdfbbn_2
