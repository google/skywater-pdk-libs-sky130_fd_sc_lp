* File: sky130_fd_sc_lp__dlrbn_2.spice
* Created: Wed Sep  2 09:46:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrbn_2.pex.spice"
.subckt sky130_fd_sc_lp__dlrbn_2  VNB VPB GATE_N D RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* GATE_N	GATE_N
* VPB	VPB
* VNB	VNB
MM1007 N_A_113_144#_M1007_d N_GATE_N_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_113_144#_M1016_g N_A_162_40#_M1016_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_392_144#_M1017_d N_D_M1017_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1025 N_A_591_155#_M1025_d N_A_113_144#_M1025_g N_A_508_155#_M1025_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_A_677_155#_M1019_d N_A_162_40#_M1019_g N_A_591_155#_M1025_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1449 AS=0.0588 PD=1.53 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_392_144#_M1014_g N_A_508_155#_M1014_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_677_155#_M1004_d N_A_942_252#_M1004_g N_VGND_M1014_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 A_1184_60# N_A_591_155#_M1027_g N_A_942_252#_M1027_s VNB NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_RESET_B_M1002_g A_1184_60# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.0882 PD=1.23 PS=1.05 NRD=5.712 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1009 N_Q_M1009_d N_A_942_252#_M1009_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1638 PD=1.12 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.1
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1022 N_Q_M1009_d N_A_942_252#_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1834 PD=1.12 PS=1.64 NRD=0 NRS=7.848 M=1 R=5.6 SA=75001.5
+ SB=75000.5 A=0.126 P=1.98 MULT=1
MM1011 N_A_1555_367#_M1011_d N_A_942_252#_M1011_g N_VGND_M1022_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0917 PD=1.37 PS=0.82 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_1555_367#_M1003_g N_Q_N_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_1555_367#_M1013_g N_Q_N_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1026 N_A_113_144#_M1026_d N_GATE_N_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_A_113_144#_M1012_g N_A_162_40#_M1012_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1392 AS=0.1696 PD=1.075 PS=1.81 NRD=19.9955 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1008 N_A_392_144#_M1008_d N_D_M1008_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1392 PD=1.81 PS=1.075 NRD=0 NRS=27.6982 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_A_591_155#_M1024_d N_A_113_144#_M1024_g N_A_606_359#_M1024_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0855057 AS=0.1113 PD=0.80434 PS=1.37 NRD=46.886
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1015 A_794_359# N_A_162_40#_M1015_g N_A_591_155#_M1024_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0672 AS=0.130294 PD=0.85 PS=1.22566 NRD=15.3857 NRS=0 M=1
+ R=4.26667 SA=75000.5 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1018 N_VPWR_M1018_d N_A_392_144#_M1018_g A_794_359# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.132226 AS=0.0672 PD=1.2317 PS=0.85 NRD=1.5366 NRS=15.3857 M=1 R=4.26667
+ SA=75000.9 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1005 N_A_606_359#_M1005_d N_A_942_252#_M1005_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0867736 PD=1.37 PS=0.808302 NRD=0 NRS=71.0973 M=1
+ R=2.8 SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_A_942_252#_M1020_d N_A_591_155#_M1020_g N_VPWR_M1020_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.8 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_RESET_B_M1006_g N_A_942_252#_M1020_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.4 A=0.189 P=2.82 MULT=1
MM1000 N_Q_M1000_d N_A_942_252#_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75001.1
+ SB=75000.9 A=0.189 P=2.82 MULT=1
MM1021 N_Q_M1000_d N_A_942_252#_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.268115 PD=1.54 PS=2.16853 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.5 A=0.189 P=2.82 MULT=1
MM1010 N_A_1555_367#_M1010_d N_A_942_252#_M1010_g N_VPWR_M1021_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.136185 PD=1.81 PS=1.10147 NRD=0 NRS=48.5605 M=1
+ R=4.26667 SA=75002 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_Q_N_M1001_d N_A_1555_367#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1023 N_Q_N_M1001_d N_A_1555_367#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=18.7859 P=23.77
*
.include "sky130_fd_sc_lp__dlrbn_2.pxi.spice"
*
.ends
*
*
