# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xor2_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__xor2_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.295000 1.900000 1.690000 ;
        RECT 1.085000 1.690000 3.265000 1.860000 ;
        RECT 2.935000 1.180000 3.265000 1.690000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.290000 1.180000 2.755000 1.510000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.417600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.215000 0.905000 1.385000 ;
        RECT 0.125000 1.385000 0.355000 2.075000 ;
        RECT 0.125000 2.075000 0.555000 3.065000 ;
        RECT 0.735000 0.575000 1.235000 1.035000 ;
        RECT 0.735000 1.035000 0.905000 1.215000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.035000 ;
      RECT 0.535000  1.565000 0.905000 1.895000 ;
      RECT 0.735000  1.895000 0.905000 2.040000 ;
      RECT 0.735000  2.040000 3.615000 2.210000 ;
      RECT 0.770000  2.390000 2.160000 2.560000 ;
      RECT 0.770000  2.560000 1.100000 3.065000 ;
      RECT 1.300000  2.740000 1.630000 3.245000 ;
      RECT 1.775000  0.085000 2.105000 0.780000 ;
      RECT 1.830000  2.560000 2.160000 3.065000 ;
      RECT 2.395000  2.210000 2.725000 3.065000 ;
      RECT 2.595000  0.320000 2.925000 0.830000 ;
      RECT 2.595000  0.830000 3.615000 1.000000 ;
      RECT 3.385000  0.085000 3.715000 0.650000 ;
      RECT 3.385000  2.390000 3.715000 3.245000 ;
      RECT 3.445000  1.000000 3.615000 2.040000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__xor2_lp
