* File: sky130_fd_sc_lp__o22ai_2.pxi.spice
* Created: Fri Aug 28 11:10:51 2020
* 
x_PM_SKY130_FD_SC_LP__O22AI_2%B1 N_B1_c_76_n N_B1_M1012_g N_B1_M1006_g
+ N_B1_c_78_n N_B1_M1013_g N_B1_M1011_g N_B1_c_87_p B1 N_B1_c_81_n
+ PM_SKY130_FD_SC_LP__O22AI_2%B1
x_PM_SKY130_FD_SC_LP__O22AI_2%B2 N_B2_M1000_g N_B2_c_118_n N_B2_M1002_g
+ N_B2_M1009_g N_B2_c_120_n N_B2_M1007_g B2 B2 N_B2_c_122_n
+ PM_SKY130_FD_SC_LP__O22AI_2%B2
x_PM_SKY130_FD_SC_LP__O22AI_2%A2 N_A2_c_168_n N_A2_M1004_g N_A2_M1001_g
+ N_A2_c_170_n N_A2_M1015_g N_A2_M1010_g A2 A2 A2 N_A2_c_173_n
+ PM_SKY130_FD_SC_LP__O22AI_2%A2
x_PM_SKY130_FD_SC_LP__O22AI_2%A1 N_A1_c_222_n N_A1_M1003_g N_A1_M1005_g
+ N_A1_c_224_n N_A1_M1008_g N_A1_M1014_g A1 A1 N_A1_c_227_n
+ PM_SKY130_FD_SC_LP__O22AI_2%A1
x_PM_SKY130_FD_SC_LP__O22AI_2%A_43_367# N_A_43_367#_M1006_s N_A_43_367#_M1011_s
+ N_A_43_367#_M1009_d N_A_43_367#_c_262_n N_A_43_367#_c_263_n
+ N_A_43_367#_c_264_n N_A_43_367#_c_279_p N_A_43_367#_c_275_n
+ N_A_43_367#_c_265_n N_A_43_367#_c_266_n PM_SKY130_FD_SC_LP__O22AI_2%A_43_367#
x_PM_SKY130_FD_SC_LP__O22AI_2%VPWR N_VPWR_M1006_d N_VPWR_M1005_s N_VPWR_c_300_n
+ N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n VPWR N_VPWR_c_304_n
+ N_VPWR_c_305_n N_VPWR_c_299_n N_VPWR_c_307_n PM_SKY130_FD_SC_LP__O22AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O22AI_2%Y N_Y_M1012_d N_Y_M1002_d N_Y_M1000_s N_Y_M1001_s
+ N_Y_c_365_n N_Y_c_375_n N_Y_c_360_n N_Y_c_361_n N_Y_c_362_n N_Y_c_393_n
+ N_Y_c_358_n Y Y Y N_Y_c_388_n Y PM_SKY130_FD_SC_LP__O22AI_2%Y
x_PM_SKY130_FD_SC_LP__O22AI_2%A_491_367# N_A_491_367#_M1001_d
+ N_A_491_367#_M1010_d N_A_491_367#_M1014_d N_A_491_367#_c_425_n
+ N_A_491_367#_c_426_n N_A_491_367#_c_430_n N_A_491_367#_c_448_n
+ N_A_491_367#_c_427_n N_A_491_367#_c_428_n N_A_491_367#_c_429_n
+ PM_SKY130_FD_SC_LP__O22AI_2%A_491_367#
x_PM_SKY130_FD_SC_LP__O22AI_2%A_43_65# N_A_43_65#_M1012_s N_A_43_65#_M1013_s
+ N_A_43_65#_M1007_s N_A_43_65#_M1015_s N_A_43_65#_M1008_s N_A_43_65#_c_460_n
+ N_A_43_65#_c_461_n N_A_43_65#_c_462_n N_A_43_65#_c_463_n N_A_43_65#_c_464_n
+ N_A_43_65#_c_475_n N_A_43_65#_c_479_n N_A_43_65#_c_465_n N_A_43_65#_c_484_n
+ N_A_43_65#_c_466_n N_A_43_65#_c_467_n N_A_43_65#_c_468_n N_A_43_65#_c_485_n
+ PM_SKY130_FD_SC_LP__O22AI_2%A_43_65#
x_PM_SKY130_FD_SC_LP__O22AI_2%VGND N_VGND_M1004_d N_VGND_M1003_d N_VGND_c_525_n
+ N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n N_VGND_c_530_n
+ VGND N_VGND_c_531_n N_VGND_c_532_n PM_SKY130_FD_SC_LP__O22AI_2%VGND
cc_1 VNB N_B1_c_76_n 0.0200925f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.275
cc_2 VNB N_B1_M1006_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_3 VNB N_B1_c_78_n 0.0170222f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.275
cc_4 VNB N_B1_M1011_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_5 VNB B1 0.021329f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_B1_c_81_n 0.0698987f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.44
cc_7 VNB N_B2_M1000_g 0.00257351f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.745
cc_8 VNB N_B2_c_118_n 0.0165307f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_9 VNB N_B2_M1009_g 0.00268533f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.745
cc_10 VNB N_B2_c_120_n 0.0187359f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_11 VNB B2 0.012451f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.48
cc_12 VNB N_B2_c_122_n 0.0457274f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.44
cc_13 VNB N_A2_c_168_n 0.0184279f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.275
cc_14 VNB N_A2_M1001_g 0.00298541f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_15 VNB N_A2_c_170_n 0.0160333f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.275
cc_16 VNB N_A2_M1010_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_17 VNB A2 0.0155099f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.44
cc_18 VNB N_A2_c_173_n 0.0536929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_222_n 0.0160333f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.275
cc_20 VNB N_A1_M1005_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_21 VNB N_A1_c_224_n 0.021262f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.275
cc_22 VNB N_A1_M1014_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_23 VNB A1 0.0419807f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.48
cc_24 VNB N_A1_c_227_n 0.0561609f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.44
cc_25 VNB N_VPWR_c_299_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_358_n 0.00228105f $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=1.295
cc_27 VNB Y 0.011422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_43_65#_c_460_n 0.0233564f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.44
cc_29 VNB N_A_43_65#_c_461_n 0.00928796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_43_65#_c_462_n 0.00655396f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.44
cc_31 VNB N_A_43_65#_c_463_n 0.00142321f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.44
cc_32 VNB N_A_43_65#_c_464_n 0.0021606f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.44
cc_33 VNB N_A_43_65#_c_465_n 0.00160609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_43_65#_c_466_n 0.0075508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_43_65#_c_467_n 0.0230663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_43_65#_c_468_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_525_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.745
cc_38 VNB N_VGND_c_526_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_39 VNB N_VGND_c_527_n 0.0666147f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.48
cc_40 VNB N_VGND_c_528_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.44
cc_41 VNB N_VGND_c_529_n 0.0144043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_530_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_43 VNB N_VGND_c_531_n 0.0261019f $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=1.48
cc_44 VNB N_VGND_c_532_n 0.288166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_B1_M1006_g 0.0262031f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_46 VPB N_B1_M1011_g 0.0193377f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_47 VPB N_B2_M1000_g 0.0195515f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.745
cc_48 VPB N_B2_M1009_g 0.0235138f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=0.745
cc_49 VPB N_A2_M1001_g 0.0237588f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_50 VPB N_A2_M1010_g 0.0195248f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_51 VPB N_A1_M1005_g 0.0185451f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_52 VPB N_A1_M1014_g 0.0243928f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_53 VPB N_A_43_367#_c_262_n 0.0427769f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_54 VPB N_A_43_367#_c_263_n 0.00653738f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.48
cc_55 VPB N_A_43_367#_c_264_n 0.00890498f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.44
cc_56 VPB N_A_43_367#_c_265_n 0.00181169f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.44
cc_57 VPB N_A_43_367#_c_266_n 0.00809879f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.44
cc_58 VPB N_VPWR_c_300_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.985 $Y2=0.745
cc_59 VPB N_VPWR_c_301_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.48
cc_60 VPB N_VPWR_c_302_n 0.0643861f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_61 VPB N_VPWR_c_303_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_304_n 0.0179216f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.44
cc_63 VPB N_VPWR_c_305_n 0.0230131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_299_n 0.0670253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_307_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_Y_c_360_n 7.46496e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_Y_c_361_n 0.00228659f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.44
cc_68 VPB N_Y_c_362_n 0.0178584f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.44
cc_69 VPB Y 0.00110672f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB Y 0.00246761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_491_367#_c_425_n 0.00181169f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=0.745
cc_72 VPB N_A_491_367#_c_426_n 0.00809951f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_73 VPB N_A_491_367#_c_427_n 0.0134556f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_74 VPB N_A_491_367#_c_428_n 0.00274866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_491_367#_c_429_n 0.0457879f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.44
cc_76 N_B1_M1011_g N_B2_M1000_g 0.0190801f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_77 N_B1_c_78_n N_B2_c_118_n 0.0302608f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_78 N_B1_c_78_n B2 0.00434752f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_79 N_B1_c_87_p B2 0.0146507f $X=0.77 $Y=1.44 $X2=0 $Y2=0
cc_80 B1 B2 0.00445101f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_B1_c_87_p N_B2_c_122_n 5.71605e-19 $X=0.77 $Y=1.44 $X2=0 $Y2=0
cc_82 N_B1_c_81_n N_B2_c_122_n 0.0190801f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_83 N_B1_M1006_g N_A_43_367#_c_263_n 0.0134039f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_84 N_B1_M1011_g N_A_43_367#_c_263_n 0.0166202f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_85 N_B1_c_87_p N_A_43_367#_c_263_n 0.0361069f $X=0.77 $Y=1.44 $X2=0 $Y2=0
cc_86 N_B1_c_81_n N_A_43_367#_c_263_n 0.00324879f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_87 B1 N_A_43_367#_c_264_n 0.0222213f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B1_c_81_n N_A_43_367#_c_264_n 0.00204992f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_89 N_B1_M1006_g N_VPWR_c_300_n 0.0159861f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_90 N_B1_M1011_g N_VPWR_c_300_n 0.0151897f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B1_M1011_g N_VPWR_c_302_n 0.00486043f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_92 N_B1_M1006_g N_VPWR_c_304_n 0.00486043f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_93 N_B1_M1006_g N_VPWR_c_299_n 0.00924722f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_94 N_B1_M1011_g N_VPWR_c_299_n 0.0082726f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_95 N_B1_c_78_n N_Y_c_365_n 0.0149928f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_96 N_B1_M1011_g N_Y_c_361_n 4.40373e-19 $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_97 N_B1_c_76_n N_Y_c_358_n 0.0119257f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_98 N_B1_c_78_n N_Y_c_358_n 0.00891785f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_99 N_B1_c_87_p N_Y_c_358_n 0.0266134f $X=0.77 $Y=1.44 $X2=0 $Y2=0
cc_100 N_B1_c_81_n N_Y_c_358_n 0.00255166f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_101 B1 N_A_43_65#_c_460_n 0.0223423f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B1_c_81_n N_A_43_65#_c_460_n 0.00169228f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_103 N_B1_c_76_n N_A_43_65#_c_468_n 0.0125492f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_104 N_B1_c_78_n N_A_43_65#_c_468_n 0.00930819f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_105 N_B1_c_76_n N_VGND_c_527_n 0.00302501f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_106 N_B1_c_78_n N_VGND_c_527_n 0.00302501f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_107 N_B1_c_76_n N_VGND_c_532_n 0.00473131f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_108 N_B1_c_78_n N_VGND_c_532_n 0.00441692f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_109 N_B2_c_120_n N_A2_c_168_n 0.00597485f $X=1.925 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_110 N_B2_c_122_n N_A2_c_173_n 0.00478178f $X=1.845 $Y=1.44 $X2=0 $Y2=0
cc_111 N_B2_M1000_g N_A_43_367#_c_263_n 4.89726e-19 $X=1.415 $Y=2.465 $X2=0
+ $Y2=0
cc_112 B2 N_A_43_367#_c_263_n 0.0127872f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B2_M1000_g N_A_43_367#_c_275_n 0.0115031f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_114 N_B2_M1009_g N_A_43_367#_c_275_n 0.0114565f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_115 N_B2_M1000_g N_VPWR_c_300_n 0.00109252f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B2_M1000_g N_VPWR_c_302_n 0.00357877f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B2_M1009_g N_VPWR_c_302_n 0.00357877f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_118 N_B2_M1000_g N_VPWR_c_299_n 0.00537654f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B2_M1009_g N_VPWR_c_299_n 0.00665089f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B2_c_118_n N_Y_c_365_n 0.0100464f $X=1.495 $Y=1.275 $X2=0 $Y2=0
cc_121 N_B2_c_120_n N_Y_c_365_n 0.0088432f $X=1.925 $Y=1.275 $X2=0 $Y2=0
cc_122 B2 N_Y_c_365_n 0.0479557f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_123 N_B2_c_122_n N_Y_c_365_n 9.45861e-19 $X=1.845 $Y=1.44 $X2=0 $Y2=0
cc_124 N_B2_M1000_g N_Y_c_375_n 0.0122296f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B2_M1009_g N_Y_c_375_n 0.0182396f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B2_M1009_g N_Y_c_360_n 0.0145067f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_127 B2 N_Y_c_360_n 0.00245623f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_128 N_B2_c_122_n N_Y_c_360_n 0.00220446f $X=1.845 $Y=1.44 $X2=0 $Y2=0
cc_129 N_B2_M1000_g N_Y_c_361_n 0.00452114f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_130 N_B2_M1009_g N_Y_c_361_n 0.00241999f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_131 B2 N_Y_c_361_n 0.0275189f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B2_c_122_n N_Y_c_361_n 0.00291181f $X=1.845 $Y=1.44 $X2=0 $Y2=0
cc_133 N_B2_c_118_n N_Y_c_358_n 0.00167699f $X=1.495 $Y=1.275 $X2=0 $Y2=0
cc_134 N_B2_c_120_n Y 0.00574783f $X=1.925 $Y=1.275 $X2=0 $Y2=0
cc_135 B2 Y 0.0260488f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B2_c_122_n Y 0.0074042f $X=1.845 $Y=1.44 $X2=0 $Y2=0
cc_137 N_B2_c_120_n N_Y_c_388_n 0.00325608f $X=1.925 $Y=1.275 $X2=0 $Y2=0
cc_138 N_B2_c_118_n N_A_43_65#_c_462_n 0.0184982f $X=1.495 $Y=1.275 $X2=0 $Y2=0
cc_139 N_B2_c_120_n N_A_43_65#_c_462_n 0.0147318f $X=1.925 $Y=1.275 $X2=0 $Y2=0
cc_140 N_B2_c_120_n N_A_43_65#_c_475_n 0.00325243f $X=1.925 $Y=1.275 $X2=0 $Y2=0
cc_141 N_B2_c_118_n N_VGND_c_527_n 0.00302501f $X=1.495 $Y=1.275 $X2=0 $Y2=0
cc_142 N_B2_c_120_n N_VGND_c_527_n 0.00302501f $X=1.925 $Y=1.275 $X2=0 $Y2=0
cc_143 N_B2_c_118_n N_VGND_c_532_n 0.00442601f $X=1.495 $Y=1.275 $X2=0 $Y2=0
cc_144 N_B2_c_120_n N_VGND_c_532_n 0.004608f $X=1.925 $Y=1.275 $X2=0 $Y2=0
cc_145 N_A2_c_170_n N_A1_c_222_n 0.0145992f $X=3.155 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_146 A2 N_A1_c_222_n 0.00413598f $X=3.515 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_147 N_A2_M1010_g N_A1_M1005_g 0.0158117f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_148 A2 N_A1_c_224_n 2.56035e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_149 A2 A1 0.0267416f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_150 A2 N_A1_c_227_n 0.0157165f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_151 N_A2_c_173_n N_A1_c_227_n 0.0256231f $X=3.225 $Y=1.44 $X2=0 $Y2=0
cc_152 N_A2_M1010_g N_VPWR_c_301_n 0.00109252f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A2_M1001_g N_VPWR_c_302_n 0.00357877f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A2_M1010_g N_VPWR_c_302_n 0.00357877f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A2_M1001_g N_VPWR_c_299_n 0.00665089f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A2_M1010_g N_VPWR_c_299_n 0.00537654f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A2_M1001_g N_Y_c_362_n 0.0156105f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A2_M1010_g N_Y_c_362_n 0.00374173f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_159 A2 N_Y_c_362_n 0.0569666f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A2_c_173_n N_Y_c_362_n 0.00760615f $X=3.225 $Y=1.44 $X2=0 $Y2=0
cc_161 N_A2_M1001_g N_Y_c_393_n 0.0182396f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A2_M1010_g N_Y_c_393_n 0.0122393f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A2_c_168_n Y 0.00338418f $X=2.725 $Y=1.275 $X2=0 $Y2=0
cc_164 N_A2_M1001_g Y 0.00234478f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_165 A2 Y 0.0246718f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_166 N_A2_c_173_n Y 0.00280543f $X=3.225 $Y=1.44 $X2=0 $Y2=0
cc_167 N_A2_M1001_g N_A_491_367#_c_430_n 0.0114565f $X=2.795 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A2_M1010_g N_A_491_367#_c_430_n 0.0115031f $X=3.225 $Y=2.465 $X2=0
+ $Y2=0
cc_169 A2 N_A_491_367#_c_427_n 0.0171849f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A2_M1010_g N_A_491_367#_c_428_n 0.00114792f $X=3.225 $Y=2.465 $X2=0
+ $Y2=0
cc_171 A2 N_A_491_367#_c_428_n 0.0167518f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_172 N_A2_c_168_n N_A_43_65#_c_464_n 8.71639e-19 $X=2.725 $Y=1.275 $X2=0 $Y2=0
cc_173 A2 N_A_43_65#_c_475_n 0.012853f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A2_c_173_n N_A_43_65#_c_475_n 4.02512e-19 $X=3.225 $Y=1.44 $X2=0 $Y2=0
cc_175 N_A2_c_168_n N_A_43_65#_c_479_n 0.0120955f $X=2.725 $Y=1.275 $X2=0 $Y2=0
cc_176 N_A2_c_170_n N_A_43_65#_c_479_n 0.0120489f $X=3.155 $Y=1.275 $X2=0 $Y2=0
cc_177 A2 N_A_43_65#_c_479_n 0.0430149f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A2_c_173_n N_A_43_65#_c_479_n 5.87177e-19 $X=3.225 $Y=1.44 $X2=0 $Y2=0
cc_179 N_A2_c_170_n N_A_43_65#_c_465_n 4.26518e-19 $X=3.155 $Y=1.275 $X2=0 $Y2=0
cc_180 A2 N_A_43_65#_c_484_n 0.018971f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_181 A2 N_A_43_65#_c_485_n 0.0149232f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A2_c_168_n N_VGND_c_525_n 0.00927214f $X=2.725 $Y=1.275 $X2=0 $Y2=0
cc_183 N_A2_c_170_n N_VGND_c_525_n 0.00888563f $X=3.155 $Y=1.275 $X2=0 $Y2=0
cc_184 N_A2_c_170_n N_VGND_c_526_n 4.78085e-19 $X=3.155 $Y=1.275 $X2=0 $Y2=0
cc_185 N_A2_c_168_n N_VGND_c_527_n 0.00414769f $X=2.725 $Y=1.275 $X2=0 $Y2=0
cc_186 N_A2_c_170_n N_VGND_c_529_n 0.00414769f $X=3.155 $Y=1.275 $X2=0 $Y2=0
cc_187 N_A2_c_168_n N_VGND_c_532_n 0.00813634f $X=2.725 $Y=1.275 $X2=0 $Y2=0
cc_188 N_A2_c_170_n N_VGND_c_532_n 0.0078848f $X=3.155 $Y=1.275 $X2=0 $Y2=0
cc_189 N_A1_M1005_g N_VPWR_c_301_n 0.0168408f $X=3.655 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A1_M1014_g N_VPWR_c_301_n 0.017681f $X=4.085 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A1_M1005_g N_VPWR_c_302_n 0.00486043f $X=3.655 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A1_M1014_g N_VPWR_c_305_n 0.00486043f $X=4.085 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A1_M1005_g N_VPWR_c_299_n 0.0082726f $X=3.655 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A1_M1014_g N_VPWR_c_299_n 0.00934144f $X=4.085 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A1_M1005_g N_A_491_367#_c_427_n 0.0135652f $X=3.655 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A1_M1014_g N_A_491_367#_c_427_n 0.0150277f $X=4.085 $Y=2.465 $X2=0
+ $Y2=0
cc_197 A1 N_A_491_367#_c_427_n 0.041904f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_198 N_A1_c_227_n N_A_491_367#_c_427_n 0.00633497f $X=4.085 $Y=1.44 $X2=0
+ $Y2=0
cc_199 N_A1_c_222_n N_A_43_65#_c_465_n 4.34092e-19 $X=3.585 $Y=1.275 $X2=0 $Y2=0
cc_200 N_A1_c_222_n N_A_43_65#_c_484_n 0.0120955f $X=3.585 $Y=1.275 $X2=0 $Y2=0
cc_201 N_A1_c_224_n N_A_43_65#_c_484_n 0.0120955f $X=4.015 $Y=1.275 $X2=0 $Y2=0
cc_202 A1 N_A_43_65#_c_484_n 0.0124985f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A1_c_227_n N_A_43_65#_c_484_n 0.00230746f $X=4.085 $Y=1.44 $X2=0 $Y2=0
cc_204 A1 N_A_43_65#_c_466_n 0.0219955f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_205 N_A1_c_227_n N_A_43_65#_c_466_n 8.68713e-19 $X=4.085 $Y=1.44 $X2=0 $Y2=0
cc_206 N_A1_c_224_n N_A_43_65#_c_467_n 0.00186805f $X=4.015 $Y=1.275 $X2=0 $Y2=0
cc_207 N_A1_c_222_n N_VGND_c_525_n 4.84056e-19 $X=3.585 $Y=1.275 $X2=0 $Y2=0
cc_208 N_A1_c_222_n N_VGND_c_526_n 0.00879717f $X=3.585 $Y=1.275 $X2=0 $Y2=0
cc_209 N_A1_c_224_n N_VGND_c_526_n 0.0112436f $X=4.015 $Y=1.275 $X2=0 $Y2=0
cc_210 N_A1_c_222_n N_VGND_c_529_n 0.00414769f $X=3.585 $Y=1.275 $X2=0 $Y2=0
cc_211 N_A1_c_224_n N_VGND_c_531_n 0.00414769f $X=4.015 $Y=1.275 $X2=0 $Y2=0
cc_212 N_A1_c_222_n N_VGND_c_532_n 0.0078848f $X=3.585 $Y=1.275 $X2=0 $Y2=0
cc_213 N_A1_c_224_n N_VGND_c_532_n 0.00830694f $X=4.015 $Y=1.275 $X2=0 $Y2=0
cc_214 N_A_43_367#_c_263_n N_VPWR_M1006_d 0.00176461f $X=1.105 $Y=1.86 $X2=-0.19
+ $Y2=1.655
cc_215 N_A_43_367#_c_263_n N_VPWR_c_300_n 0.0170777f $X=1.105 $Y=1.86 $X2=0
+ $Y2=0
cc_216 N_A_43_367#_c_279_p N_VPWR_c_302_n 0.0125234f $X=1.2 $Y=2.905 $X2=0 $Y2=0
cc_217 N_A_43_367#_c_275_n N_VPWR_c_302_n 0.0361172f $X=1.965 $Y=2.99 $X2=0
+ $Y2=0
cc_218 N_A_43_367#_c_265_n N_VPWR_c_302_n 0.0179183f $X=2.095 $Y=2.905 $X2=0
+ $Y2=0
cc_219 N_A_43_367#_c_262_n N_VPWR_c_304_n 0.0178111f $X=0.34 $Y=1.98 $X2=0 $Y2=0
cc_220 N_A_43_367#_M1006_s N_VPWR_c_299_n 0.00371702f $X=0.215 $Y=1.835 $X2=0
+ $Y2=0
cc_221 N_A_43_367#_M1011_s N_VPWR_c_299_n 0.00376627f $X=1.06 $Y=1.835 $X2=0
+ $Y2=0
cc_222 N_A_43_367#_M1009_d N_VPWR_c_299_n 0.00215161f $X=1.92 $Y=1.835 $X2=0
+ $Y2=0
cc_223 N_A_43_367#_c_262_n N_VPWR_c_299_n 0.0100304f $X=0.34 $Y=1.98 $X2=0 $Y2=0
cc_224 N_A_43_367#_c_279_p N_VPWR_c_299_n 0.00738676f $X=1.2 $Y=2.905 $X2=0
+ $Y2=0
cc_225 N_A_43_367#_c_275_n N_VPWR_c_299_n 0.023676f $X=1.965 $Y=2.99 $X2=0 $Y2=0
cc_226 N_A_43_367#_c_265_n N_VPWR_c_299_n 0.0101082f $X=2.095 $Y=2.905 $X2=0
+ $Y2=0
cc_227 N_A_43_367#_c_275_n N_Y_M1000_s 0.00332344f $X=1.965 $Y=2.99 $X2=0 $Y2=0
cc_228 N_A_43_367#_c_275_n N_Y_c_375_n 0.0159805f $X=1.965 $Y=2.99 $X2=0 $Y2=0
cc_229 N_A_43_367#_M1009_d N_Y_c_360_n 2.33864e-19 $X=1.92 $Y=1.835 $X2=0 $Y2=0
cc_230 N_A_43_367#_c_266_n N_Y_c_360_n 0.00183477f $X=2.06 $Y=2.2 $X2=0 $Y2=0
cc_231 N_A_43_367#_c_263_n N_Y_c_361_n 0.00657144f $X=1.105 $Y=1.86 $X2=0 $Y2=0
cc_232 N_A_43_367#_M1009_d Y 0.0021884f $X=1.92 $Y=1.835 $X2=0 $Y2=0
cc_233 N_A_43_367#_c_266_n Y 0.0203341f $X=2.06 $Y=2.2 $X2=0 $Y2=0
cc_234 N_A_43_367#_c_265_n N_A_491_367#_c_425_n 0.0147157f $X=2.095 $Y=2.905
+ $X2=0 $Y2=0
cc_235 N_A_43_367#_c_266_n N_A_491_367#_c_426_n 0.0645429f $X=2.06 $Y=2.2 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_299_n N_Y_M1000_s 0.00225186f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_237 N_VPWR_c_299_n N_Y_M1001_s 0.00225186f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_238 N_VPWR_c_299_n N_A_491_367#_M1001_d 0.00215161f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_239 N_VPWR_c_299_n N_A_491_367#_M1010_d 0.00376627f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_299_n N_A_491_367#_M1014_d 0.00371702f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_302_n N_A_491_367#_c_425_n 0.0179183f $X=3.705 $Y=3.33 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_299_n N_A_491_367#_c_425_n 0.0101082f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_302_n N_A_491_367#_c_430_n 0.0361172f $X=3.705 $Y=3.33 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_299_n N_A_491_367#_c_430_n 0.023676f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_c_302_n N_A_491_367#_c_448_n 0.0125234f $X=3.705 $Y=3.33 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_299_n N_A_491_367#_c_448_n 0.00738676f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_247 N_VPWR_M1005_s N_A_491_367#_c_427_n 0.00176461f $X=3.73 $Y=1.835 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_301_n N_A_491_367#_c_427_n 0.0170777f $X=3.87 $Y=2.12 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_305_n N_A_491_367#_c_429_n 0.0178111f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_299_n N_A_491_367#_c_429_n 0.0100304f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_251 N_Y_c_362_n N_A_491_367#_M1001_d 0.00234752f $X=2.845 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_252 N_Y_c_362_n N_A_491_367#_c_426_n 0.0202165f $X=2.845 $Y=1.78 $X2=0 $Y2=0
cc_253 N_Y_M1001_s N_A_491_367#_c_430_n 0.00332344f $X=2.87 $Y=1.835 $X2=0 $Y2=0
cc_254 N_Y_c_393_n N_A_491_367#_c_430_n 0.0159805f $X=3.01 $Y=1.98 $X2=0 $Y2=0
cc_255 N_Y_c_362_n N_A_491_367#_c_428_n 0.0137028f $X=2.845 $Y=1.78 $X2=0 $Y2=0
cc_256 N_Y_c_365_n N_A_43_65#_M1013_s 0.00525192f $X=2 $Y=0.925 $X2=0 $Y2=0
cc_257 Y N_A_43_65#_M1007_s 0.00247003f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_258 N_Y_c_388_n N_A_43_65#_M1007_s 0.00502944f $X=2.127 $Y=1.03 $X2=0 $Y2=0
cc_259 N_Y_M1002_d N_A_43_65#_c_462_n 0.00172792f $X=1.57 $Y=0.325 $X2=0 $Y2=0
cc_260 N_Y_c_388_n N_A_43_65#_c_462_n 0.0166088f $X=2.127 $Y=1.03 $X2=0 $Y2=0
cc_261 N_Y_c_365_n N_A_43_65#_c_463_n 0.052919f $X=2 $Y=0.925 $X2=0 $Y2=0
cc_262 N_Y_c_362_n N_A_43_65#_c_475_n 7.73326e-19 $X=2.845 $Y=1.78 $X2=0 $Y2=0
cc_263 Y N_A_43_65#_c_475_n 7.9766e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_264 N_Y_c_388_n N_A_43_65#_c_475_n 0.0184727f $X=2.127 $Y=1.03 $X2=0 $Y2=0
cc_265 N_Y_M1012_d N_A_43_65#_c_468_n 0.00176461f $X=0.63 $Y=0.325 $X2=0 $Y2=0
cc_266 N_Y_c_365_n N_A_43_65#_c_468_n 0.0037258f $X=2 $Y=0.925 $X2=0 $Y2=0
cc_267 N_Y_c_358_n N_A_43_65#_c_468_n 0.0158068f $X=0.77 $Y=0.68 $X2=0 $Y2=0
cc_268 N_A_491_367#_c_427_n N_A_43_65#_c_484_n 0.00395032f $X=4.205 $Y=1.78
+ $X2=0 $Y2=0
cc_269 N_A_43_65#_c_479_n N_VGND_M1004_d 0.003325f $X=3.285 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_270 N_A_43_65#_c_484_n N_VGND_M1003_d 0.00418232f $X=4.135 $Y=0.955 $X2=0
+ $Y2=0
cc_271 N_A_43_65#_c_464_n N_VGND_c_525_n 0.0181085f $X=2.515 $Y=0.65 $X2=0 $Y2=0
cc_272 N_A_43_65#_c_479_n N_VGND_c_525_n 0.0170777f $X=3.285 $Y=0.955 $X2=0
+ $Y2=0
cc_273 N_A_43_65#_c_465_n N_VGND_c_525_n 0.014127f $X=3.37 $Y=0.48 $X2=0 $Y2=0
cc_274 N_A_43_65#_c_465_n N_VGND_c_526_n 0.0147877f $X=3.37 $Y=0.48 $X2=0 $Y2=0
cc_275 N_A_43_65#_c_484_n N_VGND_c_526_n 0.0170777f $X=4.135 $Y=0.955 $X2=0
+ $Y2=0
cc_276 N_A_43_65#_c_467_n N_VGND_c_526_n 0.0148073f $X=4.23 $Y=0.48 $X2=0 $Y2=0
cc_277 N_A_43_65#_c_461_n N_VGND_c_527_n 0.0186386f $X=0.435 $Y=0.34 $X2=0 $Y2=0
cc_278 N_A_43_65#_c_464_n N_VGND_c_527_n 0.0129036f $X=2.515 $Y=0.65 $X2=0 $Y2=0
cc_279 N_A_43_65#_c_468_n N_VGND_c_527_n 0.13146f $X=1.105 $Y=0.452 $X2=0 $Y2=0
cc_280 N_A_43_65#_c_465_n N_VGND_c_529_n 0.00923511f $X=3.37 $Y=0.48 $X2=0 $Y2=0
cc_281 N_A_43_65#_c_467_n N_VGND_c_531_n 0.0133857f $X=4.23 $Y=0.48 $X2=0 $Y2=0
cc_282 N_A_43_65#_c_461_n N_VGND_c_532_n 0.0101082f $X=0.435 $Y=0.34 $X2=0 $Y2=0
cc_283 N_A_43_65#_c_464_n N_VGND_c_532_n 0.00699798f $X=2.515 $Y=0.65 $X2=0
+ $Y2=0
cc_284 N_A_43_65#_c_465_n N_VGND_c_532_n 0.00670918f $X=3.37 $Y=0.48 $X2=0 $Y2=0
cc_285 N_A_43_65#_c_467_n N_VGND_c_532_n 0.00972454f $X=4.23 $Y=0.48 $X2=0 $Y2=0
cc_286 N_A_43_65#_c_468_n N_VGND_c_532_n 0.0730233f $X=1.105 $Y=0.452 $X2=0
+ $Y2=0
