* File: sky130_fd_sc_lp__sdfrtp_lp2.pxi.spice
* Created: Wed Sep  2 10:34:59 2020
* 
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_81_194# N_A_81_194#_M1013_d
+ N_A_81_194#_M1023_d N_A_81_194#_M1000_g N_A_81_194#_M1030_g
+ N_A_81_194#_c_282_n N_A_81_194#_c_283_n N_A_81_194#_c_284_n
+ N_A_81_194#_c_285_n N_A_81_194#_c_286_n N_A_81_194#_c_287_n
+ N_A_81_194#_c_288_n N_A_81_194#_c_289_n N_A_81_194#_c_342_p
+ N_A_81_194#_c_290_n N_A_81_194#_c_296_n N_A_81_194#_c_291_n
+ PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_81_194#
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%D N_D_c_395_n N_D_M1001_g N_D_M1043_g D
+ PM_SKY130_FD_SC_LP__SDFRTP_LP2%D
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%SCE N_SCE_M1018_g N_SCE_M1010_g N_SCE_c_429_n
+ N_SCE_M1025_g N_SCE_M1023_g N_SCE_c_430_n N_SCE_M1013_g N_SCE_c_431_n
+ N_SCE_c_438_n N_SCE_c_432_n N_SCE_c_433_n SCE N_SCE_c_434_n N_SCE_c_442_n
+ N_SCE_c_435_n N_SCE_c_436_n PM_SKY130_FD_SC_LP__SDFRTP_LP2%SCE
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%SCD N_SCD_M1044_g N_SCD_M1041_g SCD
+ N_SCD_c_537_n PM_SKY130_FD_SC_LP__SDFRTP_LP2%SCD
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%CLK N_CLK_M1015_g N_CLK_M1031_g N_CLK_M1032_g
+ CLK N_CLK_c_574_n PM_SKY130_FD_SC_LP__SDFRTP_LP2%CLK
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_1147_408# N_A_1147_408#_M1038_d
+ N_A_1147_408#_M1016_d N_A_1147_408#_c_608_n N_A_1147_408#_c_625_n
+ N_A_1147_408#_M1019_g N_A_1147_408#_c_609_n N_A_1147_408#_M1008_g
+ N_A_1147_408#_M1039_g N_A_1147_408#_c_610_n N_A_1147_408#_c_611_n
+ N_A_1147_408#_c_612_n N_A_1147_408#_c_613_n N_A_1147_408#_c_628_n
+ N_A_1147_408#_M1037_g N_A_1147_408#_c_614_n N_A_1147_408#_c_630_n
+ N_A_1147_408#_c_615_n N_A_1147_408#_c_616_n N_A_1147_408#_c_617_n
+ N_A_1147_408#_c_618_n N_A_1147_408#_c_667_p N_A_1147_408#_c_619_n
+ N_A_1147_408#_c_620_n N_A_1147_408#_c_621_n N_A_1147_408#_c_622_n
+ N_A_1147_408#_c_623_n PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_1147_408#
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_1605_93# N_A_1605_93#_M1033_d
+ N_A_1605_93#_M1006_d N_A_1605_93#_c_782_n N_A_1605_93#_M1026_g
+ N_A_1605_93#_c_793_n N_A_1605_93#_M1045_g N_A_1605_93#_c_783_n
+ N_A_1605_93#_c_784_n N_A_1605_93#_c_785_n N_A_1605_93#_c_786_n
+ N_A_1605_93#_c_787_n N_A_1605_93#_c_812_n N_A_1605_93#_c_788_n
+ N_A_1605_93#_c_789_n N_A_1605_93#_c_796_n N_A_1605_93#_c_790_n
+ N_A_1605_93#_c_791_n N_A_1605_93#_c_797_n N_A_1605_93#_c_792_n
+ PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_1605_93#
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%RESET_B N_RESET_B_M1011_g N_RESET_B_c_907_n
+ N_RESET_B_c_908_n N_RESET_B_c_909_n N_RESET_B_c_910_n N_RESET_B_M1009_g
+ N_RESET_B_M1021_g N_RESET_B_c_912_n N_RESET_B_c_913_n N_RESET_B_M1024_g
+ N_RESET_B_M1012_g N_RESET_B_M1028_g N_RESET_B_c_915_n N_RESET_B_c_916_n
+ N_RESET_B_c_917_n N_RESET_B_c_934_n N_RESET_B_c_918_n N_RESET_B_c_919_n
+ N_RESET_B_c_920_n N_RESET_B_c_921_n N_RESET_B_c_939_n RESET_B
+ N_RESET_B_c_923_n N_RESET_B_c_924_n N_RESET_B_c_925_n N_RESET_B_c_926_n
+ N_RESET_B_c_927_n PM_SKY130_FD_SC_LP__SDFRTP_LP2%RESET_B
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_1432_119# N_A_1432_119#_M1014_d
+ N_A_1432_119#_M1019_d N_A_1432_119#_M1024_d N_A_1432_119#_c_1173_n
+ N_A_1432_119#_M1022_g N_A_1432_119#_M1033_g N_A_1432_119#_c_1174_n
+ N_A_1432_119#_c_1175_n N_A_1432_119#_M1006_g N_A_1432_119#_c_1176_n
+ N_A_1432_119#_c_1177_n N_A_1432_119#_c_1183_n N_A_1432_119#_c_1205_n
+ N_A_1432_119#_c_1184_n N_A_1432_119#_c_1185_n N_A_1432_119#_c_1186_n
+ N_A_1432_119#_c_1178_n N_A_1432_119#_c_1206_n
+ PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_1432_119#
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_876_119# N_A_876_119#_M1015_s
+ N_A_876_119#_M1031_s N_A_876_119#_M1016_g N_A_876_119#_c_1286_n
+ N_A_876_119#_M1029_g N_A_876_119#_M1038_g N_A_876_119#_c_1300_n
+ N_A_876_119#_c_1288_n N_A_876_119#_c_1301_n N_A_876_119#_c_1302_n
+ N_A_876_119#_c_1289_n N_A_876_119#_M1014_g N_A_876_119#_M1042_g
+ N_A_876_119#_c_1304_n N_A_876_119#_M1002_g N_A_876_119#_M1020_g
+ N_A_876_119#_c_1306_n N_A_876_119#_c_1292_n N_A_876_119#_c_1308_n
+ N_A_876_119#_c_1309_n N_A_876_119#_c_1293_n N_A_876_119#_c_1294_n
+ N_A_876_119#_c_1295_n N_A_876_119#_c_1296_n N_A_876_119#_c_1311_n
+ N_A_876_119#_c_1297_n N_A_876_119#_c_1298_n
+ PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_876_119#
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_2435_296# N_A_2435_296#_M1027_d
+ N_A_2435_296#_M1028_d N_A_2435_296#_M1003_g N_A_2435_296#_M1034_g
+ N_A_2435_296#_c_1472_n N_A_2435_296#_c_1473_n N_A_2435_296#_c_1474_n
+ N_A_2435_296#_c_1475_n N_A_2435_296#_c_1476_n N_A_2435_296#_c_1477_n
+ N_A_2435_296#_c_1499_n N_A_2435_296#_c_1478_n N_A_2435_296#_c_1479_n
+ N_A_2435_296#_c_1480_n PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_2435_296#
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_2092_47# N_A_2092_47#_M1039_d
+ N_A_2092_47#_M1002_d N_A_2092_47#_c_1567_n N_A_2092_47#_M1027_g
+ N_A_2092_47#_M1004_g N_A_2092_47#_c_1569_n N_A_2092_47#_c_1570_n
+ N_A_2092_47#_c_1571_n N_A_2092_47#_M1035_g N_A_2092_47#_c_1572_n
+ N_A_2092_47#_M1005_g N_A_2092_47#_c_1574_n N_A_2092_47#_M1017_g
+ N_A_2092_47#_c_1583_n N_A_2092_47#_c_1584_n N_A_2092_47#_c_1585_n
+ N_A_2092_47#_c_1575_n N_A_2092_47#_c_1576_n N_A_2092_47#_c_1577_n
+ N_A_2092_47#_c_1578_n N_A_2092_47#_c_1579_n N_A_2092_47#_c_1580_n
+ PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_2092_47#
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_2863_90# N_A_2863_90#_M1035_s
+ N_A_2863_90#_M1005_s N_A_2863_90#_M1040_g N_A_2863_90#_M1007_g
+ N_A_2863_90#_M1036_g N_A_2863_90#_c_1725_n N_A_2863_90#_c_1726_n
+ N_A_2863_90#_c_1727_n N_A_2863_90#_c_1735_n N_A_2863_90#_c_1728_n
+ N_A_2863_90#_c_1729_n N_A_2863_90#_c_1730_n N_A_2863_90#_c_1731_n
+ N_A_2863_90#_c_1732_n PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_2863_90#
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_116_419# N_A_116_419#_M1043_d
+ N_A_116_419#_M1014_s N_A_116_419#_M1001_s N_A_116_419#_M1030_d
+ N_A_116_419#_M1019_s N_A_116_419#_c_1793_n N_A_116_419#_c_1805_n
+ N_A_116_419#_c_1806_n N_A_116_419#_c_1835_n N_A_116_419#_c_1799_n
+ N_A_116_419#_c_1836_n N_A_116_419#_c_1845_n N_A_116_419#_c_1800_n
+ N_A_116_419#_c_1846_n N_A_116_419#_c_1794_n N_A_116_419#_c_1801_n
+ N_A_116_419#_c_1795_n N_A_116_419#_c_1803_n N_A_116_419#_c_1796_n
+ N_A_116_419#_c_1797_n N_A_116_419#_c_1813_n N_A_116_419#_c_1817_n
+ N_A_116_419#_c_1818_n N_A_116_419#_c_1798_n
+ PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_116_419#
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%VPWR N_VPWR_M1018_d N_VPWR_M1009_d
+ N_VPWR_M1031_d N_VPWR_M1045_d N_VPWR_M1006_s N_VPWR_M1003_d N_VPWR_M1004_d
+ N_VPWR_M1005_d N_VPWR_c_1934_n N_VPWR_c_1935_n N_VPWR_c_1936_n N_VPWR_c_1937_n
+ N_VPWR_c_1938_n N_VPWR_c_1939_n N_VPWR_c_1940_n N_VPWR_c_1941_n
+ N_VPWR_c_1942_n N_VPWR_c_1943_n N_VPWR_c_1944_n N_VPWR_c_1945_n
+ N_VPWR_c_1946_n N_VPWR_c_1947_n N_VPWR_c_1948_n VPWR N_VPWR_c_1949_n
+ N_VPWR_c_1950_n N_VPWR_c_1951_n N_VPWR_c_1952_n N_VPWR_c_1953_n
+ N_VPWR_c_1933_n N_VPWR_c_1955_n N_VPWR_c_1956_n N_VPWR_c_1957_n
+ N_VPWR_c_1958_n N_VPWR_c_1959_n PM_SKY130_FD_SC_LP__SDFRTP_LP2%VPWR
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%Q N_Q_M1036_d N_Q_M1007_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__SDFRTP_LP2%Q
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%noxref_23 N_noxref_23_M1000_s
+ N_noxref_23_M1044_d N_noxref_23_c_2134_n N_noxref_23_c_2135_n
+ N_noxref_23_c_2136_n PM_SKY130_FD_SC_LP__SDFRTP_LP2%noxref_23
x_PM_SKY130_FD_SC_LP__SDFRTP_LP2%VGND N_VGND_M1011_d N_VGND_M1032_d
+ N_VGND_M1021_d N_VGND_M1034_d N_VGND_M1017_d N_VGND_c_2163_n N_VGND_c_2164_n
+ N_VGND_c_2165_n N_VGND_c_2166_n N_VGND_c_2167_n N_VGND_c_2168_n VGND
+ N_VGND_c_2169_n N_VGND_c_2170_n N_VGND_c_2171_n N_VGND_c_2172_n
+ N_VGND_c_2173_n N_VGND_c_2174_n N_VGND_c_2175_n N_VGND_c_2176_n
+ N_VGND_c_2177_n N_VGND_c_2178_n N_VGND_c_2179_n
+ PM_SKY130_FD_SC_LP__SDFRTP_LP2%VGND
cc_1 VNB N_A_81_194#_c_282_n 0.03528f $X=-0.19 $Y=-0.245 $X2=2.435 $Y2=1.185
cc_2 VNB N_A_81_194#_c_283_n 0.00410706f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_3 VNB N_A_81_194#_c_284_n 0.017297f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_4 VNB N_A_81_194#_c_285_n 0.0190756f $X=-0.19 $Y=-0.245 $X2=3.82 $Y2=1.185
cc_5 VNB N_A_81_194#_c_286_n 0.00901596f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=0.76
cc_6 VNB N_A_81_194#_c_287_n 0.00868742f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=2.075
cc_7 VNB N_A_81_194#_c_288_n 0.0386032f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.135
cc_8 VNB N_A_81_194#_c_289_n 0.0016706f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.135
cc_9 VNB N_A_81_194#_c_290_n 0.00564402f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=1.185
cc_10 VNB N_A_81_194#_c_291_n 0.0179578f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.97
cc_11 VNB N_D_c_395_n 0.0229277f $X=-0.19 $Y=-0.245 $X2=3.845 $Y2=0.595
cc_12 VNB N_D_M1043_g 0.0484768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB D 0.00169913f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.65
cc_14 VNB N_SCE_M1010_g 0.0506883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_c_429_n 0.0157583f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.65
cc_16 VNB N_SCE_c_430_n 0.0169093f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_17 VNB N_SCE_c_431_n 0.023813f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=1.1
cc_18 VNB N_SCE_c_432_n 0.0029964f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=2.075
cc_19 VNB N_SCE_c_433_n 0.0105811f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.135
cc_20 VNB N_SCE_c_434_n 0.00802125f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.185
cc_21 VNB N_SCE_c_435_n 0.0196271f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=2.2
cc_22 VNB N_SCE_c_436_n 0.00567888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_SCD_M1044_g 0.0399378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB SCD 0.00332077f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.65
cc_25 VNB N_SCD_c_537_n 0.0159484f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=2.595
cc_26 VNB N_CLK_M1015_g 0.0205713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_CLK_M1031_g 0.0120518f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.97
cc_28 VNB N_CLK_M1032_g 0.018075f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=2.595
cc_29 VNB CLK 0.00272402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_CLK_c_574_n 0.0380381f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_31 VNB N_A_1147_408#_c_608_n 0.0123904f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.97
cc_32 VNB N_A_1147_408#_c_609_n 0.0159575f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=2.595
cc_33 VNB N_A_1147_408#_c_610_n 0.0768716f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_34 VNB N_A_1147_408#_c_611_n 0.0329701f $X=-0.19 $Y=-0.245 $X2=3.82 $Y2=1.185
cc_35 VNB N_A_1147_408#_c_612_n 0.0123448f $X=-0.19 $Y=-0.245 $X2=2.765
+ $Y2=1.185
cc_36 VNB N_A_1147_408#_c_613_n 0.00147711f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=1.1
cc_37 VNB N_A_1147_408#_c_614_n 6.61405e-19 $X=-0.19 $Y=-0.245 $X2=0.57
+ $Y2=1.135
cc_38 VNB N_A_1147_408#_c_615_n 0.0107215f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.185
cc_39 VNB N_A_1147_408#_c_616_n 0.00155339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1147_408#_c_617_n 0.053294f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=2.2
cc_41 VNB N_A_1147_408#_c_618_n 0.00703086f $X=-0.19 $Y=-0.245 $X2=0.57
+ $Y2=1.135
cc_42 VNB N_A_1147_408#_c_619_n 0.0013366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1147_408#_c_620_n 4.14555e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1147_408#_c_621_n 0.0138151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1147_408#_c_622_n 0.0349114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1147_408#_c_623_n 0.0181186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1605_93#_c_782_n 0.0168083f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.97
cc_48 VNB N_A_1605_93#_c_783_n 0.00446971f $X=-0.19 $Y=-0.245 $X2=0.735
+ $Y2=1.185
cc_49 VNB N_A_1605_93#_c_784_n 0.00139786f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_50 VNB N_A_1605_93#_c_785_n 0.0507579f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_51 VNB N_A_1605_93#_c_786_n 0.00967717f $X=-0.19 $Y=-0.245 $X2=3.82 $Y2=1.185
cc_52 VNB N_A_1605_93#_c_787_n 9.52647e-19 $X=-0.19 $Y=-0.245 $X2=2.765
+ $Y2=1.185
cc_53 VNB N_A_1605_93#_c_788_n 0.00763836f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=1.27
cc_54 VNB N_A_1605_93#_c_789_n 0.0124244f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.135
cc_55 VNB N_A_1605_93#_c_790_n 0.00499693f $X=-0.19 $Y=-0.245 $X2=4 $Y2=2.24
cc_56 VNB N_A_1605_93#_c_791_n 0.00104694f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.135
cc_57 VNB N_A_1605_93#_c_792_n 7.46876e-19 $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_58 VNB N_RESET_B_M1011_g 0.0224545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_RESET_B_c_907_n 0.495286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_RESET_B_c_908_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_RESET_B_c_909_n 0.0423859f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.97
cc_62 VNB N_RESET_B_c_910_n 0.00742257f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.65
cc_63 VNB N_RESET_B_M1021_g 0.0111631f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_64 VNB N_RESET_B_c_912_n 0.0151245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_RESET_B_c_913_n 0.0199934f $X=-0.19 $Y=-0.245 $X2=3.82 $Y2=1.185
cc_66 VNB N_RESET_B_M1012_g 0.0655005f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=1.27
cc_67 VNB N_RESET_B_c_915_n 0.0271475f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.135
cc_68 VNB N_RESET_B_c_916_n 0.00236187f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=1.185
cc_69 VNB N_RESET_B_c_917_n 7.41492e-19 $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=2.2
cc_70 VNB N_RESET_B_c_918_n 0.00986344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_RESET_B_c_919_n 0.0256008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_RESET_B_c_920_n 8.38669e-19 $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.78
cc_73 VNB N_RESET_B_c_921_n 0.00334239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB RESET_B 0.00390629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_RESET_B_c_923_n 0.0184185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_RESET_B_c_924_n 0.0016928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_RESET_B_c_925_n 0.0130433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_RESET_B_c_926_n 0.00333863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_RESET_B_c_927_n 0.00267956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1432_119#_c_1173_n 0.0296131f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=1.78
cc_81 VNB N_A_1432_119#_c_1174_n 0.0255398f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.27
cc_82 VNB N_A_1432_119#_c_1175_n 0.00721316f $X=-0.19 $Y=-0.245 $X2=2.6
+ $Y2=1.615
cc_83 VNB N_A_1432_119#_c_1176_n 0.0204536f $X=-0.19 $Y=-0.245 $X2=4.022
+ $Y2=0.76
cc_84 VNB N_A_1432_119#_c_1177_n 0.00398111f $X=-0.19 $Y=-0.245 $X2=4.14
+ $Y2=2.075
cc_85 VNB N_A_1432_119#_c_1178_n 0.046699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_876_119#_c_1286_n 0.0169027f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=2.595
cc_87 VNB N_A_876_119#_M1029_g 0.0186189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_876_119#_c_1288_n 0.0589914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_876_119#_c_1289_n 0.0192581f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=0.76
cc_90 VNB N_A_876_119#_M1002_g 0.00482222f $X=-0.19 $Y=-0.245 $X2=4 $Y2=2.2
cc_91 VNB N_A_876_119#_M1020_g 0.0298656f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=2.2
cc_92 VNB N_A_876_119#_c_1292_n 0.0142346f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_93 VNB N_A_876_119#_c_1293_n 0.00317201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_876_119#_c_1294_n 0.0638132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_876_119#_c_1295_n 0.0111047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_876_119#_c_1296_n 0.0306823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_876_119#_c_1297_n 0.00556563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_876_119#_c_1298_n 0.0345097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2435_296#_M1003_g 0.00161517f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.65
cc_100 VNB N_A_2435_296#_M1034_g 0.0347366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2435_296#_c_1472_n 0.0108744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2435_296#_c_1473_n 0.00690447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2435_296#_c_1474_n 0.00419711f $X=-0.19 $Y=-0.245 $X2=0.57
+ $Y2=1.135
cc_104 VNB N_A_2435_296#_c_1475_n 0.00988273f $X=-0.19 $Y=-0.245 $X2=0.735
+ $Y2=1.135
cc_105 VNB N_A_2435_296#_c_1476_n 0.00138697f $X=-0.19 $Y=-0.245 $X2=2.6
+ $Y2=1.185
cc_106 VNB N_A_2435_296#_c_1477_n 0.00338231f $X=-0.19 $Y=-0.245 $X2=4.022
+ $Y2=1.185
cc_107 VNB N_A_2435_296#_c_1478_n 0.00223477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2435_296#_c_1479_n 8.41942e-19 $X=-0.19 $Y=-0.245 $X2=4.14
+ $Y2=2.2
cc_109 VNB N_A_2435_296#_c_1480_n 0.0833311f $X=-0.19 $Y=-0.245 $X2=0.57
+ $Y2=1.135
cc_110 VNB N_A_2092_47#_c_1567_n 0.0193374f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.97
cc_111 VNB N_A_2092_47#_M1004_g 0.0429535f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=2.595
cc_112 VNB N_A_2092_47#_c_1569_n 0.0460167f $X=-0.19 $Y=-0.245 $X2=2.435
+ $Y2=1.185
cc_113 VNB N_A_2092_47#_c_1570_n 0.0450184f $X=-0.19 $Y=-0.245 $X2=0.735
+ $Y2=1.185
cc_114 VNB N_A_2092_47#_c_1571_n 0.0153502f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.27
cc_115 VNB N_A_2092_47#_c_1572_n 0.0196213f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_116 VNB N_A_2092_47#_M1005_g 0.0371589f $X=-0.19 $Y=-0.245 $X2=3.82 $Y2=1.185
cc_117 VNB N_A_2092_47#_c_1574_n 0.0132698f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=1.1
cc_118 VNB N_A_2092_47#_c_1575_n 0.00611448f $X=-0.19 $Y=-0.245 $X2=4 $Y2=2.24
cc_119 VNB N_A_2092_47#_c_1576_n 0.00469329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2092_47#_c_1577_n 0.0190014f $X=-0.19 $Y=-0.245 $X2=0.57
+ $Y2=1.135
cc_121 VNB N_A_2092_47#_c_1578_n 0.00475512f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.78
cc_122 VNB N_A_2092_47#_c_1579_n 0.0019942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2092_47#_c_1580_n 0.00255276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2863_90#_M1040_g 0.0194549f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.65
cc_125 VNB N_A_2863_90#_M1036_g 0.0254568f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_126 VNB N_A_2863_90#_c_1725_n 0.0255792f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=1.1
cc_127 VNB N_A_2863_90#_c_1726_n 0.0059029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_2863_90#_c_1727_n 0.0115161f $X=-0.19 $Y=-0.245 $X2=4.14
+ $Y2=2.075
cc_129 VNB N_A_2863_90#_c_1728_n 0.00796797f $X=-0.19 $Y=-0.245 $X2=4.022
+ $Y2=1.185
cc_130 VNB N_A_2863_90#_c_1729_n 0.00159225f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=2.2
cc_131 VNB N_A_2863_90#_c_1730_n 0.0267614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_2863_90#_c_1731_n 0.00428173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_2863_90#_c_1732_n 0.006901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_116_419#_c_1793_n 0.00876179f $X=-0.19 $Y=-0.245 $X2=2.6
+ $Y2=1.615
cc_135 VNB N_A_116_419#_c_1794_n 0.00561762f $X=-0.19 $Y=-0.245 $X2=4 $Y2=2.2
cc_136 VNB N_A_116_419#_c_1795_n 0.00385321f $X=-0.19 $Y=-0.245 $X2=0.57
+ $Y2=1.135
cc_137 VNB N_A_116_419#_c_1796_n 0.0423211f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_138 VNB N_A_116_419#_c_1797_n 4.16014e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_116_419#_c_1798_n 9.50902e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VPWR_c_1933_n 0.681144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB Q 0.0573351f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.97
cc_142 VNB N_noxref_23_c_2134_n 0.0251215f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.97
cc_143 VNB N_noxref_23_c_2135_n 0.00257084f $X=-0.19 $Y=-0.245 $X2=2.59
+ $Y2=2.595
cc_144 VNB N_noxref_23_c_2136_n 0.00779889f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.27
cc_145 VNB N_VGND_c_2163_n 0.00928975f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.615
cc_146 VNB N_VGND_c_2164_n 0.0191232f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=1.185
cc_147 VNB N_VGND_c_2165_n 0.0941644f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=0.76
cc_148 VNB N_VGND_c_2166_n 0.005594f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=2.075
cc_149 VNB N_VGND_c_2167_n 0.00564356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2168_n 0.0195226f $X=-0.19 $Y=-0.245 $X2=4 $Y2=2.2
cc_151 VNB N_VGND_c_2169_n 0.061839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2170_n 0.0689795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2171_n 0.0918811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2172_n 0.0578252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2173_n 0.0287523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2174_n 0.786669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2175_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2176_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2177_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2178_n 0.00631708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2179_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VPB N_A_81_194#_M1030_g 0.0342249f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=2.595
cc_163 VPB N_A_81_194#_c_283_n 7.46894e-19 $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.615
cc_164 VPB N_A_81_194#_c_284_n 0.010739f $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.615
cc_165 VPB N_A_81_194#_c_287_n 0.00869139f $X=-0.19 $Y=1.655 $X2=4.14 $Y2=2.075
cc_166 VPB N_A_81_194#_c_296_n 0.006957f $X=-0.19 $Y=1.655 $X2=4.14 $Y2=2.2
cc_167 VPB N_D_c_395_n 0.0636217f $X=-0.19 $Y=1.655 $X2=3.845 $Y2=0.595
cc_168 VPB D 0.00217111f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.65
cc_169 VPB N_SCE_M1023_g 0.0325439f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.185
cc_170 VPB N_SCE_c_438_n 0.022168f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=0.76
cc_171 VPB N_SCE_c_432_n 0.00430981f $X=-0.19 $Y=1.655 $X2=4.14 $Y2=2.075
cc_172 VPB N_SCE_c_433_n 0.019848f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.135
cc_173 VPB N_SCE_c_434_n 0.0245257f $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.185
cc_174 VPB N_SCE_c_442_n 0.0193061f $X=-0.19 $Y=1.655 $X2=4 $Y2=2.24
cc_175 VPB N_SCE_c_436_n 0.00471402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_SCD_M1041_g 0.0344486f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.97
cc_177 VPB SCD 0.00187299f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.65
cc_178 VPB N_SCD_c_537_n 0.00888613f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=2.595
cc_179 VPB N_CLK_M1031_g 0.0485364f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.97
cc_180 VPB N_A_1147_408#_c_608_n 0.0215704f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.97
cc_181 VPB N_A_1147_408#_c_625_n 0.0215383f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.65
cc_182 VPB N_A_1147_408#_c_612_n 0.0058656f $X=-0.19 $Y=1.655 $X2=2.765
+ $Y2=1.185
cc_183 VPB N_A_1147_408#_c_613_n 0.00833623f $X=-0.19 $Y=1.655 $X2=4.022 $Y2=1.1
cc_184 VPB N_A_1147_408#_c_628_n 0.0329621f $X=-0.19 $Y=1.655 $X2=4.022 $Y2=0.76
cc_185 VPB N_A_1147_408#_c_614_n 0.0110787f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.135
cc_186 VPB N_A_1147_408#_c_630_n 0.0135568f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.135
cc_187 VPB N_A_1147_408#_c_617_n 0.017323f $X=-0.19 $Y=1.655 $X2=4.14 $Y2=2.2
cc_188 VPB N_A_1147_408#_c_620_n 0.00558667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1147_408#_c_621_n 0.020354f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_1605_93#_c_793_n 0.0184849f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=2.595
cc_191 VPB N_A_1605_93#_c_783_n 0.00573561f $X=-0.19 $Y=1.655 $X2=0.735
+ $Y2=1.185
cc_192 VPB N_A_1605_93#_c_784_n 0.00151527f $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.615
cc_193 VPB N_A_1605_93#_c_796_n 0.00346344f $X=-0.19 $Y=1.655 $X2=4.022
+ $Y2=1.185
cc_194 VPB N_A_1605_93#_c_797_n 0.00251237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_1605_93#_c_792_n 0.00183665f $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.615
cc_196 VPB N_RESET_B_M1009_g 0.0352226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_RESET_B_c_913_n 0.00506436f $X=-0.19 $Y=1.655 $X2=3.82 $Y2=1.185
cc_198 VPB N_RESET_B_M1024_g 0.0261112f $X=-0.19 $Y=1.655 $X2=4.022 $Y2=1.1
cc_199 VPB N_RESET_B_M1028_g 0.0299329f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.135
cc_200 VPB N_RESET_B_c_916_n 0.00945914f $X=-0.19 $Y=1.655 $X2=4.022 $Y2=1.185
cc_201 VPB N_RESET_B_c_917_n 0.00249385f $X=-0.19 $Y=1.655 $X2=4.14 $Y2=2.2
cc_202 VPB N_RESET_B_c_934_n 0.00234029f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.97
cc_203 VPB N_RESET_B_c_918_n 0.0274408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_RESET_B_c_919_n 0.0288492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_RESET_B_c_920_n 0.00128647f $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.78
cc_206 VPB N_RESET_B_c_921_n 0.0291497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_939_n 9.59019e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB RESET_B 8.16694e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_RESET_B_c_923_n 0.00973311f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_RESET_B_c_924_n 5.08785e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_RESET_B_c_926_n 0.00372371f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_RESET_B_c_927_n 0.00820576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_1432_119#_c_1174_n 0.0175813f $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.27
cc_214 VPB N_A_1432_119#_c_1175_n 0.0203653f $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.615
cc_215 VPB N_A_1432_119#_M1006_g 0.0240243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_1432_119#_c_1177_n 2.66138e-19 $X=-0.19 $Y=1.655 $X2=4.14
+ $Y2=2.075
cc_217 VPB N_A_1432_119#_c_1183_n 0.0031176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_1432_119#_c_1184_n 0.00611774f $X=-0.19 $Y=1.655 $X2=4 $Y2=2.2
cc_219 VPB N_A_1432_119#_c_1185_n 0.0130798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_1432_119#_c_1186_n 0.0022087f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.97
cc_221 VPB N_A_876_119#_M1016_g 0.0304345f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.65
cc_222 VPB N_A_876_119#_c_1300_n 0.0785294f $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.615
cc_223 VPB N_A_876_119#_c_1301_n 0.125339f $X=-0.19 $Y=1.655 $X2=2.765 $Y2=1.185
cc_224 VPB N_A_876_119#_c_1302_n 0.0109006f $X=-0.19 $Y=1.655 $X2=4.022 $Y2=1.1
cc_225 VPB N_A_876_119#_M1042_g 0.0427198f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.135
cc_226 VPB N_A_876_119#_c_1304_n 0.22801f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.135
cc_227 VPB N_A_876_119#_M1002_g 0.0403494f $X=-0.19 $Y=1.655 $X2=4 $Y2=2.2
cc_228 VPB N_A_876_119#_c_1306_n 0.0124845f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.135
cc_229 VPB N_A_876_119#_c_1292_n 5.10071e-19 $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.615
cc_230 VPB N_A_876_119#_c_1308_n 0.0119428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_876_119#_c_1309_n 0.0162874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_876_119#_c_1294_n 0.0272392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_876_119#_c_1311_n 0.00293347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_2435_296#_M1003_g 0.0487141f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.65
cc_235 VPB N_A_2435_296#_c_1478_n 0.0029109f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_2092_47#_M1004_g 0.0477007f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=2.595
cc_237 VPB N_A_2092_47#_M1005_g 0.0359132f $X=-0.19 $Y=1.655 $X2=3.82 $Y2=1.185
cc_238 VPB N_A_2092_47#_c_1583_n 0.00182603f $X=-0.19 $Y=1.655 $X2=0.57
+ $Y2=1.135
cc_239 VPB N_A_2092_47#_c_1584_n 0.00626883f $X=-0.19 $Y=1.655 $X2=0.57
+ $Y2=1.135
cc_240 VPB N_A_2092_47#_c_1585_n 0.0150922f $X=-0.19 $Y=1.655 $X2=4.022
+ $Y2=1.185
cc_241 VPB N_A_2863_90#_M1007_g 0.0315967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_2863_90#_c_1726_n 0.00855513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_2863_90#_c_1735_n 0.0182654f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.135
cc_244 VPB N_A_2863_90#_c_1728_n 0.00353624f $X=-0.19 $Y=1.655 $X2=4.022
+ $Y2=1.185
cc_245 VPB N_A_2863_90#_c_1732_n 0.00182437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_116_419#_c_1799_n 0.0146942f $X=-0.19 $Y=1.655 $X2=4.14 $Y2=2.075
cc_247 VPB N_A_116_419#_c_1800_n 0.0231483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_116_419#_c_1801_n 0.00192193f $X=-0.19 $Y=1.655 $X2=4.14 $Y2=2.2
cc_249 VPB N_A_116_419#_c_1795_n 0.00296716f $X=-0.19 $Y=1.655 $X2=0.57
+ $Y2=1.135
cc_250 VPB N_A_116_419#_c_1803_n 0.0767979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_116_419#_c_1796_n 0.021758f $X=-0.19 $Y=1.655 $X2=2.6 $Y2=1.615
cc_252 VPB N_VPWR_c_1934_n 0.00283226f $X=-0.19 $Y=1.655 $X2=4.14 $Y2=1.27
cc_253 VPB N_VPWR_c_1935_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.135
cc_254 VPB N_VPWR_c_1936_n 0.00430263f $X=-0.19 $Y=1.655 $X2=4.022 $Y2=1.185
cc_255 VPB N_VPWR_c_1937_n 0.011031f $X=-0.19 $Y=1.655 $X2=4.14 $Y2=2.2
cc_256 VPB N_VPWR_c_1938_n 0.0325377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1939_n 0.00495263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1940_n 0.0214777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1941_n 0.0212426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1942_n 0.00766088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1943_n 0.0366879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1944_n 0.00510188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1945_n 0.0385904f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1946_n 0.0055215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1947_n 0.056191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1948_n 0.00356964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1949_n 0.0440132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1950_n 0.0870465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1951_n 0.0327942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1952_n 0.0380084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1953_n 0.0257698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1933_n 0.0867088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1955_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1956_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1957_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1958_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1959_n 0.00626055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB Q 0.0154973f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.97
cc_279 VPB Q 0.0173545f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=2.595
cc_280 VPB Q 0.0419835f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=2.595
cc_281 N_A_81_194#_c_282_n N_D_c_395_n 0.00564987f $X=2.435 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_282 N_A_81_194#_c_288_n N_D_c_395_n 0.0102465f $X=0.57 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_283 N_A_81_194#_c_289_n N_D_c_395_n 5.57265e-19 $X=0.735 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_284 N_A_81_194#_c_282_n N_D_M1043_g 0.0140793f $X=2.435 $Y=1.185 $X2=0 $Y2=0
cc_285 N_A_81_194#_c_288_n N_D_M1043_g 0.0205185f $X=0.57 $Y=1.135 $X2=0 $Y2=0
cc_286 N_A_81_194#_c_289_n N_D_M1043_g 0.0010579f $X=0.735 $Y=1.135 $X2=0 $Y2=0
cc_287 N_A_81_194#_c_291_n N_D_M1043_g 0.0366709f $X=0.57 $Y=0.97 $X2=0 $Y2=0
cc_288 N_A_81_194#_c_282_n D 0.00984194f $X=2.435 $Y=1.185 $X2=0 $Y2=0
cc_289 N_A_81_194#_c_288_n D 6.29362e-19 $X=0.57 $Y=1.135 $X2=0 $Y2=0
cc_290 N_A_81_194#_c_289_n D 0.0101398f $X=0.735 $Y=1.135 $X2=0 $Y2=0
cc_291 N_A_81_194#_c_282_n N_SCE_M1010_g 0.0138203f $X=2.435 $Y=1.185 $X2=0
+ $Y2=0
cc_292 N_A_81_194#_c_286_n N_SCE_c_429_n 0.00246975f $X=3.985 $Y=0.76 $X2=0
+ $Y2=0
cc_293 N_A_81_194#_c_287_n N_SCE_M1023_g 0.00434257f $X=4.14 $Y=2.075 $X2=0
+ $Y2=0
cc_294 N_A_81_194#_c_296_n N_SCE_M1023_g 0.00623049f $X=4.14 $Y=2.2 $X2=0 $Y2=0
cc_295 N_A_81_194#_c_286_n N_SCE_c_430_n 0.0119018f $X=3.985 $Y=0.76 $X2=0 $Y2=0
cc_296 N_A_81_194#_c_285_n N_SCE_c_431_n 0.0319768f $X=3.82 $Y=1.185 $X2=0 $Y2=0
cc_297 N_A_81_194#_c_286_n N_SCE_c_431_n 3.96313e-19 $X=3.985 $Y=0.76 $X2=0
+ $Y2=0
cc_298 N_A_81_194#_c_290_n N_SCE_c_431_n 0.00342124f $X=4.022 $Y=1.185 $X2=0
+ $Y2=0
cc_299 N_A_81_194#_M1030_g N_SCE_c_438_n 0.0148693f $X=2.59 $Y=2.595 $X2=0 $Y2=0
cc_300 N_A_81_194#_c_283_n N_SCE_c_438_n 0.0241538f $X=2.6 $Y=1.615 $X2=0 $Y2=0
cc_301 N_A_81_194#_c_284_n N_SCE_c_438_n 5.43058e-19 $X=2.6 $Y=1.615 $X2=0 $Y2=0
cc_302 N_A_81_194#_c_285_n N_SCE_c_432_n 0.0148377f $X=3.82 $Y=1.185 $X2=0 $Y2=0
cc_303 N_A_81_194#_c_287_n N_SCE_c_432_n 0.030569f $X=4.14 $Y=2.075 $X2=0 $Y2=0
cc_304 N_A_81_194#_c_290_n N_SCE_c_432_n 0.00264764f $X=4.022 $Y=1.185 $X2=0
+ $Y2=0
cc_305 N_A_81_194#_c_296_n N_SCE_c_432_n 0.00674102f $X=4.14 $Y=2.2 $X2=0 $Y2=0
cc_306 N_A_81_194#_c_285_n N_SCE_c_433_n 4.34101e-19 $X=3.82 $Y=1.185 $X2=0
+ $Y2=0
cc_307 N_A_81_194#_c_287_n N_SCE_c_433_n 0.00222857f $X=4.14 $Y=2.075 $X2=0
+ $Y2=0
cc_308 N_A_81_194#_c_290_n N_SCE_c_433_n 3.33761e-19 $X=4.022 $Y=1.185 $X2=0
+ $Y2=0
cc_309 N_A_81_194#_c_282_n N_SCE_c_434_n 0.00100875f $X=2.435 $Y=1.185 $X2=0
+ $Y2=0
cc_310 N_A_81_194#_c_285_n N_SCE_c_435_n 0.0041081f $X=3.82 $Y=1.185 $X2=0 $Y2=0
cc_311 N_A_81_194#_c_287_n N_SCE_c_435_n 0.0079456f $X=4.14 $Y=2.075 $X2=0 $Y2=0
cc_312 N_A_81_194#_c_282_n N_SCE_c_436_n 0.0338501f $X=2.435 $Y=1.185 $X2=0
+ $Y2=0
cc_313 N_A_81_194#_c_282_n N_SCD_M1044_g 0.0124896f $X=2.435 $Y=1.185 $X2=0
+ $Y2=0
cc_314 N_A_81_194#_c_283_n N_SCD_M1044_g 0.00542617f $X=2.6 $Y=1.615 $X2=0 $Y2=0
cc_315 N_A_81_194#_M1030_g N_SCD_M1041_g 0.0738992f $X=2.59 $Y=2.595 $X2=0 $Y2=0
cc_316 N_A_81_194#_c_282_n SCD 0.0254745f $X=2.435 $Y=1.185 $X2=0 $Y2=0
cc_317 N_A_81_194#_c_283_n SCD 0.0251565f $X=2.6 $Y=1.615 $X2=0 $Y2=0
cc_318 N_A_81_194#_c_284_n SCD 0.00187426f $X=2.6 $Y=1.615 $X2=0 $Y2=0
cc_319 N_A_81_194#_c_282_n N_SCD_c_537_n 0.0044775f $X=2.435 $Y=1.185 $X2=0
+ $Y2=0
cc_320 N_A_81_194#_c_283_n N_SCD_c_537_n 3.86757e-19 $X=2.6 $Y=1.615 $X2=0 $Y2=0
cc_321 N_A_81_194#_c_284_n N_SCD_c_537_n 0.0206812f $X=2.6 $Y=1.615 $X2=0 $Y2=0
cc_322 N_A_81_194#_c_286_n N_CLK_M1015_g 0.00172787f $X=3.985 $Y=0.76 $X2=0
+ $Y2=0
cc_323 N_A_81_194#_c_287_n N_CLK_M1031_g 0.00135815f $X=4.14 $Y=2.075 $X2=0
+ $Y2=0
cc_324 N_A_81_194#_c_286_n N_RESET_B_c_907_n 0.00729783f $X=3.985 $Y=0.76 $X2=0
+ $Y2=0
cc_325 N_A_81_194#_c_285_n N_RESET_B_c_909_n 0.0183561f $X=3.82 $Y=1.185 $X2=0
+ $Y2=0
cc_326 N_A_81_194#_c_342_p N_RESET_B_c_909_n 0.00938931f $X=2.6 $Y=1.185 $X2=0
+ $Y2=0
cc_327 N_A_81_194#_c_282_n N_RESET_B_c_910_n 0.00664891f $X=2.435 $Y=1.185 $X2=0
+ $Y2=0
cc_328 N_A_81_194#_c_284_n N_RESET_B_c_910_n 0.0214053f $X=2.6 $Y=1.615 $X2=0
+ $Y2=0
cc_329 N_A_81_194#_c_342_p N_RESET_B_c_910_n 0.00514747f $X=2.6 $Y=1.185 $X2=0
+ $Y2=0
cc_330 N_A_81_194#_M1030_g N_RESET_B_M1009_g 0.0340075f $X=2.59 $Y=2.595 $X2=0
+ $Y2=0
cc_331 N_A_81_194#_c_296_n N_RESET_B_M1009_g 8.49861e-19 $X=4.14 $Y=2.2 $X2=0
+ $Y2=0
cc_332 N_A_81_194#_c_285_n N_RESET_B_c_919_n 0.00938393f $X=3.82 $Y=1.185 $X2=0
+ $Y2=0
cc_333 N_A_81_194#_c_287_n N_RESET_B_c_919_n 0.0170861f $X=4.14 $Y=2.075 $X2=0
+ $Y2=0
cc_334 N_A_81_194#_c_290_n N_RESET_B_c_919_n 0.00856238f $X=4.022 $Y=1.185 $X2=0
+ $Y2=0
cc_335 N_A_81_194#_c_296_n N_RESET_B_c_919_n 0.00796292f $X=4.14 $Y=2.2 $X2=0
+ $Y2=0
cc_336 N_A_81_194#_c_283_n N_RESET_B_c_920_n 0.00611146f $X=2.6 $Y=1.615 $X2=0
+ $Y2=0
cc_337 N_A_81_194#_c_284_n N_RESET_B_c_920_n 0.00133803f $X=2.6 $Y=1.615 $X2=0
+ $Y2=0
cc_338 N_A_81_194#_c_285_n N_RESET_B_c_920_n 0.00163576f $X=3.82 $Y=1.185 $X2=0
+ $Y2=0
cc_339 N_A_81_194#_c_283_n N_RESET_B_c_923_n 9.61509e-19 $X=2.6 $Y=1.615 $X2=0
+ $Y2=0
cc_340 N_A_81_194#_c_284_n N_RESET_B_c_923_n 0.0212575f $X=2.6 $Y=1.615 $X2=0
+ $Y2=0
cc_341 N_A_81_194#_c_285_n N_RESET_B_c_923_n 0.00123532f $X=3.82 $Y=1.185 $X2=0
+ $Y2=0
cc_342 N_A_81_194#_c_283_n N_RESET_B_c_924_n 0.0177987f $X=2.6 $Y=1.615 $X2=0
+ $Y2=0
cc_343 N_A_81_194#_c_284_n N_RESET_B_c_924_n 0.00131162f $X=2.6 $Y=1.615 $X2=0
+ $Y2=0
cc_344 N_A_81_194#_c_285_n N_RESET_B_c_924_n 0.0213734f $X=3.82 $Y=1.185 $X2=0
+ $Y2=0
cc_345 N_A_81_194#_c_283_n N_RESET_B_c_925_n 0.00636019f $X=2.6 $Y=1.615 $X2=0
+ $Y2=0
cc_346 N_A_81_194#_c_285_n N_RESET_B_c_925_n 0.00355711f $X=3.82 $Y=1.185 $X2=0
+ $Y2=0
cc_347 N_A_81_194#_c_286_n N_A_876_119#_c_1292_n 0.0334652f $X=3.985 $Y=0.76
+ $X2=0 $Y2=0
cc_348 N_A_81_194#_c_287_n N_A_876_119#_c_1292_n 0.0273932f $X=4.14 $Y=2.075
+ $X2=0 $Y2=0
cc_349 N_A_81_194#_c_290_n N_A_876_119#_c_1292_n 0.0130308f $X=4.022 $Y=1.185
+ $X2=0 $Y2=0
cc_350 N_A_81_194#_c_287_n N_A_876_119#_c_1308_n 0.0158131f $X=4.14 $Y=2.075
+ $X2=0 $Y2=0
cc_351 N_A_81_194#_c_296_n N_A_876_119#_c_1308_n 0.0186811f $X=4.14 $Y=2.2 $X2=0
+ $Y2=0
cc_352 N_A_81_194#_c_287_n N_A_876_119#_c_1311_n 0.0122953f $X=4.14 $Y=2.075
+ $X2=0 $Y2=0
cc_353 N_A_81_194#_M1030_g N_A_116_419#_c_1805_n 0.0146029f $X=2.59 $Y=2.595
+ $X2=0 $Y2=0
cc_354 N_A_81_194#_c_296_n N_A_116_419#_c_1806_n 0.00180442f $X=4.14 $Y=2.2
+ $X2=0 $Y2=0
cc_355 N_A_81_194#_M1023_d N_A_116_419#_c_1799_n 0.00758169f $X=3.86 $Y=2.095
+ $X2=0 $Y2=0
cc_356 N_A_81_194#_c_296_n N_A_116_419#_c_1799_n 0.00958463f $X=4.14 $Y=2.2
+ $X2=0 $Y2=0
cc_357 N_A_81_194#_c_288_n N_A_116_419#_c_1796_n 0.00768695f $X=0.57 $Y=1.135
+ $X2=0 $Y2=0
cc_358 N_A_81_194#_c_289_n N_A_116_419#_c_1796_n 0.0243373f $X=0.735 $Y=1.135
+ $X2=0 $Y2=0
cc_359 N_A_81_194#_c_291_n N_A_116_419#_c_1796_n 0.00536188f $X=0.57 $Y=0.97
+ $X2=0 $Y2=0
cc_360 N_A_81_194#_c_282_n N_A_116_419#_c_1797_n 0.0199718f $X=2.435 $Y=1.185
+ $X2=0 $Y2=0
cc_361 N_A_81_194#_c_282_n N_A_116_419#_c_1813_n 0.0157849f $X=2.435 $Y=1.185
+ $X2=0 $Y2=0
cc_362 N_A_81_194#_c_288_n N_A_116_419#_c_1813_n 0.00373328f $X=0.57 $Y=1.135
+ $X2=0 $Y2=0
cc_363 N_A_81_194#_c_289_n N_A_116_419#_c_1813_n 0.0174476f $X=0.735 $Y=1.135
+ $X2=0 $Y2=0
cc_364 N_A_81_194#_c_291_n N_A_116_419#_c_1813_n 0.0120414f $X=0.57 $Y=0.97
+ $X2=0 $Y2=0
cc_365 N_A_81_194#_M1030_g N_A_116_419#_c_1817_n 0.00516659f $X=2.59 $Y=2.595
+ $X2=0 $Y2=0
cc_366 N_A_81_194#_M1030_g N_A_116_419#_c_1818_n 0.00837674f $X=2.59 $Y=2.595
+ $X2=0 $Y2=0
cc_367 N_A_81_194#_M1030_g N_VPWR_c_1935_n 9.35833e-19 $X=2.59 $Y=2.595 $X2=0
+ $Y2=0
cc_368 N_A_81_194#_M1030_g N_VPWR_c_1943_n 0.00939541f $X=2.59 $Y=2.595 $X2=0
+ $Y2=0
cc_369 N_A_81_194#_M1023_d N_VPWR_c_1933_n 0.00233017f $X=3.86 $Y=2.095 $X2=0
+ $Y2=0
cc_370 N_A_81_194#_M1030_g N_VPWR_c_1933_n 0.00955495f $X=2.59 $Y=2.595 $X2=0
+ $Y2=0
cc_371 N_A_81_194#_c_282_n N_noxref_23_c_2134_n 0.0145246f $X=2.435 $Y=1.185
+ $X2=0 $Y2=0
cc_372 N_A_81_194#_c_291_n N_noxref_23_c_2134_n 0.0100323f $X=0.57 $Y=0.97 $X2=0
+ $Y2=0
cc_373 N_A_81_194#_c_282_n N_noxref_23_c_2135_n 0.0225098f $X=2.435 $Y=1.185
+ $X2=0 $Y2=0
cc_374 N_A_81_194#_c_285_n N_VGND_c_2163_n 0.00799885f $X=3.82 $Y=1.185 $X2=0
+ $Y2=0
cc_375 N_A_81_194#_c_342_p N_VGND_c_2163_n 0.0146295f $X=2.6 $Y=1.185 $X2=0
+ $Y2=0
cc_376 N_A_81_194#_c_291_n N_VGND_c_2169_n 8.40037e-19 $X=0.57 $Y=0.97 $X2=0
+ $Y2=0
cc_377 N_A_81_194#_c_286_n N_VGND_c_2170_n 0.00797279f $X=3.985 $Y=0.76 $X2=0
+ $Y2=0
cc_378 N_A_81_194#_c_286_n N_VGND_c_2174_n 0.010956f $X=3.985 $Y=0.76 $X2=0
+ $Y2=0
cc_379 N_D_M1043_g N_SCE_M1010_g 0.0367658f $X=1.02 $Y=0.65 $X2=0 $Y2=0
cc_380 N_D_c_395_n N_SCE_c_434_n 0.0853247f $X=0.99 $Y=2.025 $X2=0 $Y2=0
cc_381 N_D_c_395_n N_SCE_c_436_n 0.0199402f $X=0.99 $Y=2.025 $X2=0 $Y2=0
cc_382 D N_SCE_c_436_n 0.0226408f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_383 N_D_c_395_n N_A_116_419#_c_1805_n 0.0185499f $X=0.99 $Y=2.025 $X2=0 $Y2=0
cc_384 D N_A_116_419#_c_1805_n 4.68986e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_385 N_D_c_395_n N_A_116_419#_c_1803_n 0.0322922f $X=0.99 $Y=2.025 $X2=0 $Y2=0
cc_386 D N_A_116_419#_c_1803_n 0.020679f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_387 N_D_c_395_n N_A_116_419#_c_1796_n 0.00735158f $X=0.99 $Y=2.025 $X2=0
+ $Y2=0
cc_388 N_D_M1043_g N_A_116_419#_c_1796_n 0.00422472f $X=1.02 $Y=0.65 $X2=0 $Y2=0
cc_389 D N_A_116_419#_c_1796_n 0.0156061f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_390 N_D_M1043_g N_A_116_419#_c_1797_n 5.27414e-19 $X=1.02 $Y=0.65 $X2=0 $Y2=0
cc_391 N_D_M1043_g N_A_116_419#_c_1813_n 0.0115302f $X=1.02 $Y=0.65 $X2=0 $Y2=0
cc_392 N_D_c_395_n N_VPWR_c_1934_n 0.00278628f $X=0.99 $Y=2.025 $X2=0 $Y2=0
cc_393 N_D_c_395_n N_VPWR_c_1949_n 0.00939541f $X=0.99 $Y=2.025 $X2=0 $Y2=0
cc_394 N_D_c_395_n N_VPWR_c_1933_n 0.0107661f $X=0.99 $Y=2.025 $X2=0 $Y2=0
cc_395 N_D_M1043_g N_noxref_23_c_2134_n 0.00940864f $X=1.02 $Y=0.65 $X2=0 $Y2=0
cc_396 N_D_M1043_g N_VGND_c_2169_n 8.40037e-19 $X=1.02 $Y=0.65 $X2=0 $Y2=0
cc_397 N_SCE_M1010_g N_SCD_M1044_g 0.0621785f $X=1.61 $Y=0.65 $X2=0 $Y2=0
cc_398 N_SCE_c_438_n N_SCD_M1041_g 0.0150668f $X=3.485 $Y=2.045 $X2=0 $Y2=0
cc_399 N_SCE_c_434_n N_SCD_M1041_g 0.0114963f $X=1.52 $Y=1.77 $X2=0 $Y2=0
cc_400 N_SCE_c_442_n N_SCD_M1041_g 0.0383871f $X=1.52 $Y=2.02 $X2=0 $Y2=0
cc_401 N_SCE_c_436_n N_SCD_M1041_g 0.0011946f $X=1.685 $Y=1.84 $X2=0 $Y2=0
cc_402 N_SCE_M1010_g SCD 9.55563e-19 $X=1.61 $Y=0.65 $X2=0 $Y2=0
cc_403 N_SCE_c_438_n SCD 0.025097f $X=3.485 $Y=2.045 $X2=0 $Y2=0
cc_404 N_SCE_c_436_n SCD 0.0153295f $X=1.685 $Y=1.84 $X2=0 $Y2=0
cc_405 N_SCE_M1010_g N_SCD_c_537_n 0.0208354f $X=1.61 $Y=0.65 $X2=0 $Y2=0
cc_406 N_SCE_c_438_n N_SCD_c_537_n 0.00186008f $X=3.485 $Y=2.045 $X2=0 $Y2=0
cc_407 N_SCE_c_436_n N_SCD_c_537_n 2.85665e-19 $X=1.685 $Y=1.84 $X2=0 $Y2=0
cc_408 N_SCE_c_429_n N_RESET_B_c_907_n 0.0104164f $X=3.41 $Y=1.09 $X2=0 $Y2=0
cc_409 N_SCE_c_430_n N_RESET_B_c_907_n 0.0103053f $X=3.77 $Y=1.09 $X2=0 $Y2=0
cc_410 N_SCE_c_431_n N_RESET_B_c_909_n 0.00994981f $X=3.77 $Y=1.165 $X2=0 $Y2=0
cc_411 N_SCE_M1023_g N_RESET_B_M1009_g 0.0392414f $X=3.735 $Y=2.595 $X2=0 $Y2=0
cc_412 N_SCE_c_438_n N_RESET_B_M1009_g 0.0168289f $X=3.485 $Y=2.045 $X2=0 $Y2=0
cc_413 N_SCE_c_432_n N_RESET_B_M1009_g 0.00393489f $X=3.71 $Y=1.72 $X2=0 $Y2=0
cc_414 N_SCE_c_433_n N_RESET_B_M1009_g 0.00408267f $X=3.71 $Y=1.72 $X2=0 $Y2=0
cc_415 N_SCE_c_438_n N_RESET_B_c_919_n 0.00587278f $X=3.485 $Y=2.045 $X2=0 $Y2=0
cc_416 N_SCE_c_432_n N_RESET_B_c_919_n 0.0307238f $X=3.71 $Y=1.72 $X2=0 $Y2=0
cc_417 N_SCE_c_433_n N_RESET_B_c_919_n 0.00229642f $X=3.71 $Y=1.72 $X2=0 $Y2=0
cc_418 N_SCE_c_438_n N_RESET_B_c_920_n 0.00206906f $X=3.485 $Y=2.045 $X2=0 $Y2=0
cc_419 N_SCE_c_432_n N_RESET_B_c_920_n 6.1553e-19 $X=3.71 $Y=1.72 $X2=0 $Y2=0
cc_420 N_SCE_c_438_n N_RESET_B_c_923_n 5.41421e-19 $X=3.485 $Y=2.045 $X2=0 $Y2=0
cc_421 N_SCE_c_432_n N_RESET_B_c_923_n 0.00114638f $X=3.71 $Y=1.72 $X2=0 $Y2=0
cc_422 N_SCE_c_435_n N_RESET_B_c_923_n 0.0184561f $X=3.71 $Y=1.555 $X2=0 $Y2=0
cc_423 N_SCE_c_438_n N_RESET_B_c_924_n 0.0190838f $X=3.485 $Y=2.045 $X2=0 $Y2=0
cc_424 N_SCE_c_432_n N_RESET_B_c_924_n 0.0150387f $X=3.71 $Y=1.72 $X2=0 $Y2=0
cc_425 N_SCE_c_433_n N_RESET_B_c_924_n 3.3415e-19 $X=3.71 $Y=1.72 $X2=0 $Y2=0
cc_426 N_SCE_c_435_n N_RESET_B_c_924_n 6.77823e-19 $X=3.71 $Y=1.555 $X2=0 $Y2=0
cc_427 N_SCE_c_435_n N_RESET_B_c_925_n 0.00706832f $X=3.71 $Y=1.555 $X2=0 $Y2=0
cc_428 N_SCE_c_430_n N_A_876_119#_c_1292_n 0.00130723f $X=3.77 $Y=1.09 $X2=0
+ $Y2=0
cc_429 N_SCE_M1023_g N_A_876_119#_c_1308_n 0.00494543f $X=3.735 $Y=2.595 $X2=0
+ $Y2=0
cc_430 N_SCE_c_438_n N_A_116_419#_M1030_d 0.00180746f $X=3.485 $Y=2.045 $X2=0
+ $Y2=0
cc_431 N_SCE_c_434_n N_A_116_419#_c_1805_n 3.14702e-19 $X=1.52 $Y=1.77 $X2=0
+ $Y2=0
cc_432 N_SCE_c_442_n N_A_116_419#_c_1805_n 0.0173299f $X=1.52 $Y=2.02 $X2=0
+ $Y2=0
cc_433 N_SCE_c_436_n N_A_116_419#_c_1805_n 0.0875205f $X=1.685 $Y=1.84 $X2=0
+ $Y2=0
cc_434 N_SCE_M1023_g N_A_116_419#_c_1806_n 0.0181429f $X=3.735 $Y=2.595 $X2=0
+ $Y2=0
cc_435 N_SCE_c_438_n N_A_116_419#_c_1806_n 0.0157124f $X=3.485 $Y=2.045 $X2=0
+ $Y2=0
cc_436 N_SCE_c_432_n N_A_116_419#_c_1806_n 0.00946858f $X=3.71 $Y=1.72 $X2=0
+ $Y2=0
cc_437 N_SCE_M1023_g N_A_116_419#_c_1835_n 0.00904063f $X=3.735 $Y=2.595 $X2=0
+ $Y2=0
cc_438 N_SCE_M1023_g N_A_116_419#_c_1836_n 0.00878851f $X=3.735 $Y=2.595 $X2=0
+ $Y2=0
cc_439 N_SCE_c_442_n N_A_116_419#_c_1803_n 0.00337233f $X=1.52 $Y=2.02 $X2=0
+ $Y2=0
cc_440 N_SCE_c_436_n N_A_116_419#_c_1803_n 0.0040735f $X=1.685 $Y=1.84 $X2=0
+ $Y2=0
cc_441 N_SCE_M1010_g N_A_116_419#_c_1797_n 0.00156413f $X=1.61 $Y=0.65 $X2=0
+ $Y2=0
cc_442 N_SCE_M1023_g N_A_116_419#_c_1817_n 0.00169376f $X=3.735 $Y=2.595 $X2=0
+ $Y2=0
cc_443 N_SCE_c_438_n N_A_116_419#_c_1817_n 0.0162839f $X=3.485 $Y=2.045 $X2=0
+ $Y2=0
cc_444 N_SCE_c_436_n A_223_419# 0.0014282f $X=1.685 $Y=1.84 $X2=-0.19 $Y2=-0.245
cc_445 N_SCE_c_438_n N_VPWR_M1018_d 0.00222802f $X=3.485 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_446 N_SCE_c_436_n N_VPWR_M1018_d 2.60703e-19 $X=1.685 $Y=1.84 $X2=-0.19
+ $Y2=-0.245
cc_447 N_SCE_c_438_n N_VPWR_M1009_d 0.00285834f $X=3.485 $Y=2.045 $X2=0 $Y2=0
cc_448 N_SCE_c_432_n N_VPWR_M1009_d 0.00109639f $X=3.71 $Y=1.72 $X2=0 $Y2=0
cc_449 N_SCE_c_442_n N_VPWR_c_1934_n 0.0144383f $X=1.52 $Y=2.02 $X2=0 $Y2=0
cc_450 N_SCE_M1023_g N_VPWR_c_1935_n 0.00570242f $X=3.735 $Y=2.595 $X2=0 $Y2=0
cc_451 N_SCE_M1023_g N_VPWR_c_1945_n 0.00654206f $X=3.735 $Y=2.595 $X2=0 $Y2=0
cc_452 N_SCE_c_442_n N_VPWR_c_1949_n 0.008763f $X=1.52 $Y=2.02 $X2=0 $Y2=0
cc_453 N_SCE_M1023_g N_VPWR_c_1933_n 0.00997498f $X=3.735 $Y=2.595 $X2=0 $Y2=0
cc_454 N_SCE_c_442_n N_VPWR_c_1933_n 0.00779322f $X=1.52 $Y=2.02 $X2=0 $Y2=0
cc_455 N_SCE_c_438_n A_439_419# 0.00170258f $X=3.485 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_456 N_SCE_M1010_g N_noxref_23_c_2134_n 0.0115792f $X=1.61 $Y=0.65 $X2=0 $Y2=0
cc_457 N_SCE_M1010_g N_noxref_23_c_2135_n 0.00170236f $X=1.61 $Y=0.65 $X2=0
+ $Y2=0
cc_458 N_SCE_c_429_n N_VGND_c_2163_n 0.0115205f $X=3.41 $Y=1.09 $X2=0 $Y2=0
cc_459 N_SCE_M1010_g N_VGND_c_2169_n 8.40037e-19 $X=1.61 $Y=0.65 $X2=0 $Y2=0
cc_460 N_SCE_c_429_n N_VGND_c_2174_n 9.39239e-19 $X=3.41 $Y=1.09 $X2=0 $Y2=0
cc_461 N_SCE_c_430_n N_VGND_c_2174_n 9.39239e-19 $X=3.77 $Y=1.09 $X2=0 $Y2=0
cc_462 N_SCD_M1044_g N_RESET_B_M1011_g 0.0263076f $X=2 $Y=0.65 $X2=0 $Y2=0
cc_463 N_SCD_M1041_g N_A_116_419#_c_1805_n 0.0177671f $X=2.07 $Y=2.595 $X2=0
+ $Y2=0
cc_464 N_SCD_M1041_g N_A_116_419#_c_1817_n 0.00258079f $X=2.07 $Y=2.595 $X2=0
+ $Y2=0
cc_465 N_SCD_M1041_g N_VPWR_c_1934_n 0.00568123f $X=2.07 $Y=2.595 $X2=0 $Y2=0
cc_466 N_SCD_M1041_g N_VPWR_c_1943_n 0.00975641f $X=2.07 $Y=2.595 $X2=0 $Y2=0
cc_467 N_SCD_M1041_g N_VPWR_c_1933_n 0.00980097f $X=2.07 $Y=2.595 $X2=0 $Y2=0
cc_468 N_SCD_M1044_g N_noxref_23_c_2134_n 0.0102473f $X=2 $Y=0.65 $X2=0 $Y2=0
cc_469 N_SCD_M1044_g N_noxref_23_c_2135_n 0.00889413f $X=2 $Y=0.65 $X2=0 $Y2=0
cc_470 N_SCD_M1044_g N_VGND_c_2169_n 8.58586e-19 $X=2 $Y=0.65 $X2=0 $Y2=0
cc_471 N_CLK_M1015_g N_RESET_B_c_907_n 0.0104164f $X=4.72 $Y=0.805 $X2=0 $Y2=0
cc_472 N_CLK_M1032_g N_RESET_B_c_907_n 0.0104164f $X=5.08 $Y=0.805 $X2=0 $Y2=0
cc_473 N_CLK_M1031_g N_RESET_B_c_919_n 0.00755498f $X=4.85 $Y=2.54 $X2=0 $Y2=0
cc_474 CLK N_RESET_B_c_919_n 0.0085402f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_475 N_CLK_c_574_n N_RESET_B_c_919_n 0.00733657f $X=4.99 $Y=1.335 $X2=0 $Y2=0
cc_476 N_CLK_M1031_g N_A_876_119#_M1016_g 0.0297121f $X=4.85 $Y=2.54 $X2=0 $Y2=0
cc_477 N_CLK_M1032_g N_A_876_119#_M1029_g 0.0198053f $X=5.08 $Y=0.805 $X2=0
+ $Y2=0
cc_478 N_CLK_M1015_g N_A_876_119#_c_1292_n 0.0106352f $X=4.72 $Y=0.805 $X2=0
+ $Y2=0
cc_479 CLK N_A_876_119#_c_1292_n 0.0194104f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_480 N_CLK_c_574_n N_A_876_119#_c_1292_n 0.0106775f $X=4.99 $Y=1.335 $X2=0
+ $Y2=0
cc_481 N_CLK_M1031_g N_A_876_119#_c_1308_n 0.00812807f $X=4.85 $Y=2.54 $X2=0
+ $Y2=0
cc_482 N_CLK_M1031_g N_A_876_119#_c_1309_n 0.022733f $X=4.85 $Y=2.54 $X2=0 $Y2=0
cc_483 CLK N_A_876_119#_c_1309_n 0.0196459f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_484 N_CLK_c_574_n N_A_876_119#_c_1309_n 0.00623556f $X=4.99 $Y=1.335 $X2=0
+ $Y2=0
cc_485 N_CLK_M1031_g N_A_876_119#_c_1293_n 0.00116002f $X=4.85 $Y=2.54 $X2=0
+ $Y2=0
cc_486 CLK N_A_876_119#_c_1293_n 0.0144711f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_487 N_CLK_c_574_n N_A_876_119#_c_1293_n 4.06458e-19 $X=4.99 $Y=1.335 $X2=0
+ $Y2=0
cc_488 N_CLK_M1031_g N_A_876_119#_c_1294_n 0.00827865f $X=4.85 $Y=2.54 $X2=0
+ $Y2=0
cc_489 CLK N_A_876_119#_c_1294_n 0.00150202f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_490 N_CLK_c_574_n N_A_876_119#_c_1294_n 0.0126879f $X=4.99 $Y=1.335 $X2=0
+ $Y2=0
cc_491 N_CLK_c_574_n N_A_876_119#_c_1311_n 7.86615e-19 $X=4.99 $Y=1.335 $X2=0
+ $Y2=0
cc_492 N_CLK_M1031_g N_A_116_419#_c_1799_n 0.0164635f $X=4.85 $Y=2.54 $X2=0
+ $Y2=0
cc_493 N_CLK_M1031_g N_A_116_419#_c_1845_n 0.0130064f $X=4.85 $Y=2.54 $X2=0
+ $Y2=0
cc_494 N_CLK_M1031_g N_A_116_419#_c_1846_n 0.0105353f $X=4.85 $Y=2.54 $X2=0
+ $Y2=0
cc_495 N_CLK_M1031_g N_VPWR_c_1936_n 0.00302821f $X=4.85 $Y=2.54 $X2=0 $Y2=0
cc_496 N_CLK_M1031_g N_VPWR_c_1945_n 0.00540963f $X=4.85 $Y=2.54 $X2=0 $Y2=0
cc_497 N_CLK_M1031_g N_VPWR_c_1933_n 0.00851682f $X=4.85 $Y=2.54 $X2=0 $Y2=0
cc_498 N_CLK_M1032_g N_VGND_c_2164_n 0.00456171f $X=5.08 $Y=0.805 $X2=0 $Y2=0
cc_499 N_CLK_M1015_g N_VGND_c_2174_n 9.39239e-19 $X=4.72 $Y=0.805 $X2=0 $Y2=0
cc_500 N_CLK_M1032_g N_VGND_c_2174_n 9.39239e-19 $X=5.08 $Y=0.805 $X2=0 $Y2=0
cc_501 N_A_1147_408#_c_618_n N_A_1605_93#_M1033_d 0.00358346f $X=10.21 $Y=0.71
+ $X2=-0.19 $Y2=-0.245
cc_502 N_A_1147_408#_c_609_n N_A_1605_93#_c_782_n 0.0281901f $X=7.73 $Y=1.125
+ $X2=0 $Y2=0
cc_503 N_A_1147_408#_c_616_n N_A_1605_93#_c_782_n 0.00250176f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_504 N_A_1147_408#_c_618_n N_A_1605_93#_c_782_n 0.0154524f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_505 N_A_1147_408#_c_616_n N_A_1605_93#_c_783_n 2.11641e-19 $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_506 N_A_1147_408#_c_617_n N_A_1605_93#_c_783_n 0.00275755f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_507 N_A_1147_408#_c_616_n N_A_1605_93#_c_784_n 0.0120448f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_508 N_A_1147_408#_c_617_n N_A_1605_93#_c_784_n 0.00152395f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_509 N_A_1147_408#_c_617_n N_A_1605_93#_c_785_n 0.0294077f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_510 N_A_1147_408#_c_618_n N_A_1605_93#_c_785_n 0.00171882f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_511 N_A_1147_408#_c_618_n N_A_1605_93#_c_786_n 0.0894065f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_512 N_A_1147_408#_c_616_n N_A_1605_93#_c_787_n 0.00510669f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_513 N_A_1147_408#_c_618_n N_A_1605_93#_c_787_n 0.0247499f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_514 N_A_1147_408#_c_610_n N_A_1605_93#_c_812_n 0.0040575f $X=11.455 $Y=0.805
+ $X2=0 $Y2=0
cc_515 N_A_1147_408#_c_618_n N_A_1605_93#_c_812_n 0.0239771f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_516 N_A_1147_408#_c_622_n N_A_1605_93#_c_812_n 8.73282e-19 $X=10.295 $Y=0.805
+ $X2=0 $Y2=0
cc_517 N_A_1147_408#_c_623_n N_A_1605_93#_c_812_n 0.01028f $X=10.295 $Y=0.73
+ $X2=0 $Y2=0
cc_518 N_A_1147_408#_c_610_n N_A_1605_93#_c_788_n 9.5475e-19 $X=11.455 $Y=0.805
+ $X2=0 $Y2=0
cc_519 N_A_1147_408#_c_618_n N_A_1605_93#_c_788_n 0.00591696f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_520 N_A_1147_408#_c_619_n N_A_1605_93#_c_788_n 0.0151732f $X=10.295 $Y=0.93
+ $X2=0 $Y2=0
cc_521 N_A_1147_408#_c_622_n N_A_1605_93#_c_788_n 0.00234018f $X=10.295 $Y=0.805
+ $X2=0 $Y2=0
cc_522 N_A_1147_408#_c_610_n N_A_1605_93#_c_789_n 0.0186998f $X=11.455 $Y=0.805
+ $X2=0 $Y2=0
cc_523 N_A_1147_408#_c_611_n N_A_1605_93#_c_789_n 0.00485188f $X=11.53 $Y=1.48
+ $X2=0 $Y2=0
cc_524 N_A_1147_408#_c_618_n N_A_1605_93#_c_789_n 0.0126816f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_525 N_A_1147_408#_c_619_n N_A_1605_93#_c_789_n 0.0205576f $X=10.295 $Y=0.93
+ $X2=0 $Y2=0
cc_526 N_A_1147_408#_c_622_n N_A_1605_93#_c_789_n 0.00499077f $X=10.295 $Y=0.805
+ $X2=0 $Y2=0
cc_527 N_A_1147_408#_c_623_n N_A_1605_93#_c_789_n 0.00837337f $X=10.295 $Y=0.73
+ $X2=0 $Y2=0
cc_528 N_A_1147_408#_c_618_n N_A_1605_93#_c_790_n 0.0130644f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_529 N_A_1147_408#_c_619_n N_A_1605_93#_c_790_n 0.00873157f $X=10.295 $Y=0.93
+ $X2=0 $Y2=0
cc_530 N_A_1147_408#_c_622_n N_A_1605_93#_c_790_n 8.00088e-19 $X=10.295 $Y=0.805
+ $X2=0 $Y2=0
cc_531 N_A_1147_408#_c_609_n N_RESET_B_c_907_n 0.00976871f $X=7.73 $Y=1.125
+ $X2=0 $Y2=0
cc_532 N_A_1147_408#_c_615_n N_RESET_B_c_907_n 0.0067384f $X=6.245 $Y=0.79 $X2=0
+ $Y2=0
cc_533 N_A_1147_408#_c_618_n N_RESET_B_c_907_n 0.0106121f $X=10.21 $Y=0.71 $X2=0
+ $Y2=0
cc_534 N_A_1147_408#_c_667_p N_RESET_B_c_907_n 0.00180368f $X=7.725 $Y=0.71
+ $X2=0 $Y2=0
cc_535 N_A_1147_408#_c_618_n N_RESET_B_M1021_g 0.0131738f $X=10.21 $Y=0.71 $X2=0
+ $Y2=0
cc_536 N_A_1147_408#_c_618_n N_RESET_B_c_915_n 0.0104845f $X=10.21 $Y=0.71 $X2=0
+ $Y2=0
cc_537 N_A_1147_408#_c_608_n N_RESET_B_c_919_n 0.00776635f $X=7.235 $Y=1.555
+ $X2=0 $Y2=0
cc_538 N_A_1147_408#_c_625_n N_RESET_B_c_919_n 0.00146278f $X=7.36 $Y=1.66 $X2=0
+ $Y2=0
cc_539 N_A_1147_408#_c_630_n N_RESET_B_c_919_n 0.0106121f $X=6.132 $Y=2.03 $X2=0
+ $Y2=0
cc_540 N_A_1147_408#_c_615_n N_RESET_B_c_919_n 0.00210741f $X=6.245 $Y=0.79
+ $X2=0 $Y2=0
cc_541 N_A_1147_408#_c_616_n N_RESET_B_c_919_n 0.00463772f $X=7.64 $Y=1.29 $X2=0
+ $Y2=0
cc_542 N_A_1147_408#_c_617_n N_RESET_B_c_919_n 0.0129086f $X=7.64 $Y=1.29 $X2=0
+ $Y2=0
cc_543 N_A_1147_408#_c_620_n N_RESET_B_c_919_n 0.047476f $X=6.6 $Y=1.615 $X2=0
+ $Y2=0
cc_544 N_A_1147_408#_c_621_n N_RESET_B_c_919_n 0.00452378f $X=6.6 $Y=1.555 $X2=0
+ $Y2=0
cc_545 N_A_1147_408#_c_612_n N_RESET_B_c_921_n 0.00352772f $X=11.785 $Y=1.555
+ $X2=0 $Y2=0
cc_546 N_A_1147_408#_c_613_n N_RESET_B_c_921_n 0.0029583f $X=11.605 $Y=1.555
+ $X2=0 $Y2=0
cc_547 N_A_1147_408#_c_614_n N_RESET_B_c_921_n 8.59317e-19 $X=11.81 $Y=1.87
+ $X2=0 $Y2=0
cc_548 N_A_1147_408#_c_616_n N_A_1432_119#_M1014_d 0.00199971f $X=7.64 $Y=1.29
+ $X2=-0.19 $Y2=-0.245
cc_549 N_A_1147_408#_c_667_p N_A_1432_119#_M1014_d 0.00222905f $X=7.725 $Y=0.71
+ $X2=-0.19 $Y2=-0.245
cc_550 N_A_1147_408#_c_618_n N_A_1432_119#_c_1173_n 0.0153622f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_551 N_A_1147_408#_c_623_n N_A_1432_119#_c_1173_n 0.0135159f $X=10.295 $Y=0.73
+ $X2=0 $Y2=0
cc_552 N_A_1147_408#_c_610_n N_A_1432_119#_c_1174_n 0.0013899f $X=11.455
+ $Y=0.805 $X2=0 $Y2=0
cc_553 N_A_1147_408#_c_618_n N_A_1432_119#_c_1174_n 8.78044e-19 $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_554 N_A_1147_408#_c_619_n N_A_1432_119#_c_1174_n 2.15014e-19 $X=10.295
+ $Y=0.93 $X2=0 $Y2=0
cc_555 N_A_1147_408#_c_622_n N_A_1432_119#_c_1174_n 0.0119049f $X=10.295
+ $Y=0.805 $X2=0 $Y2=0
cc_556 N_A_1147_408#_c_618_n N_A_1432_119#_c_1176_n 0.0135928f $X=10.21 $Y=0.71
+ $X2=0 $Y2=0
cc_557 N_A_1147_408#_c_619_n N_A_1432_119#_c_1176_n 0.0011094f $X=10.295 $Y=0.93
+ $X2=0 $Y2=0
cc_558 N_A_1147_408#_c_622_n N_A_1432_119#_c_1176_n 0.0213132f $X=10.295
+ $Y=0.805 $X2=0 $Y2=0
cc_559 N_A_1147_408#_c_608_n N_A_1432_119#_c_1177_n 0.00378253f $X=7.235
+ $Y=1.555 $X2=0 $Y2=0
cc_560 N_A_1147_408#_c_625_n N_A_1432_119#_c_1177_n 0.00505758f $X=7.36 $Y=1.66
+ $X2=0 $Y2=0
cc_561 N_A_1147_408#_c_609_n N_A_1432_119#_c_1177_n 0.00145899f $X=7.73 $Y=1.125
+ $X2=0 $Y2=0
cc_562 N_A_1147_408#_c_616_n N_A_1432_119#_c_1177_n 0.051337f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_563 N_A_1147_408#_c_617_n N_A_1432_119#_c_1177_n 0.0210113f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_564 N_A_1147_408#_c_667_p N_A_1432_119#_c_1177_n 0.0138308f $X=7.725 $Y=0.71
+ $X2=0 $Y2=0
cc_565 N_A_1147_408#_c_625_n N_A_1432_119#_c_1183_n 0.0270504f $X=7.36 $Y=1.66
+ $X2=0 $Y2=0
cc_566 N_A_1147_408#_c_617_n N_A_1432_119#_c_1205_n 4.22339e-19 $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_567 N_A_1147_408#_c_625_n N_A_1432_119#_c_1206_n 0.0144203f $X=7.36 $Y=1.66
+ $X2=0 $Y2=0
cc_568 N_A_1147_408#_c_616_n N_A_1432_119#_c_1206_n 0.00656632f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_569 N_A_1147_408#_c_617_n N_A_1432_119#_c_1206_n 0.00742636f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_570 N_A_1147_408#_c_630_n N_A_876_119#_M1016_g 0.0166241f $X=6.132 $Y=2.03
+ $X2=0 $Y2=0
cc_571 N_A_1147_408#_c_615_n N_A_876_119#_c_1286_n 0.0116165f $X=6.245 $Y=0.79
+ $X2=0 $Y2=0
cc_572 N_A_1147_408#_c_615_n N_A_876_119#_M1029_g 0.0026942f $X=6.245 $Y=0.79
+ $X2=0 $Y2=0
cc_573 N_A_1147_408#_c_630_n N_A_876_119#_c_1300_n 0.0204846f $X=6.132 $Y=2.03
+ $X2=0 $Y2=0
cc_574 N_A_1147_408#_c_615_n N_A_876_119#_c_1288_n 0.0155439f $X=6.245 $Y=0.79
+ $X2=0 $Y2=0
cc_575 N_A_1147_408#_c_617_n N_A_876_119#_c_1288_n 0.00753185f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_576 N_A_1147_408#_c_620_n N_A_876_119#_c_1288_n 0.00246937f $X=6.6 $Y=1.615
+ $X2=0 $Y2=0
cc_577 N_A_1147_408#_c_621_n N_A_876_119#_c_1288_n 0.0477272f $X=6.6 $Y=1.555
+ $X2=0 $Y2=0
cc_578 N_A_1147_408#_c_625_n N_A_876_119#_c_1301_n 0.0161517f $X=7.36 $Y=1.66
+ $X2=0 $Y2=0
cc_579 N_A_1147_408#_c_609_n N_A_876_119#_c_1289_n 0.0102011f $X=7.73 $Y=1.125
+ $X2=0 $Y2=0
cc_580 N_A_1147_408#_c_615_n N_A_876_119#_c_1289_n 0.00114996f $X=6.245 $Y=0.79
+ $X2=0 $Y2=0
cc_581 N_A_1147_408#_c_625_n N_A_876_119#_M1042_g 0.0175126f $X=7.36 $Y=1.66
+ $X2=0 $Y2=0
cc_582 N_A_1147_408#_c_617_n N_A_876_119#_M1042_g 0.00393108f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_583 N_A_1147_408#_c_613_n N_A_876_119#_M1002_g 0.0170607f $X=11.605 $Y=1.555
+ $X2=0 $Y2=0
cc_584 N_A_1147_408#_c_628_n N_A_876_119#_M1002_g 0.0278133f $X=11.81 $Y=1.995
+ $X2=0 $Y2=0
cc_585 N_A_1147_408#_c_614_n N_A_876_119#_M1002_g 0.00425181f $X=11.81 $Y=1.87
+ $X2=0 $Y2=0
cc_586 N_A_1147_408#_c_610_n N_A_876_119#_M1020_g 0.0111154f $X=11.455 $Y=0.805
+ $X2=0 $Y2=0
cc_587 N_A_1147_408#_c_630_n N_A_876_119#_c_1309_n 0.0123929f $X=6.132 $Y=2.03
+ $X2=0 $Y2=0
cc_588 N_A_1147_408#_c_620_n N_A_876_119#_c_1309_n 0.00739608f $X=6.6 $Y=1.615
+ $X2=0 $Y2=0
cc_589 N_A_1147_408#_c_615_n N_A_876_119#_c_1293_n 0.0143815f $X=6.245 $Y=0.79
+ $X2=0 $Y2=0
cc_590 N_A_1147_408#_c_620_n N_A_876_119#_c_1293_n 0.0171028f $X=6.6 $Y=1.615
+ $X2=0 $Y2=0
cc_591 N_A_1147_408#_c_630_n N_A_876_119#_c_1294_n 0.0110803f $X=6.132 $Y=2.03
+ $X2=0 $Y2=0
cc_592 N_A_1147_408#_c_615_n N_A_876_119#_c_1294_n 0.0148735f $X=6.245 $Y=0.79
+ $X2=0 $Y2=0
cc_593 N_A_1147_408#_c_620_n N_A_876_119#_c_1294_n 0.0203577f $X=6.6 $Y=1.615
+ $X2=0 $Y2=0
cc_594 N_A_1147_408#_c_621_n N_A_876_119#_c_1294_n 0.0215857f $X=6.6 $Y=1.555
+ $X2=0 $Y2=0
cc_595 N_A_1147_408#_c_610_n N_A_876_119#_c_1295_n 0.00600816f $X=11.455
+ $Y=0.805 $X2=0 $Y2=0
cc_596 N_A_1147_408#_c_611_n N_A_876_119#_c_1295_n 0.0184822f $X=11.53 $Y=1.48
+ $X2=0 $Y2=0
cc_597 N_A_1147_408#_c_612_n N_A_876_119#_c_1295_n 0.0053093f $X=11.785 $Y=1.555
+ $X2=0 $Y2=0
cc_598 N_A_1147_408#_c_610_n N_A_876_119#_c_1296_n 0.0197188f $X=11.455 $Y=0.805
+ $X2=0 $Y2=0
cc_599 N_A_1147_408#_c_611_n N_A_876_119#_c_1296_n 0.0170607f $X=11.53 $Y=1.48
+ $X2=0 $Y2=0
cc_600 N_A_1147_408#_c_611_n N_A_876_119#_c_1297_n 0.00240348f $X=11.53 $Y=1.48
+ $X2=0 $Y2=0
cc_601 N_A_1147_408#_c_612_n N_A_876_119#_c_1297_n 0.00126813f $X=11.785
+ $Y=1.555 $X2=0 $Y2=0
cc_602 N_A_1147_408#_c_611_n N_A_876_119#_c_1298_n 0.0212362f $X=11.53 $Y=1.48
+ $X2=0 $Y2=0
cc_603 N_A_1147_408#_c_612_n N_A_876_119#_c_1298_n 0.00662536f $X=11.785
+ $Y=1.555 $X2=0 $Y2=0
cc_604 N_A_1147_408#_c_614_n N_A_2435_296#_M1003_g 0.0495762f $X=11.81 $Y=1.87
+ $X2=0 $Y2=0
cc_605 N_A_1147_408#_c_612_n N_A_2435_296#_c_1480_n 0.0495762f $X=11.785
+ $Y=1.555 $X2=0 $Y2=0
cc_606 N_A_1147_408#_c_613_n N_A_2092_47#_c_1583_n 0.00406046f $X=11.605
+ $Y=1.555 $X2=0 $Y2=0
cc_607 N_A_1147_408#_c_628_n N_A_2092_47#_c_1584_n 0.0134257f $X=11.81 $Y=1.995
+ $X2=0 $Y2=0
cc_608 N_A_1147_408#_c_614_n N_A_2092_47#_c_1584_n 3.71594e-19 $X=11.81 $Y=1.87
+ $X2=0 $Y2=0
cc_609 N_A_1147_408#_c_612_n N_A_2092_47#_c_1585_n 0.00170621f $X=11.785
+ $Y=1.555 $X2=0 $Y2=0
cc_610 N_A_1147_408#_c_628_n N_A_2092_47#_c_1585_n 0.00262547f $X=11.81 $Y=1.995
+ $X2=0 $Y2=0
cc_611 N_A_1147_408#_c_614_n N_A_2092_47#_c_1585_n 0.0148191f $X=11.81 $Y=1.87
+ $X2=0 $Y2=0
cc_612 N_A_1147_408#_c_611_n N_A_2092_47#_c_1576_n 6.08539e-19 $X=11.53 $Y=1.48
+ $X2=0 $Y2=0
cc_613 N_A_1147_408#_c_612_n N_A_2092_47#_c_1576_n 0.00138559f $X=11.785
+ $Y=1.555 $X2=0 $Y2=0
cc_614 N_A_1147_408#_c_610_n N_A_2092_47#_c_1578_n 0.00331886f $X=11.455
+ $Y=0.805 $X2=0 $Y2=0
cc_615 N_A_1147_408#_M1016_d N_A_116_419#_c_1800_n 0.00601128f $X=5.735 $Y=2.04
+ $X2=0 $Y2=0
cc_616 N_A_1147_408#_c_630_n N_A_116_419#_c_1800_n 0.0369826f $X=6.132 $Y=2.03
+ $X2=0 $Y2=0
cc_617 N_A_1147_408#_c_621_n N_A_116_419#_c_1800_n 0.00733365f $X=6.6 $Y=1.555
+ $X2=0 $Y2=0
cc_618 N_A_1147_408#_c_615_n N_A_116_419#_c_1794_n 0.0349155f $X=6.245 $Y=0.79
+ $X2=0 $Y2=0
cc_619 N_A_1147_408#_c_625_n N_A_116_419#_c_1801_n 0.00210352f $X=7.36 $Y=1.66
+ $X2=0 $Y2=0
cc_620 N_A_1147_408#_c_608_n N_A_116_419#_c_1795_n 0.0139691f $X=7.235 $Y=1.555
+ $X2=0 $Y2=0
cc_621 N_A_1147_408#_c_625_n N_A_116_419#_c_1795_n 0.00491685f $X=7.36 $Y=1.66
+ $X2=0 $Y2=0
cc_622 N_A_1147_408#_c_630_n N_A_116_419#_c_1795_n 0.0168054f $X=6.132 $Y=2.03
+ $X2=0 $Y2=0
cc_623 N_A_1147_408#_c_615_n N_A_116_419#_c_1795_n 0.0125363f $X=6.245 $Y=0.79
+ $X2=0 $Y2=0
cc_624 N_A_1147_408#_c_617_n N_A_116_419#_c_1795_n 0.00100839f $X=7.64 $Y=1.29
+ $X2=0 $Y2=0
cc_625 N_A_1147_408#_c_620_n N_A_116_419#_c_1795_n 0.0227354f $X=6.6 $Y=1.615
+ $X2=0 $Y2=0
cc_626 N_A_1147_408#_c_621_n N_A_116_419#_c_1795_n 0.00103306f $X=6.6 $Y=1.555
+ $X2=0 $Y2=0
cc_627 N_A_1147_408#_c_621_n N_A_116_419#_c_1798_n 8.8093e-19 $X=6.6 $Y=1.555
+ $X2=0 $Y2=0
cc_628 N_A_1147_408#_c_628_n N_VPWR_c_1939_n 0.00531277f $X=11.81 $Y=1.995 $X2=0
+ $Y2=0
cc_629 N_A_1147_408#_c_628_n N_VPWR_c_1947_n 0.00975641f $X=11.81 $Y=1.995 $X2=0
+ $Y2=0
cc_630 N_A_1147_408#_c_625_n N_VPWR_c_1933_n 0.0015654f $X=7.36 $Y=1.66 $X2=0
+ $Y2=0
cc_631 N_A_1147_408#_c_628_n N_VPWR_c_1933_n 0.01748f $X=11.81 $Y=1.995 $X2=0
+ $Y2=0
cc_632 N_A_1147_408#_c_618_n N_VGND_M1021_d 0.00669475f $X=10.21 $Y=0.71 $X2=0
+ $Y2=0
cc_633 N_A_1147_408#_c_615_n N_VGND_c_2165_n 0.00749171f $X=6.245 $Y=0.79 $X2=0
+ $Y2=0
cc_634 N_A_1147_408#_c_618_n N_VGND_c_2165_n 0.0174237f $X=10.21 $Y=0.71 $X2=0
+ $Y2=0
cc_635 N_A_1147_408#_c_667_p N_VGND_c_2165_n 0.00270424f $X=7.725 $Y=0.71 $X2=0
+ $Y2=0
cc_636 N_A_1147_408#_c_618_n N_VGND_c_2166_n 0.0236119f $X=10.21 $Y=0.71 $X2=0
+ $Y2=0
cc_637 N_A_1147_408#_c_610_n N_VGND_c_2171_n 0.0131584f $X=11.455 $Y=0.805 $X2=0
+ $Y2=0
cc_638 N_A_1147_408#_c_618_n N_VGND_c_2171_n 0.0125992f $X=10.21 $Y=0.71 $X2=0
+ $Y2=0
cc_639 N_A_1147_408#_c_623_n N_VGND_c_2171_n 0.00362032f $X=10.295 $Y=0.73 $X2=0
+ $Y2=0
cc_640 N_A_1147_408#_c_609_n N_VGND_c_2174_n 9.39239e-19 $X=7.73 $Y=1.125 $X2=0
+ $Y2=0
cc_641 N_A_1147_408#_c_610_n N_VGND_c_2174_n 0.0168037f $X=11.455 $Y=0.805 $X2=0
+ $Y2=0
cc_642 N_A_1147_408#_c_615_n N_VGND_c_2174_n 0.0104008f $X=6.245 $Y=0.79 $X2=0
+ $Y2=0
cc_643 N_A_1147_408#_c_618_n N_VGND_c_2174_n 0.0520535f $X=10.21 $Y=0.71 $X2=0
+ $Y2=0
cc_644 N_A_1147_408#_c_667_p N_VGND_c_2174_n 0.00444321f $X=7.725 $Y=0.71 $X2=0
+ $Y2=0
cc_645 N_A_1147_408#_c_623_n N_VGND_c_2174_n 0.00708082f $X=10.295 $Y=0.73 $X2=0
+ $Y2=0
cc_646 N_A_1147_408#_c_618_n A_1561_119# 0.00548768f $X=10.21 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_647 N_A_1147_408#_c_618_n A_1635_119# 0.00905836f $X=10.21 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_648 N_A_1147_408#_c_618_n A_1900_47# 0.00216843f $X=10.21 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_649 N_A_1605_93#_c_782_n N_RESET_B_c_907_n 0.00976941f $X=8.1 $Y=1.125 $X2=0
+ $Y2=0
cc_650 N_A_1605_93#_c_782_n N_RESET_B_M1021_g 0.0135029f $X=8.1 $Y=1.125 $X2=0
+ $Y2=0
cc_651 N_A_1605_93#_c_782_n N_RESET_B_c_912_n 0.00151839f $X=8.1 $Y=1.125 $X2=0
+ $Y2=0
cc_652 N_A_1605_93#_c_784_n N_RESET_B_c_912_n 0.00112236f $X=8.44 $Y=1.29 $X2=0
+ $Y2=0
cc_653 N_A_1605_93#_c_785_n N_RESET_B_c_912_n 0.0135476f $X=8.44 $Y=1.29 $X2=0
+ $Y2=0
cc_654 N_A_1605_93#_c_786_n N_RESET_B_c_912_n 0.0169244f $X=9.87 $Y=1.06 $X2=0
+ $Y2=0
cc_655 N_A_1605_93#_c_783_n N_RESET_B_c_913_n 0.0135316f $X=8.5 $Y=1.605 $X2=0
+ $Y2=0
cc_656 N_A_1605_93#_c_784_n N_RESET_B_c_913_n 2.06986e-19 $X=8.44 $Y=1.29 $X2=0
+ $Y2=0
cc_657 N_A_1605_93#_c_786_n N_RESET_B_c_913_n 5.83361e-19 $X=9.87 $Y=1.06 $X2=0
+ $Y2=0
cc_658 N_A_1605_93#_c_793_n N_RESET_B_M1024_g 0.0424551f $X=8.5 $Y=1.73 $X2=0
+ $Y2=0
cc_659 N_A_1605_93#_c_783_n N_RESET_B_M1024_g 0.00116138f $X=8.5 $Y=1.605 $X2=0
+ $Y2=0
cc_660 N_A_1605_93#_c_782_n N_RESET_B_c_915_n 0.00121716f $X=8.1 $Y=1.125 $X2=0
+ $Y2=0
cc_661 N_A_1605_93#_c_786_n N_RESET_B_c_915_n 0.0055849f $X=9.87 $Y=1.06 $X2=0
+ $Y2=0
cc_662 N_A_1605_93#_c_793_n N_RESET_B_c_919_n 0.00539275f $X=8.5 $Y=1.73 $X2=0
+ $Y2=0
cc_663 N_A_1605_93#_c_783_n N_RESET_B_c_919_n 0.00215976f $X=8.5 $Y=1.605 $X2=0
+ $Y2=0
cc_664 N_A_1605_93#_c_784_n N_RESET_B_c_919_n 0.0105618f $X=8.44 $Y=1.29 $X2=0
+ $Y2=0
cc_665 N_A_1605_93#_c_785_n N_RESET_B_c_919_n 0.00323793f $X=8.44 $Y=1.29 $X2=0
+ $Y2=0
cc_666 N_A_1605_93#_c_786_n N_RESET_B_c_919_n 0.005948f $X=9.87 $Y=1.06 $X2=0
+ $Y2=0
cc_667 N_A_1605_93#_c_786_n N_RESET_B_c_921_n 0.0130781f $X=9.87 $Y=1.06 $X2=0
+ $Y2=0
cc_668 N_A_1605_93#_c_788_n N_RESET_B_c_921_n 0.0178646f $X=10.605 $Y=1.36 $X2=0
+ $Y2=0
cc_669 N_A_1605_93#_c_790_n N_RESET_B_c_921_n 0.00797415f $X=9.955 $Y=1.06 $X2=0
+ $Y2=0
cc_670 N_A_1605_93#_c_797_n N_RESET_B_c_921_n 0.0302381f $X=10.855 $Y=1.85 $X2=0
+ $Y2=0
cc_671 N_A_1605_93#_c_792_n N_RESET_B_c_921_n 0.0160577f $X=10.812 $Y=1.685
+ $X2=0 $Y2=0
cc_672 N_A_1605_93#_c_793_n N_RESET_B_c_939_n 7.33862e-19 $X=8.5 $Y=1.73 $X2=0
+ $Y2=0
cc_673 N_A_1605_93#_c_783_n N_RESET_B_c_939_n 7.15185e-19 $X=8.5 $Y=1.605 $X2=0
+ $Y2=0
cc_674 N_A_1605_93#_c_786_n N_RESET_B_c_939_n 0.00225776f $X=9.87 $Y=1.06 $X2=0
+ $Y2=0
cc_675 N_A_1605_93#_c_793_n N_RESET_B_c_926_n 0.00340134f $X=8.5 $Y=1.73 $X2=0
+ $Y2=0
cc_676 N_A_1605_93#_c_784_n N_RESET_B_c_926_n 0.0138414f $X=8.44 $Y=1.29 $X2=0
+ $Y2=0
cc_677 N_A_1605_93#_c_785_n N_RESET_B_c_926_n 0.0030242f $X=8.44 $Y=1.29 $X2=0
+ $Y2=0
cc_678 N_A_1605_93#_c_786_n N_RESET_B_c_926_n 0.0299715f $X=9.87 $Y=1.06 $X2=0
+ $Y2=0
cc_679 N_A_1605_93#_c_812_n N_A_1432_119#_c_1173_n 0.00520411f $X=10.605 $Y=0.36
+ $X2=0 $Y2=0
cc_680 N_A_1605_93#_c_788_n N_A_1432_119#_c_1174_n 0.0145911f $X=10.605 $Y=1.36
+ $X2=0 $Y2=0
cc_681 N_A_1605_93#_c_790_n N_A_1432_119#_c_1174_n 0.00580523f $X=9.955 $Y=1.06
+ $X2=0 $Y2=0
cc_682 N_A_1605_93#_c_791_n N_A_1432_119#_c_1174_n 7.66668e-19 $X=10.69 $Y=1.36
+ $X2=0 $Y2=0
cc_683 N_A_1605_93#_c_792_n N_A_1432_119#_c_1174_n 0.0071666f $X=10.812 $Y=1.685
+ $X2=0 $Y2=0
cc_684 N_A_1605_93#_c_790_n N_A_1432_119#_c_1175_n 5.92482e-19 $X=9.955 $Y=1.06
+ $X2=0 $Y2=0
cc_685 N_A_1605_93#_c_796_n N_A_1432_119#_M1006_g 0.0273113f $X=10.855 $Y=2.56
+ $X2=0 $Y2=0
cc_686 N_A_1605_93#_c_797_n N_A_1432_119#_M1006_g 0.00636443f $X=10.855 $Y=1.85
+ $X2=0 $Y2=0
cc_687 N_A_1605_93#_c_792_n N_A_1432_119#_M1006_g 0.00383851f $X=10.812 $Y=1.685
+ $X2=0 $Y2=0
cc_688 N_A_1605_93#_c_786_n N_A_1432_119#_c_1176_n 6.10118e-19 $X=9.87 $Y=1.06
+ $X2=0 $Y2=0
cc_689 N_A_1605_93#_c_793_n N_A_1432_119#_c_1205_n 0.0222983f $X=8.5 $Y=1.73
+ $X2=0 $Y2=0
cc_690 N_A_1605_93#_c_784_n N_A_1432_119#_c_1205_n 0.00539945f $X=8.44 $Y=1.29
+ $X2=0 $Y2=0
cc_691 N_A_1605_93#_c_785_n N_A_1432_119#_c_1205_n 0.00196316f $X=8.44 $Y=1.29
+ $X2=0 $Y2=0
cc_692 N_A_1605_93#_c_786_n N_A_1432_119#_c_1184_n 2.74053e-19 $X=9.87 $Y=1.06
+ $X2=0 $Y2=0
cc_693 N_A_1605_93#_c_786_n N_A_1432_119#_c_1186_n 0.0228398f $X=9.87 $Y=1.06
+ $X2=0 $Y2=0
cc_694 N_A_1605_93#_c_790_n N_A_1432_119#_c_1186_n 0.00849809f $X=9.955 $Y=1.06
+ $X2=0 $Y2=0
cc_695 N_A_1605_93#_c_786_n N_A_1432_119#_c_1178_n 0.0250657f $X=9.87 $Y=1.06
+ $X2=0 $Y2=0
cc_696 N_A_1605_93#_c_788_n N_A_1432_119#_c_1178_n 7.71134e-19 $X=10.605 $Y=1.36
+ $X2=0 $Y2=0
cc_697 N_A_1605_93#_c_790_n N_A_1432_119#_c_1178_n 0.0170039f $X=9.955 $Y=1.06
+ $X2=0 $Y2=0
cc_698 N_A_1605_93#_c_793_n N_A_876_119#_M1042_g 0.0840131f $X=8.5 $Y=1.73 $X2=0
+ $Y2=0
cc_699 N_A_1605_93#_c_785_n N_A_876_119#_M1042_g 0.0104784f $X=8.44 $Y=1.29
+ $X2=0 $Y2=0
cc_700 N_A_1605_93#_c_793_n N_A_876_119#_c_1304_n 0.0171865f $X=8.5 $Y=1.73
+ $X2=0 $Y2=0
cc_701 N_A_1605_93#_c_796_n N_A_876_119#_c_1304_n 0.00544492f $X=10.855 $Y=2.56
+ $X2=0 $Y2=0
cc_702 N_A_1605_93#_c_796_n N_A_876_119#_M1002_g 0.0135409f $X=10.855 $Y=2.56
+ $X2=0 $Y2=0
cc_703 N_A_1605_93#_c_797_n N_A_876_119#_M1002_g 0.00356504f $X=10.855 $Y=1.85
+ $X2=0 $Y2=0
cc_704 N_A_1605_93#_c_792_n N_A_876_119#_M1002_g 0.00438676f $X=10.812 $Y=1.685
+ $X2=0 $Y2=0
cc_705 N_A_1605_93#_c_789_n N_A_876_119#_c_1295_n 0.0117464f $X=10.69 $Y=1.275
+ $X2=0 $Y2=0
cc_706 N_A_1605_93#_c_791_n N_A_876_119#_c_1295_n 0.0145108f $X=10.69 $Y=1.36
+ $X2=0 $Y2=0
cc_707 N_A_1605_93#_c_797_n N_A_876_119#_c_1295_n 0.00291745f $X=10.855 $Y=1.85
+ $X2=0 $Y2=0
cc_708 N_A_1605_93#_c_789_n N_A_876_119#_c_1296_n 0.00363043f $X=10.69 $Y=1.275
+ $X2=0 $Y2=0
cc_709 N_A_1605_93#_c_791_n N_A_876_119#_c_1296_n 0.00379971f $X=10.69 $Y=1.36
+ $X2=0 $Y2=0
cc_710 N_A_1605_93#_c_797_n N_A_876_119#_c_1296_n 0.00218713f $X=10.855 $Y=1.85
+ $X2=0 $Y2=0
cc_711 N_A_1605_93#_c_812_n N_A_2092_47#_M1039_d 0.0126332f $X=10.605 $Y=0.36
+ $X2=-0.19 $Y2=-0.245
cc_712 N_A_1605_93#_c_789_n N_A_2092_47#_M1039_d 0.0110436f $X=10.69 $Y=1.275
+ $X2=-0.19 $Y2=-0.245
cc_713 N_A_1605_93#_c_797_n N_A_2092_47#_c_1583_n 0.00485083f $X=10.855 $Y=1.85
+ $X2=0 $Y2=0
cc_714 N_A_1605_93#_c_797_n N_A_2092_47#_c_1584_n 0.0232231f $X=10.855 $Y=1.85
+ $X2=0 $Y2=0
cc_715 N_A_1605_93#_c_793_n N_VPWR_c_1937_n 0.0141686f $X=8.5 $Y=1.73 $X2=0
+ $Y2=0
cc_716 N_A_1605_93#_c_788_n N_VPWR_c_1938_n 0.0143594f $X=10.605 $Y=1.36 $X2=0
+ $Y2=0
cc_717 N_A_1605_93#_c_797_n N_VPWR_c_1938_n 0.0705218f $X=10.855 $Y=1.85 $X2=0
+ $Y2=0
cc_718 N_A_1605_93#_c_796_n N_VPWR_c_1947_n 0.00877739f $X=10.855 $Y=2.56 $X2=0
+ $Y2=0
cc_719 N_A_1605_93#_c_793_n N_VPWR_c_1933_n 0.0013212f $X=8.5 $Y=1.73 $X2=0
+ $Y2=0
cc_720 N_A_1605_93#_c_796_n N_VPWR_c_1933_n 0.0110988f $X=10.855 $Y=2.56 $X2=0
+ $Y2=0
cc_721 N_A_1605_93#_c_812_n N_VGND_c_2171_n 0.04121f $X=10.605 $Y=0.36 $X2=0
+ $Y2=0
cc_722 N_A_1605_93#_M1033_d N_VGND_c_2174_n 0.00379383f $X=9.89 $Y=0.235 $X2=0
+ $Y2=0
cc_723 N_A_1605_93#_c_782_n N_VGND_c_2174_n 9.39239e-19 $X=8.1 $Y=1.125 $X2=0
+ $Y2=0
cc_724 N_A_1605_93#_c_812_n N_VGND_c_2174_n 0.0280679f $X=10.605 $Y=0.36 $X2=0
+ $Y2=0
cc_725 N_A_1605_93#_c_787_n A_1635_119# 0.00363567f $X=8.555 $Y=1.06 $X2=-0.19
+ $Y2=-0.245
cc_726 N_RESET_B_c_919_n N_A_1432_119#_M1019_d 0.0032385f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_727 N_RESET_B_c_921_n N_A_1432_119#_M1024_d 0.00141907f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_728 N_RESET_B_c_907_n N_A_1432_119#_c_1173_n 0.00704173f $X=8.645 $Y=0.18
+ $X2=0 $Y2=0
cc_729 N_RESET_B_c_921_n N_A_1432_119#_c_1175_n 0.0172836f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_730 N_RESET_B_c_921_n N_A_1432_119#_M1006_g 0.0112504f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_731 N_RESET_B_M1021_g N_A_1432_119#_c_1176_n 0.00704173f $X=8.72 $Y=0.54
+ $X2=0 $Y2=0
cc_732 N_RESET_B_c_915_n N_A_1432_119#_c_1176_n 0.00795276f $X=8.72 $Y=0.9 $X2=0
+ $Y2=0
cc_733 N_RESET_B_c_907_n N_A_1432_119#_c_1177_n 0.00327715f $X=8.645 $Y=0.18
+ $X2=0 $Y2=0
cc_734 N_RESET_B_c_919_n N_A_1432_119#_c_1177_n 0.0257126f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_735 N_RESET_B_M1024_g N_A_1432_119#_c_1205_n 0.0239542f $X=9.03 $Y=2.235
+ $X2=0 $Y2=0
cc_736 N_RESET_B_c_919_n N_A_1432_119#_c_1205_n 0.0322231f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_737 N_RESET_B_c_921_n N_A_1432_119#_c_1205_n 0.00459694f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_738 N_RESET_B_c_939_n N_A_1432_119#_c_1205_n 0.00332881f $X=9.025 $Y=1.665
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_926_n N_A_1432_119#_c_1205_n 0.0212518f $X=8.995 $Y=1.41
+ $X2=0 $Y2=0
cc_740 N_RESET_B_M1024_g N_A_1432_119#_c_1184_n 0.00731018f $X=9.03 $Y=2.235
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_921_n N_A_1432_119#_c_1184_n 0.023989f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_939_n N_A_1432_119#_c_1184_n 2.45435e-19 $X=9.025 $Y=1.665
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_926_n N_A_1432_119#_c_1184_n 0.00305529f $X=8.995 $Y=1.41
+ $X2=0 $Y2=0
cc_744 N_RESET_B_M1024_g N_A_1432_119#_c_1185_n 0.019174f $X=9.03 $Y=2.235 $X2=0
+ $Y2=0
cc_745 N_RESET_B_c_913_n N_A_1432_119#_c_1186_n 2.87181e-19 $X=9.03 $Y=1.575
+ $X2=0 $Y2=0
cc_746 N_RESET_B_M1024_g N_A_1432_119#_c_1186_n 8.44126e-19 $X=9.03 $Y=2.235
+ $X2=0 $Y2=0
cc_747 N_RESET_B_c_921_n N_A_1432_119#_c_1186_n 0.0146097f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_939_n N_A_1432_119#_c_1186_n 2.26943e-19 $X=9.025 $Y=1.665
+ $X2=0 $Y2=0
cc_749 N_RESET_B_c_926_n N_A_1432_119#_c_1186_n 0.0300703f $X=8.995 $Y=1.41
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_913_n N_A_1432_119#_c_1178_n 0.0256061f $X=9.03 $Y=1.575
+ $X2=0 $Y2=0
cc_751 N_RESET_B_c_915_n N_A_1432_119#_c_1178_n 0.0176441f $X=8.72 $Y=0.9 $X2=0
+ $Y2=0
cc_752 N_RESET_B_c_926_n N_A_1432_119#_c_1178_n 0.00157087f $X=8.995 $Y=1.41
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_919_n N_A_1432_119#_c_1206_n 0.0185207f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_907_n N_A_876_119#_c_1286_n 0.010259f $X=8.645 $Y=0.18 $X2=0
+ $Y2=0
cc_755 N_RESET_B_c_907_n N_A_876_119#_M1029_g 0.0104164f $X=8.645 $Y=0.18 $X2=0
+ $Y2=0
cc_756 N_RESET_B_c_919_n N_A_876_119#_c_1288_n 0.00141438f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_907_n N_A_876_119#_c_1289_n 0.0103053f $X=8.645 $Y=0.18 $X2=0
+ $Y2=0
cc_758 N_RESET_B_c_919_n N_A_876_119#_M1042_g 0.00628038f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_759 N_RESET_B_M1024_g N_A_876_119#_c_1304_n 0.0173232f $X=9.03 $Y=2.235 $X2=0
+ $Y2=0
cc_760 N_RESET_B_c_921_n N_A_876_119#_M1002_g 0.0137156f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_907_n N_A_876_119#_c_1292_n 0.00325143f $X=8.645 $Y=0.18
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_919_n N_A_876_119#_c_1292_n 0.014369f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_763 N_RESET_B_c_919_n N_A_876_119#_c_1309_n 0.0659037f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_919_n N_A_876_119#_c_1293_n 0.0219626f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_765 N_RESET_B_c_919_n N_A_876_119#_c_1294_n 0.00930364f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_921_n N_A_876_119#_c_1295_n 0.0266393f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_767 N_RESET_B_c_921_n N_A_876_119#_c_1296_n 0.00195965f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_768 N_RESET_B_c_919_n N_A_876_119#_c_1311_n 0.0173846f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_921_n N_A_876_119#_c_1297_n 0.00764079f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_921_n N_A_876_119#_c_1298_n 8.92391e-19 $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_771 N_RESET_B_c_917_n N_A_2435_296#_M1003_g 0.00548132f $X=13.285 $Y=1.7
+ $X2=0 $Y2=0
cc_772 N_RESET_B_c_934_n N_A_2435_296#_M1003_g 0.00193069f $X=13.32 $Y=1.77
+ $X2=0 $Y2=0
cc_773 N_RESET_B_c_921_n N_A_2435_296#_M1003_g 3.06333e-19 $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_774 N_RESET_B_c_927_n N_A_2435_296#_M1003_g 9.625e-19 $X=12.835 $Y=1.667
+ $X2=0 $Y2=0
cc_775 N_RESET_B_M1012_g N_A_2435_296#_M1034_g 0.0162661f $X=13.23 $Y=0.445
+ $X2=0 $Y2=0
cc_776 N_RESET_B_M1012_g N_A_2435_296#_c_1472_n 0.00911291f $X=13.23 $Y=0.445
+ $X2=0 $Y2=0
cc_777 N_RESET_B_c_918_n N_A_2435_296#_c_1472_n 0.00615096f $X=13.32 $Y=1.77
+ $X2=0 $Y2=0
cc_778 N_RESET_B_M1012_g N_A_2435_296#_c_1473_n 0.00105054f $X=13.23 $Y=0.445
+ $X2=0 $Y2=0
cc_779 N_RESET_B_c_916_n N_A_2435_296#_c_1476_n 0.0101401f $X=13.085 $Y=1.7
+ $X2=0 $Y2=0
cc_780 RESET_B N_A_2435_296#_c_1476_n 0.00629495f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_781 N_RESET_B_c_927_n N_A_2435_296#_c_1476_n 0.0124413f $X=12.835 $Y=1.667
+ $X2=0 $Y2=0
cc_782 N_RESET_B_M1012_g N_A_2435_296#_c_1477_n 0.00987487f $X=13.23 $Y=0.445
+ $X2=0 $Y2=0
cc_783 N_RESET_B_c_916_n N_A_2435_296#_c_1477_n 0.00540798f $X=13.085 $Y=1.7
+ $X2=0 $Y2=0
cc_784 N_RESET_B_c_917_n N_A_2435_296#_c_1477_n 0.0299106f $X=13.285 $Y=1.7
+ $X2=0 $Y2=0
cc_785 N_RESET_B_M1028_g N_A_2435_296#_c_1499_n 0.0248042f $X=13.395 $Y=2.595
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_934_n N_A_2435_296#_c_1499_n 0.0541498f $X=13.32 $Y=1.77
+ $X2=0 $Y2=0
cc_787 N_RESET_B_M1012_g N_A_2435_296#_c_1478_n 0.00304777f $X=13.23 $Y=0.445
+ $X2=0 $Y2=0
cc_788 N_RESET_B_c_917_n N_A_2435_296#_c_1478_n 0.0233777f $X=13.285 $Y=1.7
+ $X2=0 $Y2=0
cc_789 N_RESET_B_c_934_n N_A_2435_296#_c_1478_n 0.00761094f $X=13.32 $Y=1.77
+ $X2=0 $Y2=0
cc_790 N_RESET_B_c_918_n N_A_2435_296#_c_1478_n 0.00378871f $X=13.32 $Y=1.77
+ $X2=0 $Y2=0
cc_791 N_RESET_B_M1012_g N_A_2435_296#_c_1480_n 0.0262565f $X=13.23 $Y=0.445
+ $X2=0 $Y2=0
cc_792 N_RESET_B_c_916_n N_A_2435_296#_c_1480_n 0.0023221f $X=13.085 $Y=1.7
+ $X2=0 $Y2=0
cc_793 N_RESET_B_c_921_n N_A_2435_296#_c_1480_n 0.00945994f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_794 RESET_B N_A_2435_296#_c_1480_n 0.00838873f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_795 N_RESET_B_c_927_n N_A_2435_296#_c_1480_n 0.00519383f $X=12.835 $Y=1.667
+ $X2=0 $Y2=0
cc_796 N_RESET_B_c_921_n N_A_2092_47#_M1002_d 0.00205389f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_797 N_RESET_B_M1012_g N_A_2092_47#_c_1567_n 0.0365417f $X=13.23 $Y=0.445
+ $X2=0 $Y2=0
cc_798 N_RESET_B_M1012_g N_A_2092_47#_M1004_g 0.0109364f $X=13.23 $Y=0.445 $X2=0
+ $Y2=0
cc_799 N_RESET_B_c_917_n N_A_2092_47#_M1004_g 3.08338e-19 $X=13.285 $Y=1.7 $X2=0
+ $Y2=0
cc_800 N_RESET_B_c_934_n N_A_2092_47#_M1004_g 4.12812e-19 $X=13.32 $Y=1.77 $X2=0
+ $Y2=0
cc_801 N_RESET_B_c_918_n N_A_2092_47#_M1004_g 0.0379734f $X=13.32 $Y=1.77 $X2=0
+ $Y2=0
cc_802 N_RESET_B_M1012_g N_A_2092_47#_c_1570_n 0.0218037f $X=13.23 $Y=0.445
+ $X2=0 $Y2=0
cc_803 N_RESET_B_c_921_n N_A_2092_47#_c_1583_n 0.0223342f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_804 N_RESET_B_c_917_n N_A_2092_47#_c_1585_n 0.00254797f $X=13.285 $Y=1.7
+ $X2=0 $Y2=0
cc_805 N_RESET_B_c_918_n N_A_2092_47#_c_1585_n 4.85043e-19 $X=13.32 $Y=1.77
+ $X2=0 $Y2=0
cc_806 N_RESET_B_c_921_n N_A_2092_47#_c_1585_n 0.0436925f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_807 RESET_B N_A_2092_47#_c_1585_n 0.00141679f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_808 N_RESET_B_c_927_n N_A_2092_47#_c_1585_n 0.00698429f $X=12.835 $Y=1.667
+ $X2=0 $Y2=0
cc_809 N_RESET_B_c_921_n N_A_2092_47#_c_1576_n 0.0138982f $X=12.575 $Y=1.665
+ $X2=0 $Y2=0
cc_810 RESET_B N_A_2092_47#_c_1576_n 0.00136277f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_811 N_RESET_B_c_927_n N_A_2092_47#_c_1576_n 0.0085675f $X=12.835 $Y=1.667
+ $X2=0 $Y2=0
cc_812 N_RESET_B_M1012_g N_A_2092_47#_c_1577_n 0.013815f $X=13.23 $Y=0.445 $X2=0
+ $Y2=0
cc_813 N_RESET_B_M1012_g N_A_2092_47#_c_1580_n 0.00147539f $X=13.23 $Y=0.445
+ $X2=0 $Y2=0
cc_814 N_RESET_B_c_919_n N_A_116_419#_M1019_s 0.00684629f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_815 N_RESET_B_M1009_g N_A_116_419#_c_1806_n 0.0162593f $X=3.12 $Y=2.595 $X2=0
+ $Y2=0
cc_816 N_RESET_B_M1009_g N_A_116_419#_c_1835_n 6.2758e-19 $X=3.12 $Y=2.595 $X2=0
+ $Y2=0
cc_817 N_RESET_B_c_907_n N_A_116_419#_c_1794_n 0.00575488f $X=8.645 $Y=0.18
+ $X2=0 $Y2=0
cc_818 N_RESET_B_c_919_n N_A_116_419#_c_1795_n 0.0190302f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_819 N_RESET_B_M1009_g N_A_116_419#_c_1817_n 0.005519f $X=3.12 $Y=2.595 $X2=0
+ $Y2=0
cc_820 N_RESET_B_M1009_g N_A_116_419#_c_1818_n 0.00797523f $X=3.12 $Y=2.595
+ $X2=0 $Y2=0
cc_821 N_RESET_B_c_919_n N_A_116_419#_c_1798_n 0.0050568f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_822 N_RESET_B_c_919_n N_VPWR_M1045_d 9.15774e-19 $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_823 N_RESET_B_c_939_n N_VPWR_M1045_d 0.00170621f $X=9.025 $Y=1.665 $X2=0
+ $Y2=0
cc_824 N_RESET_B_c_926_n N_VPWR_M1045_d 0.00118448f $X=8.995 $Y=1.41 $X2=0 $Y2=0
cc_825 N_RESET_B_c_934_n N_VPWR_M1003_d 0.0140341f $X=13.32 $Y=1.77 $X2=0 $Y2=0
cc_826 N_RESET_B_M1009_g N_VPWR_c_1935_n 0.00950776f $X=3.12 $Y=2.595 $X2=0
+ $Y2=0
cc_827 N_RESET_B_M1024_g N_VPWR_c_1937_n 0.0143459f $X=9.03 $Y=2.235 $X2=0 $Y2=0
cc_828 N_RESET_B_c_921_n N_VPWR_c_1938_n 0.0229431f $X=12.575 $Y=1.665 $X2=0
+ $Y2=0
cc_829 N_RESET_B_M1028_g N_VPWR_c_1939_n 0.0100463f $X=13.395 $Y=2.595 $X2=0
+ $Y2=0
cc_830 N_RESET_B_c_934_n N_VPWR_c_1939_n 0.0312403f $X=13.32 $Y=1.77 $X2=0 $Y2=0
cc_831 N_RESET_B_c_921_n N_VPWR_c_1939_n 0.00567474f $X=12.575 $Y=1.665 $X2=0
+ $Y2=0
cc_832 RESET_B N_VPWR_c_1939_n 0.00302885f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_833 N_RESET_B_c_927_n N_VPWR_c_1939_n 6.9263e-19 $X=12.835 $Y=1.667 $X2=0
+ $Y2=0
cc_834 N_RESET_B_M1028_g N_VPWR_c_1940_n 0.00124663f $X=13.395 $Y=2.595 $X2=0
+ $Y2=0
cc_835 N_RESET_B_M1009_g N_VPWR_c_1943_n 0.00631431f $X=3.12 $Y=2.595 $X2=0
+ $Y2=0
cc_836 N_RESET_B_M1028_g N_VPWR_c_1952_n 0.00883214f $X=13.395 $Y=2.595 $X2=0
+ $Y2=0
cc_837 N_RESET_B_c_934_n N_VPWR_c_1952_n 0.00630371f $X=13.32 $Y=1.77 $X2=0
+ $Y2=0
cc_838 N_RESET_B_M1009_g N_VPWR_c_1933_n 0.00698085f $X=3.12 $Y=2.595 $X2=0
+ $Y2=0
cc_839 N_RESET_B_M1024_g N_VPWR_c_1933_n 0.00150904f $X=9.03 $Y=2.235 $X2=0
+ $Y2=0
cc_840 N_RESET_B_M1028_g N_VPWR_c_1933_n 0.0160775f $X=13.395 $Y=2.595 $X2=0
+ $Y2=0
cc_841 N_RESET_B_c_934_n N_VPWR_c_1933_n 0.00773033f $X=13.32 $Y=1.77 $X2=0
+ $Y2=0
cc_842 N_RESET_B_c_919_n A_1633_347# 0.00176433f $X=8.735 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_843 N_RESET_B_M1011_g N_noxref_23_c_2134_n 0.00519347f $X=2.43 $Y=0.65 $X2=0
+ $Y2=0
cc_844 N_RESET_B_M1011_g N_noxref_23_c_2135_n 0.00584187f $X=2.43 $Y=0.65 $X2=0
+ $Y2=0
cc_845 N_RESET_B_M1011_g N_VGND_c_2163_n 0.0106317f $X=2.43 $Y=0.65 $X2=0 $Y2=0
cc_846 N_RESET_B_c_907_n N_VGND_c_2163_n 0.0246054f $X=8.645 $Y=0.18 $X2=0 $Y2=0
cc_847 N_RESET_B_c_909_n N_VGND_c_2163_n 0.00648299f $X=2.975 $Y=1.165 $X2=0
+ $Y2=0
cc_848 N_RESET_B_c_907_n N_VGND_c_2164_n 0.0255538f $X=8.645 $Y=0.18 $X2=0 $Y2=0
cc_849 N_RESET_B_c_907_n N_VGND_c_2165_n 0.0926739f $X=8.645 $Y=0.18 $X2=0 $Y2=0
cc_850 N_RESET_B_c_907_n N_VGND_c_2166_n 0.00706267f $X=8.645 $Y=0.18 $X2=0
+ $Y2=0
cc_851 N_RESET_B_M1012_g N_VGND_c_2167_n 0.00959775f $X=13.23 $Y=0.445 $X2=0
+ $Y2=0
cc_852 N_RESET_B_c_908_n N_VGND_c_2169_n 0.00758518f $X=2.505 $Y=0.18 $X2=0
+ $Y2=0
cc_853 N_RESET_B_c_907_n N_VGND_c_2170_n 0.0755883f $X=8.645 $Y=0.18 $X2=0 $Y2=0
cc_854 N_RESET_B_M1012_g N_VGND_c_2172_n 0.00433016f $X=13.23 $Y=0.445 $X2=0
+ $Y2=0
cc_855 N_RESET_B_c_907_n N_VGND_c_2174_n 0.211648f $X=8.645 $Y=0.18 $X2=0 $Y2=0
cc_856 N_RESET_B_c_908_n N_VGND_c_2174_n 0.0105575f $X=2.505 $Y=0.18 $X2=0 $Y2=0
cc_857 N_RESET_B_M1012_g N_VGND_c_2174_n 0.00676843f $X=13.23 $Y=0.445 $X2=0
+ $Y2=0
cc_858 N_A_1432_119#_c_1183_n N_A_876_119#_c_1301_n 0.00727294f $X=7.625
+ $Y=2.235 $X2=0 $Y2=0
cc_859 N_A_1432_119#_c_1177_n N_A_876_119#_c_1289_n 0.00223845f $X=7.3 $Y=0.79
+ $X2=0 $Y2=0
cc_860 N_A_1432_119#_c_1177_n N_A_876_119#_M1042_g 0.00106757f $X=7.3 $Y=0.79
+ $X2=0 $Y2=0
cc_861 N_A_1432_119#_c_1205_n N_A_876_119#_M1042_g 0.0207936f $X=9.275 $Y=2.045
+ $X2=0 $Y2=0
cc_862 N_A_1432_119#_c_1206_n N_A_876_119#_M1042_g 0.0242021f $X=7.625 $Y=1.88
+ $X2=0 $Y2=0
cc_863 N_A_1432_119#_M1006_g N_A_876_119#_c_1304_n 0.0148452f $X=10.51 $Y=2.205
+ $X2=0 $Y2=0
cc_864 N_A_1432_119#_c_1185_n N_A_876_119#_c_1304_n 0.00859255f $X=9.44 $Y=2.235
+ $X2=0 $Y2=0
cc_865 N_A_1432_119#_c_1174_n N_A_876_119#_M1002_g 0.0288844f $X=10.385 $Y=1.5
+ $X2=0 $Y2=0
cc_866 N_A_1432_119#_c_1174_n N_A_876_119#_c_1296_n 0.00107671f $X=10.385 $Y=1.5
+ $X2=0 $Y2=0
cc_867 N_A_1432_119#_c_1177_n N_A_116_419#_c_1794_n 0.0884162f $X=7.3 $Y=0.79
+ $X2=0 $Y2=0
cc_868 N_A_1432_119#_c_1183_n N_A_116_419#_c_1801_n 0.012543f $X=7.625 $Y=2.235
+ $X2=0 $Y2=0
cc_869 N_A_1432_119#_c_1205_n N_VPWR_M1045_d 0.0037231f $X=9.275 $Y=2.045 $X2=0
+ $Y2=0
cc_870 N_A_1432_119#_c_1205_n N_VPWR_c_1937_n 0.0158111f $X=9.275 $Y=2.045 $X2=0
+ $Y2=0
cc_871 N_A_1432_119#_c_1185_n N_VPWR_c_1937_n 0.0198399f $X=9.44 $Y=2.235 $X2=0
+ $Y2=0
cc_872 N_A_1432_119#_c_1174_n N_VPWR_c_1938_n 0.00647868f $X=10.385 $Y=1.5 $X2=0
+ $Y2=0
cc_873 N_A_1432_119#_M1006_g N_VPWR_c_1938_n 0.0229878f $X=10.51 $Y=2.205 $X2=0
+ $Y2=0
cc_874 N_A_1432_119#_c_1184_n N_VPWR_c_1938_n 0.0200556f $X=9.487 $Y=2.13 $X2=0
+ $Y2=0
cc_875 N_A_1432_119#_c_1185_n N_VPWR_c_1938_n 0.03041f $X=9.44 $Y=2.235 $X2=0
+ $Y2=0
cc_876 N_A_1432_119#_c_1186_n N_VPWR_c_1938_n 9.43529e-19 $X=9.535 $Y=1.41 $X2=0
+ $Y2=0
cc_877 N_A_1432_119#_c_1183_n N_VPWR_c_1950_n 0.0126017f $X=7.625 $Y=2.235 $X2=0
+ $Y2=0
cc_878 N_A_1432_119#_c_1185_n N_VPWR_c_1951_n 0.00973836f $X=9.44 $Y=2.235 $X2=0
+ $Y2=0
cc_879 N_A_1432_119#_M1006_g N_VPWR_c_1933_n 0.00143131f $X=10.51 $Y=2.205 $X2=0
+ $Y2=0
cc_880 N_A_1432_119#_c_1183_n N_VPWR_c_1933_n 0.0156092f $X=7.625 $Y=2.235 $X2=0
+ $Y2=0
cc_881 N_A_1432_119#_c_1185_n N_VPWR_c_1933_n 0.011736f $X=9.44 $Y=2.235 $X2=0
+ $Y2=0
cc_882 N_A_1432_119#_c_1205_n A_1633_347# 0.00479889f $X=9.275 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_883 N_A_1432_119#_c_1177_n N_VGND_c_2165_n 0.003298f $X=7.3 $Y=0.79 $X2=0
+ $Y2=0
cc_884 N_A_1432_119#_c_1173_n N_VGND_c_2166_n 0.00797533f $X=9.425 $Y=0.73 $X2=0
+ $Y2=0
cc_885 N_A_1432_119#_c_1173_n N_VGND_c_2171_n 0.0084722f $X=9.425 $Y=0.73 $X2=0
+ $Y2=0
cc_886 N_A_1432_119#_c_1173_n N_VGND_c_2174_n 0.0127112f $X=9.425 $Y=0.73 $X2=0
+ $Y2=0
cc_887 N_A_1432_119#_c_1177_n N_VGND_c_2174_n 0.00446681f $X=7.3 $Y=0.79 $X2=0
+ $Y2=0
cc_888 N_A_876_119#_M1020_g N_A_2435_296#_M1034_g 0.023379f $X=11.92 $Y=0.445
+ $X2=0 $Y2=0
cc_889 N_A_876_119#_c_1297_n N_A_2435_296#_M1034_g 3.26261e-19 $X=11.98 $Y=1.075
+ $X2=0 $Y2=0
cc_890 N_A_876_119#_c_1298_n N_A_2435_296#_M1034_g 0.0172781f $X=11.98 $Y=1.075
+ $X2=0 $Y2=0
cc_891 N_A_876_119#_c_1297_n N_A_2435_296#_c_1480_n 0.00119061f $X=11.98
+ $Y=1.075 $X2=0 $Y2=0
cc_892 N_A_876_119#_M1002_g N_A_2092_47#_c_1583_n 0.00147089f $X=11.12 $Y=2.205
+ $X2=0 $Y2=0
cc_893 N_A_876_119#_c_1295_n N_A_2092_47#_c_1583_n 0.0160611f $X=11.815 $Y=1.285
+ $X2=0 $Y2=0
cc_894 N_A_876_119#_M1002_g N_A_2092_47#_c_1584_n 0.0163077f $X=11.12 $Y=2.205
+ $X2=0 $Y2=0
cc_895 N_A_876_119#_c_1295_n N_A_2092_47#_c_1585_n 0.00887261f $X=11.815
+ $Y=1.285 $X2=0 $Y2=0
cc_896 N_A_876_119#_c_1297_n N_A_2092_47#_c_1585_n 0.0142145f $X=11.98 $Y=1.075
+ $X2=0 $Y2=0
cc_897 N_A_876_119#_c_1298_n N_A_2092_47#_c_1585_n 0.0017104f $X=11.98 $Y=1.075
+ $X2=0 $Y2=0
cc_898 N_A_876_119#_M1020_g N_A_2092_47#_c_1575_n 0.00993283f $X=11.92 $Y=0.445
+ $X2=0 $Y2=0
cc_899 N_A_876_119#_c_1297_n N_A_2092_47#_c_1575_n 0.0156484f $X=11.98 $Y=1.075
+ $X2=0 $Y2=0
cc_900 N_A_876_119#_c_1298_n N_A_2092_47#_c_1575_n 0.00218689f $X=11.98 $Y=1.075
+ $X2=0 $Y2=0
cc_901 N_A_876_119#_c_1297_n N_A_2092_47#_c_1576_n 0.0393511f $X=11.98 $Y=1.075
+ $X2=0 $Y2=0
cc_902 N_A_876_119#_c_1298_n N_A_2092_47#_c_1576_n 0.00202895f $X=11.98 $Y=1.075
+ $X2=0 $Y2=0
cc_903 N_A_876_119#_M1020_g N_A_2092_47#_c_1578_n 4.70508e-19 $X=11.92 $Y=0.445
+ $X2=0 $Y2=0
cc_904 N_A_876_119#_c_1295_n N_A_2092_47#_c_1578_n 0.0128525f $X=11.815 $Y=1.285
+ $X2=0 $Y2=0
cc_905 N_A_876_119#_c_1297_n N_A_2092_47#_c_1578_n 0.00151785f $X=11.98 $Y=1.075
+ $X2=0 $Y2=0
cc_906 N_A_876_119#_M1020_g N_A_2092_47#_c_1579_n 0.00455611f $X=11.92 $Y=0.445
+ $X2=0 $Y2=0
cc_907 N_A_876_119#_M1031_s N_A_116_419#_c_1799_n 0.00331943f $X=4.44 $Y=2.04
+ $X2=0 $Y2=0
cc_908 N_A_876_119#_c_1308_n N_A_116_419#_c_1799_n 0.0179944f $X=4.585 $Y=2.185
+ $X2=0 $Y2=0
cc_909 N_A_876_119#_M1016_g N_A_116_419#_c_1800_n 0.0216514f $X=5.61 $Y=2.54
+ $X2=0 $Y2=0
cc_910 N_A_876_119#_c_1300_n N_A_116_419#_c_1800_n 0.0145838f $X=6.15 $Y=3.075
+ $X2=0 $Y2=0
cc_911 N_A_876_119#_c_1301_n N_A_116_419#_c_1800_n 0.00921876f $X=7.915 $Y=3.15
+ $X2=0 $Y2=0
cc_912 N_A_876_119#_c_1309_n N_A_116_419#_c_1800_n 0.0187782f $X=5.475 $Y=1.765
+ $X2=0 $Y2=0
cc_913 N_A_876_119#_c_1309_n N_A_116_419#_c_1846_n 0.00406528f $X=5.475 $Y=1.765
+ $X2=0 $Y2=0
cc_914 N_A_876_119#_c_1286_n N_A_116_419#_c_1794_n 0.00103623f $X=5.67 $Y=1.18
+ $X2=0 $Y2=0
cc_915 N_A_876_119#_c_1289_n N_A_116_419#_c_1794_n 0.00473273f $X=7.085 $Y=1.09
+ $X2=0 $Y2=0
cc_916 N_A_876_119#_c_1300_n N_A_116_419#_c_1801_n 0.00263889f $X=6.15 $Y=3.075
+ $X2=0 $Y2=0
cc_917 N_A_876_119#_c_1301_n N_A_116_419#_c_1801_n 0.00345327f $X=7.915 $Y=3.15
+ $X2=0 $Y2=0
cc_918 N_A_876_119#_c_1300_n N_A_116_419#_c_1795_n 0.0049652f $X=6.15 $Y=3.075
+ $X2=0 $Y2=0
cc_919 N_A_876_119#_c_1288_n N_A_116_419#_c_1795_n 0.00584031f $X=7.01 $Y=1.165
+ $X2=0 $Y2=0
cc_920 N_A_876_119#_c_1294_n N_A_116_419#_c_1795_n 0.00172308f $X=5.64 $Y=1.345
+ $X2=0 $Y2=0
cc_921 N_A_876_119#_c_1288_n N_A_116_419#_c_1798_n 0.00908349f $X=7.01 $Y=1.165
+ $X2=0 $Y2=0
cc_922 N_A_876_119#_c_1289_n N_A_116_419#_c_1798_n 0.0032691f $X=7.085 $Y=1.09
+ $X2=0 $Y2=0
cc_923 N_A_876_119#_M1016_g N_VPWR_c_1936_n 0.0104965f $X=5.61 $Y=2.54 $X2=0
+ $Y2=0
cc_924 N_A_876_119#_c_1300_n N_VPWR_c_1936_n 0.0017053f $X=6.15 $Y=3.075 $X2=0
+ $Y2=0
cc_925 N_A_876_119#_c_1302_n N_VPWR_c_1936_n 8.53695e-19 $X=6.225 $Y=3.15 $X2=0
+ $Y2=0
cc_926 N_A_876_119#_M1042_g N_VPWR_c_1937_n 0.00877352f $X=8.04 $Y=2.235 $X2=0
+ $Y2=0
cc_927 N_A_876_119#_c_1304_n N_VPWR_c_1937_n 0.0254328f $X=10.995 $Y=3.15 $X2=0
+ $Y2=0
cc_928 N_A_876_119#_c_1304_n N_VPWR_c_1938_n 0.0258253f $X=10.995 $Y=3.15 $X2=0
+ $Y2=0
cc_929 N_A_876_119#_M1002_g N_VPWR_c_1938_n 0.0068035f $X=11.12 $Y=2.205 $X2=0
+ $Y2=0
cc_930 N_A_876_119#_c_1304_n N_VPWR_c_1947_n 0.0261613f $X=10.995 $Y=3.15 $X2=0
+ $Y2=0
cc_931 N_A_876_119#_M1016_g N_VPWR_c_1950_n 0.00583726f $X=5.61 $Y=2.54 $X2=0
+ $Y2=0
cc_932 N_A_876_119#_c_1302_n N_VPWR_c_1950_n 0.0746654f $X=6.225 $Y=3.15 $X2=0
+ $Y2=0
cc_933 N_A_876_119#_c_1304_n N_VPWR_c_1951_n 0.0363059f $X=10.995 $Y=3.15 $X2=0
+ $Y2=0
cc_934 N_A_876_119#_M1016_g N_VPWR_c_1933_n 0.00716285f $X=5.61 $Y=2.54 $X2=0
+ $Y2=0
cc_935 N_A_876_119#_c_1301_n N_VPWR_c_1933_n 0.0543976f $X=7.915 $Y=3.15 $X2=0
+ $Y2=0
cc_936 N_A_876_119#_c_1302_n N_VPWR_c_1933_n 0.0060054f $X=6.225 $Y=3.15 $X2=0
+ $Y2=0
cc_937 N_A_876_119#_c_1304_n N_VPWR_c_1933_n 0.0968493f $X=10.995 $Y=3.15 $X2=0
+ $Y2=0
cc_938 N_A_876_119#_c_1306_n N_VPWR_c_1933_n 0.0154456f $X=8.04 $Y=3.15 $X2=0
+ $Y2=0
cc_939 N_A_876_119#_M1029_g N_VGND_c_2164_n 0.00456171f $X=5.67 $Y=0.805 $X2=0
+ $Y2=0
cc_940 N_A_876_119#_c_1293_n N_VGND_c_2164_n 0.00253443f $X=5.64 $Y=1.345 $X2=0
+ $Y2=0
cc_941 N_A_876_119#_c_1294_n N_VGND_c_2164_n 4.24337e-19 $X=5.64 $Y=1.345 $X2=0
+ $Y2=0
cc_942 N_A_876_119#_c_1292_n N_VGND_c_2170_n 0.0032269f $X=4.505 $Y=0.805 $X2=0
+ $Y2=0
cc_943 N_A_876_119#_M1020_g N_VGND_c_2171_n 0.00404693f $X=11.92 $Y=0.445 $X2=0
+ $Y2=0
cc_944 N_A_876_119#_c_1286_n N_VGND_c_2174_n 9.39239e-19 $X=5.67 $Y=1.18 $X2=0
+ $Y2=0
cc_945 N_A_876_119#_M1029_g N_VGND_c_2174_n 9.39239e-19 $X=5.67 $Y=0.805 $X2=0
+ $Y2=0
cc_946 N_A_876_119#_c_1289_n N_VGND_c_2174_n 9.39239e-19 $X=7.085 $Y=1.09 $X2=0
+ $Y2=0
cc_947 N_A_876_119#_M1020_g N_VGND_c_2174_n 0.00741786f $X=11.92 $Y=0.445 $X2=0
+ $Y2=0
cc_948 N_A_876_119#_c_1292_n N_VGND_c_2174_n 0.0044301f $X=4.505 $Y=0.805 $X2=0
+ $Y2=0
cc_949 N_A_2435_296#_c_1473_n N_A_2092_47#_c_1567_n 0.00456304f $X=14.025
+ $Y=0.402 $X2=0 $Y2=0
cc_950 N_A_2435_296#_c_1475_n N_A_2092_47#_c_1567_n 0.00433787f $X=14.11
+ $Y=1.265 $X2=0 $Y2=0
cc_951 N_A_2435_296#_c_1474_n N_A_2092_47#_M1004_g 0.0228622f $X=14.025 $Y=1.35
+ $X2=0 $Y2=0
cc_952 N_A_2435_296#_c_1475_n N_A_2092_47#_M1004_g 0.00987175f $X=14.11 $Y=1.265
+ $X2=0 $Y2=0
cc_953 N_A_2435_296#_c_1477_n N_A_2092_47#_M1004_g 7.97916e-19 $X=13.185
+ $Y=1.237 $X2=0 $Y2=0
cc_954 N_A_2435_296#_c_1499_n N_A_2092_47#_M1004_g 0.0201575f $X=13.66 $Y=2.28
+ $X2=0 $Y2=0
cc_955 N_A_2435_296#_c_1478_n N_A_2092_47#_M1004_g 0.0330617f $X=13.665 $Y=2.115
+ $X2=0 $Y2=0
cc_956 N_A_2435_296#_c_1479_n N_A_2092_47#_M1004_g 0.00407595f $X=13.75 $Y=1.35
+ $X2=0 $Y2=0
cc_957 N_A_2435_296#_c_1475_n N_A_2092_47#_c_1569_n 0.00950344f $X=14.11
+ $Y=1.265 $X2=0 $Y2=0
cc_958 N_A_2435_296#_c_1472_n N_A_2092_47#_c_1570_n 0.00379692f $X=13.665
+ $Y=1.35 $X2=0 $Y2=0
cc_959 N_A_2435_296#_c_1473_n N_A_2092_47#_c_1570_n 0.00725461f $X=14.025
+ $Y=0.402 $X2=0 $Y2=0
cc_960 N_A_2435_296#_c_1475_n N_A_2092_47#_c_1570_n 0.00565419f $X=14.11
+ $Y=1.265 $X2=0 $Y2=0
cc_961 N_A_2435_296#_c_1477_n N_A_2092_47#_c_1570_n 2.05952e-19 $X=13.185
+ $Y=1.237 $X2=0 $Y2=0
cc_962 N_A_2435_296#_c_1479_n N_A_2092_47#_c_1570_n 0.00328339f $X=13.75 $Y=1.35
+ $X2=0 $Y2=0
cc_963 N_A_2435_296#_c_1473_n N_A_2092_47#_c_1571_n 0.00365806f $X=14.025
+ $Y=0.402 $X2=0 $Y2=0
cc_964 N_A_2435_296#_c_1475_n N_A_2092_47#_c_1571_n 7.87769e-19 $X=14.11
+ $Y=1.265 $X2=0 $Y2=0
cc_965 N_A_2435_296#_M1003_g N_A_2092_47#_c_1585_n 0.0215213f $X=12.3 $Y=2.595
+ $X2=0 $Y2=0
cc_966 N_A_2435_296#_M1034_g N_A_2092_47#_c_1575_n 3.18306e-19 $X=12.46 $Y=0.445
+ $X2=0 $Y2=0
cc_967 N_A_2435_296#_M1003_g N_A_2092_47#_c_1576_n 0.0024687f $X=12.3 $Y=2.595
+ $X2=0 $Y2=0
cc_968 N_A_2435_296#_M1034_g N_A_2092_47#_c_1576_n 0.00890508f $X=12.46 $Y=0.445
+ $X2=0 $Y2=0
cc_969 N_A_2435_296#_c_1476_n N_A_2092_47#_c_1576_n 0.0235733f $X=13.015
+ $Y=1.237 $X2=0 $Y2=0
cc_970 N_A_2435_296#_c_1477_n N_A_2092_47#_c_1576_n 0.00211516f $X=13.185
+ $Y=1.237 $X2=0 $Y2=0
cc_971 N_A_2435_296#_c_1480_n N_A_2092_47#_c_1576_n 0.02592f $X=12.46 $Y=1.335
+ $X2=0 $Y2=0
cc_972 N_A_2435_296#_M1034_g N_A_2092_47#_c_1577_n 0.0105628f $X=12.46 $Y=0.445
+ $X2=0 $Y2=0
cc_973 N_A_2435_296#_c_1472_n N_A_2092_47#_c_1577_n 0.0127047f $X=13.665 $Y=1.35
+ $X2=0 $Y2=0
cc_974 N_A_2435_296#_c_1476_n N_A_2092_47#_c_1577_n 0.0404996f $X=13.015
+ $Y=1.237 $X2=0 $Y2=0
cc_975 N_A_2435_296#_c_1480_n N_A_2092_47#_c_1577_n 0.010622f $X=12.46 $Y=1.335
+ $X2=0 $Y2=0
cc_976 N_A_2435_296#_M1034_g N_A_2092_47#_c_1579_n 0.0139085f $X=12.46 $Y=0.445
+ $X2=0 $Y2=0
cc_977 N_A_2435_296#_c_1472_n N_A_2092_47#_c_1580_n 0.0108888f $X=13.665 $Y=1.35
+ $X2=0 $Y2=0
cc_978 N_A_2435_296#_c_1473_n N_A_2092_47#_c_1580_n 0.0105268f $X=14.025
+ $Y=0.402 $X2=0 $Y2=0
cc_979 N_A_2435_296#_c_1474_n N_A_2092_47#_c_1580_n 5.93443e-19 $X=14.025
+ $Y=1.35 $X2=0 $Y2=0
cc_980 N_A_2435_296#_c_1475_n N_A_2092_47#_c_1580_n 0.0282171f $X=14.11 $Y=1.265
+ $X2=0 $Y2=0
cc_981 N_A_2435_296#_c_1477_n N_A_2092_47#_c_1580_n 0.0020253f $X=13.185
+ $Y=1.237 $X2=0 $Y2=0
cc_982 N_A_2435_296#_c_1479_n N_A_2092_47#_c_1580_n 0.0138073f $X=13.75 $Y=1.35
+ $X2=0 $Y2=0
cc_983 N_A_2435_296#_c_1474_n N_A_2863_90#_c_1727_n 0.00886908f $X=14.025
+ $Y=1.35 $X2=0 $Y2=0
cc_984 N_A_2435_296#_c_1475_n N_A_2863_90#_c_1727_n 0.0162975f $X=14.11 $Y=1.265
+ $X2=0 $Y2=0
cc_985 N_A_2435_296#_c_1473_n N_A_2863_90#_c_1731_n 0.00651313f $X=14.025
+ $Y=0.402 $X2=0 $Y2=0
cc_986 N_A_2435_296#_c_1475_n N_A_2863_90#_c_1731_n 0.0283934f $X=14.11 $Y=1.265
+ $X2=0 $Y2=0
cc_987 N_A_2435_296#_M1003_g N_VPWR_c_1939_n 0.0261299f $X=12.3 $Y=2.595 $X2=0
+ $Y2=0
cc_988 N_A_2435_296#_c_1480_n N_VPWR_c_1939_n 0.00240483f $X=12.46 $Y=1.335
+ $X2=0 $Y2=0
cc_989 N_A_2435_296#_c_1474_n N_VPWR_c_1940_n 0.00602976f $X=14.025 $Y=1.35
+ $X2=0 $Y2=0
cc_990 N_A_2435_296#_c_1478_n N_VPWR_c_1940_n 0.0679117f $X=13.665 $Y=2.115
+ $X2=0 $Y2=0
cc_991 N_A_2435_296#_M1003_g N_VPWR_c_1947_n 0.008763f $X=12.3 $Y=2.595 $X2=0
+ $Y2=0
cc_992 N_A_2435_296#_c_1499_n N_VPWR_c_1952_n 0.0184348f $X=13.66 $Y=2.28 $X2=0
+ $Y2=0
cc_993 N_A_2435_296#_M1028_d N_VPWR_c_1933_n 0.00223819f $X=13.52 $Y=2.095 $X2=0
+ $Y2=0
cc_994 N_A_2435_296#_M1003_g N_VPWR_c_1933_n 0.0144563f $X=12.3 $Y=2.595 $X2=0
+ $Y2=0
cc_995 N_A_2435_296#_c_1499_n N_VPWR_c_1933_n 0.0126656f $X=13.66 $Y=2.28 $X2=0
+ $Y2=0
cc_996 N_A_2435_296#_M1034_g N_VGND_c_2167_n 0.0108659f $X=12.46 $Y=0.445 $X2=0
+ $Y2=0
cc_997 N_A_2435_296#_M1034_g N_VGND_c_2171_n 0.00420927f $X=12.46 $Y=0.445 $X2=0
+ $Y2=0
cc_998 N_A_2435_296#_c_1473_n N_VGND_c_2172_n 0.0266036f $X=14.025 $Y=0.402
+ $X2=0 $Y2=0
cc_999 N_A_2435_296#_M1027_d N_VGND_c_2174_n 0.0023412f $X=13.695 $Y=0.235 $X2=0
+ $Y2=0
cc_1000 N_A_2435_296#_M1034_g N_VGND_c_2174_n 0.00692543f $X=12.46 $Y=0.445
+ $X2=0 $Y2=0
cc_1001 N_A_2435_296#_c_1473_n N_VGND_c_2174_n 0.0193847f $X=14.025 $Y=0.402
+ $X2=0 $Y2=0
cc_1002 N_A_2092_47#_c_1574_n N_A_2863_90#_M1040_g 0.0175303f $X=15.035 $Y=0.945
+ $X2=0 $Y2=0
cc_1003 N_A_2092_47#_M1005_g N_A_2863_90#_M1007_g 0.0158144f $X=15.015 $Y=2.44
+ $X2=0 $Y2=0
cc_1004 N_A_2092_47#_c_1572_n N_A_2863_90#_c_1725_n 0.0220078f $X=15.015
+ $Y=1.095 $X2=0 $Y2=0
cc_1005 N_A_2092_47#_M1004_g N_A_2863_90#_c_1727_n 0.00510662f $X=13.925
+ $Y=2.595 $X2=0 $Y2=0
cc_1006 N_A_2092_47#_c_1569_n N_A_2863_90#_c_1727_n 0.00635851f $X=14.6 $Y=1.02
+ $X2=0 $Y2=0
cc_1007 N_A_2092_47#_c_1571_n N_A_2863_90#_c_1727_n 0.00246055f $X=14.675
+ $Y=0.945 $X2=0 $Y2=0
cc_1008 N_A_2092_47#_c_1572_n N_A_2863_90#_c_1727_n 0.00718303f $X=15.015
+ $Y=1.095 $X2=0 $Y2=0
cc_1009 N_A_2092_47#_M1005_g N_A_2863_90#_c_1727_n 0.0120439f $X=15.015 $Y=2.44
+ $X2=0 $Y2=0
cc_1010 N_A_2092_47#_c_1574_n N_A_2863_90#_c_1727_n 3.25852e-19 $X=15.035
+ $Y=0.945 $X2=0 $Y2=0
cc_1011 N_A_2092_47#_M1004_g N_A_2863_90#_c_1735_n 0.0109968f $X=13.925 $Y=2.595
+ $X2=0 $Y2=0
cc_1012 N_A_2092_47#_M1005_g N_A_2863_90#_c_1735_n 0.0259966f $X=15.015 $Y=2.44
+ $X2=0 $Y2=0
cc_1013 N_A_2092_47#_M1005_g N_A_2863_90#_c_1728_n 0.0240751f $X=15.015 $Y=2.44
+ $X2=0 $Y2=0
cc_1014 N_A_2092_47#_c_1572_n N_A_2863_90#_c_1729_n 0.00217928f $X=15.015
+ $Y=1.095 $X2=0 $Y2=0
cc_1015 N_A_2092_47#_M1005_g N_A_2863_90#_c_1730_n 0.0213924f $X=15.015 $Y=2.44
+ $X2=0 $Y2=0
cc_1016 N_A_2092_47#_c_1569_n N_A_2863_90#_c_1731_n 0.00762673f $X=14.6 $Y=1.02
+ $X2=0 $Y2=0
cc_1017 N_A_2092_47#_c_1571_n N_A_2863_90#_c_1731_n 0.0118067f $X=14.675
+ $Y=0.945 $X2=0 $Y2=0
cc_1018 N_A_2092_47#_c_1574_n N_A_2863_90#_c_1731_n 0.00142181f $X=15.035
+ $Y=0.945 $X2=0 $Y2=0
cc_1019 N_A_2092_47#_M1004_g N_A_2863_90#_c_1732_n 0.00527517f $X=13.925
+ $Y=2.595 $X2=0 $Y2=0
cc_1020 N_A_2092_47#_c_1572_n N_A_2863_90#_c_1732_n 0.00333566f $X=15.015
+ $Y=1.095 $X2=0 $Y2=0
cc_1021 N_A_2092_47#_M1005_g N_A_2863_90#_c_1732_n 0.00525478f $X=15.015 $Y=2.44
+ $X2=0 $Y2=0
cc_1022 N_A_2092_47#_c_1585_n N_VPWR_c_1939_n 0.00356713f $X=12.285 $Y=1.77
+ $X2=0 $Y2=0
cc_1023 N_A_2092_47#_M1004_g N_VPWR_c_1940_n 0.0239823f $X=13.925 $Y=2.595 $X2=0
+ $Y2=0
cc_1024 N_A_2092_47#_M1005_g N_VPWR_c_1940_n 0.00420908f $X=15.015 $Y=2.44 $X2=0
+ $Y2=0
cc_1025 N_A_2092_47#_M1005_g N_VPWR_c_1941_n 0.00817829f $X=15.015 $Y=2.44 $X2=0
+ $Y2=0
cc_1026 N_A_2092_47#_M1005_g N_VPWR_c_1942_n 0.0257173f $X=15.015 $Y=2.44 $X2=0
+ $Y2=0
cc_1027 N_A_2092_47#_c_1584_n N_VPWR_c_1947_n 0.0216625f $X=11.465 $Y=2.2 $X2=0
+ $Y2=0
cc_1028 N_A_2092_47#_M1004_g N_VPWR_c_1952_n 0.00825157f $X=13.925 $Y=2.595
+ $X2=0 $Y2=0
cc_1029 N_A_2092_47#_M1002_d N_VPWR_c_1933_n 0.00491311f $X=11.245 $Y=1.705
+ $X2=0 $Y2=0
cc_1030 N_A_2092_47#_M1004_g N_VPWR_c_1933_n 0.0132328f $X=13.925 $Y=2.595 $X2=0
+ $Y2=0
cc_1031 N_A_2092_47#_M1005_g N_VPWR_c_1933_n 0.00812777f $X=15.015 $Y=2.44 $X2=0
+ $Y2=0
cc_1032 N_A_2092_47#_c_1584_n N_VPWR_c_1933_n 0.0126859f $X=11.465 $Y=2.2 $X2=0
+ $Y2=0
cc_1033 N_A_2092_47#_M1005_g Q 2.7522e-19 $X=15.015 $Y=2.44 $X2=0 $Y2=0
cc_1034 N_A_2092_47#_c_1577_n N_VGND_c_2167_n 0.0245793f $X=13.515 $Y=0.775
+ $X2=0 $Y2=0
cc_1035 N_A_2092_47#_c_1579_n N_VGND_c_2167_n 3.54027e-19 $X=12.37 $Y=0.59 $X2=0
+ $Y2=0
cc_1036 N_A_2092_47#_c_1571_n N_VGND_c_2168_n 0.00174911f $X=14.675 $Y=0.945
+ $X2=0 $Y2=0
cc_1037 N_A_2092_47#_c_1572_n N_VGND_c_2168_n 0.00142058f $X=15.015 $Y=1.095
+ $X2=0 $Y2=0
cc_1038 N_A_2092_47#_c_1574_n N_VGND_c_2168_n 0.012411f $X=15.035 $Y=0.945 $X2=0
+ $Y2=0
cc_1039 N_A_2092_47#_c_1575_n N_VGND_c_2171_n 0.00982544f $X=12.285 $Y=0.59
+ $X2=0 $Y2=0
cc_1040 N_A_2092_47#_c_1577_n N_VGND_c_2171_n 0.0027733f $X=13.515 $Y=0.775
+ $X2=0 $Y2=0
cc_1041 N_A_2092_47#_c_1578_n N_VGND_c_2171_n 0.0193564f $X=11.675 $Y=0.47 $X2=0
+ $Y2=0
cc_1042 N_A_2092_47#_c_1579_n N_VGND_c_2171_n 0.0036116f $X=12.37 $Y=0.59 $X2=0
+ $Y2=0
cc_1043 N_A_2092_47#_c_1567_n N_VGND_c_2172_n 0.00421748f $X=13.62 $Y=0.765
+ $X2=0 $Y2=0
cc_1044 N_A_2092_47#_c_1571_n N_VGND_c_2172_n 0.00421717f $X=14.675 $Y=0.945
+ $X2=0 $Y2=0
cc_1045 N_A_2092_47#_c_1574_n N_VGND_c_2172_n 0.00432588f $X=15.035 $Y=0.945
+ $X2=0 $Y2=0
cc_1046 N_A_2092_47#_c_1577_n N_VGND_c_2172_n 0.00866747f $X=13.515 $Y=0.775
+ $X2=0 $Y2=0
cc_1047 N_A_2092_47#_c_1580_n N_VGND_c_2172_n 0.00241382f $X=13.68 $Y=0.775
+ $X2=0 $Y2=0
cc_1048 N_A_2092_47#_M1039_d N_VGND_c_2174_n 0.0199521f $X=10.46 $Y=0.235 $X2=0
+ $Y2=0
cc_1049 N_A_2092_47#_c_1567_n N_VGND_c_2174_n 0.00718403f $X=13.62 $Y=0.765
+ $X2=0 $Y2=0
cc_1050 N_A_2092_47#_c_1571_n N_VGND_c_2174_n 0.00520574f $X=14.675 $Y=0.945
+ $X2=0 $Y2=0
cc_1051 N_A_2092_47#_c_1574_n N_VGND_c_2174_n 0.00437282f $X=15.035 $Y=0.945
+ $X2=0 $Y2=0
cc_1052 N_A_2092_47#_c_1575_n N_VGND_c_2174_n 0.0132932f $X=12.285 $Y=0.59 $X2=0
+ $Y2=0
cc_1053 N_A_2092_47#_c_1577_n N_VGND_c_2174_n 0.0202802f $X=13.515 $Y=0.775
+ $X2=0 $Y2=0
cc_1054 N_A_2092_47#_c_1578_n N_VGND_c_2174_n 0.0125239f $X=11.675 $Y=0.47 $X2=0
+ $Y2=0
cc_1055 N_A_2092_47#_c_1579_n N_VGND_c_2174_n 0.00525158f $X=12.37 $Y=0.59 $X2=0
+ $Y2=0
cc_1056 N_A_2092_47#_c_1580_n N_VGND_c_2174_n 0.00411417f $X=13.68 $Y=0.775
+ $X2=0 $Y2=0
cc_1057 N_A_2092_47#_c_1575_n A_2399_47# 0.00402457f $X=12.285 $Y=0.59 $X2=-0.19
+ $Y2=-0.245
cc_1058 N_A_2092_47#_c_1579_n A_2399_47# 0.00102066f $X=12.37 $Y=0.59 $X2=-0.19
+ $Y2=-0.245
cc_1059 N_A_2863_90#_c_1735_n N_VPWR_c_1940_n 0.071546f $X=14.75 $Y=2.085 $X2=0
+ $Y2=0
cc_1060 N_A_2863_90#_c_1735_n N_VPWR_c_1941_n 0.0155423f $X=14.75 $Y=2.085 $X2=0
+ $Y2=0
cc_1061 N_A_2863_90#_M1007_g N_VPWR_c_1942_n 0.0257163f $X=15.545 $Y=2.44 $X2=0
+ $Y2=0
cc_1062 N_A_2863_90#_c_1726_n N_VPWR_c_1942_n 5.43851e-19 $X=15.515 $Y=1.74
+ $X2=0 $Y2=0
cc_1063 N_A_2863_90#_c_1735_n N_VPWR_c_1942_n 0.0692741f $X=14.75 $Y=2.085 $X2=0
+ $Y2=0
cc_1064 N_A_2863_90#_c_1728_n N_VPWR_c_1942_n 0.0266481f $X=15.35 $Y=1.655 $X2=0
+ $Y2=0
cc_1065 N_A_2863_90#_M1007_g N_VPWR_c_1953_n 0.00817829f $X=15.545 $Y=2.44 $X2=0
+ $Y2=0
cc_1066 N_A_2863_90#_M1007_g N_VPWR_c_1933_n 0.00812777f $X=15.545 $Y=2.44 $X2=0
+ $Y2=0
cc_1067 N_A_2863_90#_c_1735_n N_VPWR_c_1933_n 0.0137709f $X=14.75 $Y=2.085 $X2=0
+ $Y2=0
cc_1068 N_A_2863_90#_M1040_g Q 0.00214984f $X=15.465 $Y=0.66 $X2=0 $Y2=0
cc_1069 N_A_2863_90#_M1007_g Q 0.0067544f $X=15.545 $Y=2.44 $X2=0 $Y2=0
cc_1070 N_A_2863_90#_M1036_g Q 0.0157507f $X=15.825 $Y=0.66 $X2=0 $Y2=0
cc_1071 N_A_2863_90#_c_1725_n Q 0.00624049f $X=15.825 $Y=1.145 $X2=0 $Y2=0
cc_1072 N_A_2863_90#_c_1728_n Q 0.0128217f $X=15.35 $Y=1.655 $X2=0 $Y2=0
cc_1073 N_A_2863_90#_c_1729_n Q 0.035011f $X=15.515 $Y=1.235 $X2=0 $Y2=0
cc_1074 N_A_2863_90#_c_1730_n Q 0.00906243f $X=15.515 $Y=1.235 $X2=0 $Y2=0
cc_1075 N_A_2863_90#_M1007_g Q 0.0055764f $X=15.545 $Y=2.44 $X2=0 $Y2=0
cc_1076 N_A_2863_90#_c_1725_n Q 0.00547364f $X=15.825 $Y=1.145 $X2=0 $Y2=0
cc_1077 N_A_2863_90#_c_1728_n Q 0.00279016f $X=15.35 $Y=1.655 $X2=0 $Y2=0
cc_1078 N_A_2863_90#_M1007_g Q 0.013651f $X=15.545 $Y=2.44 $X2=0 $Y2=0
cc_1079 N_A_2863_90#_M1040_g N_VGND_c_2168_n 0.0122046f $X=15.465 $Y=0.66 $X2=0
+ $Y2=0
cc_1080 N_A_2863_90#_M1036_g N_VGND_c_2168_n 0.00180376f $X=15.825 $Y=0.66 $X2=0
+ $Y2=0
cc_1081 N_A_2863_90#_c_1725_n N_VGND_c_2168_n 3.03142e-19 $X=15.825 $Y=1.145
+ $X2=0 $Y2=0
cc_1082 N_A_2863_90#_c_1729_n N_VGND_c_2168_n 0.00526295f $X=15.515 $Y=1.235
+ $X2=0 $Y2=0
cc_1083 N_A_2863_90#_c_1731_n N_VGND_c_2168_n 0.0180446f $X=14.62 $Y=0.66 $X2=0
+ $Y2=0
cc_1084 N_A_2863_90#_c_1731_n N_VGND_c_2172_n 0.0105165f $X=14.62 $Y=0.66 $X2=0
+ $Y2=0
cc_1085 N_A_2863_90#_M1040_g N_VGND_c_2173_n 0.00432588f $X=15.465 $Y=0.66 $X2=0
+ $Y2=0
cc_1086 N_A_2863_90#_M1036_g N_VGND_c_2173_n 0.00497955f $X=15.825 $Y=0.66 $X2=0
+ $Y2=0
cc_1087 N_A_2863_90#_M1040_g N_VGND_c_2174_n 0.00437282f $X=15.465 $Y=0.66 $X2=0
+ $Y2=0
cc_1088 N_A_2863_90#_M1036_g N_VGND_c_2174_n 0.00520574f $X=15.825 $Y=0.66 $X2=0
+ $Y2=0
cc_1089 N_A_2863_90#_c_1731_n N_VGND_c_2174_n 0.0113047f $X=14.62 $Y=0.66 $X2=0
+ $Y2=0
cc_1090 N_A_116_419#_c_1805_n A_223_419# 0.00392987f $X=2.69 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_1091 N_A_116_419#_c_1805_n N_VPWR_M1018_d 0.00484953f $X=2.69 $Y=2.395
+ $X2=-0.19 $Y2=-0.245
cc_1092 N_A_116_419#_c_1806_n N_VPWR_M1009_d 0.00651692f $X=3.73 $Y=2.59 $X2=0
+ $Y2=0
cc_1093 N_A_116_419#_c_1800_n N_VPWR_M1031_d 0.014726f $X=6.865 $Y=2.545 $X2=0
+ $Y2=0
cc_1094 N_A_116_419#_c_1805_n N_VPWR_c_1934_n 0.01888f $X=2.69 $Y=2.395 $X2=0
+ $Y2=0
cc_1095 N_A_116_419#_c_1806_n N_VPWR_c_1935_n 0.0196062f $X=3.73 $Y=2.59 $X2=0
+ $Y2=0
cc_1096 N_A_116_419#_c_1835_n N_VPWR_c_1935_n 0.00279982f $X=3.815 $Y=2.895
+ $X2=0 $Y2=0
cc_1097 N_A_116_419#_c_1836_n N_VPWR_c_1935_n 0.0133991f $X=3.9 $Y=2.98 $X2=0
+ $Y2=0
cc_1098 N_A_116_419#_c_1818_n N_VPWR_c_1935_n 0.013837f $X=2.855 $Y=2.59 $X2=0
+ $Y2=0
cc_1099 N_A_116_419#_c_1799_n N_VPWR_c_1936_n 0.00800521f $X=4.84 $Y=2.98 $X2=0
+ $Y2=0
cc_1100 N_A_116_419#_c_1800_n N_VPWR_c_1936_n 0.0198761f $X=6.865 $Y=2.545 $X2=0
+ $Y2=0
cc_1101 N_A_116_419#_c_1806_n N_VPWR_c_1943_n 0.00310989f $X=3.73 $Y=2.59 $X2=0
+ $Y2=0
cc_1102 N_A_116_419#_c_1818_n N_VPWR_c_1943_n 0.0177952f $X=2.855 $Y=2.59 $X2=0
+ $Y2=0
cc_1103 N_A_116_419#_c_1806_n N_VPWR_c_1945_n 0.00243537f $X=3.73 $Y=2.59 $X2=0
+ $Y2=0
cc_1104 N_A_116_419#_c_1799_n N_VPWR_c_1945_n 0.0668459f $X=4.84 $Y=2.98 $X2=0
+ $Y2=0
cc_1105 N_A_116_419#_c_1836_n N_VPWR_c_1945_n 0.00953977f $X=3.9 $Y=2.98 $X2=0
+ $Y2=0
cc_1106 N_A_116_419#_c_1800_n N_VPWR_c_1945_n 0.00242368f $X=6.865 $Y=2.545
+ $X2=0 $Y2=0
cc_1107 N_A_116_419#_c_1803_n N_VPWR_c_1949_n 0.0514475f $X=0.725 $Y=2.24 $X2=0
+ $Y2=0
cc_1108 N_A_116_419#_c_1800_n N_VPWR_c_1950_n 0.0202786f $X=6.865 $Y=2.545 $X2=0
+ $Y2=0
cc_1109 N_A_116_419#_c_1801_n N_VPWR_c_1950_n 0.00391376f $X=6.95 $Y=2.46 $X2=0
+ $Y2=0
cc_1110 N_A_116_419#_M1001_s N_VPWR_c_1933_n 0.0023218f $X=0.58 $Y=2.095 $X2=0
+ $Y2=0
cc_1111 N_A_116_419#_M1030_d N_VPWR_c_1933_n 0.00223819f $X=2.715 $Y=2.095 $X2=0
+ $Y2=0
cc_1112 N_A_116_419#_c_1805_n N_VPWR_c_1933_n 0.0448219f $X=2.69 $Y=2.395 $X2=0
+ $Y2=0
cc_1113 N_A_116_419#_c_1806_n N_VPWR_c_1933_n 0.0106001f $X=3.73 $Y=2.59 $X2=0
+ $Y2=0
cc_1114 N_A_116_419#_c_1799_n N_VPWR_c_1933_n 0.0405319f $X=4.84 $Y=2.98 $X2=0
+ $Y2=0
cc_1115 N_A_116_419#_c_1836_n N_VPWR_c_1933_n 0.00594499f $X=3.9 $Y=2.98 $X2=0
+ $Y2=0
cc_1116 N_A_116_419#_c_1800_n N_VPWR_c_1933_n 0.0384392f $X=6.865 $Y=2.545 $X2=0
+ $Y2=0
cc_1117 N_A_116_419#_c_1801_n N_VPWR_c_1933_n 0.00471658f $X=6.95 $Y=2.46 $X2=0
+ $Y2=0
cc_1118 N_A_116_419#_c_1803_n N_VPWR_c_1933_n 0.0306938f $X=0.725 $Y=2.24 $X2=0
+ $Y2=0
cc_1119 N_A_116_419#_c_1818_n N_VPWR_c_1933_n 0.0123247f $X=2.855 $Y=2.59 $X2=0
+ $Y2=0
cc_1120 N_A_116_419#_c_1805_n A_439_419# 0.00483281f $X=2.69 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_1121 N_A_116_419#_c_1793_n N_noxref_23_M1000_s 0.00142f $X=0.26 $Y=0.705
+ $X2=-0.19 $Y2=-0.245
cc_1122 N_A_116_419#_c_1796_n N_noxref_23_M1000_s 0.00114695f $X=0.49 $Y=2.075
+ $X2=-0.19 $Y2=-0.245
cc_1123 N_A_116_419#_c_1813_n N_noxref_23_M1000_s 0.00993657f $X=1.15 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_1124 N_A_116_419#_c_1797_n N_noxref_23_c_2134_n 0.0224537f $X=1.315 $Y=0.78
+ $X2=0 $Y2=0
cc_1125 N_A_116_419#_c_1813_n N_noxref_23_c_2134_n 0.0338842f $X=1.15 $Y=0.74
+ $X2=0 $Y2=0
cc_1126 N_A_116_419#_c_1797_n N_noxref_23_c_2135_n 0.00349227f $X=1.315 $Y=0.78
+ $X2=0 $Y2=0
cc_1127 N_A_116_419#_c_1793_n N_noxref_23_c_2136_n 0.00661621f $X=0.26 $Y=0.705
+ $X2=0 $Y2=0
cc_1128 N_A_116_419#_c_1813_n N_noxref_23_c_2136_n 0.0156512f $X=1.15 $Y=0.74
+ $X2=0 $Y2=0
cc_1129 N_A_116_419#_c_1813_n noxref_24 0.00310318f $X=1.15 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_1130 N_A_116_419#_c_1794_n N_VGND_c_2165_n 0.00625348f $X=6.87 $Y=0.79 $X2=0
+ $Y2=0
cc_1131 N_A_116_419#_c_1793_n N_VGND_c_2169_n 0.00167184f $X=0.26 $Y=0.705 $X2=0
+ $Y2=0
cc_1132 N_A_116_419#_c_1793_n N_VGND_c_2174_n 0.00270497f $X=0.26 $Y=0.705 $X2=0
+ $Y2=0
cc_1133 N_A_116_419#_c_1794_n N_VGND_c_2174_n 0.00886387f $X=6.87 $Y=0.79 $X2=0
+ $Y2=0
cc_1134 A_223_419# N_VPWR_c_1933_n 0.00355777f $X=1.115 $Y=2.095 $X2=0 $Y2=0
cc_1135 N_VPWR_c_1933_n A_439_419# 0.00400249f $X=16.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1136 N_VPWR_c_1933_n A_2387_419# 0.010279f $X=16.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1137 N_VPWR_c_1942_n Q 0.0713761f $X=15.28 $Y=2.085 $X2=0 $Y2=0
cc_1138 N_VPWR_c_1953_n Q 0.0229765f $X=16.08 $Y=3.33 $X2=0 $Y2=0
cc_1139 N_VPWR_c_1933_n Q 0.0203382f $X=16.08 $Y=3.33 $X2=0 $Y2=0
cc_1140 Q N_VGND_c_2168_n 0.0153904f $X=15.995 $Y=0.47 $X2=0 $Y2=0
cc_1141 Q N_VGND_c_2173_n 0.0109928f $X=15.995 $Y=0.47 $X2=0 $Y2=0
cc_1142 Q N_VGND_c_2174_n 0.01149f $X=15.995 $Y=0.47 $X2=0 $Y2=0
cc_1143 N_noxref_23_c_2134_n N_VGND_c_2163_n 0.0136607f $X=2.05 $Y=0.35 $X2=0
+ $Y2=0
cc_1144 N_noxref_23_c_2135_n N_VGND_c_2163_n 0.0168326f $X=2.215 $Y=0.65 $X2=0
+ $Y2=0
cc_1145 N_noxref_23_c_2134_n N_VGND_c_2169_n 0.0219978f $X=2.05 $Y=0.35 $X2=0
+ $Y2=0
cc_1146 N_noxref_23_c_2136_n N_VGND_c_2169_n 0.113679f $X=0.5 $Y=0.352 $X2=0
+ $Y2=0
cc_1147 N_noxref_23_M1000_s N_VGND_c_2174_n 0.00272517f $X=0.19 $Y=0.205 $X2=0
+ $Y2=0
cc_1148 N_noxref_23_c_2134_n N_VGND_c_2174_n 0.012619f $X=2.05 $Y=0.35 $X2=0
+ $Y2=0
cc_1149 N_noxref_23_c_2136_n N_VGND_c_2174_n 0.070261f $X=0.5 $Y=0.352 $X2=0
+ $Y2=0
cc_1150 N_VGND_c_2174_n A_1900_47# 0.0027565f $X=16.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1151 N_VGND_c_2174_n A_2399_47# 0.00384968f $X=16.08 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1152 N_VGND_c_2174_n A_2661_47# 0.00297087f $X=16.08 $Y=0 $X2=-0.19
+ $Y2=-0.245
