* File: sky130_fd_sc_lp__a31oi_2.pex.spice
* Created: Wed Sep  2 09:27:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31OI_2%A3 1 3 6 8 10 12 15 17 18 25
r47 24 25 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.46
+ $X2=0.55 $Y2=1.46
r48 21 24 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.29 $Y=1.46
+ $X2=0.475 $Y2=1.46
r49 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.46 $X2=0.29 $Y2=1.46
r50 18 22 5.20967 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=1.295
+ $X2=0.272 $Y2=1.46
r51 13 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.445
+ $X2=0.905 $Y2=1.37
r52 13 15 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=0.905 $Y=1.445
+ $X2=0.905 $Y2=2.465
r53 10 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.295
+ $X2=0.905 $Y2=1.37
r54 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.905 $Y=1.295
+ $X2=0.905 $Y2=0.765
r55 8 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.37
+ $X2=0.905 $Y2=1.37
r56 8 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.37 $X2=0.55
+ $Y2=1.37
r57 4 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.625
+ $X2=0.475 $Y2=1.46
r58 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.475 $Y=1.625
+ $X2=0.475 $Y2=2.465
r59 1 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=1.46
r60 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_2%A2 1 3 6 8 10 13 15 16 23 25
c56 13 0 9.82587e-20 $X=1.845 $Y=2.465
c57 8 0 1.95662e-19 $X=1.765 $Y=1.295
r58 24 25 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=1.765 $Y=1.46
+ $X2=1.845 $Y2=1.46
r59 22 24 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=1.47 $Y=1.46
+ $X2=1.765 $Y2=1.46
r60 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.47
+ $Y=1.46 $X2=1.47 $Y2=1.46
r61 19 22 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.335 $Y=1.46
+ $X2=1.47 $Y2=1.46
r62 16 23 9.28835 $w=3.33e-07 $l=2.7e-07 $layer=LI1_cond $X=1.2 $Y=1.377
+ $X2=1.47 $Y2=1.377
r63 15 16 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.377
+ $X2=1.2 $Y2=1.377
r64 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.625
+ $X2=1.845 $Y2=1.46
r65 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.845 $Y=1.625
+ $X2=1.845 $Y2=2.465
r66 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.295
+ $X2=1.765 $Y2=1.46
r67 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.765 $Y=1.295
+ $X2=1.765 $Y2=0.765
r68 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.625
+ $X2=1.335 $Y2=1.46
r69 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.335 $Y=1.625
+ $X2=1.335 $Y2=2.465
r70 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.295
+ $X2=1.335 $Y2=1.46
r71 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.335 $Y=1.295
+ $X2=1.335 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_2%A1 3 5 6 9 11 15 19 21 22 24 28
c66 11 0 1.74935e-19 $X=3.005 $Y=1.42
r67 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.51
+ $X2=3.17 $Y2=1.675
r68 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.51 $X2=3.17 $Y2=1.51
r69 24 27 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.17 $Y=1.42 $X2=3.17
+ $Y2=1.51
r70 24 25 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.17 $Y=1.42 $X2=3.17
+ $Y2=1.345
r71 22 28 4.76343 $w=3.73e-07 $l=1.55e-07 $layer=LI1_cond $X=3.147 $Y=1.665
+ $X2=3.147 $Y2=1.51
r72 19 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.225 $Y=2.465
+ $X2=3.225 $Y2=1.675
r73 15 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.225 $Y=0.765
+ $X2=3.225 $Y2=1.345
r74 12 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.795 $Y=1.42
+ $X2=2.72 $Y2=1.42
r75 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.005 $Y=1.42
+ $X2=3.17 $Y2=1.42
r76 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.005 $Y=1.42
+ $X2=2.795 $Y2=1.42
r77 7 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.72 $Y=1.345
+ $X2=2.72 $Y2=1.42
r78 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.72 $Y=1.345 $X2=2.72
+ $Y2=0.765
r79 5 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.645 $Y=1.42
+ $X2=2.72 $Y2=1.42
r80 5 6 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.645 $Y=1.42
+ $X2=2.35 $Y2=1.42
r81 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.275 $Y=1.495
+ $X2=2.35 $Y2=1.42
r82 1 3 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.275 $Y=1.495
+ $X2=2.275 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_2%B1 3 7 11 15 17 18 19 28
r44 26 28 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.995 $Y=1.51
+ $X2=4.085 $Y2=1.51
r45 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.995
+ $Y=1.51 $X2=3.995 $Y2=1.51
r46 23 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.655 $Y=1.51
+ $X2=3.995 $Y2=1.51
r47 18 19 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.56 $Y2=1.587
r48 18 27 3.01408 $w=3.23e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=3.995 $Y2=1.587
r49 17 27 14.0066 $w=3.23e-07 $l=3.95e-07 $layer=LI1_cond $X=3.6 $Y=1.587
+ $X2=3.995 $Y2=1.587
r50 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.085 $Y=1.675
+ $X2=4.085 $Y2=1.51
r51 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.085 $Y=1.675
+ $X2=4.085 $Y2=2.465
r52 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.085 $Y=1.345
+ $X2=4.085 $Y2=1.51
r53 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.085 $Y=1.345
+ $X2=4.085 $Y2=0.765
r54 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.675
+ $X2=3.655 $Y2=1.51
r55 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.655 $Y=1.675
+ $X2=3.655 $Y2=2.465
r56 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.345
+ $X2=3.655 $Y2=1.51
r57 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.655 $Y=1.345
+ $X2=3.655 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_2%A_27_367# 1 2 3 4 5 18 22 23 26 30 38 40 42
+ 43 44 46 48 50
r61 44 54 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.335 $Y=2.905
+ $X2=4.335 $Y2=2.99
r62 44 46 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=4.335 $Y=2.905
+ $X2=4.335 $Y2=2.085
r63 42 54 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.205 $Y=2.99
+ $X2=4.335 $Y2=2.99
r64 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.205 $Y=2.99
+ $X2=3.535 $Y2=2.99
r65 41 43 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.44 $Y=2.905
+ $X2=3.535 $Y2=2.99
r66 40 52 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=2.47 $X2=3.44
+ $Y2=2.385
r67 40 41 25.3923 $w=1.88e-07 $l=4.35e-07 $layer=LI1_cond $X=3.44 $Y=2.47
+ $X2=3.44 $Y2=2.905
r68 39 50 2.45049 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=2.165 $Y=2.385
+ $X2=2.047 $Y2=2.385
r69 38 52 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.345 $Y=2.385
+ $X2=3.44 $Y2=2.385
r70 38 39 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=3.345 $Y=2.385
+ $X2=2.165 $Y2=2.385
r71 33 50 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.047 $Y=2.3
+ $X2=2.047 $Y2=2.385
r72 33 35 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.047 $Y=2.3
+ $X2=2.047 $Y2=1.96
r73 32 35 3.67801 $w=2.33e-07 $l=7.5e-08 $layer=LI1_cond $X=2.047 $Y=1.885
+ $X2=2.047 $Y2=1.96
r74 31 48 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=1.26 $Y=1.8
+ $X2=1.142 $Y2=1.8
r75 30 32 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=1.93 $Y=1.8
+ $X2=2.047 $Y2=1.885
r76 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.93 $Y=1.8 $X2=1.26
+ $Y2=1.8
r77 26 28 45.6073 $w=2.33e-07 $l=9.3e-07 $layer=LI1_cond $X=1.142 $Y=1.98
+ $X2=1.142 $Y2=2.91
r78 24 48 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.142 $Y=1.885
+ $X2=1.142 $Y2=1.8
r79 24 26 4.65881 $w=2.33e-07 $l=9.5e-08 $layer=LI1_cond $X=1.142 $Y=1.885
+ $X2=1.142 $Y2=1.98
r80 22 48 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=1.025 $Y=1.8
+ $X2=1.142 $Y2=1.8
r81 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=1.8
+ $X2=0.355 $Y2=1.8
r82 18 20 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.225 $Y=1.98
+ $X2=0.225 $Y2=2.91
r83 16 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=1.885
+ $X2=0.355 $Y2=1.8
r84 16 18 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=0.225 $Y=1.885
+ $X2=0.225 $Y2=1.98
r85 5 54 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=1.835 $X2=4.3 $Y2=2.91
r86 5 46 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=1.835 $X2=4.3 $Y2=2.085
r87 4 52 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=3.3
+ $Y=1.835 $X2=3.44 $Y2=2.465
r88 3 50 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=2.465
r89 3 35 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=1.96
r90 2 28 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.91
r91 2 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=1.98
r92 1 20 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r93 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_2%VPWR 1 2 3 12 18 23 24 25 27 42 43 46 51 57
r64 55 57 9.58177 $w=7.73e-07 $l=5.5e-08 $layer=LI1_cond $X=3.12 $Y=3.027
+ $X2=3.175 $Y2=3.027
r65 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 53 55 1.69766 $w=7.73e-07 $l=1.1e-07 $layer=LI1_cond $X=3.01 $Y=3.027
+ $X2=3.12 $Y2=3.027
r67 50 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 49 53 5.71031 $w=7.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=3.027
+ $X2=3.01 $Y2=3.027
r69 49 51 13.5944 $w=7.73e-07 $l=3.15e-07 $layer=LI1_cond $X=2.64 $Y=3.027
+ $X2=2.325 $Y2=3.027
r70 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 43 56 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 42 57 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=3.175 $Y2=3.33
r74 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 38 51 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.325 $Y2=3.33
r76 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 35 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 35 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r80 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r81 32 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r82 30 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r84 27 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r85 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r86 25 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 25 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r88 23 34 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.43 $Y=3.33 $X2=1.2
+ $Y2=3.33
r89 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.43 $Y=3.33
+ $X2=1.595 $Y2=3.33
r90 22 38 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.76 $Y=3.33 $X2=2.16
+ $Y2=3.33
r91 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.76 $Y=3.33
+ $X2=1.595 $Y2=3.33
r92 18 21 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=1.595 $Y=2.14
+ $X2=1.595 $Y2=2.95
r93 16 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.595 $Y=3.245
+ $X2=1.595 $Y2=3.33
r94 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.595 $Y=3.245
+ $X2=1.595 $Y2=2.95
r95 12 15 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=0.69 $Y=2.14
+ $X2=0.69 $Y2=2.95
r96 10 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r97 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.95
r98 3 53 300 $w=1.7e-07 $l=1.2212e-06 $layer=licon1_PDIFF $count=2 $X=2.35
+ $Y=1.835 $X2=3.01 $Y2=2.77
r99 2 21 400 $w=1.7e-07 $l=1.20395e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.595 $Y2=2.95
r100 2 18 400 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.595 $Y2=2.14
r101 1 15 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.95
r102 1 12 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.14
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_2%Y 1 2 3 4 15 17 19 23 25 31 34 35 37 38 39
c76 38 0 9.82587e-20 $X=2.64 $Y=1.665
c77 19 0 1.74935e-19 $X=3.705 $Y=2.04
c78 17 0 1.00242e-19 $X=3.345 $Y=1.17
r79 38 39 6.36053 $w=6.23e-07 $l=2.85e-07 $layer=LI1_cond $X=2.562 $Y=1.665
+ $X2=2.562 $Y2=1.95
r80 33 38 10.7778 $w=4.53e-07 $l=4.1e-07 $layer=LI1_cond $X=2.562 $Y=1.255
+ $X2=2.562 $Y2=1.665
r81 33 34 2.43256 $w=3.97e-07 $l=8.5e-08 $layer=LI1_cond $X=2.562 $Y=1.255
+ $X2=2.562 $Y2=1.17
r82 29 31 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=4.335 $Y=1.085
+ $X2=4.335 $Y2=0.49
r83 26 35 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.535 $Y=1.17
+ $X2=3.44 $Y2=1.17
r84 25 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.205 $Y=1.17
+ $X2=4.335 $Y2=1.085
r85 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.205 $Y=1.17
+ $X2=3.535 $Y2=1.17
r86 21 35 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=1.085
+ $X2=3.44 $Y2=1.17
r87 21 23 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=3.44 $Y=1.085
+ $X2=3.44 $Y2=0.49
r88 20 39 6.18715 $w=1.8e-07 $l=2.28e-07 $layer=LI1_cond $X=2.79 $Y=2.04
+ $X2=2.562 $Y2=2.04
r89 19 37 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=2.04
+ $X2=3.87 $Y2=2.04
r90 19 20 56.3788 $w=1.78e-07 $l=9.15e-07 $layer=LI1_cond $X=3.705 $Y=2.04
+ $X2=2.79 $Y2=2.04
r91 18 34 4.51935 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=2.79 $Y=1.17
+ $X2=2.562 $Y2=1.17
r92 17 35 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.345 $Y=1.17
+ $X2=3.44 $Y2=1.17
r93 17 18 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.345 $Y=1.17
+ $X2=2.79 $Y2=1.17
r94 13 34 2.43256 $w=3.97e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.505 $Y=1.085
+ $X2=2.562 $Y2=1.17
r95 13 15 13.3887 $w=3.38e-07 $l=3.95e-07 $layer=LI1_cond $X=2.505 $Y=1.085
+ $X2=2.505 $Y2=0.69
r96 4 37 300 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=2 $X=3.73
+ $Y=1.835 $X2=3.87 $Y2=2.055
r97 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.16
+ $Y=0.345 $X2=4.3 $Y2=0.49
r98 2 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.3
+ $Y=0.345 $X2=3.44 $Y2=0.49
r99 1 15 91 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=2 $X=2.375
+ $Y=0.345 $X2=2.5 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_2%A_27_69# 1 2 3 10 12 14 18 20 25 27
r42 27 29 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.98 $Y=0.7
+ $X2=1.98 $Y2=0.955
r43 21 25 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.255 $Y=0.955
+ $X2=1.14 $Y2=0.955
r44 20 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0.955
+ $X2=1.98 $Y2=0.955
r45 20 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.815 $Y=0.955
+ $X2=1.255 $Y2=0.955
r46 16 25 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.87
+ $X2=1.14 $Y2=0.955
r47 16 18 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.14 $Y=0.87
+ $X2=1.14 $Y2=0.5
r48 15 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.345 $Y=0.955
+ $X2=0.22 $Y2=0.955
r49 14 25 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.025 $Y=0.955
+ $X2=1.14 $Y2=0.955
r50 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.025 $Y=0.955
+ $X2=0.345 $Y2=0.955
r51 10 23 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.22 $Y=0.87 $X2=0.22
+ $Y2=0.955
r52 10 12 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.87
+ $X2=0.22 $Y2=0.5
r53 3 27 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.345 $X2=1.98 $Y2=0.7
r54 2 25 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.345 $X2=1.12 $Y2=0.955
r55 2 18 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.345 $X2=1.12 $Y2=0.5
r56 1 23 182 $w=1.7e-07 $l=6.69589e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.345 $X2=0.26 $Y2=0.955
r57 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.345 $X2=0.26 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_2%VGND 1 2 9 13 16 17 18 20 33 34 37
r52 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r54 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r55 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r56 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r57 27 30 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r58 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r60 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r61 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r62 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r64 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r65 18 31 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.6
+ $Y2=0
r66 18 28 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r67 16 30 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.6
+ $Y2=0
r68 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.87
+ $Y2=0
r69 15 33 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.035 $Y=0 $X2=4.56
+ $Y2=0
r70 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=0 $X2=3.87
+ $Y2=0
r71 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=0.085
+ $X2=3.87 $Y2=0
r72 11 13 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.87 $Y=0.085
+ $X2=3.87 $Y2=0.47
r73 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r74 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0.575
r75 2 13 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.73
+ $Y=0.345 $X2=3.87 $Y2=0.47
r76 1 9 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.345 $X2=0.69 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_2%A_282_69# 1 2 7 11 13
c26 13 0 1.95662e-19 $X=1.535 $Y=0.345
c27 7 0 1.00242e-19 $X=2.845 $Y=0.345
r28 13 16 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=1.535 $Y=0.345
+ $X2=1.535 $Y2=0.535
r29 9 11 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=3.01 $Y=0.435
+ $X2=3.01 $Y2=0.47
r30 8 13 1.91462 $w=1.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.645 $Y=0.345
+ $X2=1.535 $Y2=0.345
r31 7 9 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.845 $Y=0.345
+ $X2=3.01 $Y2=0.435
r32 7 8 73.9394 $w=1.78e-07 $l=1.2e-06 $layer=LI1_cond $X=2.845 $Y=0.345
+ $X2=1.645 $Y2=0.345
r33 2 11 91 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=2 $X=2.795
+ $Y=0.345 $X2=3.01 $Y2=0.47
r34 1 16 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.345 $X2=1.55 $Y2=0.535
.ends

