* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a22o_lp A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_137_409# B2 a_243_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_243_409# B1 a_137_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_225_47# B1 a_243_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_243_409# a_606_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_243_409# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_243_409# A1 a_389_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR A1 a_137_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_389_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_137_409# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_606_47# a_243_409# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
