# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a21oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a21oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.205000 1.355000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.295000 0.455000 1.605000 ;
        RECT 0.125000 1.605000 1.870000 1.675000 ;
        RECT 0.125000 1.675000 1.765000 1.785000 ;
        RECT 1.525000 1.345000 1.870000 1.605000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.040000 1.425000 2.800000 1.760000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.823200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 0.595000 1.260000 0.865000 ;
        RECT 1.025000 0.865000 2.545000 1.005000 ;
        RECT 1.025000 1.005000 3.275000 1.035000 ;
        RECT 2.285000 1.930000 3.275000 2.100000 ;
        RECT 2.285000 2.100000 2.615000 2.735000 ;
        RECT 2.335000 0.255000 2.545000 0.865000 ;
        RECT 2.345000 1.035000 3.275000 1.175000 ;
        RECT 2.970000 1.175000 3.275000 1.930000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.095000  0.085000 0.355000 1.095000 ;
      RECT 0.095000  1.955000 2.115000 2.125000 ;
      RECT 0.095000  2.125000 0.355000 3.075000 ;
      RECT 0.525000  0.255000 1.665000 0.425000 ;
      RECT 0.525000  0.425000 0.855000 1.035000 ;
      RECT 0.525000  2.295000 0.855000 3.245000 ;
      RECT 1.025000  2.125000 1.235000 3.075000 ;
      RECT 1.405000  2.295000 1.735000 3.245000 ;
      RECT 1.430000  0.425000 1.665000 0.695000 ;
      RECT 1.835000  0.085000 2.165000 0.695000 ;
      RECT 1.905000  2.125000 2.115000 2.905000 ;
      RECT 1.905000  2.905000 3.045000 3.075000 ;
      RECT 2.715000  0.085000 3.045000 0.835000 ;
      RECT 2.785000  2.270000 3.045000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__a21oi_2
END LIBRARY
