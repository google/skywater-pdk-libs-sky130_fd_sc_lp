* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfrtp_lp2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_141_88# D a_116_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_116_419# a_1147_408# a_1432_119# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VPWR RESET_B a_2435_296# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_1635_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_116_419# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_2387_419# a_2435_296# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_2863_90# a_2092_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_1432_119# a_876_119# a_1633_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_959_119# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1432_119# a_1147_408# a_1561_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_876_119# CLK a_959_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1900_47# a_1432_119# a_1605_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_116_419# D a_223_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 VPWR a_876_119# a_1147_408# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VGND a_1432_119# a_1900_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_2863_90# a_3108_90# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_223_419# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_876_119# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X18 a_116_419# SCE a_337_88# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1149_119# a_876_119# a_1147_408# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR RESET_B a_1432_119# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 a_439_419# a_81_194# a_116_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_1605_93# a_876_119# a_2092_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X23 a_337_88# SCD a_38_41# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_697_119# SCE a_81_194# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_38_41# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND a_876_119# a_1149_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_2863_90# a_2092_47# a_2950_90# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_2661_47# a_2092_47# a_2435_296# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_2950_90# a_2092_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_38_41# a_81_194# a_141_88# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VPWR a_1432_119# a_1605_93# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X32 a_1633_347# a_1605_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X33 VGND SCE a_697_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1561_119# a_1605_93# a_1635_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VGND RESET_B a_2661_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VPWR SCE a_81_194# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X37 VPWR a_2863_90# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X38 a_2092_47# a_876_119# a_2399_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VPWR SCD a_439_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X40 a_2435_296# a_2092_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X41 a_116_419# a_876_119# a_1432_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_1605_93# a_1147_408# a_2092_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 a_3108_90# a_2863_90# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_2399_47# a_2435_296# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 a_2092_47# a_1147_408# a_2387_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
