* NGSPICE file created from sky130_fd_sc_lp__o21ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_29_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=4.578e+11p pd=4.45e+06u as=3.192e+11p ps=2.44e+06u
M1001 Y A2 a_112_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=5.67e+11p pd=3.42e+06u as=2.646e+11p ps=2.94e+06u
M1002 a_112_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=6.678e+11p ps=6.1e+06u
M1003 VGND A1 a_29_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B1 a_29_47# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
.ends

