* NGSPICE file created from sky130_fd_sc_lp__inv_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__inv_1 A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=2.226e+11p ps=2.21e+06u
M1001 Y A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=3.339e+11p ps=3.05e+06u
.ends

