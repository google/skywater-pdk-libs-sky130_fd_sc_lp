* File: sky130_fd_sc_lp__ebufn_lp2.pxi.spice
* Created: Wed Sep  2 09:51:05 2020
* 
x_PM_SKY130_FD_SC_LP__EBUFN_LP2%A N_A_c_69_n N_A_M1001_g N_A_M1000_g N_A_M1007_g
+ N_A_c_71_n N_A_c_72_n A A A N_A_c_74_n PM_SKY130_FD_SC_LP__EBUFN_LP2%A
x_PM_SKY130_FD_SC_LP__EBUFN_LP2%A_27_47# N_A_27_47#_M1001_s N_A_27_47#_M1000_s
+ N_A_27_47#_c_109_n N_A_27_47#_c_110_n N_A_27_47#_M1003_g N_A_27_47#_M1004_g
+ N_A_27_47#_c_113_n N_A_27_47#_c_114_n N_A_27_47#_c_120_n N_A_27_47#_c_115_n
+ N_A_27_47#_c_122_n N_A_27_47#_c_116_n N_A_27_47#_c_124_n
+ PM_SKY130_FD_SC_LP__EBUFN_LP2%A_27_47#
x_PM_SKY130_FD_SC_LP__EBUFN_LP2%A_232_231# N_A_232_231#_M1002_d
+ N_A_232_231#_M1005_d N_A_232_231#_c_177_n N_A_232_231#_c_178_n
+ N_A_232_231#_c_179_n N_A_232_231#_M1008_g N_A_232_231#_c_181_n
+ N_A_232_231#_c_182_n N_A_232_231#_c_183_n N_A_232_231#_c_184_n
+ N_A_232_231#_c_185_n N_A_232_231#_c_186_n N_A_232_231#_c_187_n
+ N_A_232_231#_c_191_n N_A_232_231#_c_188_n N_A_232_231#_c_189_n
+ N_A_232_231#_c_190_n PM_SKY130_FD_SC_LP__EBUFN_LP2%A_232_231#
x_PM_SKY130_FD_SC_LP__EBUFN_LP2%TE_B N_TE_B_M1009_g N_TE_B_M1006_g
+ N_TE_B_M1005_g N_TE_B_M1002_g TE_B TE_B N_TE_B_c_267_n
+ PM_SKY130_FD_SC_LP__EBUFN_LP2%TE_B
x_PM_SKY130_FD_SC_LP__EBUFN_LP2%VPWR N_VPWR_M1000_d N_VPWR_M1009_d
+ N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_315_n VPWR
+ N_VPWR_c_316_n N_VPWR_c_311_n N_VPWR_c_318_n
+ PM_SKY130_FD_SC_LP__EBUFN_LP2%VPWR
x_PM_SKY130_FD_SC_LP__EBUFN_LP2%Z N_Z_M1003_s N_Z_M1004_s N_Z_c_349_n
+ N_Z_c_350_n Z Z Z Z PM_SKY130_FD_SC_LP__EBUFN_LP2%Z
x_PM_SKY130_FD_SC_LP__EBUFN_LP2%VGND N_VGND_M1007_d N_VGND_M1008_d
+ N_VGND_c_384_n N_VGND_c_385_n VGND N_VGND_c_386_n N_VGND_c_387_n
+ N_VGND_c_388_n N_VGND_c_389_n N_VGND_c_390_n N_VGND_c_391_n
+ PM_SKY130_FD_SC_LP__EBUFN_LP2%VGND
cc_1 VNB N_A_c_69_n 0.0372293f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.765
cc_2 VNB N_A_M1000_g 0.0204461f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_3 VNB N_A_c_71_n 0.0225665f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.915
cc_4 VNB N_A_c_72_n 0.0266906f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.435
cc_5 VNB A 0.002175f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_6 VNB N_A_c_74_n 0.0288115f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.93
cc_7 VNB N_A_27_47#_c_109_n 0.0367663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_110_n 0.00383763f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.765
cc_9 VNB N_A_27_47#_M1003_g 0.034322f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=0.915
cc_10 VNB N_A_27_47#_M1004_g 0.00261335f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.435
cc_11 VNB N_A_27_47#_c_113_n 0.0178293f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_A_27_47#_c_114_n 0.065636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_115_n 0.0012601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_116_n 0.00170543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_232_231#_c_177_n 0.0372338f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.765
cc_16 VNB N_A_232_231#_c_178_n 0.0616611f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_17 VNB N_A_232_231#_c_179_n 0.0108331f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_18 VNB N_A_232_231#_M1008_g 0.0232837f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.915
cc_19 VNB N_A_232_231#_c_181_n 0.00442441f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_20 VNB N_A_232_231#_c_182_n 0.0148531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_232_231#_c_183_n 0.0046752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_232_231#_c_184_n 6.17563e-19 $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.93
cc_23 VNB N_A_232_231#_c_185_n 0.0242463f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.93
cc_24 VNB N_A_232_231#_c_186_n 0.00194737f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.555
cc_25 VNB N_A_232_231#_c_187_n 0.024248f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.295
cc_26 VNB N_A_232_231#_c_188_n 0.0108904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_232_231#_c_189_n 0.0132078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_232_231#_c_190_n 0.0431782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_TE_B_M1006_g 0.0370758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_TE_B_M1002_g 0.039531f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.435
cc_31 VNB TE_B 0.00288715f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_32 VNB N_TE_B_c_267_n 0.021429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_311_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Z_c_349_n 0.00861589f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_35 VNB N_Z_c_350_n 0.0077987f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.208
cc_36 VNB Z 4.63914e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_37 VNB N_VGND_c_384_n 0.0145775f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_38 VNB N_VGND_c_385_n 0.0291248f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.915
cc_39 VNB N_VGND_c_386_n 0.0312803f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_40 VNB N_VGND_c_387_n 0.0342231f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=0.93
cc_41 VNB N_VGND_c_388_n 0.0307244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_389_n 0.244326f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.295
cc_43 VNB N_VGND_c_390_n 0.006319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_391_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A_M1000_g 0.0513237f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_46 VPB N_A_27_47#_c_110_n 0.00842711f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.765
cc_47 VPB N_A_27_47#_M1004_g 0.0299368f $X=-0.19 $Y=1.655 $X2=0.647 $Y2=1.435
cc_48 VPB N_A_27_47#_c_114_n 9.52481e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_120_n 0.0493899f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.555
cc_50 VPB N_A_27_47#_c_115_n 0.0224227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_122_n 0.0134519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_116_n 0.054253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_124_n 0.00994965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_232_231#_c_191_n 0.0291214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_232_231#_c_188_n 0.0298287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_TE_B_M1009_g 0.023206f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_57 VPB N_TE_B_M1005_g 0.0279245f $X=-0.19 $Y=1.655 $X2=0.647 $Y2=0.915
cc_58 VPB TE_B 0.00124397f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_59 VPB N_TE_B_c_267_n 0.0318952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_312_n 0.0352231f $X=-0.19 $Y=1.655 $X2=0.647 $Y2=0.915
cc_61 VPB N_VPWR_c_313_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_62 VPB N_VPWR_c_314_n 0.0540584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_315_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_316_n 0.0191606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_311_n 0.0837498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_318_n 0.0244124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB Z 0.00533f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_68 VPB Z 0.0274181f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_69 N_A_M1000_g N_A_27_47#_c_110_n 0.0109038f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_70 N_A_c_69_n N_A_27_47#_c_114_n 0.031679f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_71 A N_A_27_47#_c_114_n 0.0654014f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_72 N_A_M1000_g N_A_27_47#_c_120_n 0.0307695f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_73 N_A_M1000_g N_A_27_47#_c_115_n 0.0224651f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_74 N_A_c_72_n N_A_27_47#_c_115_n 0.0013221f $X=0.647 $Y=1.435 $X2=0 $Y2=0
cc_75 A N_A_27_47#_c_115_n 0.0197276f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_76 N_A_M1000_g N_A_27_47#_c_122_n 0.00113712f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_77 N_A_M1000_g N_A_27_47#_c_124_n 0.00513266f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_78 N_A_c_71_n N_A_232_231#_c_177_n 0.0051608f $X=0.69 $Y=0.915 $X2=0 $Y2=0
cc_79 A N_A_232_231#_c_177_n 3.64049e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_80 N_A_c_74_n N_A_232_231#_c_177_n 0.00370417f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_81 N_A_c_69_n N_A_232_231#_c_179_n 0.0051608f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_82 A N_A_232_231#_c_179_n 9.22738e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_83 N_A_M1000_g N_A_232_231#_c_181_n 2.85135e-19 $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_84 N_A_c_71_n N_A_232_231#_c_181_n 2.07712e-19 $X=0.69 $Y=0.915 $X2=0 $Y2=0
cc_85 A N_A_232_231#_c_181_n 0.0278362f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_86 N_A_c_74_n N_A_232_231#_c_181_n 0.00346263f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_87 N_A_c_69_n N_A_232_231#_c_183_n 0.00185473f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_88 A N_A_232_231#_c_183_n 0.0097312f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_89 N_A_M1000_g N_A_232_231#_c_190_n 0.00140588f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_90 A N_A_232_231#_c_190_n 0.00115096f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_91 N_A_c_74_n N_A_232_231#_c_190_n 0.0122451f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_92 N_A_M1000_g N_VPWR_c_312_n 0.0248686f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_93 N_A_M1000_g N_VPWR_c_311_n 0.014085f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_94 N_A_M1000_g N_VPWR_c_318_n 0.00769046f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_95 A A_114_47# 0.00175001f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_96 N_A_c_69_n N_VGND_c_384_n 0.0133995f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_97 A N_VGND_c_384_n 0.00779885f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_98 N_A_c_69_n N_VGND_c_386_n 0.0105812f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_99 A N_VGND_c_386_n 0.00856003f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_100 N_A_c_69_n N_VGND_c_389_n 0.0209864f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_101 A N_VGND_c_389_n 0.0109977f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_102 N_A_27_47#_M1003_g N_A_232_231#_c_177_n 0.0129854f $X=2.05 $Y=1.175 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_M1003_g N_A_232_231#_c_178_n 0.00746837f $X=2.05 $Y=1.175
+ $X2=0 $Y2=0
cc_104 N_A_27_47#_M1003_g N_A_232_231#_M1008_g 0.0140978f $X=2.05 $Y=1.175 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_110_n N_A_232_231#_c_181_n 3.72414e-19 $X=1.49 $Y=1.8 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_M1003_g N_A_232_231#_c_181_n 9.4378e-19 $X=2.05 $Y=1.175 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_115_n N_A_232_231#_c_181_n 0.0269982f $X=1.16 $Y=1.76 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_M1003_g N_A_232_231#_c_182_n 0.0090251f $X=2.05 $Y=1.175 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_M1003_g N_A_232_231#_c_184_n 0.00306209f $X=2.05 $Y=1.175
+ $X2=0 $Y2=0
cc_110 N_A_27_47#_c_113_n N_A_232_231#_c_185_n 8.88e-19 $X=2.175 $Y=1.8 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_M1003_g N_A_232_231#_c_186_n 0.00255619f $X=2.05 $Y=1.175
+ $X2=0 $Y2=0
cc_112 N_A_27_47#_c_113_n N_A_232_231#_c_186_n 0.00370096f $X=2.175 $Y=1.8 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_110_n N_A_232_231#_c_190_n 0.0255328f $X=1.49 $Y=1.8 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_115_n N_A_232_231#_c_190_n 0.0013126f $X=1.16 $Y=1.76 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_M1004_g N_TE_B_M1009_g 0.0407661f $X=2.25 $Y=2.595 $X2=0 $Y2=0
cc_116 N_A_27_47#_M1003_g TE_B 4.23194e-19 $X=2.05 $Y=1.175 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_113_n TE_B 0.00350593f $X=2.175 $Y=1.8 $X2=0 $Y2=0
cc_118 N_A_27_47#_M1003_g N_TE_B_c_267_n 0.00241356f $X=2.05 $Y=1.175 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_c_113_n N_TE_B_c_267_n 0.0407661f $X=2.175 $Y=1.8 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_120_n N_VPWR_c_312_n 0.0685263f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_115_n N_VPWR_c_312_n 0.0264018f $X=1.16 $Y=1.76 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_122_n N_VPWR_c_312_n 0.0274812f $X=1.325 $Y=1.89 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_116_n N_VPWR_c_312_n 0.0033192f $X=1.325 $Y=1.89 $X2=0 $Y2=0
cc_124 N_A_27_47#_M1004_g N_VPWR_c_313_n 0.00295152f $X=2.25 $Y=2.595 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_M1004_g N_VPWR_c_314_n 0.00751517f $X=2.25 $Y=2.595 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_M1004_g N_VPWR_c_311_n 0.0128147f $X=2.25 $Y=2.595 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_120_n N_VPWR_c_311_n 0.0125808f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_120_n N_VPWR_c_318_n 0.0220321f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_109_n N_Z_c_349_n 0.00184202f $X=1.975 $Y=1.8 $X2=0 $Y2=0
cc_130 N_A_27_47#_M1003_g N_Z_c_349_n 0.0156564f $X=2.05 $Y=1.175 $X2=0 $Y2=0
cc_131 N_A_27_47#_c_109_n N_Z_c_350_n 0.0145999f $X=1.975 $Y=1.8 $X2=0 $Y2=0
cc_132 N_A_27_47#_M1003_g N_Z_c_350_n 0.0110453f $X=2.05 $Y=1.175 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_113_n N_Z_c_350_n 0.00588611f $X=2.175 $Y=1.8 $X2=0 $Y2=0
cc_134 N_A_27_47#_c_115_n N_Z_c_350_n 0.00838339f $X=1.16 $Y=1.76 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_109_n Z 0.00494178f $X=1.975 $Y=1.8 $X2=0 $Y2=0
cc_136 N_A_27_47#_M1004_g Z 0.0133591f $X=2.25 $Y=2.595 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_113_n Z 0.00641913f $X=2.175 $Y=1.8 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_115_n Z 0.0020536f $X=1.16 $Y=1.76 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_122_n Z 0.02295f $X=1.325 $Y=1.89 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_116_n Z 0.00459135f $X=1.325 $Y=1.89 $X2=0 $Y2=0
cc_141 N_A_27_47#_M1004_g Z 0.0288445f $X=2.25 $Y=2.595 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_114_n N_VGND_c_386_n 0.0163773f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A_27_47#_M1001_s N_VGND_c_389_n 0.00427743f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_c_114_n N_VGND_c_389_n 0.00959046f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_145 N_A_232_231#_c_191_n N_TE_B_M1009_g 2.09334e-19 $X=3.535 $Y=2.495 $X2=0
+ $Y2=0
cc_146 N_A_232_231#_M1008_g N_TE_B_M1006_g 0.0155717f $X=2.525 $Y=0.975 $X2=0
+ $Y2=0
cc_147 N_A_232_231#_c_185_n N_TE_B_M1006_g 0.0151834f $X=3.395 $Y=1.34 $X2=0
+ $Y2=0
cc_148 N_A_232_231#_c_187_n N_TE_B_M1006_g 0.00182338f $X=3.56 $Y=0.975 $X2=0
+ $Y2=0
cc_149 N_A_232_231#_c_191_n N_TE_B_M1005_g 0.0140367f $X=3.535 $Y=2.495 $X2=0
+ $Y2=0
cc_150 N_A_232_231#_c_185_n N_TE_B_M1002_g 0.0144737f $X=3.395 $Y=1.34 $X2=0
+ $Y2=0
cc_151 N_A_232_231#_c_187_n N_TE_B_M1002_g 0.0115067f $X=3.56 $Y=0.975 $X2=0
+ $Y2=0
cc_152 N_A_232_231#_c_188_n N_TE_B_M1002_g 0.00900567f $X=3.547 $Y=2.33 $X2=0
+ $Y2=0
cc_153 N_A_232_231#_c_189_n N_TE_B_M1002_g 0.00496925f $X=3.56 $Y=1.34 $X2=0
+ $Y2=0
cc_154 N_A_232_231#_M1008_g TE_B 4.3524e-19 $X=2.525 $Y=0.975 $X2=0 $Y2=0
cc_155 N_A_232_231#_c_185_n TE_B 0.0529774f $X=3.395 $Y=1.34 $X2=0 $Y2=0
cc_156 N_A_232_231#_c_188_n TE_B 0.0269335f $X=3.547 $Y=2.33 $X2=0 $Y2=0
cc_157 N_A_232_231#_c_185_n N_TE_B_c_267_n 0.00850661f $X=3.395 $Y=1.34 $X2=0
+ $Y2=0
cc_158 N_A_232_231#_c_188_n N_TE_B_c_267_n 0.0148496f $X=3.547 $Y=2.33 $X2=0
+ $Y2=0
cc_159 N_A_232_231#_c_191_n N_VPWR_c_313_n 0.0486685f $X=3.535 $Y=2.495 $X2=0
+ $Y2=0
cc_160 N_A_232_231#_c_191_n N_VPWR_c_316_n 0.0214436f $X=3.535 $Y=2.495 $X2=0
+ $Y2=0
cc_161 N_A_232_231#_M1005_d N_VPWR_c_311_n 0.0023218f $X=3.395 $Y=2.095 $X2=0
+ $Y2=0
cc_162 N_A_232_231#_c_191_n N_VPWR_c_311_n 0.0134754f $X=3.535 $Y=2.495 $X2=0
+ $Y2=0
cc_163 N_A_232_231#_c_177_n N_Z_c_349_n 0.00395179f $X=1.515 $Y=1.155 $X2=0
+ $Y2=0
cc_164 N_A_232_231#_c_181_n N_Z_c_349_n 0.0310432f $X=1.325 $Y=1.32 $X2=0 $Y2=0
cc_165 N_A_232_231#_c_182_n N_Z_c_349_n 0.022977f $X=2.18 $Y=0.81 $X2=0 $Y2=0
cc_166 N_A_232_231#_c_186_n N_Z_c_349_n 0.00786608f $X=2.35 $Y=1.34 $X2=0 $Y2=0
cc_167 N_A_232_231#_c_186_n N_Z_c_350_n 0.00772283f $X=2.35 $Y=1.34 $X2=0 $Y2=0
cc_168 N_A_232_231#_c_179_n N_VGND_c_384_n 0.00323886f $X=1.59 $Y=0.52 $X2=0
+ $Y2=0
cc_169 N_A_232_231#_c_183_n N_VGND_c_384_n 0.0188101f $X=1.49 $Y=0.81 $X2=0
+ $Y2=0
cc_170 N_A_232_231#_c_190_n N_VGND_c_384_n 7.365e-19 $X=1.515 $Y=1.32 $X2=0
+ $Y2=0
cc_171 N_A_232_231#_c_178_n N_VGND_c_385_n 0.0110769f $X=2.45 $Y=0.52 $X2=0
+ $Y2=0
cc_172 N_A_232_231#_M1008_g N_VGND_c_385_n 0.0123096f $X=2.525 $Y=0.975 $X2=0
+ $Y2=0
cc_173 N_A_232_231#_c_182_n N_VGND_c_385_n 0.0113843f $X=2.18 $Y=0.81 $X2=0
+ $Y2=0
cc_174 N_A_232_231#_c_184_n N_VGND_c_385_n 0.0106821f $X=2.265 $Y=1.255 $X2=0
+ $Y2=0
cc_175 N_A_232_231#_c_185_n N_VGND_c_385_n 0.0207154f $X=3.395 $Y=1.34 $X2=0
+ $Y2=0
cc_176 N_A_232_231#_c_187_n N_VGND_c_385_n 0.0104546f $X=3.56 $Y=0.975 $X2=0
+ $Y2=0
cc_177 N_A_232_231#_c_179_n N_VGND_c_387_n 0.0236022f $X=1.59 $Y=0.52 $X2=0
+ $Y2=0
cc_178 N_A_232_231#_c_182_n N_VGND_c_387_n 0.0130994f $X=2.18 $Y=0.81 $X2=0
+ $Y2=0
cc_179 N_A_232_231#_c_183_n N_VGND_c_387_n 0.00166219f $X=1.49 $Y=0.81 $X2=0
+ $Y2=0
cc_180 N_A_232_231#_c_187_n N_VGND_c_388_n 0.00531453f $X=3.56 $Y=0.975 $X2=0
+ $Y2=0
cc_181 N_A_232_231#_c_179_n N_VGND_c_389_n 0.0321234f $X=1.59 $Y=0.52 $X2=0
+ $Y2=0
cc_182 N_A_232_231#_c_182_n N_VGND_c_389_n 0.0230971f $X=2.18 $Y=0.81 $X2=0
+ $Y2=0
cc_183 N_A_232_231#_c_183_n N_VGND_c_389_n 0.00396299f $X=1.49 $Y=0.81 $X2=0
+ $Y2=0
cc_184 N_A_232_231#_c_187_n N_VGND_c_389_n 0.00914353f $X=3.56 $Y=0.975 $X2=0
+ $Y2=0
cc_185 N_A_232_231#_c_182_n A_425_193# 0.00156358f $X=2.18 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_186 N_A_232_231#_c_184_n A_425_193# 0.00495387f $X=2.265 $Y=1.255 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_232_231#_c_185_n A_425_193# 7.30555e-19 $X=3.395 $Y=1.34 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_232_231#_c_186_n A_425_193# 6.33207e-19 $X=2.35 $Y=1.34 $X2=-0.19
+ $Y2=-0.245
cc_189 TE_B N_VPWR_M1009_d 0.00187356f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_190 N_TE_B_M1009_g N_VPWR_c_313_n 0.0215909f $X=2.74 $Y=2.595 $X2=0 $Y2=0
cc_191 N_TE_B_M1005_g N_VPWR_c_313_n 0.0200812f $X=3.27 $Y=2.595 $X2=0 $Y2=0
cc_192 TE_B N_VPWR_c_313_n 0.0177591f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_193 N_TE_B_c_267_n N_VPWR_c_313_n 4.82215e-19 $X=3.27 $Y=1.77 $X2=0 $Y2=0
cc_194 N_TE_B_M1009_g N_VPWR_c_314_n 0.008763f $X=2.74 $Y=2.595 $X2=0 $Y2=0
cc_195 N_TE_B_M1005_g N_VPWR_c_316_n 0.00840199f $X=3.27 $Y=2.595 $X2=0 $Y2=0
cc_196 N_TE_B_M1009_g N_VPWR_c_311_n 0.0144563f $X=2.74 $Y=2.595 $X2=0 $Y2=0
cc_197 N_TE_B_M1005_g N_VPWR_c_311_n 0.0145458f $X=3.27 $Y=2.595 $X2=0 $Y2=0
cc_198 TE_B N_Z_c_350_n 0.011702f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_199 N_TE_B_c_267_n N_Z_c_350_n 5.06318e-19 $X=3.27 $Y=1.77 $X2=0 $Y2=0
cc_200 N_TE_B_M1009_g Z 0.003618f $X=2.74 $Y=2.595 $X2=0 $Y2=0
cc_201 TE_B Z 0.0232372f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_202 TE_B A_475_419# 0.00199544f $X=3.035 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_203 N_TE_B_M1006_g N_VGND_c_385_n 0.00988212f $X=2.955 $Y=0.975 $X2=0 $Y2=0
cc_204 N_TE_B_M1002_g N_VGND_c_385_n 0.00147934f $X=3.345 $Y=0.975 $X2=0 $Y2=0
cc_205 N_TE_B_M1006_g N_VGND_c_388_n 0.00289826f $X=2.955 $Y=0.975 $X2=0 $Y2=0
cc_206 N_TE_B_M1002_g N_VGND_c_388_n 0.00337154f $X=3.345 $Y=0.975 $X2=0 $Y2=0
cc_207 N_TE_B_M1006_g N_VGND_c_389_n 0.00363223f $X=2.955 $Y=0.975 $X2=0 $Y2=0
cc_208 N_TE_B_M1002_g N_VGND_c_389_n 0.00432409f $X=3.345 $Y=0.975 $X2=0 $Y2=0
cc_209 N_VPWR_c_311_n N_Z_M1004_s 0.0023218f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_210 N_VPWR_c_313_n Z 0.021035f $X=3.005 $Y=2.495 $X2=0 $Y2=0
cc_211 N_VPWR_c_314_n Z 0.0277532f $X=2.84 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_311_n Z 0.0167689f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_311_n A_475_419# 0.010279f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_214 A_114_47# N_VGND_c_389_n 0.00219029f $X=0.57 $Y=0.235 $X2=0.71 $Y2=1.295
