* File: sky130_fd_sc_lp__a41oi_4.pxi.spice
* Created: Fri Aug 28 10:03:38 2020
* 
x_PM_SKY130_FD_SC_LP__A41OI_4%B1 N_B1_c_156_n N_B1_M1014_g N_B1_M1007_g
+ N_B1_c_158_n N_B1_M1021_g N_B1_M1013_g N_B1_c_160_n N_B1_M1022_g N_B1_M1023_g
+ N_B1_c_162_n N_B1_M1039_g N_B1_c_168_n N_B1_M1027_g B1 B1 B1 B1 N_B1_c_164_n
+ PM_SKY130_FD_SC_LP__A41OI_4%B1
x_PM_SKY130_FD_SC_LP__A41OI_4%A1 N_A1_M1002_g N_A1_M1010_g N_A1_M1004_g
+ N_A1_M1026_g N_A1_M1018_g N_A1_M1034_g N_A1_M1036_g N_A1_M1037_g N_A1_c_243_n
+ N_A1_c_244_n N_A1_c_245_n A1 A1 N_A1_c_246_n N_A1_c_247_n N_A1_c_248_n
+ PM_SKY130_FD_SC_LP__A41OI_4%A1
x_PM_SKY130_FD_SC_LP__A41OI_4%A2 N_A2_M1001_g N_A2_c_325_n N_A2_M1008_g
+ N_A2_M1012_g N_A2_c_327_n N_A2_M1020_g N_A2_M1017_g N_A2_c_329_n N_A2_M1028_g
+ N_A2_c_330_n N_A2_M1038_g N_A2_M1031_g A2 A2 N_A2_c_332_n N_A2_c_333_n
+ PM_SKY130_FD_SC_LP__A41OI_4%A2
x_PM_SKY130_FD_SC_LP__A41OI_4%A3 N_A3_M1003_g N_A3_M1019_g N_A3_c_422_n
+ N_A3_M1006_g N_A3_M1032_g N_A3_c_424_n N_A3_M1009_g N_A3_c_425_n N_A3_M1030_g
+ N_A3_M1033_g N_A3_c_427_n N_A3_M1035_g N_A3_c_428_n A3 N_A3_c_430_n
+ N_A3_c_431_n PM_SKY130_FD_SC_LP__A41OI_4%A3
x_PM_SKY130_FD_SC_LP__A41OI_4%A4 N_A4_M1000_g N_A4_c_512_n N_A4_M1005_g
+ N_A4_M1011_g N_A4_c_514_n N_A4_M1016_g N_A4_M1015_g N_A4_c_516_n N_A4_M1025_g
+ N_A4_M1024_g N_A4_c_518_n N_A4_M1029_g A4 A4 A4 A4 N_A4_c_520_n N_A4_c_521_n
+ PM_SKY130_FD_SC_LP__A41OI_4%A4
x_PM_SKY130_FD_SC_LP__A41OI_4%A_30_367# N_A_30_367#_M1007_d N_A_30_367#_M1013_d
+ N_A_30_367#_M1027_d N_A_30_367#_M1010_s N_A_30_367#_M1036_s
+ N_A_30_367#_M1012_d N_A_30_367#_M1031_d N_A_30_367#_M1019_d
+ N_A_30_367#_M1033_d N_A_30_367#_M1011_d N_A_30_367#_M1024_d
+ N_A_30_367#_c_587_n N_A_30_367#_c_588_n N_A_30_367#_c_603_n
+ N_A_30_367#_c_676_p N_A_30_367#_c_605_n N_A_30_367#_c_668_p
+ N_A_30_367#_c_607_n N_A_30_367#_c_609_n N_A_30_367#_c_611_n
+ N_A_30_367#_c_615_n N_A_30_367#_c_619_n N_A_30_367#_c_701_p
+ N_A_30_367#_c_589_n N_A_30_367#_c_590_n N_A_30_367#_c_628_n
+ N_A_30_367#_c_591_n N_A_30_367#_c_703_p N_A_30_367#_c_592_n
+ N_A_30_367#_c_698_p N_A_30_367#_c_593_n N_A_30_367#_c_699_p
+ N_A_30_367#_c_594_n N_A_30_367#_c_595_n N_A_30_367#_c_697_p
+ N_A_30_367#_c_674_p N_A_30_367#_c_612_n N_A_30_367#_c_631_n
+ N_A_30_367#_c_596_n N_A_30_367#_c_597_n N_A_30_367#_c_598_n
+ N_A_30_367#_c_599_n PM_SKY130_FD_SC_LP__A41OI_4%A_30_367#
x_PM_SKY130_FD_SC_LP__A41OI_4%Y N_Y_M1014_d N_Y_M1022_d N_Y_M1004_s N_Y_M1034_s
+ N_Y_M1007_s N_Y_M1023_s N_Y_c_738_n N_Y_c_832_p N_Y_c_741_n N_Y_c_745_n
+ N_Y_c_728_n N_Y_c_751_n N_Y_c_831_p N_Y_c_735_n N_Y_c_729_n N_Y_c_730_n
+ N_Y_c_731_n N_Y_c_732_n Y Y Y Y Y N_Y_c_733_n Y Y N_Y_c_734_n
+ PM_SKY130_FD_SC_LP__A41OI_4%Y
x_PM_SKY130_FD_SC_LP__A41OI_4%VPWR N_VPWR_M1002_d N_VPWR_M1026_d N_VPWR_M1001_s
+ N_VPWR_M1017_s N_VPWR_M1003_s N_VPWR_M1032_s N_VPWR_M1000_s N_VPWR_M1015_s
+ N_VPWR_c_850_n N_VPWR_c_851_n N_VPWR_c_852_n N_VPWR_c_853_n N_VPWR_c_854_n
+ N_VPWR_c_855_n N_VPWR_c_856_n N_VPWR_c_857_n N_VPWR_c_858_n N_VPWR_c_859_n
+ N_VPWR_c_860_n N_VPWR_c_861_n N_VPWR_c_862_n N_VPWR_c_863_n N_VPWR_c_864_n
+ VPWR N_VPWR_c_865_n N_VPWR_c_866_n N_VPWR_c_867_n N_VPWR_c_868_n
+ N_VPWR_c_869_n N_VPWR_c_849_n N_VPWR_c_871_n N_VPWR_c_872_n N_VPWR_c_873_n
+ N_VPWR_c_874_n N_VPWR_c_875_n PM_SKY130_FD_SC_LP__A41OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A41OI_4%VGND N_VGND_M1014_s N_VGND_M1021_s N_VGND_M1039_s
+ N_VGND_M1005_d N_VGND_M1025_d N_VGND_c_997_n N_VGND_c_998_n N_VGND_c_999_n
+ N_VGND_c_1000_n N_VGND_c_1001_n N_VGND_c_1002_n N_VGND_c_1003_n
+ N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n N_VGND_c_1007_n
+ N_VGND_c_1008_n VGND N_VGND_c_1009_n N_VGND_c_1010_n N_VGND_c_1011_n
+ N_VGND_c_1012_n PM_SKY130_FD_SC_LP__A41OI_4%VGND
x_PM_SKY130_FD_SC_LP__A41OI_4%A_478_65# N_A_478_65#_M1004_d N_A_478_65#_M1018_d
+ N_A_478_65#_M1037_d N_A_478_65#_M1020_s N_A_478_65#_M1038_s
+ N_A_478_65#_c_1114_n N_A_478_65#_c_1115_n N_A_478_65#_c_1126_n
+ N_A_478_65#_c_1116_n N_A_478_65#_c_1117_n N_A_478_65#_c_1118_n
+ N_A_478_65#_c_1119_n N_A_478_65#_c_1120_n
+ PM_SKY130_FD_SC_LP__A41OI_4%A_478_65#
x_PM_SKY130_FD_SC_LP__A41OI_4%A_921_65# N_A_921_65#_M1008_d N_A_921_65#_M1028_d
+ N_A_921_65#_M1006_s N_A_921_65#_M1030_s N_A_921_65#_c_1160_n
+ N_A_921_65#_c_1173_n N_A_921_65#_c_1166_n N_A_921_65#_c_1179_n
+ N_A_921_65#_c_1184_n PM_SKY130_FD_SC_LP__A41OI_4%A_921_65#
x_PM_SKY130_FD_SC_LP__A41OI_4%A_1291_65# N_A_1291_65#_M1006_d
+ N_A_1291_65#_M1009_d N_A_1291_65#_M1035_d N_A_1291_65#_M1016_s
+ N_A_1291_65#_M1029_s N_A_1291_65#_c_1210_n N_A_1291_65#_c_1211_n
+ N_A_1291_65#_c_1225_n N_A_1291_65#_c_1212_n N_A_1291_65#_c_1213_n
+ N_A_1291_65#_c_1214_n N_A_1291_65#_c_1215_n N_A_1291_65#_c_1216_n
+ N_A_1291_65#_c_1235_n PM_SKY130_FD_SC_LP__A41OI_4%A_1291_65#
cc_1 VNB N_B1_c_156_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_B1_M1007_g 0.0109769f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_3 VNB N_B1_c_158_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.185
cc_4 VNB N_B1_M1013_g 0.00665511f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_5 VNB N_B1_c_160_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.185
cc_6 VNB N_B1_M1023_g 0.00648053f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_7 VNB N_B1_c_162_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.185
cc_8 VNB B1 0.0111559f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_9 VNB N_B1_c_164_n 0.118672f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.455
cc_10 VNB N_A1_M1004_g 0.0231113f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_11 VNB N_A1_M1018_g 0.0182986f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_12 VNB N_A1_M1034_g 0.0184379f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_13 VNB N_A1_M1037_g 0.0188722f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_14 VNB N_A1_c_243_n 0.00201995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_244_n 0.00554835f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.455
cc_16 VNB N_A1_c_245_n 0.00105136f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.455
cc_17 VNB N_A1_c_246_n 0.00187739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_247_n 0.104543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_248_n 5.77127e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_M1001_g 0.00213574f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_21 VNB N_A2_c_325_n 0.0166882f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_22 VNB N_A2_M1012_g 0.00248458f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_23 VNB N_A2_c_327_n 0.0155792f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_24 VNB N_A2_M1017_g 0.00278413f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_25 VNB N_A2_c_329_n 0.0155811f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_26 VNB N_A2_c_330_n 0.0200848f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.185
cc_27 VNB N_A2_M1031_g 0.00286745f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_28 VNB N_A2_c_332_n 0.0150764f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.455
cc_29 VNB N_A2_c_333_n 0.0945457f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.35
cc_30 VNB N_A3_M1003_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_31 VNB N_A3_M1019_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A3_c_422_n 0.0218447f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_33 VNB N_A3_M1032_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A3_c_424_n 0.0161985f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_35 VNB N_A3_c_425_n 0.0161979f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_36 VNB N_A3_M1033_g 0.00402655f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_37 VNB N_A3_c_427_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_38 VNB N_A3_c_428_n 0.00152296f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.455
cc_39 VNB A3 0.00200247f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.455
cc_40 VNB N_A3_c_430_n 0.00179014f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.322
cc_41 VNB N_A3_c_431_n 0.126438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A4_M1000_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_43 VNB N_A4_c_512_n 0.015918f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_44 VNB N_A4_M1011_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_45 VNB N_A4_c_514_n 0.0157113f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_46 VNB N_A4_M1015_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_47 VNB N_A4_c_516_n 0.0157113f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_48 VNB N_A4_M1024_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_49 VNB N_A4_c_518_n 0.0210357f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_50 VNB A4 0.0400296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A4_c_520_n 0.0711038f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.35
cc_52 VNB N_A4_c_521_n 0.0679427f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.455
cc_53 VNB N_Y_c_728_n 0.00228659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_Y_c_729_n 0.00215668f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.455
cc_55 VNB N_Y_c_730_n 0.00367643f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.455
cc_56 VNB N_Y_c_731_n 0.00224024f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.322
cc_57 VNB N_Y_c_732_n 0.0020857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Y_c_733_n 0.0090193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_Y_c_734_n 0.00228422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VPWR_c_849_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_997_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_62 VNB N_VGND_c_998_n 0.03399f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.515
cc_63 VNB N_VGND_c_999_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.185
cc_64 VNB N_VGND_c_1000_n 0.00693495f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_65 VNB N_VGND_c_1001_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_66 VNB N_VGND_c_1002_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1003_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.35
cc_68 VNB N_VGND_c_1004_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.35
cc_69 VNB N_VGND_c_1005_n 0.148537f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.455
cc_70 VNB N_VGND_c_1006_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.455
cc_71 VNB N_VGND_c_1007_n 0.0143206f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.455
cc_72 VNB N_VGND_c_1008_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.455
cc_73 VNB N_VGND_c_1009_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.35
cc_74 VNB N_VGND_c_1010_n 0.0251472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1011_n 0.539625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1012_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_478_65#_c_1114_n 0.00864516f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.655
cc_78 VNB N_A_478_65#_c_1115_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_79 VNB N_A_478_65#_c_1116_n 0.0017696f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_80 VNB N_A_478_65#_c_1117_n 0.00462783f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_81 VNB N_A_478_65#_c_1118_n 0.00140846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_478_65#_c_1119_n 0.00221073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_478_65#_c_1120_n 0.00223571f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.35
cc_84 VNB N_A_921_65#_c_1160_n 0.0102812f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_85 VNB N_A_1291_65#_c_1210_n 0.00296443f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.655
cc_86 VNB N_A_1291_65#_c_1211_n 0.00467132f $X=-0.19 $Y=-0.245 $X2=1.35
+ $Y2=1.515
cc_87 VNB N_A_1291_65#_c_1212_n 0.00168804f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_88 VNB N_A_1291_65#_c_1213_n 0.00742396f $X=-0.19 $Y=-0.245 $X2=1.115
+ $Y2=1.21
cc_89 VNB N_A_1291_65#_c_1214_n 0.0226918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1291_65#_c_1215_n 0.00237493f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.455
cc_91 VNB N_A_1291_65#_c_1216_n 0.0016096f $X=-0.19 $Y=-0.245 $X2=0.905
+ $Y2=1.455
cc_92 VPB N_B1_M1007_g 0.0267546f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_93 VPB N_B1_M1013_g 0.0184533f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_94 VPB N_B1_M1023_g 0.0183748f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_95 VPB N_B1_c_168_n 0.0154285f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=1.725
cc_96 VPB N_B1_c_164_n 0.00438061f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.455
cc_97 VPB N_A1_M1002_g 0.0192091f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_98 VPB N_A1_M1010_g 0.0190302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A1_M1026_g 0.0223035f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.185
cc_100 VPB N_A1_M1036_g 0.0228609f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_101 VPB N_A1_c_247_n 0.0217689f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A2_M1001_g 0.0186975f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_103 VPB N_A2_M1012_g 0.0194385f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.655
cc_104 VPB N_A2_M1017_g 0.0208791f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.655
cc_105 VPB N_A2_M1031_g 0.0211037f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_106 VPB N_A3_M1003_g 0.0191445f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_107 VPB N_A3_M1019_g 0.018914f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A3_M1032_g 0.0250833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A3_M1033_g 0.0253137f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.655
cc_110 VPB N_A4_M1000_g 0.0191445f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_111 VPB N_A4_M1011_g 0.018914f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.655
cc_112 VPB N_A4_M1015_g 0.018914f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.655
cc_113 VPB N_A4_M1024_g 0.0257505f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.655
cc_114 VPB N_A_30_367#_c_587_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_30_367#_c_588_n 0.043141f $X=-0.19 $Y=1.655 $X2=0.3 $Y2=1.455
cc_116 VPB N_A_30_367#_c_589_n 0.00372464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_30_367#_c_590_n 0.00197016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_30_367#_c_591_n 0.00416497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_30_367#_c_592_n 0.00714183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_30_367#_c_593_n 0.00416497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_30_367#_c_594_n 0.0118833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_30_367#_c_595_n 0.0435297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_30_367#_c_596_n 0.00714615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_30_367#_c_597_n 0.00145388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_30_367#_c_598_n 0.00687222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_30_367#_c_599_n 0.00145388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_Y_c_735_n 0.0215161f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.455
cc_128 VPB N_Y_c_730_n 9.13216e-19 $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.455
cc_129 VPB N_Y_c_731_n 0.00491982f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.322
cc_130 VPB N_VPWR_c_850_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_131 VPB N_VPWR_c_851_n 0.00415689f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_132 VPB N_VPWR_c_852_n 0.017949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_853_n 0.00388531f $X=-0.19 $Y=1.655 $X2=0.3 $Y2=1.35
cc_134 VPB N_VPWR_c_854_n 0.00446937f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.455
cc_135 VPB N_VPWR_c_855_n 3.22457e-19 $X=-0.19 $Y=1.655 $X2=1.66 $Y2=1.35
cc_136 VPB N_VPWR_c_856_n 0.00273395f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.322
cc_137 VPB N_VPWR_c_857_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_858_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_859_n 0.0543279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_860_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_861_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_862_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_863_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_864_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_865_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_866_n 0.0183816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_867_n 0.0157463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_868_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_869_n 0.0247634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_849_n 0.0585491f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_871_n 0.0117633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_872_n 0.00420242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_873_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_874_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_875_n 0.0138973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 N_B1_c_164_n N_A1_M1002_g 0.0342449f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_157 B1 N_A1_c_246_n 0.00179429f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_158 N_B1_c_164_n N_A1_c_246_n 0.00102232f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_159 B1 N_A1_c_247_n 6.41564e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_160 N_B1_c_164_n N_A1_c_247_n 0.0196692f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_161 N_B1_M1007_g N_A_30_367#_c_588_n 0.00293325f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_162 B1 N_A_30_367#_c_588_n 0.0115406f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_163 N_B1_c_164_n N_A_30_367#_c_588_n 0.00523662f $X=1.765 $Y=1.455 $X2=0
+ $Y2=0
cc_164 N_B1_M1007_g N_A_30_367#_c_603_n 0.0115031f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_165 N_B1_M1013_g N_A_30_367#_c_603_n 0.0115031f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_166 N_B1_M1023_g N_A_30_367#_c_605_n 0.0114565f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_167 N_B1_c_168_n N_A_30_367#_c_605_n 0.0114502f $X=1.78 $Y=1.725 $X2=0 $Y2=0
cc_168 N_B1_M1007_g N_Y_c_738_n 0.0120135f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_169 N_B1_M1013_g N_Y_c_738_n 0.0116083f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_170 N_B1_M1023_g N_Y_c_738_n 6.55859e-19 $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_171 N_B1_c_158_n N_Y_c_741_n 0.0102032f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_172 N_B1_c_160_n N_Y_c_741_n 0.0101525f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_173 B1 N_Y_c_741_n 0.0400433f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_174 N_B1_c_164_n N_Y_c_741_n 0.0023741f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_175 B1 N_Y_c_745_n 0.0142048f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_176 N_B1_c_164_n N_Y_c_745_n 0.0024616f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_177 N_B1_M1007_g N_Y_c_728_n 0.0112984f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_178 N_B1_M1013_g N_Y_c_728_n 0.00300755f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_179 B1 N_Y_c_728_n 0.0268977f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_180 N_B1_c_164_n N_Y_c_728_n 0.00263213f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_181 N_B1_M1023_g N_Y_c_751_n 0.00866824f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B1_c_168_n N_Y_c_751_n 0.00985266f $X=1.78 $Y=1.725 $X2=0 $Y2=0
cc_183 N_B1_c_168_n N_Y_c_735_n 0.00562053f $X=1.78 $Y=1.725 $X2=0 $Y2=0
cc_184 B1 N_Y_c_735_n 4.1067e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_185 N_B1_M1013_g N_Y_c_731_n 0.0115646f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B1_M1023_g N_Y_c_731_n 0.0115646f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_187 B1 N_Y_c_731_n 0.0692257f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_188 N_B1_c_164_n N_Y_c_731_n 0.00253428f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_189 N_B1_M1013_g N_Y_c_732_n 4.13719e-19 $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_190 N_B1_M1023_g N_Y_c_732_n 0.00596889f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B1_c_168_n N_Y_c_732_n 0.00791428f $X=1.78 $Y=1.725 $X2=0 $Y2=0
cc_192 N_B1_c_164_n N_Y_c_732_n 0.00897097f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_193 B1 Y 0.0142048f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_194 N_B1_c_164_n Y 0.00252239f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_195 N_B1_c_162_n N_Y_c_733_n 0.0139872f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_196 B1 N_Y_c_733_n 0.0111102f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_197 N_B1_c_168_n N_VPWR_c_850_n 0.00105138f $X=1.78 $Y=1.725 $X2=0 $Y2=0
cc_198 N_B1_M1007_g N_VPWR_c_859_n 0.00357877f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_199 N_B1_M1013_g N_VPWR_c_859_n 0.00357877f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_200 N_B1_M1023_g N_VPWR_c_859_n 0.00357877f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_201 N_B1_c_168_n N_VPWR_c_859_n 0.00357877f $X=1.78 $Y=1.725 $X2=0 $Y2=0
cc_202 N_B1_M1007_g N_VPWR_c_849_n 0.00629771f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B1_M1013_g N_VPWR_c_849_n 0.0053512f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B1_M1023_g N_VPWR_c_849_n 0.0053512f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B1_c_168_n N_VPWR_c_849_n 0.00537654f $X=1.78 $Y=1.725 $X2=0 $Y2=0
cc_206 N_B1_c_156_n N_VGND_c_998_n 0.0165371f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_207 N_B1_c_158_n N_VGND_c_998_n 6.19948e-19 $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_208 B1 N_VGND_c_998_n 0.0235917f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_209 N_B1_c_164_n N_VGND_c_998_n 0.00617954f $X=1.765 $Y=1.455 $X2=0 $Y2=0
cc_210 N_B1_c_156_n N_VGND_c_999_n 5.71572e-19 $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_211 N_B1_c_158_n N_VGND_c_999_n 0.0100576f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_212 N_B1_c_160_n N_VGND_c_999_n 0.0100576f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_213 N_B1_c_162_n N_VGND_c_999_n 5.71572e-19 $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_214 N_B1_c_160_n N_VGND_c_1000_n 5.60256e-19 $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_215 N_B1_c_162_n N_VGND_c_1000_n 0.0108619f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_216 N_B1_c_160_n N_VGND_c_1003_n 0.00486043f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_217 N_B1_c_162_n N_VGND_c_1003_n 0.00486043f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_218 N_B1_c_156_n N_VGND_c_1009_n 0.00486043f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_219 N_B1_c_158_n N_VGND_c_1009_n 0.00486043f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_220 N_B1_c_156_n N_VGND_c_1011_n 0.00824727f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_221 N_B1_c_158_n N_VGND_c_1011_n 0.00457229f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_222 N_B1_c_160_n N_VGND_c_1011_n 0.00457229f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_223 N_B1_c_162_n N_VGND_c_1011_n 0.00448921f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_224 N_B1_c_162_n N_A_478_65#_c_1114_n 8.76807e-19 $X=1.765 $Y=1.185 $X2=0
+ $Y2=0
cc_225 N_A1_M1036_g N_A2_M1001_g 0.0233611f $X=3.95 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A1_c_247_n N_A2_M1001_g 0.0123265f $X=4.02 $Y=1.49 $X2=0 $Y2=0
cc_227 N_A1_M1037_g N_A2_c_325_n 0.0220367f $X=4.02 $Y=0.745 $X2=0 $Y2=0
cc_228 N_A1_M1037_g N_A2_c_333_n 0.0123265f $X=4.02 $Y=0.745 $X2=0 $Y2=0
cc_229 N_A1_M1002_g N_A_30_367#_c_607_n 0.0132511f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A1_M1010_g N_A_30_367#_c_607_n 0.0126349f $X=2.66 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A1_M1026_g N_A_30_367#_c_609_n 0.0147891f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A1_M1036_g N_A_30_367#_c_609_n 0.0130921f $X=3.95 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A1_M1036_g N_A_30_367#_c_611_n 0.014453f $X=3.95 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A1_M1036_g N_A_30_367#_c_612_n 7.54694e-19 $X=3.95 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A1_M1002_g N_Y_c_751_n 7.64429e-19 $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A1_M1002_g N_Y_c_735_n 0.0113f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A1_M1010_g N_Y_c_735_n 0.0114071f $X=2.66 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A1_M1026_g N_Y_c_735_n 0.0129765f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A1_M1036_g N_Y_c_735_n 0.0129646f $X=3.95 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A1_c_246_n N_Y_c_735_n 0.146815f $X=2.57 $Y=1.49 $X2=0 $Y2=0
cc_241 N_A1_c_247_n N_Y_c_735_n 0.0243167f $X=4.02 $Y=1.49 $X2=0 $Y2=0
cc_242 N_A1_M1037_g N_Y_c_729_n 0.0105652f $X=4.02 $Y=0.745 $X2=0 $Y2=0
cc_243 N_A1_c_245_n N_Y_c_729_n 0.00847255f $X=3.93 $Y=1.49 $X2=0 $Y2=0
cc_244 N_A1_M1036_g N_Y_c_730_n 0.00172847f $X=3.95 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A1_M1037_g N_Y_c_730_n 0.00361507f $X=4.02 $Y=0.745 $X2=0 $Y2=0
cc_246 N_A1_c_245_n N_Y_c_730_n 0.0135341f $X=3.93 $Y=1.49 $X2=0 $Y2=0
cc_247 N_A1_c_247_n N_Y_c_730_n 0.00223721f $X=4.02 $Y=1.49 $X2=0 $Y2=0
cc_248 N_A1_M1002_g N_Y_c_732_n 5.079e-19 $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A1_c_247_n N_Y_c_732_n 3.39537e-19 $X=4.02 $Y=1.49 $X2=0 $Y2=0
cc_250 N_A1_M1004_g N_Y_c_733_n 0.0126232f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_251 N_A1_M1018_g N_Y_c_733_n 0.0101305f $X=3.16 $Y=0.745 $X2=0 $Y2=0
cc_252 N_A1_M1034_g N_Y_c_733_n 0.0119183f $X=3.59 $Y=0.745 $X2=0 $Y2=0
cc_253 N_A1_c_244_n N_Y_c_733_n 0.0436708f $X=2.737 $Y=1.392 $X2=0 $Y2=0
cc_254 N_A1_c_245_n N_Y_c_733_n 0.0145161f $X=3.93 $Y=1.49 $X2=0 $Y2=0
cc_255 N_A1_c_246_n N_Y_c_733_n 0.0199897f $X=2.57 $Y=1.49 $X2=0 $Y2=0
cc_256 N_A1_c_247_n N_Y_c_733_n 0.0147621f $X=4.02 $Y=1.49 $X2=0 $Y2=0
cc_257 N_A1_M1018_g N_Y_c_734_n 0.00180143f $X=3.16 $Y=0.745 $X2=0 $Y2=0
cc_258 N_A1_M1034_g N_Y_c_734_n 0.00980621f $X=3.59 $Y=0.745 $X2=0 $Y2=0
cc_259 N_A1_M1037_g N_Y_c_734_n 0.00883369f $X=4.02 $Y=0.745 $X2=0 $Y2=0
cc_260 N_A1_c_245_n N_Y_c_734_n 0.0261135f $X=3.93 $Y=1.49 $X2=0 $Y2=0
cc_261 N_A1_c_247_n N_Y_c_734_n 0.00285928f $X=4.02 $Y=1.49 $X2=0 $Y2=0
cc_262 N_A1_c_248_n N_Y_c_734_n 8.90145e-19 $X=3.205 $Y=1.392 $X2=0 $Y2=0
cc_263 N_A1_M1002_g N_VPWR_c_850_n 0.0099879f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A1_M1010_g N_VPWR_c_850_n 0.0107197f $X=2.66 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A1_M1026_g N_VPWR_c_850_n 6.33489e-19 $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A1_M1010_g N_VPWR_c_851_n 6.13375e-19 $X=2.66 $Y=2.465 $X2=0 $Y2=0
cc_267 N_A1_M1026_g N_VPWR_c_851_n 0.0101209f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A1_M1036_g N_VPWR_c_851_n 0.00798235f $X=3.95 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A1_M1036_g N_VPWR_c_852_n 0.0054895f $X=3.95 $Y=2.465 $X2=0 $Y2=0
cc_270 N_A1_M1002_g N_VPWR_c_859_n 0.00564095f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_271 N_A1_M1010_g N_VPWR_c_865_n 0.00486043f $X=2.66 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A1_M1026_g N_VPWR_c_865_n 0.00564095f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A1_M1002_g N_VPWR_c_849_n 0.00950825f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_274 N_A1_M1010_g N_VPWR_c_849_n 0.00824727f $X=2.66 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A1_M1026_g N_VPWR_c_849_n 0.00948291f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A1_M1036_g N_VPWR_c_849_n 0.0107218f $X=3.95 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A1_M1004_g N_VGND_c_1000_n 0.00184837f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_278 N_A1_M1004_g N_VGND_c_1005_n 0.00302501f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_279 N_A1_M1018_g N_VGND_c_1005_n 0.00302501f $X=3.16 $Y=0.745 $X2=0 $Y2=0
cc_280 N_A1_M1034_g N_VGND_c_1005_n 0.00302501f $X=3.59 $Y=0.745 $X2=0 $Y2=0
cc_281 N_A1_M1037_g N_VGND_c_1005_n 0.00302501f $X=4.02 $Y=0.745 $X2=0 $Y2=0
cc_282 N_A1_M1004_g N_VGND_c_1011_n 0.0048466f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_283 N_A1_M1018_g N_VGND_c_1011_n 0.00434671f $X=3.16 $Y=0.745 $X2=0 $Y2=0
cc_284 N_A1_M1034_g N_VGND_c_1011_n 0.00433762f $X=3.59 $Y=0.745 $X2=0 $Y2=0
cc_285 N_A1_M1037_g N_VGND_c_1011_n 0.00442601f $X=4.02 $Y=0.745 $X2=0 $Y2=0
cc_286 N_A1_M1004_g N_A_478_65#_c_1114_n 0.0144613f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_287 N_A1_M1018_g N_A_478_65#_c_1114_n 0.0139603f $X=3.16 $Y=0.745 $X2=0 $Y2=0
cc_288 N_A1_M1034_g N_A_478_65#_c_1115_n 0.00913467f $X=3.59 $Y=0.745 $X2=0
+ $Y2=0
cc_289 N_A1_M1037_g N_A_478_65#_c_1115_n 0.011571f $X=4.02 $Y=0.745 $X2=0 $Y2=0
cc_290 N_A2_M1031_g N_A3_M1003_g 0.0237096f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A2_c_332_n N_A3_c_430_n 0.0191224f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_292 N_A2_c_333_n N_A3_c_430_n 3.32475e-19 $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_293 N_A2_c_332_n N_A3_c_431_n 6.45123e-19 $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_294 N_A2_c_333_n N_A3_c_431_n 0.0220316f $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_295 N_A2_M1001_g N_A_30_367#_c_611_n 0.00949266f $X=4.38 $Y=2.465 $X2=0 $Y2=0
cc_296 N_A2_M1012_g N_A_30_367#_c_611_n 6.1646e-19 $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A2_M1001_g N_A_30_367#_c_615_n 0.0113143f $X=4.38 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A2_M1012_g N_A_30_367#_c_615_n 0.0128703f $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A2_c_332_n N_A_30_367#_c_615_n 0.00617296f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_300 N_A2_c_333_n N_A_30_367#_c_615_n 0.00277058f $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_301 N_A2_M1001_g N_A_30_367#_c_619_n 8.38735e-19 $X=4.38 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A2_M1012_g N_A_30_367#_c_619_n 0.00316106f $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A2_M1017_g N_A_30_367#_c_589_n 0.0147477f $X=5.24 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A2_M1031_g N_A_30_367#_c_589_n 0.0119515f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A2_c_332_n N_A_30_367#_c_589_n 0.055998f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_306 N_A2_c_333_n N_A_30_367#_c_589_n 0.00661192f $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_307 N_A2_M1012_g N_A_30_367#_c_590_n 0.00389941f $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_308 N_A2_c_332_n N_A_30_367#_c_590_n 0.0228757f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_309 N_A2_c_333_n N_A_30_367#_c_590_n 0.0027894f $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_310 N_A2_M1017_g N_A_30_367#_c_628_n 0.00100832f $X=5.24 $Y=2.465 $X2=0 $Y2=0
cc_311 N_A2_M1031_g N_A_30_367#_c_628_n 0.0154665f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_312 N_A2_M1001_g N_A_30_367#_c_612_n 7.53639e-19 $X=4.38 $Y=2.465 $X2=0 $Y2=0
cc_313 N_A2_M1012_g N_A_30_367#_c_631_n 0.0021907f $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A2_M1031_g N_A_30_367#_c_596_n 0.0016758f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_315 N_A2_c_332_n N_A_30_367#_c_596_n 0.00799152f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_316 N_A2_c_333_n N_A_30_367#_c_596_n 0.00167044f $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_317 N_A2_M1001_g N_Y_c_735_n 0.00785493f $X=4.38 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A2_M1012_g N_Y_c_735_n 7.08049e-19 $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_319 N_A2_c_325_n N_Y_c_729_n 0.00464422f $X=4.53 $Y=1.275 $X2=0 $Y2=0
cc_320 N_A2_c_327_n N_Y_c_729_n 6.34514e-19 $X=4.96 $Y=1.275 $X2=0 $Y2=0
cc_321 N_A2_c_332_n N_Y_c_729_n 0.00339586f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_322 N_A2_M1001_g N_Y_c_730_n 0.00421425f $X=4.38 $Y=2.465 $X2=0 $Y2=0
cc_323 N_A2_c_325_n N_Y_c_730_n 3.53048e-19 $X=4.53 $Y=1.275 $X2=0 $Y2=0
cc_324 N_A2_M1012_g N_Y_c_730_n 8.74475e-19 $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_325 N_A2_c_332_n N_Y_c_730_n 0.0270831f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_326 N_A2_c_333_n N_Y_c_730_n 0.0133867f $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_327 N_A2_c_325_n N_Y_c_734_n 6.21942e-19 $X=4.53 $Y=1.275 $X2=0 $Y2=0
cc_328 N_A2_M1001_g N_VPWR_c_852_n 0.0054895f $X=4.38 $Y=2.465 $X2=0 $Y2=0
cc_329 N_A2_M1001_g N_VPWR_c_853_n 0.001552f $X=4.38 $Y=2.465 $X2=0 $Y2=0
cc_330 N_A2_M1012_g N_VPWR_c_853_n 0.00165477f $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_331 N_A2_M1017_g N_VPWR_c_854_n 0.00787607f $X=5.24 $Y=2.465 $X2=0 $Y2=0
cc_332 N_A2_M1031_g N_VPWR_c_854_n 0.00782667f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_333 N_A2_M1031_g N_VPWR_c_855_n 8.24495e-19 $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A2_M1012_g N_VPWR_c_866_n 0.00585385f $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_335 N_A2_M1017_g N_VPWR_c_866_n 0.00585385f $X=5.24 $Y=2.465 $X2=0 $Y2=0
cc_336 N_A2_M1031_g N_VPWR_c_867_n 0.0054895f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_337 N_A2_M1001_g N_VPWR_c_849_n 0.00979102f $X=4.38 $Y=2.465 $X2=0 $Y2=0
cc_338 N_A2_M1012_g N_VPWR_c_849_n 0.0105361f $X=4.81 $Y=2.465 $X2=0 $Y2=0
cc_339 N_A2_M1017_g N_VPWR_c_849_n 0.0111403f $X=5.24 $Y=2.465 $X2=0 $Y2=0
cc_340 N_A2_M1031_g N_VPWR_c_849_n 0.0103133f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_341 N_A2_c_325_n N_VGND_c_1005_n 0.00302473f $X=4.53 $Y=1.275 $X2=0 $Y2=0
cc_342 N_A2_c_327_n N_VGND_c_1005_n 0.00302501f $X=4.96 $Y=1.275 $X2=0 $Y2=0
cc_343 N_A2_c_329_n N_VGND_c_1005_n 0.00302501f $X=5.39 $Y=1.275 $X2=0 $Y2=0
cc_344 N_A2_c_330_n N_VGND_c_1005_n 0.00302501f $X=5.82 $Y=1.275 $X2=0 $Y2=0
cc_345 N_A2_c_325_n N_VGND_c_1011_n 0.004426f $X=4.53 $Y=1.275 $X2=0 $Y2=0
cc_346 N_A2_c_327_n N_VGND_c_1011_n 0.00433762f $X=4.96 $Y=1.275 $X2=0 $Y2=0
cc_347 N_A2_c_329_n N_VGND_c_1011_n 0.00434671f $X=5.39 $Y=1.275 $X2=0 $Y2=0
cc_348 N_A2_c_330_n N_VGND_c_1011_n 0.0048466f $X=5.82 $Y=1.275 $X2=0 $Y2=0
cc_349 N_A2_c_325_n N_A_478_65#_c_1126_n 0.0073239f $X=4.53 $Y=1.275 $X2=0 $Y2=0
cc_350 N_A2_c_327_n N_A_478_65#_c_1126_n 4.46945e-19 $X=4.96 $Y=1.275 $X2=0
+ $Y2=0
cc_351 N_A2_c_333_n N_A_478_65#_c_1126_n 6.02007e-19 $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_352 N_A2_c_329_n N_A_478_65#_c_1116_n 0.00904079f $X=5.39 $Y=1.275 $X2=0
+ $Y2=0
cc_353 N_A2_c_329_n N_A_478_65#_c_1117_n 0.00467288f $X=5.39 $Y=1.275 $X2=0
+ $Y2=0
cc_354 N_A2_c_330_n N_A_478_65#_c_1117_n 0.0143942f $X=5.82 $Y=1.275 $X2=0 $Y2=0
cc_355 N_A2_c_325_n N_A_478_65#_c_1119_n 0.00152212f $X=4.53 $Y=1.275 $X2=0
+ $Y2=0
cc_356 N_A2_c_325_n N_A_478_65#_c_1120_n 0.0102372f $X=4.53 $Y=1.275 $X2=0 $Y2=0
cc_357 N_A2_c_327_n N_A_478_65#_c_1120_n 0.00921399f $X=4.96 $Y=1.275 $X2=0
+ $Y2=0
cc_358 N_A2_c_327_n N_A_921_65#_c_1160_n 0.0108854f $X=4.96 $Y=1.275 $X2=0 $Y2=0
cc_359 N_A2_c_329_n N_A_921_65#_c_1160_n 0.00951259f $X=5.39 $Y=1.275 $X2=0
+ $Y2=0
cc_360 N_A2_c_330_n N_A_921_65#_c_1160_n 0.012039f $X=5.82 $Y=1.275 $X2=0 $Y2=0
cc_361 N_A2_c_332_n N_A_921_65#_c_1160_n 0.0725393f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_362 N_A2_c_333_n N_A_921_65#_c_1160_n 0.00150571f $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_363 N_A2_c_327_n N_A_921_65#_c_1166_n 0.00530459f $X=4.96 $Y=1.275 $X2=0
+ $Y2=0
cc_364 N_A2_c_329_n N_A_921_65#_c_1166_n 8.74229e-19 $X=5.39 $Y=1.275 $X2=0
+ $Y2=0
cc_365 N_A2_c_332_n N_A_921_65#_c_1166_n 0.0180857f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_366 N_A2_c_333_n N_A_921_65#_c_1166_n 6.09012e-19 $X=5.83 $Y=1.44 $X2=0 $Y2=0
cc_367 N_A2_c_330_n N_A_1291_65#_c_1215_n 9.24112e-19 $X=5.82 $Y=1.275 $X2=0
+ $Y2=0
cc_368 N_A3_M1033_g N_A4_M1000_g 0.0229538f $X=8.07 $Y=2.465 $X2=0 $Y2=0
cc_369 N_A3_c_427_n N_A4_c_512_n 0.0156839f $X=8.085 $Y=1.275 $X2=0 $Y2=0
cc_370 N_A3_c_427_n A4 0.00182063f $X=8.085 $Y=1.275 $X2=0 $Y2=0
cc_371 N_A3_c_428_n A4 0.0162683f $X=8.05 $Y=1.44 $X2=0 $Y2=0
cc_372 N_A3_c_431_n A4 9.00522e-19 $X=8.085 $Y=1.44 $X2=0 $Y2=0
cc_373 N_A3_c_428_n N_A4_c_520_n 2.83054e-19 $X=8.05 $Y=1.44 $X2=0 $Y2=0
cc_374 N_A3_c_431_n N_A4_c_520_n 0.0220943f $X=8.085 $Y=1.44 $X2=0 $Y2=0
cc_375 N_A3_M1003_g N_A_30_367#_c_591_n 0.0132004f $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_376 N_A3_M1019_g N_A_30_367#_c_591_n 0.013222f $X=6.69 $Y=2.465 $X2=0 $Y2=0
cc_377 N_A3_c_430_n N_A_30_367#_c_591_n 0.0451055f $X=7.37 $Y=1.44 $X2=0 $Y2=0
cc_378 N_A3_c_431_n N_A_30_367#_c_591_n 0.00229528f $X=8.085 $Y=1.44 $X2=0 $Y2=0
cc_379 N_A3_M1032_g N_A_30_367#_c_592_n 0.0152626f $X=7.12 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A3_M1033_g N_A_30_367#_c_592_n 0.015241f $X=8.07 $Y=2.465 $X2=0 $Y2=0
cc_381 N_A3_c_428_n N_A_30_367#_c_592_n 0.0473058f $X=8.05 $Y=1.44 $X2=0 $Y2=0
cc_382 A3 N_A_30_367#_c_592_n 0.0144903f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_383 N_A3_c_430_n N_A_30_367#_c_592_n 0.0249399f $X=7.37 $Y=1.44 $X2=0 $Y2=0
cc_384 N_A3_c_431_n N_A_30_367#_c_592_n 0.0171017f $X=8.085 $Y=1.44 $X2=0 $Y2=0
cc_385 N_A3_c_430_n N_A_30_367#_c_597_n 0.015808f $X=7.37 $Y=1.44 $X2=0 $Y2=0
cc_386 N_A3_c_431_n N_A_30_367#_c_597_n 0.0027894f $X=8.085 $Y=1.44 $X2=0 $Y2=0
cc_387 N_A3_c_428_n N_A_30_367#_c_598_n 0.00205753f $X=8.05 $Y=1.44 $X2=0 $Y2=0
cc_388 N_A3_c_431_n N_A_30_367#_c_598_n 5.96587e-19 $X=8.085 $Y=1.44 $X2=0 $Y2=0
cc_389 N_A3_M1003_g N_VPWR_c_855_n 0.0143077f $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_390 N_A3_M1019_g N_VPWR_c_855_n 0.0141279f $X=6.69 $Y=2.465 $X2=0 $Y2=0
cc_391 N_A3_M1032_g N_VPWR_c_855_n 7.24342e-19 $X=7.12 $Y=2.465 $X2=0 $Y2=0
cc_392 N_A3_M1019_g N_VPWR_c_856_n 7.37829e-19 $X=6.69 $Y=2.465 $X2=0 $Y2=0
cc_393 N_A3_M1032_g N_VPWR_c_856_n 0.0156947f $X=7.12 $Y=2.465 $X2=0 $Y2=0
cc_394 N_A3_M1033_g N_VPWR_c_856_n 0.0156947f $X=8.07 $Y=2.465 $X2=0 $Y2=0
cc_395 N_A3_M1033_g N_VPWR_c_857_n 7.24342e-19 $X=8.07 $Y=2.465 $X2=0 $Y2=0
cc_396 N_A3_M1033_g N_VPWR_c_861_n 0.00486043f $X=8.07 $Y=2.465 $X2=0 $Y2=0
cc_397 N_A3_M1003_g N_VPWR_c_867_n 0.00486043f $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_398 N_A3_M1019_g N_VPWR_c_868_n 0.00486043f $X=6.69 $Y=2.465 $X2=0 $Y2=0
cc_399 N_A3_M1032_g N_VPWR_c_868_n 0.00486043f $X=7.12 $Y=2.465 $X2=0 $Y2=0
cc_400 N_A3_M1003_g N_VPWR_c_849_n 0.0082726f $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_401 N_A3_M1019_g N_VPWR_c_849_n 0.00824727f $X=6.69 $Y=2.465 $X2=0 $Y2=0
cc_402 N_A3_M1032_g N_VPWR_c_849_n 0.00824727f $X=7.12 $Y=2.465 $X2=0 $Y2=0
cc_403 N_A3_M1033_g N_VPWR_c_849_n 0.0082726f $X=8.07 $Y=2.465 $X2=0 $Y2=0
cc_404 N_A3_c_427_n N_VGND_c_1001_n 5.15399e-19 $X=8.085 $Y=1.275 $X2=0 $Y2=0
cc_405 N_A3_c_422_n N_VGND_c_1005_n 0.00302501f $X=6.795 $Y=1.275 $X2=0 $Y2=0
cc_406 N_A3_c_424_n N_VGND_c_1005_n 0.00302501f $X=7.225 $Y=1.275 $X2=0 $Y2=0
cc_407 N_A3_c_425_n N_VGND_c_1005_n 0.00302501f $X=7.655 $Y=1.275 $X2=0 $Y2=0
cc_408 N_A3_c_427_n N_VGND_c_1005_n 0.00302501f $X=8.085 $Y=1.275 $X2=0 $Y2=0
cc_409 N_A3_c_422_n N_VGND_c_1011_n 0.00483751f $X=6.795 $Y=1.275 $X2=0 $Y2=0
cc_410 N_A3_c_424_n N_VGND_c_1011_n 0.00433762f $X=7.225 $Y=1.275 $X2=0 $Y2=0
cc_411 N_A3_c_425_n N_VGND_c_1011_n 0.00433762f $X=7.655 $Y=1.275 $X2=0 $Y2=0
cc_412 N_A3_c_427_n N_VGND_c_1011_n 0.00435646f $X=8.085 $Y=1.275 $X2=0 $Y2=0
cc_413 N_A3_c_422_n N_A_921_65#_c_1160_n 0.0131891f $X=6.795 $Y=1.275 $X2=0
+ $Y2=0
cc_414 N_A3_c_430_n N_A_921_65#_c_1160_n 0.0310279f $X=7.37 $Y=1.44 $X2=0 $Y2=0
cc_415 N_A3_c_431_n N_A_921_65#_c_1160_n 0.013036f $X=8.085 $Y=1.44 $X2=0 $Y2=0
cc_416 N_A3_c_424_n N_A_921_65#_c_1173_n 0.00960676f $X=7.225 $Y=1.275 $X2=0
+ $Y2=0
cc_417 N_A3_c_425_n N_A_921_65#_c_1173_n 0.0102376f $X=7.655 $Y=1.275 $X2=0
+ $Y2=0
cc_418 N_A3_c_428_n N_A_921_65#_c_1173_n 0.00549903f $X=8.05 $Y=1.44 $X2=0 $Y2=0
cc_419 A3 N_A_921_65#_c_1173_n 0.0130159f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_420 N_A3_c_430_n N_A_921_65#_c_1173_n 0.0061266f $X=7.37 $Y=1.44 $X2=0 $Y2=0
cc_421 N_A3_c_431_n N_A_921_65#_c_1173_n 5.20335e-19 $X=8.085 $Y=1.44 $X2=0
+ $Y2=0
cc_422 N_A3_c_422_n N_A_921_65#_c_1179_n 0.0147554f $X=6.795 $Y=1.275 $X2=0
+ $Y2=0
cc_423 N_A3_c_424_n N_A_921_65#_c_1179_n 0.00764111f $X=7.225 $Y=1.275 $X2=0
+ $Y2=0
cc_424 N_A3_c_425_n N_A_921_65#_c_1179_n 9.976e-19 $X=7.655 $Y=1.275 $X2=0 $Y2=0
cc_425 N_A3_c_430_n N_A_921_65#_c_1179_n 0.0210368f $X=7.37 $Y=1.44 $X2=0 $Y2=0
cc_426 N_A3_c_431_n N_A_921_65#_c_1179_n 0.0028345f $X=8.085 $Y=1.44 $X2=0 $Y2=0
cc_427 N_A3_c_424_n N_A_921_65#_c_1184_n 9.976e-19 $X=7.225 $Y=1.275 $X2=0 $Y2=0
cc_428 N_A3_c_425_n N_A_921_65#_c_1184_n 0.00768006f $X=7.655 $Y=1.275 $X2=0
+ $Y2=0
cc_429 N_A3_c_427_n N_A_921_65#_c_1184_n 0.00708277f $X=8.085 $Y=1.275 $X2=0
+ $Y2=0
cc_430 N_A3_c_428_n N_A_921_65#_c_1184_n 0.0175801f $X=8.05 $Y=1.44 $X2=0 $Y2=0
cc_431 N_A3_c_431_n N_A_921_65#_c_1184_n 0.00255041f $X=8.085 $Y=1.44 $X2=0
+ $Y2=0
cc_432 A3 N_A_1291_65#_M1009_d 0.00181594f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_433 N_A3_c_422_n N_A_1291_65#_c_1210_n 0.00930868f $X=6.795 $Y=1.275 $X2=0
+ $Y2=0
cc_434 N_A3_c_424_n N_A_1291_65#_c_1210_n 0.00859511f $X=7.225 $Y=1.275 $X2=0
+ $Y2=0
cc_435 N_A3_c_425_n N_A_1291_65#_c_1211_n 0.00859511f $X=7.655 $Y=1.275 $X2=0
+ $Y2=0
cc_436 N_A3_c_427_n N_A_1291_65#_c_1211_n 0.0117786f $X=8.085 $Y=1.275 $X2=0
+ $Y2=0
cc_437 N_A3_c_422_n N_A_1291_65#_c_1215_n 6.7916e-19 $X=6.795 $Y=1.275 $X2=0
+ $Y2=0
cc_438 N_A4_M1000_g N_A_30_367#_c_593_n 0.0132004f $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_439 N_A4_M1011_g N_A_30_367#_c_593_n 0.013222f $X=8.93 $Y=2.465 $X2=0 $Y2=0
cc_440 A4 N_A_30_367#_c_593_n 0.0463753f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_441 N_A4_c_520_n N_A_30_367#_c_593_n 0.00235568f $X=9.88 $Y=1.44 $X2=0 $Y2=0
cc_442 N_A4_M1015_g N_A_30_367#_c_594_n 0.013222f $X=9.36 $Y=2.465 $X2=0 $Y2=0
cc_443 N_A4_M1024_g N_A_30_367#_c_594_n 0.0138663f $X=9.79 $Y=2.465 $X2=0 $Y2=0
cc_444 A4 N_A_30_367#_c_594_n 0.0718815f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_445 N_A4_c_520_n N_A_30_367#_c_594_n 0.00342599f $X=9.88 $Y=1.44 $X2=0 $Y2=0
cc_446 N_A4_c_521_n N_A_30_367#_c_594_n 0.0062045f $X=10.29 $Y=1.44 $X2=0 $Y2=0
cc_447 A4 N_A_30_367#_c_599_n 0.0161959f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_448 N_A4_c_520_n N_A_30_367#_c_599_n 0.0024468f $X=9.88 $Y=1.44 $X2=0 $Y2=0
cc_449 N_A4_M1000_g N_VPWR_c_856_n 7.37829e-19 $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_450 N_A4_M1000_g N_VPWR_c_857_n 0.0141279f $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_451 N_A4_M1011_g N_VPWR_c_857_n 0.0141279f $X=8.93 $Y=2.465 $X2=0 $Y2=0
cc_452 N_A4_M1015_g N_VPWR_c_857_n 7.24342e-19 $X=9.36 $Y=2.465 $X2=0 $Y2=0
cc_453 N_A4_M1011_g N_VPWR_c_858_n 7.24342e-19 $X=8.93 $Y=2.465 $X2=0 $Y2=0
cc_454 N_A4_M1015_g N_VPWR_c_858_n 0.0141279f $X=9.36 $Y=2.465 $X2=0 $Y2=0
cc_455 N_A4_M1024_g N_VPWR_c_858_n 0.0161027f $X=9.79 $Y=2.465 $X2=0 $Y2=0
cc_456 N_A4_M1000_g N_VPWR_c_861_n 0.00486043f $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_457 N_A4_M1011_g N_VPWR_c_863_n 0.00486043f $X=8.93 $Y=2.465 $X2=0 $Y2=0
cc_458 N_A4_M1015_g N_VPWR_c_863_n 0.00486043f $X=9.36 $Y=2.465 $X2=0 $Y2=0
cc_459 N_A4_M1024_g N_VPWR_c_869_n 0.00486043f $X=9.79 $Y=2.465 $X2=0 $Y2=0
cc_460 N_A4_M1000_g N_VPWR_c_849_n 0.0082726f $X=8.5 $Y=2.465 $X2=0 $Y2=0
cc_461 N_A4_M1011_g N_VPWR_c_849_n 0.00824727f $X=8.93 $Y=2.465 $X2=0 $Y2=0
cc_462 N_A4_M1015_g N_VPWR_c_849_n 0.00824727f $X=9.36 $Y=2.465 $X2=0 $Y2=0
cc_463 N_A4_M1024_g N_VPWR_c_849_n 0.00936453f $X=9.79 $Y=2.465 $X2=0 $Y2=0
cc_464 N_A4_c_512_n N_VGND_c_1001_n 0.00854664f $X=8.515 $Y=1.275 $X2=0 $Y2=0
cc_465 N_A4_c_514_n N_VGND_c_1001_n 0.00857574f $X=8.945 $Y=1.275 $X2=0 $Y2=0
cc_466 N_A4_c_516_n N_VGND_c_1001_n 4.75255e-19 $X=9.375 $Y=1.275 $X2=0 $Y2=0
cc_467 N_A4_c_514_n N_VGND_c_1002_n 4.75255e-19 $X=8.945 $Y=1.275 $X2=0 $Y2=0
cc_468 N_A4_c_516_n N_VGND_c_1002_n 0.00857574f $X=9.375 $Y=1.275 $X2=0 $Y2=0
cc_469 N_A4_c_518_n N_VGND_c_1002_n 0.0110167f $X=9.805 $Y=1.275 $X2=0 $Y2=0
cc_470 N_A4_c_512_n N_VGND_c_1005_n 0.00414769f $X=8.515 $Y=1.275 $X2=0 $Y2=0
cc_471 N_A4_c_514_n N_VGND_c_1007_n 0.00414769f $X=8.945 $Y=1.275 $X2=0 $Y2=0
cc_472 N_A4_c_516_n N_VGND_c_1007_n 0.00414769f $X=9.375 $Y=1.275 $X2=0 $Y2=0
cc_473 N_A4_c_518_n N_VGND_c_1010_n 0.00414769f $X=9.805 $Y=1.275 $X2=0 $Y2=0
cc_474 N_A4_c_512_n N_VGND_c_1011_n 0.00419085f $X=8.515 $Y=1.275 $X2=0 $Y2=0
cc_475 N_A4_c_514_n N_VGND_c_1011_n 0.00418111f $X=8.945 $Y=1.275 $X2=0 $Y2=0
cc_476 N_A4_c_516_n N_VGND_c_1011_n 0.00418111f $X=9.375 $Y=1.275 $X2=0 $Y2=0
cc_477 N_A4_c_518_n N_VGND_c_1011_n 0.00460855f $X=9.805 $Y=1.275 $X2=0 $Y2=0
cc_478 N_A4_c_512_n N_A_921_65#_c_1184_n 4.9625e-19 $X=8.515 $Y=1.275 $X2=0
+ $Y2=0
cc_479 N_A4_c_512_n N_A_1291_65#_c_1211_n 5.73473e-19 $X=8.515 $Y=1.275 $X2=0
+ $Y2=0
cc_480 N_A4_c_512_n N_A_1291_65#_c_1225_n 0.00969264f $X=8.515 $Y=1.275 $X2=0
+ $Y2=0
cc_481 N_A4_c_514_n N_A_1291_65#_c_1225_n 0.00964608f $X=8.945 $Y=1.275 $X2=0
+ $Y2=0
cc_482 A4 N_A_1291_65#_c_1225_n 0.0421429f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_483 N_A4_c_520_n N_A_1291_65#_c_1225_n 5.77176e-19 $X=9.88 $Y=1.44 $X2=0
+ $Y2=0
cc_484 N_A4_c_516_n N_A_1291_65#_c_1213_n 0.00969264f $X=9.375 $Y=1.275 $X2=0
+ $Y2=0
cc_485 N_A4_c_518_n N_A_1291_65#_c_1213_n 0.00969264f $X=9.805 $Y=1.275 $X2=0
+ $Y2=0
cc_486 A4 N_A_1291_65#_c_1213_n 0.0658325f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_487 N_A4_c_520_n N_A_1291_65#_c_1213_n 5.77176e-19 $X=9.88 $Y=1.44 $X2=0
+ $Y2=0
cc_488 N_A4_c_521_n N_A_1291_65#_c_1213_n 0.00166517f $X=10.29 $Y=1.44 $X2=0
+ $Y2=0
cc_489 N_A4_c_518_n N_A_1291_65#_c_1214_n 3.18679e-19 $X=9.805 $Y=1.275 $X2=0
+ $Y2=0
cc_490 A4 N_A_1291_65#_c_1235_n 0.015637f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_491 N_A4_c_520_n N_A_1291_65#_c_1235_n 6.51443e-19 $X=9.88 $Y=1.44 $X2=0
+ $Y2=0
cc_492 N_A_30_367#_c_603_n N_Y_M1007_s 0.00332344f $X=1.04 $Y=2.99 $X2=0 $Y2=0
cc_493 N_A_30_367#_c_605_n N_Y_M1023_s 0.00332344f $X=1.9 $Y=2.99 $X2=0 $Y2=0
cc_494 N_A_30_367#_c_588_n N_Y_c_738_n 0.0345065f $X=0.275 $Y=1.99 $X2=0 $Y2=0
cc_495 N_A_30_367#_c_603_n N_Y_c_738_n 0.0159805f $X=1.04 $Y=2.99 $X2=0 $Y2=0
cc_496 N_A_30_367#_c_605_n N_Y_c_751_n 0.0159805f $X=1.9 $Y=2.99 $X2=0 $Y2=0
cc_497 N_A_30_367#_M1027_d N_Y_c_735_n 0.00177068f $X=1.855 $Y=1.835 $X2=0 $Y2=0
cc_498 N_A_30_367#_M1010_s N_Y_c_735_n 0.00177068f $X=2.735 $Y=1.835 $X2=0 $Y2=0
cc_499 N_A_30_367#_M1036_s N_Y_c_735_n 0.00177068f $X=4.025 $Y=1.835 $X2=0 $Y2=0
cc_500 N_A_30_367#_c_668_p N_Y_c_735_n 0.0136074f $X=2.005 $Y=2.285 $X2=0 $Y2=0
cc_501 N_A_30_367#_c_607_n N_Y_c_735_n 0.0342127f $X=2.78 $Y=2.195 $X2=0 $Y2=0
cc_502 N_A_30_367#_c_609_n N_Y_c_735_n 0.0626544f $X=4 $Y=2.195 $X2=0 $Y2=0
cc_503 N_A_30_367#_c_615_n N_Y_c_735_n 0.0094487f $X=4.86 $Y=2.195 $X2=0 $Y2=0
cc_504 N_A_30_367#_c_619_n N_Y_c_735_n 3.71595e-19 $X=5.025 $Y=1.98 $X2=0 $Y2=0
cc_505 N_A_30_367#_c_590_n N_Y_c_735_n 0.00710829f $X=5.13 $Y=1.84 $X2=0 $Y2=0
cc_506 N_A_30_367#_c_674_p N_Y_c_735_n 0.0136074f $X=2.875 $Y=2.27 $X2=0 $Y2=0
cc_507 N_A_30_367#_c_612_n N_Y_c_735_n 0.0175583f $X=4.165 $Y=2.22 $X2=0 $Y2=0
cc_508 N_A_30_367#_c_676_p N_Y_c_731_n 0.0146502f $X=1.135 $Y=2.125 $X2=0 $Y2=0
cc_509 N_A_30_367#_c_607_n N_VPWR_M1002_d 0.003805f $X=2.78 $Y=2.195 $X2=-0.19
+ $Y2=1.655
cc_510 N_A_30_367#_c_609_n N_VPWR_M1026_d 0.0155993f $X=4 $Y=2.195 $X2=0 $Y2=0
cc_511 N_A_30_367#_c_615_n N_VPWR_M1001_s 0.00519719f $X=4.86 $Y=2.195 $X2=0
+ $Y2=0
cc_512 N_A_30_367#_c_589_n N_VPWR_M1017_s 0.00394368f $X=5.88 $Y=1.84 $X2=0
+ $Y2=0
cc_513 N_A_30_367#_c_591_n N_VPWR_M1003_s 0.00180746f $X=6.81 $Y=1.84 $X2=0
+ $Y2=0
cc_514 N_A_30_367#_c_592_n N_VPWR_M1032_s 0.00963689f $X=8.19 $Y=1.84 $X2=0
+ $Y2=0
cc_515 N_A_30_367#_c_593_n N_VPWR_M1000_s 0.00180746f $X=9.05 $Y=1.84 $X2=0
+ $Y2=0
cc_516 N_A_30_367#_c_594_n N_VPWR_M1015_s 0.00180746f $X=9.91 $Y=1.84 $X2=0
+ $Y2=0
cc_517 N_A_30_367#_c_607_n N_VPWR_c_850_n 0.0172482f $X=2.78 $Y=2.195 $X2=0
+ $Y2=0
cc_518 N_A_30_367#_c_609_n N_VPWR_c_851_n 0.0468916f $X=4 $Y=2.195 $X2=0 $Y2=0
cc_519 N_A_30_367#_c_611_n N_VPWR_c_852_n 0.0189236f $X=4.165 $Y=2.97 $X2=0
+ $Y2=0
cc_520 N_A_30_367#_c_615_n N_VPWR_c_853_n 0.0135577f $X=4.86 $Y=2.195 $X2=0
+ $Y2=0
cc_521 N_A_30_367#_c_589_n N_VPWR_c_854_n 0.0254128f $X=5.88 $Y=1.84 $X2=0 $Y2=0
cc_522 N_A_30_367#_c_591_n N_VPWR_c_855_n 0.0163515f $X=6.81 $Y=1.84 $X2=0 $Y2=0
cc_523 N_A_30_367#_c_592_n N_VPWR_c_856_n 0.0568873f $X=8.19 $Y=1.84 $X2=0 $Y2=0
cc_524 N_A_30_367#_c_593_n N_VPWR_c_857_n 0.0163515f $X=9.05 $Y=1.84 $X2=0 $Y2=0
cc_525 N_A_30_367#_c_594_n N_VPWR_c_858_n 0.0163515f $X=9.91 $Y=1.84 $X2=0 $Y2=0
cc_526 N_A_30_367#_c_587_n N_VPWR_c_859_n 0.0179183f $X=0.24 $Y=2.905 $X2=0
+ $Y2=0
cc_527 N_A_30_367#_c_603_n N_VPWR_c_859_n 0.0361172f $X=1.04 $Y=2.99 $X2=0 $Y2=0
cc_528 N_A_30_367#_c_605_n N_VPWR_c_859_n 0.049324f $X=1.9 $Y=2.99 $X2=0 $Y2=0
cc_529 N_A_30_367#_c_697_p N_VPWR_c_859_n 0.0125234f $X=1.135 $Y=2.91 $X2=0
+ $Y2=0
cc_530 N_A_30_367#_c_698_p N_VPWR_c_861_n 0.0124525f $X=8.285 $Y=1.98 $X2=0
+ $Y2=0
cc_531 N_A_30_367#_c_699_p N_VPWR_c_863_n 0.0124525f $X=9.145 $Y=1.98 $X2=0
+ $Y2=0
cc_532 N_A_30_367#_c_674_p N_VPWR_c_865_n 0.0131621f $X=2.875 $Y=2.27 $X2=0
+ $Y2=0
cc_533 N_A_30_367#_c_701_p N_VPWR_c_866_n 0.0142265f $X=5.025 $Y=2.43 $X2=0
+ $Y2=0
cc_534 N_A_30_367#_c_628_n N_VPWR_c_867_n 0.015688f $X=6.045 $Y=1.98 $X2=0 $Y2=0
cc_535 N_A_30_367#_c_703_p N_VPWR_c_868_n 0.0124525f $X=6.905 $Y=1.98 $X2=0
+ $Y2=0
cc_536 N_A_30_367#_c_595_n N_VPWR_c_869_n 0.0178111f $X=10.005 $Y=1.98 $X2=0
+ $Y2=0
cc_537 N_A_30_367#_M1007_d N_VPWR_c_849_n 0.00215161f $X=0.15 $Y=1.835 $X2=0
+ $Y2=0
cc_538 N_A_30_367#_M1013_d N_VPWR_c_849_n 0.00223565f $X=0.995 $Y=1.835 $X2=0
+ $Y2=0
cc_539 N_A_30_367#_M1027_d N_VPWR_c_849_n 0.00307052f $X=1.855 $Y=1.835 $X2=0
+ $Y2=0
cc_540 N_A_30_367#_M1010_s N_VPWR_c_849_n 0.00467071f $X=2.735 $Y=1.835 $X2=0
+ $Y2=0
cc_541 N_A_30_367#_M1036_s N_VPWR_c_849_n 0.00223559f $X=4.025 $Y=1.835 $X2=0
+ $Y2=0
cc_542 N_A_30_367#_M1012_d N_VPWR_c_849_n 0.00362709f $X=4.885 $Y=1.835 $X2=0
+ $Y2=0
cc_543 N_A_30_367#_M1031_d N_VPWR_c_849_n 0.00380103f $X=5.905 $Y=1.835 $X2=0
+ $Y2=0
cc_544 N_A_30_367#_M1019_d N_VPWR_c_849_n 0.00536646f $X=6.765 $Y=1.835 $X2=0
+ $Y2=0
cc_545 N_A_30_367#_M1033_d N_VPWR_c_849_n 0.00536646f $X=8.145 $Y=1.835 $X2=0
+ $Y2=0
cc_546 N_A_30_367#_M1011_d N_VPWR_c_849_n 0.00536646f $X=9.005 $Y=1.835 $X2=0
+ $Y2=0
cc_547 N_A_30_367#_M1024_d N_VPWR_c_849_n 0.00371702f $X=9.865 $Y=1.835 $X2=0
+ $Y2=0
cc_548 N_A_30_367#_c_587_n N_VPWR_c_849_n 0.0101029f $X=0.24 $Y=2.905 $X2=0
+ $Y2=0
cc_549 N_A_30_367#_c_603_n N_VPWR_c_849_n 0.023676f $X=1.04 $Y=2.99 $X2=0 $Y2=0
cc_550 N_A_30_367#_c_605_n N_VPWR_c_849_n 0.0318369f $X=1.9 $Y=2.99 $X2=0 $Y2=0
cc_551 N_A_30_367#_c_611_n N_VPWR_c_849_n 0.0123859f $X=4.165 $Y=2.97 $X2=0
+ $Y2=0
cc_552 N_A_30_367#_c_701_p N_VPWR_c_849_n 0.00925289f $X=5.025 $Y=2.43 $X2=0
+ $Y2=0
cc_553 N_A_30_367#_c_628_n N_VPWR_c_849_n 0.00984745f $X=6.045 $Y=1.98 $X2=0
+ $Y2=0
cc_554 N_A_30_367#_c_703_p N_VPWR_c_849_n 0.00730901f $X=6.905 $Y=1.98 $X2=0
+ $Y2=0
cc_555 N_A_30_367#_c_698_p N_VPWR_c_849_n 0.00730901f $X=8.285 $Y=1.98 $X2=0
+ $Y2=0
cc_556 N_A_30_367#_c_699_p N_VPWR_c_849_n 0.00730901f $X=9.145 $Y=1.98 $X2=0
+ $Y2=0
cc_557 N_A_30_367#_c_595_n N_VPWR_c_849_n 0.0100304f $X=10.005 $Y=1.98 $X2=0
+ $Y2=0
cc_558 N_A_30_367#_c_697_p N_VPWR_c_849_n 0.00738676f $X=1.135 $Y=2.91 $X2=0
+ $Y2=0
cc_559 N_A_30_367#_c_674_p N_VPWR_c_849_n 0.00808656f $X=2.875 $Y=2.27 $X2=0
+ $Y2=0
cc_560 N_Y_c_735_n N_VPWR_M1002_d 0.00198885f $X=4.265 $Y=1.84 $X2=-0.19
+ $Y2=-0.245
cc_561 N_Y_c_735_n N_VPWR_M1026_d 0.00829077f $X=4.265 $Y=1.84 $X2=0 $Y2=0
cc_562 N_Y_M1007_s N_VPWR_c_849_n 0.00225186f $X=0.565 $Y=1.835 $X2=0 $Y2=0
cc_563 N_Y_M1023_s N_VPWR_c_849_n 0.00225186f $X=1.425 $Y=1.835 $X2=0 $Y2=0
cc_564 N_Y_c_741_n N_VGND_M1021_s 0.00328468f $X=1.455 $Y=0.947 $X2=0 $Y2=0
cc_565 N_Y_c_733_n N_VGND_M1039_s 0.0103623f $X=3.64 $Y=0.927 $X2=0 $Y2=0
cc_566 N_Y_c_741_n N_VGND_c_999_n 0.016817f $X=1.455 $Y=0.947 $X2=0 $Y2=0
cc_567 N_Y_c_733_n N_VGND_c_1000_n 0.0218745f $X=3.64 $Y=0.927 $X2=0 $Y2=0
cc_568 N_Y_c_831_p N_VGND_c_1003_n 0.0124525f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_569 N_Y_c_832_p N_VGND_c_1009_n 0.0124525f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_570 N_Y_M1014_d N_VGND_c_1011_n 0.00409469f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_571 N_Y_M1022_d N_VGND_c_1011_n 0.00279659f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_572 N_Y_c_832_p N_VGND_c_1011_n 0.00730901f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_573 N_Y_c_741_n N_VGND_c_1011_n 0.0108126f $X=1.455 $Y=0.947 $X2=0 $Y2=0
cc_574 N_Y_c_831_p N_VGND_c_1011_n 0.00730901f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_575 N_Y_c_733_n N_VGND_c_1011_n 0.015873f $X=3.64 $Y=0.927 $X2=0 $Y2=0
cc_576 N_Y_c_733_n N_A_478_65#_M1004_d 0.00563505f $X=3.64 $Y=0.927 $X2=-0.19
+ $Y2=-0.245
cc_577 N_Y_c_733_n N_A_478_65#_M1018_d 0.00399081f $X=3.64 $Y=0.927 $X2=0 $Y2=0
cc_578 N_Y_c_729_n N_A_478_65#_M1037_d 0.00279911f $X=4.265 $Y=1.15 $X2=0 $Y2=0
cc_579 N_Y_M1004_s N_A_478_65#_c_1114_n 0.00173964f $X=2.805 $Y=0.325 $X2=0
+ $Y2=0
cc_580 N_Y_c_733_n N_A_478_65#_c_1114_n 0.06617f $X=3.64 $Y=0.927 $X2=0 $Y2=0
cc_581 N_Y_M1034_s N_A_478_65#_c_1115_n 0.00176461f $X=3.665 $Y=0.325 $X2=0
+ $Y2=0
cc_582 N_Y_c_729_n N_A_478_65#_c_1115_n 0.00281168f $X=4.265 $Y=1.15 $X2=0 $Y2=0
cc_583 N_Y_c_733_n N_A_478_65#_c_1115_n 0.00378766f $X=3.64 $Y=0.927 $X2=0 $Y2=0
cc_584 N_Y_c_734_n N_A_478_65#_c_1115_n 0.0159058f $X=3.805 $Y=0.68 $X2=0 $Y2=0
cc_585 N_Y_c_729_n N_A_478_65#_c_1126_n 0.0210495f $X=4.265 $Y=1.15 $X2=0 $Y2=0
cc_586 N_VGND_c_1000_n N_A_478_65#_c_1114_n 0.0300763f $X=1.98 $Y=0.505 $X2=0
+ $Y2=0
cc_587 N_VGND_c_1005_n N_A_478_65#_c_1114_n 0.11839f $X=8.565 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_1011_n N_A_478_65#_c_1114_n 0.0657262f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_c_1005_n N_A_478_65#_c_1119_n 0.0234617f $X=8.565 $Y=0 $X2=0 $Y2=0
cc_590 N_VGND_c_1011_n N_A_478_65#_c_1119_n 0.012695f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_591 N_VGND_c_1005_n N_A_478_65#_c_1120_n 0.109255f $X=8.565 $Y=0 $X2=0 $Y2=0
cc_592 N_VGND_c_1011_n N_A_478_65#_c_1120_n 0.0605417f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_593 N_VGND_c_1011_n N_A_921_65#_c_1160_n 0.014901f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_c_1011_n N_A_921_65#_c_1173_n 0.00124588f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_595 N_VGND_c_1005_n N_A_1291_65#_c_1210_n 0.042287f $X=8.565 $Y=0 $X2=0 $Y2=0
cc_596 N_VGND_c_1011_n N_A_1291_65#_c_1210_n 0.0238254f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_597 N_VGND_c_1001_n N_A_1291_65#_c_1211_n 0.00962585f $X=8.73 $Y=0.565 $X2=0
+ $Y2=0
cc_598 N_VGND_c_1005_n N_A_1291_65#_c_1211_n 0.0558056f $X=8.565 $Y=0 $X2=0
+ $Y2=0
cc_599 N_VGND_c_1011_n N_A_1291_65#_c_1211_n 0.0311953f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_600 N_VGND_M1005_d N_A_1291_65#_c_1225_n 0.00330692f $X=8.59 $Y=0.325 $X2=0
+ $Y2=0
cc_601 N_VGND_c_1001_n N_A_1291_65#_c_1225_n 0.0167297f $X=8.73 $Y=0.565 $X2=0
+ $Y2=0
cc_602 N_VGND_c_1011_n N_A_1291_65#_c_1225_n 0.0107397f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1001_n N_A_1291_65#_c_1212_n 0.0144153f $X=8.73 $Y=0.565 $X2=0
+ $Y2=0
cc_604 N_VGND_c_1002_n N_A_1291_65#_c_1212_n 0.0144153f $X=9.59 $Y=0.565 $X2=0
+ $Y2=0
cc_605 N_VGND_c_1007_n N_A_1291_65#_c_1212_n 0.00979032f $X=9.425 $Y=0 $X2=0
+ $Y2=0
cc_606 N_VGND_c_1011_n N_A_1291_65#_c_1212_n 0.00709742f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_607 N_VGND_M1025_d N_A_1291_65#_c_1213_n 0.00330692f $X=9.45 $Y=0.325 $X2=0
+ $Y2=0
cc_608 N_VGND_c_1002_n N_A_1291_65#_c_1213_n 0.0167297f $X=9.59 $Y=0.565 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1011_n N_A_1291_65#_c_1213_n 0.0107397f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1002_n N_A_1291_65#_c_1214_n 0.0144321f $X=9.59 $Y=0.565 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1010_n N_A_1291_65#_c_1214_n 0.0134357f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1011_n N_A_1291_65#_c_1214_n 0.00974008f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_613 N_VGND_c_1005_n N_A_1291_65#_c_1215_n 0.0136191f $X=8.565 $Y=0 $X2=0
+ $Y2=0
cc_614 N_VGND_c_1011_n N_A_1291_65#_c_1215_n 0.0075906f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1005_n N_A_1291_65#_c_1216_n 0.0129313f $X=8.565 $Y=0 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1011_n N_A_1291_65#_c_1216_n 0.00720724f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_617 N_A_478_65#_c_1120_n N_A_921_65#_M1008_d 0.00176461f $X=5.07 $Y=0.45
+ $X2=-0.19 $Y2=-0.245
cc_618 N_A_478_65#_c_1117_n N_A_921_65#_M1028_d 0.00172844f $X=6.035 $Y=0.47
+ $X2=0 $Y2=0
cc_619 N_A_478_65#_M1020_s N_A_921_65#_c_1160_n 0.00332844f $X=5.035 $Y=0.325
+ $X2=0 $Y2=0
cc_620 N_A_478_65#_M1038_s N_A_921_65#_c_1160_n 0.0108086f $X=5.895 $Y=0.325
+ $X2=0 $Y2=0
cc_621 N_A_478_65#_c_1116_n N_A_921_65#_c_1160_n 0.0611031f $X=5.46 $Y=0.45
+ $X2=0 $Y2=0
cc_622 N_A_478_65#_c_1120_n N_A_921_65#_c_1160_n 0.00407346f $X=5.07 $Y=0.45
+ $X2=0 $Y2=0
cc_623 N_A_478_65#_c_1120_n N_A_921_65#_c_1166_n 0.0131301f $X=5.07 $Y=0.45
+ $X2=0 $Y2=0
cc_624 N_A_478_65#_c_1117_n N_A_1291_65#_c_1215_n 0.0195814f $X=6.035 $Y=0.47
+ $X2=0 $Y2=0
cc_625 N_A_921_65#_c_1160_n N_A_1291_65#_M1006_d 0.00561779f $X=6.845 $Y=0.92
+ $X2=-0.19 $Y2=-0.245
cc_626 N_A_921_65#_c_1173_n N_A_1291_65#_M1009_d 0.00331295f $X=7.705 $Y=0.9
+ $X2=0 $Y2=0
cc_627 N_A_921_65#_M1006_s N_A_1291_65#_c_1210_n 0.00184993f $X=6.87 $Y=0.325
+ $X2=0 $Y2=0
cc_628 N_A_921_65#_c_1160_n N_A_1291_65#_c_1210_n 0.00377044f $X=6.845 $Y=0.92
+ $X2=0 $Y2=0
cc_629 N_A_921_65#_c_1173_n N_A_1291_65#_c_1210_n 0.00371875f $X=7.705 $Y=0.9
+ $X2=0 $Y2=0
cc_630 N_A_921_65#_c_1179_n N_A_1291_65#_c_1210_n 0.0142317f $X=7.01 $Y=0.7
+ $X2=0 $Y2=0
cc_631 N_A_921_65#_M1030_s N_A_1291_65#_c_1211_n 0.00184993f $X=7.73 $Y=0.325
+ $X2=0 $Y2=0
cc_632 N_A_921_65#_c_1173_n N_A_1291_65#_c_1211_n 0.00371875f $X=7.705 $Y=0.9
+ $X2=0 $Y2=0
cc_633 N_A_921_65#_c_1184_n N_A_1291_65#_c_1211_n 0.0142317f $X=7.87 $Y=0.7
+ $X2=0 $Y2=0
cc_634 N_A_921_65#_c_1160_n N_A_1291_65#_c_1215_n 0.0143909f $X=6.845 $Y=0.92
+ $X2=0 $Y2=0
cc_635 N_A_921_65#_c_1173_n N_A_1291_65#_c_1216_n 0.0125904f $X=7.705 $Y=0.9
+ $X2=0 $Y2=0
