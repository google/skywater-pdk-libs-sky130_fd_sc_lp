* File: sky130_fd_sc_lp__nand3_lp.pxi.spice
* Created: Wed Sep  2 10:04:31 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3_LP%C N_C_M1000_g N_C_M1004_g N_C_c_45_n N_C_c_46_n C
+ C N_C_c_48_n PM_SKY130_FD_SC_LP__NAND3_LP%C
x_PM_SKY130_FD_SC_LP__NAND3_LP%B N_B_M1005_g N_B_c_74_n N_B_M1003_g N_B_c_76_n
+ N_B_c_77_n B B B N_B_c_79_n PM_SKY130_FD_SC_LP__NAND3_LP%B
x_PM_SKY130_FD_SC_LP__NAND3_LP%A N_A_M1001_g N_A_M1002_g N_A_c_124_n N_A_c_125_n
+ A N_A_c_126_n N_A_c_127_n PM_SKY130_FD_SC_LP__NAND3_LP%A
x_PM_SKY130_FD_SC_LP__NAND3_LP%VPWR N_VPWR_M1000_s N_VPWR_M1003_d N_VPWR_c_160_n
+ N_VPWR_c_161_n N_VPWR_c_162_n N_VPWR_c_163_n N_VPWR_c_164_n VPWR
+ N_VPWR_c_165_n N_VPWR_c_159_n PM_SKY130_FD_SC_LP__NAND3_LP%VPWR
x_PM_SKY130_FD_SC_LP__NAND3_LP%Y N_Y_M1001_d N_Y_M1000_d N_Y_M1002_d N_Y_c_188_n
+ N_Y_c_189_n N_Y_c_190_n N_Y_c_186_n N_Y_c_187_n N_Y_c_192_n Y Y Y
+ PM_SKY130_FD_SC_LP__NAND3_LP%Y
x_PM_SKY130_FD_SC_LP__NAND3_LP%VGND N_VGND_M1004_s N_VGND_c_232_n N_VGND_c_233_n
+ N_VGND_c_234_n VGND N_VGND_c_235_n N_VGND_c_236_n
+ PM_SKY130_FD_SC_LP__NAND3_LP%VGND
cc_1 VNB N_C_M1000_g 0.0123316f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.545
cc_2 VNB N_C_M1004_g 0.0278914f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.445
cc_3 VNB N_C_c_45_n 0.025421f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.36
cc_4 VNB N_C_c_46_n 0.016913f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.525
cc_5 VNB C 0.049118f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_C_c_48_n 0.0170897f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.02
cc_7 VNB N_B_c_74_n 0.0138849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_M1003_g 0.0142945f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.445
cc_9 VNB N_B_c_76_n 0.0167692f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.02
cc_10 VNB N_B_c_77_n 0.0238826f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.855
cc_11 VNB B 0.00202451f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.36
cc_12 VNB N_B_c_79_n 0.0167997f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.02
cc_13 VNB N_A_M1001_g 0.0274943f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.545
cc_14 VNB N_A_M1002_g 0.00914525f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.445
cc_15 VNB N_A_c_124_n 0.023974f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.36
cc_16 VNB N_A_c_125_n 0.0141141f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.525
cc_17 VNB N_A_c_126_n 0.0168121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_c_127_n 0.00789325f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.02
cc_19 VNB N_VPWR_c_159_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_186_n 0.0469445f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.02
cc_21 VNB N_Y_c_187_n 0.0279443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_232_n 0.021704f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.445
cc_23 VNB N_VGND_c_233_n 0.0123263f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.02
cc_24 VNB N_VGND_c_234_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.855
cc_25 VNB N_VGND_c_235_n 0.0502847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_236_n 0.155834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_C_M1000_g 0.0523987f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.545
cc_28 VPB N_B_M1003_g 0.0377496f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.445
cc_29 VPB N_A_M1002_g 0.0471146f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.445
cc_30 VPB N_VPWR_c_160_n 0.012566f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.445
cc_31 VPB N_VPWR_c_161_n 0.049112f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.02
cc_32 VPB N_VPWR_c_162_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_163_n 0.0220628f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.19
cc_34 VPB N_VPWR_c_164_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_165_n 0.0223858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_159_n 0.0578664f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_Y_c_188_n 0.0107084f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.855
cc_38 VPB N_Y_c_189_n 0.00824007f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.36
cc_39 VPB N_Y_c_190_n 0.0563339f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_40 VPB N_Y_c_186_n 0.00230012f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.02
cc_41 VPB N_Y_c_192_n 0.0163622f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.19
cc_42 VPB Y 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 N_C_c_46_n N_B_c_74_n 0.0175101f $X=0.61 $Y=1.525 $X2=0 $Y2=0
cc_44 N_C_c_46_n N_B_M1003_g 0.0355188f $X=0.61 $Y=1.525 $X2=0 $Y2=0
cc_45 C N_B_M1003_g 0.00233426f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_46 N_C_M1004_g N_B_c_76_n 0.0175101f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_47 N_C_c_45_n N_B_c_77_n 0.0175101f $X=0.61 $Y=1.36 $X2=0 $Y2=0
cc_48 N_C_M1004_g B 0.00198258f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_49 C B 0.0468687f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_50 N_C_c_48_n B 6.51932e-19 $X=0.61 $Y=1.02 $X2=0 $Y2=0
cc_51 C N_B_c_79_n 0.00379022f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_52 N_C_c_48_n N_B_c_79_n 0.0175101f $X=0.61 $Y=1.02 $X2=0 $Y2=0
cc_53 N_C_M1000_g N_VPWR_c_161_n 0.00758316f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_54 C N_VPWR_c_161_n 0.0109253f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_55 N_C_M1000_g N_VPWR_c_162_n 9.30781e-19 $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_56 N_C_M1000_g N_VPWR_c_163_n 0.00658484f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_57 N_C_M1000_g N_VPWR_c_159_n 0.0111188f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_58 N_C_M1000_g N_Y_c_189_n 0.014769f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_59 C N_Y_c_189_n 0.019027f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_60 N_C_M1000_g Y 0.0364935f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_61 N_C_M1004_g N_VGND_c_232_n 0.0142538f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_62 C N_VGND_c_232_n 0.0275544f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_63 N_C_c_48_n N_VGND_c_232_n 0.0048437f $X=0.61 $Y=1.02 $X2=0 $Y2=0
cc_64 N_C_M1004_g N_VGND_c_235_n 0.00486043f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_65 N_C_M1004_g N_VGND_c_236_n 0.00456945f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_66 C N_VGND_c_236_n 0.014985f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B_c_76_n N_A_M1001_g 0.017898f $X=1.18 $Y=0.765 $X2=0 $Y2=0
cc_68 B N_A_M1001_g 0.00466138f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_69 N_B_c_79_n N_A_M1001_g 0.0119135f $X=1.18 $Y=0.93 $X2=0 $Y2=0
cc_70 N_B_c_74_n N_A_c_124_n 0.0119135f $X=1.18 $Y=1.435 $X2=0 $Y2=0
cc_71 N_B_M1003_g N_A_c_125_n 0.0350619f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_72 N_B_c_77_n N_A_c_126_n 0.0119135f $X=1.18 $Y=1.27 $X2=0 $Y2=0
cc_73 B N_A_c_126_n 7.12343e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_74 N_B_M1003_g N_A_c_127_n 0.00195423f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_75 B N_A_c_127_n 0.0379791f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_76 N_B_c_79_n N_A_c_127_n 0.00355018f $X=1.18 $Y=0.93 $X2=0 $Y2=0
cc_77 N_B_M1003_g N_VPWR_c_162_n 0.0217134f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_78 N_B_M1003_g N_VPWR_c_163_n 0.00769046f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_79 N_B_M1003_g N_VPWR_c_159_n 0.0134474f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_80 N_B_c_74_n N_Y_c_188_n 2.46944e-19 $X=1.18 $Y=1.435 $X2=0 $Y2=0
cc_81 N_B_M1003_g N_Y_c_188_n 0.018626f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_82 B N_Y_c_188_n 0.0139985f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_83 N_B_c_74_n N_Y_c_189_n 2.89032e-19 $X=1.18 $Y=1.435 $X2=0 $Y2=0
cc_84 N_B_M1003_g N_Y_c_189_n 0.00286413f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_85 B N_Y_c_189_n 0.00391311f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_86 N_B_M1003_g N_Y_c_190_n 0.00101079f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_87 N_B_c_76_n N_Y_c_187_n 0.0010022f $X=1.18 $Y=0.765 $X2=0 $Y2=0
cc_88 B N_Y_c_187_n 0.0104887f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_89 N_B_M1003_g Y 0.0233221f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_90 N_B_c_76_n N_VGND_c_232_n 0.00272611f $X=1.18 $Y=0.765 $X2=0 $Y2=0
cc_91 B N_VGND_c_232_n 0.00954636f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_92 N_B_c_76_n N_VGND_c_235_n 0.00394642f $X=1.18 $Y=0.765 $X2=0 $Y2=0
cc_93 B N_VGND_c_235_n 0.00930091f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_94 N_B_c_79_n N_VGND_c_235_n 4.68308e-19 $X=1.18 $Y=0.93 $X2=0 $Y2=0
cc_95 N_B_c_76_n N_VGND_c_236_n 0.00586352f $X=1.18 $Y=0.765 $X2=0 $Y2=0
cc_96 B N_VGND_c_236_n 0.0106938f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_97 B A_233_47# 0.00428579f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_98 N_A_M1002_g N_VPWR_c_162_n 0.0229651f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_99 N_A_M1002_g N_VPWR_c_165_n 0.00769046f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_100 N_A_M1002_g N_VPWR_c_159_n 0.0141575f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_101 N_A_M1002_g N_Y_c_188_n 0.0178513f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_102 N_A_c_127_n N_Y_c_188_n 0.0178533f $X=1.75 $Y=1.02 $X2=0 $Y2=0
cc_103 N_A_M1002_g N_Y_c_190_n 0.0251588f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_104 N_A_M1001_g N_Y_c_186_n 0.00362326f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_M1002_g N_Y_c_186_n 0.00427061f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_106 N_A_c_126_n N_Y_c_186_n 0.0148853f $X=1.75 $Y=1.02 $X2=0 $Y2=0
cc_107 N_A_c_127_n N_Y_c_186_n 0.0483772f $X=1.75 $Y=1.02 $X2=0 $Y2=0
cc_108 N_A_M1001_g N_Y_c_187_n 0.00830224f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_c_126_n N_Y_c_187_n 0.0013229f $X=1.75 $Y=1.02 $X2=0 $Y2=0
cc_110 N_A_c_127_n N_Y_c_187_n 0.0161733f $X=1.75 $Y=1.02 $X2=0 $Y2=0
cc_111 N_A_M1002_g N_Y_c_192_n 0.00448409f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_112 N_A_c_125_n N_Y_c_192_n 6.14058e-19 $X=1.75 $Y=1.525 $X2=0 $Y2=0
cc_113 N_A_c_127_n N_Y_c_192_n 0.00875454f $X=1.75 $Y=1.02 $X2=0 $Y2=0
cc_114 N_A_M1002_g Y 0.00101008f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_115 N_A_M1001_g N_VGND_c_235_n 0.0054778f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_M1001_g N_VGND_c_236_n 0.00791832f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_c_127_n N_VGND_c_236_n 0.00494663f $X=1.75 $Y=1.02 $X2=0 $Y2=0
cc_118 N_VPWR_c_162_n N_Y_c_188_n 0.0207154f $X=1.445 $Y=2.22 $X2=0 $Y2=0
cc_119 N_VPWR_c_162_n N_Y_c_190_n 0.0682253f $X=1.445 $Y=2.22 $X2=0 $Y2=0
cc_120 N_VPWR_c_165_n N_Y_c_190_n 0.0304602f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_121 N_VPWR_c_159_n N_Y_c_190_n 0.0174175f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_122 N_VPWR_c_161_n Y 0.0778156f $X=0.34 $Y=2.19 $X2=0 $Y2=0
cc_123 N_VPWR_c_162_n Y 0.0684559f $X=1.445 $Y=2.22 $X2=0 $Y2=0
cc_124 N_VPWR_c_163_n Y 0.0312234f $X=1.28 $Y=3.33 $X2=0 $Y2=0
cc_125 N_VPWR_c_159_n Y 0.0174129f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_126 N_Y_c_187_n N_VGND_c_235_n 0.0252817f $X=1.875 $Y=0.47 $X2=0 $Y2=0
cc_127 N_Y_M1001_d N_VGND_c_236_n 0.0023218f $X=1.735 $Y=0.235 $X2=0 $Y2=0
cc_128 N_Y_c_187_n N_VGND_c_236_n 0.0198916f $X=1.875 $Y=0.47 $X2=0 $Y2=0
cc_129 N_VGND_c_236_n A_155_47# 0.00860318f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
cc_130 N_VGND_c_236_n A_233_47# 0.0114018f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
