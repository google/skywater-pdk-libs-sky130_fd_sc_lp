* File: sky130_fd_sc_lp__or3_m.pxi.spice
* Created: Wed Sep  2 10:30:56 2020
* 
x_PM_SKY130_FD_SC_LP__OR3_M%C N_C_M1002_g N_C_c_62_n N_C_c_63_n N_C_c_69_n
+ N_C_c_70_n N_C_M1005_g N_C_c_64_n C C C N_C_c_66_n N_C_c_67_n
+ PM_SKY130_FD_SC_LP__OR3_M%C
x_PM_SKY130_FD_SC_LP__OR3_M%B N_B_M1001_g N_B_M1007_g N_B_c_106_n N_B_c_107_n
+ N_B_c_108_n B B N_B_c_110_n PM_SKY130_FD_SC_LP__OR3_M%B
x_PM_SKY130_FD_SC_LP__OR3_M%A N_A_M1006_g N_A_M1004_g N_A_c_150_n N_A_c_151_n A
+ N_A_c_152_n N_A_c_153_n PM_SKY130_FD_SC_LP__OR3_M%A
x_PM_SKY130_FD_SC_LP__OR3_M%A_43_47# N_A_43_47#_M1002_s N_A_43_47#_M1001_d
+ N_A_43_47#_M1005_s N_A_43_47#_c_198_n N_A_43_47#_M1003_g N_A_43_47#_M1000_g
+ N_A_43_47#_c_193_n N_A_43_47#_c_201_n N_A_43_47#_c_202_n N_A_43_47#_c_203_n
+ N_A_43_47#_c_204_n N_A_43_47#_c_205_n N_A_43_47#_c_194_n N_A_43_47#_c_206_n
+ N_A_43_47#_c_195_n N_A_43_47#_c_196_n N_A_43_47#_c_197_n N_A_43_47#_c_219_n
+ N_A_43_47#_c_208_n N_A_43_47#_c_209_n PM_SKY130_FD_SC_LP__OR3_M%A_43_47#
x_PM_SKY130_FD_SC_LP__OR3_M%VPWR N_VPWR_M1006_d N_VPWR_c_289_n N_VPWR_c_290_n
+ N_VPWR_c_291_n VPWR N_VPWR_c_292_n N_VPWR_c_288_n
+ PM_SKY130_FD_SC_LP__OR3_M%VPWR
x_PM_SKY130_FD_SC_LP__OR3_M%X N_X_M1003_d N_X_M1000_d X X X X X X X X X
+ N_X_c_315_n PM_SKY130_FD_SC_LP__OR3_M%X
x_PM_SKY130_FD_SC_LP__OR3_M%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_c_334_n
+ N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n VGND N_VGND_c_338_n
+ N_VGND_c_339_n N_VGND_c_340_n N_VGND_c_341_n PM_SKY130_FD_SC_LP__OR3_M%VGND
cc_1 VNB N_C_c_62_n 0.0234759f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.248
cc_2 VNB N_C_c_63_n 0.0105712f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.675
cc_3 VNB N_C_c_64_n 0.0177363f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.435
cc_4 VNB C 0.00285959f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB N_C_c_66_n 0.0217807f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.93
cc_6 VNB N_C_c_67_n 0.0213139f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=0.765
cc_7 VNB N_B_M1007_g 0.016371f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.435
cc_8 VNB N_B_c_106_n 0.0188694f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.75
cc_9 VNB N_B_c_107_n 0.0187137f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.825
cc_10 VNB N_B_c_108_n 0.0182204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB B 0.00403377f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.435
cc_12 VNB N_B_c_110_n 0.0260289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_M1004_g 0.0279611f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.675
cc_14 VNB N_A_c_150_n 0.0189756f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.195
cc_15 VNB N_A_c_151_n 0.00950329f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.195
cc_16 VNB N_A_c_152_n 0.0150415f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_17 VNB N_A_c_153_n 0.00842727f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_18 VNB N_A_43_47#_M1003_g 0.0645913f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.435
cc_19 VNB N_A_43_47#_c_193_n 0.0482227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_43_47#_c_194_n 0.00136178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_43_47#_c_195_n 0.0108561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_43_47#_c_196_n 0.00615618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_43_47#_c_197_n 0.00562888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_288_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.93
cc_25 VNB X 0.0101162f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.675
cc_26 VNB X 0.0543694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_334_n 0.0027661f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.75
cc_28 VNB N_VGND_c_335_n 0.00433998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_336_n 0.0153555f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_30 VNB N_VGND_c_337_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_31 VNB N_VGND_c_338_n 0.030783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_339_n 0.0220412f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.295
cc_33 VNB N_VGND_c_340_n 0.176337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_341_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_C_c_63_n 7.76949e-19 $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.675
cc_36 VPB N_C_c_69_n 0.032637f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.75
cc_37 VPB N_C_c_70_n 0.0104381f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.75
cc_38 VPB N_C_M1005_g 0.0252423f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.195
cc_39 VPB N_B_M1007_g 0.0217819f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.435
cc_40 VPB N_A_M1006_g 0.0254213f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.445
cc_41 VPB N_A_c_151_n 0.00527662f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.195
cc_42 VPB N_A_43_47#_c_198_n 0.0529065f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=1.825
cc_43 VPB N_A_43_47#_M1003_g 0.0429591f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.435
cc_44 VPB N_A_43_47#_c_193_n 0.00644978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_43_47#_c_201_n 0.0107183f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.93
cc_46 VPB N_A_43_47#_c_202_n 0.0149891f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.93
cc_47 VPB N_A_43_47#_c_203_n 7.87255e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_43_47#_c_204_n 0.0102925f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.925
cc_49 VPB N_A_43_47#_c_205_n 0.0117398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_43_47#_c_206_n 0.0139038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_43_47#_c_197_n 0.00155037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_43_47#_c_208_n 0.00661647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_43_47#_c_209_n 0.0513783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_289_n 0.020532f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.435
cc_55 VPB N_VPWR_c_290_n 0.056758f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.75
cc_56 VPB N_VPWR_c_291_n 0.00632158f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=1.825
cc_57 VPB N_VPWR_c_292_n 0.023333f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=0.93
cc_58 VPB N_VPWR_c_288_n 0.102204f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.93
cc_59 VPB X 0.0222134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB X 0.026731f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_X_c_315_n 0.00874805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 N_C_c_63_n N_B_M1007_g 0.00137928f $X=0.555 $Y=1.675 $X2=0 $Y2=0
cc_63 N_C_c_69_n N_B_M1007_g 0.0526703f $X=0.93 $Y=1.75 $X2=0 $Y2=0
cc_64 C N_B_c_106_n 0.00437248f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_65 N_C_c_67_n N_B_c_106_n 0.00584737f $X=0.667 $Y=0.765 $X2=0 $Y2=0
cc_66 C N_B_c_107_n 0.00226188f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_67 N_C_c_66_n N_B_c_107_n 0.0140104f $X=0.69 $Y=0.93 $X2=0 $Y2=0
cc_68 N_C_c_69_n N_B_c_108_n 0.00101013f $X=0.93 $Y=1.75 $X2=0 $Y2=0
cc_69 N_C_c_64_n N_B_c_108_n 0.0140104f $X=0.667 $Y=1.435 $X2=0 $Y2=0
cc_70 C B 0.0287056f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_71 N_C_c_66_n B 0.00229005f $X=0.69 $Y=0.93 $X2=0 $Y2=0
cc_72 N_C_c_62_n N_B_c_110_n 0.0140104f $X=0.667 $Y=1.248 $X2=0 $Y2=0
cc_73 C N_A_43_47#_c_193_n 0.0605595f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_74 N_C_c_67_n N_A_43_47#_c_193_n 0.0366174f $X=0.667 $Y=0.765 $X2=0 $Y2=0
cc_75 N_C_c_69_n N_A_43_47#_c_201_n 0.00168051f $X=0.93 $Y=1.75 $X2=0 $Y2=0
cc_76 N_C_c_70_n N_A_43_47#_c_201_n 0.00960287f $X=0.63 $Y=1.75 $X2=0 $Y2=0
cc_77 C N_A_43_47#_c_201_n 0.00324953f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_78 N_C_M1005_g N_A_43_47#_c_203_n 5.07566e-19 $X=1.005 $Y=2.195 $X2=0 $Y2=0
cc_79 N_C_c_69_n N_A_43_47#_c_204_n 0.00793547f $X=0.93 $Y=1.75 $X2=0 $Y2=0
cc_80 N_C_M1005_g N_A_43_47#_c_204_n 0.0128061f $X=1.005 $Y=2.195 $X2=0 $Y2=0
cc_81 N_C_M1005_g N_A_43_47#_c_205_n 0.00272023f $X=1.005 $Y=2.195 $X2=0 $Y2=0
cc_82 N_C_c_69_n N_A_43_47#_c_219_n 0.00912276f $X=0.93 $Y=1.75 $X2=0 $Y2=0
cc_83 N_C_c_64_n N_A_43_47#_c_219_n 4.22351e-19 $X=0.667 $Y=1.435 $X2=0 $Y2=0
cc_84 C N_A_43_47#_c_219_n 0.00536356f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_85 N_C_M1005_g N_VPWR_c_288_n 0.00393927f $X=1.005 $Y=2.195 $X2=0 $Y2=0
cc_86 C N_VGND_M1002_d 0.00448587f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_87 C N_VGND_c_334_n 0.00111151f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_88 N_C_c_67_n N_VGND_c_334_n 0.00544326f $X=0.667 $Y=0.765 $X2=0 $Y2=0
cc_89 C N_VGND_c_338_n 0.0049248f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_90 N_C_c_66_n N_VGND_c_338_n 0.00146872f $X=0.69 $Y=0.93 $X2=0 $Y2=0
cc_91 N_C_c_67_n N_VGND_c_338_n 0.00555499f $X=0.667 $Y=0.765 $X2=0 $Y2=0
cc_92 C N_VGND_c_340_n 0.00664343f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_93 N_C_c_66_n N_VGND_c_340_n 0.00134702f $X=0.69 $Y=0.93 $X2=0 $Y2=0
cc_94 N_C_c_67_n N_VGND_c_340_n 0.011951f $X=0.667 $Y=0.765 $X2=0 $Y2=0
cc_95 N_B_c_106_n N_A_M1004_g 0.0204633f $X=1.252 $Y=0.765 $X2=0 $Y2=0
cc_96 B N_A_M1004_g 6.10683e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_97 N_B_c_110_n N_A_M1004_g 0.00328357f $X=1.23 $Y=0.93 $X2=0 $Y2=0
cc_98 N_B_c_108_n N_A_c_150_n 0.0382316f $X=1.252 $Y=1.435 $X2=0 $Y2=0
cc_99 N_B_M1007_g N_A_c_151_n 0.0382316f $X=1.365 $Y=2.195 $X2=0 $Y2=0
cc_100 B N_A_c_152_n 8.38169e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_101 N_B_c_110_n N_A_c_152_n 0.0147262f $X=1.23 $Y=0.93 $X2=0 $Y2=0
cc_102 N_B_c_108_n N_A_c_153_n 0.00470309f $X=1.252 $Y=1.435 $X2=0 $Y2=0
cc_103 B N_A_c_153_n 0.0192112f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_104 N_B_c_110_n N_A_c_153_n 0.00154322f $X=1.23 $Y=0.93 $X2=0 $Y2=0
cc_105 N_B_M1007_g N_A_43_47#_c_204_n 0.00156812f $X=1.365 $Y=2.195 $X2=0 $Y2=0
cc_106 N_B_c_108_n N_A_43_47#_c_204_n 0.002331f $X=1.252 $Y=1.435 $X2=0 $Y2=0
cc_107 B N_A_43_47#_c_204_n 0.00808774f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_108 N_B_M1007_g N_A_43_47#_c_205_n 0.0190742f $X=1.365 $Y=2.195 $X2=0 $Y2=0
cc_109 N_B_c_106_n N_A_43_47#_c_194_n 0.001666f $X=1.252 $Y=0.765 $X2=0 $Y2=0
cc_110 N_B_c_106_n N_A_43_47#_c_196_n 0.00246608f $X=1.252 $Y=0.765 $X2=0 $Y2=0
cc_111 B N_A_43_47#_c_196_n 0.0101535f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_112 N_B_M1007_g N_A_43_47#_c_208_n 0.0106648f $X=1.365 $Y=2.195 $X2=0 $Y2=0
cc_113 B N_A_43_47#_c_208_n 8.75347e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_114 N_B_M1007_g N_A_43_47#_c_209_n 0.00802091f $X=1.365 $Y=2.195 $X2=0 $Y2=0
cc_115 N_B_c_106_n N_VGND_c_334_n 0.00825083f $X=1.252 $Y=0.765 $X2=0 $Y2=0
cc_116 N_B_c_107_n N_VGND_c_334_n 0.00315899f $X=1.252 $Y=0.915 $X2=0 $Y2=0
cc_117 B N_VGND_c_334_n 0.00871739f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_118 N_B_c_106_n N_VGND_c_336_n 0.00486043f $X=1.252 $Y=0.765 $X2=0 $Y2=0
cc_119 N_B_c_106_n N_VGND_c_340_n 0.00838234f $X=1.252 $Y=0.765 $X2=0 $Y2=0
cc_120 B N_VGND_c_340_n 9.30845e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_121 N_A_M1006_g N_A_43_47#_c_198_n 0.00971367f $X=1.725 $Y=2.195 $X2=0 $Y2=0
cc_122 N_A_M1006_g N_A_43_47#_M1003_g 0.0183501f $X=1.725 $Y=2.195 $X2=0 $Y2=0
cc_123 N_A_M1004_g N_A_43_47#_M1003_g 0.0210898f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A_c_152_n N_A_43_47#_M1003_g 0.0428645f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_c_153_n N_A_43_47#_M1003_g 6.05484e-19 $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_M1006_g N_A_43_47#_c_205_n 0.00287053f $X=1.725 $Y=2.195 $X2=0 $Y2=0
cc_127 N_A_M1004_g N_A_43_47#_c_194_n 0.00170909f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_128 N_A_M1006_g N_A_43_47#_c_206_n 0.0150385f $X=1.725 $Y=2.195 $X2=0 $Y2=0
cc_129 N_A_c_151_n N_A_43_47#_c_206_n 0.00501678f $X=1.815 $Y=1.665 $X2=0 $Y2=0
cc_130 N_A_c_153_n N_A_43_47#_c_206_n 0.0230466f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_M1004_g N_A_43_47#_c_195_n 0.0119958f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A_c_152_n N_A_43_47#_c_195_n 0.00411815f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_c_153_n N_A_43_47#_c_195_n 0.0213608f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_c_152_n N_A_43_47#_c_196_n 0.00103578f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_153_n N_A_43_47#_c_196_n 0.00761077f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_M1006_g N_A_43_47#_c_197_n 0.00223388f $X=1.725 $Y=2.195 $X2=0 $Y2=0
cc_137 N_A_M1004_g N_A_43_47#_c_197_n 0.00180664f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_138 N_A_c_151_n N_A_43_47#_c_197_n 0.00163398f $X=1.815 $Y=1.665 $X2=0 $Y2=0
cc_139 N_A_c_152_n N_A_43_47#_c_197_n 0.00313912f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_c_153_n N_A_43_47#_c_197_n 0.0371013f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_c_153_n N_A_43_47#_c_208_n 0.00236015f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_M1006_g N_VPWR_c_289_n 0.00129574f $X=1.725 $Y=2.195 $X2=0 $Y2=0
cc_143 N_A_M1004_g N_VGND_c_334_n 7.58747e-19 $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A_M1004_g N_VGND_c_335_n 0.0015506f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_145 N_A_M1004_g N_VGND_c_336_n 0.00437852f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_M1004_g N_VGND_c_340_n 0.00614167f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_43_47#_c_198_n N_VPWR_c_289_n 0.0258133f $X=2.19 $Y=2.85 $X2=0 $Y2=0
cc_148 N_A_43_47#_M1003_g N_VPWR_c_289_n 0.00796314f $X=2.265 $Y=0.445 $X2=0
+ $Y2=0
cc_149 N_A_43_47#_c_205_n N_VPWR_c_289_n 0.0478384f $X=1.46 $Y=2.94 $X2=0 $Y2=0
cc_150 N_A_43_47#_c_206_n N_VPWR_c_289_n 0.0228627f $X=2.16 $Y=1.88 $X2=0 $Y2=0
cc_151 N_A_43_47#_c_209_n N_VPWR_c_289_n 0.00524695f $X=1.46 $Y=2.85 $X2=0 $Y2=0
cc_152 N_A_43_47#_c_198_n N_VPWR_c_290_n 0.00445258f $X=2.19 $Y=2.85 $X2=0 $Y2=0
cc_153 N_A_43_47#_c_205_n N_VPWR_c_290_n 0.0167839f $X=1.46 $Y=2.94 $X2=0 $Y2=0
cc_154 N_A_43_47#_c_209_n N_VPWR_c_290_n 0.0059602f $X=1.46 $Y=2.85 $X2=0 $Y2=0
cc_155 N_A_43_47#_c_198_n N_VPWR_c_292_n 0.00581074f $X=2.19 $Y=2.85 $X2=0 $Y2=0
cc_156 N_A_43_47#_c_198_n N_VPWR_c_288_n 0.0111595f $X=2.19 $Y=2.85 $X2=0 $Y2=0
cc_157 N_A_43_47#_c_205_n N_VPWR_c_288_n 0.0108843f $X=1.46 $Y=2.94 $X2=0 $Y2=0
cc_158 N_A_43_47#_c_209_n N_VPWR_c_288_n 0.00813556f $X=1.46 $Y=2.85 $X2=0 $Y2=0
cc_159 N_A_43_47#_M1003_g X 0.0031553f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_43_47#_c_195_n X 8.02648e-19 $X=2.16 $Y=0.81 $X2=0 $Y2=0
cc_161 N_A_43_47#_M1003_g X 0.033579f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_43_47#_c_206_n X 0.0109915f $X=2.16 $Y=1.88 $X2=0 $Y2=0
cc_163 N_A_43_47#_c_195_n X 0.0109915f $X=2.16 $Y=0.81 $X2=0 $Y2=0
cc_164 N_A_43_47#_c_197_n X 0.0521626f $X=2.245 $Y=1.795 $X2=0 $Y2=0
cc_165 N_A_43_47#_c_198_n X 0.00352547f $X=2.19 $Y=2.85 $X2=0 $Y2=0
cc_166 N_A_43_47#_M1003_g X 0.012309f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A_43_47#_M1003_g N_X_c_315_n 0.00283907f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_43_47#_c_206_n N_X_c_315_n 0.00108594f $X=2.16 $Y=1.88 $X2=0 $Y2=0
cc_169 N_A_43_47#_M1003_g N_VGND_c_335_n 0.00452264f $X=2.265 $Y=0.445 $X2=0
+ $Y2=0
cc_170 N_A_43_47#_c_195_n N_VGND_c_335_n 0.0148498f $X=2.16 $Y=0.81 $X2=0 $Y2=0
cc_171 N_A_43_47#_c_194_n N_VGND_c_336_n 0.00776392f $X=1.58 $Y=0.51 $X2=0 $Y2=0
cc_172 N_A_43_47#_c_195_n N_VGND_c_336_n 0.00305343f $X=2.16 $Y=0.81 $X2=0 $Y2=0
cc_173 N_A_43_47#_c_193_n N_VGND_c_338_n 0.00831216f $X=0.34 $Y=0.51 $X2=0 $Y2=0
cc_174 N_A_43_47#_M1003_g N_VGND_c_339_n 0.00425102f $X=2.265 $Y=0.445 $X2=0
+ $Y2=0
cc_175 N_A_43_47#_c_195_n N_VGND_c_339_n 0.00301865f $X=2.16 $Y=0.81 $X2=0 $Y2=0
cc_176 N_A_43_47#_M1002_s N_VGND_c_340_n 0.00489501f $X=0.215 $Y=0.235 $X2=0
+ $Y2=0
cc_177 N_A_43_47#_M1001_d N_VGND_c_340_n 0.00442034f $X=1.44 $Y=0.235 $X2=0
+ $Y2=0
cc_178 N_A_43_47#_M1003_g N_VGND_c_340_n 0.00705503f $X=2.265 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_A_43_47#_c_193_n N_VGND_c_340_n 0.0069578f $X=0.34 $Y=0.51 $X2=0 $Y2=0
cc_180 N_A_43_47#_c_194_n N_VGND_c_340_n 0.00690901f $X=1.58 $Y=0.51 $X2=0 $Y2=0
cc_181 N_A_43_47#_c_195_n N_VGND_c_340_n 0.0108681f $X=2.16 $Y=0.81 $X2=0 $Y2=0
cc_182 N_VPWR_c_292_n X 0.0121896f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_288_n X 0.0139254f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_289_n N_X_c_315_n 0.0438388f $X=1.97 $Y=2.26 $X2=0 $Y2=0
cc_185 X N_VGND_c_335_n 0.0140547f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_186 X N_VGND_c_335_n 0.00219104f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_187 X N_VGND_c_339_n 0.0219946f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_188 N_X_M1003_d N_VGND_c_340_n 0.00215867f $X=2.34 $Y=0.235 $X2=0 $Y2=0
cc_189 X N_VGND_c_340_n 0.0151186f $X=2.555 $Y=0.47 $X2=0 $Y2=0
