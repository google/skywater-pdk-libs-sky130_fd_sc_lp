* File: sky130_fd_sc_lp__ebufn_4.spice
* Created: Fri Aug 28 10:31:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ebufn_4.pex.spice"
.subckt sky130_fd_sc_lp__ebufn_4  VNB VPB TE_B A Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1000 N_Z_M1000_d N_A_84_21#_M1000_g N_A_27_47#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1003 N_Z_M1000_d N_A_84_21#_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.6
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1004 N_Z_M1004_d N_A_84_21#_M1004_g N_A_27_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1018 N_Z_M1004_d N_A_84_21#_M1018_g N_A_27_47#_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A_456_21#_M1008_g N_A_27_47#_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1008_d N_A_456_21#_M1010_g N_A_27_47#_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_456_21#_M1013_g N_A_27_47#_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1013_d N_A_456_21#_M1014_g N_A_27_47#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75003.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_TE_B_M1012_g N_A_456_21#_M1012_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1764 AS=0.2394 PD=1.26 PS=2.25 NRD=9.996 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1019 N_A_84_21#_M1019_d N_A_M1019_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1764 PD=2.25 PS=1.26 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_Z_M1001_d N_A_84_21#_M1001_g N_A_27_367#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1006 N_Z_M1001_d N_A_84_21#_M1006_g N_A_27_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2205 PD=1.54 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1011 N_Z_M1011_d N_A_84_21#_M1011_g N_A_27_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75002.8 A=0.189 P=2.82 MULT=1
MM1015 N_Z_M1011_d N_A_84_21#_M1015_g N_A_27_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75001.6 SB=75002.3 A=0.189 P=2.82 MULT=1
MM1007 N_A_27_367#_M1015_s N_TE_B_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2646 PD=1.61 PS=1.68 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75002.1 SB=75001.8 A=0.189 P=2.82 MULT=1
MM1009 N_A_27_367#_M1009_d N_TE_B_M1009_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2646 PD=1.54 PS=1.68 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75002.7 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1016 N_A_27_367#_M1009_d N_TE_B_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2898 PD=1.54 PS=1.72 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75003.1 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1017 N_A_27_367#_M1017_d N_TE_B_M1017_g N_VPWR_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.2898 PD=3.09 PS=1.72 NRD=0 NRS=17.1981 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_TE_B_M1002_g N_A_456_21#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.5185 PD=1.61 PS=3.42 NRD=0 NRS=17.9664 M=1 R=8.4
+ SA=75000.3 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1005 N_A_84_21#_M1005_d N_A_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.2205 PD=3.09 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4 SA=75000.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3883 P=17.07
c_75 VNB 0 2.71838e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__ebufn_4.pxi.spice"
*
.ends
*
*
