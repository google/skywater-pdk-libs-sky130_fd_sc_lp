* File: sky130_fd_sc_lp__or2b_lp.pex.spice
* Created: Wed Sep  2 10:30:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2B_LP%B_N 3 7 11 15 17 18 19 23
r37 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=1.295
+ $X2=0.725 $Y2=1.665
r38 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=1.34 $X2=0.725 $Y2=1.34
r39 16 23 33.9804 $w=4.55e-07 $l=2.78e-07 $layer=POLY_cond $X=0.662 $Y=1.618
+ $X2=0.662 $Y2=1.34
r40 16 17 38.953 $w=4.55e-07 $l=2.27e-07 $layer=POLY_cond $X=0.662 $Y=1.618
+ $X2=0.662 $Y2=1.845
r41 15 23 1.83347 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=0.662 $Y=1.325
+ $X2=0.662 $Y2=1.34
r42 7 17 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.56 $Y=2.545 $X2=0.56
+ $Y2=1.845
r43 1 15 24.7927 $w=4.55e-07 $l=1.5e-07 $layer=POLY_cond $X=0.69 $Y=1.175
+ $X2=0.69 $Y2=1.325
r44 1 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.87 $Y=1.175
+ $X2=0.87 $Y2=0.495
r45 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.51 $Y=1.175 $X2=0.51
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_LP%A_30_57# 1 2 7 9 10 12 15 19 23 27 31 33 37
c65 33 0 5.81057e-20 $X=1.35 $Y=0.99
r66 34 37 31.0968 $w=5.27e-07 $l=3.4e-07 $layer=POLY_cond $X=1.35 $Y=1.16
+ $X2=1.69 $Y2=1.16
r67 34 35 4.57305 $w=5.27e-07 $l=5e-08 $layer=POLY_cond $X=1.35 $Y=1.16 $X2=1.3
+ $Y2=1.16
r68 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=0.99 $X2=1.35 $Y2=0.99
r69 28 31 3.3199 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=0.91
+ $X2=0.295 $Y2=0.91
r70 27 33 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=0.91
+ $X2=1.35 $Y2=0.91
r71 27 28 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.185 $Y=0.91
+ $X2=0.46 $Y2=0.91
r72 23 25 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.255 $Y=2.19
+ $X2=0.255 $Y2=2.9
r73 21 31 3.24686 $w=2.9e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.255 $Y=0.995
+ $X2=0.295 $Y2=0.91
r74 21 23 55.0868 $w=2.48e-07 $l=1.195e-06 $layer=LI1_cond $X=0.255 $Y=0.995
+ $X2=0.255 $Y2=2.19
r75 17 31 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.295 $Y=0.825
+ $X2=0.295 $Y2=0.91
r76 17 19 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.295 $Y=0.825
+ $X2=0.295 $Y2=0.495
r77 13 37 15.5484 $w=5.27e-07 $l=4.11309e-07 $layer=POLY_cond $X=1.86 $Y=1.495
+ $X2=1.69 $Y2=1.16
r78 13 15 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.86 $Y=1.495
+ $X2=1.86 $Y2=2.545
r79 10 37 32.7418 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.69 $Y=0.825
+ $X2=1.69 $Y2=1.16
r80 10 12 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.69 $Y=0.825
+ $X2=1.69 $Y2=0.495
r81 7 35 32.7418 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.3 $Y=0.825 $X2=1.3
+ $Y2=1.16
r82 7 9 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.3 $Y=0.825 $X2=1.3
+ $Y2=0.495
r83 2 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.045 $X2=0.295 $Y2=2.9
r84 2 23 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.045 $X2=0.295 $Y2=2.19
r85 1 19 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.285 $X2=0.295 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_LP%A 1 3 4 5 8 10 12 16 17 18 19 20 21 22 23 29
+ 30
c64 5 0 5.81057e-20 $X=2.195 $Y=0.855
r65 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.39
+ $Y=1.38 $X2=2.39 $Y2=1.38
r66 22 23 8.67743 $w=5.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.3 $Y=2.405 $X2=2.3
+ $Y2=2.775
r67 21 22 8.67743 $w=5.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.3 $Y=2.035 $X2=2.3
+ $Y2=2.405
r68 20 21 8.67743 $w=5.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.3 $Y=1.665 $X2=2.3
+ $Y2=2.035
r69 20 30 6.68397 $w=5.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.3 $Y=1.665
+ $X2=2.3 $Y2=1.38
r70 17 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.39 $Y=1.72
+ $X2=2.39 $Y2=1.38
r71 17 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.39 $Y=1.72
+ $X2=2.39 $Y2=1.885
r72 16 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.39 $Y=1.215
+ $X2=2.39 $Y2=1.38
r73 13 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.48 $Y=0.93
+ $X2=2.48 $Y2=0.855
r74 13 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.48 $Y=0.93
+ $X2=2.48 $Y2=1.215
r75 10 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.48 $Y=0.78
+ $X2=2.48 $Y2=0.855
r76 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.48 $Y=0.78 $X2=2.48
+ $Y2=0.495
r77 8 18 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.35 $Y=2.545
+ $X2=2.35 $Y2=1.885
r78 4 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.405 $Y=0.855
+ $X2=2.48 $Y2=0.855
r79 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.405 $Y=0.855
+ $X2=2.195 $Y2=0.855
r80 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=0.78
+ $X2=2.195 $Y2=0.855
r81 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.12 $Y=0.78 $X2=2.12
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_LP%A_290_409# 1 2 9 13 17 23 25 28 32 36 41 42
+ 43 45 46
r86 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3 $Y=1.03
+ $X2=3 $Y2=1.03
r87 41 42 8.80985 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=1.647 $Y=2.19
+ $X2=1.647 $Y2=2.025
r88 37 43 3.08518 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=2.07 $Y=0.95
+ $X2=1.882 $Y2=0.95
r89 36 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=0.95 $X2=3
+ $Y2=0.95
r90 36 37 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.835 $Y=0.95
+ $X2=2.07 $Y2=0.95
r91 34 43 3.43356 $w=2.72e-07 $l=1.38109e-07 $layer=LI1_cond $X=1.78 $Y=1.035
+ $X2=1.882 $Y2=0.95
r92 34 42 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.78 $Y=1.035
+ $X2=1.78 $Y2=2.025
r93 30 43 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=1.882 $Y=0.865
+ $X2=1.882 $Y2=0.95
r94 30 32 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.882 $Y=0.865
+ $X2=1.882 $Y2=0.495
r95 26 41 1.37763 $w=4.33e-07 $l=5.2e-08 $layer=LI1_cond $X=1.647 $Y=2.242
+ $X2=1.647 $Y2=2.19
r96 26 28 17.4324 $w=4.33e-07 $l=6.58e-07 $layer=LI1_cond $X=1.647 $Y=2.242
+ $X2=1.647 $Y2=2.9
r97 25 46 53.3155 $w=3.55e-07 $l=3.28e-07 $layer=POLY_cond $X=3.012 $Y=1.358
+ $X2=3.012 $Y2=1.03
r98 22 46 2.43821 $w=3.55e-07 $l=1.5e-08 $layer=POLY_cond $X=3.012 $Y=1.015
+ $X2=3.012 $Y2=1.03
r99 22 23 147.677 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=3.012 $Y=0.94
+ $X2=3.3 $Y2=0.94
r100 19 22 52.3021 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=2.91 $Y=0.94
+ $X2=3.012 $Y2=0.94
r101 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.3 $Y=0.865
+ $X2=3.3 $Y2=0.94
r102 15 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.3 $Y=0.865
+ $X2=3.3 $Y2=0.495
r103 11 25 46.8051 $w=3.11e-07 $l=3.70689e-07 $layer=POLY_cond $X=3.165 $Y=1.66
+ $X2=3.012 $Y2=1.358
r104 11 13 219.881 $w=2.5e-07 $l=8.85e-07 $layer=POLY_cond $X=3.165 $Y=1.66
+ $X2=3.165 $Y2=2.545
r105 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.91 $Y=0.865
+ $X2=2.91 $Y2=0.94
r106 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.91 $Y=0.865
+ $X2=2.91 $Y2=0.495
r107 2 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=2.045 $X2=1.595 $Y2=2.19
r108 2 28 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=2.045 $X2=1.595 $Y2=2.9
r109 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.285 $X2=1.905 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_LP%VPWR 1 2 11 17 22 23 24 34 35 38
r37 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r39 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r40 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 29 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 26 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.825 $Y2=3.33
r45 26 28 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 24 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 24 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 22 31 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 22 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.9 $Y2=3.33
r50 21 34 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=3.6 $Y2=3.33
r51 21 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=2.9 $Y2=3.33
r52 17 20 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.9 $Y=2.19 $X2=2.9
+ $Y2=2.9
r53 15 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=3.245 $X2=2.9
+ $Y2=3.33
r54 15 20 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.9 $Y=3.245
+ $X2=2.9 $Y2=2.9
r55 11 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.825 $Y=2.19
+ $X2=0.825 $Y2=2.9
r56 9 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=3.33
r57 9 14 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=2.9
r58 2 20 400 $w=1.7e-07 $l=1.04614e-06 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=2.045 $X2=2.9 $Y2=2.9
r59 2 17 400 $w=1.7e-07 $l=4.92189e-07 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=2.045 $X2=2.9 $Y2=2.19
r60 1 14 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.045 $X2=0.825 $Y2=2.9
r61 1 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.045 $X2=0.825 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_LP%X 1 2 7 8 9 10 11 12 13 43
r18 43 44 0.727651 $w=4.48e-07 $l=1e-08 $layer=LI1_cond $X=3.49 $Y=2.035
+ $X2=3.49 $Y2=2.025
r19 34 47 1.59477 $w=4.48e-07 $l=6e-08 $layer=LI1_cond $X=3.49 $Y=2.25 $X2=3.49
+ $Y2=2.19
r20 13 40 3.32244 $w=4.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.49 $Y=2.775
+ $X2=3.49 $Y2=2.9
r21 12 13 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.49 $Y=2.405
+ $X2=3.49 $Y2=2.775
r22 12 34 4.11983 $w=4.48e-07 $l=1.55e-07 $layer=LI1_cond $X=3.49 $Y=2.405
+ $X2=3.49 $Y2=2.25
r23 11 47 3.13638 $w=4.48e-07 $l=1.18e-07 $layer=LI1_cond $X=3.49 $Y=2.072
+ $X2=3.49 $Y2=2.19
r24 11 43 0.983442 $w=4.48e-07 $l=3.7e-08 $layer=LI1_cond $X=3.49 $Y=2.072
+ $X2=3.49 $Y2=2.035
r25 11 44 1.1998 $w=3.63e-07 $l=3.8e-08 $layer=LI1_cond $X=3.532 $Y=1.987
+ $X2=3.532 $Y2=2.025
r26 10 11 10.1668 $w=3.63e-07 $l=3.22e-07 $layer=LI1_cond $X=3.532 $Y=1.665
+ $X2=3.532 $Y2=1.987
r27 9 10 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.532 $Y=1.295
+ $X2=3.532 $Y2=1.665
r28 8 9 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.532 $Y=0.925
+ $X2=3.532 $Y2=1.295
r29 7 8 13.5767 $w=3.63e-07 $l=4.3e-07 $layer=LI1_cond $X=3.532 $Y=0.495
+ $X2=3.532 $Y2=0.925
r30 2 47 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=2.045 $X2=3.43 $Y2=2.19
r31 2 40 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=2.045 $X2=3.43 $Y2=2.9
r32 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.285 $X2=3.515 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r52 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r53 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r55 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r56 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.695
+ $Y2=0
r57 27 29 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=3.6
+ $Y2=0
r58 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r59 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r60 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.085
+ $Y2=0
r61 23 25 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=2.16
+ $Y2=0
r62 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.695
+ $Y2=0
r63 22 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.16
+ $Y2=0
r64 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r65 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=1.085
+ $Y2=0
r67 17 19 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=0.72
+ $Y2=0
r68 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r69 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r70 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0.085
+ $X2=2.695 $Y2=0
r71 11 13 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.695 $Y=0.085
+ $X2=2.695 $Y2=0.475
r72 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=0.085
+ $X2=1.085 $Y2=0
r73 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.085 $Y=0.085
+ $X2=1.085 $Y2=0.455
r74 2 13 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.285 $X2=2.695 $Y2=0.475
r75 1 9 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=0.945
+ $Y=0.285 $X2=1.085 $Y2=0.455
.ends

