* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_86_275# D1 a_427_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_427_367# C1 a_499_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_86_275# A1 a_715_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND a_86_275# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_715_49# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND D1 a_86_275# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_86_275# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VGND B1 a_86_275# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR a_86_275# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR A2 a_607_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 X a_86_275# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 X a_86_275# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_607_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_499_367# B1 a_607_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
