* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_614_93# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_33_463# a_202_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR a_486_119# a_614_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR a_1175_417# a_1329_65# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR SET_B a_1175_417# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND D a_400_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_486_119# a_202_463# a_572_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_486_119# a_33_463# a_582_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_582_463# a_614_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1832_131# a_1175_417# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_614_93# a_486_119# a_853_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1287_91# a_1329_65# a_1359_91# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1175_417# a_33_463# a_985_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 VPWR a_1832_131# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_853_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1832_131# a_1175_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_1092_417# a_202_463# a_1175_417# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 VPWR a_486_119# a_985_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 a_1110_47# a_202_463# a_1175_417# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_1175_417# a_33_463# a_1287_91# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1359_91# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_33_463# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_33_463# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_1175_417# a_1329_65# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_33_463# a_202_463# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_1092_417# a_1329_65# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_400_119# a_33_463# a_486_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VGND a_486_119# a_1110_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 VGND a_1832_131# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 VPWR D a_400_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 a_400_119# a_202_463# a_486_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_572_119# a_614_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
