* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o221ai_m A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 Y C1 a_148_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_234_47# B2 a_148_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_148_47# B1 a_234_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_441_463# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR B1 a_245_480# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND A1 a_234_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 Y A2 a_441_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_234_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_245_480# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
