* File: sky130_fd_sc_lp__o211ai_m.spice
* Created: Fri Aug 28 11:03:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o211ai_m.pex.spice"
.subckt sky130_fd_sc_lp__o211ai_m  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A1_M1007_g N_A_29_47#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_A_29_47#_M1002_d N_A2_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 A_292_47# N_B1_M1005_g N_A_29_47#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_C1_M1006_g A_292_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 A_148_535# N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A2_M1004_g A_148_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_C1_M1001_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=9.3772 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
c_31 VNB 0 9.47829e-20 $X=0 $Y=0
c_56 VPB 0 1.69038e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o211ai_m.pxi.spice"
*
.ends
*
*
