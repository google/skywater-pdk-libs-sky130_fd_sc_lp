* File: sky130_fd_sc_lp__xor2_4.pxi.spice
* Created: Wed Sep  2 10:41:22 2020
* 
x_PM_SKY130_FD_SC_LP__XOR2_4%A N_A_M1012_g N_A_M1000_g N_A_M1020_g N_A_M1004_g
+ N_A_M1030_g N_A_M1014_g N_A_M1039_g N_A_M1037_g N_A_M1008_g N_A_M1006_g
+ N_A_M1017_g N_A_M1021_g N_A_M1018_g N_A_M1027_g N_A_M1034_g N_A_M1036_g
+ N_A_c_176_n N_A_c_177_n N_A_c_240_p N_A_c_178_n N_A_c_179_n N_A_c_180_n
+ N_A_c_181_n N_A_c_182_n N_A_c_183_n A N_A_c_185_n N_A_c_186_n N_A_c_187_n
+ N_A_c_188_n PM_SKY130_FD_SC_LP__XOR2_4%A
x_PM_SKY130_FD_SC_LP__XOR2_4%B N_B_M1007_g N_B_M1003_g N_B_M1016_g N_B_M1009_g
+ N_B_M1019_g N_B_M1025_g N_B_M1033_g N_B_M1032_g N_B_M1002_g N_B_M1001_g
+ N_B_M1015_g N_B_M1011_g N_B_M1028_g N_B_M1023_g N_B_M1029_g N_B_M1038_g
+ N_B_c_423_n N_B_c_424_n N_B_c_425_n N_B_c_438_n B N_B_c_440_n N_B_c_427_n
+ N_B_c_428_n PM_SKY130_FD_SC_LP__XOR2_4%B
x_PM_SKY130_FD_SC_LP__XOR2_4%A_776_255# N_A_776_255#_M1008_d
+ N_A_776_255#_M1018_d N_A_776_255#_M1002_s N_A_776_255#_M1028_s
+ N_A_776_255#_M1001_d N_A_776_255#_M1023_d N_A_776_255#_M1005_g
+ N_A_776_255#_M1013_g N_A_776_255#_M1010_g N_A_776_255#_M1024_g
+ N_A_776_255#_M1022_g N_A_776_255#_M1026_g N_A_776_255#_M1035_g
+ N_A_776_255#_M1031_g N_A_776_255#_c_634_n N_A_776_255#_c_635_n
+ N_A_776_255#_c_636_n N_A_776_255#_c_673_n N_A_776_255#_c_801_p
+ N_A_776_255#_c_826_p N_A_776_255#_c_677_n N_A_776_255#_c_822_p
+ N_A_776_255#_c_637_n N_A_776_255#_c_823_p N_A_776_255#_c_709_n
+ N_A_776_255#_c_638_n N_A_776_255#_c_649_n N_A_776_255#_c_650_n
+ N_A_776_255#_c_820_p N_A_776_255#_c_725_n N_A_776_255#_c_639_n
+ N_A_776_255#_c_651_n N_A_776_255#_c_640_n N_A_776_255#_c_686_n
+ N_A_776_255#_c_641_n N_A_776_255#_c_642_n N_A_776_255#_c_643_n
+ N_A_776_255#_c_653_n N_A_776_255#_c_644_n
+ PM_SKY130_FD_SC_LP__XOR2_4%A_776_255#
x_PM_SKY130_FD_SC_LP__XOR2_4%A_27_367# N_A_27_367#_M1000_s N_A_27_367#_M1004_s
+ N_A_27_367#_M1003_s N_A_27_367#_M1025_s N_A_27_367#_M1037_s
+ N_A_27_367#_M1010_d N_A_27_367#_M1035_d N_A_27_367#_c_850_n
+ N_A_27_367#_c_851_n N_A_27_367#_c_852_n N_A_27_367#_c_908_p
+ N_A_27_367#_c_860_n N_A_27_367#_c_909_p N_A_27_367#_c_875_n
+ N_A_27_367#_c_906_p N_A_27_367#_c_863_n N_A_27_367#_c_866_n
+ N_A_27_367#_c_911_p N_A_27_367#_c_892_n N_A_27_367#_c_853_n
+ N_A_27_367#_c_854_n N_A_27_367#_c_855_n N_A_27_367#_c_886_n
+ N_A_27_367#_c_888_n PM_SKY130_FD_SC_LP__XOR2_4%A_27_367#
x_PM_SKY130_FD_SC_LP__XOR2_4%VPWR N_VPWR_M1000_d N_VPWR_M1014_d N_VPWR_M1009_d
+ N_VPWR_M1032_d N_VPWR_M1006_d N_VPWR_M1027_d N_VPWR_c_940_n N_VPWR_c_941_n
+ N_VPWR_c_942_n N_VPWR_c_943_n N_VPWR_c_944_n N_VPWR_c_945_n N_VPWR_c_946_n
+ N_VPWR_c_947_n N_VPWR_c_948_n N_VPWR_c_949_n N_VPWR_c_950_n VPWR
+ N_VPWR_c_951_n N_VPWR_c_952_n N_VPWR_c_953_n N_VPWR_c_954_n N_VPWR_c_939_n
+ N_VPWR_c_956_n N_VPWR_c_957_n N_VPWR_c_958_n N_VPWR_c_959_n
+ PM_SKY130_FD_SC_LP__XOR2_4%VPWR
x_PM_SKY130_FD_SC_LP__XOR2_4%X N_X_M1007_d N_X_M1019_d N_X_M1013_s N_X_M1026_s
+ N_X_M1005_s N_X_M1022_s N_X_c_1082_n N_X_c_1105_n N_X_c_1078_n N_X_c_1145_p
+ N_X_c_1079_n N_X_c_1118_n N_X_c_1102_n N_X_c_1153_p N_X_c_1080_n X X X
+ N_X_c_1103_n PM_SKY130_FD_SC_LP__XOR2_4%X
x_PM_SKY130_FD_SC_LP__XOR2_4%A_1199_367# N_A_1199_367#_M1006_s
+ N_A_1199_367#_M1021_s N_A_1199_367#_M1036_s N_A_1199_367#_M1011_s
+ N_A_1199_367#_M1038_s N_A_1199_367#_c_1161_n N_A_1199_367#_c_1165_n
+ N_A_1199_367#_c_1162_n N_A_1199_367#_c_1207_n N_A_1199_367#_c_1170_n
+ N_A_1199_367#_c_1211_n N_A_1199_367#_c_1181_n N_A_1199_367#_c_1191_n
+ N_A_1199_367#_c_1183_n N_A_1199_367#_c_1163_n N_A_1199_367#_c_1164_n
+ N_A_1199_367#_c_1174_n N_A_1199_367#_c_1219_n
+ PM_SKY130_FD_SC_LP__XOR2_4%A_1199_367#
x_PM_SKY130_FD_SC_LP__XOR2_4%VGND N_VGND_M1012_s N_VGND_M1020_s N_VGND_M1039_s
+ N_VGND_M1024_d N_VGND_M1031_d N_VGND_M1017_s N_VGND_M1034_s N_VGND_M1015_d
+ N_VGND_M1029_d N_VGND_c_1221_n N_VGND_c_1222_n N_VGND_c_1223_n N_VGND_c_1224_n
+ N_VGND_c_1225_n N_VGND_c_1226_n N_VGND_c_1227_n N_VGND_c_1228_n
+ N_VGND_c_1229_n N_VGND_c_1230_n N_VGND_c_1231_n N_VGND_c_1232_n
+ N_VGND_c_1233_n N_VGND_c_1234_n N_VGND_c_1235_n N_VGND_c_1236_n
+ N_VGND_c_1237_n VGND N_VGND_c_1238_n N_VGND_c_1239_n N_VGND_c_1240_n
+ N_VGND_c_1241_n N_VGND_c_1242_n N_VGND_c_1243_n N_VGND_c_1244_n
+ N_VGND_c_1245_n N_VGND_c_1246_n N_VGND_c_1247_n N_VGND_c_1248_n
+ PM_SKY130_FD_SC_LP__XOR2_4%VGND
x_PM_SKY130_FD_SC_LP__XOR2_4%A_110_47# N_A_110_47#_M1012_d N_A_110_47#_M1030_d
+ N_A_110_47#_M1016_s N_A_110_47#_M1033_s N_A_110_47#_c_1393_n
+ N_A_110_47#_c_1428_n N_A_110_47#_c_1400_n N_A_110_47#_c_1406_n
+ N_A_110_47#_c_1407_n N_A_110_47#_c_1412_n PM_SKY130_FD_SC_LP__XOR2_4%A_110_47#
cc_1 VNB N_A_M1012_g 0.028051f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A_M1000_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_A_M1020_g 0.0207288f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_4 VNB N_A_M1004_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_5 VNB N_A_M1030_g 0.0196233f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_6 VNB N_A_M1014_g 0.00256887f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_7 VNB N_A_M1037_g 0.0070956f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=2.465
cc_8 VNB N_A_M1008_g 0.0235727f $X=-0.19 $Y=-0.245 $X2=6.265 $Y2=0.655
cc_9 VNB N_A_M1006_g 0.00309338f $X=-0.19 $Y=-0.245 $X2=6.335 $Y2=2.465
cc_10 VNB N_A_M1017_g 0.019861f $X=-0.19 $Y=-0.245 $X2=6.695 $Y2=0.655
cc_11 VNB N_A_M1021_g 0.00209543f $X=-0.19 $Y=-0.245 $X2=6.765 $Y2=2.465
cc_12 VNB N_A_M1018_g 0.0202259f $X=-0.19 $Y=-0.245 $X2=7.125 $Y2=0.655
cc_13 VNB N_A_M1027_g 0.00209543f $X=-0.19 $Y=-0.245 $X2=7.195 $Y2=2.465
cc_14 VNB N_A_M1034_g 0.0197943f $X=-0.19 $Y=-0.245 $X2=7.555 $Y2=0.655
cc_15 VNB N_A_M1036_g 0.00211543f $X=-0.19 $Y=-0.245 $X2=7.625 $Y2=2.465
cc_16 VNB N_A_c_176_n 0.0101004f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.4
cc_17 VNB N_A_c_177_n 0.0215617f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=1.16
cc_18 VNB N_A_c_178_n 0.00496906f $X=-0.19 $Y=-0.245 $X2=1.407 $Y2=1.16
cc_19 VNB N_A_c_179_n 0.00222881f $X=-0.19 $Y=-0.245 $X2=6.908 $Y2=1.367
cc_20 VNB N_A_c_180_n 0.00131986f $X=-0.19 $Y=-0.245 $X2=7.075 $Y2=1.367
cc_21 VNB N_A_c_181_n 0.0121773f $X=-0.19 $Y=-0.245 $X2=6.335 $Y2=1.295
cc_22 VNB N_A_c_182_n 0.00154102f $X=-0.19 $Y=-0.245 $X2=3.745 $Y2=1.295
cc_23 VNB N_A_c_183_n 0.00421727f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=1.295
cc_24 VNB A 0.00197311f $X=-0.19 $Y=-0.245 $X2=6.395 $Y2=1.21
cc_25 VNB N_A_c_185_n 0.0617134f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.44
cc_26 VNB N_A_c_186_n 0.0303956f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.35
cc_27 VNB N_A_c_187_n 0.0160285f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.185
cc_28 VNB N_A_c_188_n 0.0868856f $X=-0.19 $Y=-0.245 $X2=7.625 $Y2=1.44
cc_29 VNB N_B_M1007_g 0.0221857f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_30 VNB N_B_M1016_g 0.0220935f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_31 VNB N_B_M1019_g 0.0220935f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_32 VNB N_B_M1033_g 0.0217136f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=0.655
cc_33 VNB N_B_M1002_g 0.0197997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_M1001_g 0.00229065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_M1015_g 0.0196295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_M1011_g 0.00248813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_M1028_g 0.0196295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_B_M1023_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_M1029_g 0.0240669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_B_M1038_g 0.00287449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_B_c_423_n 0.00167151f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.44
cc_42 VNB N_B_c_424_n 0.0991105f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.44
cc_43 VNB N_B_c_425_n 0.00535061f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.16
cc_44 VNB B 0.00113317f $X=-0.19 $Y=-0.245 $X2=1.407 $Y2=1.16
cc_45 VNB N_B_c_427_n 0.0689381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_B_c_428_n 0.00333044f $X=-0.19 $Y=-0.245 $X2=6.695 $Y2=1.44
cc_47 VNB N_A_776_255#_M1005_g 0.00212819f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=1.605
cc_48 VNB N_A_776_255#_M1013_g 0.0202016f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=1.185
cc_49 VNB N_A_776_255#_M1010_g 0.00209543f $X=-0.19 $Y=-0.245 $X2=3.515
+ $Y2=2.465
cc_50 VNB N_A_776_255#_M1024_g 0.0191498f $X=-0.19 $Y=-0.245 $X2=6.265 $Y2=0.655
cc_51 VNB N_A_776_255#_M1022_g 0.00209543f $X=-0.19 $Y=-0.245 $X2=6.335
+ $Y2=2.465
cc_52 VNB N_A_776_255#_M1026_g 0.0192139f $X=-0.19 $Y=-0.245 $X2=6.695 $Y2=0.655
cc_53 VNB N_A_776_255#_M1035_g 0.00309338f $X=-0.19 $Y=-0.245 $X2=6.765
+ $Y2=2.465
cc_54 VNB N_A_776_255#_M1031_g 0.0246947f $X=-0.19 $Y=-0.245 $X2=7.125 $Y2=0.655
cc_55 VNB N_A_776_255#_c_634_n 0.00368483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_776_255#_c_635_n 0.0613877f $X=-0.19 $Y=-0.245 $X2=7.555 $Y2=0.655
cc_57 VNB N_A_776_255#_c_636_n 0.00435356f $X=-0.19 $Y=-0.245 $X2=7.625
+ $Y2=1.605
cc_58 VNB N_A_776_255#_c_637_n 0.00375136f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.16
cc_59 VNB N_A_776_255#_c_638_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=6.908
+ $Y2=1.367
cc_60 VNB N_A_776_255#_c_639_n 0.0270824f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.44
cc_61 VNB N_A_776_255#_c_640_n 0.0246478f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.35
cc_62 VNB N_A_776_255#_c_641_n 0.00248817f $X=-0.19 $Y=-0.245 $X2=3.505
+ $Y2=1.515
cc_63 VNB N_A_776_255#_c_642_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=6.335 $Y2=1.44
cc_64 VNB N_A_776_255#_c_643_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=6.47 $Y2=1.44
cc_65 VNB N_A_776_255#_c_644_n 0.0781208f $X=-0.19 $Y=-0.245 $X2=6.47 $Y2=1.44
cc_66 VNB N_VPWR_c_939_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_X_c_1078_n 0.00166317f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.515
cc_68 VNB N_X_c_1079_n 0.00497019f $X=-0.19 $Y=-0.245 $X2=6.265 $Y2=0.655
cc_69 VNB N_X_c_1080_n 4.28853e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1221_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.515
cc_71 VNB N_VGND_c_1222_n 0.0408474f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=2.465
cc_72 VNB N_VGND_c_1223_n 0.0043494f $X=-0.19 $Y=-0.245 $X2=6.265 $Y2=0.655
cc_73 VNB N_VGND_c_1224_n 0.00269335f $X=-0.19 $Y=-0.245 $X2=6.335 $Y2=2.465
cc_74 VNB N_VGND_c_1225_n 3.08929e-19 $X=-0.19 $Y=-0.245 $X2=6.695 $Y2=0.655
cc_75 VNB N_VGND_c_1226_n 0.00199238f $X=-0.19 $Y=-0.245 $X2=6.765 $Y2=2.465
cc_76 VNB N_VGND_c_1227_n 3.08929e-19 $X=-0.19 $Y=-0.245 $X2=7.125 $Y2=0.655
cc_77 VNB N_VGND_c_1228_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=7.195 $Y2=2.465
cc_78 VNB N_VGND_c_1229_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=7.555 $Y2=0.655
cc_79 VNB N_VGND_c_1230_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=7.625 $Y2=1.605
cc_80 VNB N_VGND_c_1231_n 0.0264919f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.4
cc_81 VNB N_VGND_c_1232_n 0.0547364f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.44
cc_82 VNB N_VGND_c_1233_n 0.00510143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1234_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.44
cc_84 VNB N_VGND_c_1235_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.44
cc_85 VNB N_VGND_c_1236_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=1.16
cc_86 VNB N_VGND_c_1237_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.16
cc_87 VNB N_VGND_c_1238_n 0.0139945f $X=-0.19 $Y=-0.245 $X2=7.49 $Y2=1.44
cc_88 VNB N_VGND_c_1239_n 0.012251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1240_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1241_n 0.0156676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1242_n 0.480575f $X=-0.19 $Y=-0.245 $X2=6.335 $Y2=1.44
cc_92 VNB N_VGND_c_1243_n 0.00439334f $X=-0.19 $Y=-0.245 $X2=6.81 $Y2=1.44
cc_93 VNB N_VGND_c_1244_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=7.125 $Y2=1.44
cc_94 VNB N_VGND_c_1245_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=7.625 $Y2=1.44
cc_95 VNB N_VGND_c_1246_n 0.0176477f $X=-0.19 $Y=-0.245 $X2=3.512 $Y2=1.295
cc_96 VNB N_VGND_c_1247_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=6.48 $Y2=1.295
cc_97 VNB N_VGND_c_1248_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_110_47#_c_1393_n 0.00184664f $X=-0.19 $Y=-0.245 $X2=0.905
+ $Y2=1.605
cc_99 VPB N_A_M1000_g 0.0243928f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_100 VPB N_A_M1004_g 0.0184123f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_101 VPB N_A_M1014_g 0.0198547f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_102 VPB N_A_M1037_g 0.0199867f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=2.465
cc_103 VPB N_A_M1006_g 0.0258837f $X=-0.19 $Y=1.655 $X2=6.335 $Y2=2.465
cc_104 VPB N_A_M1021_g 0.0189697f $X=-0.19 $Y=1.655 $X2=6.765 $Y2=2.465
cc_105 VPB N_A_M1027_g 0.018968f $X=-0.19 $Y=1.655 $X2=7.195 $Y2=2.465
cc_106 VPB N_A_M1036_g 0.0192041f $X=-0.19 $Y=1.655 $X2=7.625 $Y2=2.465
cc_107 VPB N_B_M1003_g 0.0183924f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_108 VPB N_B_M1009_g 0.0177297f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_109 VPB N_B_M1025_g 0.0176811f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_110 VPB N_B_M1032_g 0.0185221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_B_M1001_g 0.019292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_B_M1011_g 0.018687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_B_M1023_g 0.0186909f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_B_M1038_g 0.0236764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_B_c_425_n 0.035284f $X=-0.19 $Y=1.655 $X2=1.555 $Y2=1.16
cc_116 VPB N_B_c_438_n 0.0011832f $X=-0.19 $Y=1.655 $X2=7.075 $Y2=1.445
cc_117 VPB B 0.00104138f $X=-0.19 $Y=1.655 $X2=1.407 $Y2=1.16
cc_118 VPB N_B_c_440_n 0.00698679f $X=-0.19 $Y=1.655 $X2=6.395 $Y2=1.21
cc_119 VPB N_B_c_427_n 0.0123334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_B_c_428_n 0.004546f $X=-0.19 $Y=1.655 $X2=6.695 $Y2=1.44
cc_121 VPB N_A_776_255#_M1005_g 0.0190996f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.605
cc_122 VPB N_A_776_255#_M1010_g 0.0191366f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=2.465
cc_123 VPB N_A_776_255#_M1022_g 0.019163f $X=-0.19 $Y=1.655 $X2=6.335 $Y2=2.465
cc_124 VPB N_A_776_255#_M1035_g 0.0258905f $X=-0.19 $Y=1.655 $X2=6.765 $Y2=2.465
cc_125 VPB N_A_776_255#_c_649_n 0.00223864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_776_255#_c_650_n 0.00276981f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_776_255#_c_651_n 0.0234352f $X=-0.19 $Y=1.655 $X2=1.245 $Y2=1.44
cc_128 VPB N_A_776_255#_c_640_n 0.00269647f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=1.35
cc_129 VPB N_A_776_255#_c_653_n 0.00228829f $X=-0.19 $Y=1.655 $X2=6.47 $Y2=1.44
cc_130 VPB N_A_27_367#_c_850_n 0.0457879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_27_367#_c_851_n 0.00362418f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=1.515
cc_132 VPB N_A_27_367#_c_852_n 0.0118541f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=2.465
cc_133 VPB N_A_27_367#_c_853_n 0.00370134f $X=-0.19 $Y=1.655 $X2=7.195 $Y2=2.465
cc_134 VPB N_A_27_367#_c_854_n 0.0133259f $X=-0.19 $Y=1.655 $X2=7.555 $Y2=1.275
cc_135 VPB N_A_27_367#_c_855_n 0.00314784f $X=-0.19 $Y=1.655 $X2=7.555 $Y2=0.655
cc_136 VPB N_VPWR_c_940_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.605
cc_137 VPB N_VPWR_c_941_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=3.485 $Y2=0.655
cc_138 VPB N_VPWR_c_942_n 3.11777e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_943_n 0.013276f $X=-0.19 $Y=1.655 $X2=6.265 $Y2=0.655
cc_140 VPB N_VPWR_c_944_n 4.01796e-19 $X=-0.19 $Y=1.655 $X2=6.335 $Y2=2.465
cc_141 VPB N_VPWR_c_945_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=6.695 $Y2=0.655
cc_142 VPB N_VPWR_c_946_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=6.765 $Y2=2.465
cc_143 VPB N_VPWR_c_947_n 0.0129398f $X=-0.19 $Y=1.655 $X2=7.125 $Y2=1.275
cc_144 VPB N_VPWR_c_948_n 0.00436868f $X=-0.19 $Y=1.655 $X2=7.125 $Y2=0.655
cc_145 VPB N_VPWR_c_949_n 0.0129398f $X=-0.19 $Y=1.655 $X2=7.125 $Y2=0.655
cc_146 VPB N_VPWR_c_950_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_951_n 0.0153759f $X=-0.19 $Y=1.655 $X2=7.195 $Y2=2.465
cc_148 VPB N_VPWR_c_952_n 0.0694907f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.44
cc_149 VPB N_VPWR_c_953_n 0.0129398f $X=-0.19 $Y=1.655 $X2=7.075 $Y2=1.445
cc_150 VPB N_VPWR_c_954_n 0.061676f $X=-0.19 $Y=1.655 $X2=7.075 $Y2=1.367
cc_151 VPB N_VPWR_c_939_n 0.0711167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_956_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.745 $Y2=1.295
cc_153 VPB N_VPWR_c_957_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.6 $Y2=1.295
cc_154 VPB N_VPWR_c_958_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_959_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.44
cc_156 VPB N_X_c_1078_n 0.00209795f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=1.515
cc_157 VPB N_A_1199_367#_c_1161_n 0.0106879f $X=-0.19 $Y=1.655 $X2=1.335
+ $Y2=0.655
cc_158 VPB N_A_1199_367#_c_1162_n 0.00237364f $X=-0.19 $Y=1.655 $X2=1.335
+ $Y2=2.465
cc_159 VPB N_A_1199_367#_c_1163_n 0.00746637f $X=-0.19 $Y=1.655 $X2=6.695
+ $Y2=0.655
cc_160 VPB N_A_1199_367#_c_1164_n 0.032697f $X=-0.19 $Y=1.655 $X2=6.765
+ $Y2=1.605
cc_161 N_A_M1030_g N_B_M1007_g 0.0263035f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A_c_177_n N_B_M1007_g 0.0110396f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_c_178_n N_B_M1007_g 0.00460636f $X=1.407 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_c_183_n N_B_M1007_g 0.00123709f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_165 N_A_M1014_g N_B_M1003_g 0.0263035f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A_c_177_n N_B_M1016_g 0.00952628f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_c_183_n N_B_M1016_g 0.00122391f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_168 N_A_c_177_n N_B_M1019_g 0.00952628f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_c_183_n N_B_M1019_g 0.00122391f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_170 N_A_c_177_n N_B_M1033_g 0.0117228f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_c_183_n N_B_M1033_g 0.00110395f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_172 N_A_c_186_n N_B_M1033_g 0.022994f $X=3.505 $Y=1.35 $X2=0 $Y2=0
cc_173 N_A_c_187_n N_B_M1033_g 0.0356721f $X=3.505 $Y=1.185 $X2=0 $Y2=0
cc_174 N_A_M1034_g N_B_M1002_g 0.0205379f $X=7.555 $Y=0.655 $X2=0 $Y2=0
cc_175 N_A_M1036_g N_B_M1001_g 0.0249865f $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_c_188_n N_B_c_424_n 0.0232454f $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_177 N_A_M1037_g N_B_c_425_n 0.00509513f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_M1006_g N_B_c_425_n 0.00517919f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A_M1021_g N_B_c_425_n 0.0038895f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_M1027_g N_B_c_425_n 0.0038895f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A_M1036_g N_B_c_425_n 0.00391464f $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A_c_177_n N_B_c_425_n 0.00572269f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_c_179_n N_B_c_425_n 0.0333091f $X=6.908 $Y=1.367 $X2=0 $Y2=0
cc_184 N_A_c_181_n N_B_c_425_n 0.188841f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_185 N_A_c_182_n N_B_c_425_n 0.0244797f $X=3.745 $Y=1.295 $X2=0 $Y2=0
cc_186 N_A_c_183_n N_B_c_425_n 0.0498264f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_187 A N_B_c_425_n 0.0239851f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A_c_186_n N_B_c_425_n 0.00303998f $X=3.505 $Y=1.35 $X2=0 $Y2=0
cc_189 N_A_c_188_n N_B_c_425_n 0.0160603f $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_190 N_A_c_177_n N_B_c_438_n 3.30608e-19 $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_c_183_n N_B_c_438_n 0.0239841f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_192 N_A_M1036_g B 7.34611e-19 $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A_c_188_n B 7.62495e-19 $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_194 N_A_M1037_g N_B_c_440_n 0.00194885f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A_c_177_n N_B_c_440_n 0.0871971f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_c_178_n N_B_c_440_n 0.0086846f $X=1.407 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_c_183_n N_B_c_440_n 0.0234993f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_198 N_A_c_185_n N_B_c_440_n 0.00141108f $X=1.335 $Y=1.44 $X2=0 $Y2=0
cc_199 N_A_c_186_n N_B_c_440_n 5.69001e-19 $X=3.505 $Y=1.35 $X2=0 $Y2=0
cc_200 N_A_M1037_g N_B_c_427_n 0.0418802f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_201 N_A_c_177_n N_B_c_427_n 0.00565725f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A_c_183_n N_B_c_427_n 0.0150086f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_203 N_A_c_185_n N_B_c_427_n 0.0263035f $X=1.335 $Y=1.44 $X2=0 $Y2=0
cc_204 N_A_c_240_p N_B_c_428_n 0.0143389f $X=7.49 $Y=1.44 $X2=0 $Y2=0
cc_205 N_A_c_188_n N_B_c_428_n 0.00619014f $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_206 N_A_c_177_n N_A_776_255#_M1013_g 0.00129174f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_c_181_n N_A_776_255#_M1013_g 0.00118055f $X=6.335 $Y=1.295 $X2=0
+ $Y2=0
cc_208 N_A_c_182_n N_A_776_255#_M1013_g 6.79515e-19 $X=3.745 $Y=1.295 $X2=0
+ $Y2=0
cc_209 N_A_c_186_n N_A_776_255#_M1013_g 0.00484934f $X=3.505 $Y=1.35 $X2=0 $Y2=0
cc_210 N_A_c_187_n N_A_776_255#_M1013_g 0.0297276f $X=3.505 $Y=1.185 $X2=0 $Y2=0
cc_211 N_A_c_181_n N_A_776_255#_M1024_g 0.00198208f $X=6.335 $Y=1.295 $X2=0
+ $Y2=0
cc_212 N_A_c_181_n N_A_776_255#_M1026_g 0.0020293f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_213 N_A_c_181_n N_A_776_255#_M1031_g 0.0066385f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_214 N_A_c_179_n N_A_776_255#_c_634_n 0.0154027f $X=6.908 $Y=1.367 $X2=0 $Y2=0
cc_215 N_A_c_181_n N_A_776_255#_c_634_n 0.0351699f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_216 A N_A_776_255#_c_634_n 3.51154e-19 $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_217 N_A_c_188_n N_A_776_255#_c_634_n 0.00179045f $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_218 N_A_c_179_n N_A_776_255#_c_635_n 2.30261e-19 $X=6.908 $Y=1.367 $X2=0
+ $Y2=0
cc_219 N_A_c_181_n N_A_776_255#_c_635_n 0.00417412f $X=6.335 $Y=1.295 $X2=0
+ $Y2=0
cc_220 N_A_c_188_n N_A_776_255#_c_635_n 0.0161402f $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_221 N_A_M1008_g N_A_776_255#_c_636_n 0.00812351f $X=6.265 $Y=0.655 $X2=0
+ $Y2=0
cc_222 N_A_c_179_n N_A_776_255#_c_636_n 0.0107931f $X=6.908 $Y=1.367 $X2=0 $Y2=0
cc_223 N_A_c_181_n N_A_776_255#_c_636_n 0.0152409f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_224 A N_A_776_255#_c_636_n 0.00114706f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_225 N_A_M1008_g N_A_776_255#_c_673_n 0.0114563f $X=6.265 $Y=0.655 $X2=0 $Y2=0
cc_226 N_A_c_179_n N_A_776_255#_c_673_n 0.00385582f $X=6.908 $Y=1.367 $X2=0
+ $Y2=0
cc_227 N_A_c_181_n N_A_776_255#_c_673_n 0.00685668f $X=6.335 $Y=1.295 $X2=0
+ $Y2=0
cc_228 A N_A_776_255#_c_673_n 0.00137504f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_229 N_A_M1017_g N_A_776_255#_c_677_n 0.00967899f $X=6.695 $Y=0.655 $X2=0
+ $Y2=0
cc_230 N_A_M1018_g N_A_776_255#_c_677_n 0.0104705f $X=7.125 $Y=0.655 $X2=0 $Y2=0
cc_231 N_A_c_240_p N_A_776_255#_c_677_n 0.0053926f $X=7.49 $Y=1.44 $X2=0 $Y2=0
cc_232 N_A_c_179_n N_A_776_255#_c_677_n 0.0310252f $X=6.908 $Y=1.367 $X2=0 $Y2=0
cc_233 A N_A_776_255#_c_677_n 0.00137504f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_234 N_A_c_188_n N_A_776_255#_c_677_n 5.91523e-19 $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_235 N_A_M1034_g N_A_776_255#_c_637_n 0.0126915f $X=7.555 $Y=0.655 $X2=0 $Y2=0
cc_236 N_A_c_240_p N_A_776_255#_c_637_n 0.0144914f $X=7.49 $Y=1.44 $X2=0 $Y2=0
cc_237 N_A_c_188_n N_A_776_255#_c_637_n 0.00276121f $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_238 N_A_c_179_n N_A_776_255#_c_686_n 0.0128846f $X=6.908 $Y=1.367 $X2=0 $Y2=0
cc_239 A N_A_776_255#_c_686_n 0.0055226f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_240 N_A_c_188_n N_A_776_255#_c_686_n 6.47713e-19 $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_241 N_A_M1018_g N_A_776_255#_c_641_n 0.00269527f $X=7.125 $Y=0.655 $X2=0
+ $Y2=0
cc_242 N_A_M1034_g N_A_776_255#_c_641_n 2.39567e-19 $X=7.555 $Y=0.655 $X2=0
+ $Y2=0
cc_243 N_A_c_240_p N_A_776_255#_c_641_n 0.0143841f $X=7.49 $Y=1.44 $X2=0 $Y2=0
cc_244 N_A_c_188_n N_A_776_255#_c_641_n 0.00286879f $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_245 N_A_M1037_g N_A_776_255#_c_644_n 0.0261443f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A_c_177_n N_A_776_255#_c_644_n 9.70067e-19 $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_c_181_n N_A_776_255#_c_644_n 0.00559541f $X=6.335 $Y=1.295 $X2=0
+ $Y2=0
cc_248 N_A_c_182_n N_A_776_255#_c_644_n 7.28461e-19 $X=3.745 $Y=1.295 $X2=0
+ $Y2=0
cc_249 N_A_c_186_n N_A_776_255#_c_644_n 0.0167337f $X=3.505 $Y=1.35 $X2=0 $Y2=0
cc_250 N_A_M1000_g N_A_27_367#_c_851_n 0.0150277f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A_M1004_g N_A_27_367#_c_851_n 0.0128944f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_252 N_A_c_176_n N_A_27_367#_c_851_n 0.0448757f $X=1.26 $Y=1.4 $X2=0 $Y2=0
cc_253 N_A_c_185_n N_A_27_367#_c_851_n 0.00246472f $X=1.335 $Y=1.44 $X2=0 $Y2=0
cc_254 N_A_M1014_g N_A_27_367#_c_860_n 0.0134728f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_255 N_A_c_178_n N_A_27_367#_c_860_n 0.0089841f $X=1.407 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A_c_183_n N_A_27_367#_c_860_n 0.00697024f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_257 N_A_M1037_g N_A_27_367#_c_863_n 0.0142193f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A_c_177_n N_A_27_367#_c_863_n 0.00309534f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_c_186_n N_A_27_367#_c_863_n 0.00179192f $X=3.505 $Y=1.35 $X2=0 $Y2=0
cc_260 N_A_c_177_n N_A_27_367#_c_866_n 7.43166e-19 $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_c_186_n N_A_27_367#_c_866_n 8.08263e-19 $X=3.505 $Y=1.35 $X2=0 $Y2=0
cc_262 N_A_M1006_g N_A_27_367#_c_854_n 0.00388976f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A_M1004_g N_A_27_367#_c_855_n 3.05538e-19 $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A_M1014_g N_A_27_367#_c_855_n 0.00247677f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A_c_176_n N_A_27_367#_c_855_n 0.0163587f $X=1.26 $Y=1.4 $X2=0 $Y2=0
cc_266 N_A_c_185_n N_A_27_367#_c_855_n 0.00256759f $X=1.335 $Y=1.44 $X2=0 $Y2=0
cc_267 N_A_M1000_g N_VPWR_c_940_n 0.0174402f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A_M1004_g N_VPWR_c_940_n 0.0154271f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A_M1014_g N_VPWR_c_940_n 7.21796e-19 $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_270 N_A_M1004_g N_VPWR_c_941_n 6.73419e-19 $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_271 N_A_M1014_g N_VPWR_c_941_n 0.0142626f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A_M1037_g N_VPWR_c_944_n 0.0146175f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A_M1006_g N_VPWR_c_945_n 0.0156533f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_274 N_A_M1021_g N_VPWR_c_945_n 0.0137908f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A_M1027_g N_VPWR_c_945_n 6.66346e-19 $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A_M1021_g N_VPWR_c_946_n 6.66346e-19 $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A_M1027_g N_VPWR_c_946_n 0.0137908f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_278 N_A_M1036_g N_VPWR_c_946_n 0.0149637f $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_279 N_A_M1004_g N_VPWR_c_947_n 0.00486043f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_280 N_A_M1014_g N_VPWR_c_947_n 0.00486043f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_281 N_A_M1000_g N_VPWR_c_951_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_282 N_A_M1037_g N_VPWR_c_952_n 0.00544582f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_283 N_A_M1006_g N_VPWR_c_952_n 0.00486043f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_284 N_A_M1021_g N_VPWR_c_953_n 0.00486043f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_285 N_A_M1027_g N_VPWR_c_953_n 0.00486043f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A_M1036_g N_VPWR_c_954_n 0.00486043f $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A_M1000_g N_VPWR_c_939_n 0.00917987f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_288 N_A_M1004_g N_VPWR_c_939_n 0.00824727f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_289 N_A_M1014_g N_VPWR_c_939_n 0.00824727f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_290 N_A_M1037_g N_VPWR_c_939_n 0.0092234f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A_M1006_g N_VPWR_c_939_n 0.00954696f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A_M1021_g N_VPWR_c_939_n 0.00824727f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A_M1027_g N_VPWR_c_939_n 0.00824727f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A_M1036_g N_VPWR_c_939_n 0.0082726f $X=7.625 $Y=2.465 $X2=0 $Y2=0
cc_295 N_A_c_177_n N_X_c_1082_n 0.111937f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_c_181_n N_X_c_1082_n 0.00936877f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_297 N_A_c_182_n N_X_c_1082_n 0.00398601f $X=3.745 $Y=1.295 $X2=0 $Y2=0
cc_298 N_A_c_183_n N_X_c_1082_n 0.00878377f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_299 N_A_c_186_n N_X_c_1082_n 7.55146e-19 $X=3.505 $Y=1.35 $X2=0 $Y2=0
cc_300 N_A_c_187_n N_X_c_1082_n 0.0136918f $X=3.505 $Y=1.185 $X2=0 $Y2=0
cc_301 N_A_M1037_g N_X_c_1078_n 0.00244561f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A_c_181_n N_X_c_1078_n 0.0296506f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_303 N_A_c_182_n N_X_c_1078_n 0.00124833f $X=3.745 $Y=1.295 $X2=0 $Y2=0
cc_304 N_A_c_186_n N_X_c_1078_n 8.12771e-19 $X=3.505 $Y=1.35 $X2=0 $Y2=0
cc_305 N_A_c_181_n N_X_c_1079_n 0.0271594f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_306 N_A_c_177_n N_X_c_1080_n 0.0147052f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_307 N_A_c_181_n N_X_c_1080_n 0.00114401f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_308 N_A_c_182_n N_X_c_1080_n 0.00124463f $X=3.745 $Y=1.295 $X2=0 $Y2=0
cc_309 N_A_c_187_n N_X_c_1080_n 0.00108173f $X=3.505 $Y=1.185 $X2=0 $Y2=0
cc_310 N_A_M1006_g N_A_1199_367#_c_1165_n 0.0143192f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A_M1021_g N_A_1199_367#_c_1165_n 0.0134161f $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_312 N_A_c_179_n N_A_1199_367#_c_1165_n 0.00816101f $X=6.908 $Y=1.367 $X2=0
+ $Y2=0
cc_313 N_A_c_188_n N_A_1199_367#_c_1165_n 0.00147896f $X=7.625 $Y=1.44 $X2=0
+ $Y2=0
cc_314 N_A_c_188_n N_A_1199_367#_c_1162_n 5.45485e-19 $X=7.625 $Y=1.44 $X2=0
+ $Y2=0
cc_315 N_A_M1027_g N_A_1199_367#_c_1170_n 0.0133695f $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_316 N_A_M1036_g N_A_1199_367#_c_1170_n 0.0136351f $X=7.625 $Y=2.465 $X2=0
+ $Y2=0
cc_317 N_A_c_240_p N_A_1199_367#_c_1170_n 0.00773808f $X=7.49 $Y=1.44 $X2=0
+ $Y2=0
cc_318 N_A_c_188_n N_A_1199_367#_c_1170_n 0.00147896f $X=7.625 $Y=1.44 $X2=0
+ $Y2=0
cc_319 N_A_c_179_n N_A_1199_367#_c_1174_n 0.00339029f $X=6.908 $Y=1.367 $X2=0
+ $Y2=0
cc_320 N_A_c_188_n N_A_1199_367#_c_1174_n 0.00162f $X=7.625 $Y=1.44 $X2=0 $Y2=0
cc_321 N_A_c_177_n N_VGND_M1039_s 0.00134915f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A_M1012_g N_VGND_c_1222_n 0.0175764f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_323 N_A_M1020_g N_VGND_c_1222_n 5.98206e-19 $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_324 N_A_c_176_n N_VGND_c_1222_n 0.00179347f $X=1.26 $Y=1.4 $X2=0 $Y2=0
cc_325 N_A_M1020_g N_VGND_c_1223_n 0.001584f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_326 N_A_M1030_g N_VGND_c_1223_n 0.00285858f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_327 N_A_c_187_n N_VGND_c_1224_n 0.00457506f $X=3.505 $Y=1.185 $X2=0 $Y2=0
cc_328 N_A_M1008_g N_VGND_c_1226_n 0.0042091f $X=6.265 $Y=0.655 $X2=0 $Y2=0
cc_329 N_A_c_181_n N_VGND_c_1226_n 0.00938257f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_330 N_A_M1008_g N_VGND_c_1227_n 5.72576e-19 $X=6.265 $Y=0.655 $X2=0 $Y2=0
cc_331 N_A_M1017_g N_VGND_c_1227_n 0.0103386f $X=6.695 $Y=0.655 $X2=0 $Y2=0
cc_332 N_A_M1018_g N_VGND_c_1227_n 0.0103489f $X=7.125 $Y=0.655 $X2=0 $Y2=0
cc_333 N_A_M1034_g N_VGND_c_1227_n 5.72987e-19 $X=7.555 $Y=0.655 $X2=0 $Y2=0
cc_334 N_A_M1018_g N_VGND_c_1228_n 6.16837e-19 $X=7.125 $Y=0.655 $X2=0 $Y2=0
cc_335 N_A_M1034_g N_VGND_c_1228_n 0.0102423f $X=7.555 $Y=0.655 $X2=0 $Y2=0
cc_336 N_A_M1030_g N_VGND_c_1232_n 0.00425616f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_337 N_A_c_187_n N_VGND_c_1232_n 0.00421077f $X=3.505 $Y=1.185 $X2=0 $Y2=0
cc_338 N_A_M1018_g N_VGND_c_1234_n 0.00486043f $X=7.125 $Y=0.655 $X2=0 $Y2=0
cc_339 N_A_M1034_g N_VGND_c_1234_n 0.00486043f $X=7.555 $Y=0.655 $X2=0 $Y2=0
cc_340 N_A_M1012_g N_VGND_c_1238_n 0.00486043f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_341 N_A_M1020_g N_VGND_c_1238_n 0.00439206f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_342 N_A_M1008_g N_VGND_c_1240_n 0.00486043f $X=6.265 $Y=0.655 $X2=0 $Y2=0
cc_343 N_A_M1017_g N_VGND_c_1240_n 0.00486043f $X=6.695 $Y=0.655 $X2=0 $Y2=0
cc_344 N_A_M1012_g N_VGND_c_1242_n 0.00824727f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_345 N_A_M1020_g N_VGND_c_1242_n 0.00586174f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_346 N_A_M1030_g N_VGND_c_1242_n 0.00586053f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_347 N_A_M1008_g N_VGND_c_1242_n 0.00456312f $X=6.265 $Y=0.655 $X2=0 $Y2=0
cc_348 N_A_M1017_g N_VGND_c_1242_n 0.00458264f $X=6.695 $Y=0.655 $X2=0 $Y2=0
cc_349 N_A_M1018_g N_VGND_c_1242_n 0.00458264f $X=7.125 $Y=0.655 $X2=0 $Y2=0
cc_350 N_A_M1034_g N_VGND_c_1242_n 0.00824727f $X=7.555 $Y=0.655 $X2=0 $Y2=0
cc_351 N_A_c_187_n N_VGND_c_1242_n 0.00605278f $X=3.505 $Y=1.185 $X2=0 $Y2=0
cc_352 N_A_M1008_g N_VGND_c_1246_n 0.0136172f $X=6.265 $Y=0.655 $X2=0 $Y2=0
cc_353 N_A_M1017_g N_VGND_c_1246_n 5.8953e-19 $X=6.695 $Y=0.655 $X2=0 $Y2=0
cc_354 N_A_c_181_n N_VGND_c_1246_n 0.0053631f $X=6.335 $Y=1.295 $X2=0 $Y2=0
cc_355 N_A_c_178_n N_A_110_47#_M1030_d 0.0015736f $X=1.407 $Y=1.16 $X2=0 $Y2=0
cc_356 N_A_c_177_n N_A_110_47#_M1033_s 7.50739e-19 $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_357 N_A_M1020_g N_A_110_47#_c_1393_n 2.2122e-19 $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_358 N_A_c_176_n N_A_110_47#_c_1393_n 0.0150652f $X=1.26 $Y=1.4 $X2=0 $Y2=0
cc_359 N_A_c_178_n N_A_110_47#_c_1393_n 6.7581e-19 $X=1.407 $Y=1.16 $X2=0 $Y2=0
cc_360 N_A_c_185_n N_A_110_47#_c_1393_n 0.00231808f $X=1.335 $Y=1.44 $X2=0 $Y2=0
cc_361 N_A_M1020_g N_A_110_47#_c_1400_n 0.0112498f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_362 N_A_M1030_g N_A_110_47#_c_1400_n 0.00873255f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_363 N_A_c_176_n N_A_110_47#_c_1400_n 0.0146728f $X=1.26 $Y=1.4 $X2=0 $Y2=0
cc_364 N_A_c_178_n N_A_110_47#_c_1400_n 0.0084836f $X=1.407 $Y=1.16 $X2=0 $Y2=0
cc_365 N_A_c_183_n N_A_110_47#_c_1400_n 6.67853e-19 $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_366 N_A_c_185_n N_A_110_47#_c_1400_n 0.00194014f $X=1.335 $Y=1.44 $X2=0 $Y2=0
cc_367 N_A_M1030_g N_A_110_47#_c_1406_n 0.00294618f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_368 N_A_M1020_g N_A_110_47#_c_1407_n 4.55047e-19 $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_369 N_A_M1030_g N_A_110_47#_c_1407_n 0.00417357f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_370 N_A_c_177_n N_A_110_47#_c_1407_n 0.00643428f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_371 N_A_c_178_n N_A_110_47#_c_1407_n 0.0113221f $X=1.407 $Y=1.16 $X2=0 $Y2=0
cc_372 N_A_c_183_n N_A_110_47#_c_1407_n 0.00160826f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_373 N_A_c_177_n N_A_110_47#_c_1412_n 0.004087f $X=3.34 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A_c_187_n N_A_110_47#_c_1412_n 0.00329243f $X=3.505 $Y=1.185 $X2=0
+ $Y2=0
cc_375 N_B_c_425_n N_A_776_255#_M1005_g 0.00569712f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_376 N_B_c_425_n N_A_776_255#_M1010_g 0.00419064f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_377 N_B_c_425_n N_A_776_255#_M1022_g 0.00441105f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_378 N_B_c_425_n N_A_776_255#_M1035_g 0.00911556f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_379 N_B_c_425_n N_A_776_255#_c_634_n 0.0334539f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_380 N_B_c_425_n N_A_776_255#_c_635_n 0.0093254f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_381 N_B_M1002_g N_A_776_255#_c_637_n 0.0134807f $X=7.985 $Y=0.655 $X2=0 $Y2=0
cc_382 N_B_c_423_n N_A_776_255#_c_637_n 0.00606602f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_383 N_B_c_425_n N_A_776_255#_c_637_n 0.00450496f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_384 B N_A_776_255#_c_637_n 0.00299608f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_385 N_B_c_428_n N_A_776_255#_c_637_n 0.0137551f $X=7.92 $Y=1.445 $X2=0 $Y2=0
cc_386 N_B_M1011_g N_A_776_255#_c_709_n 0.012262f $X=8.485 $Y=2.465 $X2=0 $Y2=0
cc_387 N_B_M1023_g N_A_776_255#_c_709_n 6.32357e-19 $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_388 N_B_M1015_g N_A_776_255#_c_638_n 0.0135734f $X=8.415 $Y=0.655 $X2=0 $Y2=0
cc_389 N_B_M1028_g N_A_776_255#_c_638_n 0.0135734f $X=8.845 $Y=0.655 $X2=0 $Y2=0
cc_390 N_B_c_423_n N_A_776_255#_c_638_n 0.0469271f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_391 N_B_c_424_n N_A_776_255#_c_638_n 0.00276559f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_392 N_B_M1011_g N_A_776_255#_c_649_n 0.01115f $X=8.485 $Y=2.465 $X2=0 $Y2=0
cc_393 N_B_M1023_g N_A_776_255#_c_649_n 0.0111034f $X=8.915 $Y=2.465 $X2=0 $Y2=0
cc_394 N_B_c_423_n N_A_776_255#_c_649_n 0.0370651f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_395 N_B_c_424_n N_A_776_255#_c_649_n 0.00273301f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_396 N_B_M1001_g N_A_776_255#_c_650_n 0.00184744f $X=8.055 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_B_M1011_g N_A_776_255#_c_650_n 0.00192937f $X=8.485 $Y=2.465 $X2=0
+ $Y2=0
cc_398 N_B_c_423_n N_A_776_255#_c_650_n 0.0201351f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_399 N_B_c_424_n N_A_776_255#_c_650_n 0.00283411f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_400 B N_A_776_255#_c_650_n 0.00219466f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_401 N_B_c_428_n N_A_776_255#_c_650_n 0.00685781f $X=7.92 $Y=1.445 $X2=0 $Y2=0
cc_402 N_B_M1011_g N_A_776_255#_c_725_n 6.30056e-19 $X=8.485 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_B_M1023_g N_A_776_255#_c_725_n 0.0102493f $X=8.915 $Y=2.465 $X2=0 $Y2=0
cc_404 N_B_M1038_g N_A_776_255#_c_725_n 0.0150032f $X=9.345 $Y=2.465 $X2=0 $Y2=0
cc_405 N_B_M1029_g N_A_776_255#_c_639_n 0.0155199f $X=9.275 $Y=0.655 $X2=0 $Y2=0
cc_406 N_B_c_423_n N_A_776_255#_c_639_n 0.0313612f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_407 N_B_c_424_n N_A_776_255#_c_639_n 0.00646267f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_408 N_B_M1038_g N_A_776_255#_c_651_n 0.0130252f $X=9.345 $Y=2.465 $X2=0 $Y2=0
cc_409 N_B_c_423_n N_A_776_255#_c_651_n 0.0214032f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_410 N_B_c_424_n N_A_776_255#_c_651_n 0.00438376f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_411 N_B_M1029_g N_A_776_255#_c_640_n 0.00241875f $X=9.275 $Y=0.655 $X2=0
+ $Y2=0
cc_412 N_B_M1038_g N_A_776_255#_c_640_n 0.00289347f $X=9.345 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_B_c_423_n N_A_776_255#_c_640_n 0.0145177f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_414 N_B_c_424_n N_A_776_255#_c_640_n 0.00774881f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_415 N_B_c_423_n N_A_776_255#_c_642_n 0.015388f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_416 N_B_c_424_n N_A_776_255#_c_642_n 0.00286879f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_417 N_B_c_423_n N_A_776_255#_c_643_n 0.015388f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_418 N_B_c_424_n N_A_776_255#_c_643_n 0.00286879f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_419 N_B_M1023_g N_A_776_255#_c_653_n 0.00229961f $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_420 N_B_M1038_g N_A_776_255#_c_653_n 0.00229961f $X=9.345 $Y=2.465 $X2=0
+ $Y2=0
cc_421 N_B_c_423_n N_A_776_255#_c_653_n 0.0265023f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_422 N_B_c_424_n N_A_776_255#_c_653_n 0.00283411f $X=9.435 $Y=1.44 $X2=0 $Y2=0
cc_423 N_B_c_425_n N_A_776_255#_c_644_n 0.0108357f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_424 N_B_M1003_g N_A_27_367#_c_860_n 0.0126616f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_425 N_B_c_440_n N_A_27_367#_c_860_n 0.0092301f $X=2.92 $Y=1.51 $X2=0 $Y2=0
cc_426 N_B_M1009_g N_A_27_367#_c_875_n 0.0122531f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_427 N_B_M1025_g N_A_27_367#_c_875_n 0.0121795f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_428 N_B_c_438_n N_A_27_367#_c_875_n 0.00625646f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_429 N_B_c_440_n N_A_27_367#_c_875_n 0.0401825f $X=2.92 $Y=1.51 $X2=0 $Y2=0
cc_430 N_B_c_427_n N_A_27_367#_c_875_n 5.45297e-19 $X=3.055 $Y=1.51 $X2=0 $Y2=0
cc_431 N_B_M1032_g N_A_27_367#_c_863_n 0.0129116f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_432 N_B_c_425_n N_A_27_367#_c_863_n 0.0190864f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_433 N_B_c_440_n N_A_27_367#_c_863_n 0.00817045f $X=2.92 $Y=1.51 $X2=0 $Y2=0
cc_434 N_B_c_425_n N_A_27_367#_c_866_n 0.00889582f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_435 N_B_c_425_n N_A_27_367#_c_854_n 0.00816414f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_436 N_B_c_440_n N_A_27_367#_c_855_n 0.00276363f $X=2.92 $Y=1.51 $X2=0 $Y2=0
cc_437 N_B_c_440_n N_A_27_367#_c_886_n 0.0151123f $X=2.92 $Y=1.51 $X2=0 $Y2=0
cc_438 N_B_c_427_n N_A_27_367#_c_886_n 6.16419e-19 $X=3.055 $Y=1.51 $X2=0 $Y2=0
cc_439 N_B_c_425_n N_A_27_367#_c_888_n 0.00128847f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_440 N_B_c_438_n N_A_27_367#_c_888_n 0.00114299f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_441 N_B_c_440_n N_A_27_367#_c_888_n 0.0145874f $X=2.92 $Y=1.51 $X2=0 $Y2=0
cc_442 N_B_c_427_n N_A_27_367#_c_888_n 6.16419e-19 $X=3.055 $Y=1.51 $X2=0 $Y2=0
cc_443 N_B_M1003_g N_VPWR_c_941_n 0.0142626f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_444 N_B_M1009_g N_VPWR_c_941_n 6.73419e-19 $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_445 N_B_M1003_g N_VPWR_c_942_n 6.73419e-19 $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_446 N_B_M1009_g N_VPWR_c_942_n 0.0143455f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_447 N_B_M1025_g N_VPWR_c_942_n 0.0143786f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_448 N_B_M1032_g N_VPWR_c_942_n 6.79552e-19 $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_449 N_B_M1025_g N_VPWR_c_943_n 0.00486043f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_450 N_B_M1032_g N_VPWR_c_943_n 0.00544582f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_451 N_B_M1025_g N_VPWR_c_944_n 6.54139e-19 $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_452 N_B_M1032_g N_VPWR_c_944_n 0.0133914f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_453 N_B_M1001_g N_VPWR_c_946_n 0.00109252f $X=8.055 $Y=2.465 $X2=0 $Y2=0
cc_454 N_B_M1003_g N_VPWR_c_949_n 0.00486043f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_455 N_B_M1009_g N_VPWR_c_949_n 0.00486043f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_456 N_B_M1001_g N_VPWR_c_954_n 0.00357877f $X=8.055 $Y=2.465 $X2=0 $Y2=0
cc_457 N_B_M1011_g N_VPWR_c_954_n 0.00357877f $X=8.485 $Y=2.465 $X2=0 $Y2=0
cc_458 N_B_M1023_g N_VPWR_c_954_n 0.00357877f $X=8.915 $Y=2.465 $X2=0 $Y2=0
cc_459 N_B_M1038_g N_VPWR_c_954_n 0.00357877f $X=9.345 $Y=2.465 $X2=0 $Y2=0
cc_460 N_B_M1003_g N_VPWR_c_939_n 0.00824727f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_461 N_B_M1009_g N_VPWR_c_939_n 0.00824727f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_462 N_B_M1025_g N_VPWR_c_939_n 0.00824727f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_463 N_B_M1032_g N_VPWR_c_939_n 0.009174f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_464 N_B_M1001_g N_VPWR_c_939_n 0.00537654f $X=8.055 $Y=2.465 $X2=0 $Y2=0
cc_465 N_B_M1011_g N_VPWR_c_939_n 0.0053512f $X=8.485 $Y=2.465 $X2=0 $Y2=0
cc_466 N_B_M1023_g N_VPWR_c_939_n 0.0053512f $X=8.915 $Y=2.465 $X2=0 $Y2=0
cc_467 N_B_M1038_g N_VPWR_c_939_n 0.00645423f $X=9.345 $Y=2.465 $X2=0 $Y2=0
cc_468 N_B_M1007_g N_X_c_1082_n 0.00276183f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_469 N_B_M1016_g N_X_c_1082_n 0.00946563f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_470 N_B_M1019_g N_X_c_1082_n 0.00946563f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_471 N_B_M1033_g N_X_c_1082_n 0.00940797f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_472 N_B_c_425_n N_X_c_1078_n 0.0324501f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_473 N_B_c_425_n N_X_c_1102_n 0.00995652f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_474 N_B_c_425_n N_X_c_1103_n 0.017827f $X=7.775 $Y=1.665 $X2=0 $Y2=0
cc_475 N_B_c_425_n N_A_1199_367#_c_1165_n 0.0178672f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_476 N_B_c_425_n N_A_1199_367#_c_1162_n 0.00912651f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_477 N_B_c_425_n N_A_1199_367#_c_1170_n 0.0193276f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_478 B N_A_1199_367#_c_1170_n 0.00362863f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_479 N_B_c_428_n N_A_1199_367#_c_1170_n 0.00838371f $X=7.92 $Y=1.445 $X2=0
+ $Y2=0
cc_480 N_B_M1001_g N_A_1199_367#_c_1181_n 0.012237f $X=8.055 $Y=2.465 $X2=0
+ $Y2=0
cc_481 N_B_M1011_g N_A_1199_367#_c_1181_n 0.0114565f $X=8.485 $Y=2.465 $X2=0
+ $Y2=0
cc_482 N_B_M1023_g N_A_1199_367#_c_1183_n 0.0115031f $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_483 N_B_M1038_g N_A_1199_367#_c_1183_n 0.0115031f $X=9.345 $Y=2.465 $X2=0
+ $Y2=0
cc_484 N_B_c_425_n N_A_1199_367#_c_1174_n 0.00546674f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_485 N_B_M1002_g N_VGND_c_1228_n 0.0102423f $X=7.985 $Y=0.655 $X2=0 $Y2=0
cc_486 N_B_M1015_g N_VGND_c_1228_n 6.16837e-19 $X=8.415 $Y=0.655 $X2=0 $Y2=0
cc_487 N_B_M1002_g N_VGND_c_1229_n 6.16837e-19 $X=7.985 $Y=0.655 $X2=0 $Y2=0
cc_488 N_B_M1015_g N_VGND_c_1229_n 0.010278f $X=8.415 $Y=0.655 $X2=0 $Y2=0
cc_489 N_B_M1028_g N_VGND_c_1229_n 0.010278f $X=8.845 $Y=0.655 $X2=0 $Y2=0
cc_490 N_B_M1029_g N_VGND_c_1229_n 6.16837e-19 $X=9.275 $Y=0.655 $X2=0 $Y2=0
cc_491 N_B_M1028_g N_VGND_c_1230_n 0.00486043f $X=8.845 $Y=0.655 $X2=0 $Y2=0
cc_492 N_B_M1029_g N_VGND_c_1230_n 0.00486043f $X=9.275 $Y=0.655 $X2=0 $Y2=0
cc_493 N_B_M1028_g N_VGND_c_1231_n 6.16837e-19 $X=8.845 $Y=0.655 $X2=0 $Y2=0
cc_494 N_B_M1029_g N_VGND_c_1231_n 0.0113415f $X=9.275 $Y=0.655 $X2=0 $Y2=0
cc_495 N_B_M1007_g N_VGND_c_1232_n 0.00357877f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_496 N_B_M1016_g N_VGND_c_1232_n 0.00357877f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_497 N_B_M1019_g N_VGND_c_1232_n 0.00357877f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_498 N_B_M1033_g N_VGND_c_1232_n 0.00357877f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_499 N_B_M1002_g N_VGND_c_1236_n 0.00486043f $X=7.985 $Y=0.655 $X2=0 $Y2=0
cc_500 N_B_M1015_g N_VGND_c_1236_n 0.00486043f $X=8.415 $Y=0.655 $X2=0 $Y2=0
cc_501 N_B_M1007_g N_VGND_c_1242_n 0.00537654f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_502 N_B_M1016_g N_VGND_c_1242_n 0.0053512f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_503 N_B_M1019_g N_VGND_c_1242_n 0.0053512f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_504 N_B_M1033_g N_VGND_c_1242_n 0.00537654f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_505 N_B_M1002_g N_VGND_c_1242_n 0.00824727f $X=7.985 $Y=0.655 $X2=0 $Y2=0
cc_506 N_B_M1015_g N_VGND_c_1242_n 0.00824727f $X=8.415 $Y=0.655 $X2=0 $Y2=0
cc_507 N_B_M1028_g N_VGND_c_1242_n 0.00824727f $X=8.845 $Y=0.655 $X2=0 $Y2=0
cc_508 N_B_M1029_g N_VGND_c_1242_n 0.00824727f $X=9.275 $Y=0.655 $X2=0 $Y2=0
cc_509 N_B_M1007_g N_A_110_47#_c_1412_n 0.0118957f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_510 N_B_M1016_g N_A_110_47#_c_1412_n 0.0103254f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_511 N_B_M1019_g N_A_110_47#_c_1412_n 0.0103254f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_512 N_B_M1033_g N_A_110_47#_c_1412_n 0.0103254f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_513 N_A_776_255#_M1005_g N_A_27_367#_c_892_n 0.0148836f $X=3.955 $Y=2.465
+ $X2=0 $Y2=0
cc_514 N_A_776_255#_M1010_g N_A_27_367#_c_892_n 0.0110316f $X=4.385 $Y=2.465
+ $X2=0 $Y2=0
cc_515 N_A_776_255#_M1022_g N_A_27_367#_c_892_n 0.0111131f $X=4.815 $Y=2.465
+ $X2=0 $Y2=0
cc_516 N_A_776_255#_M1035_g N_A_27_367#_c_892_n 0.01523f $X=5.245 $Y=2.465 $X2=0
+ $Y2=0
cc_517 N_A_776_255#_M1035_g N_A_27_367#_c_854_n 0.00448354f $X=5.245 $Y=2.465
+ $X2=0 $Y2=0
cc_518 N_A_776_255#_c_634_n N_A_27_367#_c_854_n 0.00873746f $X=5.825 $Y=1.445
+ $X2=0 $Y2=0
cc_519 N_A_776_255#_c_635_n N_A_27_367#_c_854_n 0.00471729f $X=5.74 $Y=1.44
+ $X2=0 $Y2=0
cc_520 N_A_776_255#_M1005_g N_VPWR_c_944_n 0.00104719f $X=3.955 $Y=2.465 $X2=0
+ $Y2=0
cc_521 N_A_776_255#_M1005_g N_VPWR_c_952_n 0.00357877f $X=3.955 $Y=2.465 $X2=0
+ $Y2=0
cc_522 N_A_776_255#_M1010_g N_VPWR_c_952_n 0.00357877f $X=4.385 $Y=2.465 $X2=0
+ $Y2=0
cc_523 N_A_776_255#_M1022_g N_VPWR_c_952_n 0.00357877f $X=4.815 $Y=2.465 $X2=0
+ $Y2=0
cc_524 N_A_776_255#_M1035_g N_VPWR_c_952_n 0.00357877f $X=5.245 $Y=2.465 $X2=0
+ $Y2=0
cc_525 N_A_776_255#_M1001_d N_VPWR_c_939_n 0.00225186f $X=8.13 $Y=1.835 $X2=0
+ $Y2=0
cc_526 N_A_776_255#_M1023_d N_VPWR_c_939_n 0.00225186f $X=8.99 $Y=1.835 $X2=0
+ $Y2=0
cc_527 N_A_776_255#_M1005_g N_VPWR_c_939_n 0.0054006f $X=3.955 $Y=2.465 $X2=0
+ $Y2=0
cc_528 N_A_776_255#_M1010_g N_VPWR_c_939_n 0.0053512f $X=4.385 $Y=2.465 $X2=0
+ $Y2=0
cc_529 N_A_776_255#_M1022_g N_VPWR_c_939_n 0.0053512f $X=4.815 $Y=2.465 $X2=0
+ $Y2=0
cc_530 N_A_776_255#_M1035_g N_VPWR_c_939_n 0.00665089f $X=5.245 $Y=2.465 $X2=0
+ $Y2=0
cc_531 N_A_776_255#_M1013_g N_X_c_1082_n 0.00874807f $X=3.985 $Y=0.655 $X2=0
+ $Y2=0
cc_532 N_A_776_255#_M1005_g N_X_c_1105_n 0.00389289f $X=3.955 $Y=2.465 $X2=0
+ $Y2=0
cc_533 N_A_776_255#_M1005_g N_X_c_1078_n 0.0135226f $X=3.955 $Y=2.465 $X2=0
+ $Y2=0
cc_534 N_A_776_255#_M1013_g N_X_c_1078_n 0.0019661f $X=3.985 $Y=0.655 $X2=0
+ $Y2=0
cc_535 N_A_776_255#_M1010_g N_X_c_1078_n 0.00595244f $X=4.385 $Y=2.465 $X2=0
+ $Y2=0
cc_536 N_A_776_255#_M1024_g N_X_c_1078_n 0.00206138f $X=4.415 $Y=0.655 $X2=0
+ $Y2=0
cc_537 N_A_776_255#_c_634_n N_X_c_1078_n 0.0139245f $X=5.825 $Y=1.445 $X2=0
+ $Y2=0
cc_538 N_A_776_255#_c_644_n N_X_c_1078_n 0.0250141f $X=5.35 $Y=1.44 $X2=0 $Y2=0
cc_539 N_A_776_255#_M1024_g N_X_c_1079_n 0.0127308f $X=4.415 $Y=0.655 $X2=0
+ $Y2=0
cc_540 N_A_776_255#_M1026_g N_X_c_1079_n 0.0131284f $X=4.845 $Y=0.655 $X2=0
+ $Y2=0
cc_541 N_A_776_255#_M1031_g N_X_c_1079_n 0.00159113f $X=5.275 $Y=0.655 $X2=0
+ $Y2=0
cc_542 N_A_776_255#_c_634_n N_X_c_1079_n 0.0445847f $X=5.825 $Y=1.445 $X2=0
+ $Y2=0
cc_543 N_A_776_255#_c_636_n N_X_c_1079_n 0.00265947f $X=5.98 $Y=1.355 $X2=0
+ $Y2=0
cc_544 N_A_776_255#_c_644_n N_X_c_1079_n 0.00413685f $X=5.35 $Y=1.44 $X2=0 $Y2=0
cc_545 N_A_776_255#_M1022_g N_X_c_1118_n 0.00123811f $X=4.815 $Y=2.465 $X2=0
+ $Y2=0
cc_546 N_A_776_255#_M1035_g N_X_c_1118_n 0.00389531f $X=5.245 $Y=2.465 $X2=0
+ $Y2=0
cc_547 N_A_776_255#_M1010_g N_X_c_1102_n 0.00134152f $X=4.385 $Y=2.465 $X2=0
+ $Y2=0
cc_548 N_A_776_255#_M1022_g N_X_c_1102_n 0.0102121f $X=4.815 $Y=2.465 $X2=0
+ $Y2=0
cc_549 N_A_776_255#_M1035_g N_X_c_1102_n 0.00677322f $X=5.245 $Y=2.465 $X2=0
+ $Y2=0
cc_550 N_A_776_255#_c_634_n N_X_c_1102_n 0.00739597f $X=5.825 $Y=1.445 $X2=0
+ $Y2=0
cc_551 N_A_776_255#_c_644_n N_X_c_1102_n 0.00181199f $X=5.35 $Y=1.44 $X2=0 $Y2=0
cc_552 N_A_776_255#_M1013_g N_X_c_1080_n 0.01036f $X=3.985 $Y=0.655 $X2=0 $Y2=0
cc_553 N_A_776_255#_M1024_g N_X_c_1080_n 2.39785e-19 $X=4.415 $Y=0.655 $X2=0
+ $Y2=0
cc_554 N_A_776_255#_M1010_g N_X_c_1103_n 0.0139317f $X=4.385 $Y=2.465 $X2=0
+ $Y2=0
cc_555 N_A_776_255#_M1022_g N_X_c_1103_n 0.0122214f $X=4.815 $Y=2.465 $X2=0
+ $Y2=0
cc_556 N_A_776_255#_c_644_n N_X_c_1103_n 0.00179283f $X=5.35 $Y=1.44 $X2=0 $Y2=0
cc_557 N_A_776_255#_c_649_n N_A_1199_367#_M1011_s 0.00176461f $X=8.965 $Y=1.79
+ $X2=0 $Y2=0
cc_558 N_A_776_255#_c_651_n N_A_1199_367#_M1038_s 0.00239457f $X=9.77 $Y=1.79
+ $X2=0 $Y2=0
cc_559 N_A_776_255#_c_634_n N_A_1199_367#_c_1162_n 0.00406983f $X=5.825 $Y=1.445
+ $X2=0 $Y2=0
cc_560 N_A_776_255#_M1001_d N_A_1199_367#_c_1181_n 0.00332344f $X=8.13 $Y=1.835
+ $X2=0 $Y2=0
cc_561 N_A_776_255#_c_709_n N_A_1199_367#_c_1181_n 0.0143076f $X=8.27 $Y=1.96
+ $X2=0 $Y2=0
cc_562 N_A_776_255#_c_649_n N_A_1199_367#_c_1191_n 0.0135055f $X=8.965 $Y=1.79
+ $X2=0 $Y2=0
cc_563 N_A_776_255#_M1023_d N_A_1199_367#_c_1183_n 0.00332344f $X=8.99 $Y=1.835
+ $X2=0 $Y2=0
cc_564 N_A_776_255#_c_725_n N_A_1199_367#_c_1183_n 0.0159805f $X=9.13 $Y=1.96
+ $X2=0 $Y2=0
cc_565 N_A_776_255#_c_651_n N_A_1199_367#_c_1164_n 0.0202165f $X=9.77 $Y=1.79
+ $X2=0 $Y2=0
cc_566 N_A_776_255#_c_636_n N_VGND_M1031_d 8.69174e-19 $X=5.98 $Y=1.355 $X2=0
+ $Y2=0
cc_567 N_A_776_255#_c_801_p N_VGND_M1031_d 0.00677731f $X=6.135 $Y=0.945 $X2=0
+ $Y2=0
cc_568 N_A_776_255#_c_677_n N_VGND_M1017_s 0.00328191f $X=7.245 $Y=0.945 $X2=0
+ $Y2=0
cc_569 N_A_776_255#_c_637_n N_VGND_M1034_s 0.00176461f $X=8.105 $Y=1.1 $X2=0
+ $Y2=0
cc_570 N_A_776_255#_c_638_n N_VGND_M1015_d 0.00176461f $X=8.965 $Y=1.1 $X2=0
+ $Y2=0
cc_571 N_A_776_255#_c_639_n N_VGND_M1029_d 0.00248866f $X=9.77 $Y=1.1 $X2=0
+ $Y2=0
cc_572 N_A_776_255#_M1013_g N_VGND_c_1224_n 0.00705068f $X=3.985 $Y=0.655 $X2=0
+ $Y2=0
cc_573 N_A_776_255#_M1024_g N_VGND_c_1224_n 5.26307e-19 $X=4.415 $Y=0.655 $X2=0
+ $Y2=0
cc_574 N_A_776_255#_M1013_g N_VGND_c_1225_n 6.35001e-19 $X=3.985 $Y=0.655 $X2=0
+ $Y2=0
cc_575 N_A_776_255#_M1024_g N_VGND_c_1225_n 0.0102659f $X=4.415 $Y=0.655 $X2=0
+ $Y2=0
cc_576 N_A_776_255#_M1026_g N_VGND_c_1225_n 0.0102635f $X=4.845 $Y=0.655 $X2=0
+ $Y2=0
cc_577 N_A_776_255#_M1031_g N_VGND_c_1225_n 6.16426e-19 $X=5.275 $Y=0.655 $X2=0
+ $Y2=0
cc_578 N_A_776_255#_M1031_g N_VGND_c_1226_n 0.0063572f $X=5.275 $Y=0.655 $X2=0
+ $Y2=0
cc_579 N_A_776_255#_c_634_n N_VGND_c_1226_n 0.01403f $X=5.825 $Y=1.445 $X2=0
+ $Y2=0
cc_580 N_A_776_255#_c_635_n N_VGND_c_1226_n 0.0056629f $X=5.74 $Y=1.44 $X2=0
+ $Y2=0
cc_581 N_A_776_255#_c_636_n N_VGND_c_1226_n 0.00603927f $X=5.98 $Y=1.355 $X2=0
+ $Y2=0
cc_582 N_A_776_255#_c_801_p N_VGND_c_1226_n 0.0144778f $X=6.135 $Y=0.945 $X2=0
+ $Y2=0
cc_583 N_A_776_255#_c_677_n N_VGND_c_1227_n 0.0167297f $X=7.245 $Y=0.945 $X2=0
+ $Y2=0
cc_584 N_A_776_255#_c_637_n N_VGND_c_1228_n 0.0170777f $X=8.105 $Y=1.1 $X2=0
+ $Y2=0
cc_585 N_A_776_255#_c_638_n N_VGND_c_1229_n 0.0170777f $X=8.965 $Y=1.1 $X2=0
+ $Y2=0
cc_586 N_A_776_255#_c_820_p N_VGND_c_1230_n 0.0124525f $X=9.06 $Y=0.42 $X2=0
+ $Y2=0
cc_587 N_A_776_255#_c_639_n N_VGND_c_1231_n 0.0220026f $X=9.77 $Y=1.1 $X2=0
+ $Y2=0
cc_588 N_A_776_255#_c_822_p N_VGND_c_1234_n 0.0124525f $X=7.34 $Y=0.42 $X2=0
+ $Y2=0
cc_589 N_A_776_255#_c_823_p N_VGND_c_1236_n 0.0124525f $X=8.2 $Y=0.42 $X2=0
+ $Y2=0
cc_590 N_A_776_255#_M1013_g N_VGND_c_1239_n 0.00361616f $X=3.985 $Y=0.655 $X2=0
+ $Y2=0
cc_591 N_A_776_255#_M1024_g N_VGND_c_1239_n 0.00486043f $X=4.415 $Y=0.655 $X2=0
+ $Y2=0
cc_592 N_A_776_255#_c_826_p N_VGND_c_1240_n 0.0124525f $X=6.48 $Y=0.42 $X2=0
+ $Y2=0
cc_593 N_A_776_255#_M1008_d N_VGND_c_1242_n 0.00282948f $X=6.34 $Y=0.235 $X2=0
+ $Y2=0
cc_594 N_A_776_255#_M1018_d N_VGND_c_1242_n 0.00409797f $X=7.2 $Y=0.235 $X2=0
+ $Y2=0
cc_595 N_A_776_255#_M1002_s N_VGND_c_1242_n 0.00536646f $X=8.06 $Y=0.235 $X2=0
+ $Y2=0
cc_596 N_A_776_255#_M1028_s N_VGND_c_1242_n 0.00536646f $X=8.92 $Y=0.235 $X2=0
+ $Y2=0
cc_597 N_A_776_255#_M1013_g N_VGND_c_1242_n 0.00422438f $X=3.985 $Y=0.655 $X2=0
+ $Y2=0
cc_598 N_A_776_255#_M1024_g N_VGND_c_1242_n 0.00824727f $X=4.415 $Y=0.655 $X2=0
+ $Y2=0
cc_599 N_A_776_255#_M1026_g N_VGND_c_1242_n 0.00824727f $X=4.845 $Y=0.655 $X2=0
+ $Y2=0
cc_600 N_A_776_255#_M1031_g N_VGND_c_1242_n 0.00819843f $X=5.275 $Y=0.655 $X2=0
+ $Y2=0
cc_601 N_A_776_255#_c_673_n N_VGND_c_1242_n 0.00504665f $X=6.385 $Y=0.945 $X2=0
+ $Y2=0
cc_602 N_A_776_255#_c_801_p N_VGND_c_1242_n 0.00109435f $X=6.135 $Y=0.945 $X2=0
+ $Y2=0
cc_603 N_A_776_255#_c_826_p N_VGND_c_1242_n 0.00730901f $X=6.48 $Y=0.42 $X2=0
+ $Y2=0
cc_604 N_A_776_255#_c_677_n N_VGND_c_1242_n 0.0106723f $X=7.245 $Y=0.945 $X2=0
+ $Y2=0
cc_605 N_A_776_255#_c_822_p N_VGND_c_1242_n 0.00730901f $X=7.34 $Y=0.42 $X2=0
+ $Y2=0
cc_606 N_A_776_255#_c_823_p N_VGND_c_1242_n 0.00730901f $X=8.2 $Y=0.42 $X2=0
+ $Y2=0
cc_607 N_A_776_255#_c_820_p N_VGND_c_1242_n 0.00730901f $X=9.06 $Y=0.42 $X2=0
+ $Y2=0
cc_608 N_A_776_255#_M1026_g N_VGND_c_1245_n 0.00486043f $X=4.845 $Y=0.655 $X2=0
+ $Y2=0
cc_609 N_A_776_255#_M1031_g N_VGND_c_1245_n 0.00486043f $X=5.275 $Y=0.655 $X2=0
+ $Y2=0
cc_610 N_A_776_255#_M1026_g N_VGND_c_1246_n 5.8953e-19 $X=4.845 $Y=0.655 $X2=0
+ $Y2=0
cc_611 N_A_776_255#_M1031_g N_VGND_c_1246_n 0.0128133f $X=5.275 $Y=0.655 $X2=0
+ $Y2=0
cc_612 N_A_776_255#_c_634_n N_VGND_c_1246_n 0.00212874f $X=5.825 $Y=1.445 $X2=0
+ $Y2=0
cc_613 N_A_776_255#_c_635_n N_VGND_c_1246_n 0.00233628f $X=5.74 $Y=1.44 $X2=0
+ $Y2=0
cc_614 N_A_776_255#_c_673_n N_VGND_c_1246_n 0.00175175f $X=6.385 $Y=0.945 $X2=0
+ $Y2=0
cc_615 N_A_776_255#_c_801_p N_VGND_c_1246_n 0.0261577f $X=6.135 $Y=0.945 $X2=0
+ $Y2=0
cc_616 N_A_27_367#_c_851_n N_VPWR_M1000_d 0.00176461f $X=1.025 $Y=1.78 $X2=-0.19
+ $Y2=1.655
cc_617 N_A_27_367#_c_860_n N_VPWR_M1014_d 0.00464713f $X=1.885 $Y=2.03 $X2=0
+ $Y2=0
cc_618 N_A_27_367#_c_875_n N_VPWR_M1009_d 0.00331377f $X=2.745 $Y=2.03 $X2=0
+ $Y2=0
cc_619 N_A_27_367#_c_863_n N_VPWR_M1032_d 0.00468694f $X=3.625 $Y=2.03 $X2=0
+ $Y2=0
cc_620 N_A_27_367#_c_851_n N_VPWR_c_940_n 0.0170777f $X=1.025 $Y=1.78 $X2=0
+ $Y2=0
cc_621 N_A_27_367#_c_860_n N_VPWR_c_941_n 0.0170777f $X=1.885 $Y=2.03 $X2=0
+ $Y2=0
cc_622 N_A_27_367#_c_875_n N_VPWR_c_942_n 0.0170111f $X=2.745 $Y=2.03 $X2=0
+ $Y2=0
cc_623 N_A_27_367#_c_906_p N_VPWR_c_943_n 0.0129847f $X=2.84 $Y=2.48 $X2=0 $Y2=0
cc_624 N_A_27_367#_c_863_n N_VPWR_c_944_n 0.0166824f $X=3.625 $Y=2.03 $X2=0
+ $Y2=0
cc_625 N_A_27_367#_c_908_p N_VPWR_c_947_n 0.0124525f $X=1.12 $Y=2.44 $X2=0 $Y2=0
cc_626 N_A_27_367#_c_909_p N_VPWR_c_949_n 0.0124525f $X=1.98 $Y=2.48 $X2=0 $Y2=0
cc_627 N_A_27_367#_c_850_n N_VPWR_c_951_n 0.0178111f $X=0.26 $Y=1.98 $X2=0 $Y2=0
cc_628 N_A_27_367#_c_911_p N_VPWR_c_952_n 0.0132266f $X=3.725 $Y=2.775 $X2=0
+ $Y2=0
cc_629 N_A_27_367#_c_892_n N_VPWR_c_952_n 0.0866227f $X=5.365 $Y=2.925 $X2=0
+ $Y2=0
cc_630 N_A_27_367#_c_853_n N_VPWR_c_952_n 0.0179183f $X=5.495 $Y=2.775 $X2=0
+ $Y2=0
cc_631 N_A_27_367#_M1000_s N_VPWR_c_939_n 0.00371702f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_632 N_A_27_367#_M1004_s N_VPWR_c_939_n 0.00536646f $X=0.98 $Y=1.835 $X2=0
+ $Y2=0
cc_633 N_A_27_367#_M1003_s N_VPWR_c_939_n 0.00536646f $X=1.84 $Y=1.835 $X2=0
+ $Y2=0
cc_634 N_A_27_367#_M1025_s N_VPWR_c_939_n 0.00484465f $X=2.7 $Y=1.835 $X2=0
+ $Y2=0
cc_635 N_A_27_367#_M1037_s N_VPWR_c_939_n 0.00349882f $X=3.59 $Y=1.835 $X2=0
+ $Y2=0
cc_636 N_A_27_367#_M1010_d N_VPWR_c_939_n 0.00223577f $X=4.46 $Y=1.835 $X2=0
+ $Y2=0
cc_637 N_A_27_367#_M1035_d N_VPWR_c_939_n 0.00215161f $X=5.32 $Y=1.835 $X2=0
+ $Y2=0
cc_638 N_A_27_367#_c_850_n N_VPWR_c_939_n 0.0100304f $X=0.26 $Y=1.98 $X2=0 $Y2=0
cc_639 N_A_27_367#_c_908_p N_VPWR_c_939_n 0.00730901f $X=1.12 $Y=2.44 $X2=0
+ $Y2=0
cc_640 N_A_27_367#_c_909_p N_VPWR_c_939_n 0.00730901f $X=1.98 $Y=2.48 $X2=0
+ $Y2=0
cc_641 N_A_27_367#_c_906_p N_VPWR_c_939_n 0.00789217f $X=2.84 $Y=2.48 $X2=0
+ $Y2=0
cc_642 N_A_27_367#_c_911_p N_VPWR_c_939_n 0.00776497f $X=3.725 $Y=2.775 $X2=0
+ $Y2=0
cc_643 N_A_27_367#_c_892_n N_VPWR_c_939_n 0.055599f $X=5.365 $Y=2.925 $X2=0
+ $Y2=0
cc_644 N_A_27_367#_c_853_n N_VPWR_c_939_n 0.0101029f $X=5.495 $Y=2.775 $X2=0
+ $Y2=0
cc_645 N_A_27_367#_c_892_n N_X_M1005_s 0.00338208f $X=5.365 $Y=2.925 $X2=0 $Y2=0
cc_646 N_A_27_367#_c_892_n N_X_M1022_s 0.00338208f $X=5.365 $Y=2.925 $X2=0 $Y2=0
cc_647 N_A_27_367#_c_892_n N_X_c_1105_n 0.0160685f $X=5.365 $Y=2.925 $X2=0 $Y2=0
cc_648 N_A_27_367#_c_892_n N_X_c_1118_n 0.0172102f $X=5.365 $Y=2.925 $X2=0 $Y2=0
cc_649 N_A_27_367#_M1010_d N_X_c_1103_n 0.00412038f $X=4.46 $Y=1.835 $X2=0 $Y2=0
cc_650 N_A_27_367#_c_892_n N_X_c_1103_n 0.0321645f $X=5.365 $Y=2.925 $X2=0 $Y2=0
cc_651 N_A_27_367#_c_853_n N_A_1199_367#_c_1161_n 0.0164532f $X=5.495 $Y=2.775
+ $X2=0 $Y2=0
cc_652 N_A_27_367#_c_854_n N_A_1199_367#_c_1161_n 0.0321754f $X=5.46 $Y=1.98
+ $X2=0 $Y2=0
cc_653 N_A_27_367#_c_854_n N_A_1199_367#_c_1162_n 0.0093235f $X=5.46 $Y=1.98
+ $X2=0 $Y2=0
cc_654 N_A_27_367#_c_851_n N_VGND_c_1222_n 0.00156123f $X=1.025 $Y=1.78 $X2=0
+ $Y2=0
cc_655 N_A_27_367#_c_852_n N_VGND_c_1222_n 0.0100387f $X=0.355 $Y=1.78 $X2=0
+ $Y2=0
cc_656 N_VPWR_c_939_n N_X_M1005_s 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_657 N_VPWR_c_939_n N_X_M1022_s 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_658 N_VPWR_c_939_n N_A_1199_367#_M1006_s 0.00371702f $X=9.84 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_659 N_VPWR_c_939_n N_A_1199_367#_M1021_s 0.00536646f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_660 N_VPWR_c_939_n N_A_1199_367#_M1036_s 0.00376627f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_661 N_VPWR_c_939_n N_A_1199_367#_M1011_s 0.00223565f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_662 N_VPWR_c_939_n N_A_1199_367#_M1038_s 0.00215161f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_952_n N_A_1199_367#_c_1161_n 0.0178111f $X=6.385 $Y=3.33 $X2=0
+ $Y2=0
cc_664 N_VPWR_c_939_n N_A_1199_367#_c_1161_n 0.0100304f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_665 N_VPWR_M1006_d N_A_1199_367#_c_1165_n 0.00393074f $X=6.41 $Y=1.835 $X2=0
+ $Y2=0
cc_666 N_VPWR_c_945_n N_A_1199_367#_c_1165_n 0.0165807f $X=6.55 $Y=2.415 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_953_n N_A_1199_367#_c_1207_n 0.0124525f $X=7.245 $Y=3.33 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_939_n N_A_1199_367#_c_1207_n 0.00730901f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_669 N_VPWR_M1027_d N_A_1199_367#_c_1170_n 0.00393074f $X=7.27 $Y=1.835 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_946_n N_A_1199_367#_c_1170_n 0.0165807f $X=7.41 $Y=2.415 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_954_n N_A_1199_367#_c_1211_n 0.0125234f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_672 N_VPWR_c_939_n N_A_1199_367#_c_1211_n 0.00738676f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_954_n N_A_1199_367#_c_1181_n 0.0361172f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_674 N_VPWR_c_939_n N_A_1199_367#_c_1181_n 0.023676f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_675 N_VPWR_c_954_n N_A_1199_367#_c_1183_n 0.0361172f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_939_n N_A_1199_367#_c_1183_n 0.023676f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_677 N_VPWR_c_954_n N_A_1199_367#_c_1163_n 0.0179183f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_678 N_VPWR_c_939_n N_A_1199_367#_c_1163_n 0.0101082f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_679 N_VPWR_c_954_n N_A_1199_367#_c_1219_n 0.0125234f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_680 N_VPWR_c_939_n N_A_1199_367#_c_1219_n 0.00738676f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_681 N_X_c_1082_n N_VGND_M1039_s 0.00562262f $X=3.995 $Y=0.8 $X2=0 $Y2=0
cc_682 N_X_c_1079_n N_VGND_M1024_d 0.00176461f $X=4.965 $Y=1.1 $X2=0 $Y2=0
cc_683 N_X_c_1082_n N_VGND_c_1224_n 0.0202946f $X=3.995 $Y=0.8 $X2=0 $Y2=0
cc_684 N_X_c_1079_n N_VGND_c_1225_n 0.0160814f $X=4.965 $Y=1.1 $X2=0 $Y2=0
cc_685 N_X_c_1079_n N_VGND_c_1226_n 0.00474502f $X=4.965 $Y=1.1 $X2=0 $Y2=0
cc_686 N_X_c_1082_n N_VGND_c_1232_n 0.00217533f $X=3.995 $Y=0.8 $X2=0 $Y2=0
cc_687 N_X_c_1082_n N_VGND_c_1239_n 8.58939e-19 $X=3.995 $Y=0.8 $X2=0 $Y2=0
cc_688 N_X_c_1145_p N_VGND_c_1239_n 0.0124525f $X=4.2 $Y=0.42 $X2=0 $Y2=0
cc_689 N_X_c_1080_n N_VGND_c_1239_n 0.00138195f $X=4.145 $Y=0.8 $X2=0 $Y2=0
cc_690 N_X_M1007_d N_VGND_c_1242_n 0.00225186f $X=1.84 $Y=0.235 $X2=0 $Y2=0
cc_691 N_X_M1019_d N_VGND_c_1242_n 0.00225186f $X=2.7 $Y=0.235 $X2=0 $Y2=0
cc_692 N_X_M1013_s N_VGND_c_1242_n 0.00398877f $X=4.06 $Y=0.235 $X2=0 $Y2=0
cc_693 N_X_M1026_s N_VGND_c_1242_n 0.00536646f $X=4.92 $Y=0.235 $X2=0 $Y2=0
cc_694 N_X_c_1082_n N_VGND_c_1242_n 0.00957098f $X=3.995 $Y=0.8 $X2=0 $Y2=0
cc_695 N_X_c_1145_p N_VGND_c_1242_n 0.00730901f $X=4.2 $Y=0.42 $X2=0 $Y2=0
cc_696 N_X_c_1153_p N_VGND_c_1242_n 0.00730901f $X=5.06 $Y=0.42 $X2=0 $Y2=0
cc_697 N_X_c_1080_n N_VGND_c_1242_n 0.00278726f $X=4.145 $Y=0.8 $X2=0 $Y2=0
cc_698 N_X_c_1153_p N_VGND_c_1245_n 0.0124525f $X=5.06 $Y=0.42 $X2=0 $Y2=0
cc_699 N_X_c_1082_n N_A_110_47#_M1016_s 0.00328308f $X=3.995 $Y=0.8 $X2=0 $Y2=0
cc_700 N_X_c_1082_n N_A_110_47#_M1033_s 0.00338154f $X=3.995 $Y=0.8 $X2=0 $Y2=0
cc_701 N_X_M1007_d N_A_110_47#_c_1412_n 0.00337551f $X=1.84 $Y=0.235 $X2=0 $Y2=0
cc_702 N_X_M1019_d N_A_110_47#_c_1412_n 0.00337551f $X=2.7 $Y=0.235 $X2=0 $Y2=0
cc_703 N_X_c_1082_n N_A_110_47#_c_1412_n 0.0825734f $X=3.995 $Y=0.8 $X2=0 $Y2=0
cc_704 N_VGND_c_1242_n N_A_110_47#_M1012_d 0.00386382f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_705 N_VGND_c_1242_n N_A_110_47#_M1030_d 0.00223562f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_706 N_VGND_c_1242_n N_A_110_47#_M1016_s 0.00223577f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_707 N_VGND_c_1242_n N_A_110_47#_M1033_s 0.00223577f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_708 N_VGND_c_1222_n N_A_110_47#_c_1393_n 0.0143034f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_709 N_VGND_c_1238_n N_A_110_47#_c_1428_n 0.0135169f $X=0.985 $Y=0 $X2=0 $Y2=0
cc_710 N_VGND_c_1242_n N_A_110_47#_c_1428_n 0.008474f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_711 N_VGND_M1020_s N_A_110_47#_c_1400_n 0.00399804f $X=0.98 $Y=0.235 $X2=0
+ $Y2=0
cc_712 N_VGND_c_1223_n N_A_110_47#_c_1400_n 0.0130182f $X=1.12 $Y=0.4 $X2=0
+ $Y2=0
cc_713 N_VGND_c_1232_n N_A_110_47#_c_1400_n 0.00196209f $X=3.605 $Y=0 $X2=0
+ $Y2=0
cc_714 N_VGND_c_1238_n N_A_110_47#_c_1400_n 0.00210007f $X=0.985 $Y=0 $X2=0
+ $Y2=0
cc_715 N_VGND_c_1242_n N_A_110_47#_c_1400_n 0.00833451f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_716 N_VGND_c_1232_n N_A_110_47#_c_1406_n 0.0157478f $X=3.605 $Y=0 $X2=0 $Y2=0
cc_717 N_VGND_c_1242_n N_A_110_47#_c_1406_n 0.00990873f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_718 N_VGND_c_1232_n N_A_110_47#_c_1412_n 0.100607f $X=3.605 $Y=0 $X2=0 $Y2=0
cc_719 N_VGND_c_1242_n N_A_110_47#_c_1412_n 0.0647738f $X=9.84 $Y=0 $X2=0 $Y2=0
