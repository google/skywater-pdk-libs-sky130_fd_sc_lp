* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4_lp A B C D VGND VNB VPB VPWR Y
X0 a_454_57# B Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 Y A a_612_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND C a_138_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 Y D a_296_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_409# C a_134_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_570_409# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_134_409# B a_570_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_612_57# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_296_57# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND B a_454_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 Y D a_27_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_138_57# C Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
