* File: sky130_fd_sc_lp__bufkapwr_4.pxi.spice
* Created: Wed Sep  2 09:36:08 2020
* 
x_PM_SKY130_FD_SC_LP__BUFKAPWR_4%A N_A_M1004_g N_A_M1009_g A N_A_c_51_n
+ N_A_c_52_n PM_SKY130_FD_SC_LP__BUFKAPWR_4%A
x_PM_SKY130_FD_SC_LP__BUFKAPWR_4%A_27_47# N_A_27_47#_M1004_s N_A_27_47#_M1009_s
+ N_A_27_47#_M1000_g N_A_27_47#_M1001_g N_A_27_47#_M1003_g N_A_27_47#_M1002_g
+ N_A_27_47#_M1006_g N_A_27_47#_M1005_g N_A_27_47#_M1008_g N_A_27_47#_M1007_g
+ N_A_27_47#_c_90_n N_A_27_47#_c_91_n N_A_27_47#_c_110_n N_A_27_47#_c_130_p
+ N_A_27_47#_c_92_n N_A_27_47#_c_93_n N_A_27_47#_c_94_n N_A_27_47#_c_95_n
+ PM_SKY130_FD_SC_LP__BUFKAPWR_4%A_27_47#
x_PM_SKY130_FD_SC_LP__BUFKAPWR_4%KAPWR N_KAPWR_M1009_d N_KAPWR_M1003_d
+ N_KAPWR_M1008_d KAPWR N_KAPWR_c_186_n N_KAPWR_c_199_p N_KAPWR_c_204_p
+ N_KAPWR_c_185_n KAPWR PM_SKY130_FD_SC_LP__BUFKAPWR_4%KAPWR
x_PM_SKY130_FD_SC_LP__BUFKAPWR_4%X N_X_M1001_d N_X_M1005_d N_X_M1000_s
+ N_X_M1006_s N_X_c_219_n N_X_c_232_n N_X_c_220_n N_X_c_221_n N_X_c_225_n
+ N_X_c_226_n N_X_c_222_n N_X_c_252_n X X X X PM_SKY130_FD_SC_LP__BUFKAPWR_4%X
x_PM_SKY130_FD_SC_LP__BUFKAPWR_4%VGND N_VGND_M1004_d N_VGND_M1002_s
+ N_VGND_M1007_s N_VGND_c_292_n N_VGND_c_293_n N_VGND_c_294_n N_VGND_c_295_n
+ N_VGND_c_296_n N_VGND_c_297_n VGND N_VGND_c_298_n N_VGND_c_299_n
+ N_VGND_c_300_n N_VGND_c_301_n PM_SKY130_FD_SC_LP__BUFKAPWR_4%VGND
x_PM_SKY130_FD_SC_LP__BUFKAPWR_4%VPWR VPWR N_VPWR_c_338_n VPWR
+ PM_SKY130_FD_SC_LP__BUFKAPWR_4%VPWR
cc_1 VNB N_A_M1009_g 0.0324163f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB A 0.00476547f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_3 VNB N_A_c_51_n 0.0314602f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.94
cc_4 VNB N_A_c_52_n 0.0206597f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.775
cc_5 VNB N_A_27_47#_M1000_g 0.00646593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_M1001_g 0.0391347f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.775
cc_7 VNB N_A_27_47#_M1003_g 0.00605191f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.94
cc_8 VNB N_A_27_47#_M1002_g 0.036407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1006_g 0.00604073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1005_g 0.0363926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1008_g 0.00738123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_M1007_g 0.0484726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_90_n 0.0313161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_91_n 0.00614616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_92_n 0.0132114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_93_n 0.0137262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_94_n 0.00875186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_95_n 0.0805965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_X_c_219_n 0.00246622f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.94
cc_20 VNB N_X_c_220_n 0.00543963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_221_n 0.00466661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_X_c_222_n 0.00276625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB X 0.0244059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB X 0.032052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_292_n 0.00475331f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.94
cc_26 VNB N_VGND_c_293_n 0.00404131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_294_n 0.0160143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_295_n 0.00474766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_296_n 0.0181274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_297_n 0.00487935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_298_n 0.0170407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_299_n 0.0168545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_300_n 0.00526407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_301_n 0.170308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB VPWR 0.123877f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.775
cc_36 VPB N_A_M1009_g 0.0240578f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_37 VPB N_A_27_47#_M1000_g 0.0207069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_M1003_g 0.0188623f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.94
cc_39 VPB N_A_27_47#_M1006_g 0.0188382f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_M1008_g 0.0239324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_91_n 0.0517803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_KAPWR_c_185_n 0.0298389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_X_c_225_n 0.0024786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_X_c_226_n 0.00359947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB X 0.0046916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB X 0.0187478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB VPWR 0.0439515f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.775
cc_48 VPB N_VPWR_c_338_n 0.0806132f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_49 N_A_M1009_g N_A_27_47#_M1001_g 0.00389195f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_50 A N_A_27_47#_M1001_g 0.00391122f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_51 N_A_c_51_n N_A_27_47#_M1001_g 0.0193356f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_52 N_A_c_52_n N_A_27_47#_M1001_g 0.0105633f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_53 N_A_M1009_g N_A_27_47#_c_90_n 0.00594476f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_54 A N_A_27_47#_c_90_n 0.025039f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_55 N_A_c_51_n N_A_27_47#_c_90_n 0.00816168f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_56 N_A_c_52_n N_A_27_47#_c_90_n 0.00544175f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_57 N_A_M1009_g N_A_27_47#_c_91_n 0.0138405f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_58 N_A_M1009_g N_A_27_47#_c_110_n 2.89127e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A_c_51_n N_A_27_47#_c_93_n 0.00165146f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_60 N_A_M1009_g N_A_27_47#_c_94_n 0.0222055f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_61 A N_A_27_47#_c_94_n 0.0295536f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_62 N_A_c_51_n N_A_27_47#_c_94_n 0.00300839f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_63 N_A_M1009_g N_A_27_47#_c_95_n 0.031642f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A_M1009_g N_KAPWR_c_186_n 7.52435e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_65 N_A_M1009_g N_KAPWR_c_185_n 0.00759753f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_66 A N_X_c_221_n 0.017502f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_67 A N_VGND_c_292_n 0.018208f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_68 N_A_c_51_n N_VGND_c_292_n 0.00261478f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_69 N_A_c_52_n N_VGND_c_292_n 0.00328447f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_70 N_A_c_51_n N_VGND_c_298_n 3.61504e-19 $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_71 N_A_c_52_n N_VGND_c_298_n 0.00585385f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_72 A N_VGND_c_301_n 0.00494628f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_73 N_A_c_51_n N_VGND_c_301_n 4.44682e-19 $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_74 N_A_c_52_n N_VGND_c_301_n 0.00798939f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_75 N_A_M1009_g VPWR 0.00642934f $X=0.475 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_76 N_A_M1009_g N_VPWR_c_338_n 0.00585385f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A_27_47#_M1000_g N_KAPWR_c_186_n 7.7142e-19 $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_78 N_A_27_47#_c_91_n N_KAPWR_c_186_n 0.00916602f $X=0.26 $Y=2.04 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_94_n N_KAPWR_c_186_n 0.013485f $X=1.075 $Y=1.37 $X2=0 $Y2=0
cc_80 N_A_27_47#_M1000_g N_KAPWR_c_185_n 0.00753148f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_81 N_A_27_47#_M1003_g N_KAPWR_c_185_n 0.00741597f $X=1.385 $Y=2.465 $X2=0
+ $Y2=0
cc_82 N_A_27_47#_M1006_g N_KAPWR_c_185_n 0.00741597f $X=1.815 $Y=2.465 $X2=0
+ $Y2=0
cc_83 N_A_27_47#_M1008_g N_KAPWR_c_185_n 0.00741597f $X=2.245 $Y=2.465 $X2=0
+ $Y2=0
cc_84 N_A_27_47#_c_91_n N_KAPWR_c_185_n 0.03569f $X=0.26 $Y=2.04 $X2=0 $Y2=0
cc_85 N_A_27_47#_M1001_g N_X_c_219_n 0.00333577f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A_27_47#_M1002_g N_X_c_219_n 0.00180205f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_27_47#_M1000_g N_X_c_232_n 6.92982e-19 $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_88 N_A_27_47#_M1003_g N_X_c_232_n 7.10691e-19 $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_27_47#_M1002_g N_X_c_220_n 0.0145209f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_90 N_A_27_47#_M1005_g N_X_c_220_n 0.0149582f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_130_p N_X_c_220_n 0.056586f $X=1.92 $Y=1.37 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_95_n N_X_c_220_n 0.00226821f $X=2.25 $Y=1.37 $X2=0 $Y2=0
cc_93 N_A_27_47#_M1001_g N_X_c_221_n 0.00262782f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_110_n N_X_c_221_n 0.0185462f $X=1.24 $Y=1.37 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_94_n N_X_c_221_n 0.00184173f $X=1.075 $Y=1.37 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_95_n N_X_c_221_n 0.00233759f $X=2.25 $Y=1.37 $X2=0 $Y2=0
cc_97 N_A_27_47#_M1003_g N_X_c_225_n 0.0143084f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_27_47#_M1006_g N_X_c_225_n 0.014515f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_130_p N_X_c_225_n 0.052712f $X=1.92 $Y=1.37 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_95_n N_X_c_225_n 0.00223239f $X=2.25 $Y=1.37 $X2=0 $Y2=0
cc_101 N_A_27_47#_M1000_g N_X_c_226_n 0.001967f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_91_n N_X_c_226_n 0.00367816f $X=0.26 $Y=2.04 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_94_n N_X_c_226_n 0.0200667f $X=1.075 $Y=1.37 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_95_n N_X_c_226_n 0.00232558f $X=2.25 $Y=1.37 $X2=0 $Y2=0
cc_105 N_A_27_47#_M1005_g N_X_c_222_n 0.00181183f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_27_47#_M1007_g N_X_c_222_n 0.00335855f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_27_47#_M1006_g N_X_c_252_n 7.02482e-19 $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_27_47#_M1008_g N_X_c_252_n 7.10691e-19 $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_27_47#_M1007_g X 0.0193193f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_95_n X 0.00226821f $X=2.25 $Y=1.37 $X2=0 $Y2=0
cc_111 N_A_27_47#_M1006_g X 9.88575e-19 $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_27_47#_M1005_g X 9.45451e-19 $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_27_47#_M1008_g X 0.00854578f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A_27_47#_M1007_g X 0.0081772f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_130_p X 0.0270337f $X=1.92 $Y=1.37 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_95_n X 0.0141672f $X=2.25 $Y=1.37 $X2=0 $Y2=0
cc_117 N_A_27_47#_M1008_g X 0.0180802f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_95_n X 0.0022548f $X=2.25 $Y=1.37 $X2=0 $Y2=0
cc_119 N_A_27_47#_M1001_g N_VGND_c_292_n 0.00163339f $X=0.96 $Y=0.445 $X2=0
+ $Y2=0
cc_120 N_A_27_47#_c_94_n N_VGND_c_292_n 7.37231e-19 $X=1.075 $Y=1.37 $X2=0 $Y2=0
cc_121 N_A_27_47#_M1002_g N_VGND_c_293_n 0.0017325f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_27_47#_M1005_g N_VGND_c_293_n 0.00165702f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_M1007_g N_VGND_c_295_n 0.00361578f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_M1001_g N_VGND_c_296_n 0.00585385f $X=0.96 $Y=0.445 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_M1002_g N_VGND_c_296_n 0.00585385f $X=1.39 $Y=0.445 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_c_92_n N_VGND_c_298_n 0.016561f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_127 N_A_27_47#_M1005_g N_VGND_c_299_n 0.00585385f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_128 N_A_27_47#_M1007_g N_VGND_c_299_n 0.00585385f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_M1004_s N_VGND_c_301_n 0.00232366f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_130 N_A_27_47#_M1001_g N_VGND_c_301_n 0.0109324f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_27_47#_M1002_g N_VGND_c_301_n 0.00609696f $X=1.39 $Y=0.445 $X2=0
+ $Y2=0
cc_132 N_A_27_47#_M1005_g N_VGND_c_301_n 0.00611063f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_M1007_g N_VGND_c_301_n 0.00722757f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_134 N_A_27_47#_c_92_n N_VGND_c_301_n 0.0113221f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_135 N_A_27_47#_M1009_s VPWR 0.0011275f $X=0.135 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_136 N_A_27_47#_M1000_g VPWR 0.00546086f $X=0.955 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_27_47#_M1003_g VPWR 0.00528318f $X=1.385 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_27_47#_M1006_g VPWR 0.00528318f $X=1.815 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_139 N_A_27_47#_M1008_g VPWR 0.00633597f $X=2.245 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_27_47#_c_91_n VPWR 0.00293051f $X=0.26 $Y=2.04 $X2=-0.19 $Y2=-0.245
cc_141 N_A_27_47#_M1000_g N_VPWR_c_338_n 0.00585385f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_M1003_g N_VPWR_c_338_n 0.00585385f $X=1.385 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_M1006_g N_VPWR_c_338_n 0.00585385f $X=1.815 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_M1008_g N_VPWR_c_338_n 0.00585385f $X=2.245 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_c_91_n N_VPWR_c_338_n 0.0182083f $X=0.26 $Y=2.04 $X2=0 $Y2=0
cc_146 N_KAPWR_c_185_n N_X_M1000_s 6.27314e-19 $X=2.475 $Y=2.81 $X2=0 $Y2=0
cc_147 N_KAPWR_c_185_n N_X_M1006_s 6.27314e-19 $X=2.475 $Y=2.81 $X2=0 $Y2=0
cc_148 N_KAPWR_c_186_n N_X_c_232_n 0.00914075f $X=0.69 $Y=2.04 $X2=0 $Y2=0
cc_149 N_KAPWR_c_199_p N_X_c_232_n 0.0091127f $X=1.6 $Y=2.23 $X2=0 $Y2=0
cc_150 N_KAPWR_c_185_n N_X_c_232_n 0.0289849f $X=2.475 $Y=2.81 $X2=0 $Y2=0
cc_151 N_KAPWR_M1003_d N_X_c_225_n 0.00176461f $X=1.46 $Y=1.835 $X2=0 $Y2=0
cc_152 N_KAPWR_c_199_p N_X_c_225_n 0.0135055f $X=1.6 $Y=2.23 $X2=0 $Y2=0
cc_153 N_KAPWR_c_199_p N_X_c_252_n 0.00885226f $X=1.6 $Y=2.23 $X2=0 $Y2=0
cc_154 N_KAPWR_c_204_p N_X_c_252_n 0.00912866f $X=2.46 $Y=2.23 $X2=0 $Y2=0
cc_155 N_KAPWR_c_185_n N_X_c_252_n 0.0290477f $X=2.475 $Y=2.81 $X2=0 $Y2=0
cc_156 N_KAPWR_M1008_d X 0.00296439f $X=2.32 $Y=1.835 $X2=0 $Y2=0
cc_157 N_KAPWR_c_204_p X 0.0196888f $X=2.46 $Y=2.23 $X2=0 $Y2=0
cc_158 N_KAPWR_M1009_d VPWR 0.00142085f $X=0.55 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_159 N_KAPWR_M1003_d VPWR 0.00123505f $X=1.46 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_160 N_KAPWR_M1008_d VPWR 0.00131667f $X=2.32 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_161 N_KAPWR_c_186_n VPWR 0.00293051f $X=0.69 $Y=2.04 $X2=-0.19 $Y2=1.655
cc_162 N_KAPWR_c_199_p VPWR 0.00237745f $X=1.6 $Y=2.23 $X2=-0.19 $Y2=1.655
cc_163 N_KAPWR_c_204_p VPWR 0.00265936f $X=2.46 $Y=2.23 $X2=-0.19 $Y2=1.655
cc_164 N_KAPWR_c_185_n VPWR 0.283742f $X=2.475 $Y=2.81 $X2=-0.19 $Y2=1.655
cc_165 N_KAPWR_c_186_n N_VPWR_c_338_n 0.0168497f $X=0.69 $Y=2.04 $X2=0 $Y2=0
cc_166 N_KAPWR_c_199_p N_VPWR_c_338_n 0.0147587f $X=1.6 $Y=2.23 $X2=0 $Y2=0
cc_167 N_KAPWR_c_204_p N_VPWR_c_338_n 0.0184704f $X=2.46 $Y=2.23 $X2=0 $Y2=0
cc_168 N_KAPWR_c_185_n N_VPWR_c_338_n 0.00654195f $X=2.475 $Y=2.81 $X2=0 $Y2=0
cc_169 N_X_c_220_n N_VGND_c_293_n 0.0169757f $X=1.905 $Y=0.9 $X2=0 $Y2=0
cc_170 X N_VGND_c_295_n 0.0208839f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_171 N_X_c_219_n N_VGND_c_296_n 0.0132609f $X=1.175 $Y=0.44 $X2=0 $Y2=0
cc_172 N_X_c_222_n N_VGND_c_299_n 0.0130349f $X=2.035 $Y=0.44 $X2=0 $Y2=0
cc_173 N_X_M1001_d N_VGND_c_301_n 0.00263279f $X=1.035 $Y=0.235 $X2=0 $Y2=0
cc_174 N_X_M1005_d N_VGND_c_301_n 0.0023552f $X=1.895 $Y=0.235 $X2=0 $Y2=0
cc_175 N_X_c_219_n N_VGND_c_301_n 0.00993371f $X=1.175 $Y=0.44 $X2=0 $Y2=0
cc_176 N_X_c_220_n N_VGND_c_301_n 0.016916f $X=1.905 $Y=0.9 $X2=0 $Y2=0
cc_177 N_X_c_222_n N_VGND_c_301_n 0.00984975f $X=2.035 $Y=0.44 $X2=0 $Y2=0
cc_178 X N_VGND_c_301_n 0.00671905f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_179 N_X_M1000_s VPWR 0.00121654f $X=1.03 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_180 N_X_M1006_s VPWR 0.00121654f $X=1.89 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_181 N_X_c_232_n VPWR 0.00245478f $X=1.17 $Y=2.04 $X2=-0.19 $Y2=-0.245
cc_182 N_X_c_252_n VPWR 0.00245478f $X=2.03 $Y=2.04 $X2=-0.19 $Y2=-0.245
cc_183 N_X_c_232_n N_VPWR_c_338_n 0.0136436f $X=1.17 $Y=2.04 $X2=0 $Y2=0
cc_184 N_X_c_252_n N_VPWR_c_338_n 0.0136436f $X=2.03 $Y=2.04 $X2=0 $Y2=0
