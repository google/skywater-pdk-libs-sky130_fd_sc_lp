* File: sky130_fd_sc_lp__nand4_0.pxi.spice
* Created: Fri Aug 28 10:50:31 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4_0%D N_D_M1004_g N_D_M1001_g N_D_c_62_n N_D_c_67_n D
+ D D D N_D_c_64_n PM_SKY130_FD_SC_LP__NAND4_0%D
x_PM_SKY130_FD_SC_LP__NAND4_0%C N_C_M1005_g N_C_M1006_g N_C_c_95_n N_C_c_96_n
+ N_C_c_97_n C C C C N_C_c_99_n PM_SKY130_FD_SC_LP__NAND4_0%C
x_PM_SKY130_FD_SC_LP__NAND4_0%B N_B_M1007_g N_B_M1003_g N_B_c_142_n N_B_c_143_n
+ N_B_c_144_n B B B B N_B_c_146_n PM_SKY130_FD_SC_LP__NAND4_0%B
x_PM_SKY130_FD_SC_LP__NAND4_0%A N_A_M1000_g N_A_M1002_g N_A_c_191_n N_A_c_198_n
+ N_A_c_192_n N_A_c_193_n A A A N_A_c_195_n PM_SKY130_FD_SC_LP__NAND4_0%A
x_PM_SKY130_FD_SC_LP__NAND4_0%VPWR N_VPWR_M1001_s N_VPWR_M1006_d N_VPWR_M1000_d
+ N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n
+ N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n VPWR
+ N_VPWR_c_243_n N_VPWR_c_233_n PM_SKY130_FD_SC_LP__NAND4_0%VPWR
x_PM_SKY130_FD_SC_LP__NAND4_0%Y N_Y_M1002_d N_Y_M1001_d N_Y_M1003_d N_Y_c_271_n
+ N_Y_c_272_n N_Y_c_273_n N_Y_c_269_n N_Y_c_275_n N_Y_c_276_n N_Y_c_270_n
+ N_Y_c_277_n Y Y Y PM_SKY130_FD_SC_LP__NAND4_0%Y
x_PM_SKY130_FD_SC_LP__NAND4_0%VGND N_VGND_M1004_s N_VGND_c_321_n N_VGND_c_322_n
+ N_VGND_c_323_n VGND N_VGND_c_324_n N_VGND_c_325_n
+ PM_SKY130_FD_SC_LP__NAND4_0%VGND
cc_1 VNB N_D_M1004_g 0.0466367f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.445
cc_2 VNB N_D_c_62_n 0.0285917f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_3 VNB D 0.0479844f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_4 VNB N_D_c_64_n 0.0185785f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_5 VNB N_C_M1006_g 0.0116035f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.63
cc_6 VNB N_C_c_95_n 0.0167706f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_7 VNB N_C_c_96_n 0.0238991f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.155
cc_8 VNB N_C_c_97_n 0.0167753f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.675
cc_9 VNB C 0.00241433f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_10 VNB N_C_c_99_n 0.0169494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_M1003_g 0.0101297f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.63
cc_12 VNB N_B_c_142_n 0.0176842f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_13 VNB N_B_c_143_n 0.021756f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.155
cc_14 VNB N_B_c_144_n 0.0160811f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.675
cc_15 VNB B 0.00885055f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_16 VNB N_B_c_146_n 0.0164392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_M1002_g 0.0251516f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.63
cc_18 VNB N_A_c_191_n 0.00886083f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.155
cc_19 VNB N_A_c_192_n 0.023629f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_20 VNB N_A_c_193_n 0.0172574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A 0.0109226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_c_195_n 0.016546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_233_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_269_n 0.0509824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_270_n 0.0170756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_321_n 0.0175269f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.63
cc_27 VNB N_VGND_c_322_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_28 VNB N_VGND_c_323_n 0.00510915f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.155
cc_29 VNB N_VGND_c_324_n 0.0619965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_325_n 0.172119f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_31 VPB N_D_M1001_g 0.0427627f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.63
cc_32 VPB N_D_c_62_n 0.00166729f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_33 VPB N_D_c_67_n 0.0321045f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.825
cc_34 VPB D 0.0445907f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_35 VPB N_C_M1006_g 0.0434257f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.63
cc_36 VPB C 0.00238326f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_37 VPB N_B_M1003_g 0.0428836f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.63
cc_38 VPB B 0.00288995f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_39 VPB N_A_M1000_g 0.0435375f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.445
cc_40 VPB N_A_c_191_n 0.00116914f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.155
cc_41 VPB N_A_c_198_n 0.0158467f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.825
cc_42 VPB A 0.00287133f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_234_n 0.0407451f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_44 VPB N_VPWR_c_235_n 0.0103017f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_45 VPB N_VPWR_c_236_n 0.0401575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_237_n 0.0174178f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.32
cc_47 VPB N_VPWR_c_238_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.32
cc_48 VPB N_VPWR_c_239_n 0.0170916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_240_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_241_n 0.0170916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_242_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.32
cc_52 VPB N_VPWR_c_243_n 0.013281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_233_n 0.0879491f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_Y_c_271_n 0.00703579f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.155
cc_55 VPB N_Y_c_272_n 0.00611905f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_56 VPB N_Y_c_273_n 0.00556397f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_57 VPB N_Y_c_269_n 0.0136633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_Y_c_275_n 0.0104711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_Y_c_276_n 0.00564143f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.32
cc_60 VPB N_Y_c_277_n 0.0307503f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.295
cc_61 N_D_c_62_n N_C_M1006_g 0.00584442f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_62 N_D_c_67_n N_C_M1006_g 0.0314245f $X=0.7 $Y=1.825 $X2=0 $Y2=0
cc_63 D N_C_M1006_g 5.7795e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_64 N_D_M1004_g N_C_c_95_n 0.0229844f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_65 N_D_c_62_n N_C_c_96_n 0.0229844f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_66 N_D_M1004_g C 0.00444194f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_67 N_D_c_62_n C 0.00213136f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_68 N_D_c_67_n C 7.58509e-19 $X=0.7 $Y=1.825 $X2=0 $Y2=0
cc_69 D C 0.0443454f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_70 D N_C_c_99_n 0.00192631f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_71 N_D_c_64_n N_C_c_99_n 0.0229844f $X=0.63 $Y=1.32 $X2=0 $Y2=0
cc_72 N_D_M1001_g N_VPWR_c_234_n 0.00432564f $X=0.86 $Y=2.63 $X2=0 $Y2=0
cc_73 N_D_c_67_n N_VPWR_c_234_n 0.00309196f $X=0.7 $Y=1.825 $X2=0 $Y2=0
cc_74 D N_VPWR_c_234_n 0.0218313f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_75 N_D_M1001_g N_VPWR_c_239_n 0.00570944f $X=0.86 $Y=2.63 $X2=0 $Y2=0
cc_76 N_D_M1001_g N_VPWR_c_233_n 0.00542671f $X=0.86 $Y=2.63 $X2=0 $Y2=0
cc_77 N_D_M1001_g N_Y_c_271_n 0.00237954f $X=0.86 $Y=2.63 $X2=0 $Y2=0
cc_78 D N_Y_c_271_n 0.0149808f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_79 N_D_M1001_g N_Y_c_272_n 0.00459558f $X=0.86 $Y=2.63 $X2=0 $Y2=0
cc_80 N_D_M1004_g N_VGND_c_321_n 0.0124262f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_81 D N_VGND_c_321_n 0.0207459f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_82 N_D_c_64_n N_VGND_c_321_n 6.21319e-19 $X=0.63 $Y=1.32 $X2=0 $Y2=0
cc_83 N_D_M1004_g N_VGND_c_324_n 0.00486043f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_84 N_D_M1004_g N_VGND_c_325_n 0.00693889f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_85 D N_VGND_c_325_n 0.012864f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_86 N_C_M1006_g N_B_M1003_g 0.0426691f $X=1.29 $Y=2.63 $X2=0 $Y2=0
cc_87 C N_B_M1003_g 3.18478e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_88 N_C_c_95_n N_B_c_142_n 0.0189742f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_89 C N_B_c_142_n 0.00123044f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_90 N_C_c_96_n N_B_c_143_n 0.011703f $X=1.2 $Y=1.27 $X2=0 $Y2=0
cc_91 N_C_c_97_n N_B_c_144_n 0.011703f $X=1.2 $Y=1.435 $X2=0 $Y2=0
cc_92 N_C_c_95_n B 0.00103717f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_93 C B 0.109213f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_94 N_C_c_99_n B 0.00607693f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_95 C N_B_c_146_n 7.02226e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_96 N_C_c_99_n N_B_c_146_n 0.011703f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_97 N_C_M1006_g N_VPWR_c_235_n 0.00188237f $X=1.29 $Y=2.63 $X2=0 $Y2=0
cc_98 N_C_M1006_g N_VPWR_c_239_n 0.00570944f $X=1.29 $Y=2.63 $X2=0 $Y2=0
cc_99 N_C_M1006_g N_VPWR_c_233_n 0.00542671f $X=1.29 $Y=2.63 $X2=0 $Y2=0
cc_100 N_C_c_97_n N_Y_c_271_n 6.74187e-19 $X=1.2 $Y=1.435 $X2=0 $Y2=0
cc_101 C N_Y_c_271_n 0.0158347f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_102 N_C_M1006_g N_Y_c_272_n 0.00259305f $X=1.29 $Y=2.63 $X2=0 $Y2=0
cc_103 N_C_M1006_g N_Y_c_275_n 0.0167942f $X=1.29 $Y=2.63 $X2=0 $Y2=0
cc_104 C N_Y_c_275_n 0.0111761f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_105 N_C_c_95_n N_VGND_c_321_n 0.00240392f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_106 C N_VGND_c_321_n 0.00951248f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_107 N_C_c_95_n N_VGND_c_324_n 0.00382867f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_108 C N_VGND_c_324_n 0.0110208f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_109 N_C_c_99_n N_VGND_c_324_n 7.20442e-19 $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_110 N_C_c_95_n N_VGND_c_325_n 0.00576641f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_111 C N_VGND_c_325_n 0.0106581f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_112 N_C_c_99_n N_VGND_c_325_n 4.27572e-19 $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_113 C A_237_47# 0.00379429f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_114 N_B_c_142_n N_A_M1002_g 0.017727f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_115 B N_A_M1002_g 0.00576247f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_116 N_B_c_146_n N_A_M1002_g 0.0115976f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_117 N_B_M1003_g N_A_c_198_n 0.0331581f $X=1.72 $Y=2.63 $X2=0 $Y2=0
cc_118 B N_A_c_198_n 2.33878e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_119 N_B_c_144_n N_A_c_192_n 0.0115976f $X=1.77 $Y=1.435 $X2=0 $Y2=0
cc_120 N_B_M1003_g N_A_c_193_n 0.00712579f $X=1.72 $Y=2.63 $X2=0 $Y2=0
cc_121 B N_A_c_193_n 6.40753e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_122 N_B_M1003_g A 0.00104882f $X=1.72 $Y=2.63 $X2=0 $Y2=0
cc_123 B A 0.0792574f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_124 N_B_c_146_n A 0.00472668f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_125 N_B_c_143_n N_A_c_195_n 0.0115976f $X=1.77 $Y=1.27 $X2=0 $Y2=0
cc_126 N_B_M1003_g N_VPWR_c_235_n 0.00188237f $X=1.72 $Y=2.63 $X2=0 $Y2=0
cc_127 N_B_M1003_g N_VPWR_c_241_n 0.00570944f $X=1.72 $Y=2.63 $X2=0 $Y2=0
cc_128 N_B_M1003_g N_VPWR_c_233_n 0.00542671f $X=1.72 $Y=2.63 $X2=0 $Y2=0
cc_129 N_B_M1003_g N_Y_c_273_n 0.00259305f $X=1.72 $Y=2.63 $X2=0 $Y2=0
cc_130 N_B_M1003_g N_Y_c_275_n 0.0166561f $X=1.72 $Y=2.63 $X2=0 $Y2=0
cc_131 B N_Y_c_275_n 0.023039f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_132 N_B_c_144_n N_Y_c_276_n 0.00298798f $X=1.77 $Y=1.435 $X2=0 $Y2=0
cc_133 B N_Y_c_276_n 0.00459114f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_134 N_B_c_142_n N_Y_c_270_n 6.66953e-19 $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_135 B N_Y_c_270_n 0.00928808f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 N_B_c_142_n N_VGND_c_324_n 0.00381508f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_137 B N_VGND_c_324_n 0.0107555f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_138 N_B_c_146_n N_VGND_c_324_n 0.00183241f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_139 N_B_c_142_n N_VGND_c_325_n 0.00620791f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_140 B N_VGND_c_325_n 0.0113807f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_141 N_B_c_146_n N_VGND_c_325_n 0.00213938f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_142 B A_237_47# 0.00288588f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_143 B A_351_47# 0.00430623f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_144 N_A_M1000_g N_VPWR_c_236_n 0.00408958f $X=2.15 $Y=2.63 $X2=0 $Y2=0
cc_145 N_A_M1000_g N_VPWR_c_241_n 0.00570944f $X=2.15 $Y=2.63 $X2=0 $Y2=0
cc_146 N_A_M1000_g N_VPWR_c_233_n 0.00542671f $X=2.15 $Y=2.63 $X2=0 $Y2=0
cc_147 N_A_M1000_g N_Y_c_273_n 0.00478965f $X=2.15 $Y=2.63 $X2=0 $Y2=0
cc_148 N_A_M1000_g N_Y_c_269_n 0.00265293f $X=2.15 $Y=2.63 $X2=0 $Y2=0
cc_149 N_A_M1002_g N_Y_c_269_n 0.00520665f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_c_191_n N_Y_c_269_n 0.00133173f $X=2.25 $Y=1.675 $X2=0 $Y2=0
cc_151 N_A_c_198_n N_Y_c_269_n 0.00249223f $X=2.25 $Y=1.75 $X2=0 $Y2=0
cc_152 A N_Y_c_269_n 0.0760885f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_153 N_A_c_195_n N_Y_c_269_n 0.0165356f $X=2.34 $Y=1.005 $X2=0 $Y2=0
cc_154 A N_Y_c_276_n 0.00365421f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_Y_c_270_n 0.00728652f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_156 A N_Y_c_270_n 0.00946419f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_157 N_A_c_195_n N_Y_c_270_n 0.003828f $X=2.34 $Y=1.005 $X2=0 $Y2=0
cc_158 N_A_M1000_g N_Y_c_277_n 0.0190282f $X=2.15 $Y=2.63 $X2=0 $Y2=0
cc_159 N_A_c_198_n N_Y_c_277_n 0.00288879f $X=2.25 $Y=1.75 $X2=0 $Y2=0
cc_160 N_A_c_193_n N_Y_c_277_n 0.00304381f $X=2.34 $Y=1.51 $X2=0 $Y2=0
cc_161 A N_Y_c_277_n 0.0290106f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_162 N_A_M1002_g N_VGND_c_324_n 0.00518687f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_M1002_g N_VGND_c_325_n 0.00757642f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_164 A N_VGND_c_325_n 0.0100177f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_165 N_VPWR_c_234_n N_Y_c_272_n 0.00226893f $X=0.645 $Y=2.455 $X2=0 $Y2=0
cc_166 N_VPWR_c_235_n N_Y_c_272_n 0.00144465f $X=1.505 $Y=2.465 $X2=0 $Y2=0
cc_167 N_VPWR_c_239_n N_Y_c_272_n 0.0106557f $X=1.375 $Y=3.33 $X2=0 $Y2=0
cc_168 N_VPWR_c_233_n N_Y_c_272_n 0.00941316f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_169 N_VPWR_c_235_n N_Y_c_273_n 0.00144465f $X=1.505 $Y=2.465 $X2=0 $Y2=0
cc_170 N_VPWR_c_236_n N_Y_c_273_n 0.0014586f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_171 N_VPWR_c_241_n N_Y_c_273_n 0.0106557f $X=2.235 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_233_n N_Y_c_273_n 0.00941316f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_173 N_VPWR_c_235_n N_Y_c_275_n 0.0221091f $X=1.505 $Y=2.465 $X2=0 $Y2=0
cc_174 N_VPWR_c_236_n N_Y_c_277_n 0.0251083f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_175 N_Y_c_270_n N_VGND_c_324_n 0.0280566f $X=2.695 $Y=0.445 $X2=0 $Y2=0
cc_176 N_Y_M1002_d N_VGND_c_325_n 0.00233781f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_177 N_Y_c_270_n N_VGND_c_325_n 0.019163f $X=2.695 $Y=0.445 $X2=0 $Y2=0
cc_178 N_VGND_c_325_n A_159_47# 0.010279f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_179 N_VGND_c_325_n A_237_47# 0.00913729f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_180 N_VGND_c_325_n A_351_47# 0.00841618f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
