* File: sky130_fd_sc_lp__nand2b_2.spice
* Created: Fri Aug 28 10:48:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2b_2.pex.spice"
.subckt sky130_fd_sc_lp__nand2b_2  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_N_M1008_g N_A_27_131#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1113 PD=0.856667 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1008_d N_B_M1000_g N_A_229_47#_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2184 AS=0.1365 PD=1.71333 PS=1.165 NRD=11.784 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_27_131#_M1003_g N_A_229_47#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1323 AS=0.1365 PD=1.155 PS=1.165 NRD=4.992 NRS=6.42 M=1 R=5.6
+ SA=75001 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1003_d N_A_27_131#_M1005_g N_A_229_47#_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1323 AS=0.1176 PD=1.155 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g N_A_229_47#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_A_N_M1001_g N_A_27_131#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.095025 AS=0.1197 PD=0.8175 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1001_d N_B_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=4.9447 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A_27_131#_M1004_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1004_d N_A_27_131#_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_B_M1007_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__nand2b_2.pxi.spice"
*
.ends
*
*
