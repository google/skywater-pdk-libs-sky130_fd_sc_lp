# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrtn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.375000 0.815000 2.005000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.573300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.075000 2.640000 6.635000 2.970000 ;
        RECT 6.090000 0.255000 6.635000 1.095000 ;
        RECT 6.370000 1.095000 6.635000 2.640000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.425000 0.840000 5.740000 2.130000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.800000 1.325000 2.005000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.195000  0.300000 0.455000 2.175000 ;
      RECT 0.195000  2.175000 1.235000 2.345000 ;
      RECT 0.195000  2.345000 0.465000 2.985000 ;
      RECT 0.685000  2.515000 0.895000 3.245000 ;
      RECT 0.985000  0.085000 1.205000 0.605000 ;
      RECT 1.065000  2.345000 1.235000 2.815000 ;
      RECT 1.065000  2.815000 2.045000 2.985000 ;
      RECT 1.375000  0.300000 1.705000 0.630000 ;
      RECT 1.405000  2.305000 1.705000 2.635000 ;
      RECT 1.495000  0.630000 1.705000 2.305000 ;
      RECT 1.875000  2.315000 2.990000 2.485000 ;
      RECT 1.875000  2.485000 2.045000 2.815000 ;
      RECT 1.915000  0.685000 2.245000 1.095000 ;
      RECT 1.915000  1.095000 3.460000 1.265000 ;
      RECT 1.915000  1.265000 2.245000 2.145000 ;
      RECT 2.425000  0.085000 2.755000 0.925000 ;
      RECT 2.500000  2.655000 2.830000 3.245000 ;
      RECT 2.660000  1.435000 2.990000 2.315000 ;
      RECT 2.925000  0.255000 3.890000 0.495000 ;
      RECT 2.925000  0.495000 3.145000 1.095000 ;
      RECT 3.200000  1.265000 3.460000 2.075000 ;
      RECT 3.325000  0.665000 3.800000 0.925000 ;
      RECT 3.340000  2.245000 3.800000 2.885000 ;
      RECT 3.630000  0.925000 3.800000 1.065000 ;
      RECT 3.630000  1.065000 4.905000 1.235000 ;
      RECT 3.630000  1.235000 3.800000 2.245000 ;
      RECT 4.100000  1.405000 4.430000 1.685000 ;
      RECT 4.100000  1.685000 5.255000 1.855000 ;
      RECT 4.100000  1.855000 4.430000 2.075000 ;
      RECT 4.225000  0.085000 4.555000 0.895000 ;
      RECT 4.295000  2.285000 4.915000 3.245000 ;
      RECT 4.650000  2.025000 4.915000 2.285000 ;
      RECT 4.655000  1.235000 4.905000 1.515000 ;
      RECT 4.745000  0.325000 5.255000 0.875000 ;
      RECT 5.075000  0.875000 5.255000 1.685000 ;
      RECT 5.085000  1.855000 5.255000 2.300000 ;
      RECT 5.085000  2.300000 6.200000 2.470000 ;
      RECT 5.085000  2.470000 5.385000 3.075000 ;
      RECT 5.575000  2.640000 5.905000 3.245000 ;
      RECT 5.590000  0.085000 5.920000 0.670000 ;
      RECT 5.950000  1.345000 6.200000 2.300000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrtn_1
