* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__maj3_2 A B C VGND VNB VPB VPWR X
X0 VPWR A a_310_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_59_491# C a_154_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_318_49# B a_59_491# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_59_491# B a_482_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 X a_59_491# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_474_491# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VPWR a_59_491# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_310_491# B a_59_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VGND A a_318_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_59_491# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_59_491# B a_474_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_59_491# C a_146_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_154_49# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_146_491# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_482_49# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_59_491# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
