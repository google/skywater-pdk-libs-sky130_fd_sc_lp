* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21bai_0 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 VGND A1 a_320_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_39_51# Y VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 Y A2 a_406_473# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_39_51# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_39_51# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_406_473# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 Y a_39_51# a_320_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_320_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
