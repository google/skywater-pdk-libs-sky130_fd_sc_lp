* File: sky130_fd_sc_lp__bufkapwr_8.pex.spice
* Created: Wed Sep  2 09:36:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_8%A 3 7 11 15 17 18 26
r41 25 26 34.3377 $w=6.7e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.905 $Y2=1.235
r42 22 25 16.3703 $w=6.7e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.235
+ $X2=0.475 $Y2=1.235
r43 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.065 $X2=0.27 $Y2=1.065
r44 18 23 8.41466 $w=3.13e-07 $l=2.3e-07 $layer=LI1_cond $X=0.242 $Y=1.295
+ $X2=0.242 $Y2=1.065
r45 17 23 5.12197 $w=3.13e-07 $l=1.4e-07 $layer=LI1_cond $X=0.242 $Y=0.925
+ $X2=0.242 $Y2=1.065
r46 13 26 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.905 $Y=1.57
+ $X2=0.905 $Y2=1.235
r47 13 15 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=0.905 $Y=1.57
+ $X2=0.905 $Y2=2.465
r48 9 26 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=1.235
r49 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=0.445
r50 5 25 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.475 $Y=1.57
+ $X2=0.475 $Y2=1.235
r51 5 7 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=0.475 $Y=1.57
+ $X2=0.475 $Y2=2.465
r52 1 25 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=1.235
r53 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_8%A_110_47# 1 2 9 13 17 21 25 29 33 37 41
+ 45 49 53 57 61 65 69 73 77 86 89 100
r169 99 100 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.915 $Y=1.32
+ $X2=4.345 $Y2=1.32
r170 98 99 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.485 $Y=1.32
+ $X2=3.915 $Y2=1.32
r171 95 96 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.625 $Y=1.32
+ $X2=3.055 $Y2=1.32
r172 94 95 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.195 $Y=1.32
+ $X2=2.625 $Y2=1.32
r173 93 94 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.765 $Y=1.32
+ $X2=2.195 $Y2=1.32
r174 87 98 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.245 $Y=1.32
+ $X2=3.485 $Y2=1.32
r175 87 96 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.245 $Y=1.32
+ $X2=3.055 $Y2=1.32
r176 86 87 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.245
+ $Y=1.32 $X2=3.245 $Y2=1.32
r177 84 93 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.545 $Y=1.32
+ $X2=1.765 $Y2=1.32
r178 84 90 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.545 $Y=1.32
+ $X2=1.335 $Y2=1.32
r179 83 86 59.3683 $w=3.28e-07 $l=1.7e-06 $layer=LI1_cond $X=1.545 $Y=1.32
+ $X2=3.245 $Y2=1.32
r180 83 84 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=1.545
+ $Y=1.32 $X2=1.545 $Y2=1.32
r181 81 89 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=1.32
+ $X2=0.695 $Y2=1.32
r182 81 83 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=0.82 $Y=1.32
+ $X2=1.545 $Y2=1.32
r183 77 79 39.1831 $w=2.48e-07 $l=8.5e-07 $layer=LI1_cond $X=0.695 $Y=2.04
+ $X2=0.695 $Y2=2.89
r184 75 89 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=1.485
+ $X2=0.695 $Y2=1.32
r185 75 77 25.5842 $w=2.48e-07 $l=5.55e-07 $layer=LI1_cond $X=0.695 $Y=1.485
+ $X2=0.695 $Y2=2.04
r186 71 89 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=1.155
+ $X2=0.695 $Y2=1.32
r187 71 73 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.695 $Y=1.155
+ $X2=0.695 $Y2=0.445
r188 67 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.485
+ $X2=4.345 $Y2=1.32
r189 67 69 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.345 $Y=1.485
+ $X2=4.345 $Y2=2.465
r190 63 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.155
+ $X2=4.345 $Y2=1.32
r191 63 65 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.345 $Y=1.155
+ $X2=4.345 $Y2=0.445
r192 59 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.485
+ $X2=3.915 $Y2=1.32
r193 59 61 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.915 $Y=1.485
+ $X2=3.915 $Y2=2.465
r194 55 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.155
+ $X2=3.915 $Y2=1.32
r195 55 57 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.915 $Y=1.155
+ $X2=3.915 $Y2=0.445
r196 51 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.485
+ $X2=3.485 $Y2=1.32
r197 51 53 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.485 $Y=1.485
+ $X2=3.485 $Y2=2.465
r198 47 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.155
+ $X2=3.485 $Y2=1.32
r199 47 49 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.485 $Y=1.155
+ $X2=3.485 $Y2=0.445
r200 43 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.485
+ $X2=3.055 $Y2=1.32
r201 43 45 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.055 $Y=1.485
+ $X2=3.055 $Y2=2.465
r202 39 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.155
+ $X2=3.055 $Y2=1.32
r203 39 41 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.055 $Y=1.155
+ $X2=3.055 $Y2=0.445
r204 35 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.485
+ $X2=2.625 $Y2=1.32
r205 35 37 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.625 $Y=1.485
+ $X2=2.625 $Y2=2.465
r206 31 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.155
+ $X2=2.625 $Y2=1.32
r207 31 33 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.625 $Y=1.155
+ $X2=2.625 $Y2=0.445
r208 27 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.485
+ $X2=2.195 $Y2=1.32
r209 27 29 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.195 $Y=1.485
+ $X2=2.195 $Y2=2.465
r210 23 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.155
+ $X2=2.195 $Y2=1.32
r211 23 25 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.195 $Y=1.155
+ $X2=2.195 $Y2=0.445
r212 19 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.485
+ $X2=1.765 $Y2=1.32
r213 19 21 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.765 $Y=1.485
+ $X2=1.765 $Y2=2.465
r214 15 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.155
+ $X2=1.765 $Y2=1.32
r215 15 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.765 $Y=1.155
+ $X2=1.765 $Y2=0.445
r216 11 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.485
+ $X2=1.335 $Y2=1.32
r217 11 13 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.335 $Y=1.485
+ $X2=1.335 $Y2=2.465
r218 7 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.155
+ $X2=1.335 $Y2=1.32
r219 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.335 $Y=1.155
+ $X2=1.335 $Y2=0.445
r220 2 79 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.89
r221 2 77 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.04
r222 1 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_8%KAPWR 1 2 3 4 5 6 19 22 30 38 46 54 62 66
+ 75
r69 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.575 $Y=2.81
+ $X2=4.575 $Y2=2.81
r70 62 65 22.6582 $w=2.93e-07 $l=5.8e-07 $layer=LI1_cond $X=4.577 $Y=2.23
+ $X2=4.577 $Y2=2.81
r71 58 66 0.512151 $w=2.55e-07 $l=8.85e-07 $layer=MET1_cond $X=3.69 $Y=2.817
+ $X2=4.575 $Y2=2.817
r72 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.69 $Y=2.81
+ $X2=3.69 $Y2=2.81
r73 54 57 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=3.7 $Y=2.23 $X2=3.7
+ $Y2=2.81
r74 50 58 0.49479 $w=2.55e-07 $l=8.55e-07 $layer=MET1_cond $X=2.835 $Y=2.817
+ $X2=3.69 $Y2=2.817
r75 50 75 0.109953 $w=2.55e-07 $l=1.9e-07 $layer=MET1_cond $X=2.835 $Y=2.817
+ $X2=2.645 $Y2=2.817
r76 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.835 $Y=2.81
+ $X2=2.835 $Y2=2.81
r77 46 49 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=2.84 $Y=2.23
+ $X2=2.84 $Y2=2.81
r78 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.975 $Y=2.81
+ $X2=1.975 $Y2=2.81
r79 38 41 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=1.98 $Y=2.23
+ $X2=1.98 $Y2=2.81
r80 34 42 0.491897 $w=2.55e-07 $l=8.5e-07 $layer=MET1_cond $X=1.125 $Y=2.817
+ $X2=1.975 $Y2=2.817
r81 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.125 $Y=2.81
+ $X2=1.125 $Y2=2.81
r82 30 33 34.13 $w=2.58e-07 $l=7.7e-07 $layer=LI1_cond $X=1.12 $Y=2.04 $X2=1.12
+ $Y2=2.81
r83 26 34 0.506364 $w=2.55e-07 $l=8.75e-07 $layer=MET1_cond $X=0.25 $Y=2.817
+ $X2=1.125 $Y2=2.817
r84 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.25 $Y=2.81
+ $X2=0.25 $Y2=2.81
r85 22 25 30.0807 $w=2.93e-07 $l=7.7e-07 $layer=LI1_cond $X=0.242 $Y=2.04
+ $X2=0.242 $Y2=2.81
r86 19 75 0.00289351 $w=2.55e-07 $l=5e-09 $layer=MET1_cond $X=2.64 $Y=2.817
+ $X2=2.645 $Y2=2.817
r87 19 42 0.384837 $w=2.55e-07 $l=6.65e-07 $layer=MET1_cond $X=2.64 $Y=2.817
+ $X2=1.975 $Y2=2.817
r88 6 65 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.835 $X2=4.56 $Y2=2.91
r89 6 62 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.835 $X2=4.56 $Y2=2.23
r90 5 57 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.91
r91 5 54 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.23
r92 4 49 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.91
r93 4 46 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.23
r94 3 41 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.91
r95 3 38 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.23
r96 2 33 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.89
r97 2 30 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.04
r98 1 25 400 $w=1.7e-07 $l=1.11575e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.89
r99 1 22 400 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_8%X 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45
+ 49 51 55 59 63 65 69 73 77 78 79 80 81 82 83
r151 83 98 2.23356 $w=6.15e-07 $l=1.2e-07 $layer=LI1_cond $X=4.245 $Y=1.775
+ $X2=4.245 $Y2=1.655
r152 83 98 0.477938 $w=9.68e-07 $l=3.8e-08 $layer=LI1_cond $X=4.245 $Y=1.617
+ $X2=4.245 $Y2=1.655
r153 82 83 4.0499 $w=9.68e-07 $l=3.22e-07 $layer=LI1_cond $X=4.245 $Y=1.295
+ $X2=4.245 $Y2=1.617
r154 81 97 2.23356 $w=6.15e-07 $l=1.2e-07 $layer=LI1_cond $X=4.245 $Y=0.855
+ $X2=4.245 $Y2=0.975
r155 81 82 3.81093 $w=9.68e-07 $l=3.03e-07 $layer=LI1_cond $X=4.245 $Y=0.992
+ $X2=4.245 $Y2=1.295
r156 81 97 0.213814 $w=9.68e-07 $l=1.7e-08 $layer=LI1_cond $X=4.245 $Y=0.992
+ $X2=4.245 $Y2=0.975
r157 73 75 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=4.13 $Y=2.04
+ $X2=4.13 $Y2=2.89
r158 71 83 2.23356 $w=6.15e-07 $l=1.67929e-07 $layer=LI1_cond $X=4.13 $Y=1.895
+ $X2=4.245 $Y2=1.775
r159 71 73 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=4.13 $Y=1.895
+ $X2=4.13 $Y2=2.04
r160 67 81 2.23356 $w=6.15e-07 $l=1.67929e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.245 $Y2=0.855
r161 67 69 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.13 $Y2=0.445
r162 66 80 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=1.775
+ $X2=3.27 $Y2=1.775
r163 65 83 4.87019 $w=2.4e-07 $l=4.85e-07 $layer=LI1_cond $X=3.76 $Y=1.775
+ $X2=4.245 $Y2=1.775
r164 65 66 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=3.76 $Y=1.775
+ $X2=3.4 $Y2=1.775
r165 64 79 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=0.855
+ $X2=3.27 $Y2=0.855
r166 63 81 4.87019 $w=2.4e-07 $l=4.85e-07 $layer=LI1_cond $X=3.76 $Y=0.855
+ $X2=4.245 $Y2=0.855
r167 63 64 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=3.76 $Y=0.855
+ $X2=3.4 $Y2=0.855
r168 59 61 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=3.27 $Y=2.04
+ $X2=3.27 $Y2=2.89
r169 57 80 1.05597 $w=2.6e-07 $l=1.2e-07 $layer=LI1_cond $X=3.27 $Y=1.895
+ $X2=3.27 $Y2=1.775
r170 57 59 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=3.27 $Y=1.895
+ $X2=3.27 $Y2=2.04
r171 53 79 1.05597 $w=2.6e-07 $l=1.2e-07 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.855
r172 53 55 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.445
r173 52 78 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=1.775
+ $X2=2.41 $Y2=1.775
r174 51 80 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=1.775
+ $X2=3.27 $Y2=1.775
r175 51 52 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=1.775
+ $X2=2.54 $Y2=1.775
r176 50 77 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=0.855
+ $X2=2.41 $Y2=0.855
r177 49 79 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=0.855
+ $X2=3.27 $Y2=0.855
r178 49 50 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=0.855
+ $X2=2.54 $Y2=0.855
r179 45 47 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=2.41 $Y=2.04
+ $X2=2.41 $Y2=2.89
r180 43 78 1.05597 $w=2.6e-07 $l=1.2e-07 $layer=LI1_cond $X=2.41 $Y=1.895
+ $X2=2.41 $Y2=1.775
r181 43 45 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=2.41 $Y=1.895
+ $X2=2.41 $Y2=2.04
r182 39 77 1.05597 $w=2.6e-07 $l=1.2e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.855
r183 39 41 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.445
r184 37 78 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=1.775
+ $X2=2.41 $Y2=1.775
r185 37 38 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=2.28 $Y=1.775
+ $X2=1.68 $Y2=1.775
r186 35 77 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=0.855
+ $X2=2.41 $Y2=0.855
r187 35 36 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=2.28 $Y=0.855
+ $X2=1.68 $Y2=0.855
r188 31 33 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=1.55 $Y=2.04
+ $X2=1.55 $Y2=2.89
r189 29 38 6.83069 $w=2.4e-07 $l=1.80278e-07 $layer=LI1_cond $X=1.55 $Y=1.895
+ $X2=1.68 $Y2=1.775
r190 29 31 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.55 $Y=1.895
+ $X2=1.55 $Y2=2.04
r191 25 36 6.83069 $w=2.4e-07 $l=1.80278e-07 $layer=LI1_cond $X=1.55 $Y=0.735
+ $X2=1.68 $Y2=0.855
r192 25 27 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=1.55 $Y=0.735
+ $X2=1.55 $Y2=0.445
r193 8 75 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.835 $X2=4.13 $Y2=2.89
r194 8 73 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.835 $X2=4.13 $Y2=2.04
r195 7 61 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.89
r196 7 59 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.04
r197 6 47 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.89
r198 6 45 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.04
r199 5 33 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.89
r200 5 31 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.04
r201 4 69 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.235 $X2=4.13 $Y2=0.445
r202 3 55 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.445
r203 2 41 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.445
r204 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_8%VGND 1 2 3 4 5 6 19 21 25 29 33 35 39 43
+ 46 47 49 50 51 52 53 65 72 73 79 82
r83 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r84 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r85 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r86 73 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r87 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r88 70 82 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.58
+ $Y2=0
r89 70 72 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=5.04
+ $Y2=0
r90 69 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r91 69 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r92 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r93 66 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.7
+ $Y2=0
r94 66 68 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=4.08
+ $Y2=0
r95 65 82 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.58
+ $Y2=0
r96 65 68 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.08
+ $Y2=0
r97 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r98 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r99 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r100 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r101 55 76 3.93884 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r102 55 57 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.72
+ $Y2=0
r103 53 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r104 53 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r105 53 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r106 51 63 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.64
+ $Y2=0
r107 51 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.84
+ $Y2=0
r108 49 60 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.68
+ $Y2=0
r109 49 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.98
+ $Y2=0
r110 48 63 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.64
+ $Y2=0
r111 48 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=1.98
+ $Y2=0
r112 46 57 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r113 46 47 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.12
+ $Y2=0
r114 45 60 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.68
+ $Y2=0
r115 45 47 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.12
+ $Y2=0
r116 41 82 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0
r117 41 43 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0.4
r118 37 79 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0
r119 37 39 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.4
r120 36 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=2.84
+ $Y2=0
r121 35 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.7
+ $Y2=0
r122 35 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=2.97
+ $Y2=0
r123 31 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r124 31 33 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.4
r125 27 50 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r126 27 29 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.4
r127 23 47 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r128 23 25 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.445
r129 19 76 3.17127 $w=2.45e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.195 $Y2=0
r130 19 21 16.9339 $w=2.43e-07 $l=3.6e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.267 $Y2=0.445
r131 6 43 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.235 $X2=4.565 $Y2=0.4
r132 5 39 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.4
r133 4 33 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.4
r134 3 29 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.4
r135 2 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.445
r136 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_8%VPWR 1 8 14
r58 5 14 0.00288826 $w=5.28e-06 $l=1.22e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.208
r59 5 8 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r60 4 8 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=5.04
+ $Y2=3.33
r61 4 5 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 1 14 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=3.207
+ $X2=2.64 $Y2=3.208
.ends

