* File: sky130_fd_sc_lp__dlrbn_1.spice
* Created: Fri Aug 28 10:25:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrbn_1.pex.spice"
.subckt sky130_fd_sc_lp__dlrbn_1  VNB VPB GATE_N D RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* GATE_N	GATE_N
* VPB	VPB
* VNB	VNB
MM1009 N_A_112_70#_M1009_d N_GATE_N_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_112_70#_M1001_g N_A_207_40#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_437_144#_M1017_d N_D_M1017_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1016 N_A_630_167#_M1016_d N_A_112_70#_M1016_g N_A_547_167#_M1016_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_716_167#_M1007_d N_A_207_40#_M1007_g N_A_630_167#_M1016_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_437_144#_M1019_g N_A_547_167#_M1019_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1021 N_A_716_167#_M1021_d N_A_955_271#_M1021_g N_VGND_M1019_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 A_1211_47# N_A_630_167#_M1008_g N_A_955_271#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_RESET_B_M1010_g A_1211_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2464 AS=0.0882 PD=1.94 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1023 N_A_1394_367#_M1023_d N_A_955_271#_M1023_g N_VGND_M1010_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1512 AS=0.1232 PD=1.56 PS=0.97 NRD=27.132 NRS=68.088 M=1
+ R=2.8 SA=75001.3 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_1394_367#_M1002_g N_Q_N_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.2226 PD=1.37 PS=2.21 NRD=35.712 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1006 N_Q_M1006_d N_A_955_271#_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.2226 PD=2.25 PS=1.37 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_A_112_70#_M1011_d N_GATE_N_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A_112_70#_M1005_g N_A_207_40#_M1005_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1392 AS=0.1696 PD=1.075 PS=1.81 NRD=23.0687 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1018 N_A_437_144#_M1018_d N_D_M1018_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1392 PD=1.81 PS=1.075 NRD=0 NRS=24.6053 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_A_630_167#_M1000_d N_A_112_70#_M1000_g N_A_625_377#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0855057 AS=0.1113 PD=0.80434 PS=1.37 NRD=69.6789 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1013 A_813_377# N_A_207_40#_M1013_g N_A_630_167#_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0672 AS=0.130294 PD=0.85 PS=1.22566 NRD=15.3857 NRS=0 M=1
+ R=4.26667 SA=75000.5 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1015 N_VPWR_M1015_d N_A_437_144#_M1015_g A_813_377# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.130294 AS=0.0672 PD=1.22566 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75000.9 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1004 N_A_625_377#_M1004_d N_A_955_271#_M1004_g N_VPWR_M1015_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0855057 PD=1.37 PS=0.80434 NRD=0 NRS=46.886 M=1
+ R=2.8 SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_955_271#_M1012_d N_A_630_167#_M1012_g N_VPWR_M1012_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_RESET_B_M1003_g N_A_955_271#_M1012_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.268115 AS=0.1764 PD=2.16853 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1020 N_A_1394_367#_M1020_d N_A_955_271#_M1020_g N_VPWR_M1003_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.136185 PD=1.81 PS=1.10147 NRD=0 NRS=20.7638 M=1
+ R=4.26667 SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1022 N_VPWR_M1022_d N_A_1394_367#_M1022_g N_Q_N_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_Q_M1014_d N_A_955_271#_M1014_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=18.6777 P=23.77
c_191 VPB 0 6.36774e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlrbn_1.pxi.spice"
*
.ends
*
*
