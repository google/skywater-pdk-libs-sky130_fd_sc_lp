# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a311oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a311oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.290000 1.425000 3.685000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.385000 1.415000 2.735000 1.585000 ;
        RECT 1.940000 1.585000 2.735000 1.750000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.415000 1.105000 1.585000 ;
        RECT 0.155000 1.585000 0.550000 1.750000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.900000 1.425000 4.230000 1.750000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.425000 5.675000 1.750000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.352400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.920000 5.195000 2.120000 ;
        RECT 2.655000 0.595000 2.995000 1.085000 ;
        RECT 2.655000 1.085000 5.665000 1.245000 ;
        RECT 2.905000 1.245000 5.665000 1.255000 ;
        RECT 2.905000 1.255000 3.075000 1.920000 ;
        RECT 3.665000 0.305000 3.855000 1.085000 ;
        RECT 4.525000 0.305000 4.715000 1.085000 ;
        RECT 4.920000 2.120000 5.195000 2.735000 ;
        RECT 5.385000 0.305000 5.665000 1.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.220000  0.325000 0.480000 1.075000 ;
      RECT 0.220000  1.075000 2.350000 1.245000 ;
      RECT 0.220000  1.920000 0.550000 3.245000 ;
      RECT 0.650000  0.085000 0.980000 0.905000 ;
      RECT 0.720000  1.755000 1.770000 1.925000 ;
      RECT 0.720000  1.925000 0.900000 3.075000 ;
      RECT 1.080000  2.095000 1.410000 3.245000 ;
      RECT 1.150000  0.325000 1.340000 1.075000 ;
      RECT 1.510000  0.255000 3.495000 0.425000 ;
      RECT 1.510000  0.425000 1.840000 0.905000 ;
      RECT 1.580000  1.925000 1.770000 2.290000 ;
      RECT 1.580000  2.290000 4.320000 2.460000 ;
      RECT 1.580000  2.460000 1.840000 3.075000 ;
      RECT 2.010000  0.595000 2.350000 1.075000 ;
      RECT 2.060000  2.630000 2.390000 3.245000 ;
      RECT 2.605000  2.460000 2.865000 3.075000 ;
      RECT 3.035000  2.630000 3.365000 3.245000 ;
      RECT 3.165000  0.425000 3.495000 0.895000 ;
      RECT 3.595000  2.800000 4.750000 2.905000 ;
      RECT 3.595000  2.905000 5.645000 3.075000 ;
      RECT 4.025000  0.085000 4.355000 0.915000 ;
      RECT 4.025000  2.460000 4.320000 2.630000 ;
      RECT 4.490000  2.290000 4.750000 2.800000 ;
      RECT 4.885000  0.085000 5.215000 0.915000 ;
      RECT 5.365000  1.920000 5.645000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__a311oi_2
