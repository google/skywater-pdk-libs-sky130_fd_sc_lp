* File: sky130_fd_sc_lp__xor2_lp.pxi.spice
* Created: Wed Sep  2 10:41:29 2020
* 
x_PM_SKY130_FD_SC_LP__XOR2_LP%A_84_93# N_A_84_93#_M1003_d N_A_84_93#_M1010_s
+ N_A_84_93#_M1002_g N_A_84_93#_M1004_g N_A_84_93#_M1012_g N_A_84_93#_c_85_n
+ N_A_84_93#_c_86_n N_A_84_93#_c_147_p N_A_84_93#_c_87_n N_A_84_93#_c_79_n
+ N_A_84_93#_c_88_n N_A_84_93#_c_80_n N_A_84_93#_c_81_n N_A_84_93#_c_82_n
+ N_A_84_93#_c_83_n N_A_84_93#_c_91_n N_A_84_93#_c_92_n
+ PM_SKY130_FD_SC_LP__XOR2_LP%A_84_93#
x_PM_SKY130_FD_SC_LP__XOR2_LP%A N_A_c_197_n N_A_M1001_g N_A_c_186_n N_A_c_187_n
+ N_A_M1006_g N_A_M1008_g N_A_M1011_g N_A_M1009_g N_A_c_192_n N_A_c_200_n
+ N_A_c_193_n A A N_A_c_194_n N_A_c_195_n N_A_c_196_n
+ PM_SKY130_FD_SC_LP__XOR2_LP%A
x_PM_SKY130_FD_SC_LP__XOR2_LP%B N_B_M1000_g N_B_c_292_n N_B_c_293_n N_B_c_301_n
+ N_B_M1005_g N_B_c_302_n N_B_c_303_n N_B_M1007_g N_B_c_295_n N_B_c_305_n
+ N_B_c_296_n N_B_M1003_g N_B_c_306_n N_B_M1010_g N_B_c_297_n N_B_c_307_n B
+ N_B_c_299_n N_B_c_300_n PM_SKY130_FD_SC_LP__XOR2_LP%B
x_PM_SKY130_FD_SC_LP__XOR2_LP%X N_X_M1012_d N_X_M1004_s N_X_c_377_n N_X_c_378_n
+ N_X_c_379_n N_X_c_380_n X X X X X PM_SKY130_FD_SC_LP__XOR2_LP%X
x_PM_SKY130_FD_SC_LP__XOR2_LP%A_159_419# N_A_159_419#_M1004_d
+ N_A_159_419#_M1005_d N_A_159_419#_c_425_n N_A_159_419#_c_426_n
+ N_A_159_419#_c_421_n PM_SKY130_FD_SC_LP__XOR2_LP%A_159_419#
x_PM_SKY130_FD_SC_LP__XOR2_LP%VPWR N_VPWR_M1001_d N_VPWR_M1011_d N_VPWR_c_452_n
+ N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n VPWR
+ N_VPWR_c_457_n N_VPWR_c_451_n PM_SKY130_FD_SC_LP__XOR2_LP%VPWR
x_PM_SKY130_FD_SC_LP__XOR2_LP%VGND N_VGND_M1002_s N_VGND_M1006_d N_VGND_M1009_d
+ N_VGND_c_495_n N_VGND_c_496_n N_VGND_c_497_n N_VGND_c_498_n N_VGND_c_499_n
+ N_VGND_c_500_n N_VGND_c_501_n VGND N_VGND_c_502_n N_VGND_c_503_n
+ PM_SKY130_FD_SC_LP__XOR2_LP%VGND
cc_1 VNB N_A_84_93#_M1002_g 0.0456751f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_2 VNB N_A_84_93#_M1012_g 0.0393457f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.805
cc_3 VNB N_A_84_93#_c_79_n 0.00228193f $X=-0.19 $Y=-0.245 $X2=2.76 $Y2=0.55
cc_4 VNB N_A_84_93#_c_80_n 0.0155442f $X=-0.19 $Y=-0.245 $X2=3.445 $Y2=0.915
cc_5 VNB N_A_84_93#_c_81_n 0.00719818f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=0.915
cc_6 VNB N_A_84_93#_c_82_n 0.0299904f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.04
cc_7 VNB N_A_84_93#_c_83_n 0.00947449f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.73
cc_8 VNB N_A_c_186_n 0.0173331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_187_n 0.0068954f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.565
cc_10 VNB N_A_M1006_g 0.0295893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_M1008_g 0.0296397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_M1011_g 0.0104987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_M1009_g 0.0363412f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.125
cc_14 VNB N_A_c_192_n 0.00163592f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.9
cc_15 VNB N_A_c_193_n 0.00229623f $X=-0.19 $Y=-0.245 $X2=2.76 $Y2=0.55
cc_16 VNB N_A_c_194_n 0.0320125f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.73
cc_17 VNB N_A_c_195_n 0.0400158f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.73
cc_18 VNB N_A_c_196_n 0.0183941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_M1000_g 0.0358484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_c_292_n 0.0624425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_293_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_M1007_g 0.0084304f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.565
cc_23 VNB N_B_c_295_n 0.0102f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.895
cc_24 VNB N_B_c_296_n 0.0144954f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.125
cc_25 VNB N_B_c_297_n 0.0281827f $X=-0.19 $Y=-0.245 $X2=3.445 $Y2=2.125
cc_26 VNB B 0.00791867f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=0.915
cc_27 VNB N_B_c_299_n 0.0248428f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.73
cc_28 VNB N_B_c_300_n 0.0142062f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.73
cc_29 VNB N_X_c_377_n 0.0102865f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.565
cc_30 VNB N_X_c_378_n 0.00984489f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_31 VNB N_X_c_379_n 0.0018379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_380_n 0.0116206f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.565
cc_33 VNB X 0.0133278f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.805
cc_34 VNB N_VPWR_c_451_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.04
cc_35 VNB N_VGND_c_495_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_496_n 0.0491446f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.595
cc_37 VNB N_VGND_c_497_n 0.00903781f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.805
cc_38 VNB N_VGND_c_498_n 0.0121187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_499_n 0.0208932f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.04
cc_40 VNB N_VGND_c_500_n 0.0387104f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.21
cc_41 VNB N_VGND_c_501_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.9
cc_42 VNB N_VGND_c_502_n 0.0365488f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=0.915
cc_43 VNB N_VGND_c_503_n 0.236089f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.73
cc_44 VPB N_A_84_93#_M1004_g 0.0310647f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.595
cc_45 VPB N_A_84_93#_c_85_n 0.0015051f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.04
cc_46 VPB N_A_84_93#_c_86_n 0.0205898f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=2.125
cc_47 VPB N_A_84_93#_c_87_n 0.0110041f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.9
cc_48 VPB N_A_84_93#_c_88_n 0.00355229f $X=-0.19 $Y=1.655 $X2=3.445 $Y2=2.125
cc_49 VPB N_A_84_93#_c_82_n 0.0174505f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=2.04
cc_50 VPB N_A_84_93#_c_83_n 0.0283036f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.73
cc_51 VPB N_A_84_93#_c_91_n 0.00144641f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.73
cc_52 VPB N_A_84_93#_c_92_n 0.00233943f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.205
cc_53 VPB N_A_c_197_n 0.026482f $X=-0.19 $Y=1.655 $X2=2.62 $Y2=0.34
cc_54 VPB N_A_M1011_g 0.0446064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_c_192_n 0.0168875f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.9
cc_56 VPB N_A_c_200_n 0.0230537f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.9
cc_57 VPB N_A_c_193_n 4.71068e-19 $X=-0.19 $Y=1.655 $X2=2.76 $Y2=0.55
cc_58 VPB N_A_c_196_n 0.00499601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_B_c_301_n 0.0267958f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.565
cc_60 VPB N_B_c_302_n 0.0257658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_B_c_303_n 0.00936306f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.895
cc_62 VPB N_B_c_295_n 0.00984047f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.895
cc_63 VPB N_B_c_305_n 0.0254665f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.04
cc_64 VPB N_B_c_306_n 0.0242879f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.9
cc_65 VPB N_B_c_307_n 0.00613356f $X=-0.19 $Y=1.655 $X2=3.445 $Y2=0.915
cc_66 VPB X 0.0213318f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.805
cc_67 VPB X 0.0133383f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB X 0.034084f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.895
cc_69 VPB N_A_159_419#_c_421_n 0.00631557f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.805
cc_70 VPB N_VPWR_c_452_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.805
cc_71 VPB N_VPWR_c_453_n 0.0115621f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.895
cc_72 VPB N_VPWR_c_454_n 0.030732f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.595
cc_73 VPB N_VPWR_c_455_n 0.0354905f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.805
cc_74 VPB N_VPWR_c_456_n 0.00436844f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.805
cc_75 VPB N_VPWR_c_457_n 0.0478688f $X=-0.19 $Y=1.655 $X2=2.76 $Y2=0.83
cc_76 VPB N_VPWR_c_451_n 0.0682666f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=2.04
cc_77 N_A_84_93#_M1004_g N_A_c_197_n 0.0254707f $X=0.67 $Y=2.595 $X2=-0.19
+ $Y2=-0.245
cc_78 N_A_84_93#_c_85_n N_A_c_197_n 0.00177549f $X=0.82 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_79 N_A_84_93#_c_86_n N_A_c_197_n 0.0145638f $X=2.395 $Y=2.125 $X2=-0.19
+ $Y2=-0.245
cc_80 N_A_84_93#_c_86_n N_A_c_186_n 0.00116015f $X=2.395 $Y=2.125 $X2=0 $Y2=0
cc_81 N_A_84_93#_M1012_g N_A_c_187_n 0.00612329f $X=0.855 $Y=0.805 $X2=0 $Y2=0
cc_82 N_A_84_93#_M1012_g N_A_M1006_g 0.00481307f $X=0.855 $Y=0.805 $X2=0 $Y2=0
cc_83 N_A_84_93#_c_79_n N_A_M1008_g 0.00996701f $X=2.76 $Y=0.55 $X2=0 $Y2=0
cc_84 N_A_84_93#_c_80_n N_A_M1008_g 0.0083362f $X=3.445 $Y=0.915 $X2=0 $Y2=0
cc_85 N_A_84_93#_c_81_n N_A_M1008_g 0.00355688f $X=2.925 $Y=0.915 $X2=0 $Y2=0
cc_86 N_A_84_93#_c_87_n N_A_M1011_g 0.00255408f $X=2.56 $Y=2.9 $X2=0 $Y2=0
cc_87 N_A_84_93#_c_88_n N_A_M1011_g 0.0267847f $X=3.445 $Y=2.125 $X2=0 $Y2=0
cc_88 N_A_84_93#_c_79_n N_A_M1009_g 0.00179788f $X=2.76 $Y=0.55 $X2=0 $Y2=0
cc_89 N_A_84_93#_c_80_n N_A_M1009_g 0.0166982f $X=3.445 $Y=0.915 $X2=0 $Y2=0
cc_90 N_A_84_93#_c_82_n N_A_M1009_g 0.0329558f $X=3.53 $Y=2.04 $X2=0 $Y2=0
cc_91 N_A_84_93#_M1004_g N_A_c_192_n 0.00160606f $X=0.67 $Y=2.595 $X2=0 $Y2=0
cc_92 N_A_84_93#_c_85_n N_A_c_192_n 0.00114816f $X=0.82 $Y=2.04 $X2=0 $Y2=0
cc_93 N_A_84_93#_c_83_n N_A_c_192_n 0.013166f $X=0.7 $Y=1.73 $X2=0 $Y2=0
cc_94 N_A_84_93#_c_91_n N_A_c_192_n 0.00119217f $X=0.82 $Y=1.73 $X2=0 $Y2=0
cc_95 N_A_84_93#_c_88_n N_A_c_200_n 0.0392523f $X=3.445 $Y=2.125 $X2=0 $Y2=0
cc_96 N_A_84_93#_c_82_n N_A_c_200_n 0.0130054f $X=3.53 $Y=2.04 $X2=0 $Y2=0
cc_97 N_A_84_93#_c_92_n N_A_c_200_n 0.0253273f $X=2.56 $Y=2.205 $X2=0 $Y2=0
cc_98 N_A_84_93#_c_80_n N_A_c_193_n 0.0246548f $X=3.445 $Y=0.915 $X2=0 $Y2=0
cc_99 N_A_84_93#_c_82_n N_A_c_193_n 0.0366358f $X=3.53 $Y=2.04 $X2=0 $Y2=0
cc_100 N_A_84_93#_c_86_n N_A_c_194_n 2.36812e-19 $X=2.395 $Y=2.125 $X2=0 $Y2=0
cc_101 N_A_84_93#_c_88_n N_A_c_195_n 7.15305e-19 $X=3.445 $Y=2.125 $X2=0 $Y2=0
cc_102 N_A_84_93#_c_80_n N_A_c_195_n 2.07958e-19 $X=3.445 $Y=0.915 $X2=0 $Y2=0
cc_103 N_A_84_93#_M1012_g N_A_c_196_n 0.00734446f $X=0.855 $Y=0.805 $X2=0 $Y2=0
cc_104 N_A_84_93#_c_86_n N_A_c_196_n 0.0947494f $X=2.395 $Y=2.125 $X2=0 $Y2=0
cc_105 N_A_84_93#_c_83_n N_A_c_196_n 5.41107e-19 $X=0.7 $Y=1.73 $X2=0 $Y2=0
cc_106 N_A_84_93#_c_91_n N_A_c_196_n 0.0245693f $X=0.82 $Y=1.73 $X2=0 $Y2=0
cc_107 N_A_84_93#_M1012_g N_B_M1000_g 0.0136624f $X=0.855 $Y=0.805 $X2=0 $Y2=0
cc_108 N_A_84_93#_c_86_n N_B_c_301_n 0.0168568f $X=2.395 $Y=2.125 $X2=0 $Y2=0
cc_109 N_A_84_93#_c_87_n N_B_c_301_n 0.00439175f $X=2.56 $Y=2.9 $X2=0 $Y2=0
cc_110 N_A_84_93#_c_86_n N_B_c_302_n 0.0107804f $X=2.395 $Y=2.125 $X2=0 $Y2=0
cc_111 N_A_84_93#_c_79_n N_B_M1007_g 0.00154695f $X=2.76 $Y=0.55 $X2=0 $Y2=0
cc_112 N_A_84_93#_c_79_n N_B_c_296_n 0.0101124f $X=2.76 $Y=0.55 $X2=0 $Y2=0
cc_113 N_A_84_93#_c_87_n N_B_c_306_n 0.0180874f $X=2.56 $Y=2.9 $X2=0 $Y2=0
cc_114 N_A_84_93#_c_88_n N_B_c_306_n 0.0180811f $X=3.445 $Y=2.125 $X2=0 $Y2=0
cc_115 N_A_84_93#_c_92_n N_B_c_306_n 0.00122348f $X=2.56 $Y=2.205 $X2=0 $Y2=0
cc_116 N_A_84_93#_c_81_n N_B_c_297_n 0.00947779f $X=2.925 $Y=0.915 $X2=0 $Y2=0
cc_117 N_A_84_93#_c_92_n N_B_c_307_n 0.00534957f $X=2.56 $Y=2.205 $X2=0 $Y2=0
cc_118 N_A_84_93#_c_81_n B 0.0133736f $X=2.925 $Y=0.915 $X2=0 $Y2=0
cc_119 N_A_84_93#_c_81_n N_B_c_299_n 0.00128556f $X=2.925 $Y=0.915 $X2=0 $Y2=0
cc_120 N_A_84_93#_M1002_g N_X_c_377_n 0.0184891f $X=0.495 $Y=0.805 $X2=0 $Y2=0
cc_121 N_A_84_93#_M1012_g N_X_c_377_n 0.00752751f $X=0.855 $Y=0.805 $X2=0 $Y2=0
cc_122 N_A_84_93#_c_83_n N_X_c_377_n 7.85225e-19 $X=0.7 $Y=1.73 $X2=0 $Y2=0
cc_123 N_A_84_93#_c_91_n N_X_c_377_n 0.0267293f $X=0.82 $Y=1.73 $X2=0 $Y2=0
cc_124 N_A_84_93#_M1002_g N_X_c_379_n 0.00358826f $X=0.495 $Y=0.805 $X2=0 $Y2=0
cc_125 N_A_84_93#_M1012_g N_X_c_379_n 0.00598504f $X=0.855 $Y=0.805 $X2=0 $Y2=0
cc_126 N_A_84_93#_M1002_g N_X_c_380_n 0.00135797f $X=0.495 $Y=0.805 $X2=0 $Y2=0
cc_127 N_A_84_93#_M1012_g N_X_c_380_n 0.012363f $X=0.855 $Y=0.805 $X2=0 $Y2=0
cc_128 N_A_84_93#_M1002_g X 0.0162943f $X=0.495 $Y=0.805 $X2=0 $Y2=0
cc_129 N_A_84_93#_M1004_g X 0.00415669f $X=0.67 $Y=2.595 $X2=0 $Y2=0
cc_130 N_A_84_93#_c_85_n X 0.00580618f $X=0.82 $Y=2.04 $X2=0 $Y2=0
cc_131 N_A_84_93#_c_147_p X 0.00153788f $X=0.905 $Y=2.125 $X2=0 $Y2=0
cc_132 N_A_84_93#_c_91_n X 0.0244853f $X=0.82 $Y=1.73 $X2=0 $Y2=0
cc_133 N_A_84_93#_M1004_g X 0.00410317f $X=0.67 $Y=2.595 $X2=0 $Y2=0
cc_134 N_A_84_93#_c_147_p X 0.0104916f $X=0.905 $Y=2.125 $X2=0 $Y2=0
cc_135 N_A_84_93#_c_83_n X 0.00577539f $X=0.7 $Y=1.73 $X2=0 $Y2=0
cc_136 N_A_84_93#_c_91_n X 0.00149385f $X=0.82 $Y=1.73 $X2=0 $Y2=0
cc_137 N_A_84_93#_M1004_g X 0.018775f $X=0.67 $Y=2.595 $X2=0 $Y2=0
cc_138 N_A_84_93#_c_86_n N_A_159_419#_M1004_d 0.00121949f $X=2.395 $Y=2.125
+ $X2=-0.19 $Y2=-0.245
cc_139 N_A_84_93#_c_147_p N_A_159_419#_M1004_d 5.75827e-19 $X=0.905 $Y=2.125
+ $X2=-0.19 $Y2=-0.245
cc_140 N_A_84_93#_c_86_n N_A_159_419#_M1005_d 0.00314508f $X=2.395 $Y=2.125
+ $X2=0 $Y2=0
cc_141 N_A_84_93#_c_86_n N_A_159_419#_c_425_n 0.0406254f $X=2.395 $Y=2.125 $X2=0
+ $Y2=0
cc_142 N_A_84_93#_M1004_g N_A_159_419#_c_426_n 0.0128526f $X=0.67 $Y=2.595 $X2=0
+ $Y2=0
cc_143 N_A_84_93#_c_86_n N_A_159_419#_c_426_n 0.0105458f $X=2.395 $Y=2.125 $X2=0
+ $Y2=0
cc_144 N_A_84_93#_c_147_p N_A_159_419#_c_426_n 0.00619993f $X=0.905 $Y=2.125
+ $X2=0 $Y2=0
cc_145 N_A_84_93#_c_83_n N_A_159_419#_c_426_n 2.33532e-19 $X=0.7 $Y=1.73 $X2=0
+ $Y2=0
cc_146 N_A_84_93#_c_86_n N_A_159_419#_c_421_n 0.021161f $X=2.395 $Y=2.125 $X2=0
+ $Y2=0
cc_147 N_A_84_93#_c_87_n N_A_159_419#_c_421_n 0.0454923f $X=2.56 $Y=2.9 $X2=0
+ $Y2=0
cc_148 N_A_84_93#_c_86_n N_VPWR_M1001_d 0.00181172f $X=2.395 $Y=2.125 $X2=-0.19
+ $Y2=-0.245
cc_149 N_A_84_93#_c_88_n N_VPWR_M1011_d 0.00865209f $X=3.445 $Y=2.125 $X2=0
+ $Y2=0
cc_150 N_A_84_93#_M1004_g N_VPWR_c_452_n 9.35833e-19 $X=0.67 $Y=2.595 $X2=0
+ $Y2=0
cc_151 N_A_84_93#_c_87_n N_VPWR_c_454_n 0.0163111f $X=2.56 $Y=2.9 $X2=0 $Y2=0
cc_152 N_A_84_93#_c_88_n N_VPWR_c_454_n 0.0144877f $X=3.445 $Y=2.125 $X2=0 $Y2=0
cc_153 N_A_84_93#_M1004_g N_VPWR_c_455_n 0.00926003f $X=0.67 $Y=2.595 $X2=0
+ $Y2=0
cc_154 N_A_84_93#_c_87_n N_VPWR_c_457_n 0.0220321f $X=2.56 $Y=2.9 $X2=0 $Y2=0
cc_155 N_A_84_93#_M1004_g N_VPWR_c_451_n 0.0168687f $X=0.67 $Y=2.595 $X2=0 $Y2=0
cc_156 N_A_84_93#_c_87_n N_VPWR_c_451_n 0.0125808f $X=2.56 $Y=2.9 $X2=0 $Y2=0
cc_157 N_A_84_93#_c_88_n A_590_412# 0.00366293f $X=3.445 $Y=2.125 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A_84_93#_M1002_g N_VGND_c_496_n 0.0122529f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_159 N_A_84_93#_M1012_g N_VGND_c_496_n 0.00100791f $X=0.855 $Y=0.805 $X2=0
+ $Y2=0
cc_160 N_A_84_93#_c_79_n N_VGND_c_497_n 0.0145731f $X=2.76 $Y=0.55 $X2=0 $Y2=0
cc_161 N_A_84_93#_c_79_n N_VGND_c_499_n 0.0110409f $X=2.76 $Y=0.55 $X2=0 $Y2=0
cc_162 N_A_84_93#_c_80_n N_VGND_c_499_n 0.0164042f $X=3.445 $Y=0.915 $X2=0 $Y2=0
cc_163 N_A_84_93#_M1002_g N_VGND_c_500_n 0.0035863f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_164 N_A_84_93#_M1012_g N_VGND_c_500_n 0.0032894f $X=0.855 $Y=0.805 $X2=0
+ $Y2=0
cc_165 N_A_84_93#_c_79_n N_VGND_c_502_n 0.0164809f $X=2.76 $Y=0.55 $X2=0 $Y2=0
cc_166 N_A_84_93#_M1002_g N_VGND_c_503_n 0.00401353f $X=0.495 $Y=0.805 $X2=0
+ $Y2=0
cc_167 N_A_84_93#_M1012_g N_VGND_c_503_n 0.00477801f $X=0.855 $Y=0.805 $X2=0
+ $Y2=0
cc_168 N_A_84_93#_c_79_n N_VGND_c_503_n 0.0121f $X=2.76 $Y=0.55 $X2=0 $Y2=0
cc_169 N_A_84_93#_c_80_n N_VGND_c_503_n 0.0150883f $X=3.445 $Y=0.915 $X2=0 $Y2=0
cc_170 N_A_c_187_n N_B_M1000_g 0.00543192f $X=1.325 $Y=1.55 $X2=0 $Y2=0
cc_171 N_A_M1006_g N_B_M1000_g 0.041275f $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_172 N_A_c_196_n N_B_M1000_g 0.00389065f $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_173 N_A_M1006_g N_B_c_292_n 0.0104164f $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_174 N_A_c_197_n N_B_c_301_n 0.0250885f $X=1.2 $Y=2.08 $X2=0 $Y2=0
cc_175 N_A_c_200_n N_B_c_302_n 0.0111922f $X=2.935 $Y=1.775 $X2=0 $Y2=0
cc_176 N_A_c_196_n N_B_c_302_n 0.00115687f $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_177 N_A_c_192_n N_B_c_303_n 0.0250885f $X=1.2 $Y=1.955 $X2=0 $Y2=0
cc_178 N_A_c_194_n N_B_c_303_n 0.0192159f $X=1.735 $Y=1.46 $X2=0 $Y2=0
cc_179 N_A_c_196_n N_B_c_303_n 0.0068601f $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_180 N_A_M1006_g N_B_M1007_g 0.0132889f $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_181 N_A_M1011_g N_B_c_295_n 0.00307129f $X=3.285 $Y=2.56 $X2=0 $Y2=0
cc_182 N_A_c_200_n N_B_c_295_n 0.00847177f $X=2.935 $Y=1.775 $X2=0 $Y2=0
cc_183 N_A_c_193_n N_B_c_295_n 0.00332237f $X=3.1 $Y=1.345 $X2=0 $Y2=0
cc_184 N_A_c_196_n N_B_c_295_n 0.00211629f $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_185 N_A_M1011_g N_B_c_305_n 0.0890886f $X=3.285 $Y=2.56 $X2=0 $Y2=0
cc_186 N_A_c_200_n N_B_c_305_n 0.0143817f $X=2.935 $Y=1.775 $X2=0 $Y2=0
cc_187 N_A_c_195_n N_B_c_305_n 0.00188854f $X=3.335 $Y=1.345 $X2=0 $Y2=0
cc_188 N_A_M1008_g N_B_c_296_n 0.0216025f $X=2.975 $Y=0.55 $X2=0 $Y2=0
cc_189 N_A_c_200_n N_B_c_307_n 0.00164963f $X=2.935 $Y=1.775 $X2=0 $Y2=0
cc_190 N_A_M1006_g B 5.76577e-19 $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_191 N_A_c_200_n B 0.0334701f $X=2.935 $Y=1.775 $X2=0 $Y2=0
cc_192 N_A_c_193_n B 0.0256788f $X=3.1 $Y=1.345 $X2=0 $Y2=0
cc_193 N_A_c_194_n B 2.64371e-19 $X=1.735 $Y=1.46 $X2=0 $Y2=0
cc_194 N_A_c_195_n B 0.00252696f $X=3.335 $Y=1.345 $X2=0 $Y2=0
cc_195 N_A_c_196_n B 0.00891413f $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_196 N_A_M1006_g N_B_c_299_n 0.00476118f $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_197 N_A_c_193_n N_B_c_299_n 3.14114e-19 $X=3.1 $Y=1.345 $X2=0 $Y2=0
cc_198 N_A_c_194_n N_B_c_299_n 0.00934542f $X=1.735 $Y=1.46 $X2=0 $Y2=0
cc_199 N_A_c_195_n N_B_c_299_n 0.0216025f $X=3.335 $Y=1.345 $X2=0 $Y2=0
cc_200 N_A_c_196_n N_B_c_299_n 2.63338e-19 $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_201 N_A_c_200_n N_B_c_300_n 0.00137043f $X=2.935 $Y=1.775 $X2=0 $Y2=0
cc_202 N_A_c_196_n N_B_c_300_n 6.63365e-19 $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_203 N_A_M1006_g N_X_c_377_n 3.72893e-19 $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_204 N_A_c_196_n N_X_c_377_n 0.007597f $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_205 N_A_M1006_g N_X_c_379_n 4.43984e-19 $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_206 N_A_M1006_g N_X_c_380_n 0.00184703f $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_207 N_A_c_196_n N_X_c_380_n 0.00981319f $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_208 N_A_c_197_n X 7.66595e-19 $X=1.2 $Y=2.08 $X2=0 $Y2=0
cc_209 N_A_c_197_n N_A_159_419#_c_425_n 0.0133988f $X=1.2 $Y=2.08 $X2=0 $Y2=0
cc_210 N_A_c_197_n N_A_159_419#_c_426_n 0.010006f $X=1.2 $Y=2.08 $X2=0 $Y2=0
cc_211 N_A_c_197_n N_A_159_419#_c_421_n 7.5175e-19 $X=1.2 $Y=2.08 $X2=0 $Y2=0
cc_212 N_A_c_197_n N_VPWR_c_452_n 0.0113662f $X=1.2 $Y=2.08 $X2=0 $Y2=0
cc_213 N_A_M1011_g N_VPWR_c_454_n 0.0206572f $X=3.285 $Y=2.56 $X2=0 $Y2=0
cc_214 N_A_c_197_n N_VPWR_c_455_n 0.00840199f $X=1.2 $Y=2.08 $X2=0 $Y2=0
cc_215 N_A_M1011_g N_VPWR_c_457_n 0.00823892f $X=3.285 $Y=2.56 $X2=0 $Y2=0
cc_216 N_A_c_197_n N_VPWR_c_451_n 0.0073633f $X=1.2 $Y=2.08 $X2=0 $Y2=0
cc_217 N_A_M1011_g N_VPWR_c_451_n 0.0142593f $X=3.285 $Y=2.56 $X2=0 $Y2=0
cc_218 N_A_M1006_g N_VGND_c_497_n 0.00434651f $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_219 N_A_c_194_n N_VGND_c_497_n 0.00229259f $X=1.735 $Y=1.46 $X2=0 $Y2=0
cc_220 N_A_c_196_n N_VGND_c_497_n 0.00446503f $X=1.9 $Y=1.577 $X2=0 $Y2=0
cc_221 N_A_M1008_g N_VGND_c_499_n 0.0015698f $X=2.975 $Y=0.55 $X2=0 $Y2=0
cc_222 N_A_M1009_g N_VGND_c_499_n 0.010742f $X=3.335 $Y=0.55 $X2=0 $Y2=0
cc_223 N_A_M1008_g N_VGND_c_502_n 0.00457319f $X=2.975 $Y=0.55 $X2=0 $Y2=0
cc_224 N_A_M1009_g N_VGND_c_502_n 0.0040395f $X=3.335 $Y=0.55 $X2=0 $Y2=0
cc_225 N_A_M1006_g N_VGND_c_503_n 9.39239e-19 $X=1.645 $Y=0.805 $X2=0 $Y2=0
cc_226 N_A_M1008_g N_VGND_c_503_n 0.00493169f $X=2.975 $Y=0.55 $X2=0 $Y2=0
cc_227 N_A_M1009_g N_VGND_c_503_n 0.00396826f $X=3.335 $Y=0.55 $X2=0 $Y2=0
cc_228 N_B_M1000_g N_X_c_379_n 6.59698e-19 $X=1.285 $Y=0.805 $X2=0 $Y2=0
cc_229 N_B_M1000_g N_X_c_380_n 0.00969965f $X=1.285 $Y=0.805 $X2=0 $Y2=0
cc_230 N_B_c_301_n N_A_159_419#_c_425_n 0.0133988f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_231 N_B_c_301_n N_A_159_419#_c_426_n 7.5175e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_232 N_B_c_301_n N_A_159_419#_c_421_n 0.010006f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_233 N_B_c_306_n N_A_159_419#_c_421_n 8.95699e-19 $X=2.825 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_B_c_301_n N_VPWR_c_452_n 0.0120984f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_235 N_B_c_306_n N_VPWR_c_454_n 0.00260219f $X=2.825 $Y=1.985 $X2=0 $Y2=0
cc_236 N_B_c_301_n N_VPWR_c_457_n 0.00840199f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_237 N_B_c_306_n N_VPWR_c_457_n 0.00883132f $X=2.825 $Y=1.985 $X2=0 $Y2=0
cc_238 N_B_c_301_n N_VPWR_c_451_n 0.00865707f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_239 N_B_c_306_n N_VPWR_c_451_n 0.0168579f $X=2.825 $Y=1.985 $X2=0 $Y2=0
cc_240 N_B_M1000_g N_VGND_c_497_n 0.00478595f $X=1.285 $Y=0.805 $X2=0 $Y2=0
cc_241 N_B_c_292_n N_VGND_c_497_n 0.02199f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_242 N_B_M1007_g N_VGND_c_497_n 0.0119975f $X=2.155 $Y=0.55 $X2=0 $Y2=0
cc_243 N_B_c_296_n N_VGND_c_497_n 0.00195521f $X=2.545 $Y=0.835 $X2=0 $Y2=0
cc_244 N_B_c_293_n N_VGND_c_500_n 0.0205169f $X=1.36 $Y=0.18 $X2=0 $Y2=0
cc_245 N_B_c_292_n N_VGND_c_502_n 0.00486043f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_246 N_B_c_296_n N_VGND_c_502_n 0.00457319f $X=2.545 $Y=0.835 $X2=0 $Y2=0
cc_247 N_B_c_292_n N_VGND_c_503_n 0.029163f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_248 N_B_c_293_n N_VGND_c_503_n 0.0107545f $X=1.36 $Y=0.18 $X2=0 $Y2=0
cc_249 N_B_c_296_n N_VGND_c_503_n 0.00872815f $X=2.545 $Y=0.835 $X2=0 $Y2=0
cc_250 N_B_c_297_n N_VGND_c_503_n 0.0015396f $X=2.545 $Y=0.91 $X2=0 $Y2=0
cc_251 X N_A_159_419#_c_426_n 0.0434813f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_252 X N_VPWR_c_455_n 0.026532f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_253 N_X_M1004_s N_VPWR_c_451_n 0.00244761f $X=0.245 $Y=2.095 $X2=0 $Y2=0
cc_254 X N_VPWR_c_451_n 0.0164464f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_255 N_X_c_377_n N_VGND_c_496_n 0.00698135f $X=0.735 $Y=1.3 $X2=0 $Y2=0
cc_256 N_X_c_378_n N_VGND_c_496_n 0.0206891f $X=0.355 $Y=1.3 $X2=0 $Y2=0
cc_257 N_X_c_380_n N_VGND_c_496_n 0.0123476f $X=1.07 $Y=0.805 $X2=0 $Y2=0
cc_258 N_X_c_380_n N_VGND_c_497_n 0.00349948f $X=1.07 $Y=0.805 $X2=0 $Y2=0
cc_259 N_X_c_380_n N_VGND_c_500_n 0.010776f $X=1.07 $Y=0.805 $X2=0 $Y2=0
cc_260 N_X_c_380_n N_VGND_c_503_n 0.0152747f $X=1.07 $Y=0.805 $X2=0 $Y2=0
cc_261 N_A_159_419#_c_425_n N_VPWR_M1001_d 0.00358238f $X=1.83 $Y=2.475
+ $X2=-0.19 $Y2=1.655
cc_262 N_A_159_419#_c_425_n N_VPWR_c_452_n 0.0157965f $X=1.83 $Y=2.475 $X2=0
+ $Y2=0
cc_263 N_A_159_419#_c_426_n N_VPWR_c_452_n 0.0214145f $X=0.935 $Y=2.555 $X2=0
+ $Y2=0
cc_264 N_A_159_419#_c_421_n N_VPWR_c_452_n 0.0214145f $X=1.995 $Y=2.555 $X2=0
+ $Y2=0
cc_265 N_A_159_419#_c_426_n N_VPWR_c_455_n 0.0177877f $X=0.935 $Y=2.555 $X2=0
+ $Y2=0
cc_266 N_A_159_419#_c_421_n N_VPWR_c_457_n 0.0197484f $X=1.995 $Y=2.555 $X2=0
+ $Y2=0
cc_267 N_A_159_419#_M1004_d N_VPWR_c_451_n 0.00223819f $X=0.795 $Y=2.095 $X2=0
+ $Y2=0
cc_268 N_A_159_419#_M1005_d N_VPWR_c_451_n 0.0023218f $X=1.855 $Y=2.095 $X2=0
+ $Y2=0
cc_269 N_A_159_419#_c_425_n N_VPWR_c_451_n 0.0130057f $X=1.83 $Y=2.475 $X2=0
+ $Y2=0
cc_270 N_A_159_419#_c_426_n N_VPWR_c_451_n 0.0123222f $X=0.935 $Y=2.555 $X2=0
+ $Y2=0
cc_271 N_A_159_419#_c_421_n N_VPWR_c_451_n 0.0125055f $X=1.995 $Y=2.555 $X2=0
+ $Y2=0
