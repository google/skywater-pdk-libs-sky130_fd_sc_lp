* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__maj3_0 A B C VGND VNB VPB VPWR X
X0 a_477_57# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND a_28_431# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_313_57# B a_28_431# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR A a_319_431# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_28_431# C a_149_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_28_431# B a_477_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_149_57# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_28_431# B a_477_431# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_477_431# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_319_431# B a_28_431# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR a_28_431# X VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VGND A a_313_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_115_431# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_28_431# C a_115_431# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
