* File: sky130_fd_sc_lp__ebufn_4.pex.spice
* Created: Fri Aug 28 10:31:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EBUFN_4%A_84_21# 1 2 9 13 17 21 25 29 33 37 39 44 45
+ 46 47 48 54 55 56 57 61 65 70 73 78 79 81
c162 70 0 1.17434e-19 $X=1.72 $Y=1.48
c163 55 0 9.69886e-20 $X=4.325 $Y=2.1
c164 54 0 1.77381e-19 $X=2.13 $Y=2.015
r165 79 81 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=6.06 $Y=1.95
+ $X2=6.06 $Y2=1.135
r166 78 79 8.80985 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=5.927 $Y=2.115
+ $X2=5.927 $Y2=1.95
r167 73 75 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.41 $Y=2.1
+ $X2=4.41 $Y2=2.27
r168 70 72 22.4305 $w=2.23e-07 $l=4.1e-07 $layer=LI1_cond $X=1.72 $Y=1.48
+ $X2=2.13 $Y2=1.48
r169 70 71 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.48 $X2=1.72 $Y2=1.48
r170 63 81 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=5.962 $Y=0.953
+ $X2=5.962 $Y2=1.135
r171 63 65 16.8288 $w=3.63e-07 $l=5.33e-07 $layer=LI1_cond $X=5.962 $Y=0.953
+ $X2=5.962 $Y2=0.42
r172 59 61 14.7036 $w=4.33e-07 $l=5.55e-07 $layer=LI1_cond $X=5.927 $Y=2.355
+ $X2=5.927 $Y2=2.91
r173 58 75 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=2.27
+ $X2=4.41 $Y2=2.27
r174 57 59 2.2519 $w=4.33e-07 $l=8.5e-08 $layer=LI1_cond $X=5.927 $Y=2.27
+ $X2=5.927 $Y2=2.355
r175 57 78 4.10641 $w=4.33e-07 $l=1.55e-07 $layer=LI1_cond $X=5.927 $Y=2.27
+ $X2=5.927 $Y2=2.115
r176 57 58 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=5.71 $Y=2.27
+ $X2=4.495 $Y2=2.27
r177 55 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.325 $Y=2.1
+ $X2=4.41 $Y2=2.1
r178 55 56 137.658 $w=1.68e-07 $l=2.11e-06 $layer=LI1_cond $X=4.325 $Y=2.1
+ $X2=2.215 $Y2=2.1
r179 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=2.015
+ $X2=2.215 $Y2=2.1
r180 53 72 2.32876 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.13 $Y=1.645
+ $X2=2.13 $Y2=1.48
r181 53 54 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.13 $Y=1.645
+ $X2=2.13 $Y2=2.015
r182 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.48 $X2=1.04 $Y2=1.48
r183 48 70 1.28872 $w=3.3e-07 $l=1.31364e-07 $layer=LI1_cond $X=1.72 $Y=1.48
+ $X2=1.72 $Y2=1.48
r184 48 50 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.72 $Y=1.48
+ $X2=1.04 $Y2=1.48
r185 46 71 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.85 $Y=1.48
+ $X2=1.72 $Y2=1.48
r186 46 47 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.85 $Y=1.48
+ $X2=1.925 $Y2=1.48
r187 44 51 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=1.35 $Y=1.48
+ $X2=1.04 $Y2=1.48
r188 44 45 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.35 $Y=1.48
+ $X2=1.425 $Y2=1.48
r189 43 71 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.5 $Y=1.48
+ $X2=1.72 $Y2=1.48
r190 43 45 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.5 $Y=1.48
+ $X2=1.425 $Y2=1.48
r191 40 42 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.925 $Y2=1.48
r192 39 51 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1 $Y=1.48 $X2=1.04
+ $Y2=1.48
r193 39 42 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1 $Y=1.48 $X2=0.925
+ $Y2=1.48
r194 35 47 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.645
+ $X2=1.925 $Y2=1.48
r195 35 37 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.925 $Y=1.645
+ $X2=1.925 $Y2=2.465
r196 31 47 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.315
+ $X2=1.925 $Y2=1.48
r197 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.925 $Y=1.315
+ $X2=1.925 $Y2=0.655
r198 27 45 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.645
+ $X2=1.425 $Y2=1.48
r199 27 29 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.425 $Y=1.645
+ $X2=1.425 $Y2=2.465
r200 23 45 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.315
+ $X2=1.425 $Y2=1.48
r201 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.425 $Y=1.315
+ $X2=1.425 $Y2=0.655
r202 19 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.645
+ $X2=0.925 $Y2=1.48
r203 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.925 $Y=1.645
+ $X2=0.925 $Y2=2.465
r204 15 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.315
+ $X2=0.925 $Y2=1.48
r205 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.925 $Y=1.315
+ $X2=0.925 $Y2=0.655
r206 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.645
+ $X2=0.495 $Y2=1.48
r207 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.495 $Y=1.645
+ $X2=0.495 $Y2=2.465
r208 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.315
+ $X2=0.495 $Y2=1.48
r209 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.315
+ $X2=0.495 $Y2=0.655
r210 2 78 400 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.835 $X2=5.875 $Y2=2.115
r211 2 61 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.835 $X2=5.875 $Y2=2.91
r212 1 65 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.805
+ $Y=0.275 $X2=5.945 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_4%A_456_21# 1 2 7 9 10 11 12 14 15 17 19 20 22
+ 24 25 28 29 30 31 33 34 39 42 44
c109 39 0 7.68297e-20 $X=5.025 $Y=1.765
c110 25 0 1.4047e-19 $X=4.08 $Y=1.26
c111 11 0 1.17434e-19 $X=2.43 $Y=1.26
c112 7 0 5.58653e-20 $X=2.355 $Y=1.185
r113 44 45 1.39429 $w=7e-07 $l=8e-08 $layer=LI1_cond $X=4.945 $Y=0.632 $X2=5.025
+ $Y2=0.632
r114 41 44 10.1957 $w=7e-07 $l=5.85e-07 $layer=LI1_cond $X=4.36 $Y=0.632
+ $X2=4.945 $Y2=0.632
r115 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.36
+ $Y=0.505 $X2=4.36 $Y2=0.505
r116 38 45 9.32152 $w=1.7e-07 $l=3.78e-07 $layer=LI1_cond $X=5.025 $Y=1.01
+ $X2=5.025 $Y2=0.632
r117 38 39 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=5.025 $Y=1.01
+ $X2=5.025 $Y2=1.765
r118 34 39 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.94 $Y=1.89
+ $X2=5.025 $Y2=1.765
r119 34 36 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=4.94 $Y=1.89
+ $X2=4.83 $Y2=1.89
r120 32 42 35.3689 $w=4.45e-07 $l=2.83e-07 $layer=POLY_cond $X=4.302 $Y=0.788
+ $X2=4.302 $Y2=0.505
r121 32 33 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=4.302 $Y=0.788
+ $X2=4.302 $Y2=1.01
r122 28 33 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.155 $Y=1.185
+ $X2=4.155 $Y2=1.01
r123 26 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.72 $Y=1.26
+ $X2=3.645 $Y2=1.26
r124 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.08 $Y=1.26
+ $X2=4.155 $Y2=1.185
r125 25 26 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.08 $Y=1.26
+ $X2=3.72 $Y2=1.26
r126 22 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.645 $Y=1.185
+ $X2=3.645 $Y2=1.26
r127 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.645 $Y=1.185
+ $X2=3.645 $Y2=0.655
r128 21 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.29 $Y=1.26
+ $X2=3.215 $Y2=1.26
r129 20 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.57 $Y=1.26
+ $X2=3.645 $Y2=1.26
r130 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.57 $Y=1.26
+ $X2=3.29 $Y2=1.26
r131 17 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.215 $Y=1.185
+ $X2=3.215 $Y2=1.26
r132 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.215 $Y=1.185
+ $X2=3.215 $Y2=0.655
r133 16 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.86 $Y=1.26
+ $X2=2.785 $Y2=1.26
r134 15 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.14 $Y=1.26
+ $X2=3.215 $Y2=1.26
r135 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.14 $Y=1.26
+ $X2=2.86 $Y2=1.26
r136 12 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.785 $Y=1.185
+ $X2=2.785 $Y2=1.26
r137 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.785 $Y=1.185
+ $X2=2.785 $Y2=0.655
r138 10 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.71 $Y=1.26
+ $X2=2.785 $Y2=1.26
r139 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.71 $Y=1.26
+ $X2=2.43 $Y2=1.26
r140 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.43 $Y2=1.26
r141 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=0.655
r142 2 36 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.685
+ $Y=1.785 $X2=4.83 $Y2=1.93
r143 1 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.8
+ $Y=0.275 $X2=4.945 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_4%TE_B 1 3 4 5 6 8 9 11 13 14 16 18 19 21 25
+ 29 31 32 33 34 35 36 37 41 48
c132 37 0 4.34819e-20 $X=4.56 $Y=1.295
r133 44 46 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.605 $Y=1.43
+ $X2=4.605 $Y2=1.62
r134 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.605
+ $Y=1.43 $X2=4.605 $Y2=1.43
r135 41 44 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.605 $Y=1.34
+ $X2=4.605 $Y2=1.43
r136 37 45 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.605 $Y=1.295
+ $X2=4.605 $Y2=1.43
r137 37 48 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=1.295
+ $X2=4.44 $Y2=1.295
r138 36 48 18.0382 $w=2.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.08 $Y=1.295
+ $X2=4.44 $Y2=1.295
r139 35 36 24.051 $w=2.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.295
+ $X2=4.08 $Y2=1.295
r140 27 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.16 $Y=1.415
+ $X2=5.16 $Y2=1.34
r141 27 29 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=5.16 $Y=1.415
+ $X2=5.16 $Y2=2.465
r142 23 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.16 $Y=1.265
+ $X2=5.16 $Y2=1.34
r143 23 25 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.16 $Y=1.265
+ $X2=5.16 $Y2=0.695
r144 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.34
+ $X2=4.605 $Y2=1.34
r145 21 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.085 $Y=1.34
+ $X2=5.16 $Y2=1.34
r146 21 22 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=5.085 $Y=1.34
+ $X2=4.77 $Y2=1.34
r147 20 33 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=4.11 $Y=1.62
+ $X2=4.035 $Y2=1.635
r148 19 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.44 $Y=1.62
+ $X2=4.605 $Y2=1.62
r149 19 20 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.44 $Y=1.62
+ $X2=4.11 $Y2=1.62
r150 16 33 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.035 $Y=1.725
+ $X2=4.035 $Y2=1.635
r151 16 18 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.035 $Y=1.725
+ $X2=4.035 $Y2=2.465
r152 15 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.5 $Y=1.65
+ $X2=3.425 $Y2=1.65
r153 14 33 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=3.96 $Y=1.65
+ $X2=4.035 $Y2=1.635
r154 14 15 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.96 $Y=1.65
+ $X2=3.5 $Y2=1.65
r155 11 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.425 $Y=1.725
+ $X2=3.425 $Y2=1.65
r156 11 13 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.425 $Y=1.725
+ $X2=3.425 $Y2=2.465
r157 10 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.07 $Y=1.65
+ $X2=2.995 $Y2=1.65
r158 9 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.35 $Y=1.65
+ $X2=3.425 $Y2=1.65
r159 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.35 $Y=1.65
+ $X2=3.07 $Y2=1.65
r160 6 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.995 $Y=1.725
+ $X2=2.995 $Y2=1.65
r161 6 8 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.995 $Y=1.725
+ $X2=2.995 $Y2=2.465
r162 4 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.92 $Y=1.65
+ $X2=2.995 $Y2=1.65
r163 4 5 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.92 $Y=1.65 $X2=2.5
+ $Y2=1.65
r164 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.425 $Y=1.725
+ $X2=2.5 $Y2=1.65
r165 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.425 $Y=1.725
+ $X2=2.425 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_4%A 3 7 9 12 13
c36 3 0 7.68297e-20 $X=5.66 $Y=2.465
r37 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.64 $Y=1.51
+ $X2=5.64 $Y2=1.675
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.64 $Y=1.51
+ $X2=5.64 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=1.51 $X2=5.64 $Y2=1.51
r40 9 13 4.46572 $w=3.98e-07 $l=1.55e-07 $layer=LI1_cond $X=5.605 $Y=1.665
+ $X2=5.605 $Y2=1.51
r41 7 14 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=5.73 $Y=0.695
+ $X2=5.73 $Y2=1.345
r42 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.66 $Y=2.465
+ $X2=5.66 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_4%A_27_367# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 34 38 43 46 50
r76 49 50 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.21 $Y=2.52 $X2=3.21
+ $Y2=2.61
r77 46 49 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.21 $Y=2.44 $X2=3.21
+ $Y2=2.52
r78 36 38 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.25 $Y=2.695
+ $X2=4.25 $Y2=2.8
r79 35 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=2.61
+ $X2=3.21 $Y2=2.61
r80 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.085 $Y=2.61
+ $X2=4.25 $Y2=2.695
r81 34 35 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.085 $Y=2.61
+ $X2=3.375 $Y2=2.61
r82 31 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=2.44
+ $X2=2.21 $Y2=2.44
r83 30 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=2.44
+ $X2=3.21 $Y2=2.44
r84 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.045 $Y=2.44
+ $X2=2.375 $Y2=2.44
r85 28 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=2.525 $X2=2.21
+ $Y2=2.44
r86 28 29 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.21 $Y=2.525
+ $X2=2.21 $Y2=2.905
r87 27 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=2.99
+ $X2=1.21 $Y2=2.99
r88 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=2.21 $Y2=2.905
r89 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=1.375 $Y2=2.99
r90 22 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=2.905
+ $X2=1.21 $Y2=2.99
r91 22 24 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.21 $Y=2.905
+ $X2=1.21 $Y2=2.24
r92 21 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.99
+ $X2=0.24 $Y2=2.99
r93 20 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=2.99
+ $X2=1.21 $Y2=2.99
r94 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=2.99
+ $X2=0.365 $Y2=2.99
r95 16 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.905
+ $X2=0.24 $Y2=2.99
r96 16 18 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=0.24 $Y=2.905
+ $X2=0.24 $Y2=1.98
r97 5 38 600 $w=1.7e-07 $l=1.03263e-06 $layer=licon1_PDIFF $count=1 $X=4.11
+ $Y=1.835 $X2=4.25 $Y2=2.8
r98 4 49 300 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_PDIFF $count=2 $X=3.07
+ $Y=1.835 $X2=3.21 $Y2=2.52
r99 3 45 300 $w=1.7e-07 $l=7.82991e-07 $layer=licon1_PDIFF $count=2 $X=2
+ $Y=1.835 $X2=2.21 $Y2=2.52
r100 2 43 400 $w=1.7e-07 $l=1.21547e-06 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.21 $Y2=2.95
r101 2 24 400 $w=1.7e-07 $l=4.99074e-07 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.21 $Y2=2.24
r102 1 41 400 $w=1.7e-07 $l=1.14521e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=2.91
r103 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_4%Z 1 2 3 4 15 17 18 21 23 27 33 35 37 38
c65 21 0 5.58653e-20 $X=1.545 $Y=1.06
c66 18 0 9.44575e-20 $X=0.62 $Y=1.815
r67 33 38 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=1.295
+ $X2=0.24 $Y2=1.295
r68 32 33 0.873046 $w=2.3e-07 $l=1.7e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.535 $Y2=1.295
r69 31 32 12.1483 $w=2.36e-07 $l=2.35e-07 $layer=LI1_cond $X=0.705 $Y=1.06
+ $X2=0.705 $Y2=1.295
r70 25 27 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.71 $Y=0.975
+ $X2=1.71 $Y2=0.805
r71 24 35 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.875 $Y=1.9
+ $X2=0.705 $Y2=1.9
r72 23 37 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.9
+ $X2=1.71 $Y2=1.9
r73 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.545 $Y=1.9
+ $X2=0.875 $Y2=1.9
r74 22 31 2.65936 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.875 $Y=1.06
+ $X2=0.705 $Y2=1.06
r75 21 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.545 $Y=1.06
+ $X2=1.71 $Y2=0.975
r76 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.545 $Y=1.06
+ $X2=0.875 $Y2=1.06
r77 18 35 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.62 $Y=1.815
+ $X2=0.705 $Y2=1.9
r78 17 32 6.91891 $w=2.36e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.62 $Y=1.41
+ $X2=0.705 $Y2=1.295
r79 17 18 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.62 $Y=1.41
+ $X2=0.62 $Y2=1.815
r80 13 31 4.20344 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.975
+ $X2=0.705 $Y2=1.06
r81 13 15 5.76222 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.705 $Y=0.975
+ $X2=0.705 $Y2=0.805
r82 4 37 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.835 $X2=1.71 $Y2=1.98
r83 3 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=1.98
r84 2 27 182 $w=1.7e-07 $l=6.66783e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.235 $X2=1.71 $Y2=0.805
r85 1 15 182 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_4%VPWR 1 2 3 12 14 18 22 25 26 27 29 45 46 49
+ 52
r74 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r75 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r76 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r77 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r78 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r79 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r80 40 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r81 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=5.04
+ $Y2=3.33
r82 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r83 37 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.71 $Y2=3.33
r84 37 39 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.08 $Y2=3.33
r85 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r86 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r87 32 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r88 31 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r89 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r90 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.71 $Y2=3.33
r91 29 35 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.16 $Y2=3.33
r92 27 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r93 27 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 25 42 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.375 $Y2=3.33
r96 24 45 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.54 $Y=3.33 $X2=6
+ $Y2=3.33
r97 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=3.33
+ $X2=5.375 $Y2=3.33
r98 20 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=3.245
+ $X2=5.375 $Y2=3.33
r99 20 22 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=5.375 $Y=3.245
+ $X2=5.375 $Y2=2.82
r100 16 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=3.33
r101 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=2.95
r102 15 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=2.71 $Y2=3.33
r103 14 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=3.71 $Y2=3.33
r104 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=2.875 $Y2=3.33
r105 10 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=3.245
+ $X2=2.71 $Y2=3.33
r106 10 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.71 $Y=3.245
+ $X2=2.71 $Y2=2.905
r107 3 22 600 $w=1.7e-07 $l=1.05268e-06 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.835 $X2=5.375 $Y2=2.82
r108 2 18 600 $w=1.7e-07 $l=1.21547e-06 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.835 $X2=3.71 $Y2=2.95
r109 1 12 600 $w=1.7e-07 $l=1.1703e-06 $layer=licon1_PDIFF $count=1 $X=2.5
+ $Y=1.835 $X2=2.71 $Y2=2.905
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_4%A_27_47# 1 2 3 4 5 18 22 24 25 26 27 30 32
+ 36 39 41 45
r75 45 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3 $Y=0.925 $X2=3
+ $Y2=1.22
r76 34 36 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=3.86 $Y=0.84
+ $X2=3.86 $Y2=0.42
r77 33 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.925 $X2=3
+ $Y2=0.925
r78 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.695 $Y=0.925
+ $X2=3.86 $Y2=0.84
r79 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.695 $Y=0.925
+ $X2=3.085 $Y2=0.925
r80 28 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=0.84 $X2=3
+ $Y2=0.925
r81 28 30 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3 $Y=0.84 $X2=3
+ $Y2=0.42
r82 26 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=1.22 $X2=3
+ $Y2=1.22
r83 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.915 $Y=1.22
+ $X2=2.225 $Y2=1.22
r84 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=1.135
+ $X2=2.225 $Y2=1.22
r85 24 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.34
r86 24 25 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=1.135
r87 23 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.34
+ $X2=1.21 $Y2=0.34
r88 22 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.34
+ $X2=2.14 $Y2=0.34
r89 22 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.055 $Y=0.34
+ $X2=1.375 $Y2=0.34
r90 19 39 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=0.34
+ $X2=0.24 $Y2=0.34
r91 18 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.21 $Y2=0.34
r92 18 19 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.365 $Y2=0.34
r93 5 36 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.72
+ $Y=0.235 $X2=3.86 $Y2=0.42
r94 4 45 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=2.86
+ $Y=0.235 $X2=3 $Y2=0.93
r95 4 30 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.86
+ $Y=0.235 $X2=3 $Y2=0.42
r96 3 43 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.235
+ $X2=2.14 $Y2=0.42
r97 2 41 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.235
+ $X2=1.21 $Y2=0.38
r98 1 39 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_4%VGND 1 2 3 12 16 20 23 24 25 27 39 48 49 52
+ 55
r77 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r78 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r79 49 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r80 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r81 46 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.445
+ $Y2=0
r82 46 48 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=6
+ $Y2=0
r83 45 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r84 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r85 42 45 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r86 41 44 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r87 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r88 39 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.28 $Y=0 $X2=5.445
+ $Y2=0
r89 39 44 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.28 $Y=0 $X2=5.04
+ $Y2=0
r90 35 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.57
+ $Y2=0
r91 35 37 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=3.12
+ $Y2=0
r92 34 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r93 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r94 30 34 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r95 29 33 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r96 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r97 27 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.57
+ $Y2=0
r98 27 33 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.16
+ $Y2=0
r99 25 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r100 25 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r101 25 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r102 23 37 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=0
+ $X2=3.12 $Y2=0
r103 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.39
+ $Y2=0
r104 22 41 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.6
+ $Y2=0
r105 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.39
+ $Y2=0
r106 18 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=0.085
+ $X2=5.445 $Y2=0
r107 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.445 $Y=0.085
+ $X2=5.445 $Y2=0.42
r108 14 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.39 $Y2=0
r109 14 16 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.39 $Y2=0.44
r110 10 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=0.085
+ $X2=2.57 $Y2=0
r111 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.57 $Y=0.085
+ $X2=2.57 $Y2=0.38
r112 3 20 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.235
+ $Y=0.275 $X2=5.445 $Y2=0.42
r113 2 16 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.235 $X2=3.43 $Y2=0.44
r114 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.43
+ $Y=0.235 $X2=2.57 $Y2=0.38
.ends

