* File: sky130_fd_sc_lp__a41o_4.spice
* Created: Wed Sep  2 09:29:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41o_4.pex.spice"
.subckt sky130_fd_sc_lp__a41o_4  VNB VPB B1 A1 A2 A3 A4 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_100_23#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_100_23#_M1004_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1004_d N_A_100_23#_M1016_g N_X_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1024_d N_A_100_23#_M1024_g N_X_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1013 N_A_100_23#_M1013_d N_B1_M1013_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1022 N_A_100_23#_M1013_d N_B1_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1017 N_A_667_47#_M1017_d N_A1_M1017_g N_A_100_23#_M1017_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1025 N_A_667_47#_M1025_d N_A1_M1025_g N_A_100_23#_M1017_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1003 N_A_667_47#_M1025_d N_A2_M1003_g N_A_922_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1018 N_A_667_47#_M1018_d N_A2_M1018_g N_A_922_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_A_1115_47#_M1011_d N_A3_M1011_g N_A_922_47#_M1011_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1026 N_A_1115_47#_M1026_d N_A3_M1026_g N_A_922_47#_M1011_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1009 N_A_1115_47#_M1026_d N_A4_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1019 N_A_1115_47#_M1019_d N_A4_M1019_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_X_M1000_d N_A_100_23#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_X_M1000_d N_A_100_23#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1015 N_X_M1015_d N_A_100_23#_M1015_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1020 N_X_M1015_d N_A_100_23#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1007 N_A_100_23#_M1007_d N_B1_M1007_g N_A_495_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1023 N_A_100_23#_M1007_d N_B1_M1023_g N_A_495_367#_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1001 N_A_495_367#_M1023_s N_A1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1012 N_A_495_367#_M1012_d N_A1_M1012_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_495_367#_M1012_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.20475 AS=0.1764 PD=1.585 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1027 N_VPWR_M1008_d N_A2_M1027_g N_A_495_367#_M1027_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.20475 AS=0.1764 PD=1.585 PS=1.54 NRD=3.9006 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1005 N_A_495_367#_M1027_s N_A3_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1014 N_A_495_367#_M1014_d N_A3_M1014_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1010 N_A_495_367#_M1014_d N_A4_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1021 N_A_495_367#_M1021_d N_A4_M1021_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.0319 P=19.85
*
.include "sky130_fd_sc_lp__a41o_4.pxi.spice"
*
.ends
*
*
