* File: sky130_fd_sc_lp__fahcin_1.spice
* Created: Fri Aug 28 10:35:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__fahcin_1.pex.spice"
.subckt sky130_fd_sc_lp__fahcin_1  VNB VPB A B CIN VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CIN	CIN
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_A_M1016_g N_A_29_47#_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.232135 AS=0.2394 PD=1.57784 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1005 N_A_256_87#_M1005_d N_A_29_47#_M1005_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1728 AS=0.176865 PD=1.82 PS=1.20216 NRD=0 NRS=51.552 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1026 N_A_29_47#_M1026_d N_A_439_47#_M1026_g N_A_364_73#_M1026_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.37515 PD=0.92 PS=3.05 NRD=0 NRS=99.588 M=1
+ R=4.26667 SA=75000.3 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1006 N_A_555_73#_M1006_d N_B_M1006_g N_A_29_47#_M1026_d VNB NSHORT L=0.15
+ W=0.64 AD=0.17405 AS=0.0896 PD=1.45 PS=0.92 NRD=50.616 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001 A=0.096 P=1.58 MULT=1
MM1009 N_A_256_87#_M1009_d N_A_439_47#_M1009_g N_A_555_73#_M1006_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1744 AS=0.17405 PD=1.185 PS=1.45 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1000 N_A_364_73#_M1000_d N_B_M1000_g N_A_256_87#_M1009_d VNB NSHORT L=0.15
+ W=0.64 AD=0.176 AS=0.1744 PD=1.83 PS=1.185 NRD=0.936 NRS=49.68 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_A_439_47#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.244849 AS=0.231 PD=1.58919 PS=2.23 NRD=11.424 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1015 N_A_1152_389#_M1015_d N_A_439_47#_M1015_g N_VGND_M1004_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.186551 PD=0.92 PS=1.21081 NRD=0 NRS=37.5 M=1
+ R=4.26667 SA=75000.9 SB=75004.6 A=0.096 P=1.58 MULT=1
MM1027 N_COUT_M1027_d N_A_364_73#_M1027_g N_A_1152_389#_M1015_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.3328 AS=0.0896 PD=1.68 PS=0.92 NRD=14.988 NRS=0 M=1
+ R=4.26667 SA=75001.3 SB=75004.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_1500_63#_M1008_d N_A_555_73#_M1008_g N_COUT_M1027_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1728 AS=0.3328 PD=1.18 PS=1.68 NRD=48.744 NRS=127.5 M=1 R=4.26667
+ SA=75002.5 SB=75003 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_CIN_M1011_g N_A_1500_63#_M1008_d VNB NSHORT L=0.15
+ W=0.64 AD=0.227805 AS=0.1728 PD=1.37081 PS=1.18 NRD=14.988 NRS=0 M=1 R=4.26667
+ SA=75003.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1022 N_A_1774_367#_M1022_d N_CIN_M1022_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.84 AD=0.184573 AS=0.298995 PD=1.58351 PS=1.79919 NRD=16.428 NRS=54.996 M=1
+ R=5.6 SA=75003.2 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1031 N_A_1926_135#_M1031_d N_A_555_73#_M1031_g N_A_1774_367#_M1022_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.176 AS=0.140627 PD=1.19 PS=1.20649 NRD=50.616 NRS=0
+ M=1 R=4.26667 SA=75002.3 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1028 N_A_1883_395#_M1028_d N_A_364_73#_M1028_g N_A_1926_135#_M1031_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1748 AS=0.176 PD=1.23 PS=1.19 NRD=21.552 NRS=0 M=1
+ R=4.26667 SA=75003 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1017 N_VGND_M1017_d N_A_1774_367#_M1017_g N_A_1883_395#_M1028_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.228065 AS=0.1748 PD=1.34054 PS=1.23 NRD=142.5 NRS=10.932
+ M=1 R=4.26667 SA=75003.5 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_SUM_M1001_d N_A_1926_135#_M1001_g N_VGND_M1017_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.299335 PD=2.25 PS=1.75946 NRD=0 NRS=11.424 M=1 R=5.6
+ SA=75003.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g N_A_29_47#_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.392551 AS=0.3591 PD=2.10743 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1007 N_A_256_87#_M1007_d N_A_29_47#_M1007_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=1 AD=0.285 AS=0.311549 PD=2.57 PS=1.67257 NRD=0 NRS=69.2652 M=1 R=6.66667
+ SA=75001 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1021 N_A_256_87#_M1021_d N_A_439_47#_M1021_g N_A_364_73#_M1021_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1010 N_A_555_73#_M1010_d N_B_M1010_g N_A_256_87#_M1021_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2345 AS=0.1176 PD=1.49 PS=1.12 NRD=27.5406 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1002 N_A_29_47#_M1002_d N_A_439_47#_M1002_g N_A_555_73#_M1010_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2268 AS=0.2345 PD=1.38 PS=1.49 NRD=0 NRS=26.9693 M=1 R=5.6
+ SA=75001.1 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1014 N_A_364_73#_M1014_d N_B_M1014_g N_A_29_47#_M1002_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.2268 PD=2.27 PS=1.38 NRD=2.3443 NRS=60.9715 M=1 R=5.6
+ SA=75001.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_B_M1013_g N_A_439_47#_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.286622 AS=0.3591 PD=1.89558 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1019 N_A_1152_389#_M1019_d N_A_439_47#_M1019_g N_VPWR_M1013_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.205109 AS=0.227478 PD=1.5163 PS=1.50442 NRD=0 NRS=32.4853 M=1
+ R=6.66667 SA=75000.8 SB=75002.8 A=0.15 P=2.3 MULT=1
MM1030 N_COUT_M1030_d N_A_555_73#_M1030_g N_A_1152_389#_M1019_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.4494 AS=0.172291 PD=1.91 PS=1.2737 NRD=57.4452 NRS=26.9693
+ M=1 R=5.6 SA=75001.3 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1029 N_A_1500_63#_M1029_d N_A_364_73#_M1029_g N_COUT_M1030_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.172291 AS=0.4494 PD=1.2737 PS=1.91 NRD=26.9693 NRS=127.814
+ M=1 R=5.6 SA=75002.6 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_CIN_M1003_g N_A_1500_63#_M1029_d VPB PHIGHVT L=0.15 W=1
+ AD=0.320398 AS=0.205109 PD=1.69027 PS=1.5163 NRD=73.2052 NRS=0 M=1 R=6.66667
+ SA=75002.6 SB=75001 A=0.15 P=2.3 MULT=1
MM1023 N_A_1774_367#_M1023_d N_CIN_M1023_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3465 AS=0.403702 PD=3.07 PS=2.12973 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1020 N_A_1926_135#_M1020_d N_A_555_73#_M1020_g N_A_1883_395#_M1020_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1176 AS=0.2352 PD=1.12 PS=2.24 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1024 N_A_1774_367#_M1024_d N_A_364_73#_M1024_g N_A_1926_135#_M1020_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.392 AS=0.1176 PD=2.92 PS=1.12 NRD=96.53 NRS=0 M=1
+ R=5.6 SA=75000.6 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1025 N_VPWR_M1025_d N_A_1774_367#_M1025_g N_A_1883_395#_M1025_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.27615 AS=0.28 PD=1.60177 PS=2.56 NRD=53.5052 NRS=0 M=1
+ R=6.66667 SA=75000.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1018 N_SUM_M1018_d N_A_1926_135#_M1018_g N_VPWR_M1025_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3528 AS=0.34795 PD=3.08 PS=2.01823 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.8 SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=23.7299 P=29.85
*
.include "sky130_fd_sc_lp__fahcin_1.pxi.spice"
*
.ends
*
*
