* File: sky130_fd_sc_lp__a221o_1.pxi.spice
* Created: Wed Sep  2 09:21:10 2020
* 
x_PM_SKY130_FD_SC_LP__A221O_1%A_80_21# N_A_80_21#_M1009_d N_A_80_21#_M1003_d
+ N_A_80_21#_M1000_d N_A_80_21#_M1001_g N_A_80_21#_M1011_g N_A_80_21#_c_67_n
+ N_A_80_21#_c_68_n N_A_80_21#_c_74_n N_A_80_21#_c_131_p N_A_80_21#_c_69_n
+ N_A_80_21#_c_76_n N_A_80_21#_c_104_p N_A_80_21#_c_77_n N_A_80_21#_c_70_n
+ N_A_80_21#_c_71_n N_A_80_21#_c_101_p N_A_80_21#_c_78_n
+ PM_SKY130_FD_SC_LP__A221O_1%A_80_21#
x_PM_SKY130_FD_SC_LP__A221O_1%A2 N_A2_M1007_g N_A2_M1008_g A2 A2 A2 N_A2_c_176_n
+ N_A2_c_177_n PM_SKY130_FD_SC_LP__A221O_1%A2
x_PM_SKY130_FD_SC_LP__A221O_1%A1 N_A1_M1009_g N_A1_M1002_g A1 A1 A1 N_A1_c_214_n
+ N_A1_c_215_n PM_SKY130_FD_SC_LP__A221O_1%A1
x_PM_SKY130_FD_SC_LP__A221O_1%B1 N_B1_M1010_g N_B1_M1005_g B1 N_B1_c_249_n
+ N_B1_c_250_n N_B1_c_252_n PM_SKY130_FD_SC_LP__A221O_1%B1
x_PM_SKY130_FD_SC_LP__A221O_1%B2 N_B2_c_282_n N_B2_M1004_g N_B2_c_283_n
+ N_B2_M1006_g B2 PM_SKY130_FD_SC_LP__A221O_1%B2
x_PM_SKY130_FD_SC_LP__A221O_1%C1 N_C1_M1003_g N_C1_M1000_g C1 C1 N_C1_c_318_n
+ N_C1_c_319_n PM_SKY130_FD_SC_LP__A221O_1%C1
x_PM_SKY130_FD_SC_LP__A221O_1%X N_X_M1001_s N_X_M1011_s X X X X X X X
+ N_X_c_341_n X PM_SKY130_FD_SC_LP__A221O_1%X
x_PM_SKY130_FD_SC_LP__A221O_1%VPWR N_VPWR_M1011_d N_VPWR_M1002_d N_VPWR_c_357_n
+ N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n VPWR N_VPWR_c_361_n
+ N_VPWR_c_362_n N_VPWR_c_356_n N_VPWR_c_364_n PM_SKY130_FD_SC_LP__A221O_1%VPWR
x_PM_SKY130_FD_SC_LP__A221O_1%A_264_367# N_A_264_367#_M1008_d
+ N_A_264_367#_M1005_d N_A_264_367#_c_414_n N_A_264_367#_c_426_n
+ N_A_264_367#_c_411_n N_A_264_367#_c_418_n N_A_264_367#_c_423_n
+ PM_SKY130_FD_SC_LP__A221O_1%A_264_367#
x_PM_SKY130_FD_SC_LP__A221O_1%A_458_367# N_A_458_367#_M1005_s
+ N_A_458_367#_M1006_d N_A_458_367#_c_434_n N_A_458_367#_c_441_n
+ N_A_458_367#_c_435_n N_A_458_367#_c_453_n N_A_458_367#_c_438_n
+ PM_SKY130_FD_SC_LP__A221O_1%A_458_367#
x_PM_SKY130_FD_SC_LP__A221O_1%VGND N_VGND_M1001_d N_VGND_M1004_d N_VGND_c_459_n
+ N_VGND_c_460_n N_VGND_c_461_n N_VGND_c_462_n VGND N_VGND_c_463_n
+ N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n PM_SKY130_FD_SC_LP__A221O_1%VGND
cc_1 VNB N_A_80_21#_M1001_g 0.0292456f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A_80_21#_c_67_n 0.00431751f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.47
cc_3 VNB N_A_80_21#_c_68_n 0.0347239f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.47
cc_4 VNB N_A_80_21#_c_69_n 0.0119004f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.685
cc_5 VNB N_A_80_21#_c_70_n 0.00795955f $X=-0.19 $Y=-0.245 $X2=3.835 $Y2=0.835
cc_6 VNB N_A_80_21#_c_71_n 0.0221734f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=0.42
cc_7 VNB N_A2_M1008_g 0.00815345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A2 0.0022149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A2 0.00575153f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.305
cc_10 VNB N_A2_c_176_n 0.0356216f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_11 VNB N_A2_c_177_n 0.0177067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_M1002_g 0.00866721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A1 0.00184062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A1 0.006935f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.305
cc_15 VNB N_A1_c_214_n 0.0351098f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_16 VNB N_A1_c_215_n 0.0196659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB B1 0.00346295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_249_n 0.0443357f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.305
cc_19 VNB N_B1_c_250_n 0.0192477f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_20 VNB N_B2_c_282_n 0.0173739f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=0.235
cc_21 VNB N_B2_c_283_n 0.0335076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B2_M1006_g 0.00805065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB B2 0.00620096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C1_M1000_g 0.0115272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB C1 0.0362302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C1_c_318_n 0.0357983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C1_c_319_n 0.0237062f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_28 VNB X 0.029776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_341_n 0.0258088f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.77
cc_30 VNB X 0.00666696f $X=-0.19 $Y=-0.245 $X2=2.257 $Y2=1.015
cc_31 VNB N_VPWR_c_356_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_459_n 0.00564356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_460_n 0.00563065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_461_n 0.0594237f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_35 VNB N_VGND_c_462_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_463_n 0.0184065f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.47
cc_37 VNB N_VGND_c_464_n 0.026989f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.98
cc_38 VNB N_VGND_c_465_n 0.239261f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=2.91
cc_39 VNB N_VGND_c_466_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.835 $Y2=0.835
cc_40 VPB N_A_80_21#_M1011_g 0.0237672f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_41 VPB N_A_80_21#_c_68_n 0.0078414f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.47
cc_42 VPB N_A_80_21#_c_74_n 0.0158681f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=1.77
cc_43 VPB N_A_80_21#_c_69_n 6.70288e-19 $X=-0.19 $Y=1.655 $X2=2.115 $Y2=1.685
cc_44 VPB N_A_80_21#_c_76_n 0.0199642f $X=-0.19 $Y=1.655 $X2=3.64 $Y2=1.77
cc_45 VPB N_A_80_21#_c_77_n 0.0474727f $X=-0.19 $Y=1.655 $X2=3.805 $Y2=1.98
cc_46 VPB N_A_80_21#_c_78_n 0.00229695f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=1.77
cc_47 VPB N_A2_M1008_g 0.0213006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A1_M1002_g 0.0227442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B1_c_249_n 0.013102f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.305
cc_50 VPB N_B1_c_252_n 0.0203226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B2_M1006_g 0.0199179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_C1_M1000_g 0.0247075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB X 0.0567012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_357_n 0.00183427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_358_n 0.00974806f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_56 VPB N_VPWR_c_359_n 0.0130519f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.685
cc_57 VPB N_VPWR_c_360_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.47
cc_58 VPB N_VPWR_c_361_n 0.0153759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_362_n 0.0590673f $X=-0.19 $Y=1.655 $X2=3.805 $Y2=2.91
cc_60 VPB N_VPWR_c_356_n 0.0633364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_364_n 0.0104351f $X=-0.19 $Y=1.655 $X2=3.805 $Y2=0.42
cc_62 VPB N_A_264_367#_c_411_n 0.0114475f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_63 VPB N_A_458_367#_c_434_n 0.0051799f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_458_367#_c_435_n 0.00182193f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_65 N_A_80_21#_M1011_g N_A2_M1008_g 0.00615779f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_67_n N_A2_M1008_g 0.00109182f $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_67 N_A_80_21#_c_68_n N_A2_M1008_g 0.00525516f $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_74_n N_A2_M1008_g 0.0156049f $X=2.025 $Y=1.77 $X2=0 $Y2=0
cc_69 N_A_80_21#_M1001_g A2 0.0019208f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_70 N_A_80_21#_M1001_g A2 5.86648e-19 $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_67_n A2 0.0100194f $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_68_n A2 6.61114e-19 $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_74_n A2 0.023994f $X=2.025 $Y=1.77 $X2=0 $Y2=0
cc_74 N_A_80_21#_M1001_g N_A2_c_176_n 0.00318644f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_67_n N_A2_c_176_n 7.83826e-19 $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_68_n N_A2_c_176_n 0.0131303f $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_74_n N_A2_c_176_n 0.00384651f $X=2.025 $Y=1.77 $X2=0 $Y2=0
cc_78 N_A_80_21#_M1001_g N_A2_c_177_n 0.0134806f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_74_n N_A1_M1002_g 0.0122918f $X=2.025 $Y=1.77 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_69_n N_A1_M1002_g 0.00350319f $X=2.115 $Y=1.685 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_69_n A1 0.00785433f $X=2.115 $Y=1.685 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_74_n A1 0.0247751f $X=2.025 $Y=1.77 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_69_n A1 0.0248494f $X=2.115 $Y=1.685 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_74_n N_A1_c_214_n 0.00374077f $X=2.025 $Y=1.77 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_69_n N_A1_c_214_n 0.00283446f $X=2.115 $Y=1.685 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_69_n N_A1_c_215_n 0.00108516f $X=2.115 $Y=1.685 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_101_p N_A1_c_215_n 0.00829042f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_69_n B1 0.0241746f $X=2.115 $Y=1.685 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_76_n B1 0.0291949f $X=3.64 $Y=1.77 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_104_p B1 0.0131373f $X=3.7 $Y=0.925 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_101_p B1 0.0133542f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_69_n N_B1_c_249_n 0.00758205f $X=2.115 $Y=1.685 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_76_n N_B1_c_249_n 0.0134291f $X=3.64 $Y=1.77 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_101_p N_B1_c_249_n 0.00680255f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_69_n N_B1_c_250_n 0.00453093f $X=2.115 $Y=1.685 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_104_p N_B1_c_250_n 0.00898084f $X=3.7 $Y=0.925 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_101_p N_B1_c_250_n 0.0124524f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_76_n N_B1_c_252_n 0.00876406f $X=3.64 $Y=1.77 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_104_p N_B2_c_282_n 0.0131558f $X=3.7 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_80_21#_c_101_p N_B2_c_282_n 0.00208942f $X=2.415 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_80_21#_c_76_n N_B2_c_283_n 0.00227942f $X=3.64 $Y=1.77 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_104_p N_B2_c_283_n 0.00134633f $X=3.7 $Y=0.925 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_76_n N_B2_M1006_g 0.0150591f $X=3.64 $Y=1.77 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_77_n N_B2_M1006_g 9.88871e-19 $X=3.805 $Y=1.98 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_76_n B2 0.0246472f $X=3.64 $Y=1.77 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_104_p B2 0.0225117f $X=3.7 $Y=0.925 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_76_n N_C1_M1000_g 0.0154616f $X=3.64 $Y=1.77 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_77_n N_C1_M1000_g 0.0170021f $X=3.805 $Y=1.98 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_76_n C1 0.0305384f $X=3.64 $Y=1.77 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_104_p C1 0.0139424f $X=3.7 $Y=0.925 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_70_n C1 0.0214512f $X=3.835 $Y=0.835 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_76_n N_C1_c_318_n 0.00442554f $X=3.64 $Y=1.77 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_70_n N_C1_c_318_n 0.00331083f $X=3.835 $Y=0.835 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_104_p N_C1_c_319_n 0.0110744f $X=3.7 $Y=0.925 $X2=0 $Y2=0
cc_115 N_A_80_21#_M1001_g X 0.0255503f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_67_n X 0.0288424f $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_131_p X 0.0131656f $X=0.765 $Y=1.77 $X2=0 $Y2=0
cc_118 N_A_80_21#_M1001_g N_X_c_341_n 0.0106142f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_119 N_A_80_21#_M1001_g X 0.00503192f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_74_n N_VPWR_M1011_d 0.00373705f $X=2.025 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_80_21#_c_131_p N_VPWR_M1011_d 0.00172619f $X=0.765 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_80_21#_c_74_n N_VPWR_M1002_d 0.00230586f $X=2.025 $Y=1.77 $X2=0 $Y2=0
cc_123 N_A_80_21#_M1011_g N_VPWR_c_357_n 0.0194251f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_124 N_A_80_21#_c_68_n N_VPWR_c_357_n 9.86686e-19 $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_74_n N_VPWR_c_357_n 0.0300624f $X=2.025 $Y=1.77 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_131_p N_VPWR_c_357_n 0.0159833f $X=0.765 $Y=1.77 $X2=0 $Y2=0
cc_127 N_A_80_21#_M1011_g N_VPWR_c_361_n 0.00486043f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_A_80_21#_c_77_n N_VPWR_c_362_n 0.0210467f $X=3.805 $Y=1.98 $X2=0 $Y2=0
cc_129 N_A_80_21#_M1000_d N_VPWR_c_356_n 0.00215158f $X=3.665 $Y=1.835 $X2=0
+ $Y2=0
cc_130 N_A_80_21#_M1011_g N_VPWR_c_356_n 0.00917987f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_A_80_21#_c_77_n N_VPWR_c_356_n 0.0125689f $X=3.805 $Y=1.98 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_74_n N_A_264_367#_M1008_d 0.00181776f $X=2.025 $Y=1.77
+ $X2=-0.19 $Y2=-0.245
cc_133 N_A_80_21#_c_76_n N_A_264_367#_M1005_d 0.00261503f $X=3.64 $Y=1.77 $X2=0
+ $Y2=0
cc_134 N_A_80_21#_c_74_n N_A_264_367#_c_414_n 0.0139123f $X=2.025 $Y=1.77 $X2=0
+ $Y2=0
cc_135 N_A_80_21#_c_74_n N_A_264_367#_c_411_n 0.0255797f $X=2.025 $Y=1.77 $X2=0
+ $Y2=0
cc_136 N_A_80_21#_c_76_n N_A_264_367#_c_411_n 0.0316376f $X=3.64 $Y=1.77 $X2=0
+ $Y2=0
cc_137 N_A_80_21#_c_78_n N_A_264_367#_c_411_n 0.0151096f $X=2.115 $Y=1.77 $X2=0
+ $Y2=0
cc_138 N_A_80_21#_c_76_n N_A_264_367#_c_418_n 0.0211892f $X=3.64 $Y=1.77 $X2=0
+ $Y2=0
cc_139 N_A_80_21#_c_76_n N_A_458_367#_M1005_s 0.00221647f $X=3.64 $Y=1.77
+ $X2=-0.19 $Y2=-0.245
cc_140 N_A_80_21#_c_76_n N_A_458_367#_M1006_d 0.00197722f $X=3.64 $Y=1.77 $X2=0
+ $Y2=0
cc_141 N_A_80_21#_c_76_n N_A_458_367#_c_438_n 0.0151327f $X=3.64 $Y=1.77 $X2=0
+ $Y2=0
cc_142 N_A_80_21#_c_104_p N_VGND_M1004_d 0.00927245f $X=3.7 $Y=0.925 $X2=0 $Y2=0
cc_143 N_A_80_21#_M1001_g N_VGND_c_459_n 0.0124534f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_144 N_A_80_21#_c_67_n N_VGND_c_459_n 0.00842919f $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_145 N_A_80_21#_c_68_n N_VGND_c_459_n 0.00109583f $X=0.6 $Y=1.47 $X2=0 $Y2=0
cc_146 N_A_80_21#_c_74_n N_VGND_c_459_n 0.00542444f $X=2.025 $Y=1.77 $X2=0 $Y2=0
cc_147 N_A_80_21#_c_104_p N_VGND_c_460_n 0.0261077f $X=3.7 $Y=0.925 $X2=0 $Y2=0
cc_148 N_A_80_21#_c_101_p N_VGND_c_460_n 0.0133153f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_149 N_A_80_21#_c_101_p N_VGND_c_461_n 0.0431415f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_150 N_A_80_21#_M1001_g N_VGND_c_463_n 0.0054895f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_151 N_A_80_21#_c_71_n N_VGND_c_464_n 0.0181659f $X=3.805 $Y=0.42 $X2=0 $Y2=0
cc_152 N_A_80_21#_M1009_d N_VGND_c_465_n 0.0125587f $X=1.755 $Y=0.235 $X2=0
+ $Y2=0
cc_153 N_A_80_21#_M1003_d N_VGND_c_465_n 0.00236652f $X=3.665 $Y=0.235 $X2=0
+ $Y2=0
cc_154 N_A_80_21#_M1001_g N_VGND_c_465_n 0.0115508f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_155 N_A_80_21#_c_104_p N_VGND_c_465_n 0.0255174f $X=3.7 $Y=0.925 $X2=0 $Y2=0
cc_156 N_A_80_21#_c_71_n N_VGND_c_465_n 0.0104192f $X=3.805 $Y=0.42 $X2=0 $Y2=0
cc_157 N_A_80_21#_c_101_p N_VGND_c_465_n 0.0248154f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_158 N_A_80_21#_c_104_p A_541_47# 0.00364351f $X=3.7 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A2_M1008_g N_A1_M1002_g 0.0307444f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_160 A2 A1 0.0320963f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_161 N_A2_c_177_n A1 0.00179244f $X=1.147 $Y=1.185 $X2=0 $Y2=0
cc_162 A2 A1 0.0320963f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A2_c_176_n A1 0.00179244f $X=1.14 $Y=1.35 $X2=0 $Y2=0
cc_164 A2 N_A1_c_214_n 9.23157e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A2_c_176_n N_A1_c_214_n 0.0307444f $X=1.14 $Y=1.35 $X2=0 $Y2=0
cc_166 A2 N_A1_c_215_n 9.23157e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_167 N_A2_c_177_n N_A1_c_215_n 0.0307444f $X=1.147 $Y=1.185 $X2=0 $Y2=0
cc_168 N_A2_M1008_g N_VPWR_c_357_n 0.0170993f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A2_M1008_g N_VPWR_c_358_n 6.47631e-19 $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A2_M1008_g N_VPWR_c_359_n 0.00486043f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A2_M1008_g N_VPWR_c_356_n 0.00828469f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A2_c_177_n N_VGND_c_459_n 0.00726963f $X=1.147 $Y=1.185 $X2=0 $Y2=0
cc_173 A2 N_VGND_c_461_n 0.00923851f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_174 N_A2_c_177_n N_VGND_c_461_n 0.00372875f $X=1.147 $Y=1.185 $X2=0 $Y2=0
cc_175 A2 N_VGND_c_465_n 0.00855134f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_176 N_A2_c_177_n N_VGND_c_465_n 0.00618949f $X=1.147 $Y=1.185 $X2=0 $Y2=0
cc_177 N_A1_M1002_g N_B1_c_249_n 0.00304509f $X=1.68 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A1_c_214_n N_B1_c_249_n 0.00881334f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_179 N_A1_M1002_g N_VPWR_c_357_n 7.07902e-19 $X=1.68 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A1_M1002_g N_VPWR_c_358_n 0.0141948f $X=1.68 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A1_M1002_g N_VPWR_c_359_n 0.00486043f $X=1.68 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A1_M1002_g N_VPWR_c_356_n 0.00828469f $X=1.68 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A1_M1002_g N_A_264_367#_c_411_n 0.0143f $X=1.68 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A1_M1002_g N_A_458_367#_c_434_n 0.00102588f $X=1.68 $Y=2.465 $X2=0
+ $Y2=0
cc_185 A1 N_VGND_c_461_n 0.00901346f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_186 N_A1_c_215_n N_VGND_c_461_n 0.00372875f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_187 A1 N_VGND_c_465_n 0.00780391f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_188 N_A1_c_215_n N_VGND_c_465_n 0.00689865f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_189 A1 A_264_47# 0.00653283f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_190 N_B1_c_250_n N_B2_c_282_n 0.0382234f $X=2.505 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_191 B1 N_B2_c_283_n 0.00206146f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_192 N_B1_c_249_n N_B2_c_283_n 0.047714f $X=2.47 $Y=1.35 $X2=0 $Y2=0
cc_193 N_B1_c_249_n N_B2_M1006_g 0.0439426f $X=2.47 $Y=1.35 $X2=0 $Y2=0
cc_194 B1 B2 0.026516f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_195 N_B1_c_249_n B2 3.38201e-19 $X=2.47 $Y=1.35 $X2=0 $Y2=0
cc_196 N_B1_c_252_n N_VPWR_c_358_n 0.00359061f $X=2.505 $Y=1.725 $X2=0 $Y2=0
cc_197 N_B1_c_252_n N_VPWR_c_362_n 0.00357842f $X=2.505 $Y=1.725 $X2=0 $Y2=0
cc_198 N_B1_c_252_n N_VPWR_c_356_n 0.00687291f $X=2.505 $Y=1.725 $X2=0 $Y2=0
cc_199 N_B1_c_249_n N_A_264_367#_c_411_n 0.00116726f $X=2.47 $Y=1.35 $X2=0 $Y2=0
cc_200 N_B1_c_252_n N_A_264_367#_c_411_n 0.0167616f $X=2.505 $Y=1.725 $X2=0
+ $Y2=0
cc_201 N_B1_c_252_n N_A_458_367#_c_434_n 0.00912841f $X=2.505 $Y=1.725 $X2=0
+ $Y2=0
cc_202 N_B1_c_252_n N_A_458_367#_c_441_n 0.0109018f $X=2.505 $Y=1.725 $X2=0
+ $Y2=0
cc_203 N_B1_c_252_n N_A_458_367#_c_435_n 5.81207e-19 $X=2.505 $Y=1.725 $X2=0
+ $Y2=0
cc_204 N_B1_c_250_n N_VGND_c_461_n 0.0054895f $X=2.505 $Y=1.185 $X2=0 $Y2=0
cc_205 N_B1_c_250_n N_VGND_c_465_n 0.00738979f $X=2.505 $Y=1.185 $X2=0 $Y2=0
cc_206 N_B2_M1006_g N_C1_M1000_g 0.0270981f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B2_c_283_n C1 9.28985e-19 $X=3.14 $Y=1.515 $X2=0 $Y2=0
cc_208 B2 C1 0.0219546f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_209 N_B2_c_283_n N_C1_c_318_n 0.0180163f $X=3.14 $Y=1.515 $X2=0 $Y2=0
cc_210 B2 N_C1_c_318_n 0.00253543f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_211 N_B2_c_282_n N_C1_c_319_n 0.0257801f $X=2.99 $Y=1.185 $X2=0 $Y2=0
cc_212 N_B2_M1006_g N_VPWR_c_362_n 0.00357877f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_213 N_B2_M1006_g N_VPWR_c_356_n 0.00564628f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_214 N_B2_M1006_g N_A_264_367#_c_418_n 0.00180335f $X=3.14 $Y=2.465 $X2=0
+ $Y2=0
cc_215 N_B2_M1006_g N_A_264_367#_c_423_n 0.00683714f $X=3.14 $Y=2.465 $X2=0
+ $Y2=0
cc_216 N_B2_M1006_g N_A_458_367#_c_434_n 4.47609e-19 $X=3.14 $Y=2.465 $X2=0
+ $Y2=0
cc_217 N_B2_M1006_g N_A_458_367#_c_441_n 0.0121902f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B2_c_282_n N_VGND_c_460_n 0.00961532f $X=2.99 $Y=1.185 $X2=0 $Y2=0
cc_219 N_B2_c_282_n N_VGND_c_461_n 0.00585385f $X=2.99 $Y=1.185 $X2=0 $Y2=0
cc_220 N_B2_c_282_n N_VGND_c_465_n 0.00666997f $X=2.99 $Y=1.185 $X2=0 $Y2=0
cc_221 N_C1_M1000_g N_VPWR_c_362_n 0.0054895f $X=3.59 $Y=2.465 $X2=0 $Y2=0
cc_222 N_C1_M1000_g N_VPWR_c_356_n 0.0110868f $X=3.59 $Y=2.465 $X2=0 $Y2=0
cc_223 N_C1_c_319_n N_VGND_c_460_n 0.00584406f $X=3.68 $Y=1.185 $X2=0 $Y2=0
cc_224 N_C1_c_319_n N_VGND_c_464_n 0.00585385f $X=3.68 $Y=1.185 $X2=0 $Y2=0
cc_225 N_C1_c_319_n N_VGND_c_465_n 0.00783339f $X=3.68 $Y=1.185 $X2=0 $Y2=0
cc_226 X N_VPWR_c_361_n 0.0181731f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_227 N_X_M1011_s N_VPWR_c_356_n 0.0040649f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_228 X N_VPWR_c_356_n 0.0100252f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_229 N_X_c_341_n N_VGND_c_459_n 0.0542326f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_230 N_X_c_341_n N_VGND_c_463_n 0.0217635f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_231 N_X_M1001_s N_VGND_c_465_n 0.00215158f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_232 N_X_c_341_n N_VGND_c_465_n 0.0129577f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_233 N_VPWR_c_356_n N_A_264_367#_M1008_d 0.00540667f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_234 N_VPWR_c_356_n N_A_264_367#_M1005_d 0.00289524f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_359_n N_A_264_367#_c_426_n 0.012804f $X=1.73 $Y=3.33 $X2=0 $Y2=0
cc_236 N_VPWR_c_356_n N_A_264_367#_c_426_n 0.00750339f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_237 N_VPWR_M1002_d N_A_264_367#_c_411_n 0.00507577f $X=1.755 $Y=1.835 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_358_n N_A_264_367#_c_411_n 0.0220026f $X=1.895 $Y=2.48 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_356_n N_A_458_367#_M1005_s 0.00215158f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_240 N_VPWR_c_356_n N_A_458_367#_M1006_d 0.0039271f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_358_n N_A_458_367#_c_434_n 0.0415428f $X=1.895 $Y=2.48 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_362_n N_A_458_367#_c_441_n 0.0377104f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_356_n N_A_458_367#_c_441_n 0.023861f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_358_n N_A_458_367#_c_435_n 0.0139f $X=1.895 $Y=2.48 $X2=0 $Y2=0
cc_245 N_VPWR_c_362_n N_A_458_367#_c_435_n 0.0212472f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_356_n N_A_458_367#_c_435_n 0.0126566f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_362_n N_A_458_367#_c_453_n 0.0142845f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_356_n N_A_458_367#_c_453_n 0.00855309f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_249 N_A_264_367#_c_411_n N_A_458_367#_M1005_s 0.00485898f $X=2.75 $Y=2.11
+ $X2=-0.19 $Y2=1.655
cc_250 N_A_264_367#_c_411_n N_A_458_367#_c_434_n 0.0220808f $X=2.75 $Y=2.11
+ $X2=0 $Y2=0
cc_251 N_A_264_367#_M1005_d N_A_458_367#_c_441_n 0.0049251f $X=2.705 $Y=1.835
+ $X2=0 $Y2=0
cc_252 N_A_264_367#_c_423_n N_A_458_367#_c_441_n 0.0197499f $X=2.915 $Y=2.625
+ $X2=0 $Y2=0
cc_253 N_VGND_c_465_n A_264_47# 0.00830005f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_254 N_VGND_c_465_n A_541_47# 0.00306596f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
