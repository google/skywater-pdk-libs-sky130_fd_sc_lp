* File: sky130_fd_sc_lp__a22o_1.pex.spice
* Created: Fri Aug 28 09:54:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22O_1%A_80_246# 1 2 9 11 13 17 18 19 20 21 22 25 27
+ 29
c67 22 0 3.30696e-20 $X=0.845 $Y=1.735
c68 11 0 5.53362e-20 $X=0.555 $Y=1.23
r69 33 35 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=0.475 $Y=1.395
+ $X2=0.555 $Y2=1.395
r70 27 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=0.87 $X2=2.06
+ $Y2=0.955
r71 27 29 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.06 $Y=0.87
+ $X2=2.06 $Y2=0.42
r72 23 25 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.64 $Y=1.82 $X2=1.64
+ $Y2=1.98
r73 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.475 $Y=1.735
+ $X2=1.64 $Y2=1.82
r74 21 22 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.475 $Y=1.735
+ $X2=0.845 $Y2=1.735
r75 19 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=0.955
+ $X2=2.06 $Y2=0.955
r76 19 20 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=1.895 $Y=0.955
+ $X2=0.845 $Y2=0.955
r77 18 35 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.71 $Y=1.395
+ $X2=0.555 $Y2=1.395
r78 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.395 $X2=0.71 $Y2=1.395
r79 15 22 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.725 $Y=1.65
+ $X2=0.845 $Y2=1.735
r80 15 17 12.2447 $w=2.38e-07 $l=2.55e-07 $layer=LI1_cond $X=0.725 $Y=1.65
+ $X2=0.725 $Y2=1.395
r81 14 20 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.725 $Y=1.04
+ $X2=0.845 $Y2=0.955
r82 14 17 17.0466 $w=2.38e-07 $l=3.55e-07 $layer=LI1_cond $X=0.725 $Y=1.04
+ $X2=0.725 $Y2=1.395
r83 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.23
+ $X2=0.555 $Y2=1.395
r84 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.555 $Y=1.23
+ $X2=0.555 $Y2=0.7
r85 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.56
+ $X2=0.475 $Y2=1.395
r86 7 9 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=0.475 $Y=1.56
+ $X2=0.475 $Y2=2.465
r87 2 25 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=1.98
r88 1 32 182 $w=1.7e-07 $l=7.68521e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.28 $X2=2.06 $Y2=0.955
r89 1 29 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.28 $X2=2.06 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_1%B2 1 3 6 8 13
c33 8 0 5.53362e-20 $X=1.2 $Y=1.295
r34 13 14 4.57595 $w=3.16e-07 $l=3e-08 $layer=POLY_cond $X=1.395 $Y=1.395
+ $X2=1.425 $Y2=1.395
r35 11 13 22.1171 $w=3.16e-07 $l=1.45e-07 $layer=POLY_cond $X=1.25 $Y=1.395
+ $X2=1.395 $Y2=1.395
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.395 $X2=1.25 $Y2=1.395
r37 8 12 2.88111 $w=3.98e-07 $l=1e-07 $layer=LI1_cond $X=1.215 $Y=1.295
+ $X2=1.215 $Y2=1.395
r38 4 14 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.56
+ $X2=1.425 $Y2=1.395
r39 4 6 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.425 $Y=1.56
+ $X2=1.425 $Y2=2.465
r40 1 13 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.23
+ $X2=1.395 $Y2=1.395
r41 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.395 $Y=1.23
+ $X2=1.395 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_1%B1 3 6 8 11 12 13
c36 13 0 1.63009e-20 $X=1.875 $Y=1.23
c37 12 0 1.53057e-19 $X=1.875 $Y=1.395
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.395
+ $X2=1.875 $Y2=1.23
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.875
+ $Y=1.395 $X2=1.875 $Y2=1.395
r40 8 12 8.3232 $w=2.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.68 $Y=1.345
+ $X2=1.875 $Y2=1.345
r41 4 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.56
+ $X2=1.875 $Y2=1.395
r42 4 6 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.875 $Y=1.56
+ $X2=1.875 $Y2=2.465
r43 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.785 $Y=0.7
+ $X2=1.785 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_1%A1 3 6 8 9 10 16 18
c38 18 0 1.65551e-19 $X=2.415 $Y=1.23
c39 10 0 1.63009e-20 $X=2.64 $Y=1.295
r40 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.395
+ $X2=2.415 $Y2=1.56
r41 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.395
+ $X2=2.415 $Y2=1.23
r42 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.395 $X2=2.415 $Y2=1.395
r43 10 17 2.84554 $w=4.03e-07 $l=1e-07 $layer=LI1_cond $X=2.532 $Y=1.295
+ $X2=2.532 $Y2=1.395
r44 9 10 9.15279 $w=4.53e-07 $l=2.85e-07 $layer=LI1_cond $X=2.592 $Y=0.925
+ $X2=2.592 $Y2=1.21
r45 8 9 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.592 $Y=0.555
+ $X2=2.592 $Y2=0.925
r46 6 19 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=2.325 $Y=2.465
+ $X2=2.325 $Y2=1.56
r47 3 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.325 $Y=0.7
+ $X2=2.325 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_1%A2 3 6 8 11 13
c25 8 0 1.24942e-20 $X=3.12 $Y=1.295
r26 11 14 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.972 $Y=1.395
+ $X2=2.972 $Y2=1.56
r27 11 13 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.972 $Y=1.395
+ $X2=2.972 $Y2=1.23
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.395 $X2=2.99 $Y2=1.395
r29 8 12 4.2805 $w=3.48e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.385 $X2=2.99
+ $Y2=1.385
r30 6 14 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=2.865 $Y=2.465
+ $X2=2.865 $Y2=1.56
r31 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.865 $Y=0.7
+ $X2=2.865 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_1%X 1 2 7 8 9 10 11 12 13 24 30
r17 22 30 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=0.265 $Y=0.97
+ $X2=0.265 $Y2=0.925
r18 13 44 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.23 $Y=2.775
+ $X2=0.23 $Y2=2.91
r19 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=2.405
+ $X2=0.23 $Y2=2.775
r20 11 12 16.6464 $w=2.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.23 $Y=2.015
+ $X2=0.23 $Y2=2.405
r21 10 11 14.9391 $w=2.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.23 $Y=1.665
+ $X2=0.23 $Y2=2.015
r22 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.665
r23 9 47 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.14
r24 8 47 5.60547 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.265 $Y=0.99
+ $X2=0.265 $Y2=1.14
r25 8 22 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=0.265 $Y=0.99
+ $X2=0.265 $Y2=0.97
r26 8 30 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=0.265 $Y=0.905
+ $X2=0.265 $Y2=0.925
r27 7 8 11.8634 $w=3.38e-07 $l=3.5e-07 $layer=LI1_cond $X=0.265 $Y=0.555
+ $X2=0.265 $Y2=0.905
r28 7 24 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.265 $Y=0.555
+ $X2=0.265 $Y2=0.425
r29 2 44 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r30 2 11 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.015
r31 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.215
+ $Y=0.28 $X2=0.34 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_1%VPWR 1 2 9 15 19 21 26 36 37 40 43
r45 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 37 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 34 43 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=2.595 $Y2=3.33
r50 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r55 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 27 40 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 26 43 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=2.595 $Y2=3.33
r59 26 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 21 40 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 21 23 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 19 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 19 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 15 18 26.9468 $w=3.38e-07 $l=7.95e-07 $layer=LI1_cond $X=2.595 $Y=2.155
+ $X2=2.595 $Y2=2.95
r67 13 43 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=3.33
r68 13 18 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=2.95
r69 9 12 33.933 $w=2.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.72 $Y=2.155
+ $X2=0.72 $Y2=2.95
r70 7 40 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r71 7 12 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.95
r72 2 18 400 $w=1.7e-07 $l=1.21088e-06 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.835 $X2=2.6 $Y2=2.95
r73 2 15 400 $w=1.7e-07 $l=4.07922e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.835 $X2=2.6 $Y2=2.155
r74 1 12 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.95
r75 1 9 400 $w=1.7e-07 $l=3.83667e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_1%A_217_367# 1 2 3 10 12 14 17 19 20 21 24
r42 24 26 34.5733 $w=3.08e-07 $l=9.3e-07 $layer=LI1_cond $X=3.09 $Y=1.98
+ $X2=3.09 $Y2=2.91
r43 22 24 2.97405 $w=3.08e-07 $l=8e-08 $layer=LI1_cond $X=3.09 $Y=1.9 $X2=3.09
+ $Y2=1.98
r44 20 22 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.935 $Y=1.815
+ $X2=3.09 $Y2=1.9
r45 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.935 $Y=1.815
+ $X2=2.255 $Y2=1.815
r46 17 31 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=2.905
+ $X2=2.115 $Y2=2.99
r47 17 19 38.0718 $w=2.78e-07 $l=9.25e-07 $layer=LI1_cond $X=2.115 $Y=2.905
+ $X2=2.115 $Y2=1.98
r48 16 21 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.115 $Y=1.9
+ $X2=2.255 $Y2=1.815
r49 16 19 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=2.115 $Y=1.9 $X2=2.115
+ $Y2=1.98
r50 15 29 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.305 $Y=2.99
+ $X2=1.175 $Y2=2.99
r51 14 31 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.975 $Y=2.99
+ $X2=2.115 $Y2=2.99
r52 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=2.99
+ $X2=1.305 $Y2=2.99
r53 10 29 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=2.905
+ $X2=1.175 $Y2=2.99
r54 10 12 33.2435 $w=2.58e-07 $l=7.5e-07 $layer=LI1_cond $X=1.175 $Y=2.905
+ $X2=1.175 $Y2=2.155
r55 3 26 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=2.91
r56 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=1.98
r57 2 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.835 $X2=2.09 $Y2=2.91
r58 2 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.835 $X2=2.09 $Y2=1.98
r59 1 29 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.21 $Y2=2.91
r60 1 12 400 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.21 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_1%VGND 1 2 7 9 11 13 18 28 37
r37 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r38 29 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r39 28 33 9.29385 $w=7.38e-07 $l=5.75e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.975 $Y2=0.575
r40 28 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 25 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r43 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 21 24 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r45 19 28 9.68893 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=0.975
+ $Y2=0
r46 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.68
+ $Y2=0
r47 18 36 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r48 18 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r49 16 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r50 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 13 28 9.68893 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.975
+ $Y2=0
r52 13 15 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.24
+ $Y2=0
r53 11 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r54 11 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r55 11 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 7 36 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r57 7 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.08 $Y=0.085 $X2=3.08
+ $Y2=0.425
r58 2 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.28 $X2=3.08 $Y2=0.425
r59 1 33 91 $w=1.7e-07 $l=6.81726e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.28 $X2=1.18 $Y2=0.575
.ends

