* File: sky130_fd_sc_lp__a31o_m.spice
* Created: Wed Sep  2 09:26:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a31o_m.pex.spice"
.subckt sky130_fd_sc_lp__a31o_m  VNB VPB A3 A2 A1 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_86_172#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.1113 PD=0.77 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1003 A_282_66# N_A3_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0735 PD=0.63 PS=0.77 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.7 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1004 A_354_66# N_A2_M1004_g A_282_66# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.1 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_86_172#_M1001_d N_A1_M1001_g A_354_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_B1_M1006_g N_A_86_172#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_86_172#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_274_512#_M1008_d N_A3_M1008_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_274_512#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_A_274_512#_M1009_d N_A1_M1009_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_86_172#_M1007_d N_B1_M1007_g N_A_274_512#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a31o_m.pxi.spice"
*
.ends
*
*
