* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_345_367# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR A2 a_345_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_345_367# B2 a_108_267# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_631_47# A2 a_739_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND B2 a_432_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_739_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_432_47# B1 a_108_267# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_345_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_108_267# B1 a_345_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR a_108_267# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 X a_108_267# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND a_108_267# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_108_267# A1 a_631_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 X a_108_267# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
