* File: sky130_fd_sc_lp__o2111a_lp.spice
* Created: Wed Sep  2 10:12:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o2111a_lp  VNB VPB A1 A2 B1 C1 D1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D1	D1
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A1_M1012_g N_A_29_51#_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1197 PD=0.78 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_29_51#_M1010_d N_A2_M1010_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0756 PD=0.81 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 A_326_51# N_B1_M1005_g N_A_29_51#_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=31.428 M=1 R=2.8 SA=75001.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_404_51# N_C1_M1003_g A_326_51# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_232_419#_M1004_d N_D1_M1004_g A_404_51# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_708_47# N_A_232_419#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_232_419#_M1001_g A_708_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 A_134_419# N_A1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1000 N_A_232_419#_M1000_d N_A2_M1000_g A_134_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.16 AS=0.12 PD=1.32 PS=1.24 NRD=7.8603 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_B1_M1009_g N_A_232_419#_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.3 AS=0.16 PD=1.6 PS=1.32 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1007 N_A_232_419#_M1007_d N_C1_M1007_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.15 AS=0.3 PD=1.3 PS=1.6 NRD=3.9203 NRS=63.04 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_D1_M1008_g N_A_232_419#_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.15 PD=1.28 PS=1.3 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1002 N_X_M1002_d N_A_232_419#_M1002_g N_VPWR_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__o2111a_lp.pxi.spice"
*
.ends
*
*
