* File: sky130_fd_sc_lp__nand3b_m.spice
* Created: Wed Sep  2 10:05:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand3b_m.pex.spice"
.subckt sky130_fd_sc_lp__nand3b_m  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_N_M1001_g N_A_37_47#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.10605 AS=0.1113 PD=0.925 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 A_251_47# N_C_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.10605 PD=0.63 PS=0.925 NRD=14.28 NRS=64.284 M=1 R=2.8 SA=75000.8
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1004 A_323_47# N_B_M1004_g A_251_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_A_37_47#_M1005_g A_323_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1218 AS=0.0441 PD=1.42 PS=0.63 NRD=7.14 NRS=14.28 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_37_47#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_C_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A_37_47#_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__nand3b_m.pxi.spice"
*
.ends
*
*
