* NGSPICE file created from sky130_fd_sc_lp__o31ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=6.678e+11p pd=6.1e+06u as=8.001e+11p ps=3.79e+06u
M1001 Y B1 a_110_47# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=5.292e+11p ps=4.62e+06u
M1002 Y A3 a_182_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=4.914e+11p ps=3.3e+06u
M1003 a_110_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=7.434e+11p ps=5.13e+06u
M1004 a_110_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_110_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_182_367# A2 a_110_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1007 a_110_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

