* File: sky130_fd_sc_lp__dlrtp_1.spice
* Created: Wed Sep  2 09:47:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrtp_1.pex.spice"
.subckt sky130_fd_sc_lp__dlrtp_1  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_D_M1000_g N_A_41_464#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.09135 AS=0.1113 PD=0.855 PS=1.37 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1013 N_A_249_70#_M1013_d N_GATE_M1013_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.09135 PD=1.37 PS=0.855 NRD=0 NRS=21.42 M=1 R=2.8
+ SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_249_70#_M1012_g N_A_371_473#_M1012_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1003 A_587_47# N_A_41_464#_M1003_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_A_659_47#_M1005_d N_A_371_473#_M1005_g A_587_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 A_767_47# N_A_249_70#_M1009_g N_A_659_47#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_809_21#_M1010_g A_767_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1512 AS=0.0441 PD=1.56 PS=0.63 NRD=27.132 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1006 A_1056_73# N_A_659_47#_M1006_g N_A_809_21#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1019_d N_RESET_B_M1019_g A_1056_73# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.0882 PD=1.23 PS=1.05 NRD=15.708 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1011 N_Q_M1011_d N_A_809_21#_M1011_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 N_VPWR_M1015_d N_D_M1015_g N_A_41_464#_M1015_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.152 AS=0.1696 PD=1.115 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1014 N_A_249_70#_M1014_d N_GATE_M1014_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2048 AS=0.152 PD=1.92 PS=1.115 NRD=16.9223 NRS=60.0062 M=1
+ R=4.26667 SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A_249_70#_M1001_g N_A_371_473#_M1001_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2224 AS=0.1696 PD=1.335 PS=1.81 NRD=90.7973 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1002 A_623_473# N_A_41_464#_M1002_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.2224 PD=0.85 PS=1.335 NRD=15.3857 NRS=36.9178 M=1 R=4.26667
+ SA=75001 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1007 N_A_659_47#_M1007_d N_A_249_70#_M1007_g A_623_473# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.130294 AS=0.0672 PD=1.22566 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.4 SB=75002 A=0.096 P=1.58 MULT=1
MM1017 A_800_473# N_A_371_473#_M1017_g N_A_659_47#_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0855057 PD=0.66 PS=0.80434 NRD=30.4759 NRS=44.5417 M=1
+ R=2.8 SA=75001.9 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_809_21#_M1008_g A_800_473# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.13335 AS=0.0504 PD=1 PS=0.66 NRD=109.04 NRS=30.4759 M=1 R=2.8 SA=75002.3
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1004 N_A_809_21#_M1004_d N_A_659_47#_M1004_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.40005 PD=1.54 PS=3 NRD=0 NRS=35.9525 M=1 R=8.4
+ SA=75001.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_RESET_B_M1016_g N_A_809_21#_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.22365 AS=0.1764 PD=1.615 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75001.6 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1018 N_Q_M1018_d N_A_809_21#_M1018_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.22365 PD=3.05 PS=1.615 NRD=0 NRS=5.4569 M=1 R=8.4 SA=75002.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=13.2415 P=17.93
*
.include "sky130_fd_sc_lp__dlrtp_1.pxi.spice"
*
.ends
*
*
