* File: sky130_fd_sc_lp__o41ai_1.pex.spice
* Created: Fri Aug 28 11:20:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41AI_1%B1 3 7 9 10 11 15
c38 15 0 9.09918e-20 $X=0.29 $Y=1.46
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.46 $X2=0.29 $Y2=1.46
r40 11 15 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=1.46
r41 9 14 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.63 $Y=1.46 $X2=0.29
+ $Y2=1.46
r42 9 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.63 $Y=1.46
+ $X2=0.705 $Y2=1.46
r43 5 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.705 $Y=1.625
+ $X2=0.705 $Y2=1.46
r44 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.705 $Y=1.625
+ $X2=0.705 $Y2=2.465
r45 1 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=1.46
r46 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_1%A4 3 7 9 12 13
c38 13 0 2.55912e-20 $X=1.155 $Y=1.51
c39 12 0 6.54007e-20 $X=1.155 $Y=1.51
r40 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.51
+ $X2=1.155 $Y2=1.675
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.51
+ $X2=1.155 $Y2=1.345
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.51 $X2=1.155 $Y2=1.51
r43 9 13 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.215 $Y=1.665
+ $X2=1.215 $Y2=1.51
r44 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.245 $Y=2.465
+ $X2=1.245 $Y2=1.675
r45 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.235 $Y=0.665
+ $X2=1.235 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_1%A3 3 7 9 10 11 12 18 19
r34 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.51
+ $X2=1.695 $Y2=1.675
r35 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.51
+ $X2=1.695 $Y2=1.345
r36 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.695
+ $Y=1.51 $X2=1.695 $Y2=1.51
r37 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=2.405
+ $X2=1.695 $Y2=2.775
r38 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=2.035
+ $X2=1.695 $Y2=2.405
r39 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=2.035
r40 9 19 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.51
r41 7 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.685 $Y=0.665
+ $X2=1.685 $Y2=1.345
r42 3 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.605 $Y=2.465
+ $X2=1.605 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_1%A2 3 7 9 10 11 12 18 19
r41 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.51
+ $X2=2.235 $Y2=1.675
r42 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.51
+ $X2=2.235 $Y2=1.345
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.51 $X2=2.235 $Y2=1.51
r44 11 12 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.215 $Y=2.405
+ $X2=2.215 $Y2=2.775
r45 10 11 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.215 $Y=2.035
+ $X2=2.215 $Y2=2.405
r46 9 10 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.215 $Y=1.665
+ $X2=2.215 $Y2=2.035
r47 9 19 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.215 $Y=1.665
+ $X2=2.215 $Y2=1.51
r48 7 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.145 $Y=2.465
+ $X2=2.145 $Y2=1.675
r49 3 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.145 $Y=0.665
+ $X2=2.145 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_1%A1 3 5 7 8 9 16
r28 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.375 $X2=2.99 $Y2=1.375
r29 14 16 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.705 $Y=1.375
+ $X2=2.99 $Y2=1.375
r30 12 14 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.685 $Y=1.375
+ $X2=2.705 $Y2=1.375
r31 9 17 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.375
r32 8 17 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.375
r33 5 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.21
+ $X2=2.705 $Y2=1.375
r34 5 7 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.705 $Y=1.21
+ $X2=2.705 $Y2=0.665
r35 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.685 $Y=1.54
+ $X2=2.685 $Y2=1.375
r36 1 3 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.685 $Y=1.54
+ $X2=2.685 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_1%VPWR 1 2 9 12 15 20 23 24 25 26 27 28 42
r45 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 39 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 38 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 35 38 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 32 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 28 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 28 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 26 38 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 26 27 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.88 $Y2=3.33
r56 25 41 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 25 27 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=2.88 $Y2=3.33
r58 23 31 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.31 $Y=3.33 $X2=0.24
+ $Y2=3.33
r59 23 24 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.31 $Y=3.33
+ $X2=0.502 $Y2=3.33
r60 22 35 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.695 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 22 24 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.695 $Y=3.33
+ $X2=0.502 $Y2=3.33
r62 20 21 6.35386 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.502 $Y=2.505
+ $X2=0.502 $Y2=2.34
r63 15 18 29.2783 $w=3.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.88 $Y=2.01
+ $X2=2.88 $Y2=2.95
r64 13 27 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=3.33
r65 13 18 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=2.95
r66 12 24 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.502 $Y=3.245
+ $X2=0.502 $Y2=3.33
r67 11 20 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=0.502 $Y=2.532
+ $X2=0.502 $Y2=2.505
r68 11 12 21.3426 $w=3.83e-07 $l=7.13e-07 $layer=LI1_cond $X=0.502 $Y=2.532
+ $X2=0.502 $Y2=3.245
r69 9 21 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=0.435 $Y=2.09
+ $X2=0.435 $Y2=2.34
r70 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=1.835 $X2=2.9 $Y2=2.95
r71 2 15 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=1.835 $X2=2.9 $Y2=2.01
r72 1 20 300 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=2 $X=0.35
+ $Y=1.835 $X2=0.49 $Y2=2.505
r73 1 9 600 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=0.35
+ $Y=1.835 $X2=0.475 $Y2=2.09
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_1%Y 1 2 7 8 13 17 20 21 23 24
r41 23 24 7.80969 $w=5.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.44 $Y=0.555
+ $X2=0.44 $Y2=0.925
r42 23 28 2.84948 $w=5.78e-07 $l=1.35e-07 $layer=LI1_cond $X=0.44 $Y=0.555
+ $X2=0.44 $Y2=0.42
r43 20 22 4.69647 $w=4.33e-07 $l=1.35e-07 $layer=LI1_cond $X=0.947 $Y=2.035
+ $X2=0.947 $Y2=2.17
r44 20 21 6.69042 $w=4.33e-07 $l=8.5e-08 $layer=LI1_cond $X=0.947 $Y=2.035
+ $X2=0.947 $Y2=1.95
r45 15 17 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.71 $Y=1.43
+ $X2=0.815 $Y2=1.43
r46 13 22 11.5244 $w=2.98e-07 $l=3e-07 $layer=LI1_cond $X=1.015 $Y=2.47
+ $X2=1.015 $Y2=2.17
r47 9 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=1.515
+ $X2=0.815 $Y2=1.43
r48 9 21 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.815 $Y=1.515
+ $X2=0.815 $Y2=1.95
r49 8 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.345
+ $X2=0.71 $Y2=1.43
r50 7 24 12.4294 $w=5.78e-07 $l=3.81838e-07 $layer=LI1_cond $X=0.71 $Y=1.195
+ $X2=0.44 $Y2=0.925
r51 7 8 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.71 $Y=1.195 $X2=0.71
+ $Y2=1.345
r52 2 20 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=0.78
+ $Y=1.835 $X2=1 $Y2=2.035
r53 2 13 300 $w=1.7e-07 $l=7.36834e-07 $layer=licon1_PDIFF $count=2 $X=0.78
+ $Y=1.835 $X2=1 $Y2=2.47
r54 1 28 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=0.365
+ $Y=0.245 $X2=0.49 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_1%A_156_49# 1 2 3 12 15 16 17 20 22 26 28 29
r45 24 26 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.92 $Y=0.87
+ $X2=2.92 $Y2=0.39
r46 23 29 5.91114 $w=2.37e-07 $l=1.4e-07 $layer=LI1_cond $X=2.085 $Y=1.022
+ $X2=1.945 $Y2=1.022
r47 22 24 16.2597 $w=1.33e-07 $l=4.05947e-07 $layer=LI1_cond $X=2.583 $Y=1.022
+ $X2=2.92 $Y2=0.87
r48 22 23 18.8169 $w=3.03e-07 $l=4.98e-07 $layer=LI1_cond $X=2.583 $Y=1.022
+ $X2=2.085 $Y2=1.022
r49 18 29 0.757028 $w=2.8e-07 $l=1.52e-07 $layer=LI1_cond $X=1.945 $Y=0.87
+ $X2=1.945 $Y2=1.022
r50 18 20 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=1.945 $Y=0.87
+ $X2=1.945 $Y2=0.42
r51 16 29 5.91114 $w=2.37e-07 $l=1.70646e-07 $layer=LI1_cond $X=1.805 $Y=1.09
+ $X2=1.945 $Y2=1.022
r52 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.805 $Y=1.09
+ $X2=1.135 $Y2=1.09
r53 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=1.005
+ $X2=1.135 $Y2=1.09
r54 15 28 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.05 $Y=1.005
+ $X2=1.05 $Y2=0.855
r55 10 28 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0.69
+ $X2=0.97 $Y2=0.855
r56 10 12 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.97 $Y=0.69
+ $X2=0.97 $Y2=0.4
r57 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.78
+ $Y=0.245 $X2=2.92 $Y2=0.39
r58 2 20 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.76
+ $Y=0.245 $X2=1.9 $Y2=0.42
r59 1 12 91 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=2 $X=0.78
+ $Y=0.245 $X2=0.97 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r40 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r42 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r43 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r45 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r46 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r48 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r49 19 31 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.16
+ $Y2=0
r50 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.42
+ $Y2=0
r51 18 34 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.585 $Y=0 $X2=3.12
+ $Y2=0
r52 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.42
+ $Y2=0
r53 16 28 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.2
+ $Y2=0
r54 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.47
+ $Y2=0
r55 15 31 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.635 $Y=0 $X2=2.16
+ $Y2=0
r56 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.635 $Y=0 $X2=1.47
+ $Y2=0
r57 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=0.085
+ $X2=2.42 $Y2=0
r58 11 13 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.42 $Y=0.085
+ $X2=2.42 $Y2=0.575
r59 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.47 $Y=0.085 $X2=1.47
+ $Y2=0
r60 7 9 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.47 $Y=0.085
+ $X2=1.47 $Y2=0.41
r61 2 13 182 $w=1.7e-07 $l=4.1821e-07 $layer=licon1_NDIFF $count=1 $X=2.22
+ $Y=0.245 $X2=2.42 $Y2=0.575
r62 1 9 91 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=2 $X=1.31
+ $Y=0.245 $X2=1.47 $Y2=0.41
.ends

