# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__ebufn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__ebufn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.305000 3.895000 2.150000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.537000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995000 1.305000 3.325000 2.150000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.596400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.955000 0.945000 1.125000 ;
        RECT 0.125000 1.125000 0.355000 1.795000 ;
        RECT 0.125000 1.795000 0.855000 1.965000 ;
        RECT 0.615000 0.595000 0.945000 0.955000 ;
        RECT 0.685000 1.965000 0.855000 2.735000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.255000 1.445000 0.425000 ;
      RECT 0.115000  0.425000 0.445000 0.785000 ;
      RECT 0.175000  2.135000 0.505000 2.905000 ;
      RECT 0.175000  2.905000 1.365000 3.075000 ;
      RECT 0.740000  1.295000 2.485000 1.625000 ;
      RECT 1.035000  1.815000 2.145000 1.985000 ;
      RECT 1.035000  1.985000 1.365000 2.905000 ;
      RECT 1.115000  0.425000 1.445000 0.955000 ;
      RECT 1.115000  0.955000 2.375000 1.125000 ;
      RECT 1.545000  2.155000 1.715000 3.245000 ;
      RECT 1.625000  0.085000 1.875000 0.785000 ;
      RECT 1.895000  1.985000 2.145000 3.075000 ;
      RECT 2.045000  0.255000 2.375000 0.955000 ;
      RECT 2.315000  1.625000 2.485000 2.615000 ;
      RECT 2.315000  2.615000 3.165000 2.785000 ;
      RECT 2.605000  0.255000 3.200000 0.585000 ;
      RECT 2.655000  0.585000 3.200000 1.135000 ;
      RECT 2.655000  1.135000 2.825000 2.445000 ;
      RECT 2.995000  2.445000 4.235000 2.615000 ;
      RECT 3.335000  2.785000 3.665000 3.245000 ;
      RECT 3.370000  0.085000 3.700000 1.135000 ;
      RECT 3.835000  2.435000 4.235000 2.445000 ;
      RECT 3.835000  2.615000 4.235000 3.075000 ;
      RECT 3.870000  0.675000 4.235000 1.135000 ;
      RECT 4.065000  1.135000 4.235000 2.435000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__ebufn_2
END LIBRARY
