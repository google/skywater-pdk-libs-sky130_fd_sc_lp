* NGSPICE file created from sky130_fd_sc_lp__mux2i_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
M1000 VPWR S a_126_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.16955e+12p pd=1.619e+07u as=1.4364e+12p ps=1.236e+07u
M1001 Y A0 a_126_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.7262e+12p pd=1.534e+07u as=0p ps=0u
M1002 Y A1 a_470_69# VNB nshort w=840000u l=150000u
+  ad=1.2348e+12p pd=1.134e+07u as=1.2734e+12p ps=1.004e+07u
M1003 a_1418_21# S VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=1.1634e+12p ps=1.117e+07u
M1004 VPWR S a_126_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_110_69# A0 Y VNB nshort w=840000u l=150000u
+  ad=9.408e+11p pd=8.96e+06u as=0p ps=0u
M1006 VGND a_1418_21# a_110_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A1 a_470_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.4112e+12p ps=1.232e+07u
M1008 VPWR a_1418_21# a_470_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_110_69# a_1418_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND S a_470_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_1418_21# a_470_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND S a_470_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A1 a_470_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_126_367# A0 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1418_21# S VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1016 a_126_367# A0 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_126_367# S VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_470_69# A1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A1 a_470_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A0 a_110_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_470_367# a_1418_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_470_367# a_1418_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_470_367# A1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_110_69# A0 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A0 a_126_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_126_367# S VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_1418_21# a_110_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_110_69# a_1418_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A0 a_110_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_470_69# A1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_470_69# S VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_470_367# A1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_470_69# S VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

