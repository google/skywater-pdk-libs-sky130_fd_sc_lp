* File: sky130_fd_sc_lp__buflp_2.pex.spice
* Created: Wed Sep  2 09:36:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFLP_2%A_98_21# 1 2 9 13 15 19 23 25 29 33 35 39 43
+ 45 46 47 49 50 51 54 58 64 66
c116 43 0 1.82654e-19 $X=1.995 $Y=0.655
r117 62 70 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.967 $Y=1.43
+ $X2=1.967 $Y2=1.595
r118 61 64 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.99 $Y=1.43
+ $X2=2.2 $Y2=1.43
r119 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=1.43 $X2=1.99 $Y2=1.43
r120 56 66 3.22182 $w=2.92e-07 $l=1.01833e-07 $layer=LI1_cond $X=3.117 $Y=0.885
+ $X2=3.08 $Y2=0.8
r121 56 58 51.747 $w=2.53e-07 $l=1.145e-06 $layer=LI1_cond $X=3.117 $Y=0.885
+ $X2=3.117 $Y2=2.03
r122 52 66 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.715
+ $X2=3.08 $Y2=0.8
r123 52 54 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.08 $Y=0.715
+ $X2=3.08 $Y2=0.465
r124 50 66 3.35233 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0.8
+ $X2=3.08 $Y2=0.8
r125 50 51 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.915 $Y=0.8
+ $X2=2.285 $Y2=0.8
r126 49 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.2 $Y=1.265
+ $X2=2.2 $Y2=1.43
r127 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.2 $Y=0.885
+ $X2=2.285 $Y2=0.8
r128 48 49 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.2 $Y=0.885
+ $X2=2.2 $Y2=1.265
r129 43 68 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.995 $Y=0.655
+ $X2=1.995 $Y2=1.265
r130 39 70 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.855 $Y=2.465
+ $X2=1.855 $Y2=1.595
r131 36 47 12.05 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.57 $Y=1.34 $X2=1.46
+ $Y2=1.34
r132 35 62 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=1.967 $Y=1.34
+ $X2=1.967 $Y2=1.43
r133 35 68 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=1.967 $Y=1.34
+ $X2=1.967 $Y2=1.265
r134 35 36 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.78 $Y=1.34
+ $X2=1.57 $Y2=1.34
r135 31 47 12.05 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.495 $Y=1.265
+ $X2=1.46 $Y2=1.34
r136 31 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=1.265
+ $X2=1.495 $Y2=0.655
r137 27 47 12.05 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.425 $Y=1.415
+ $X2=1.46 $Y2=1.34
r138 27 29 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.425 $Y=1.415
+ $X2=1.425 $Y2=2.465
r139 26 46 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.07 $Y=1.34 $X2=0.995
+ $Y2=1.34
r140 25 47 12.05 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.35 $Y=1.34 $X2=1.46
+ $Y2=1.34
r141 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.35 $Y=1.34
+ $X2=1.07 $Y2=1.34
r142 21 46 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.995 $Y=1.415
+ $X2=0.995 $Y2=1.34
r143 21 23 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.995 $Y=1.415
+ $X2=0.995 $Y2=2.465
r144 17 46 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.995 $Y=1.265
+ $X2=0.995 $Y2=1.34
r145 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.265
+ $X2=0.995 $Y2=0.655
r146 16 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.64 $Y=1.34
+ $X2=0.565 $Y2=1.34
r147 15 46 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.92 $Y=1.34 $X2=0.995
+ $Y2=1.34
r148 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.92 $Y=1.34
+ $X2=0.64 $Y2=1.34
r149 11 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.565 $Y=1.415
+ $X2=0.565 $Y2=1.34
r150 11 13 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.565 $Y=1.415
+ $X2=0.565 $Y2=2.465
r151 7 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.565 $Y=1.265
+ $X2=0.565 $Y2=1.34
r152 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.565 $Y=1.265
+ $X2=0.565 $Y2=0.655
r153 2 58 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.885 $X2=3.075 $Y2=2.03
r154 1 54 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_2%A 3 7 11 14 18 19 20 21 22 23 24 36
r46 34 36 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=2.64 $Y=1.22
+ $X2=2.865 $Y2=1.22
r47 32 34 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.505 $Y=1.22
+ $X2=2.64 $Y2=1.22
r48 30 32 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.47 $Y=1.22
+ $X2=2.505 $Y2=1.22
r49 23 24 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=2.405
+ $X2=2.64 $Y2=2.775
r50 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=2.035
+ $X2=2.64 $Y2=2.405
r51 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=2.035
r52 20 21 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.64 $Y=1.22
+ $X2=2.64 $Y2=1.665
r53 20 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.64
+ $Y=1.22 $X2=2.64 $Y2=1.22
r54 18 19 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=2.862 $Y=1.625
+ $X2=2.862 $Y2=1.775
r55 16 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.385
+ $X2=2.865 $Y2=1.22
r56 16 18 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.865 $Y=1.385
+ $X2=2.865 $Y2=1.625
r57 12 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.055
+ $X2=2.865 $Y2=1.22
r58 12 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.865 $Y=1.055
+ $X2=2.865 $Y2=0.445
r59 11 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.86 $Y=2.205
+ $X2=2.86 $Y2=1.775
r60 5 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=1.055
+ $X2=2.505 $Y2=1.22
r61 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.505 $Y=1.055
+ $X2=2.505 $Y2=0.445
r62 1 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=1.385
+ $X2=2.47 $Y2=1.22
r63 1 3 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.47 $Y=1.385 $X2=2.47
+ $Y2=2.205
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_2%VPWR 1 2 7 9 15 19 21 31 32 38
r40 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 32 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.14 $Y2=3.33
r45 29 31 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 25 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r48 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 22 35 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r50 22 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 21 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=2.14 $Y2=3.33
r52 21 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 19 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 19 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 19 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 15 18 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=2.14 $Y=1.98
+ $X2=2.14 $Y2=2.465
r57 13 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=3.245
+ $X2=2.14 $Y2=3.33
r58 13 18 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.14 $Y=3.245
+ $X2=2.14 $Y2=2.465
r59 9 12 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=0.28 $Y=1.98 $X2=0.28
+ $Y2=2.95
r60 7 35 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r61 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.95
r62 2 18 300 $w=1.7e-07 $l=7.27461e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.835 $X2=2.14 $Y2=2.465
r63 2 15 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.835 $X2=2.14 $Y2=1.98
r64 1 12 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=2.95
r65 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_2%A_128_367# 1 2 7 9 11 13 15
r26 13 20 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.905
+ $X2=1.68 $Y2=2.99
r27 13 15 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=1.68 $Y=2.905
+ $X2=1.68 $Y2=1.98
r28 12 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.865 $Y=2.99
+ $X2=0.74 $Y2=2.99
r29 11 20 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=2.99
+ $X2=1.68 $Y2=2.99
r30 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.555 $Y=2.99
+ $X2=0.865 $Y2=2.99
r31 7 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=2.905 $X2=0.74
+ $Y2=2.99
r32 7 9 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=0.74 $Y=2.905
+ $X2=0.74 $Y2=1.98
r33 2 20 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=2.91
r34 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=1.98
r35 1 18 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.835 $X2=0.78 $Y2=2.91
r36 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.835 $X2=0.78 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_2%X 1 2 9 13 14 15 16 30 32
c27 9 0 1.82654e-19 $X=1.28 $Y=0.845
r28 21 32 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.21 $Y=1.715 $X2=1.21
+ $Y2=1.665
r29 15 16 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.21 $Y=1.98
+ $X2=1.21 $Y2=2.405
r30 14 32 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=1.21 $Y=1.647
+ $X2=1.21 $Y2=1.665
r31 14 30 3.93806 $w=3.28e-07 $l=9.7e-08 $layer=LI1_cond $X=1.21 $Y=1.647
+ $X2=1.21 $Y2=1.55
r32 14 15 8.66078 $w=3.28e-07 $l=2.48e-07 $layer=LI1_cond $X=1.21 $Y=1.732
+ $X2=1.21 $Y2=1.98
r33 14 21 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=1.21 $Y=1.732
+ $X2=1.21 $Y2=1.715
r34 13 30 20.1678 $w=2.58e-07 $l=4.55e-07 $layer=LI1_cond $X=1.245 $Y=1.095
+ $X2=1.245 $Y2=1.55
r35 7 13 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=0.93
+ $X2=1.28 $Y2=1.095
r36 7 9 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.93 $X2=1.28
+ $Y2=0.845
r37 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.835 $X2=1.21 $Y2=1.98
r38 1 9 182 $w=1.7e-07 $l=7.07248e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.28 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_2%VGND 1 2 7 9 13 15 17 24 25 31
r46 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r47 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 25 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r49 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.28
+ $Y2=0
r51 22 24 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=3.12
+ $Y2=0
r52 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r53 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r54 18 28 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r55 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r56 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.28
+ $Y2=0
r57 17 20 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=0.72 $Y2=0
r58 15 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r59 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r60 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r61 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.38
r62 7 28 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r63 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.38
r64 2 13 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.235 $X2=2.28 $Y2=0.38
r65 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_2%A_128_47# 1 2 9 14 16
r27 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0.34
+ $X2=0.78 $Y2=0.34
r28 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0.34
+ $X2=1.78 $Y2=0.34
r29 9 10 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0.34
+ $X2=0.945 $Y2=0.34
r30 2 16 91 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.235 $X2=1.78 $Y2=0.42
r31 1 14 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.235 $X2=0.78 $Y2=0.42
.ends

