* File: sky130_fd_sc_lp__o211a_lp.pex.spice
* Created: Fri Aug 28 11:02:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211A_LP%A1 3 7 9 10 11 12 16 17
r35 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.405 $Y=1.56
+ $X2=0.405 $Y2=1.725
r36 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.405 $Y=1.56
+ $X2=0.405 $Y2=1.395
r37 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.56 $X2=0.405 $Y2=1.56
r38 11 12 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.342 $Y=1.665
+ $X2=0.342 $Y2=2.035
r39 11 17 2.76018 $w=4.53e-07 $l=1.05e-07 $layer=LI1_cond $X=0.342 $Y=1.665
+ $X2=0.342 $Y2=1.56
r40 10 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.495 $Y=1.965
+ $X2=0.495 $Y2=1.725
r41 7 10 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.545 $Y=2.09
+ $X2=0.545 $Y2=1.965
r42 7 9 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.545 $Y=2.09
+ $X2=0.545 $Y2=2.595
r43 3 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.495 $Y=0.93
+ $X2=0.495 $Y2=1.395
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_LP%A2 3 7 9 10 14 15
r37 14 17 30.6595 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.56
+ $X2=0.97 $Y2=1.725
r38 14 16 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.56
+ $X2=0.97 $Y2=1.395
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.945
+ $Y=1.56 $X2=0.945 $Y2=1.56
r40 9 10 6.91483 $w=6.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.1 $Y=1.665 $X2=1.1
+ $Y2=2.035
r41 9 15 1.96232 $w=6.38e-07 $l=1.05e-07 $layer=LI1_cond $X=1.1 $Y=1.665 $X2=1.1
+ $Y2=1.56
r42 7 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.085 $Y=0.93
+ $X2=1.085 $Y2=1.395
r43 3 17 216.155 $w=2.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.035 $Y=2.595
+ $X2=1.035 $Y2=1.725
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_LP%B1 3 7 9 10 17
c35 7 0 2.9391e-19 $X=1.565 $Y=2.595
r36 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.705
+ $Y=1.77 $X2=1.705 $Y2=1.77
r37 15 17 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.565 $Y=1.77
+ $X2=1.705 $Y2=1.77
r38 13 15 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.515 $Y=1.77
+ $X2=1.565 $Y2=1.77
r39 10 18 10.9071 $w=2.78e-07 $l=2.65e-07 $layer=LI1_cond $X=1.73 $Y=2.035
+ $X2=1.73 $Y2=1.77
r40 9 18 4.32166 $w=2.78e-07 $l=1.05e-07 $layer=LI1_cond $X=1.73 $Y=1.665
+ $X2=1.73 $Y2=1.77
r41 5 15 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.565 $Y=1.935
+ $X2=1.565 $Y2=1.77
r42 5 7 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.565 $Y=1.935
+ $X2=1.565 $Y2=2.595
r43 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.605
+ $X2=1.515 $Y2=1.77
r44 1 3 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.515 $Y=1.605
+ $X2=1.515 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_LP%C1 1 3 6 8 11 12 16
c43 1 0 1.69062e-19 $X=1.905 $Y=1.215
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.51 $X2=2.69 $Y2=1.51
r45 12 17 11.392 $w=4.33e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=1.562
+ $X2=2.69 $Y2=1.562
r46 11 17 1.32465 $w=4.33e-07 $l=5e-08 $layer=LI1_cond $X=2.64 $Y=1.562 $X2=2.69
+ $Y2=1.562
r47 8 16 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.33 $Y=1.51 $X2=2.69
+ $Y2=1.51
r48 8 10 18.6134 $w=3.3e-07 $l=1.5411e-07 $layer=POLY_cond $X=2.33 $Y=1.51
+ $X2=2.205 $Y2=1.445
r49 4 10 7.52206 $w=2.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.205 $Y=1.675
+ $X2=2.205 $Y2=1.445
r50 4 6 228.577 $w=2.5e-07 $l=9.2e-07 $layer=POLY_cond $X=2.205 $Y=1.675
+ $X2=2.205 $Y2=2.595
r51 1 10 47.4098 $w=3.05e-07 $l=3.98748e-07 $layer=POLY_cond $X=1.905 $Y=1.215
+ $X2=2.205 $Y2=1.445
r52 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.905 $Y=1.215
+ $X2=1.905 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_LP%A_232_419# 1 2 3 12 14 16 19 23 26 32 34 38
+ 43 44 45 49
c77 45 0 1.12223e-19 $X=2.405 $Y=2.395
c78 44 0 1.81687e-19 $X=2.405 $Y=2.075
r79 43 45 4.03026 $w=4.58e-07 $l=1.55e-07 $layer=LI1_cond $X=2.405 $Y=2.24
+ $X2=2.405 $Y2=2.395
r80 43 44 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=2.24
+ $X2=2.405 $Y2=2.075
r81 40 41 3.8382 $w=4.45e-07 $l=1.4e-07 $layer=LI1_cond $X=2.12 $Y=0.93 $X2=2.26
+ $Y2=0.93
r82 35 49 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=3.045 $Y=0.96
+ $X2=3.345 $Y2=0.96
r83 35 46 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.045 $Y=0.96
+ $X2=2.955 $Y2=0.96
r84 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.045
+ $Y=0.96 $X2=3.045 $Y2=0.96
r85 32 41 3.17052 $w=4.45e-07 $l=9.88686e-08 $layer=LI1_cond $X=2.345 $Y=0.96
+ $X2=2.26 $Y2=0.93
r86 32 34 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.345 $Y=0.96
+ $X2=3.045 $Y2=0.96
r87 28 41 6.43131 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.26 $Y=1.16 $X2=2.26
+ $Y2=0.93
r88 28 44 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.26 $Y=1.16
+ $X2=2.26 $Y2=2.075
r89 27 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.395
+ $X2=1.3 $Y2=2.395
r90 26 45 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.175 $Y=2.395
+ $X2=2.405 $Y2=2.395
r91 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.175 $Y=2.395
+ $X2=1.465 $Y2=2.395
r92 21 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.125
+ $X2=3.345 $Y2=0.96
r93 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.345 $Y=1.125
+ $X2=3.345 $Y2=1.915
r94 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=0.795
+ $X2=3.345 $Y2=0.96
r95 17 19 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.345 $Y=0.795
+ $X2=3.345 $Y2=0.445
r96 14 23 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=3.295 $Y=2.04
+ $X2=3.295 $Y2=1.915
r97 14 16 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.295 $Y=2.04
+ $X2=3.295 $Y2=2.545
r98 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=0.795
+ $X2=2.955 $Y2=0.96
r99 10 12 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.955 $Y=0.795
+ $X2=2.955 $Y2=0.445
r100 3 43 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.33
+ $Y=2.095 $X2=2.47 $Y2=2.24
r101 2 38 300 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.16
+ $Y=2.095 $X2=1.3 $Y2=2.475
r102 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.72 $X2=2.12 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_LP%VPWR 1 2 3 10 12 16 20 25 26 27 29 39 40 46
r50 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.83 $Y2=3.33
r56 34 36 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 33 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 30 43 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r61 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=1.83 $Y2=3.33
r63 29 32 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 27 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 27 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 25 36 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=3.03 $Y2=3.33
r68 24 39 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.03 $Y2=3.33
r70 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.03 $Y=2.19 $X2=3.03
+ $Y2=2.9
r71 18 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=3.33
r72 18 23 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=2.9
r73 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=3.245
+ $X2=1.83 $Y2=3.33
r74 14 16 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.83 $Y=3.245
+ $X2=1.83 $Y2=2.885
r75 10 43 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r76 10 12 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.475
r77 3 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.885
+ $Y=2.045 $X2=3.03 $Y2=2.9
r78 3 20 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.885
+ $Y=2.045 $X2=3.03 $Y2=2.19
r79 2 16 600 $w=1.7e-07 $l=8.57146e-07 $layer=licon1_PDIFF $count=1 $X=1.69
+ $Y=2.095 $X2=1.83 $Y2=2.885
r80 1 12 300 $w=1.7e-07 $l=4.46654e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_LP%X 1 2 7 8 9 10 11 12 13
r15 13 37 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.6 $Y=2.775
+ $X2=3.6 $Y2=2.9
r16 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=2.405 $X2=3.6
+ $Y2=2.775
r17 12 31 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=3.6 $Y=2.405
+ $X2=3.6 $Y2=2.19
r18 11 31 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=3.6 $Y=2.035
+ $X2=3.6 $Y2=2.19
r19 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=1.665 $X2=3.6
+ $Y2=2.035
r20 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=1.295 $X2=3.6
+ $Y2=1.665
r21 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=0.925 $X2=3.6
+ $Y2=1.295
r22 8 43 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=3.6 $Y=0.925 $X2=3.6
+ $Y2=0.675
r23 7 43 7.86378 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.56 $Y=0.47
+ $X2=3.56 $Y2=0.675
r24 2 37 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=2.045 $X2=3.56 $Y2=2.9
r25 2 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=2.045 $X2=3.56 $Y2=2.19
r26 1 7 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.235 $X2=3.56 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_LP%A_27_144# 1 2 7 11 14
c26 7 0 1.69062e-19 $X=1.135 $Y=1.185
r27 14 16 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.24 $Y=1.015
+ $X2=0.24 $Y2=1.185
r28 9 11 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.3 $Y=1.1 $X2=1.3
+ $Y2=0.93
r29 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.185
+ $X2=0.24 $Y2=1.185
r30 7 9 16.8978 $w=1.14e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.135 $Y=1.185
+ $X2=1.3 $Y2=1.1
r31 7 8 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=1.185
+ $X2=0.365 $Y2=1.185
r32 2 11 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.72 $X2=1.3 $Y2=0.93
r33 1 14 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.72 $X2=0.28 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r41 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.74
+ $Y2=0
r46 27 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.6
+ $Y2=0
r47 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r50 23 25 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r51 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.74
+ $Y2=0
r52 22 25 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.575 $Y=0 $X2=1.2
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r56 17 19 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r57 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r58 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r59 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0
r60 11 13 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0.415
r61 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085 $X2=0.79
+ $Y2=0
r62 7 9 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.79 $Y=0.085 $X2=0.79
+ $Y2=0.845
r63 2 13 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.235 $X2=2.74 $Y2=0.415
r64 1 9 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.57 $Y=0.72
+ $X2=0.79 $Y2=0.845
.ends

