* File: sky130_fd_sc_lp__o311ai_4.pxi.spice
* Created: Wed Sep  2 10:23:59 2020
* 
x_PM_SKY130_FD_SC_LP__O311AI_4%A1 N_A1_c_146_n N_A1_M1002_g N_A1_M1005_g
+ N_A1_c_148_n N_A1_M1016_g N_A1_M1013_g N_A1_c_150_n N_A1_M1018_g N_A1_M1027_g
+ N_A1_c_152_n N_A1_M1028_g N_A1_M1030_g A1 A1 A1 A1 N_A1_c_155_n
+ PM_SKY130_FD_SC_LP__O311AI_4%A1
x_PM_SKY130_FD_SC_LP__O311AI_4%A2 N_A2_c_224_n N_A2_M1000_g N_A2_M1001_g
+ N_A2_c_226_n N_A2_M1015_g N_A2_M1019_g N_A2_c_228_n N_A2_M1023_g N_A2_M1024_g
+ N_A2_c_230_n N_A2_M1039_g N_A2_M1035_g A2 A2 A2 A2 N_A2_c_233_n
+ PM_SKY130_FD_SC_LP__O311AI_4%A2
x_PM_SKY130_FD_SC_LP__O311AI_4%A3 N_A3_M1007_g N_A3_c_319_n N_A3_M1009_g
+ N_A3_M1014_g N_A3_M1026_g N_A3_M1020_g N_A3_M1037_g N_A3_M1031_g N_A3_M1036_g
+ A3 A3 A3 A3 N_A3_c_324_n N_A3_c_325_n PM_SKY130_FD_SC_LP__O311AI_4%A3
x_PM_SKY130_FD_SC_LP__O311AI_4%B1 N_B1_c_416_n N_B1_M1003_g N_B1_M1010_g
+ N_B1_c_417_n N_B1_M1025_g N_B1_M1011_g N_B1_c_418_n N_B1_M1032_g N_B1_M1029_g
+ N_B1_c_419_n N_B1_M1038_g N_B1_M1034_g B1 B1 B1 N_B1_c_414_n N_B1_c_415_n
+ PM_SKY130_FD_SC_LP__O311AI_4%B1
x_PM_SKY130_FD_SC_LP__O311AI_4%C1 N_C1_c_488_n N_C1_M1004_g N_C1_M1008_g
+ N_C1_c_489_n N_C1_M1006_g N_C1_M1012_g N_C1_c_490_n N_C1_M1021_g N_C1_M1017_g
+ N_C1_c_491_n N_C1_M1033_g N_C1_M1022_g C1 C1 C1 C1 C1 N_C1_c_487_n
+ PM_SKY130_FD_SC_LP__O311AI_4%C1
x_PM_SKY130_FD_SC_LP__O311AI_4%A_30_367# N_A_30_367#_M1005_d N_A_30_367#_M1013_d
+ N_A_30_367#_M1030_d N_A_30_367#_M1019_s N_A_30_367#_M1035_s
+ N_A_30_367#_c_569_n N_A_30_367#_c_561_n N_A_30_367#_c_562_n
+ N_A_30_367#_c_572_n N_A_30_367#_c_563_n N_A_30_367#_c_574_n
+ N_A_30_367#_c_564_n N_A_30_367#_c_576_n N_A_30_367#_c_565_n
+ N_A_30_367#_c_578_n N_A_30_367#_c_566_n N_A_30_367#_c_567_n
+ N_A_30_367#_c_568_n PM_SKY130_FD_SC_LP__O311AI_4%A_30_367#
x_PM_SKY130_FD_SC_LP__O311AI_4%VPWR N_VPWR_M1005_s N_VPWR_M1027_s N_VPWR_M1003_d
+ N_VPWR_M1032_d N_VPWR_M1004_s N_VPWR_M1021_s N_VPWR_c_638_n N_VPWR_c_639_n
+ N_VPWR_c_640_n N_VPWR_c_641_n N_VPWR_c_642_n N_VPWR_c_643_n N_VPWR_c_644_n
+ N_VPWR_c_645_n N_VPWR_c_646_n N_VPWR_c_647_n N_VPWR_c_648_n N_VPWR_c_649_n
+ N_VPWR_c_650_n VPWR N_VPWR_c_651_n N_VPWR_c_652_n N_VPWR_c_653_n
+ N_VPWR_c_637_n N_VPWR_c_655_n N_VPWR_c_656_n N_VPWR_c_657_n
+ PM_SKY130_FD_SC_LP__O311AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O311AI_4%A_457_367# N_A_457_367#_M1001_d
+ N_A_457_367#_M1024_d N_A_457_367#_M1014_s N_A_457_367#_M1031_s
+ N_A_457_367#_c_775_n N_A_457_367#_c_777_n N_A_457_367#_c_780_n
+ N_A_457_367#_c_782_n N_A_457_367#_c_774_n N_A_457_367#_c_789_n
+ N_A_457_367#_c_792_n N_A_457_367#_c_795_n N_A_457_367#_c_786_n
+ N_A_457_367#_c_798_n PM_SKY130_FD_SC_LP__O311AI_4%A_457_367#
x_PM_SKY130_FD_SC_LP__O311AI_4%Y N_Y_M1008_s N_Y_M1017_s N_Y_M1014_d N_Y_M1020_d
+ N_Y_M1036_d N_Y_M1025_s N_Y_M1038_s N_Y_M1006_d N_Y_M1033_d N_Y_c_830_n
+ N_Y_c_836_n N_Y_c_831_n N_Y_c_832_n N_Y_c_921_n N_Y_c_876_n N_Y_c_925_n
+ N_Y_c_890_n N_Y_c_961_p N_Y_c_833_n N_Y_c_929_n N_Y_c_899_n N_Y_c_903_n
+ N_Y_c_837_n N_Y_c_838_n N_Y_c_839_n N_Y_c_880_n N_Y_c_884_n N_Y_c_886_n
+ N_Y_c_834_n N_Y_c_908_n Y Y Y N_Y_c_862_n N_Y_c_866_n N_Y_c_946_n N_Y_c_937_n
+ PM_SKY130_FD_SC_LP__O311AI_4%Y
x_PM_SKY130_FD_SC_LP__O311AI_4%VGND N_VGND_M1002_s N_VGND_M1016_s N_VGND_M1028_s
+ N_VGND_M1015_s N_VGND_M1039_s N_VGND_M1009_s N_VGND_M1037_s N_VGND_c_969_n
+ N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n N_VGND_c_974_n
+ N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n N_VGND_c_978_n N_VGND_c_979_n
+ N_VGND_c_980_n N_VGND_c_981_n VGND N_VGND_c_982_n N_VGND_c_983_n
+ N_VGND_c_984_n N_VGND_c_985_n N_VGND_c_986_n N_VGND_c_987_n N_VGND_c_988_n
+ N_VGND_c_989_n N_VGND_c_990_n PM_SKY130_FD_SC_LP__O311AI_4%VGND
x_PM_SKY130_FD_SC_LP__O311AI_4%A_113_47# N_A_113_47#_M1002_d N_A_113_47#_M1018_d
+ N_A_113_47#_M1000_d N_A_113_47#_M1023_d N_A_113_47#_M1007_d
+ N_A_113_47#_M1026_d N_A_113_47#_M1010_s N_A_113_47#_M1029_s
+ N_A_113_47#_c_1161_n N_A_113_47#_c_1115_n N_A_113_47#_c_1119_n
+ N_A_113_47#_c_1166_n N_A_113_47#_c_1121_n N_A_113_47#_c_1171_n
+ N_A_113_47#_c_1127_n N_A_113_47#_c_1176_n N_A_113_47#_c_1131_n
+ N_A_113_47#_c_1182_n N_A_113_47#_c_1138_n N_A_113_47#_c_1133_n
+ N_A_113_47#_c_1193_n N_A_113_47#_c_1114_n N_A_113_47#_c_1123_n
+ N_A_113_47#_c_1134_n N_A_113_47#_c_1136_n N_A_113_47#_c_1154_n
+ PM_SKY130_FD_SC_LP__O311AI_4%A_113_47#
x_PM_SKY130_FD_SC_LP__O311AI_4%A_1166_65# N_A_1166_65#_M1010_d
+ N_A_1166_65#_M1011_d N_A_1166_65#_M1034_d N_A_1166_65#_M1012_d
+ N_A_1166_65#_M1022_d N_A_1166_65#_c_1205_n N_A_1166_65#_c_1206_n
+ N_A_1166_65#_c_1219_n N_A_1166_65#_c_1207_n N_A_1166_65#_c_1208_n
+ N_A_1166_65#_c_1209_n N_A_1166_65#_c_1210_n
+ PM_SKY130_FD_SC_LP__O311AI_4%A_1166_65#
cc_1 VNB N_A1_c_146_n 0.0210214f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.185
cc_2 VNB N_A1_M1005_g 0.0100771f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_3 VNB N_A1_c_148_n 0.0159015f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.185
cc_4 VNB N_A1_M1013_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_5 VNB N_A1_c_150_n 0.0159015f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.185
cc_6 VNB N_A1_M1027_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_7 VNB N_A1_c_152_n 0.0160911f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.185
cc_8 VNB N_A1_M1030_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_9 VNB A1 0.0258007f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_10 VNB N_A1_c_155_n 0.104237f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.35
cc_11 VNB N_A2_c_224_n 0.0160911f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.185
cc_12 VNB N_A2_M1001_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_13 VNB N_A2_c_226_n 0.0159015f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.185
cc_14 VNB N_A2_M1019_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_15 VNB N_A2_c_228_n 0.0159015f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.185
cc_16 VNB N_A2_M1024_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_17 VNB N_A2_c_230_n 0.0160871f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.185
cc_18 VNB N_A2_M1035_g 0.00841695f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_19 VNB A2 0.0174681f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_20 VNB N_A2_c_233_n 0.0761197f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.35
cc_21 VNB N_A3_M1007_g 0.0243989f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_22 VNB N_A3_c_319_n 0.0129075f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_23 VNB N_A3_M1009_g 0.0223448f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.655
cc_24 VNB N_A3_M1026_g 0.0227151f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_25 VNB N_A3_M1037_g 0.0302894f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.515
cc_26 VNB A3 0.00450904f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.35
cc_27 VNB N_A3_c_324_n 0.0172383f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.35
cc_28 VNB N_A3_c_325_n 0.0774649f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.307
cc_29 VNB N_B1_M1010_g 0.0252071f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_30 VNB N_B1_M1011_g 0.0190066f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_31 VNB N_B1_M1029_g 0.0197273f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_32 VNB N_B1_M1034_g 0.0200465f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_33 VNB N_B1_c_414_n 0.00143057f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.35
cc_34 VNB N_B1_c_415_n 0.0683021f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.35
cc_35 VNB N_C1_M1008_g 0.0206807f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_36 VNB N_C1_M1012_g 0.020608f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_37 VNB N_C1_M1017_g 0.0200852f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_38 VNB N_C1_M1022_g 0.0272763f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_39 VNB C1 0.0161608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_C1_c_487_n 0.104689f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.35
cc_41 VNB N_A_30_367#_c_561_n 0.00289786f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.185
cc_42 VNB N_A_30_367#_c_562_n 0.00395544f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_43 VNB N_A_30_367#_c_563_n 0.00330382f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_44 VNB N_A_30_367#_c_564_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.35
cc_45 VNB N_A_30_367#_c_565_n 0.00650216f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.35
cc_46 VNB N_A_30_367#_c_566_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.35
cc_47 VNB N_A_30_367#_c_567_n 0.00268362f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.35
cc_48 VNB N_A_30_367#_c_568_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.35
cc_49 VNB N_VPWR_c_637_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_Y_c_830_n 0.00244581f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_51 VNB N_Y_c_831_n 0.033814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_Y_c_832_n 0.00352222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_Y_c_833_n 0.00524921f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.35
cc_54 VNB N_Y_c_834_n 0.00244469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_969_n 0.0108441f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.185
cc_56 VNB N_VGND_c_970_n 0.032872f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_57 VNB N_VGND_c_971_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_972_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_59 VNB N_VGND_c_973_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_974_n 0.0123241f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.35
cc_61 VNB N_VGND_c_975_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.35
cc_62 VNB N_VGND_c_976_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.35
cc_63 VNB N_VGND_c_977_n 0.00619278f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.35
cc_64 VNB N_VGND_c_978_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_979_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.307
cc_66 VNB N_VGND_c_980_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_981_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_982_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_983_n 0.0117072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_984_n 0.0116838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_985_n 0.104723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_986_n 0.495754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_987_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_988_n 0.00436768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_989_n 0.00436768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_990_n 0.00510637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_113_47#_c_1114_n 0.00726499f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.307
cc_78 VNB N_A_1166_65#_c_1205_n 0.0116927f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_79 VNB N_A_1166_65#_c_1206_n 0.00295012f $X=-0.19 $Y=-0.245 $X2=1.78
+ $Y2=0.655
cc_80 VNB N_A_1166_65#_c_1207_n 0.00787259f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_81 VNB N_A_1166_65#_c_1208_n 0.00299464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1166_65#_c_1209_n 0.00211003f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.35
cc_83 VNB N_A_1166_65#_c_1210_n 0.00218279f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.35
cc_84 VPB N_A1_M1005_g 0.0232847f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_85 VPB N_A1_M1013_g 0.0185652f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_86 VPB N_A1_M1027_g 0.0185652f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_87 VPB N_A1_M1030_g 0.018727f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_88 VPB N_A2_M1001_g 0.0189261f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_89 VPB N_A2_M1019_g 0.0187643f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_90 VPB N_A2_M1024_g 0.0187643f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_91 VPB N_A2_M1035_g 0.0233896f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_92 VPB N_A3_M1014_g 0.0217292f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_93 VPB N_A3_M1020_g 0.0181349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A3_M1031_g 0.0181378f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_95 VPB N_A3_M1036_g 0.0183424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB A3 0.011112f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.35
cc_97 VPB N_A3_c_325_n 0.0153062f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.307
cc_98 VPB N_B1_c_416_n 0.016229f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.185
cc_99 VPB N_B1_c_417_n 0.015814f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.185
cc_100 VPB N_B1_c_418_n 0.015814f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.185
cc_101 VPB N_B1_c_419_n 0.016015f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=1.185
cc_102 VPB N_B1_c_414_n 0.00908534f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.35
cc_103 VPB N_B1_c_415_n 0.0236623f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.35
cc_104 VPB N_C1_c_488_n 0.016015f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.185
cc_105 VPB N_C1_c_489_n 0.015814f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.185
cc_106 VPB N_C1_c_490_n 0.015814f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.185
cc_107 VPB N_C1_c_491_n 0.0213619f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=1.185
cc_108 VPB C1 0.0312304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_C1_c_487_n 0.0402339f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=1.35
cc_110 VPB N_A_30_367#_c_569_n 0.0498589f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.515
cc_111 VPB N_A_30_367#_c_561_n 0.00559032f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=1.185
cc_112 VPB N_A_30_367#_c_562_n 0.0054421f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=0.655
cc_113 VPB N_A_30_367#_c_572_n 9.96097e-19 $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_114 VPB N_A_30_367#_c_563_n 0.00559032f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_115 VPB N_A_30_367#_c_574_n 9.96097e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_30_367#_c_564_n 0.00559032f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.35
cc_117 VPB N_A_30_367#_c_576_n 9.96097e-19 $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.35
cc_118 VPB N_A_30_367#_c_565_n 0.00706527f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.35
cc_119 VPB N_A_30_367#_c_578_n 0.00968f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.35
cc_120 VPB N_VPWR_c_638_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_639_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_122 VPB N_VPWR_c_640_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_641_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.35
cc_124 VPB N_VPWR_c_642_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.35
cc_125 VPB N_VPWR_c_643_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.35
cc_126 VPB N_VPWR_c_644_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.35
cc_127 VPB N_VPWR_c_645_n 0.104084f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.35
cc_128 VPB N_VPWR_c_646_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.35
cc_129 VPB N_VPWR_c_647_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_648_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.307
cc_131 VPB N_VPWR_c_649_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_650_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_651_n 0.0158404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_652_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_653_n 0.028582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_637_n 0.0661721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_655_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_656_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_657_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_457_367#_c_774_n 0.0113537f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=0.655
cc_141 VPB N_Y_c_830_n 0.00349393f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_142 VPB N_Y_c_836_n 0.00588761f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_143 VPB N_Y_c_837_n 0.00743012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_Y_c_838_n 0.0373194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_Y_c_839_n 0.00184265f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 N_A1_c_152_n N_A2_c_224_n 0.024785f $X=1.78 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_147 A1 N_A2_c_224_n 7.86898e-19 $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_148 N_A1_M1030_g N_A2_M1001_g 0.024785f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A1_c_152_n A2 9.92942e-19 $X=1.78 $Y=1.185 $X2=0 $Y2=0
cc_150 A1 A2 0.0236984f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_151 N_A1_c_155_n N_A2_c_233_n 0.024785f $X=1.78 $Y=1.35 $X2=0 $Y2=0
cc_152 N_A1_M1005_g N_A_30_367#_c_569_n 0.0046421f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A1_M1005_g N_A_30_367#_c_561_n 0.0157274f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A1_M1013_g N_A_30_367#_c_561_n 0.0143398f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_155 A1 N_A_30_367#_c_561_n 0.0481851f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A1_c_155_n N_A_30_367#_c_561_n 0.00357126f $X=1.78 $Y=1.35 $X2=0 $Y2=0
cc_157 A1 N_A_30_367#_c_562_n 0.0217644f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A1_c_155_n N_A_30_367#_c_562_n 0.00526356f $X=1.78 $Y=1.35 $X2=0 $Y2=0
cc_159 N_A1_M1013_g N_A_30_367#_c_572_n 0.0014373f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A1_M1027_g N_A_30_367#_c_572_n 0.0014373f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A1_M1027_g N_A_30_367#_c_563_n 0.0143398f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A1_M1030_g N_A_30_367#_c_563_n 0.0142932f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_163 A1 N_A_30_367#_c_563_n 0.0452949f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A1_c_155_n N_A_30_367#_c_563_n 0.00246472f $X=1.78 $Y=1.35 $X2=0 $Y2=0
cc_165 N_A1_M1030_g N_A_30_367#_c_574_n 0.0014373f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_166 A1 N_A_30_367#_c_566_n 0.0157467f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_167 N_A1_c_155_n N_A_30_367#_c_566_n 0.00256759f $X=1.78 $Y=1.35 $X2=0 $Y2=0
cc_168 N_A1_M1005_g N_VPWR_c_638_n 0.0194824f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A1_M1013_g N_VPWR_c_638_n 0.01742f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A1_M1027_g N_VPWR_c_638_n 7.69607e-19 $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A1_M1013_g N_VPWR_c_639_n 7.69607e-19 $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A1_M1027_g N_VPWR_c_639_n 0.01742f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A1_M1030_g N_VPWR_c_639_n 0.0186126f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A1_M1030_g N_VPWR_c_645_n 0.00486043f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A1_M1005_g N_VPWR_c_651_n 0.00486043f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A1_M1013_g N_VPWR_c_652_n 0.00486043f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A1_M1027_g N_VPWR_c_652_n 0.00486043f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A1_M1005_g N_VPWR_c_637_n 0.00919377f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A1_M1013_g N_VPWR_c_637_n 0.00824727f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A1_M1027_g N_VPWR_c_637_n 0.00824727f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A1_M1030_g N_VPWR_c_637_n 0.0082726f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A1_c_146_n N_VGND_c_970_n 0.0152201f $X=0.49 $Y=1.185 $X2=0 $Y2=0
cc_183 N_A1_c_148_n N_VGND_c_970_n 6.15704e-19 $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_184 A1 N_VGND_c_970_n 0.0252165f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A1_c_155_n N_VGND_c_970_n 0.00178271f $X=1.78 $Y=1.35 $X2=0 $Y2=0
cc_186 N_A1_c_146_n N_VGND_c_971_n 5.67328e-19 $X=0.49 $Y=1.185 $X2=0 $Y2=0
cc_187 N_A1_c_148_n N_VGND_c_971_n 0.00990604f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_188 N_A1_c_150_n N_VGND_c_971_n 0.00990604f $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_189 N_A1_c_152_n N_VGND_c_971_n 5.67328e-19 $X=1.78 $Y=1.185 $X2=0 $Y2=0
cc_190 N_A1_c_150_n N_VGND_c_972_n 5.67328e-19 $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_191 N_A1_c_152_n N_VGND_c_972_n 0.00983814f $X=1.78 $Y=1.185 $X2=0 $Y2=0
cc_192 N_A1_c_150_n N_VGND_c_978_n 0.00486043f $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_193 N_A1_c_152_n N_VGND_c_978_n 0.00486043f $X=1.78 $Y=1.185 $X2=0 $Y2=0
cc_194 N_A1_c_146_n N_VGND_c_982_n 0.00486043f $X=0.49 $Y=1.185 $X2=0 $Y2=0
cc_195 N_A1_c_148_n N_VGND_c_982_n 0.00486043f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_196 N_A1_c_146_n N_VGND_c_986_n 0.00824727f $X=0.49 $Y=1.185 $X2=0 $Y2=0
cc_197 N_A1_c_148_n N_VGND_c_986_n 0.00454119f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_198 N_A1_c_150_n N_VGND_c_986_n 0.00454119f $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_199 N_A1_c_152_n N_VGND_c_986_n 0.00454119f $X=1.78 $Y=1.185 $X2=0 $Y2=0
cc_200 N_A1_c_148_n N_A_113_47#_c_1115_n 0.00973732f $X=0.92 $Y=1.185 $X2=0
+ $Y2=0
cc_201 N_A1_c_150_n N_A_113_47#_c_1115_n 0.00969075f $X=1.35 $Y=1.185 $X2=0
+ $Y2=0
cc_202 A1 N_A_113_47#_c_1115_n 0.0417635f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A1_c_155_n N_A_113_47#_c_1115_n 6.95778e-19 $X=1.78 $Y=1.35 $X2=0 $Y2=0
cc_204 A1 N_A_113_47#_c_1119_n 0.0150898f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_205 N_A1_c_155_n N_A_113_47#_c_1119_n 7.81868e-19 $X=1.78 $Y=1.35 $X2=0 $Y2=0
cc_206 N_A1_c_152_n N_A_113_47#_c_1121_n 0.00969075f $X=1.78 $Y=1.185 $X2=0
+ $Y2=0
cc_207 A1 N_A_113_47#_c_1121_n 0.012462f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_208 A1 N_A_113_47#_c_1123_n 0.0150898f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_209 N_A1_c_155_n N_A_113_47#_c_1123_n 7.81868e-19 $X=1.78 $Y=1.35 $X2=0 $Y2=0
cc_210 N_A2_c_230_n N_A3_M1007_g 0.0226619f $X=3.5 $Y=1.185 $X2=0 $Y2=0
cc_211 A2 N_A3_M1007_g 0.00274906f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_212 N_A2_c_233_n N_A3_c_319_n 0.0226619f $X=3.5 $Y=1.35 $X2=0 $Y2=0
cc_213 N_A2_c_233_n N_A3_c_325_n 0.00179648f $X=3.5 $Y=1.35 $X2=0 $Y2=0
cc_214 N_A2_M1001_g N_A_30_367#_c_574_n 0.0014373f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A2_M1001_g N_A_30_367#_c_564_n 0.0142932f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A2_M1019_g N_A_30_367#_c_564_n 0.0143398f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_217 A2 N_A_30_367#_c_564_n 0.0483649f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_218 N_A2_c_233_n N_A_30_367#_c_564_n 0.00246472f $X=3.5 $Y=1.35 $X2=0 $Y2=0
cc_219 N_A2_M1019_g N_A_30_367#_c_576_n 0.00165214f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A2_M1024_g N_A_30_367#_c_576_n 0.00165214f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A2_M1024_g N_A_30_367#_c_565_n 0.0143398f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A2_M1035_g N_A_30_367#_c_565_n 0.0155114f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_223 A2 N_A_30_367#_c_565_n 0.0635656f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_224 N_A2_c_233_n N_A_30_367#_c_565_n 0.00246472f $X=3.5 $Y=1.35 $X2=0 $Y2=0
cc_225 N_A2_M1035_g N_A_30_367#_c_578_n 0.00561046f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_226 A2 N_A_30_367#_c_567_n 0.00521166f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_227 A2 N_A_30_367#_c_568_n 0.0157467f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A2_c_233_n N_A_30_367#_c_568_n 0.00256759f $X=3.5 $Y=1.35 $X2=0 $Y2=0
cc_229 N_A2_M1001_g N_VPWR_c_639_n 0.00141193f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A2_M1001_g N_VPWR_c_645_n 0.00547432f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A2_M1019_g N_VPWR_c_645_n 0.00357842f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A2_M1024_g N_VPWR_c_645_n 0.00357842f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A2_M1035_g N_VPWR_c_645_n 0.00357842f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A2_M1001_g N_VPWR_c_637_n 0.00990114f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A2_M1019_g N_VPWR_c_637_n 0.00535118f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A2_M1024_g N_VPWR_c_637_n 0.00535118f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A2_M1035_g N_VPWR_c_637_n 0.00675085f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A2_M1001_g N_A_457_367#_c_775_n 0.00193114f $X=2.21 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A2_M1019_g N_A_457_367#_c_775_n 5.89773e-19 $X=2.64 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_A2_M1001_g N_A_457_367#_c_777_n 0.0117092f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_241 N_A2_M1019_g N_A_457_367#_c_777_n 0.0129502f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_242 N_A2_M1024_g N_A_457_367#_c_777_n 6.58347e-19 $X=3.07 $Y=2.465 $X2=0
+ $Y2=0
cc_243 N_A2_M1019_g N_A_457_367#_c_780_n 0.0105205f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A2_M1024_g N_A_457_367#_c_780_n 0.0105205f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A2_M1019_g N_A_457_367#_c_782_n 6.58347e-19 $X=2.64 $Y=2.465 $X2=0
+ $Y2=0
cc_246 N_A2_M1024_g N_A_457_367#_c_782_n 0.0129502f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_247 N_A2_M1035_g N_A_457_367#_c_782_n 0.0177589f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A2_M1035_g N_A_457_367#_c_774_n 0.0125611f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A2_M1024_g N_A_457_367#_c_786_n 5.89773e-19 $X=3.07 $Y=2.465 $X2=0
+ $Y2=0
cc_250 N_A2_M1035_g N_A_457_367#_c_786_n 5.89773e-19 $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A2_M1035_g N_Y_c_830_n 7.48373e-19 $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_252 A2 N_Y_c_830_n 0.0103113f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_253 N_A2_c_233_n N_Y_c_830_n 0.00226299f $X=3.5 $Y=1.35 $X2=0 $Y2=0
cc_254 A2 N_Y_c_832_n 0.00481566f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_255 N_A2_c_224_n N_VGND_c_972_n 0.00983814f $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_256 N_A2_c_226_n N_VGND_c_972_n 5.67328e-19 $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_257 N_A2_c_224_n N_VGND_c_973_n 5.67328e-19 $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_258 N_A2_c_226_n N_VGND_c_973_n 0.00990604f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_259 N_A2_c_228_n N_VGND_c_973_n 0.00990604f $X=3.07 $Y=1.185 $X2=0 $Y2=0
cc_260 N_A2_c_230_n N_VGND_c_973_n 5.67328e-19 $X=3.5 $Y=1.185 $X2=0 $Y2=0
cc_261 N_A2_c_228_n N_VGND_c_974_n 0.00486043f $X=3.07 $Y=1.185 $X2=0 $Y2=0
cc_262 N_A2_c_230_n N_VGND_c_974_n 0.00366311f $X=3.5 $Y=1.185 $X2=0 $Y2=0
cc_263 N_A2_c_228_n N_VGND_c_975_n 5.40452e-19 $X=3.07 $Y=1.185 $X2=0 $Y2=0
cc_264 N_A2_c_230_n N_VGND_c_975_n 0.00776046f $X=3.5 $Y=1.185 $X2=0 $Y2=0
cc_265 N_A2_c_224_n N_VGND_c_980_n 0.00486043f $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_266 N_A2_c_226_n N_VGND_c_980_n 0.00486043f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_267 N_A2_c_224_n N_VGND_c_986_n 0.00454119f $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_268 N_A2_c_226_n N_VGND_c_986_n 0.00454119f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_269 N_A2_c_228_n N_VGND_c_986_n 0.00454119f $X=3.07 $Y=1.185 $X2=0 $Y2=0
cc_270 N_A2_c_230_n N_VGND_c_986_n 0.00434326f $X=3.5 $Y=1.185 $X2=0 $Y2=0
cc_271 N_A2_c_224_n N_A_113_47#_c_1121_n 0.00969075f $X=2.21 $Y=1.185 $X2=0
+ $Y2=0
cc_272 A2 N_A_113_47#_c_1121_n 0.0182093f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_273 N_A2_c_226_n N_A_113_47#_c_1127_n 0.00973732f $X=2.64 $Y=1.185 $X2=0
+ $Y2=0
cc_274 N_A2_c_228_n N_A_113_47#_c_1127_n 0.00973732f $X=3.07 $Y=1.185 $X2=0
+ $Y2=0
cc_275 A2 N_A_113_47#_c_1127_n 0.0417635f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_276 N_A2_c_233_n N_A_113_47#_c_1127_n 6.95778e-19 $X=3.5 $Y=1.35 $X2=0 $Y2=0
cc_277 N_A2_c_230_n N_A_113_47#_c_1131_n 0.0123724f $X=3.5 $Y=1.185 $X2=0 $Y2=0
cc_278 A2 N_A_113_47#_c_1131_n 0.0263744f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_279 A2 N_A_113_47#_c_1133_n 0.00134701f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_280 A2 N_A_113_47#_c_1134_n 0.0150898f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_281 N_A2_c_233_n N_A_113_47#_c_1134_n 7.81868e-19 $X=3.5 $Y=1.35 $X2=0 $Y2=0
cc_282 A2 N_A_113_47#_c_1136_n 0.0150898f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_283 N_A2_c_233_n N_A_113_47#_c_1136_n 7.81868e-19 $X=3.5 $Y=1.35 $X2=0 $Y2=0
cc_284 N_A3_M1036_g N_B1_c_416_n 0.0114566f $X=5.75 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_285 A3 N_B1_c_414_n 0.0289001f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_286 A3 N_B1_c_415_n 0.00345042f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_287 N_A3_c_325_n N_B1_c_415_n 0.0228959f $X=5.75 $Y=1.51 $X2=0 $Y2=0
cc_288 N_A3_c_319_n N_A_30_367#_c_565_n 8.9861e-19 $X=4.005 $Y=1.42 $X2=0 $Y2=0
cc_289 N_A3_c_325_n N_A_30_367#_c_565_n 2.27638e-19 $X=5.75 $Y=1.51 $X2=0 $Y2=0
cc_290 N_A3_M1036_g N_VPWR_c_640_n 0.00131432f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A3_M1014_g N_VPWR_c_645_n 0.00357842f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A3_M1020_g N_VPWR_c_645_n 0.00357842f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A3_M1031_g N_VPWR_c_645_n 0.00357842f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A3_M1036_g N_VPWR_c_645_n 0.00547432f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_295 N_A3_M1014_g N_VPWR_c_637_n 0.00675085f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_296 N_A3_M1020_g N_VPWR_c_637_n 0.00535118f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A3_M1031_g N_VPWR_c_637_n 0.00535118f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A3_M1036_g N_VPWR_c_637_n 0.00990114f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A3_M1014_g N_A_457_367#_c_774_n 0.0125611f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A3_M1014_g N_A_457_367#_c_789_n 0.0141439f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A3_M1020_g N_A_457_367#_c_789_n 0.00952429f $X=4.89 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_A3_M1031_g N_A_457_367#_c_789_n 5.60744e-19 $X=5.32 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A3_M1020_g N_A_457_367#_c_792_n 0.0105205f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A3_M1031_g N_A_457_367#_c_792_n 0.0111103f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A3_M1036_g N_A_457_367#_c_792_n 0.00193114f $X=5.75 $Y=2.465 $X2=0
+ $Y2=0
cc_306 N_A3_M1020_g N_A_457_367#_c_795_n 5.60744e-19 $X=4.89 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A3_M1031_g N_A_457_367#_c_795_n 0.00952429f $X=5.32 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A3_M1036_g N_A_457_367#_c_795_n 0.00828328f $X=5.75 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A3_M1014_g N_A_457_367#_c_798_n 5.89773e-19 $X=4.46 $Y=2.465 $X2=0
+ $Y2=0
cc_310 N_A3_M1020_g N_A_457_367#_c_798_n 5.89773e-19 $X=4.89 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A3_M1007_g N_Y_c_830_n 7.56191e-19 $X=3.93 $Y=0.655 $X2=0 $Y2=0
cc_312 N_A3_M1009_g N_Y_c_830_n 0.00220818f $X=4.36 $Y=0.655 $X2=0 $Y2=0
cc_313 N_A3_M1014_g N_Y_c_830_n 0.00652606f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A3_M1026_g N_Y_c_830_n 4.21966e-19 $X=4.79 $Y=0.655 $X2=0 $Y2=0
cc_315 A3 N_Y_c_830_n 0.0252521f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_316 N_A3_c_324_n N_Y_c_830_n 0.0120123f $X=4.285 $Y=1.51 $X2=0 $Y2=0
cc_317 N_A3_c_325_n N_Y_c_830_n 0.010376f $X=5.75 $Y=1.51 $X2=0 $Y2=0
cc_318 N_A3_M1009_g N_Y_c_831_n 0.00974903f $X=4.36 $Y=0.655 $X2=0 $Y2=0
cc_319 N_A3_M1026_g N_Y_c_831_n 0.010446f $X=4.79 $Y=0.655 $X2=0 $Y2=0
cc_320 N_A3_M1037_g N_Y_c_831_n 0.0125331f $X=5.22 $Y=0.655 $X2=0 $Y2=0
cc_321 A3 N_Y_c_831_n 0.122352f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_322 N_A3_c_325_n N_Y_c_831_n 0.0207003f $X=5.75 $Y=1.51 $X2=0 $Y2=0
cc_323 N_A3_M1007_g N_Y_c_832_n 0.00369874f $X=3.93 $Y=0.655 $X2=0 $Y2=0
cc_324 N_A3_M1009_g N_Y_c_832_n 0.00177864f $X=4.36 $Y=0.655 $X2=0 $Y2=0
cc_325 N_A3_c_325_n N_Y_c_839_n 0.00128908f $X=5.75 $Y=1.51 $X2=0 $Y2=0
cc_326 A3 Y 0.0153757f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_327 N_A3_c_325_n Y 6.4545e-19 $X=5.75 $Y=1.51 $X2=0 $Y2=0
cc_328 A3 Y 0.0153758f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_329 N_A3_M1014_g N_Y_c_862_n 0.0143082f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_330 N_A3_M1020_g N_Y_c_862_n 0.0131606f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_331 A3 N_Y_c_862_n 0.0355229f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_332 N_A3_c_325_n N_Y_c_862_n 5.78018e-19 $X=5.75 $Y=1.51 $X2=0 $Y2=0
cc_333 N_A3_M1031_g N_Y_c_866_n 0.0131606f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A3_M1036_g N_Y_c_866_n 0.0131606f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_335 A3 N_Y_c_866_n 0.043132f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_336 N_A3_c_325_n N_Y_c_866_n 5.8554e-19 $X=5.75 $Y=1.51 $X2=0 $Y2=0
cc_337 N_A3_M1007_g N_VGND_c_975_n 0.00775945f $X=3.93 $Y=0.655 $X2=0 $Y2=0
cc_338 N_A3_M1009_g N_VGND_c_975_n 5.40452e-19 $X=4.36 $Y=0.655 $X2=0 $Y2=0
cc_339 N_A3_M1007_g N_VGND_c_976_n 5.40452e-19 $X=3.93 $Y=0.655 $X2=0 $Y2=0
cc_340 N_A3_M1009_g N_VGND_c_976_n 0.00780203f $X=4.36 $Y=0.655 $X2=0 $Y2=0
cc_341 N_A3_M1026_g N_VGND_c_976_n 0.00780203f $X=4.79 $Y=0.655 $X2=0 $Y2=0
cc_342 N_A3_M1037_g N_VGND_c_976_n 5.40452e-19 $X=5.22 $Y=0.655 $X2=0 $Y2=0
cc_343 N_A3_M1026_g N_VGND_c_977_n 5.34794e-19 $X=4.79 $Y=0.655 $X2=0 $Y2=0
cc_344 N_A3_M1037_g N_VGND_c_977_n 0.00863329f $X=5.22 $Y=0.655 $X2=0 $Y2=0
cc_345 N_A3_M1007_g N_VGND_c_983_n 0.003662f $X=3.93 $Y=0.655 $X2=0 $Y2=0
cc_346 N_A3_M1009_g N_VGND_c_983_n 0.00366311f $X=4.36 $Y=0.655 $X2=0 $Y2=0
cc_347 N_A3_M1026_g N_VGND_c_984_n 0.00366311f $X=4.79 $Y=0.655 $X2=0 $Y2=0
cc_348 N_A3_M1037_g N_VGND_c_984_n 0.00364083f $X=5.22 $Y=0.655 $X2=0 $Y2=0
cc_349 N_A3_M1007_g N_VGND_c_986_n 0.00434118f $X=3.93 $Y=0.655 $X2=0 $Y2=0
cc_350 N_A3_M1009_g N_VGND_c_986_n 0.00434326f $X=4.36 $Y=0.655 $X2=0 $Y2=0
cc_351 N_A3_M1026_g N_VGND_c_986_n 0.00434326f $X=4.79 $Y=0.655 $X2=0 $Y2=0
cc_352 N_A3_M1037_g N_VGND_c_986_n 0.00430165f $X=5.22 $Y=0.655 $X2=0 $Y2=0
cc_353 N_A3_M1009_g N_A_113_47#_c_1138_n 0.0099311f $X=4.36 $Y=0.655 $X2=0 $Y2=0
cc_354 N_A3_M1026_g N_A_113_47#_c_1138_n 0.00993147f $X=4.79 $Y=0.655 $X2=0
+ $Y2=0
cc_355 N_A3_M1007_g N_A_113_47#_c_1133_n 0.016986f $X=3.93 $Y=0.655 $X2=0 $Y2=0
cc_356 N_A3_c_324_n N_A_113_47#_c_1133_n 4.46852e-19 $X=4.285 $Y=1.51 $X2=0
+ $Y2=0
cc_357 N_A3_M1037_g N_A_113_47#_c_1114_n 0.0126834f $X=5.22 $Y=0.655 $X2=0 $Y2=0
cc_358 N_B1_c_419_n N_C1_c_488_n 0.0092982f $X=7.47 $Y=1.725 $X2=-0.19
+ $Y2=-0.245
cc_359 N_B1_M1034_g N_C1_M1008_g 0.0203165f $X=7.54 $Y=0.745 $X2=0 $Y2=0
cc_360 N_B1_c_414_n C1 0.0291311f $X=7.45 $Y=1.51 $X2=0 $Y2=0
cc_361 N_B1_c_415_n C1 0.00118521f $X=7.47 $Y=1.535 $X2=0 $Y2=0
cc_362 N_B1_c_414_n N_C1_c_487_n 5.48153e-19 $X=7.45 $Y=1.51 $X2=0 $Y2=0
cc_363 N_B1_c_415_n N_C1_c_487_n 0.0323575f $X=7.47 $Y=1.535 $X2=0 $Y2=0
cc_364 N_B1_c_416_n N_VPWR_c_640_n 0.0156682f $X=6.18 $Y=1.725 $X2=0 $Y2=0
cc_365 N_B1_c_417_n N_VPWR_c_640_n 0.0144755f $X=6.61 $Y=1.725 $X2=0 $Y2=0
cc_366 N_B1_c_418_n N_VPWR_c_640_n 6.72004e-19 $X=7.04 $Y=1.725 $X2=0 $Y2=0
cc_367 N_B1_c_417_n N_VPWR_c_641_n 6.80491e-19 $X=6.61 $Y=1.725 $X2=0 $Y2=0
cc_368 N_B1_c_418_n N_VPWR_c_641_n 0.0151398f $X=7.04 $Y=1.725 $X2=0 $Y2=0
cc_369 N_B1_c_419_n N_VPWR_c_641_n 0.0151398f $X=7.47 $Y=1.725 $X2=0 $Y2=0
cc_370 N_B1_c_419_n N_VPWR_c_642_n 6.80491e-19 $X=7.47 $Y=1.725 $X2=0 $Y2=0
cc_371 N_B1_c_416_n N_VPWR_c_645_n 0.00486043f $X=6.18 $Y=1.725 $X2=0 $Y2=0
cc_372 N_B1_c_417_n N_VPWR_c_647_n 0.00486043f $X=6.61 $Y=1.725 $X2=0 $Y2=0
cc_373 N_B1_c_418_n N_VPWR_c_647_n 0.00486043f $X=7.04 $Y=1.725 $X2=0 $Y2=0
cc_374 N_B1_c_419_n N_VPWR_c_649_n 0.00486043f $X=7.47 $Y=1.725 $X2=0 $Y2=0
cc_375 N_B1_c_416_n N_VPWR_c_637_n 0.0082726f $X=6.18 $Y=1.725 $X2=0 $Y2=0
cc_376 N_B1_c_417_n N_VPWR_c_637_n 0.00824727f $X=6.61 $Y=1.725 $X2=0 $Y2=0
cc_377 N_B1_c_418_n N_VPWR_c_637_n 0.00824727f $X=7.04 $Y=1.725 $X2=0 $Y2=0
cc_378 N_B1_c_419_n N_VPWR_c_637_n 0.0082726f $X=7.47 $Y=1.725 $X2=0 $Y2=0
cc_379 N_B1_M1010_g N_Y_c_831_n 0.0147266f $X=6.19 $Y=0.745 $X2=0 $Y2=0
cc_380 N_B1_M1011_g N_Y_c_831_n 0.0104926f $X=6.62 $Y=0.745 $X2=0 $Y2=0
cc_381 N_B1_M1029_g N_Y_c_831_n 0.0108341f $X=7.05 $Y=0.745 $X2=0 $Y2=0
cc_382 N_B1_M1034_g N_Y_c_831_n 0.012434f $X=7.54 $Y=0.745 $X2=0 $Y2=0
cc_383 N_B1_c_414_n N_Y_c_831_n 0.0996643f $X=7.45 $Y=1.51 $X2=0 $Y2=0
cc_384 N_B1_c_415_n N_Y_c_831_n 0.00971487f $X=7.47 $Y=1.535 $X2=0 $Y2=0
cc_385 N_B1_c_418_n N_Y_c_876_n 0.0122595f $X=7.04 $Y=1.725 $X2=0 $Y2=0
cc_386 N_B1_c_419_n N_Y_c_876_n 0.0122595f $X=7.47 $Y=1.725 $X2=0 $Y2=0
cc_387 N_B1_c_414_n N_Y_c_876_n 0.0427275f $X=7.45 $Y=1.51 $X2=0 $Y2=0
cc_388 N_B1_c_415_n N_Y_c_876_n 6.55157e-19 $X=7.47 $Y=1.535 $X2=0 $Y2=0
cc_389 N_B1_c_416_n N_Y_c_880_n 0.0152789f $X=6.18 $Y=1.725 $X2=0 $Y2=0
cc_390 N_B1_c_417_n N_Y_c_880_n 0.0131606f $X=6.61 $Y=1.725 $X2=0 $Y2=0
cc_391 N_B1_c_414_n N_Y_c_880_n 0.0300546f $X=7.45 $Y=1.51 $X2=0 $Y2=0
cc_392 N_B1_c_415_n N_Y_c_880_n 6.63131e-19 $X=7.47 $Y=1.535 $X2=0 $Y2=0
cc_393 N_B1_c_414_n N_Y_c_884_n 0.0153756f $X=7.45 $Y=1.51 $X2=0 $Y2=0
cc_394 N_B1_c_415_n N_Y_c_884_n 7.3774e-19 $X=7.47 $Y=1.535 $X2=0 $Y2=0
cc_395 N_B1_c_414_n N_Y_c_886_n 0.00162626f $X=7.45 $Y=1.51 $X2=0 $Y2=0
cc_396 N_B1_M1010_g N_VGND_c_977_n 0.0016998f $X=6.19 $Y=0.745 $X2=0 $Y2=0
cc_397 N_B1_M1010_g N_VGND_c_985_n 0.00302501f $X=6.19 $Y=0.745 $X2=0 $Y2=0
cc_398 N_B1_M1011_g N_VGND_c_985_n 0.00302501f $X=6.62 $Y=0.745 $X2=0 $Y2=0
cc_399 N_B1_M1029_g N_VGND_c_985_n 0.00302501f $X=7.05 $Y=0.745 $X2=0 $Y2=0
cc_400 N_B1_M1034_g N_VGND_c_985_n 0.00302484f $X=7.54 $Y=0.745 $X2=0 $Y2=0
cc_401 N_B1_M1010_g N_VGND_c_986_n 0.0048466f $X=6.19 $Y=0.745 $X2=0 $Y2=0
cc_402 N_B1_M1011_g N_VGND_c_986_n 0.00434671f $X=6.62 $Y=0.745 $X2=0 $Y2=0
cc_403 N_B1_M1029_g N_VGND_c_986_n 0.00440366f $X=7.05 $Y=0.745 $X2=0 $Y2=0
cc_404 N_B1_M1034_g N_VGND_c_986_n 0.00442265f $X=7.54 $Y=0.745 $X2=0 $Y2=0
cc_405 N_B1_M1010_g N_A_113_47#_c_1114_n 0.0112524f $X=6.19 $Y=0.745 $X2=0 $Y2=0
cc_406 N_B1_M1011_g N_A_113_47#_c_1114_n 0.0089689f $X=6.62 $Y=0.745 $X2=0 $Y2=0
cc_407 N_B1_M1029_g N_A_113_47#_c_1114_n 0.0089689f $X=7.05 $Y=0.745 $X2=0 $Y2=0
cc_408 N_B1_M1010_g N_A_1166_65#_c_1205_n 0.0121603f $X=6.19 $Y=0.745 $X2=0
+ $Y2=0
cc_409 N_B1_M1011_g N_A_1166_65#_c_1205_n 0.0115987f $X=6.62 $Y=0.745 $X2=0
+ $Y2=0
cc_410 N_B1_M1029_g N_A_1166_65#_c_1205_n 0.0122044f $X=7.05 $Y=0.745 $X2=0
+ $Y2=0
cc_411 N_B1_M1034_g N_A_1166_65#_c_1205_n 0.0122882f $X=7.54 $Y=0.745 $X2=0
+ $Y2=0
cc_412 N_B1_M1029_g N_A_1166_65#_c_1209_n 5.64826e-19 $X=7.05 $Y=0.745 $X2=0
+ $Y2=0
cc_413 N_B1_M1034_g N_A_1166_65#_c_1209_n 0.00642323f $X=7.54 $Y=0.745 $X2=0
+ $Y2=0
cc_414 N_C1_c_488_n N_VPWR_c_641_n 6.80491e-19 $X=7.9 $Y=1.725 $X2=0 $Y2=0
cc_415 N_C1_c_488_n N_VPWR_c_642_n 0.0151398f $X=7.9 $Y=1.725 $X2=0 $Y2=0
cc_416 N_C1_c_489_n N_VPWR_c_642_n 0.0151398f $X=8.33 $Y=1.725 $X2=0 $Y2=0
cc_417 N_C1_c_490_n N_VPWR_c_642_n 6.80491e-19 $X=8.76 $Y=1.725 $X2=0 $Y2=0
cc_418 N_C1_c_489_n N_VPWR_c_643_n 0.00486043f $X=8.33 $Y=1.725 $X2=0 $Y2=0
cc_419 N_C1_c_490_n N_VPWR_c_643_n 0.00486043f $X=8.76 $Y=1.725 $X2=0 $Y2=0
cc_420 N_C1_c_489_n N_VPWR_c_644_n 6.80491e-19 $X=8.33 $Y=1.725 $X2=0 $Y2=0
cc_421 N_C1_c_490_n N_VPWR_c_644_n 0.0151398f $X=8.76 $Y=1.725 $X2=0 $Y2=0
cc_422 N_C1_c_491_n N_VPWR_c_644_n 0.0170297f $X=9.19 $Y=1.725 $X2=0 $Y2=0
cc_423 N_C1_c_488_n N_VPWR_c_649_n 0.00486043f $X=7.9 $Y=1.725 $X2=0 $Y2=0
cc_424 N_C1_c_491_n N_VPWR_c_653_n 0.00486043f $X=9.19 $Y=1.725 $X2=0 $Y2=0
cc_425 N_C1_c_488_n N_VPWR_c_637_n 0.0082726f $X=7.9 $Y=1.725 $X2=0 $Y2=0
cc_426 N_C1_c_489_n N_VPWR_c_637_n 0.00824727f $X=8.33 $Y=1.725 $X2=0 $Y2=0
cc_427 N_C1_c_490_n N_VPWR_c_637_n 0.00824727f $X=8.76 $Y=1.725 $X2=0 $Y2=0
cc_428 N_C1_c_491_n N_VPWR_c_637_n 0.00954696f $X=9.19 $Y=1.725 $X2=0 $Y2=0
cc_429 N_C1_M1008_g N_Y_c_831_n 0.0129936f $X=7.98 $Y=0.745 $X2=0 $Y2=0
cc_430 C1 N_Y_c_831_n 0.0232124f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_431 N_C1_c_487_n N_Y_c_831_n 0.00231562f $X=9.48 $Y=1.535 $X2=0 $Y2=0
cc_432 N_C1_c_488_n N_Y_c_890_n 0.0122595f $X=7.9 $Y=1.725 $X2=0 $Y2=0
cc_433 N_C1_c_489_n N_Y_c_890_n 0.0122595f $X=8.33 $Y=1.725 $X2=0 $Y2=0
cc_434 C1 N_Y_c_890_n 0.0425198f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_435 N_C1_c_487_n N_Y_c_890_n 6.5019e-19 $X=9.48 $Y=1.535 $X2=0 $Y2=0
cc_436 N_C1_M1012_g N_Y_c_833_n 0.0120547f $X=8.53 $Y=0.745 $X2=0 $Y2=0
cc_437 N_C1_M1017_g N_Y_c_833_n 0.0128627f $X=8.98 $Y=0.745 $X2=0 $Y2=0
cc_438 N_C1_M1022_g N_Y_c_833_n 0.0058102f $X=9.48 $Y=0.745 $X2=0 $Y2=0
cc_439 C1 N_Y_c_833_n 0.0767221f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_440 N_C1_c_487_n N_Y_c_833_n 0.00834269f $X=9.48 $Y=1.535 $X2=0 $Y2=0
cc_441 N_C1_c_490_n N_Y_c_899_n 0.0122595f $X=8.76 $Y=1.725 $X2=0 $Y2=0
cc_442 N_C1_c_491_n N_Y_c_899_n 0.0122595f $X=9.19 $Y=1.725 $X2=0 $Y2=0
cc_443 C1 N_Y_c_899_n 0.0427275f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_444 N_C1_c_487_n N_Y_c_899_n 6.48771e-19 $X=9.48 $Y=1.535 $X2=0 $Y2=0
cc_445 N_C1_M1022_g N_Y_c_903_n 0.00553704f $X=9.48 $Y=0.745 $X2=0 $Y2=0
cc_446 C1 N_Y_c_837_n 0.0220461f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_447 N_C1_c_487_n N_Y_c_837_n 0.00164811f $X=9.48 $Y=1.535 $X2=0 $Y2=0
cc_448 C1 N_Y_c_834_n 0.0277326f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_449 N_C1_c_487_n N_Y_c_834_n 0.0065082f $X=9.48 $Y=1.535 $X2=0 $Y2=0
cc_450 C1 N_Y_c_908_n 0.0153756f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_451 N_C1_c_487_n N_Y_c_908_n 7.31333e-19 $X=9.48 $Y=1.535 $X2=0 $Y2=0
cc_452 N_C1_M1008_g N_VGND_c_985_n 0.00302473f $X=7.98 $Y=0.745 $X2=0 $Y2=0
cc_453 N_C1_M1012_g N_VGND_c_985_n 0.00302495f $X=8.53 $Y=0.745 $X2=0 $Y2=0
cc_454 N_C1_M1017_g N_VGND_c_985_n 0.00302473f $X=8.98 $Y=0.745 $X2=0 $Y2=0
cc_455 N_C1_M1022_g N_VGND_c_985_n 0.00302501f $X=9.48 $Y=0.745 $X2=0 $Y2=0
cc_456 N_C1_M1008_g N_VGND_c_986_n 0.00447339f $X=7.98 $Y=0.745 $X2=0 $Y2=0
cc_457 N_C1_M1012_g N_VGND_c_986_n 0.00447412f $X=8.53 $Y=0.745 $X2=0 $Y2=0
cc_458 N_C1_M1017_g N_VGND_c_986_n 0.00443223f $X=8.98 $Y=0.745 $X2=0 $Y2=0
cc_459 N_C1_M1022_g N_VGND_c_986_n 0.00480917f $X=9.48 $Y=0.745 $X2=0 $Y2=0
cc_460 N_C1_M1008_g N_A_1166_65#_c_1206_n 0.0089388f $X=7.98 $Y=0.745 $X2=0
+ $Y2=0
cc_461 N_C1_M1012_g N_A_1166_65#_c_1206_n 0.00995493f $X=8.53 $Y=0.745 $X2=0
+ $Y2=0
cc_462 N_C1_M1008_g N_A_1166_65#_c_1219_n 5.77295e-19 $X=7.98 $Y=0.745 $X2=0
+ $Y2=0
cc_463 N_C1_M1012_g N_A_1166_65#_c_1219_n 0.00604173f $X=8.53 $Y=0.745 $X2=0
+ $Y2=0
cc_464 N_C1_M1017_g N_A_1166_65#_c_1219_n 0.00697855f $X=8.98 $Y=0.745 $X2=0
+ $Y2=0
cc_465 N_C1_M1022_g N_A_1166_65#_c_1219_n 2.75259e-19 $X=9.48 $Y=0.745 $X2=0
+ $Y2=0
cc_466 N_C1_M1017_g N_A_1166_65#_c_1207_n 0.00869988f $X=8.98 $Y=0.745 $X2=0
+ $Y2=0
cc_467 N_C1_M1022_g N_A_1166_65#_c_1207_n 0.0129425f $X=9.48 $Y=0.745 $X2=0
+ $Y2=0
cc_468 N_C1_M1022_g N_A_1166_65#_c_1208_n 0.00375448f $X=9.48 $Y=0.745 $X2=0
+ $Y2=0
cc_469 C1 N_A_1166_65#_c_1208_n 0.0170788f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_470 N_C1_c_487_n N_A_1166_65#_c_1208_n 0.00630056f $X=9.48 $Y=1.535 $X2=0
+ $Y2=0
cc_471 N_C1_M1008_g N_A_1166_65#_c_1209_n 0.00842595f $X=7.98 $Y=0.745 $X2=0
+ $Y2=0
cc_472 N_C1_M1012_g N_A_1166_65#_c_1209_n 2.36317e-19 $X=8.53 $Y=0.745 $X2=0
+ $Y2=0
cc_473 N_C1_M1012_g N_A_1166_65#_c_1210_n 9.44044e-19 $X=8.53 $Y=0.745 $X2=0
+ $Y2=0
cc_474 N_C1_M1017_g N_A_1166_65#_c_1210_n 0.0014148f $X=8.98 $Y=0.745 $X2=0
+ $Y2=0
cc_475 N_A_30_367#_c_561_n N_VPWR_c_638_n 0.0216087f $X=1.04 $Y=1.69 $X2=0 $Y2=0
cc_476 N_A_30_367#_c_563_n N_VPWR_c_639_n 0.0216087f $X=1.9 $Y=1.69 $X2=0 $Y2=0
cc_477 N_A_30_367#_c_574_n N_VPWR_c_645_n 0.0124525f $X=1.995 $Y=1.98 $X2=0
+ $Y2=0
cc_478 N_A_30_367#_c_569_n N_VPWR_c_651_n 0.0178111f $X=0.275 $Y=1.98 $X2=0
+ $Y2=0
cc_479 N_A_30_367#_c_572_n N_VPWR_c_652_n 0.0124525f $X=1.135 $Y=1.98 $X2=0
+ $Y2=0
cc_480 N_A_30_367#_M1005_d N_VPWR_c_637_n 0.00371702f $X=0.15 $Y=1.835 $X2=0
+ $Y2=0
cc_481 N_A_30_367#_M1013_d N_VPWR_c_637_n 0.00536646f $X=0.995 $Y=1.835 $X2=0
+ $Y2=0
cc_482 N_A_30_367#_M1030_d N_VPWR_c_637_n 0.00536646f $X=1.855 $Y=1.835 $X2=0
+ $Y2=0
cc_483 N_A_30_367#_M1019_s N_VPWR_c_637_n 0.00225186f $X=2.715 $Y=1.835 $X2=0
+ $Y2=0
cc_484 N_A_30_367#_M1035_s N_VPWR_c_637_n 0.0021598f $X=3.575 $Y=1.835 $X2=0
+ $Y2=0
cc_485 N_A_30_367#_c_569_n N_VPWR_c_637_n 0.0100304f $X=0.275 $Y=1.98 $X2=0
+ $Y2=0
cc_486 N_A_30_367#_c_572_n N_VPWR_c_637_n 0.00730901f $X=1.135 $Y=1.98 $X2=0
+ $Y2=0
cc_487 N_A_30_367#_c_574_n N_VPWR_c_637_n 0.00730901f $X=1.995 $Y=1.98 $X2=0
+ $Y2=0
cc_488 N_A_30_367#_c_564_n N_A_457_367#_c_777_n 0.0216087f $X=2.76 $Y=1.69 $X2=0
+ $Y2=0
cc_489 N_A_30_367#_M1019_s N_A_457_367#_c_780_n 0.00332344f $X=2.715 $Y=1.835
+ $X2=0 $Y2=0
cc_490 N_A_30_367#_c_576_n N_A_457_367#_c_780_n 0.0126348f $X=2.855 $Y=1.98
+ $X2=0 $Y2=0
cc_491 N_A_30_367#_c_565_n N_A_457_367#_c_782_n 0.0216087f $X=3.62 $Y=1.69 $X2=0
+ $Y2=0
cc_492 N_A_30_367#_M1035_s N_A_457_367#_c_774_n 0.00495471f $X=3.575 $Y=1.835
+ $X2=0 $Y2=0
cc_493 N_A_30_367#_c_578_n N_A_457_367#_c_774_n 0.0189128f $X=3.715 $Y=1.98
+ $X2=0 $Y2=0
cc_494 N_A_30_367#_c_565_n N_Y_c_830_n 0.0130093f $X=3.62 $Y=1.69 $X2=0 $Y2=0
cc_495 N_A_30_367#_c_578_n N_Y_c_830_n 0.010172f $X=3.715 $Y=1.98 $X2=0 $Y2=0
cc_496 N_A_30_367#_c_578_n N_Y_c_836_n 0.0440331f $X=3.715 $Y=1.98 $X2=0 $Y2=0
cc_497 N_A_30_367#_c_578_n N_Y_c_839_n 0.0155096f $X=3.715 $Y=1.98 $X2=0 $Y2=0
cc_498 N_A_30_367#_c_567_n N_A_113_47#_c_1121_n 0.0042147f $X=1.995 $Y=1.69
+ $X2=0 $Y2=0
cc_499 N_A_30_367#_c_565_n N_A_113_47#_c_1133_n 0.00201962f $X=3.62 $Y=1.69
+ $X2=0 $Y2=0
cc_500 N_VPWR_c_637_n N_A_457_367#_M1001_d 0.00223559f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_501 N_VPWR_c_637_n N_A_457_367#_M1024_d 0.00223559f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_637_n N_A_457_367#_M1014_s 0.00223559f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_637_n N_A_457_367#_M1031_s 0.00223559f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_645_n N_A_457_367#_c_775_n 0.01906f $X=6.23 $Y=3.33 $X2=0 $Y2=0
cc_505 N_VPWR_c_637_n N_A_457_367#_c_775_n 0.0124545f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_645_n N_A_457_367#_c_780_n 0.0298674f $X=6.23 $Y=3.33 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_637_n N_A_457_367#_c_780_n 0.0187823f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_645_n N_A_457_367#_c_774_n 0.0637509f $X=6.23 $Y=3.33 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_637_n N_A_457_367#_c_774_n 0.0387091f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_645_n N_A_457_367#_c_792_n 0.0489273f $X=6.23 $Y=3.33 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_637_n N_A_457_367#_c_792_n 0.0312368f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_645_n N_A_457_367#_c_786_n 0.01906f $X=6.23 $Y=3.33 $X2=0 $Y2=0
cc_513 N_VPWR_c_637_n N_A_457_367#_c_786_n 0.0124545f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_514 N_VPWR_c_645_n N_A_457_367#_c_798_n 0.01906f $X=6.23 $Y=3.33 $X2=0 $Y2=0
cc_515 N_VPWR_c_637_n N_A_457_367#_c_798_n 0.0124545f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_637_n N_Y_M1014_d 0.0021598f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_517 N_VPWR_c_637_n N_Y_M1020_d 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_518 N_VPWR_c_637_n N_Y_M1036_d 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_519 N_VPWR_c_637_n N_Y_M1025_s 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_520 N_VPWR_c_637_n N_Y_M1038_s 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_521 N_VPWR_c_637_n N_Y_M1006_d 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_522 N_VPWR_c_637_n N_Y_M1033_d 0.00371702f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_523 N_VPWR_c_647_n N_Y_c_921_n 0.0124525f $X=7.09 $Y=3.33 $X2=0 $Y2=0
cc_524 N_VPWR_c_637_n N_Y_c_921_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_525 N_VPWR_M1032_d N_Y_c_876_n 0.00331217f $X=7.115 $Y=1.835 $X2=0 $Y2=0
cc_526 N_VPWR_c_641_n N_Y_c_876_n 0.0170777f $X=7.255 $Y=2.345 $X2=0 $Y2=0
cc_527 N_VPWR_c_649_n N_Y_c_925_n 0.0124525f $X=7.95 $Y=3.33 $X2=0 $Y2=0
cc_528 N_VPWR_c_637_n N_Y_c_925_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_529 N_VPWR_M1004_s N_Y_c_890_n 0.00331217f $X=7.975 $Y=1.835 $X2=0 $Y2=0
cc_530 N_VPWR_c_642_n N_Y_c_890_n 0.0170777f $X=8.115 $Y=2.345 $X2=0 $Y2=0
cc_531 N_VPWR_c_643_n N_Y_c_929_n 0.0124525f $X=8.81 $Y=3.33 $X2=0 $Y2=0
cc_532 N_VPWR_c_637_n N_Y_c_929_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_533 N_VPWR_M1021_s N_Y_c_899_n 0.00331217f $X=8.835 $Y=1.835 $X2=0 $Y2=0
cc_534 N_VPWR_c_644_n N_Y_c_899_n 0.0170777f $X=8.975 $Y=2.345 $X2=0 $Y2=0
cc_535 N_VPWR_c_653_n N_Y_c_838_n 0.0178111f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_536 N_VPWR_c_637_n N_Y_c_838_n 0.0100304f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_537 N_VPWR_M1003_d N_Y_c_880_n 0.00332882f $X=6.255 $Y=1.835 $X2=0 $Y2=0
cc_538 N_VPWR_c_640_n N_Y_c_880_n 0.0172684f $X=6.395 $Y=2.375 $X2=0 $Y2=0
cc_539 N_VPWR_c_645_n N_Y_c_937_n 0.0124525f $X=6.23 $Y=3.33 $X2=0 $Y2=0
cc_540 N_VPWR_c_637_n N_Y_c_937_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_541 N_A_457_367#_c_774_n N_Y_M1014_d 0.00495471f $X=4.51 $Y=2.99 $X2=0 $Y2=0
cc_542 N_A_457_367#_c_792_n N_Y_M1020_d 0.00332344f $X=5.37 $Y=2.99 $X2=0 $Y2=0
cc_543 N_A_457_367#_c_774_n N_Y_c_836_n 0.0189128f $X=4.51 $Y=2.99 $X2=0 $Y2=0
cc_544 N_A_457_367#_M1014_s N_Y_c_862_n 0.00334509f $X=4.535 $Y=1.835 $X2=0
+ $Y2=0
cc_545 N_A_457_367#_c_789_n N_Y_c_862_n 0.0172684f $X=4.675 $Y=2.375 $X2=0 $Y2=0
cc_546 N_A_457_367#_M1031_s N_Y_c_866_n 0.00334509f $X=5.395 $Y=1.835 $X2=0
+ $Y2=0
cc_547 N_A_457_367#_c_795_n N_Y_c_866_n 0.0172684f $X=5.535 $Y=2.375 $X2=0 $Y2=0
cc_548 N_A_457_367#_c_792_n N_Y_c_946_n 0.0126348f $X=5.37 $Y=2.99 $X2=0 $Y2=0
cc_549 N_Y_c_831_n N_A_113_47#_M1010_s 0.00176891f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_550 N_Y_c_831_n N_A_113_47#_M1029_s 0.00240828f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_551 N_Y_c_831_n N_A_113_47#_c_1138_n 0.0378535f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_552 N_Y_c_832_n N_A_113_47#_c_1138_n 0.00282707f $X=4.295 $Y=1.17 $X2=0 $Y2=0
cc_553 N_Y_c_832_n N_A_113_47#_c_1133_n 0.0141383f $X=4.295 $Y=1.17 $X2=0 $Y2=0
cc_554 N_Y_c_831_n N_A_113_47#_c_1114_n 0.138308f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_555 N_Y_c_831_n N_A_113_47#_c_1154_n 0.014601f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_556 N_Y_c_831_n N_A_1166_65#_M1010_d 0.00288872f $X=8.1 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_557 N_Y_c_831_n N_A_1166_65#_M1011_d 0.00176891f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_558 N_Y_c_831_n N_A_1166_65#_M1034_d 0.00187091f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_559 N_Y_c_833_n N_A_1166_65#_M1012_d 0.00197722f $X=9.1 $Y=1.17 $X2=0 $Y2=0
cc_560 N_Y_c_831_n N_A_1166_65#_c_1205_n 0.0037567f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_561 N_Y_M1008_s N_A_1166_65#_c_1206_n 0.00325942f $X=8.055 $Y=0.325 $X2=0
+ $Y2=0
cc_562 N_Y_c_831_n N_A_1166_65#_c_1206_n 0.00272017f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_563 N_Y_c_961_p N_A_1166_65#_c_1206_n 0.0217182f $X=8.265 $Y=0.68 $X2=0 $Y2=0
cc_564 N_Y_c_833_n N_A_1166_65#_c_1206_n 0.00314622f $X=9.1 $Y=1.17 $X2=0 $Y2=0
cc_565 N_Y_c_833_n N_A_1166_65#_c_1219_n 0.0171395f $X=9.1 $Y=1.17 $X2=0 $Y2=0
cc_566 N_Y_M1017_s N_A_1166_65#_c_1207_n 0.00250873f $X=9.055 $Y=0.325 $X2=0
+ $Y2=0
cc_567 N_Y_c_833_n N_A_1166_65#_c_1207_n 0.00272017f $X=9.1 $Y=1.17 $X2=0 $Y2=0
cc_568 N_Y_c_903_n N_A_1166_65#_c_1207_n 0.0195903f $X=9.265 $Y=0.68 $X2=0 $Y2=0
cc_569 N_Y_c_833_n N_A_1166_65#_c_1208_n 0.0053902f $X=9.1 $Y=1.17 $X2=0 $Y2=0
cc_570 N_Y_c_831_n N_A_1166_65#_c_1209_n 0.0170877f $X=8.1 $Y=1.17 $X2=0 $Y2=0
cc_571 N_VGND_c_986_n N_A_113_47#_M1002_d 0.00408483f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_572 N_VGND_c_986_n N_A_113_47#_M1018_d 0.0028032f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_c_986_n N_A_113_47#_M1000_d 0.0028032f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_574 N_VGND_c_986_n N_A_113_47#_M1023_d 0.00274056f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_575 N_VGND_c_986_n N_A_113_47#_M1007_d 0.00267726f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_576 N_VGND_c_986_n N_A_113_47#_M1026_d 0.00266477f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_577 N_VGND_c_982_n N_A_113_47#_c_1161_n 0.0124525f $X=0.97 $Y=0 $X2=0 $Y2=0
cc_578 N_VGND_c_986_n N_A_113_47#_c_1161_n 0.00730901f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_579 N_VGND_M1016_s N_A_113_47#_c_1115_n 0.00328233f $X=0.995 $Y=0.235 $X2=0
+ $Y2=0
cc_580 N_VGND_c_971_n N_A_113_47#_c_1115_n 0.0167019f $X=1.135 $Y=0.545 $X2=0
+ $Y2=0
cc_581 N_VGND_c_986_n N_A_113_47#_c_1115_n 0.0108944f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_582 N_VGND_c_978_n N_A_113_47#_c_1166_n 0.0124525f $X=1.83 $Y=0 $X2=0 $Y2=0
cc_583 N_VGND_c_986_n N_A_113_47#_c_1166_n 0.00730901f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_584 N_VGND_M1028_s N_A_113_47#_c_1121_n 0.00458879f $X=1.855 $Y=0.235 $X2=0
+ $Y2=0
cc_585 N_VGND_c_972_n N_A_113_47#_c_1121_n 0.0167019f $X=1.995 $Y=0.545 $X2=0
+ $Y2=0
cc_586 N_VGND_c_986_n N_A_113_47#_c_1121_n 0.0108944f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_980_n N_A_113_47#_c_1171_n 0.0124525f $X=2.69 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_986_n N_A_113_47#_c_1171_n 0.00730901f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_M1015_s N_A_113_47#_c_1127_n 0.00328233f $X=2.715 $Y=0.235 $X2=0
+ $Y2=0
cc_590 N_VGND_c_973_n N_A_113_47#_c_1127_n 0.0167019f $X=2.855 $Y=0.545 $X2=0
+ $Y2=0
cc_591 N_VGND_c_986_n N_A_113_47#_c_1127_n 0.0108944f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_592 N_VGND_c_974_n N_A_113_47#_c_1176_n 0.0124525f $X=3.55 $Y=0 $X2=0 $Y2=0
cc_593 N_VGND_c_986_n N_A_113_47#_c_1176_n 0.00730901f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_M1039_s N_A_113_47#_c_1131_n 0.0030939f $X=3.575 $Y=0.235 $X2=0
+ $Y2=0
cc_595 N_VGND_c_974_n N_A_113_47#_c_1131_n 0.00196714f $X=3.55 $Y=0 $X2=0 $Y2=0
cc_596 N_VGND_c_975_n N_A_113_47#_c_1131_n 0.0135609f $X=3.715 $Y=0.45 $X2=0
+ $Y2=0
cc_597 N_VGND_c_986_n N_A_113_47#_c_1131_n 0.00475742f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_c_983_n N_A_113_47#_c_1182_n 0.0124269f $X=4.41 $Y=0 $X2=0 $Y2=0
cc_599 N_VGND_c_986_n N_A_113_47#_c_1182_n 0.00730326f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_600 N_VGND_M1009_s N_A_113_47#_c_1138_n 0.00335318f $X=4.435 $Y=0.235 $X2=0
+ $Y2=0
cc_601 N_VGND_c_976_n N_A_113_47#_c_1138_n 0.0165001f $X=4.575 $Y=0.45 $X2=0
+ $Y2=0
cc_602 N_VGND_c_983_n N_A_113_47#_c_1138_n 0.00191958f $X=4.41 $Y=0 $X2=0 $Y2=0
cc_603 N_VGND_c_984_n N_A_113_47#_c_1138_n 0.00191958f $X=5.27 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_986_n N_A_113_47#_c_1138_n 0.00882814f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_605 N_VGND_M1039_s N_A_113_47#_c_1133_n 3.93454e-19 $X=3.575 $Y=0.235 $X2=0
+ $Y2=0
cc_606 N_VGND_c_975_n N_A_113_47#_c_1133_n 0.00341623f $X=3.715 $Y=0.45 $X2=0
+ $Y2=0
cc_607 N_VGND_c_983_n N_A_113_47#_c_1133_n 0.00193642f $X=4.41 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_c_986_n N_A_113_47#_c_1133_n 0.00422043f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_609 N_VGND_c_984_n N_A_113_47#_c_1193_n 0.0124269f $X=5.27 $Y=0 $X2=0 $Y2=0
cc_610 N_VGND_c_986_n N_A_113_47#_c_1193_n 0.00730326f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_M1037_s N_A_113_47#_c_1114_n 0.00497837f $X=5.295 $Y=0.235 $X2=0
+ $Y2=0
cc_612 N_VGND_c_977_n N_A_113_47#_c_1114_n 0.0213079f $X=5.435 $Y=0.44 $X2=0
+ $Y2=0
cc_613 N_VGND_c_984_n N_A_113_47#_c_1114_n 0.00201785f $X=5.27 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_c_985_n N_A_113_47#_c_1114_n 0.00321199f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_615 N_VGND_c_986_n N_A_113_47#_c_1114_n 0.0134585f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_616 N_VGND_c_977_n N_A_1166_65#_c_1205_n 0.0227137f $X=5.435 $Y=0.44 $X2=0
+ $Y2=0
cc_617 N_VGND_c_985_n N_A_1166_65#_c_1205_n 0.118137f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_618 N_VGND_c_986_n N_A_1166_65#_c_1205_n 0.0654774f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_c_985_n N_A_1166_65#_c_1206_n 0.0423218f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_620 N_VGND_c_986_n N_A_1166_65#_c_1206_n 0.0239549f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_621 N_VGND_c_985_n N_A_1166_65#_c_1207_n 0.0609429f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_622 N_VGND_c_986_n N_A_1166_65#_c_1207_n 0.0340398f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_623 N_VGND_c_985_n N_A_1166_65#_c_1209_n 0.0234634f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_624 N_VGND_c_986_n N_A_1166_65#_c_1209_n 0.0126366f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_625 N_VGND_c_985_n N_A_1166_65#_c_1210_n 0.0234984f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_626 N_VGND_c_986_n N_A_1166_65#_c_1210_n 0.0126823f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_627 N_A_113_47#_c_1114_n N_A_1166_65#_M1010_d 0.00590758f $X=7.265 $Y=0.82
+ $X2=-0.19 $Y2=-0.245
cc_628 N_A_113_47#_c_1114_n N_A_1166_65#_M1011_d 0.00336447f $X=7.265 $Y=0.82
+ $X2=0 $Y2=0
cc_629 N_A_113_47#_M1010_s N_A_1166_65#_c_1205_n 0.00180013f $X=6.265 $Y=0.325
+ $X2=0 $Y2=0
cc_630 N_A_113_47#_M1029_s N_A_1166_65#_c_1205_n 0.00245078f $X=7.125 $Y=0.325
+ $X2=0 $Y2=0
cc_631 N_A_113_47#_c_1114_n N_A_1166_65#_c_1205_n 0.0901911f $X=7.265 $Y=0.82
+ $X2=0 $Y2=0
