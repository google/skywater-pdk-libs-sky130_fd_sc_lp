* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfxtp_2 CLK D VGND VNB VPB VPWR Q
X0 a_679_93# a_110_62# a_1004_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 a_637_119# a_679_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR a_1175_93# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_1004_379# a_240_443# a_1163_379# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_1163_379# a_1175_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_551_119# a_679_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_1004_379# a_110_62# a_1133_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR D a_432_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND D a_432_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR CLK a_110_62# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_240_443# a_110_62# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 Q a_1175_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND CLK a_110_62# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_679_93# a_240_443# a_1004_379# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_432_119# a_240_443# a_551_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_1133_119# a_1175_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_1004_379# a_1175_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 a_551_119# a_240_443# a_637_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_551_119# a_110_62# a_705_443# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_705_443# a_679_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VPWR a_551_119# a_679_93# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 VGND a_1175_93# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 Q a_1175_93# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_240_443# a_110_62# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_1004_379# a_1175_93# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 a_432_119# a_110_62# a_551_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
