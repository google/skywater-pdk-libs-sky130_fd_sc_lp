# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfrbp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfrbp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.24000 BY  3.330000 ;
  SYMMETRY R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.189000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.440000 2.315000 1.460000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.785000 0.265000 18.115000 3.065000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.515000 0.265000 15.845000 3.065000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.567000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.055000 1.550000  1.345000 1.595000 ;
        RECT  1.055000 1.595000 12.385000 1.735000 ;
        RECT  1.055000 1.735000  1.345000 1.780000 ;
        RECT  4.895000 1.550000  5.185000 1.595000 ;
        RECT  4.895000 1.735000  5.185000 1.780000 ;
        RECT 12.095000 1.550000 12.385000 1.595000 ;
        RECT 12.095000 1.735000 12.385000 1.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 13.565000 1.080000 14.275000 1.410000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 18.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 18.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.240000 0.085000 ;
      RECT  0.000000  3.245000 18.240000 3.415000 ;
      RECT  0.100000  2.265000  0.350000 2.895000 ;
      RECT  0.100000  2.895000  1.210000 3.065000 ;
      RECT  0.530000  1.960000  2.985000 2.130000 ;
      RECT  0.530000  2.130000  0.860000 2.715000 ;
      RECT  0.985000  1.110000  1.315000 1.780000 ;
      RECT  1.040000  2.310000  2.185000 2.480000 ;
      RECT  1.040000  2.480000  1.210000 2.895000 ;
      RECT  1.055000  0.085000  1.385000 0.700000 ;
      RECT  1.055000  0.700000  1.315000 0.940000 ;
      RECT  1.425000  2.660000  1.755000 3.245000 ;
      RECT  1.935000  2.480000  2.185000 2.910000 ;
      RECT  2.385000  2.310000  2.635000 2.895000 ;
      RECT  2.385000  2.895000  4.385000 3.065000 ;
      RECT  2.495000  0.580000  2.825000 1.960000 ;
      RECT  2.815000  2.130000  2.985000 2.545000 ;
      RECT  2.815000  2.545000  3.845000 2.715000 ;
      RECT  3.005000  0.580000  3.335000 1.000000 ;
      RECT  3.165000  1.000000  3.335000 1.685000 ;
      RECT  3.165000  1.685000  4.195000 1.855000 ;
      RECT  3.165000  1.855000  3.335000 2.365000 ;
      RECT  3.515000  0.750000  5.395000 0.920000 ;
      RECT  3.515000  0.920000  3.845000 1.460000 ;
      RECT  3.515000  2.035000  3.845000 2.545000 ;
      RECT  4.025000  1.100000  5.870000 1.270000 ;
      RECT  4.025000  1.270000  4.195000 1.685000 ;
      RECT  4.025000  1.855000  4.195000 2.310000 ;
      RECT  4.025000  2.310000  5.850000 2.480000 ;
      RECT  4.055000  2.660000  4.385000 2.895000 ;
      RECT  4.375000  1.455000  4.705000 1.960000 ;
      RECT  4.375000  1.960000  6.380000 2.045000 ;
      RECT  4.375000  2.045000  8.440000 2.130000 ;
      RECT  4.660000  2.660000  4.990000 3.245000 ;
      RECT  4.715000  0.085000  5.045000 0.570000 ;
      RECT  4.925000  1.450000  5.275000 1.780000 ;
      RECT  5.225000  0.265000  6.730000 0.435000 ;
      RECT  5.225000  0.435000  5.395000 0.750000 ;
      RECT  5.520000  2.480000  5.850000 2.725000 ;
      RECT  5.540000  1.270000  5.870000 1.770000 ;
      RECT  6.050000  0.615000  6.380000 1.960000 ;
      RECT  6.050000  2.130000  8.440000 2.215000 ;
      RECT  6.050000  2.215000  6.380000 2.725000 ;
      RECT  6.560000  0.435000  6.730000 1.175000 ;
      RECT  6.560000  1.175000  8.740000 1.345000 ;
      RECT  6.840000  2.395000  7.170000 3.245000 ;
      RECT  6.910000  0.085000  7.240000 0.995000 ;
      RECT  7.815000  0.535000  8.145000 1.175000 ;
      RECT  7.815000  1.345000  8.090000 1.865000 ;
      RECT  8.270000  1.525000  9.250000 1.695000 ;
      RECT  8.270000  1.695000  8.440000 2.045000 ;
      RECT  8.410000  0.675000  8.740000 1.175000 ;
      RECT  8.620000  1.875000  8.870000 2.895000 ;
      RECT  8.620000  2.895000 10.455000 3.065000 ;
      RECT  8.920000  0.265000  9.250000 1.525000 ;
      RECT  9.075000  2.385000 10.105000 2.715000 ;
      RECT  9.080000  1.695000  9.250000 1.875000 ;
      RECT  9.080000  1.875000  9.755000 2.205000 ;
      RECT  9.430000  0.265000  9.760000 1.525000 ;
      RECT  9.430000  1.525000 11.585000 1.695000 ;
      RECT  9.935000  1.695000 10.105000 2.385000 ;
      RECT  9.940000  0.665000 11.315000 0.835000 ;
      RECT  9.940000  0.835000 10.270000 1.345000 ;
      RECT 10.285000  2.655000 10.455000 2.895000 ;
      RECT 10.510000  1.015000 11.935000 1.185000 ;
      RECT 10.510000  1.185000 10.840000 1.345000 ;
      RECT 10.635000  0.085000 10.965000 0.485000 ;
      RECT 10.635000  2.655000 10.885000 3.245000 ;
      RECT 10.905000  1.965000 11.235000 2.425000 ;
      RECT 11.065000  2.425000 11.235000 2.895000 ;
      RECT 11.065000  2.895000 12.635000 3.065000 ;
      RECT 11.145000  0.265000 14.000000 0.435000 ;
      RECT 11.145000  0.435000 11.315000 0.665000 ;
      RECT 11.215000  1.365000 11.585000 1.525000 ;
      RECT 11.415000  1.695000 11.585000 2.545000 ;
      RECT 11.415000  2.545000 12.285000 2.715000 ;
      RECT 11.765000  0.615000 13.275000 0.865000 ;
      RECT 11.765000  0.865000 11.935000 1.015000 ;
      RECT 11.765000  1.185000 11.935000 2.365000 ;
      RECT 12.115000  1.960000 13.370000 2.130000 ;
      RECT 12.115000  2.130000 12.285000 2.545000 ;
      RECT 12.125000  1.110000 12.455000 1.780000 ;
      RECT 12.465000  2.310000 13.495000 2.480000 ;
      RECT 12.465000  2.480000 12.635000 2.895000 ;
      RECT 12.815000  2.660000 12.985000 3.245000 ;
      RECT 13.040000  1.590000 14.985000 1.760000 ;
      RECT 13.040000  1.760000 13.370000 1.960000 ;
      RECT 13.165000  2.480000 13.495000 2.990000 ;
      RECT 13.670000  0.435000 14.000000 0.730000 ;
      RECT 13.670000  0.730000 15.335000 0.900000 ;
      RECT 13.700000  1.940000 15.335000 2.110000 ;
      RECT 13.700000  2.110000 14.030000 2.495000 ;
      RECT 14.490000  0.085000 14.820000 0.550000 ;
      RECT 14.715000  2.290000 15.045000 3.245000 ;
      RECT 14.725000  1.345000 14.985000 1.590000 ;
      RECT 15.165000  0.900000 15.335000 1.940000 ;
      RECT 16.090000  0.665000 16.420000 1.305000 ;
      RECT 16.090000  1.305000 17.605000 1.635000 ;
      RECT 16.090000  1.635000 16.420000 2.495000 ;
      RECT 16.995000  0.085000 17.325000 1.125000 ;
      RECT 16.995000  1.815000 17.325000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.580000  1.285000 1.750000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.580000  5.125000 1.750000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  1.580000 12.325000 1.750000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.245000 18.085000 3.415000 ;
  END
END sky130_fd_sc_lp__dfrbp_lp
END LIBRARY
