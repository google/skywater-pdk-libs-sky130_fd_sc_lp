* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
X0 a_185_23# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_27_133# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_516_125# a_558_99# a_588_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR B_N a_558_99# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_696_125# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR C a_185_23# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_27_133# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_185_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_185_23# a_27_133# a_516_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_27_133# a_185_23# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VGND a_185_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_588_125# C a_696_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 X a_185_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VGND B_N a_558_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 X a_185_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_185_23# a_558_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
