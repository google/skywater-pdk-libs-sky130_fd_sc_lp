* File: sky130_fd_sc_lp__o32ai_1.pex.spice
* Created: Wed Sep  2 10:26:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32AI_1%B1 1 3 6 8 9 10 18 20
r34 15 18 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.5 $Y=1.46 $X2=0.72
+ $Y2=1.46
r35 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.5
+ $Y=1.46 $X2=0.5 $Y2=1.46
r36 10 16 4.71531 $w=5.18e-07 $l=2.05e-07 $layer=LI1_cond $X=0.345 $Y=1.665
+ $X2=0.345 $Y2=1.46
r37 9 16 3.79525 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=0.345 $Y=1.295
+ $X2=0.345 $Y2=1.46
r38 9 20 2.30015 $w=5.18e-07 $l=1e-07 $layer=LI1_cond $X=0.345 $Y=1.295
+ $X2=0.345 $Y2=1.195
r39 8 20 6.33462 $w=5.2e-07 $l=2.7e-07 $layer=LI1_cond $X=0.345 $Y=0.925
+ $X2=0.345 $Y2=1.195
r40 4 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.625
+ $X2=0.72 $Y2=1.46
r41 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.72 $Y=1.625 $X2=0.72
+ $Y2=2.465
r42 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.295
+ $X2=0.72 $Y2=1.46
r43 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.72 $Y=1.295 $X2=0.72
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_1%B2 3 7 9 12 13
c36 3 0 1.81973e-19 $X=1.08 $Y=2.465
r37 12 15 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.51
+ $X2=1.185 $Y2=1.675
r38 12 14 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.51
+ $X2=1.185 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.51 $X2=1.2 $Y2=1.51
r40 9 13 5.95429 $w=2.98e-07 $l=1.55e-07 $layer=LI1_cond $X=1.265 $Y=1.665
+ $X2=1.265 $Y2=1.51
r41 7 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.2 $Y=0.765 $X2=1.2
+ $Y2=1.345
r42 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.08 $Y=2.465
+ $X2=1.08 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_1%A3 1 3 6 8 9 17
c35 8 0 4.48966e-19 $X=1.68 $Y=1.295
r36 15 17 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.76 $Y=1.46
+ $X2=1.92 $Y2=1.46
r37 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.76
+ $Y=1.46 $X2=1.76 $Y2=1.46
r38 12 15 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.65 $Y=1.46
+ $X2=1.76 $Y2=1.46
r39 9 16 8.43753 $w=2.78e-07 $l=2.05e-07 $layer=LI1_cond $X=1.725 $Y=1.665
+ $X2=1.725 $Y2=1.46
r40 8 16 6.79118 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=1.295
+ $X2=1.725 $Y2=1.46
r41 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.625
+ $X2=1.92 $Y2=1.46
r42 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.92 $Y=1.625 $X2=1.92
+ $Y2=2.465
r43 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=1.295
+ $X2=1.65 $Y2=1.46
r44 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.65 $Y=1.295 $X2=1.65
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_1%A2 3 7 8 10 17 19
c31 19 0 3.80786e-19 $X=2.37 $Y=1.295
c32 3 0 8.89057e-20 $X=2.37 $Y=2.465
r33 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.46
+ $X2=2.37 $Y2=1.295
r34 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=1.46 $X2=2.37 $Y2=1.46
r35 10 18 5.20873 $w=6.18e-07 $l=2.7e-07 $layer=LI1_cond $X=2.64 $Y=1.52
+ $X2=2.37 $Y2=1.52
r36 8 18 4.05123 $w=6.18e-07 $l=2.1e-07 $layer=LI1_cond $X=2.16 $Y=1.52 $X2=2.37
+ $Y2=1.52
r37 7 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.42 $Y=0.765
+ $X2=2.42 $Y2=1.295
r38 1 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.625
+ $X2=2.37 $Y2=1.46
r39 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.37 $Y=1.625 $X2=2.37
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_1%A1 3 7 8 9 13 15
c24 15 0 1.41268e-19 $X=2.95 $Y=1.295
c25 8 0 6.143e-20 $X=3.12 $Y=1.295
r26 13 16 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.46
+ $X2=2.95 $Y2=1.625
r27 13 15 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.46
+ $X2=2.95 $Y2=1.295
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.46 $X2=2.99 $Y2=1.46
r29 9 14 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.46
r30 8 14 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.46
r31 7 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.85 $Y=0.765
+ $X2=2.85 $Y2=1.295
r32 3 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.82 $Y=2.465
+ $X2=2.82 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_1%VPWR 1 2 9 13 15 20 21 22 28 37
r31 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 34 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r33 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 30 33 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 28 36 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.87 $Y=3.33
+ $X2=3.115 $Y2=3.33
r37 28 33 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.87 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 26 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 22 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 22 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 20 25 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.34 $Y=3.33 $X2=0.24
+ $Y2=3.33
r43 20 21 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=0.34 $Y=3.33
+ $X2=0.472 $Y2=3.33
r44 19 30 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 19 21 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.472 $Y2=3.33
r46 15 18 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=3.035 $Y=2.005
+ $X2=3.035 $Y2=2.95
r47 13 36 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.035 $Y=3.245
+ $X2=3.115 $Y2=3.33
r48 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.035 $Y=3.245
+ $X2=3.035 $Y2=2.95
r49 9 12 37.6175 $w=2.63e-07 $l=8.65e-07 $layer=LI1_cond $X=0.472 $Y=2.085
+ $X2=0.472 $Y2=2.95
r50 7 21 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.472 $Y=3.245
+ $X2=0.472 $Y2=3.33
r51 7 12 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.472 $Y=3.245
+ $X2=0.472 $Y2=2.95
r52 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=1.835 $X2=3.035 $Y2=2.95
r53 2 15 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=1.835 $X2=3.035 $Y2=2.005
r54 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.38
+ $Y=1.835 $X2=0.505 $Y2=2.95
r55 1 9 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.38
+ $Y=1.835 $X2=0.505 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_1%Y 1 2 8 12 15 16 17 18 29 30
r30 29 30 12.4766 $w=1.093e-06 $l=8.5e-08 $layer=LI1_cond $X=1.322 $Y=2.005
+ $X2=1.322 $Y2=1.92
r31 18 41 1.94977 $w=1.093e-06 $l=1.75e-07 $layer=LI1_cond $X=1.322 $Y=2.775
+ $X2=1.322 $Y2=2.95
r32 17 18 4.12237 $w=1.093e-06 $l=3.7e-07 $layer=LI1_cond $X=1.322 $Y=2.405
+ $X2=1.322 $Y2=2.775
r33 16 17 4.12237 $w=1.093e-06 $l=3.7e-07 $layer=LI1_cond $X=1.322 $Y=2.035
+ $X2=1.322 $Y2=2.405
r34 16 29 0.334247 $w=1.093e-06 $l=3e-08 $layer=LI1_cond $X=1.322 $Y=2.035
+ $X2=1.322 $Y2=2.005
r35 15 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.86 $Y=1.175
+ $X2=0.86 $Y2=1.92
r36 12 14 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.935 $Y=0.72
+ $X2=0.935 $Y2=0.765
r37 8 15 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=0.937 $Y=1.013
+ $X2=0.937 $Y2=1.175
r38 8 14 8.79403 $w=3.23e-07 $l=2.48e-07 $layer=LI1_cond $X=0.937 $Y=1.013
+ $X2=0.937 $Y2=0.765
r39 2 41 200 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=3 $X=1.155
+ $Y=1.835 $X2=1.295 $Y2=2.95
r40 2 29 200 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=3 $X=1.155
+ $Y=1.835 $X2=1.295 $Y2=2.005
r41 1 12 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=0.795
+ $Y=0.345 $X2=0.935 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_1%A_76_69# 1 2 3 10 15 16 17 20 22
c34 20 0 2.82536e-19 $X=2.635 $Y=0.49
r35 22 25 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=0.47 $Y=0.34
+ $X2=0.47 $Y2=0.49
r36 18 20 22.1818 $w=1.88e-07 $l=3.8e-07 $layer=LI1_cond $X=2.635 $Y=0.87
+ $X2=2.635 $Y2=0.49
r37 16 18 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.54 $Y=0.955
+ $X2=2.635 $Y2=0.87
r38 16 17 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.54 $Y=0.955
+ $X2=1.53 $Y2=0.955
r39 13 17 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.4 $Y=0.87
+ $X2=1.53 $Y2=0.955
r40 13 15 16.8434 $w=2.58e-07 $l=3.8e-07 $layer=LI1_cond $X=1.4 $Y=0.87 $X2=1.4
+ $Y2=0.49
r41 12 15 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=1.4 $Y=0.425 $X2=1.4
+ $Y2=0.49
r42 11 22 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.6 $Y=0.34 $X2=0.47
+ $Y2=0.34
r43 10 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.27 $Y=0.34
+ $X2=1.4 $Y2=0.425
r44 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.27 $Y=0.34 $X2=0.6
+ $Y2=0.34
r45 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.495
+ $Y=0.345 $X2=2.635 $Y2=0.49
r46 2 15 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.275
+ $Y=0.345 $X2=1.435 $Y2=0.49
r47 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.38
+ $Y=0.345 $X2=0.505 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_1%VGND 1 2 7 9 11 13 21 28 35
r36 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r37 28 31 10.2649 $w=6.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.035 $Y=0
+ $X2=2.035 $Y2=0.575
r38 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r40 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r41 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 22 28 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.035
+ $Y2=0
r43 22 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.64
+ $Y2=0
r44 21 34 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=3.13
+ $Y2=0
r45 21 24 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=2.64
+ $Y2=0
r46 15 19 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r47 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 13 28 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.7 $Y=0 $X2=2.035
+ $Y2=0
r49 13 19 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.68
+ $Y2=0
r50 11 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r51 11 16 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r52 11 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 7 34 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.13 $Y2=0
r54 7 9 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.065 $Y2=0.49
r55 2 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.925
+ $Y=0.345 $X2=3.065 $Y2=0.49
r56 1 31 91 $w=1.7e-07 $l=5.83781e-07 $layer=licon1_NDIFF $count=2 $X=1.725
+ $Y=0.345 $X2=2.205 $Y2=0.575
.ends

