# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrtn_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465000 0.840000 0.835000 1.790000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.905000 0.255000 6.115000 2.145000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945000 0.375000 5.185000 0.685000 ;
        RECT 4.945000 0.685000 5.520000 0.855000 ;
        RECT 5.260000 0.855000 5.520000 1.515000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 0.840000 1.295000 1.790000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  0.395000 0.530000 0.670000 ;
      RECT 0.115000  0.670000 0.285000 1.960000 ;
      RECT 0.115000  1.960000 1.145000 2.130000 ;
      RECT 0.115000  2.130000 0.410000 2.970000 ;
      RECT 0.580000  2.300000 0.805000 3.245000 ;
      RECT 0.700000  0.085000 0.940000 0.670000 ;
      RECT 0.975000  2.130000 1.145000 2.810000 ;
      RECT 0.975000  2.810000 1.985000 2.980000 ;
      RECT 1.110000  0.340000 1.635000 0.670000 ;
      RECT 1.325000  2.300000 1.635000 2.630000 ;
      RECT 1.465000  0.670000 1.635000 1.155000 ;
      RECT 1.465000  1.155000 1.755000 1.825000 ;
      RECT 1.465000  1.825000 1.635000 2.300000 ;
      RECT 1.815000  2.425000 2.910000 2.595000 ;
      RECT 1.815000  2.595000 1.985000 2.810000 ;
      RECT 1.820000  1.995000 2.150000 2.255000 ;
      RECT 1.885000  0.670000 2.145000 0.995000 ;
      RECT 1.925000  0.995000 2.145000 1.125000 ;
      RECT 1.925000  1.125000 3.380000 1.295000 ;
      RECT 1.925000  1.295000 2.150000 1.995000 ;
      RECT 2.315000  0.085000 2.645000 0.955000 ;
      RECT 2.400000  2.765000 2.730000 3.245000 ;
      RECT 2.580000  1.515000 2.910000 2.425000 ;
      RECT 2.815000  0.255000 3.670000 0.500000 ;
      RECT 2.815000  0.500000 2.985000 1.125000 ;
      RECT 3.120000  1.295000 3.380000 2.205000 ;
      RECT 3.175000  0.670000 3.720000 0.955000 ;
      RECT 3.265000  2.375000 3.720000 3.015000 ;
      RECT 3.550000  0.955000 3.720000 1.365000 ;
      RECT 3.550000  1.365000 4.750000 1.550000 ;
      RECT 3.550000  1.550000 3.720000 2.375000 ;
      RECT 4.005000  0.085000 4.335000 1.000000 ;
      RECT 4.025000  1.720000 5.540000 1.890000 ;
      RECT 4.025000  1.890000 4.355000 2.190000 ;
      RECT 4.150000  2.410000 4.855000 3.245000 ;
      RECT 4.525000  0.255000 4.775000 1.025000 ;
      RECT 4.525000  1.025000 5.090000 1.195000 ;
      RECT 4.525000  2.060000 4.855000 2.410000 ;
      RECT 4.920000  1.195000 5.090000 1.720000 ;
      RECT 5.025000  1.890000 5.540000 2.315000 ;
      RECT 5.025000  2.315000 6.615000 2.485000 ;
      RECT 5.025000  2.485000 5.235000 3.075000 ;
      RECT 5.355000  0.085000 5.685000 0.515000 ;
      RECT 5.405000  2.655000 5.735000 3.245000 ;
      RECT 6.285000  0.085000 6.615000 1.095000 ;
      RECT 6.285000  2.655000 6.615000 3.245000 ;
      RECT 6.345000  1.295000 6.615000 2.315000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrtn_2
END LIBRARY
