# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a21boi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a21boi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 1.425000 3.315000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.250000 1.425000 2.595000 1.595000 ;
        RECT 2.425000 1.595000 2.595000 1.925000 ;
        RECT 2.425000 1.925000 3.745000 2.120000 ;
        RECT 3.515000 1.355000 4.060000 1.645000 ;
        RECT 3.515000 1.645000 3.745000 1.925000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.320000 0.470000 2.490000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.890400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 0.285000 1.805000 1.075000 ;
        RECT 1.545000 1.075000 3.325000 1.245000 ;
        RECT 1.545000 1.245000 1.795000 1.820000 ;
        RECT 1.545000 1.820000 1.875000 2.730000 ;
        RECT 2.995000 0.605000 3.325000 1.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.140000  2.660000 0.470000 3.245000 ;
      RECT 0.640000  0.370000 0.920000 1.340000 ;
      RECT 0.640000  1.340000 1.165000 1.605000 ;
      RECT 0.640000  1.605000 0.900000 2.875000 ;
      RECT 1.115000  0.085000 1.375000 1.170000 ;
      RECT 1.115000  1.830000 1.375000 2.905000 ;
      RECT 1.115000  2.905000 2.315000 3.075000 ;
      RECT 1.975000  0.085000 2.305000 0.905000 ;
      RECT 2.045000  1.830000 2.245000 2.290000 ;
      RECT 2.045000  2.290000 4.185000 2.460000 ;
      RECT 2.045000  2.460000 2.315000 2.905000 ;
      RECT 2.485000  0.265000 3.720000 0.435000 ;
      RECT 2.485000  0.435000 2.815000 0.905000 ;
      RECT 2.485000  2.640000 2.815000 3.245000 ;
      RECT 2.985000  2.460000 3.255000 2.970000 ;
      RECT 3.425000  2.630000 3.755000 3.245000 ;
      RECT 3.495000  0.435000 3.720000 1.185000 ;
      RECT 3.890000  0.085000 4.185000 1.185000 ;
      RECT 3.915000  1.815000 4.185000 2.290000 ;
      RECT 3.925000  2.460000 4.185000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__a21boi_2
END LIBRARY
