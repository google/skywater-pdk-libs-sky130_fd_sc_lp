* File: sky130_fd_sc_lp__clkinv_4.pex.spice
* Created: Fri Aug 28 10:18:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKINV_4%A 3 7 11 15 19 23 27 31 35 39 41 42 43 44
+ 45 69 70
r86 69 71 12.0818 $w=3.79e-07 $l=9.5e-08 $layer=POLY_cond $X=2.7 $Y=1.485
+ $X2=2.795 $Y2=1.485
r87 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7
+ $Y=1.46 $X2=2.7 $Y2=1.46
r88 67 69 42.6042 $w=3.79e-07 $l=3.35e-07 $layer=POLY_cond $X=2.365 $Y=1.485
+ $X2=2.7 $Y2=1.485
r89 65 67 0.635884 $w=3.79e-07 $l=5e-09 $layer=POLY_cond $X=2.36 $Y=1.485
+ $X2=2.365 $Y2=1.485
r90 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.36
+ $Y=1.46 $X2=2.36 $Y2=1.46
r91 63 65 54.0501 $w=3.79e-07 $l=4.25e-07 $layer=POLY_cond $X=1.935 $Y=1.485
+ $X2=2.36 $Y2=1.485
r92 61 63 32.4301 $w=3.79e-07 $l=2.55e-07 $layer=POLY_cond $X=1.68 $Y=1.485
+ $X2=1.935 $Y2=1.485
r93 59 61 22.2559 $w=3.79e-07 $l=1.75e-07 $layer=POLY_cond $X=1.505 $Y=1.485
+ $X2=1.68 $Y2=1.485
r94 57 59 20.9842 $w=3.79e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.485
+ $X2=1.505 $Y2=1.485
r95 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.34
+ $Y=1.46 $X2=1.34 $Y2=1.46
r96 55 57 33.7018 $w=3.79e-07 $l=2.65e-07 $layer=POLY_cond $X=1.075 $Y=1.485
+ $X2=1.34 $Y2=1.485
r97 53 55 9.53826 $w=3.79e-07 $l=7.5e-08 $layer=POLY_cond $X=1 $Y=1.485
+ $X2=1.075 $Y2=1.485
r98 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.46
+ $X2=1 $Y2=1.46
r99 51 53 45.1478 $w=3.79e-07 $l=3.55e-07 $layer=POLY_cond $X=0.645 $Y=1.485
+ $X2=1 $Y2=1.485
r100 45 70 2.06408 $w=3.33e-07 $l=6e-08 $layer=LI1_cond $X=2.64 $Y=1.377 $X2=2.7
+ $Y2=1.377
r101 45 66 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=2.64 $Y=1.377
+ $X2=2.36 $Y2=1.377
r102 44 66 6.88026 $w=3.33e-07 $l=2e-07 $layer=LI1_cond $X=2.16 $Y=1.377
+ $X2=2.36 $Y2=1.377
r103 43 44 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.377
+ $X2=2.16 $Y2=1.377
r104 43 58 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=1.68 $Y=1.377
+ $X2=1.34 $Y2=1.377
r105 43 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.46 $X2=1.68 $Y2=1.46
r106 42 58 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.377
+ $X2=1.34 $Y2=1.377
r107 42 54 6.88026 $w=3.33e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=1.377 $X2=1
+ $Y2=1.377
r108 41 54 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=0.72 $Y=1.377 $X2=1
+ $Y2=1.377
r109 37 71 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.795 $Y=1.675
+ $X2=2.795 $Y2=1.485
r110 37 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.795 $Y=1.675
+ $X2=2.795 $Y2=2.465
r111 33 67 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.365 $Y=1.675
+ $X2=2.365 $Y2=1.485
r112 33 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.365 $Y=1.675
+ $X2=2.365 $Y2=2.465
r113 29 67 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.365 $Y=1.295
+ $X2=2.365 $Y2=1.485
r114 29 31 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=2.365 $Y=1.295
+ $X2=2.365 $Y2=0.56
r115 25 63 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.935 $Y=1.675
+ $X2=1.935 $Y2=1.485
r116 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.935 $Y=1.675
+ $X2=1.935 $Y2=2.465
r117 21 63 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.935 $Y=1.295
+ $X2=1.935 $Y2=1.485
r118 21 23 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.935 $Y=1.295
+ $X2=1.935 $Y2=0.56
r119 17 59 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.505 $Y=1.675
+ $X2=1.505 $Y2=1.485
r120 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.505 $Y=1.675
+ $X2=1.505 $Y2=2.465
r121 13 59 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.505 $Y=1.295
+ $X2=1.505 $Y2=1.485
r122 13 15 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.505 $Y=1.295
+ $X2=1.505 $Y2=0.56
r123 9 55 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.075 $Y=1.675
+ $X2=1.075 $Y2=1.485
r124 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.075 $Y=1.675
+ $X2=1.075 $Y2=2.465
r125 5 55 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.075 $Y=1.295
+ $X2=1.075 $Y2=1.485
r126 5 7 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.075 $Y=1.295
+ $X2=1.075 $Y2=0.56
r127 1 51 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.645 $Y=1.675
+ $X2=0.645 $Y2=1.485
r128 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.645 $Y=1.675
+ $X2=0.645 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_4%VPWR 1 2 3 4 15 19 23 29 33 35 39 40 41 46
+ 51 57 60 64
r53 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 55 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 55 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 52 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=3.33 $X2=2.15
+ $Y2=3.33
r60 52 54 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 51 63 3.93273 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=3.33 $X2=3.12
+ $Y2=3.33
r62 51 54 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 47 57 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.42 $Y=3.33 $X2=1.29
+ $Y2=3.33
r64 47 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.42 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 46 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.02 $Y=3.33 $X2=2.15
+ $Y2=3.33
r66 46 49 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.02 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 45 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 41 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 41 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r71 41 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 39 44 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=0.3 $Y=3.33 $X2=0.24
+ $Y2=3.33
r73 39 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.3 $Y=3.33 $X2=0.43
+ $Y2=3.33
r74 35 38 31.4097 $w=2.53e-07 $l=6.95e-07 $layer=LI1_cond $X=3.007 $Y=2.22
+ $X2=3.007 $Y2=2.915
r75 33 63 3.2445 $w=2.55e-07 $l=1.49579e-07 $layer=LI1_cond $X=3.007 $Y=3.245
+ $X2=3.12 $Y2=3.33
r76 33 38 14.914 $w=2.53e-07 $l=3.3e-07 $layer=LI1_cond $X=3.007 $Y=3.245
+ $X2=3.007 $Y2=2.915
r77 29 32 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=2.15 $Y=2.22
+ $X2=2.15 $Y2=2.915
r78 27 60 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r79 27 32 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.915
r80 23 26 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=1.29 $Y=2.22
+ $X2=1.29 $Y2=2.915
r81 21 57 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.29 $Y=3.245
+ $X2=1.29 $Y2=3.33
r82 21 26 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=1.29 $Y=3.245
+ $X2=1.29 $Y2=2.915
r83 20 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.43
+ $Y2=3.33
r84 19 57 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.16 $Y=3.33 $X2=1.29
+ $Y2=3.33
r85 19 20 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.16 $Y=3.33 $X2=0.56
+ $Y2=3.33
r86 15 18 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=0.43 $Y=2.22
+ $X2=0.43 $Y2=2.915
r87 13 40 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.43 $Y=3.245
+ $X2=0.43 $Y2=3.33
r88 13 18 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=0.43 $Y=3.245
+ $X2=0.43 $Y2=2.915
r89 4 38 400 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.835 $X2=3.01 $Y2=2.915
r90 4 35 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.835 $X2=3.01 $Y2=2.22
r91 3 32 400 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.15 $Y2=2.915
r92 3 29 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.15 $Y2=2.22
r93 2 26 400 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=1.835 $X2=1.29 $Y2=2.915
r94 2 23 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=1.835 $X2=1.29 $Y2=2.22
r95 1 18 400 $w=1.7e-07 $l=1.14315e-06 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.835 $X2=0.43 $Y2=2.915
r96 1 15 400 $w=1.7e-07 $l=4.45281e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.835 $X2=0.43 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_4%Y 1 2 3 4 5 17 18 19 20 21 24 28 32 34 38
+ 42 46 50 54 55 56 58 60 61 62 63 70 71 76
r98 71 76 2.99754 $w=1.83e-07 $l=5e-08 $layer=LI1_cond $X=3.127 $Y=1.715
+ $X2=3.127 $Y2=1.665
r99 63 71 3.28106 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.127 $Y=1.8
+ $X2=3.127 $Y2=1.715
r100 63 76 1.07912 $w=1.83e-07 $l=1.8e-08 $layer=LI1_cond $X=3.127 $Y=1.647
+ $X2=3.127 $Y2=1.665
r101 62 63 21.1027 $w=1.83e-07 $l=3.52e-07 $layer=LI1_cond $X=3.127 $Y=1.295
+ $X2=3.127 $Y2=1.647
r102 62 70 15.2875 $w=1.83e-07 $l=2.55e-07 $layer=LI1_cond $X=3.127 $Y=1.295
+ $X2=3.127 $Y2=1.04
r103 61 70 3.55727 $w=1.85e-07 $l=1e-07 $layer=LI1_cond $X=3.127 $Y=0.94
+ $X2=3.127 $Y2=1.04
r104 59 63 17.9392 $w=2.03e-07 $l=3.25e-07 $layer=LI1_cond $X=2.71 $Y=1.8
+ $X2=3.035 $Y2=1.8
r105 59 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=1.8 $X2=2.58
+ $Y2=1.8
r106 57 61 24.9971 $w=3.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.275 $Y=0.94
+ $X2=3.035 $Y2=0.94
r107 57 58 6.29182 $w=2e-07 $l=1.28e-07 $layer=LI1_cond $X=2.275 $Y=0.94
+ $X2=2.147 $Y2=0.94
r108 50 52 39.0058 $w=2.58e-07 $l=8.8e-07 $layer=LI1_cond $X=2.58 $Y=2 $X2=2.58
+ $Y2=2.88
r109 48 60 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=1.885
+ $X2=2.58 $Y2=1.8
r110 48 50 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=2.58 $Y=1.885
+ $X2=2.58 $Y2=2
r111 44 58 0.484182 $w=2.55e-07 $l=1e-07 $layer=LI1_cond $X=2.147 $Y=0.84
+ $X2=2.147 $Y2=0.94
r112 44 46 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=2.147 $Y=0.84
+ $X2=2.147 $Y2=0.56
r113 43 56 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.85 $Y=1.8
+ $X2=1.722 $Y2=1.8
r114 42 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.45 $Y=1.8 $X2=2.58
+ $Y2=1.8
r115 42 43 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.45 $Y=1.8 $X2=1.85
+ $Y2=1.8
r116 38 40 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=1.722 $Y=2
+ $X2=1.722 $Y2=2.88
r117 36 56 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.722 $Y=1.885
+ $X2=1.722 $Y2=1.8
r118 36 38 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=1.722 $Y=1.885
+ $X2=1.722 $Y2=2
r119 35 55 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.42 $Y=0.94 $X2=1.29
+ $Y2=0.94
r120 34 58 6.29182 $w=2e-07 $l=1.27e-07 $layer=LI1_cond $X=2.02 $Y=0.94
+ $X2=2.147 $Y2=0.94
r121 34 35 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=2.02 $Y=0.94 $X2=1.42
+ $Y2=0.94
r122 30 55 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=1.29 $Y=0.84 $X2=1.29
+ $Y2=0.94
r123 30 32 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=1.29 $Y=0.84
+ $X2=1.29 $Y2=0.56
r124 29 54 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.99 $Y=1.8
+ $X2=0.862 $Y2=1.8
r125 28 56 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.595 $Y=1.8
+ $X2=1.722 $Y2=1.8
r126 28 29 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.595 $Y=1.8
+ $X2=0.99 $Y2=1.8
r127 24 26 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=0.862 $Y=2
+ $X2=0.862 $Y2=2.88
r128 22 54 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.862 $Y=1.885
+ $X2=0.862 $Y2=1.8
r129 22 24 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=0.862 $Y=1.885
+ $X2=0.862 $Y2=2
r130 20 54 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.735 $Y=1.8
+ $X2=0.862 $Y2=1.8
r131 20 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.735 $Y=1.8
+ $X2=0.4 $Y2=1.8
r132 18 55 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.16 $Y=0.94 $X2=1.29
+ $Y2=0.94
r133 18 19 42.1455 $w=1.98e-07 $l=7.6e-07 $layer=LI1_cond $X=1.16 $Y=0.94
+ $X2=0.4 $Y2=0.94
r134 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.315 $Y=1.715
+ $X2=0.4 $Y2=1.8
r135 16 19 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.315 $Y=1.04
+ $X2=0.4 $Y2=0.94
r136 16 17 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.315 $Y=1.04
+ $X2=0.315 $Y2=1.715
r137 5 52 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.835 $X2=2.58 $Y2=2.88
r138 5 50 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.835 $X2=2.58 $Y2=2
r139 4 40 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.835 $X2=1.72 $Y2=2.88
r140 4 38 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.835 $X2=1.72 $Y2=2
r141 3 26 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.835 $X2=0.86 $Y2=2.88
r142 3 24 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.835 $X2=0.86 $Y2=2
r143 2 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.01
+ $Y=0.35 $X2=2.15 $Y2=0.56
r144 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.15
+ $Y=0.35 $X2=1.29 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_4%VGND 1 2 3 14 18 22 24 26 31 38 39 42 45 48
r34 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 39 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r37 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r38 36 48 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.595
+ $Y2=0
r39 36 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=3.12
+ $Y2=0
r40 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 32 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.72
+ $Y2=0
r43 32 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.16
+ $Y2=0
r44 31 48 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.595
+ $Y2=0
r45 31 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.16
+ $Y2=0
r46 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r47 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r48 27 42 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.842
+ $Y2=0
r49 27 29 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r50 26 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.59 $Y=0 $X2=1.72
+ $Y2=0
r51 26 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.59 $Y=0 $X2=1.2
+ $Y2=0
r52 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r53 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 24 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 20 48 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0
r56 20 22 16.1342 $w=2.98e-07 $l=4.2e-07 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0.505
r57 16 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0
r58 16 18 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0.505
r59 12 42 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0
r60 12 14 16.4077 $w=2.93e-07 $l=4.2e-07 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0.505
r61 3 22 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.35 $X2=2.58 $Y2=0.505
r62 2 18 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.58
+ $Y=0.35 $X2=1.72 $Y2=0.505
r63 1 14 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.735
+ $Y=0.35 $X2=0.86 $Y2=0.505
.ends

