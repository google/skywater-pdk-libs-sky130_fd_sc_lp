* NGSPICE file created from sky130_fd_sc_lp__tapvgnd_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__tapvgnd_1 VGND VPB VPWR
.ends

