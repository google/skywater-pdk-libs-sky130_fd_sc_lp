* File: sky130_fd_sc_lp__nor3_2.pxi.spice
* Created: Fri Aug 28 10:55:33 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3_2%A N_A_M1000_g N_A_c_59_n N_A_M1004_g N_A_c_60_n
+ N_A_M1006_g N_A_M1009_g A A N_A_c_62_n N_A_c_63_n PM_SKY130_FD_SC_LP__NOR3_2%A
x_PM_SKY130_FD_SC_LP__NOR3_2%B N_B_M1010_g N_B_M1002_g N_B_c_106_n N_B_M1011_g
+ N_B_M1005_g N_B_c_108_n N_B_c_109_n B B N_B_c_111_n N_B_c_112_n N_B_c_113_n B
+ PM_SKY130_FD_SC_LP__NOR3_2%B
x_PM_SKY130_FD_SC_LP__NOR3_2%C N_C_c_183_n N_C_M1003_g N_C_c_187_n N_C_M1001_g
+ N_C_c_184_n N_C_M1007_g N_C_c_188_n N_C_M1008_g C C N_C_c_186_n
+ PM_SKY130_FD_SC_LP__NOR3_2%C
x_PM_SKY130_FD_SC_LP__NOR3_2%A_36_367# N_A_36_367#_M1000_s N_A_36_367#_M1009_s
+ N_A_36_367#_M1005_d N_A_36_367#_c_234_n N_A_36_367#_c_235_n
+ N_A_36_367#_c_236_n N_A_36_367#_c_244_n N_A_36_367#_c_246_n
+ N_A_36_367#_c_262_p N_A_36_367#_c_267_p N_A_36_367#_c_247_n
+ N_A_36_367#_c_248_n N_A_36_367#_c_249_n N_A_36_367#_c_252_n
+ N_A_36_367#_c_237_n N_A_36_367#_c_238_n N_A_36_367#_c_298_p
+ PM_SKY130_FD_SC_LP__NOR3_2%A_36_367#
x_PM_SKY130_FD_SC_LP__NOR3_2%VPWR N_VPWR_M1000_d N_VPWR_c_307_n VPWR
+ N_VPWR_c_303_n N_VPWR_c_302_n N_VPWR_c_305_n N_VPWR_c_306_n
+ PM_SKY130_FD_SC_LP__NOR3_2%VPWR
x_PM_SKY130_FD_SC_LP__NOR3_2%A_360_367# N_A_360_367#_M1002_s
+ N_A_360_367#_M1008_s N_A_360_367#_c_351_n N_A_360_367#_c_353_n
+ PM_SKY130_FD_SC_LP__NOR3_2%A_360_367#
x_PM_SKY130_FD_SC_LP__NOR3_2%Y N_Y_M1004_d N_Y_M1010_s N_Y_M1007_s N_Y_M1001_d
+ N_Y_c_372_n N_Y_c_379_n N_Y_c_387_n N_Y_c_429_p N_Y_c_391_n Y Y Y N_Y_c_395_n
+ N_Y_c_380_n Y N_Y_c_427_p N_Y_c_428_p PM_SKY130_FD_SC_LP__NOR3_2%Y
x_PM_SKY130_FD_SC_LP__NOR3_2%VGND N_VGND_M1004_s N_VGND_M1006_s N_VGND_M1003_d
+ N_VGND_M1011_d N_VGND_c_439_n N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n
+ N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_446_n N_VGND_c_447_n
+ N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n VGND N_VGND_c_451_n
+ N_VGND_c_452_n PM_SKY130_FD_SC_LP__NOR3_2%VGND
cc_1 VNB N_A_M1000_g 0.0127772f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.465
cc_2 VNB N_A_c_59_n 0.0214009f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.185
cc_3 VNB N_A_c_60_n 0.0157453f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.185
cc_4 VNB N_A_M1009_g 0.00764983f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=2.465
cc_5 VNB N_A_c_62_n 0.0281911f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.35
cc_6 VNB N_A_c_63_n 0.0686847f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.35
cc_7 VNB N_B_M1010_g 0.0257518f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.465
cc_8 VNB N_B_c_106_n 0.021801f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=0.655
cc_9 VNB N_B_M1005_g 0.00259123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_108_n 8.06644e-19 $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.35
cc_11 VNB N_B_c_109_n 0.0263444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB B 0.0154206f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.35
cc_13 VNB N_B_c_111_n 0.0952637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_c_112_n 0.00380378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_113_n 0.00589554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C_c_183_n 0.0166908f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.515
cc_17 VNB N_C_c_184_n 0.0162434f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.655
cc_18 VNB C 0.00627714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_C_c_186_n 0.0462038f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.35
cc_20 VNB N_VPWR_c_302_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_372_n 0.0043013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_439_n 0.0329366f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB N_VGND_c_440_n 3.21238e-19 $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.35
cc_24 VNB N_VGND_c_441_n 3.23802e-19 $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.35
cc_25 VNB N_VGND_c_442_n 0.0395733f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.35
cc_26 VNB N_VGND_c_443_n 0.0169405f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_27 VNB N_VGND_c_444_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_445_n 0.0133881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_446_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_447_n 0.0140605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_448_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_449_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_450_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_451_n 0.014713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_452_n 0.235075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_A_M1000_g 0.0272056f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.465
cc_37 VPB N_A_M1009_g 0.0218828f $X=-0.19 $Y=1.655 $X2=1.295 $Y2=2.465
cc_38 VPB N_B_M1002_g 0.0192514f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.655
cc_39 VPB N_B_M1005_g 0.0277868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_B_c_108_n 8.76453e-19 $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.35
cc_41 VPB N_B_c_109_n 0.00649147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB B 0.0090301f $X=-0.19 $Y=1.655 $X2=1.295 $Y2=1.35
cc_43 VPB N_B_c_112_n 0.00233975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_B_c_113_n 0.00875732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_C_c_187_n 0.0163164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_C_c_188_n 0.0180209f $X=-0.19 $Y=1.655 $X2=1.295 $Y2=0.655
cc_47 VPB N_C_c_186_n 0.00965699f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=1.35
cc_48 VPB N_A_36_367#_c_234_n 0.046369f $X=-0.19 $Y=1.655 $X2=1.295 $Y2=2.465
cc_49 VPB N_A_36_367#_c_235_n 0.00694896f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_50 VPB N_A_36_367#_c_236_n 0.0106522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_36_367#_c_237_n 0.00747071f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=1.35
cc_52 VPB N_A_36_367#_c_238_n 0.0360021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_303_n 0.063095f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_302_n 0.0469319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_305_n 0.0170261f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.35
cc_56 VPB N_VPWR_c_306_n 0.0123786f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=1.35
cc_57 VPB N_Y_c_372_n 0.00123934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 N_A_c_60_n N_B_M1010_g 0.0365681f $X=1.295 $Y=1.185 $X2=0 $Y2=0
cc_59 N_A_M1009_g N_B_M1002_g 0.035892f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_60 N_A_c_63_n N_B_c_108_n 3.90305e-19 $X=1.295 $Y=1.35 $X2=0 $Y2=0
cc_61 N_A_c_63_n N_B_c_109_n 0.0204229f $X=1.295 $Y=1.35 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_A_36_367#_c_235_n 0.0167816f $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_63 N_A_M1009_g N_A_36_367#_c_235_n 0.00202336f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A_c_62_n N_A_36_367#_c_235_n 0.0574372f $X=1.075 $Y=1.35 $X2=0 $Y2=0
cc_65 N_A_c_63_n N_A_36_367#_c_235_n 0.0110431f $X=1.295 $Y=1.35 $X2=0 $Y2=0
cc_66 N_A_c_62_n N_A_36_367#_c_236_n 0.0225577f $X=1.075 $Y=1.35 $X2=0 $Y2=0
cc_67 N_A_M1000_g N_A_36_367#_c_244_n 0.00134061f $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A_M1009_g N_A_36_367#_c_244_n 0.00942692f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_69 N_A_M1009_g N_A_36_367#_c_246_n 0.0139204f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_M1000_g N_VPWR_c_307_n 0.00810008f $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_71 N_A_M1009_g N_VPWR_c_307_n 0.00240418f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_72 N_A_M1009_g N_VPWR_c_303_n 0.00359504f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A_M1000_g N_VPWR_c_302_n 0.00978874f $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_74 N_A_M1009_g N_VPWR_c_302_n 0.00422763f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_VPWR_c_305_n 0.00525069f $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_76 N_A_M1000_g N_VPWR_c_306_n 0.00889278f $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A_M1009_g N_VPWR_c_306_n 0.00925331f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_c_59_n N_Y_c_372_n 7.19472e-19 $X=0.845 $Y=1.185 $X2=0 $Y2=0
cc_79 N_A_c_60_n N_Y_c_372_n 0.00364053f $X=1.295 $Y=1.185 $X2=0 $Y2=0
cc_80 N_A_M1009_g N_Y_c_372_n 0.0131076f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_81 N_A_c_62_n N_Y_c_372_n 0.0249855f $X=1.075 $Y=1.35 $X2=0 $Y2=0
cc_82 N_A_c_63_n N_Y_c_372_n 0.00766262f $X=1.295 $Y=1.35 $X2=0 $Y2=0
cc_83 N_A_M1009_g N_Y_c_379_n 0.00831302f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_84 N_A_c_60_n N_Y_c_380_n 0.0135942f $X=1.295 $Y=1.185 $X2=0 $Y2=0
cc_85 N_A_c_62_n N_Y_c_380_n 0.0155648f $X=1.075 $Y=1.35 $X2=0 $Y2=0
cc_86 N_A_c_63_n N_Y_c_380_n 0.00279548f $X=1.295 $Y=1.35 $X2=0 $Y2=0
cc_87 N_A_c_59_n N_VGND_c_439_n 0.0163739f $X=0.845 $Y=1.185 $X2=0 $Y2=0
cc_88 N_A_c_60_n N_VGND_c_439_n 6.04604e-19 $X=1.295 $Y=1.185 $X2=0 $Y2=0
cc_89 N_A_c_62_n N_VGND_c_439_n 0.0244884f $X=1.075 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A_c_63_n N_VGND_c_439_n 0.00777197f $X=1.295 $Y=1.35 $X2=0 $Y2=0
cc_91 N_A_c_59_n N_VGND_c_440_n 5.59014e-19 $X=0.845 $Y=1.185 $X2=0 $Y2=0
cc_92 N_A_c_60_n N_VGND_c_440_n 0.00989876f $X=1.295 $Y=1.185 $X2=0 $Y2=0
cc_93 N_A_c_59_n N_VGND_c_445_n 0.00486043f $X=0.845 $Y=1.185 $X2=0 $Y2=0
cc_94 N_A_c_60_n N_VGND_c_445_n 0.00486043f $X=1.295 $Y=1.185 $X2=0 $Y2=0
cc_95 N_A_c_59_n N_VGND_c_452_n 0.00829853f $X=0.845 $Y=1.185 $X2=0 $Y2=0
cc_96 N_A_c_60_n N_VGND_c_452_n 0.00459037f $X=1.295 $Y=1.185 $X2=0 $Y2=0
cc_97 N_B_M1010_g N_C_c_183_n 0.0185609f $X=1.725 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_98 N_B_c_113_n N_C_c_187_n 0.00426107f $X=2.94 $Y=1.535 $X2=0 $Y2=0
cc_99 N_B_c_106_n N_C_c_184_n 0.0174719f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_100 N_B_c_113_n N_C_c_188_n 0.00819707f $X=2.94 $Y=1.535 $X2=0 $Y2=0
cc_101 N_B_M1010_g C 0.00143894f $X=1.725 $Y=0.655 $X2=0 $Y2=0
cc_102 N_B_c_108_n C 0.00729286f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_103 N_B_c_109_n C 6.05664e-19 $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_104 N_B_c_111_n C 0.00255216f $X=3.57 $Y=1.45 $X2=0 $Y2=0
cc_105 N_B_c_112_n C 0.0133662f $X=3.19 $Y=1.535 $X2=0 $Y2=0
cc_106 N_B_c_113_n C 0.0511694f $X=2.94 $Y=1.535 $X2=0 $Y2=0
cc_107 N_B_M1002_g N_C_c_186_n 0.0469311f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_108 N_B_M1005_g N_C_c_186_n 0.0207414f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_109 N_B_c_108_n N_C_c_186_n 0.00136637f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_110 N_B_c_109_n N_C_c_186_n 0.0222753f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_111 N_B_c_111_n N_C_c_186_n 0.0174719f $X=3.57 $Y=1.45 $X2=0 $Y2=0
cc_112 N_B_c_112_n N_C_c_186_n 0.00510435f $X=3.19 $Y=1.535 $X2=0 $Y2=0
cc_113 N_B_c_113_n N_C_c_186_n 0.0194016f $X=2.94 $Y=1.535 $X2=0 $Y2=0
cc_114 N_B_M1002_g N_A_36_367#_c_247_n 0.0102629f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_115 N_B_M1005_g N_A_36_367#_c_248_n 0.0012546f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B_M1005_g N_A_36_367#_c_249_n 0.0134452f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B_c_111_n N_A_36_367#_c_249_n 0.00131854f $X=3.57 $Y=1.45 $X2=0 $Y2=0
cc_118 N_B_c_113_n N_A_36_367#_c_249_n 0.046139f $X=2.94 $Y=1.535 $X2=0 $Y2=0
cc_119 N_B_c_113_n N_A_36_367#_c_252_n 0.0113369f $X=2.94 $Y=1.535 $X2=0 $Y2=0
cc_120 B N_A_36_367#_c_237_n 0.022776f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_121 N_B_c_111_n N_A_36_367#_c_237_n 0.00129585f $X=3.57 $Y=1.45 $X2=0 $Y2=0
cc_122 N_B_M1002_g N_VPWR_c_303_n 0.00419907f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B_M1005_g N_VPWR_c_303_n 0.00547432f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B_M1002_g N_VPWR_c_302_n 0.00604645f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B_M1005_g N_VPWR_c_302_n 0.0115112f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B_M1002_g N_VPWR_c_306_n 0.00122463f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B_M1002_g N_A_360_367#_c_351_n 0.00316013f $X=1.725 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_B_M1005_g N_A_360_367#_c_351_n 0.00795998f $X=3.365 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_B_M1005_g N_A_360_367#_c_353_n 0.00828986f $X=3.365 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_B_M1010_g N_Y_c_372_n 0.00490411f $X=1.725 $Y=0.655 $X2=0 $Y2=0
cc_131 N_B_M1002_g N_Y_c_372_n 0.00442674f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_132 N_B_c_108_n N_Y_c_372_n 0.0318105f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_133 N_B_c_109_n N_Y_c_372_n 0.00209765f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_134 N_B_M1002_g N_Y_c_387_n 0.0178114f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_135 N_B_c_108_n N_Y_c_387_n 0.0128592f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_136 N_B_c_109_n N_Y_c_387_n 0.002022f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_137 N_B_c_113_n N_Y_c_387_n 0.0421147f $X=2.94 $Y=1.535 $X2=0 $Y2=0
cc_138 N_B_c_113_n N_Y_c_391_n 0.00599467f $X=2.94 $Y=1.535 $X2=0 $Y2=0
cc_139 N_B_c_108_n Y 9.43718e-19 $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_140 N_B_c_109_n Y 0.0013844f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_141 N_B_c_113_n Y 0.00572783f $X=2.94 $Y=1.535 $X2=0 $Y2=0
cc_142 N_B_M1010_g N_Y_c_395_n 0.0117896f $X=1.725 $Y=0.655 $X2=0 $Y2=0
cc_143 N_B_c_108_n N_Y_c_395_n 0.00708316f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_144 N_B_c_109_n N_Y_c_395_n 0.00142837f $X=1.755 $Y=1.51 $X2=0 $Y2=0
cc_145 N_B_M1010_g N_VGND_c_440_n 0.00998942f $X=1.725 $Y=0.655 $X2=0 $Y2=0
cc_146 N_B_M1010_g N_VGND_c_441_n 5.45796e-19 $X=1.725 $Y=0.655 $X2=0 $Y2=0
cc_147 N_B_c_106_n N_VGND_c_441_n 5.81548e-19 $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_148 N_B_c_106_n N_VGND_c_442_n 0.00745762f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_149 N_B_c_111_n N_VGND_c_442_n 0.00847824f $X=3.57 $Y=1.45 $X2=0 $Y2=0
cc_150 N_B_c_112_n N_VGND_c_442_n 0.0233497f $X=3.19 $Y=1.535 $X2=0 $Y2=0
cc_151 N_B_M1010_g N_VGND_c_447_n 0.00486043f $X=1.725 $Y=0.655 $X2=0 $Y2=0
cc_152 N_B_c_106_n N_VGND_c_449_n 0.00585385f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_153 N_B_M1010_g N_VGND_c_452_n 0.00468261f $X=1.725 $Y=0.655 $X2=0 $Y2=0
cc_154 N_B_c_106_n N_VGND_c_452_n 0.0116669f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_155 N_C_c_187_n N_A_36_367#_c_247_n 0.0110611f $X=2.205 $Y=1.725 $X2=0 $Y2=0
cc_156 N_C_c_188_n N_A_36_367#_c_247_n 0.0139732f $X=2.635 $Y=1.725 $X2=0 $Y2=0
cc_157 N_C_c_187_n N_A_36_367#_c_248_n 7.86653e-19 $X=2.205 $Y=1.725 $X2=0 $Y2=0
cc_158 N_C_c_188_n N_A_36_367#_c_248_n 0.00901818f $X=2.635 $Y=1.725 $X2=0 $Y2=0
cc_159 N_C_c_188_n N_A_36_367#_c_252_n 0.00569832f $X=2.635 $Y=1.725 $X2=0 $Y2=0
cc_160 N_C_c_187_n N_VPWR_c_303_n 0.00357877f $X=2.205 $Y=1.725 $X2=0 $Y2=0
cc_161 N_C_c_188_n N_VPWR_c_303_n 0.00357877f $X=2.635 $Y=1.725 $X2=0 $Y2=0
cc_162 N_C_c_187_n N_VPWR_c_302_n 0.00549262f $X=2.205 $Y=1.725 $X2=0 $Y2=0
cc_163 N_C_c_188_n N_VPWR_c_302_n 0.00593812f $X=2.635 $Y=1.725 $X2=0 $Y2=0
cc_164 N_C_c_187_n N_A_360_367#_c_351_n 0.0100622f $X=2.205 $Y=1.725 $X2=0 $Y2=0
cc_165 N_C_c_188_n N_A_360_367#_c_351_n 0.0100608f $X=2.635 $Y=1.725 $X2=0 $Y2=0
cc_166 N_C_c_188_n N_A_360_367#_c_353_n 0.00444992f $X=2.635 $Y=1.725 $X2=0
+ $Y2=0
cc_167 C N_Y_c_372_n 0.00504819f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_168 N_C_c_187_n N_Y_c_387_n 0.0132325f $X=2.205 $Y=1.725 $X2=0 $Y2=0
cc_169 N_C_c_186_n N_Y_c_387_n 6.24178e-19 $X=2.635 $Y=1.455 $X2=0 $Y2=0
cc_170 N_C_c_183_n N_Y_c_391_n 0.0105357f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_171 N_C_c_184_n N_Y_c_391_n 0.0105906f $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_172 C N_Y_c_391_n 0.04059f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_173 N_C_c_186_n N_Y_c_391_n 0.00256473f $X=2.635 $Y=1.455 $X2=0 $Y2=0
cc_174 C Y 0.00325646f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_175 N_C_c_183_n N_VGND_c_440_n 5.45796e-19 $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_176 N_C_c_183_n N_VGND_c_441_n 0.0100573f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_177 N_C_c_184_n N_VGND_c_441_n 0.00998663f $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_178 N_C_c_183_n N_VGND_c_447_n 0.00486043f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_179 N_C_c_184_n N_VGND_c_449_n 0.00486043f $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_180 N_C_c_183_n N_VGND_c_452_n 0.00468261f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_181 N_C_c_184_n N_VGND_c_452_n 0.00456652f $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_182 N_A_36_367#_c_235_n N_VPWR_M1000_d 0.00883341f $X=0.99 $Y=1.77 $X2=-0.19
+ $Y2=1.655
cc_183 N_A_36_367#_c_244_n N_VPWR_M1000_d 0.0161459f $X=1.075 $Y=2.465 $X2=-0.19
+ $Y2=1.655
cc_184 N_A_36_367#_c_262_p N_VPWR_M1000_d 0.00403699f $X=1.16 $Y=2.555 $X2=-0.19
+ $Y2=1.655
cc_185 N_A_36_367#_c_235_n N_VPWR_c_307_n 0.0146112f $X=0.99 $Y=1.77 $X2=0 $Y2=0
cc_186 N_A_36_367#_c_244_n N_VPWR_c_307_n 0.0327694f $X=1.075 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_36_367#_c_262_p N_VPWR_c_307_n 0.0149926f $X=1.16 $Y=2.555 $X2=0
+ $Y2=0
cc_188 N_A_36_367#_c_246_n N_VPWR_c_303_n 0.00220098f $X=1.415 $Y=2.555 $X2=0
+ $Y2=0
cc_189 N_A_36_367#_c_267_p N_VPWR_c_303_n 0.0123601f $X=1.51 $Y=2.91 $X2=0 $Y2=0
cc_190 N_A_36_367#_c_247_n N_VPWR_c_303_n 0.00220957f $X=2.675 $Y=2.555 $X2=0
+ $Y2=0
cc_191 N_A_36_367#_c_238_n N_VPWR_c_303_n 0.0178111f $X=3.58 $Y=2.495 $X2=0
+ $Y2=0
cc_192 N_A_36_367#_M1000_s N_VPWR_c_302_n 0.00336915f $X=0.18 $Y=1.835 $X2=0
+ $Y2=0
cc_193 N_A_36_367#_M1009_s N_VPWR_c_302_n 0.00259937f $X=1.37 $Y=1.835 $X2=0
+ $Y2=0
cc_194 N_A_36_367#_M1005_d N_VPWR_c_302_n 0.00371702f $X=3.44 $Y=1.835 $X2=0
+ $Y2=0
cc_195 N_A_36_367#_c_234_n N_VPWR_c_302_n 0.0104192f $X=0.305 $Y=1.98 $X2=0
+ $Y2=0
cc_196 N_A_36_367#_c_246_n N_VPWR_c_302_n 0.00433773f $X=1.415 $Y=2.555 $X2=0
+ $Y2=0
cc_197 N_A_36_367#_c_262_p N_VPWR_c_302_n 7.93477e-19 $X=1.16 $Y=2.555 $X2=0
+ $Y2=0
cc_198 N_A_36_367#_c_267_p N_VPWR_c_302_n 0.00728824f $X=1.51 $Y=2.91 $X2=0
+ $Y2=0
cc_199 N_A_36_367#_c_247_n N_VPWR_c_302_n 0.00554022f $X=2.675 $Y=2.555 $X2=0
+ $Y2=0
cc_200 N_A_36_367#_c_238_n N_VPWR_c_302_n 0.0100304f $X=3.58 $Y=2.495 $X2=0
+ $Y2=0
cc_201 N_A_36_367#_c_234_n N_VPWR_c_305_n 0.0181659f $X=0.305 $Y=1.98 $X2=0
+ $Y2=0
cc_202 N_A_36_367#_c_246_n N_VPWR_c_306_n 0.00189815f $X=1.415 $Y=2.555 $X2=0
+ $Y2=0
cc_203 N_A_36_367#_c_262_p N_VPWR_c_306_n 0.0144549f $X=1.16 $Y=2.555 $X2=0
+ $Y2=0
cc_204 N_A_36_367#_c_247_n N_A_360_367#_M1002_s 0.00454108f $X=2.675 $Y=2.555
+ $X2=-0.19 $Y2=1.655
cc_205 N_A_36_367#_c_247_n N_A_360_367#_M1008_s 0.00258127f $X=2.675 $Y=2.555
+ $X2=0 $Y2=0
cc_206 N_A_36_367#_c_248_n N_A_360_367#_M1008_s 0.00422024f $X=2.76 $Y=2.465
+ $X2=0 $Y2=0
cc_207 N_A_36_367#_c_249_n N_A_360_367#_M1008_s 0.0145455f $X=3.485 $Y=2.04
+ $X2=0 $Y2=0
cc_208 N_A_36_367#_c_252_n N_A_360_367#_M1008_s 8.65676e-19 $X=2.845 $Y=2.04
+ $X2=0 $Y2=0
cc_209 N_A_36_367#_c_247_n N_A_360_367#_c_351_n 0.0558083f $X=2.675 $Y=2.555
+ $X2=0 $Y2=0
cc_210 N_A_36_367#_c_247_n N_A_360_367#_c_353_n 0.015227f $X=2.675 $Y=2.555
+ $X2=0 $Y2=0
cc_211 N_A_36_367#_c_248_n N_A_360_367#_c_353_n 0.012859f $X=2.76 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_A_36_367#_c_249_n N_A_360_367#_c_353_n 0.0194409f $X=3.485 $Y=2.04
+ $X2=0 $Y2=0
cc_213 N_A_36_367#_c_247_n N_Y_M1001_d 0.0034899f $X=2.675 $Y=2.555 $X2=0 $Y2=0
cc_214 N_A_36_367#_M1009_s N_Y_c_372_n 0.00147732f $X=1.37 $Y=1.835 $X2=0 $Y2=0
cc_215 N_A_36_367#_c_235_n N_Y_c_372_n 0.0136794f $X=0.99 $Y=1.77 $X2=0 $Y2=0
cc_216 N_A_36_367#_c_244_n N_Y_c_372_n 0.00765223f $X=1.075 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_36_367#_M1009_s N_Y_c_379_n 7.96769e-19 $X=1.37 $Y=1.835 $X2=0 $Y2=0
cc_218 N_A_36_367#_c_244_n N_Y_c_379_n 0.0259373f $X=1.075 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A_36_367#_c_246_n N_Y_c_379_n 0.00298257f $X=1.415 $Y=2.555 $X2=0 $Y2=0
cc_220 N_A_36_367#_c_298_p N_Y_c_379_n 0.00648413f $X=1.51 $Y=2.55 $X2=0 $Y2=0
cc_221 N_A_36_367#_M1009_s N_Y_c_387_n 0.00444344f $X=1.37 $Y=1.835 $X2=0 $Y2=0
cc_222 N_A_36_367#_c_247_n N_Y_c_387_n 0.0507545f $X=2.675 $Y=2.555 $X2=0 $Y2=0
cc_223 N_A_36_367#_c_298_p N_Y_c_387_n 0.00781324f $X=1.51 $Y=2.55 $X2=0 $Y2=0
cc_224 N_VPWR_c_302_n N_A_360_367#_M1002_s 0.00263789f $X=3.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_225 N_VPWR_c_302_n N_A_360_367#_M1008_s 0.0047303f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_226 N_VPWR_c_303_n N_A_360_367#_c_351_n 0.090655f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_227 N_VPWR_c_302_n N_A_360_367#_c_351_n 0.0569047f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_228 N_VPWR_c_302_n N_Y_M1001_d 0.00225186f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_229 N_A_360_367#_c_351_n N_Y_M1001_d 0.0033716f $X=3.015 $Y=2.945 $X2=0 $Y2=0
cc_230 N_A_360_367#_M1002_s N_Y_c_387_n 0.00462002f $X=1.8 $Y=1.835 $X2=1.87
+ $Y2=1.695
cc_231 N_Y_c_372_n N_VGND_M1006_s 3.8937e-19 $X=1.415 $Y=1.965 $X2=0 $Y2=0
cc_232 N_Y_c_395_n N_VGND_M1006_s 0.00421502f $X=1.845 $Y=0.94 $X2=0 $Y2=0
cc_233 N_Y_c_380_n N_VGND_M1006_s 7.96865e-19 $X=1.5 $Y=0.94 $X2=0 $Y2=0
cc_234 N_Y_c_391_n N_VGND_M1003_d 0.0032907f $X=2.755 $Y=0.94 $X2=0 $Y2=0
cc_235 N_Y_c_395_n N_VGND_c_440_n 0.00921043f $X=1.845 $Y=0.94 $X2=0 $Y2=0
cc_236 N_Y_c_380_n N_VGND_c_440_n 0.00836355f $X=1.5 $Y=0.94 $X2=0 $Y2=0
cc_237 N_Y_c_391_n N_VGND_c_441_n 0.0168833f $X=2.755 $Y=0.94 $X2=0 $Y2=0
cc_238 N_Y_c_427_p N_VGND_c_445_n 0.0138587f $X=1.06 $Y=0.42 $X2=0 $Y2=0
cc_239 N_Y_c_428_p N_VGND_c_447_n 0.0159681f $X=1.965 $Y=0.42 $X2=0 $Y2=0
cc_240 N_Y_c_429_p N_VGND_c_449_n 0.0136943f $X=2.85 $Y=0.42 $X2=0 $Y2=0
cc_241 N_Y_M1004_d N_VGND_c_452_n 0.00424501f $X=0.92 $Y=0.235 $X2=0 $Y2=0
cc_242 N_Y_M1010_s N_VGND_c_452_n 0.00320529f $X=1.8 $Y=0.235 $X2=0 $Y2=0
cc_243 N_Y_M1007_s N_VGND_c_452_n 0.00286727f $X=2.71 $Y=0.235 $X2=0 $Y2=0
cc_244 N_Y_c_429_p N_VGND_c_452_n 0.00866972f $X=2.85 $Y=0.42 $X2=0 $Y2=0
cc_245 N_Y_c_391_n N_VGND_c_452_n 0.0110625f $X=2.755 $Y=0.94 $X2=0 $Y2=0
cc_246 N_Y_c_395_n N_VGND_c_452_n 0.0055623f $X=1.845 $Y=0.94 $X2=0 $Y2=0
cc_247 N_Y_c_380_n N_VGND_c_452_n 0.00557171f $X=1.5 $Y=0.94 $X2=0 $Y2=0
cc_248 N_Y_c_427_p N_VGND_c_452_n 0.00808656f $X=1.06 $Y=0.42 $X2=0 $Y2=0
cc_249 N_Y_c_428_p N_VGND_c_452_n 0.00925289f $X=1.965 $Y=0.42 $X2=0 $Y2=0
