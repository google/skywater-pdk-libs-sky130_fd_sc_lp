* File: sky130_fd_sc_lp__dlrbp_2.spice
* Created: Wed Sep  2 09:46:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrbp_2.pex.spice"
.subckt sky130_fd_sc_lp__dlrbp_2  VNB VPB RESET_B D GATE VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* GATE	GATE
* D	D
* RESET_B	RESET_B
* VPB	VPB
* VNB	VNB
MM1007 N_Q_N_M1007_d N_A_80_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1012 N_Q_N_M1007_d N_A_80_21#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_432_109#_M1009_g N_A_80_21#_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.1113 PD=0.876667 PS=1.37 NRD=64.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1011 N_Q_M1011_d N_A_432_109#_M1011_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2352 PD=1.12 PS=1.75333 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1025 N_Q_M1011_d N_A_432_109#_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1638 PD=1.12 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1002 A_781_51# N_RESET_B_M1002_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1638 PD=1.05 PS=1.23 NRD=7.14 NRS=5.712 M=1 R=5.6 SA=75001.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_A_432_109#_M1005_d N_A_823_25#_M1005_g A_781_51# VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1019 A_1067_119# N_A_432_109#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1013 N_A_823_25#_M1013_d N_A_1109_21#_M1013_g A_1067_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1018 A_1225_119# N_A_1023_405#_M1018_g N_A_823_25#_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_1246_339#_M1024_g A_1225_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75001.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1026 N_A_1246_339#_M1026_d N_D_M1026_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1109_21#_M1010_g N_A_1023_405#_M1010_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_A_1109_21#_M1020_d N_GATE_M1020_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_80_21#_M1006_g N_Q_N_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.17955 PD=3.05 PS=1.545 NRD=0 NRS=0.7683 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_VPWR_M1027_d N_A_80_21#_M1027_g N_Q_N_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.17955 PD=3.05 PS=1.545 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1021_d N_A_432_109#_M1021_g N_A_80_21#_M1021_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.144674 AS=0.1824 PD=1.11495 PS=1.85 NRD=52.6384 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1001 N_Q_M1001_d N_A_432_109#_M1001_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.284826 PD=1.54 PS=2.19505 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75000.5
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1014 N_Q_M1001_d N_A_432_109#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.27405 PD=1.54 PS=1.695 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75000.9
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1003 N_A_432_109#_M1003_d N_RESET_B_M1003_g N_VPWR_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.27405 PD=1.54 PS=1.695 NRD=0 NRS=12.4898 M=1 R=8.4
+ SA=75001.5 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_A_823_25#_M1022_g N_A_432_109#_M1003_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1015 A_981_503# N_A_432_109#_M1015_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0924 AS=0.095025 PD=0.86 PS=0.8175 NRD=77.3816 NRS=46.886 M=1 R=2.8
+ SA=75002.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_823_25#_M1000_d N_A_1023_405#_M1000_g A_981_503# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0855057 AS=0.0924 PD=0.80434 PS=0.86 NRD=46.886 NRS=77.3816 M=1
+ R=2.8 SA=75002.8 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1016 A_1204_459# N_A_1109_21#_M1016_g N_A_823_25#_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0672 AS=0.130294 PD=0.85 PS=1.22566 NRD=15.3857 NRS=0 M=1
+ R=4.26667 SA=75002.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1023 N_VPWR_M1023_d N_A_1246_339#_M1023_g A_1204_459# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1952 AS=0.0672 PD=1.25 PS=0.85 NRD=3.0732 NRS=15.3857 M=1
+ R=4.26667 SA=75002.6 SB=75001 A=0.096 P=1.58 MULT=1
MM1017 N_A_1246_339#_M1017_d N_D_M1017_g N_VPWR_M1023_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1952 PD=1.85 PS=1.25 NRD=6.1464 NRS=98.5 M=1 R=4.26667
+ SA=75003.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1004_d N_A_1109_21#_M1004_g N_A_1023_405#_M1004_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_1109_21#_M1008_d N_GATE_M1008_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=1.5366 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.7175 P=22.73
*
.include "sky130_fd_sc_lp__dlrbp_2.pxi.spice"
*
.ends
*
*
