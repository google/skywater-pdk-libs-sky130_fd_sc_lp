* File: sky130_fd_sc_lp__nand3b_m.pxi.spice
* Created: Wed Sep  2 10:05:13 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3B_M%A_N N_A_N_M1001_g N_A_N_M1000_g N_A_N_c_58_n
+ N_A_N_c_59_n A_N A_N A_N N_A_N_c_61_n PM_SKY130_FD_SC_LP__NAND3B_M%A_N
x_PM_SKY130_FD_SC_LP__NAND3B_M%C N_C_M1002_g N_C_M1007_g N_C_c_99_n N_C_c_100_n
+ N_C_c_101_n C C C N_C_c_103_n PM_SKY130_FD_SC_LP__NAND3B_M%C
x_PM_SKY130_FD_SC_LP__NAND3B_M%B N_B_M1006_g N_B_M1004_g N_B_c_141_n N_B_c_146_n
+ B B B N_B_c_143_n PM_SKY130_FD_SC_LP__NAND3B_M%B
x_PM_SKY130_FD_SC_LP__NAND3B_M%A_37_47# N_A_37_47#_M1001_s N_A_37_47#_M1000_s
+ N_A_37_47#_c_184_n N_A_37_47#_c_179_n N_A_37_47#_M1005_g N_A_37_47#_M1003_g
+ N_A_37_47#_c_180_n N_A_37_47#_c_181_n N_A_37_47#_c_187_n N_A_37_47#_c_182_n
+ N_A_37_47#_c_188_n N_A_37_47#_c_183_n N_A_37_47#_c_190_n N_A_37_47#_c_191_n
+ N_A_37_47#_c_192_n PM_SKY130_FD_SC_LP__NAND3B_M%A_37_47#
x_PM_SKY130_FD_SC_LP__NAND3B_M%VPWR N_VPWR_M1000_d N_VPWR_M1006_d N_VPWR_c_258_n
+ N_VPWR_c_247_n N_VPWR_c_248_n N_VPWR_c_249_n N_VPWR_c_282_p N_VPWR_c_250_n
+ N_VPWR_c_251_n N_VPWR_c_252_n N_VPWR_c_253_n N_VPWR_c_254_n VPWR
+ N_VPWR_c_255_n N_VPWR_c_246_n N_VPWR_c_257_n PM_SKY130_FD_SC_LP__NAND3B_M%VPWR
x_PM_SKY130_FD_SC_LP__NAND3B_M%Y N_Y_M1005_d N_Y_M1002_d N_Y_M1003_d Y Y
+ N_Y_c_283_n Y Y PM_SKY130_FD_SC_LP__NAND3B_M%Y
x_PM_SKY130_FD_SC_LP__NAND3B_M%VGND N_VGND_M1001_d N_VGND_c_312_n VGND
+ N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n PM_SKY130_FD_SC_LP__NAND3B_M%VGND
cc_1 VNB N_A_N_M1001_g 0.0257625f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.445
cc_2 VNB N_A_N_M1000_g 0.00834029f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.165
cc_3 VNB N_A_N_c_58_n 0.0232589f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.345
cc_4 VNB N_A_N_c_59_n 0.0172748f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.51
cc_5 VNB A_N 0.0101883f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_A_N_c_61_n 0.0163756f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.005
cc_7 VNB N_C_M1002_g 0.012187f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.445
cc_8 VNB N_C_c_99_n 0.016341f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.005
cc_9 VNB N_C_c_100_n 0.0209401f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.84
cc_10 VNB N_C_c_101_n 0.0168991f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.345
cc_11 VNB C 0.0080575f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.51
cc_12 VNB N_C_c_103_n 0.0163822f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.005
cc_13 VNB N_B_M1004_g 0.0324122f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.165
cc_14 VNB N_B_c_141_n 0.0121465f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.345
cc_15 VNB B 0.00315826f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_16 VNB N_B_c_143_n 0.0323419f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.005
cc_17 VNB N_A_37_47#_c_179_n 0.0187532f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.005
cc_18 VNB N_A_37_47#_c_180_n 0.0416114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_37_47#_c_181_n 0.025688f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.005
cc_20 VNB N_A_37_47#_c_182_n 0.00933277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_37_47#_c_183_n 0.0489036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_246_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_283_n 0.0503499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB Y 0.00775605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_312_n 0.00472864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_313_n 0.0461976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_314_n 0.149504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_315_n 0.023669f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.005
cc_29 VPB N_A_N_M1000_g 0.0281702f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.165
cc_30 VPB A_N 0.00581397f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_31 VPB N_C_M1002_g 0.0229678f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.445
cc_32 VPB N_B_M1006_g 0.0139846f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.445
cc_33 VPB N_B_c_141_n 0.0012422f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.345
cc_34 VPB N_B_c_146_n 0.0111688f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.51
cc_35 VPB N_A_37_47#_c_184_n 0.0889886f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.165
cc_36 VPB N_A_37_47#_M1003_g 0.0501051f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_37 VPB N_A_37_47#_c_180_n 0.00173387f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_37_47#_c_187_n 0.0219321f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_37_47#_c_188_n 0.0160879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_37_47#_c_183_n 0.023488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_37_47#_c_190_n 0.0173667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_37_47#_c_191_n 0.0419335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_37_47#_c_192_n 0.0171676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_247_n 0.0134523f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.51
cc_45 VPB N_VPWR_c_248_n 0.00629305f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_46 VPB N_VPWR_c_249_n 0.0185522f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_47 VPB N_VPWR_c_250_n 0.0139051f $X=-0.19 $Y=1.655 $X2=0.632 $Y2=0.925
cc_48 VPB N_VPWR_c_251_n 0.00205435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_252_n 0.0258981f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_253_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0.632 $Y2=1.005
cc_51 VPB N_VPWR_c_254_n 0.00210201f $X=-0.19 $Y=1.655 $X2=0.632 $Y2=1.295
cc_52 VPB N_VPWR_c_255_n 0.0213956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_246_n 0.0802488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_257_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB Y 0.0341839f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 N_A_N_c_59_n N_C_M1002_g 0.0309871f $X=0.545 $Y=1.51 $X2=0 $Y2=0
cc_57 A_N N_C_M1002_g 0.00679089f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_58 N_A_N_M1001_g N_C_c_99_n 0.00955783f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_59 N_A_N_c_58_n N_C_c_100_n 0.0119097f $X=0.545 $Y=1.345 $X2=0 $Y2=0
cc_60 N_A_N_c_59_n N_C_c_101_n 0.0119097f $X=0.545 $Y=1.51 $X2=0 $Y2=0
cc_61 N_A_N_M1001_g C 0.00379541f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_62 A_N C 0.0412837f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_63 N_A_N_c_61_n C 5.54644e-19 $X=0.545 $Y=1.005 $X2=0 $Y2=0
cc_64 N_A_N_M1001_g N_C_c_103_n 0.00278948f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_65 A_N N_C_c_103_n 0.00403425f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_66 N_A_N_c_61_n N_C_c_103_n 0.0119097f $X=0.545 $Y=1.005 $X2=0 $Y2=0
cc_67 N_A_N_M1001_g N_A_37_47#_c_182_n 0.00379512f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_68 A_N N_A_37_47#_c_182_n 8.15844e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_69 N_A_N_c_61_n N_A_37_47#_c_182_n 0.00179161f $X=0.545 $Y=1.005 $X2=0 $Y2=0
cc_70 N_A_N_M1000_g N_A_37_47#_c_188_n 0.00268538f $X=0.635 $Y=2.165 $X2=0 $Y2=0
cc_71 N_A_N_c_59_n N_A_37_47#_c_188_n 0.00275567f $X=0.545 $Y=1.51 $X2=0 $Y2=0
cc_72 A_N N_A_37_47#_c_188_n 0.00477326f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_73 N_A_N_M1001_g N_A_37_47#_c_183_n 0.00701047f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_N_M1000_g N_A_37_47#_c_183_n 0.0107179f $X=0.635 $Y=2.165 $X2=0 $Y2=0
cc_75 A_N N_A_37_47#_c_183_n 0.0666584f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_76 N_A_N_c_61_n N_A_37_47#_c_183_n 0.0163648f $X=0.545 $Y=1.005 $X2=0 $Y2=0
cc_77 N_A_N_M1000_g N_A_37_47#_c_190_n 8.78795e-19 $X=0.635 $Y=2.165 $X2=0 $Y2=0
cc_78 N_A_N_M1000_g N_A_37_47#_c_191_n 0.0101002f $X=0.635 $Y=2.165 $X2=0 $Y2=0
cc_79 N_A_N_M1000_g N_A_37_47#_c_192_n 0.00458034f $X=0.635 $Y=2.165 $X2=0 $Y2=0
cc_80 A_N N_VPWR_c_258_n 0.00215917f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_81 N_A_N_M1000_g N_VPWR_c_251_n 0.00107303f $X=0.635 $Y=2.165 $X2=0 $Y2=0
cc_82 N_A_N_M1000_g Y 0.00154119f $X=0.635 $Y=2.165 $X2=0 $Y2=0
cc_83 A_N Y 0.00187765f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A_N_M1001_g N_VGND_c_312_n 0.0030202f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_85 A_N N_VGND_c_312_n 0.00803394f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_86 N_A_N_c_61_n N_VGND_c_312_n 3.85626e-19 $X=0.545 $Y=1.005 $X2=0 $Y2=0
cc_87 N_A_N_M1001_g N_VGND_c_314_n 0.00769505f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_88 A_N N_VGND_c_314_n 0.00659976f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_89 N_A_N_M1001_g N_VGND_c_315_n 0.00552362f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_90 N_C_c_99_n N_B_M1004_g 0.0410294f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_91 C N_B_M1004_g 0.00548494f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_92 N_C_M1002_g N_B_c_146_n 0.0217434f $X=1.065 $Y=2.165 $X2=0 $Y2=0
cc_93 N_C_c_99_n B 0.00107684f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_94 C B 0.0608089f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_95 N_C_M1002_g N_B_c_143_n 0.00929001f $X=1.065 $Y=2.165 $X2=0 $Y2=0
cc_96 N_C_c_100_n N_B_c_143_n 0.0410294f $X=1.09 $Y=1.27 $X2=0 $Y2=0
cc_97 N_C_M1002_g N_A_37_47#_c_184_n 0.00415463f $X=1.065 $Y=2.165 $X2=0 $Y2=0
cc_98 C N_A_37_47#_c_182_n 0.00220043f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_99 N_C_c_101_n N_VPWR_c_258_n 2.53281e-19 $X=1.09 $Y=1.435 $X2=0 $Y2=0
cc_100 N_C_M1002_g N_VPWR_c_248_n 0.00696628f $X=1.065 $Y=2.165 $X2=0 $Y2=0
cc_101 N_C_M1002_g N_VPWR_c_251_n 0.0051066f $X=1.065 $Y=2.165 $X2=0 $Y2=0
cc_102 N_C_M1002_g Y 0.0121261f $X=1.065 $Y=2.165 $X2=0 $Y2=0
cc_103 N_C_c_101_n Y 8.11051e-19 $X=1.09 $Y=1.435 $X2=0 $Y2=0
cc_104 C Y 0.0101154f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_105 C N_VGND_M1001_d 0.0029947f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_106 N_C_c_99_n N_VGND_c_312_n 0.00675011f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_107 C N_VGND_c_312_n 0.00542328f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_108 N_C_c_99_n N_VGND_c_313_n 0.00398598f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_109 C N_VGND_c_313_n 0.00665758f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_110 N_C_c_103_n N_VGND_c_313_n 0.00185892f $X=1.09 $Y=0.93 $X2=0 $Y2=0
cc_111 N_C_c_99_n N_VGND_c_314_n 0.00600116f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_112 C N_VGND_c_314_n 0.0087435f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_113 N_C_c_103_n N_VGND_c_314_n 0.00214436f $X=1.09 $Y=0.93 $X2=0 $Y2=0
cc_114 N_B_M1006_g N_A_37_47#_c_184_n 0.00404438f $X=1.495 $Y=2.165 $X2=0 $Y2=0
cc_115 N_B_M1004_g N_A_37_47#_c_179_n 0.0506303f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_116 B N_A_37_47#_c_179_n 0.00256773f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_117 N_B_M1004_g N_A_37_47#_c_180_n 0.00306742f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_118 N_B_c_141_n N_A_37_47#_c_180_n 0.00363384f $X=1.517 $Y=1.675 $X2=0 $Y2=0
cc_119 B N_A_37_47#_c_180_n 7.02187e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_120 N_B_c_143_n N_A_37_47#_c_180_n 0.017344f $X=1.63 $Y=1.29 $X2=0 $Y2=0
cc_121 N_B_M1006_g N_A_37_47#_c_187_n 0.0139218f $X=1.495 $Y=2.165 $X2=0 $Y2=0
cc_122 N_B_c_146_n N_A_37_47#_c_187_n 0.00731964f $X=1.517 $Y=1.825 $X2=0 $Y2=0
cc_123 N_B_M1006_g N_VPWR_c_248_n 0.00986173f $X=1.495 $Y=2.165 $X2=0 $Y2=0
cc_124 N_B_c_146_n N_VPWR_c_248_n 2.21149e-19 $X=1.517 $Y=1.825 $X2=0 $Y2=0
cc_125 N_B_M1004_g N_Y_c_283_n 8.64744e-19 $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_126 N_B_c_141_n N_Y_c_283_n 0.00246305f $X=1.517 $Y=1.675 $X2=0 $Y2=0
cc_127 B N_Y_c_283_n 0.0635992f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_128 N_B_c_143_n N_Y_c_283_n 0.00329787f $X=1.63 $Y=1.29 $X2=0 $Y2=0
cc_129 N_B_M1006_g Y 0.0102999f $X=1.495 $Y=2.165 $X2=0 $Y2=0
cc_130 N_B_c_141_n Y 0.00424754f $X=1.517 $Y=1.675 $X2=0 $Y2=0
cc_131 N_B_c_146_n Y 0.0111003f $X=1.517 $Y=1.825 $X2=0 $Y2=0
cc_132 B Y 0.020506f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_133 N_B_c_143_n Y 0.00441557f $X=1.63 $Y=1.29 $X2=0 $Y2=0
cc_134 N_B_M1004_g N_VGND_c_313_n 0.00399843f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_135 B N_VGND_c_313_n 0.00814594f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 N_B_M1004_g N_VGND_c_314_n 0.00531224f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_137 B N_VGND_c_314_n 0.0104566f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_138 B A_323_47# 0.00139886f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_139 N_A_37_47#_c_184_n N_VPWR_c_247_n 0.0154483f $X=1.85 $Y=2.97 $X2=0 $Y2=0
cc_140 N_A_37_47#_c_190_n N_VPWR_c_247_n 0.0248188f $X=0.575 $Y=2.88 $X2=0 $Y2=0
cc_141 N_A_37_47#_c_191_n N_VPWR_c_247_n 0.00423018f $X=0.575 $Y=2.88 $X2=0
+ $Y2=0
cc_142 N_A_37_47#_c_192_n N_VPWR_c_247_n 0.00936092f $X=0.477 $Y=2.715 $X2=0
+ $Y2=0
cc_143 N_A_37_47#_c_184_n N_VPWR_c_248_n 0.0138228f $X=1.85 $Y=2.97 $X2=0 $Y2=0
cc_144 N_A_37_47#_c_184_n N_VPWR_c_249_n 0.0171156f $X=1.85 $Y=2.97 $X2=0 $Y2=0
cc_145 N_A_37_47#_c_184_n N_VPWR_c_250_n 0.0197724f $X=1.85 $Y=2.97 $X2=0 $Y2=0
cc_146 N_A_37_47#_M1003_g N_VPWR_c_250_n 0.0135453f $X=1.925 $Y=2.165 $X2=0
+ $Y2=0
cc_147 N_A_37_47#_c_184_n N_VPWR_c_251_n 0.00338061f $X=1.85 $Y=2.97 $X2=0 $Y2=0
cc_148 N_A_37_47#_c_192_n N_VPWR_c_251_n 0.0138527f $X=0.477 $Y=2.715 $X2=0
+ $Y2=0
cc_149 N_A_37_47#_c_190_n N_VPWR_c_252_n 0.025398f $X=0.575 $Y=2.88 $X2=0 $Y2=0
cc_150 N_A_37_47#_c_191_n N_VPWR_c_252_n 0.00692277f $X=0.575 $Y=2.88 $X2=0
+ $Y2=0
cc_151 N_A_37_47#_M1003_g N_VPWR_c_254_n 0.00595032f $X=1.925 $Y=2.165 $X2=0
+ $Y2=0
cc_152 N_A_37_47#_c_184_n N_VPWR_c_255_n 0.00703326f $X=1.85 $Y=2.97 $X2=0 $Y2=0
cc_153 N_A_37_47#_c_190_n N_VPWR_c_246_n 0.0166926f $X=0.575 $Y=2.88 $X2=0 $Y2=0
cc_154 N_A_37_47#_c_191_n N_VPWR_c_246_n 0.0284278f $X=0.575 $Y=2.88 $X2=0 $Y2=0
cc_155 N_A_37_47#_c_179_n N_Y_c_283_n 0.00261673f $X=1.9 $Y=0.765 $X2=0 $Y2=0
cc_156 N_A_37_47#_c_180_n N_Y_c_283_n 0.0235911f $X=2.11 $Y=1.695 $X2=0 $Y2=0
cc_157 N_A_37_47#_c_181_n N_Y_c_283_n 0.0125605f $X=2.11 $Y=0.84 $X2=0 $Y2=0
cc_158 N_A_37_47#_M1003_g Y 0.0130995f $X=1.925 $Y=2.165 $X2=0 $Y2=0
cc_159 N_A_37_47#_c_180_n Y 0.00390941f $X=2.11 $Y=1.695 $X2=0 $Y2=0
cc_160 N_A_37_47#_c_181_n Y 0.00409795f $X=2.11 $Y=0.84 $X2=0 $Y2=0
cc_161 N_A_37_47#_c_187_n Y 0.0162157f $X=2.11 $Y=1.77 $X2=0 $Y2=0
cc_162 N_A_37_47#_c_179_n N_VGND_c_313_n 0.00585385f $X=1.9 $Y=0.765 $X2=0 $Y2=0
cc_163 N_A_37_47#_c_181_n N_VGND_c_313_n 5.32744e-19 $X=2.11 $Y=0.84 $X2=0 $Y2=0
cc_164 N_A_37_47#_M1001_s N_VGND_c_314_n 0.00236056f $X=0.185 $Y=0.235 $X2=0
+ $Y2=0
cc_165 N_A_37_47#_c_179_n N_VGND_c_314_n 0.0118418f $X=1.9 $Y=0.765 $X2=0 $Y2=0
cc_166 N_A_37_47#_c_182_n N_VGND_c_314_n 0.0123647f $X=0.31 $Y=0.51 $X2=0 $Y2=0
cc_167 N_A_37_47#_c_182_n N_VGND_c_315_n 0.011147f $X=0.31 $Y=0.51 $X2=0 $Y2=0
cc_168 N_VPWR_c_248_n Y 0.0254895f $X=1.625 $Y=2.46 $X2=0 $Y2=0
cc_169 N_VPWR_c_282_p Y 0.0138662f $X=1.71 $Y=2.23 $X2=0 $Y2=0
cc_170 N_Y_c_283_n N_VGND_c_313_n 0.0107327f $X=2.14 $Y=0.51 $X2=0 $Y2=0
cc_171 N_Y_M1005_d N_VGND_c_314_n 0.0025776f $X=1.975 $Y=0.235 $X2=0 $Y2=0
cc_172 N_Y_c_283_n N_VGND_c_314_n 0.011704f $X=2.14 $Y=0.51 $X2=0 $Y2=0
cc_173 N_VGND_c_314_n A_251_47# 0.00802611f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
cc_174 N_VGND_c_314_n A_323_47# 0.00301913f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
