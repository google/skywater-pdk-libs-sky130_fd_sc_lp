* File: sky130_fd_sc_lp__and3b_m.pex.spice
* Created: Wed Sep  2 09:32:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3B_M%A_N 2 5 9 11 12 13 14 15 16 23
r29 23 25 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.327 $Y=1.005
+ $X2=0.327 $Y2=0.84
r30 15 16 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r31 14 15 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r32 13 14 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r33 12 13 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.295
r34 12 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r35 9 11 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=0.475 $Y=2.77
+ $X2=0.475 $Y2=1.51
r36 5 25 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.475 $Y=0.475
+ $X2=0.475 $Y2=0.84
r37 2 11 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=0.327 $Y=1.288
+ $X2=0.327 $Y2=1.51
r38 1 23 7.12377 $w=4.45e-07 $l=5.7e-08 $layer=POLY_cond $X=0.327 $Y=1.062
+ $X2=0.327 $Y2=1.005
r39 1 2 28.2451 $w=4.45e-07 $l=2.26e-07 $layer=POLY_cond $X=0.327 $Y=1.062
+ $X2=0.327 $Y2=1.288
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_M%A_110_53# 1 2 8 9 11 12 15 19 22 25 29 32 33
r56 32 35 16.7741 $w=4.53e-07 $l=5.05e-07 $layer=LI1_cond $X=0.812 $Y=0.96
+ $X2=0.812 $Y2=1.465
r57 32 34 7.83639 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.812 $Y=0.96
+ $X2=0.812 $Y2=0.795
r58 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=0.96 $X2=0.955 $Y2=0.96
r59 29 35 72.355 $w=2.08e-07 $l=1.37e-06 $layer=LI1_cond $X=0.69 $Y=2.835
+ $X2=0.69 $Y2=1.465
r60 25 34 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=0.69 $Y=0.495 $X2=0.69
+ $Y2=0.795
r61 21 33 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.955 $Y=1.315
+ $X2=0.955 $Y2=0.96
r62 21 22 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=0.955 $Y=1.315
+ $X2=0.955 $Y2=1.39
r63 17 19 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.445 $Y=1.315
+ $X2=1.445 $Y2=0.475
r64 13 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.44 $Y=1.855
+ $X2=1.44 $Y2=2.225
r65 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.365 $Y=1.78
+ $X2=1.44 $Y2=1.855
r66 11 12 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.365 $Y=1.78
+ $X2=1.12 $Y2=1.78
r67 10 22 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.39
+ $X2=0.955 $Y2=1.39
r68 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.37 $Y=1.39
+ $X2=1.445 $Y2=1.315
r69 9 10 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.37 $Y=1.39 $X2=1.12
+ $Y2=1.39
r70 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.045 $Y=1.705
+ $X2=1.12 $Y2=1.78
r71 7 22 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.045 $Y=1.465
+ $X2=0.955 $Y2=1.39
r72 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.045 $Y=1.465
+ $X2=1.045 $Y2=1.705
r73 2 29 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.56 $X2=0.69 $Y2=2.835
r74 1 25 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.265 $X2=0.69 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_M%B 3 6 9 10 11 12 13 14 19
r44 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.895
+ $Y=0.96 $X2=1.895 $Y2=0.96
r45 14 20 10.0278 $w=3.83e-07 $l=3.35e-07 $layer=LI1_cond $X=1.787 $Y=1.295
+ $X2=1.787 $Y2=0.96
r46 13 20 1.04768 $w=3.83e-07 $l=3.5e-08 $layer=LI1_cond $X=1.787 $Y=0.925
+ $X2=1.787 $Y2=0.96
r47 12 13 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.787 $Y=0.555
+ $X2=1.787 $Y2=0.925
r48 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.895 $Y=1.3
+ $X2=1.895 $Y2=0.96
r49 10 11 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.3
+ $X2=1.895 $Y2=1.465
r50 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=0.795
+ $X2=1.895 $Y2=0.96
r51 6 11 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.87 $Y=2.225
+ $X2=1.87 $Y2=1.465
r52 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.805 $Y=0.475
+ $X2=1.805 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_M%C 3 7 10 11 14 15 16 21
r42 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.435
+ $Y=1.35 $X2=2.435 $Y2=1.35
r43 16 22 9.68052 $w=3.73e-07 $l=3.15e-07 $layer=LI1_cond $X=2.537 $Y=1.665
+ $X2=2.537 $Y2=1.35
r44 15 22 1.69025 $w=3.73e-07 $l=5.5e-08 $layer=LI1_cond $X=2.537 $Y=1.295
+ $X2=2.537 $Y2=1.35
r45 14 15 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.537 $Y=0.925
+ $X2=2.537 $Y2=1.295
r46 13 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.185
+ $X2=2.435 $Y2=1.35
r47 10 21 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.435 $Y=1.705
+ $X2=2.435 $Y2=1.35
r48 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.412 $Y=1.705
+ $X2=2.412 $Y2=1.855
r49 7 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.345 $Y=0.475
+ $X2=2.345 $Y2=1.185
r50 3 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.3 $Y=2.225 $X2=2.3
+ $Y2=1.855
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_M%A_220_53# 1 2 3 10 12 14 18 20 21 26 30 32
+ 37 38
r71 38 42 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.145 $Y=2.94
+ $X2=2.145 $Y2=3.03
r72 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.145
+ $Y=2.94 $X2=2.145 $Y2=2.94
r73 32 34 15.3138 $w=2.39e-07 $l=3e-07 $layer=LI1_cond $X=1.255 $Y=1.86
+ $X2=1.255 $Y2=2.16
r74 28 30 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.225 $Y=0.51
+ $X2=1.305 $Y2=0.51
r75 24 37 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=2.855
+ $X2=2.075 $Y2=2.94
r76 24 26 40.5694 $w=1.88e-07 $l=6.95e-07 $layer=LI1_cond $X=2.075 $Y=2.855
+ $X2=2.075 $Y2=2.16
r77 23 26 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=2.075 $Y=1.945
+ $X2=2.075 $Y2=2.16
r78 22 32 2.73298 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.39 $Y=1.86
+ $X2=1.255 $Y2=1.86
r79 21 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.98 $Y=1.86
+ $X2=2.075 $Y2=1.945
r80 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.98 $Y=1.86 $X2=1.39
+ $Y2=1.86
r81 20 32 5.37298 $w=2.39e-07 $l=1.07121e-07 $layer=LI1_cond $X=1.305 $Y=1.775
+ $X2=1.255 $Y2=1.86
r82 19 30 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.305 $Y=0.615
+ $X2=1.305 $Y2=0.51
r83 19 20 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=1.305 $Y=0.615
+ $X2=1.305 $Y2=1.775
r84 16 18 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.885 $Y=2.955
+ $X2=2.885 $Y2=2.225
r85 15 18 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=2.885 $Y=1.095
+ $X2=2.885 $Y2=2.225
r86 12 15 61.5319 $w=2.35e-07 $l=3.50714e-07 $layer=POLY_cond $X=2.775 $Y=0.795
+ $X2=2.885 $Y2=1.095
r87 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.775 $Y=0.795
+ $X2=2.775 $Y2=0.475
r88 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=3.03
+ $X2=2.145 $Y2=3.03
r89 10 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.81 $Y=3.03
+ $X2=2.885 $Y2=2.955
r90 10 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.81 $Y=3.03 $X2=2.31
+ $Y2=3.03
r91 3 26 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=2.015 $X2=2.085 $Y2=2.16
r92 2 34 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=2.015 $X2=1.225 $Y2=2.16
r93 1 28 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.265 $X2=1.225 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_M%VPWR 1 2 3 10 12 16 20 23 24 26 27 28 38 39
r46 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 33 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 30 42 3.52379 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=3.33
+ $X2=0.172 $Y2=3.33
r53 30 32 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=0.345 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 28 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 26 35 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 26 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.595 $Y2=3.33
r58 25 38 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.7 $Y=3.33 $X2=3.12
+ $Y2=3.33
r59 25 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.7 $Y=3.33
+ $X2=2.595 $Y2=3.33
r60 23 32 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 23 24 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=1.665 $Y2=3.33
r62 22 35 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.76 $Y=3.33 $X2=2.16
+ $Y2=3.33
r63 22 24 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.76 $Y=3.33
+ $X2=1.665 $Y2=3.33
r64 18 27 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=3.33
r65 18 20 50.4372 $w=2.08e-07 $l=9.55e-07 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=2.29
r66 14 24 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=3.245
+ $X2=1.665 $Y2=3.33
r67 14 16 55.7464 $w=1.88e-07 $l=9.55e-07 $layer=LI1_cond $X=1.665 $Y=3.245
+ $X2=1.665 $Y2=2.29
r68 10 42 3.3201 $w=1.9e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.25 $Y=3.245
+ $X2=0.172 $Y2=3.33
r69 10 12 23.933 $w=1.88e-07 $l=4.1e-07 $layer=LI1_cond $X=0.25 $Y=3.245
+ $X2=0.25 $Y2=2.835
r70 3 20 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=2.015 $X2=2.595 $Y2=2.29
r71 2 16 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=2.015 $X2=1.655 $Y2=2.29
r72 1 12 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.56 $X2=0.26 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_M%X 1 2 7 8 9 10 11 12 20
r12 12 33 3.68142 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=3.085 $Y=2.405
+ $X2=3.085 $Y2=2.29
r13 11 33 8.16314 $w=3.58e-07 $l=2.55e-07 $layer=LI1_cond $X=3.085 $Y=2.035
+ $X2=3.085 $Y2=2.29
r14 10 11 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.085 $Y=1.665
+ $X2=3.085 $Y2=2.035
r15 9 10 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.085 $Y=1.295
+ $X2=3.085 $Y2=1.665
r16 8 9 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.085 $Y=0.925
+ $X2=3.085 $Y2=1.295
r17 7 8 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.085 $Y=0.555
+ $X2=3.085 $Y2=0.925
r18 7 20 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=3.085 $Y=0.555
+ $X2=3.085 $Y2=0.54
r19 2 33 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=2.015 $X2=3.1 $Y2=2.29
r20 1 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.265 $X2=2.99 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_M%VGND 1 2 7 9 13 15 17 27 28 34
r40 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r42 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r43 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.56
+ $Y2=0
r45 25 27 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=3.12
+ $Y2=0
r46 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r47 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r49 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r50 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r51 18 31 3.65746 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r52 18 20 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r53 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.56
+ $Y2=0
r54 17 23 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.16
+ $Y2=0
r55 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r56 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r57 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r58 11 13 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.41
r59 7 31 3.25773 $w=2.1e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.182 $Y2=0
r60 7 9 17.1645 $w=2.08e-07 $l=3.25e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.41
r61 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.42
+ $Y=0.265 $X2=2.56 $Y2=0.41
r62 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.41
.ends

