* File: sky130_fd_sc_lp__srsdfxtp_1.pxi.spice
* Created: Wed Sep  2 10:39:30 2020
* 
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%SCE N_SCE_c_292_n N_SCE_c_302_n N_SCE_M1030_g
+ N_SCE_M1040_g N_SCE_c_303_n N_SCE_c_304_n N_SCE_c_305_n N_SCE_M1000_g
+ N_SCE_M1018_g N_SCE_c_295_n N_SCE_c_296_n N_SCE_c_297_n SCE N_SCE_c_299_n
+ N_SCE_c_300_n PM_SKY130_FD_SC_LP__SRSDFXTP_1%SCE
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_31_477# N_A_31_477#_M1040_s
+ N_A_31_477#_M1030_s N_A_31_477#_M1037_g N_A_31_477#_M1004_g
+ N_A_31_477#_c_395_n N_A_31_477#_c_401_n N_A_31_477#_c_402_n
+ N_A_31_477#_c_403_n N_A_31_477#_c_404_n N_A_31_477#_c_396_n
+ N_A_31_477#_c_405_n N_A_31_477#_c_397_n N_A_31_477#_c_398_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_31_477#
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%D N_D_M1021_g N_D_M1003_g D N_D_c_487_n
+ N_D_c_488_n PM_SKY130_FD_SC_LP__SRSDFXTP_1%D
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%SCD N_SCD_M1039_g N_SCD_M1016_g N_SCD_c_522_n
+ SCD N_SCD_c_525_n N_SCD_c_526_n N_SCD_c_523_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%SCD
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_570_47# N_A_570_47#_M1025_d
+ N_A_570_47#_M1027_d N_A_570_47#_c_576_n N_A_570_47#_c_601_n
+ N_A_570_47#_M1008_g N_A_570_47#_c_602_n N_A_570_47#_M1035_g
+ N_A_570_47#_c_578_n N_A_570_47#_M1028_g N_A_570_47#_c_579_n
+ N_A_570_47#_M1012_g N_A_570_47#_c_603_n N_A_570_47#_M1001_g
+ N_A_570_47#_c_604_n N_A_570_47#_c_580_n N_A_570_47#_c_606_n
+ N_A_570_47#_c_607_n N_A_570_47#_c_608_n N_A_570_47#_c_581_n
+ N_A_570_47#_c_582_n N_A_570_47#_c_583_n N_A_570_47#_c_584_n
+ N_A_570_47#_c_633_p N_A_570_47#_c_585_n N_A_570_47#_c_586_n
+ N_A_570_47#_c_587_n N_A_570_47#_c_588_n N_A_570_47#_c_589_n
+ N_A_570_47#_c_590_n N_A_570_47#_c_591_n N_A_570_47#_c_592_n
+ N_A_570_47#_c_593_n N_A_570_47#_c_594_n N_A_570_47#_c_595_n
+ N_A_570_47#_c_596_n N_A_570_47#_c_597_n N_A_570_47#_c_598_n
+ N_A_570_47#_c_599_n N_A_570_47#_c_611_n N_A_570_47#_c_600_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_570_47#
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_914_245# N_A_914_245#_M1038_d
+ N_A_914_245#_M1023_d N_A_914_245#_M1034_g N_A_914_245#_M1036_g
+ N_A_914_245#_c_823_n N_A_914_245#_c_824_n N_A_914_245#_c_825_n
+ N_A_914_245#_c_842_n N_A_914_245#_c_844_n N_A_914_245#_c_826_n
+ N_A_914_245#_c_831_n N_A_914_245#_c_832_n N_A_914_245#_c_833_n
+ N_A_914_245#_c_827_n N_A_914_245#_c_834_n N_A_914_245#_c_828_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_914_245#
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_786_139# N_A_786_139#_M1005_d
+ N_A_786_139#_M1035_d N_A_786_139#_M1038_g N_A_786_139#_c_929_n
+ N_A_786_139#_M1023_g N_A_786_139#_c_930_n N_A_786_139#_c_931_n
+ N_A_786_139#_c_926_n N_A_786_139#_c_933_n N_A_786_139#_c_934_n
+ N_A_786_139#_c_935_n N_A_786_139#_c_936_n N_A_786_139#_c_937_n
+ N_A_786_139#_c_927_n N_A_786_139#_c_939_n N_A_786_139#_c_940_n
+ N_A_786_139#_c_941_n N_A_786_139#_c_942_n N_A_786_139#_c_943_n
+ N_A_786_139#_c_944_n N_A_786_139#_c_928_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_786_139#
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_540_21# N_A_540_21#_M1013_s
+ N_A_540_21#_M1010_d N_A_540_21#_M1025_g N_A_540_21#_c_1069_n
+ N_A_540_21#_M1027_g N_A_540_21#_c_1085_n N_A_540_21#_M1005_g
+ N_A_540_21#_c_1087_n N_A_540_21#_M1022_g N_A_540_21#_c_1089_n
+ N_A_540_21#_c_1071_n N_A_540_21#_c_1091_n N_A_540_21#_M1009_g
+ N_A_540_21#_c_1072_n N_A_540_21#_c_1093_n N_A_540_21#_M1014_g
+ N_A_540_21#_M1026_g N_A_540_21#_c_1074_n N_A_540_21#_c_1075_n
+ N_A_540_21#_c_1095_n N_A_540_21#_c_1096_n N_A_540_21#_c_1097_n
+ N_A_540_21#_c_1076_n N_A_540_21#_c_1077_n N_A_540_21#_c_1078_n
+ N_A_540_21#_c_1101_n N_A_540_21#_c_1102_n N_A_540_21#_c_1103_n
+ N_A_540_21#_c_1079_n N_A_540_21#_c_1080_n N_A_540_21#_c_1105_n
+ N_A_540_21#_c_1106_n N_A_540_21#_c_1107_n N_A_540_21#_c_1108_n
+ N_A_540_21#_c_1081_n N_A_540_21#_c_1082_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_540_21#
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_1319_69# N_A_1319_69#_M1012_d
+ N_A_1319_69#_M1014_d N_A_1319_69#_M1001_s N_A_1319_69#_M1020_g
+ N_A_1319_69#_M1007_g N_A_1319_69#_c_1326_n N_A_1319_69#_M1029_g
+ N_A_1319_69#_c_1327_n N_A_1319_69#_c_1328_n N_A_1319_69#_c_1314_n
+ N_A_1319_69#_c_1315_n N_A_1319_69#_M1032_g N_A_1319_69#_c_1330_n
+ N_A_1319_69#_M1011_g N_A_1319_69#_c_1317_n N_A_1319_69#_c_1318_n
+ N_A_1319_69#_c_1319_n N_A_1319_69#_c_1320_n N_A_1319_69#_c_1321_n
+ N_A_1319_69#_c_1322_n N_A_1319_69#_c_1323_n N_A_1319_69#_c_1334_n
+ N_A_1319_69#_c_1335_n N_A_1319_69#_c_1358_n N_A_1319_69#_c_1336_n
+ N_A_1319_69#_c_1337_n N_A_1319_69#_c_1338_n N_A_1319_69#_c_1339_n
+ N_A_1319_69#_c_1401_n N_A_1319_69#_c_1402_n N_A_1319_69#_c_1448_p
+ N_A_1319_69#_c_1477_p N_A_1319_69#_c_1340_n N_A_1319_69#_c_1341_n
+ N_A_1319_69#_c_1359_n N_A_1319_69#_c_1324_n N_A_1319_69#_c_1342_n
+ N_A_1319_69#_c_1325_n N_A_1319_69#_c_1344_n N_A_1319_69#_c_1345_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_1319_69#
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_1493_21# N_A_1493_21#_M1007_d
+ N_A_1493_21#_M1029_d N_A_1493_21#_M1019_g N_A_1493_21#_c_1529_n
+ N_A_1493_21#_c_1530_n N_A_1493_21#_M1006_g N_A_1493_21#_c_1532_n
+ N_A_1493_21#_c_1533_n N_A_1493_21#_c_1546_n N_A_1493_21#_M1017_g
+ N_A_1493_21#_c_1534_n N_A_1493_21#_c_1535_n N_A_1493_21#_c_1536_n
+ N_A_1493_21#_c_1537_n N_A_1493_21#_c_1538_n N_A_1493_21#_c_1539_n
+ N_A_1493_21#_c_1549_n N_A_1493_21#_c_1583_n N_A_1493_21#_c_1550_n
+ N_A_1493_21#_c_1540_n N_A_1493_21#_c_1541_n N_A_1493_21#_c_1542_n
+ N_A_1493_21#_c_1543_n N_A_1493_21#_c_1544_n N_A_1493_21#_c_1545_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_1493_21#
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%SLEEP_B N_SLEEP_B_M1010_g N_SLEEP_B_M1002_g
+ N_SLEEP_B_c_1684_n N_SLEEP_B_M1033_g N_SLEEP_B_c_1685_n N_SLEEP_B_c_1686_n
+ N_SLEEP_B_c_1687_n SLEEP_B N_SLEEP_B_c_1688_n N_SLEEP_B_c_1689_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%SLEEP_B
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%CLK N_CLK_M1015_g N_CLK_M1013_g CLK CLK CLK
+ N_CLK_c_1750_n PM_SKY130_FD_SC_LP__SRSDFXTP_1%CLK
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_2504_57# N_A_2504_57#_M1032_s
+ N_A_2504_57#_M1011_s N_A_2504_57#_M1031_g N_A_2504_57#_M1024_g
+ N_A_2504_57#_c_1799_n N_A_2504_57#_c_1804_n N_A_2504_57#_c_1800_n
+ N_A_2504_57#_c_1801_n N_A_2504_57#_c_1802_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_2504_57#
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%VPWR N_VPWR_M1030_d N_VPWR_M1039_d
+ N_VPWR_M1036_d N_VPWR_M1011_d N_VPWR_c_1855_n N_VPWR_c_1856_n N_VPWR_c_1857_n
+ N_VPWR_c_1858_n VPWR N_VPWR_c_1859_n N_VPWR_c_1860_n N_VPWR_c_1861_n
+ N_VPWR_c_1862_n N_VPWR_c_1854_n N_VPWR_c_1864_n N_VPWR_c_1865_n
+ N_VPWR_c_1866_n N_VPWR_c_1867_n VPWR PM_SKY130_FD_SC_LP__SRSDFXTP_1%VPWR
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_282_477# N_A_282_477#_M1003_d
+ N_A_282_477#_M1005_s N_A_282_477#_M1021_d N_A_282_477#_M1035_s
+ N_A_282_477#_c_2003_n N_A_282_477#_c_2004_n N_A_282_477#_c_2005_n
+ N_A_282_477#_c_1995_n N_A_282_477#_c_1996_n N_A_282_477#_c_1997_n
+ N_A_282_477#_c_1998_n N_A_282_477#_c_1999_n N_A_282_477#_c_2053_n
+ N_A_282_477#_c_2007_n N_A_282_477#_c_2008_n N_A_282_477#_c_2000_n
+ N_A_282_477#_c_2010_n N_A_282_477#_c_2011_n N_A_282_477#_c_2012_n
+ N_A_282_477#_c_2001_n N_A_282_477#_c_2013_n N_A_282_477#_c_2002_n
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_282_477#
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%KAPWR N_KAPWR_M1017_d N_KAPWR_M1015_d KAPWR
+ N_KAPWR_c_2176_n N_KAPWR_c_2214_n N_KAPWR_c_2164_n KAPWR
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%KAPWR
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%Q N_Q_M1031_d N_Q_M1024_d N_Q_c_2286_n
+ N_Q_c_2287_n N_Q_c_2283_n Q Q N_Q_c_2285_n Q PM_SKY130_FD_SC_LP__SRSDFXTP_1%Q
x_PM_SKY130_FD_SC_LP__SRSDFXTP_1%VGND N_VGND_M1040_d N_VGND_M1016_d
+ N_VGND_M1034_d N_VGND_M1006_d N_VGND_M1033_d N_VGND_M1032_d N_VGND_c_2305_n
+ N_VGND_c_2306_n N_VGND_c_2307_n N_VGND_c_2308_n N_VGND_c_2309_n
+ N_VGND_c_2310_n N_VGND_c_2311_n N_VGND_c_2312_n N_VGND_c_2313_n
+ N_VGND_c_2314_n VGND N_VGND_c_2315_n N_VGND_c_2316_n N_VGND_c_2317_n
+ N_VGND_c_2318_n N_VGND_c_2319_n N_VGND_c_2320_n N_VGND_c_2321_n
+ N_VGND_c_2322_n N_VGND_c_2323_n N_VGND_c_2324_n VGND
+ PM_SKY130_FD_SC_LP__SRSDFXTP_1%VGND
cc_1 VNB N_SCE_c_292_n 0.0210431f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=2.125
cc_2 VNB N_SCE_M1040_g 0.0312114f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_3 VNB N_SCE_M1018_g 0.0393518f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=0.445
cc_4 VNB N_SCE_c_295_n 0.0222231f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.925
cc_5 VNB N_SCE_c_296_n 0.00189563f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.18
cc_6 VNB N_SCE_c_297_n 0.00938349f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.925
cc_7 VNB SCE 0.00709151f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_8 VNB N_SCE_c_299_n 0.04845f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.15
cc_9 VNB N_SCE_c_300_n 0.0343409f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.345
cc_10 VNB N_A_31_477#_M1037_g 0.0564082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_31_477#_c_395_n 0.0376644f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=0.445
cc_12 VNB N_A_31_477#_c_396_n 0.0204683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_31_477#_c_397_n 0.00367141f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.15
cc_14 VNB N_A_31_477#_c_398_n 0.0156424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_D_M1021_g 0.0114233f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.275
cc_16 VNB N_D_M1003_g 0.0386033f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_17 VNB N_D_c_487_n 0.0272535f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.275
cc_18 VNB N_D_c_488_n 0.00862439f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.705
cc_19 VNB N_SCD_M1016_g 0.0186162f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_20 VNB N_SCD_c_522_n 0.0159206f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.705
cc_21 VNB N_SCD_c_523_n 0.0420279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_570_47#_c_576_n 0.0545682f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_23 VNB N_A_570_47#_M1008_g 0.0327453f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.705
cc_24 VNB N_A_570_47#_c_578_n 0.0168531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_570_47#_c_579_n 0.0187475f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.2
cc_26 VNB N_A_570_47#_c_580_n 0.0122224f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_27 VNB N_A_570_47#_c_581_n 0.0132004f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.18
cc_28 VNB N_A_570_47#_c_582_n 0.00647552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_570_47#_c_583_n 0.0011449f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.345
cc_30 VNB N_A_570_47#_c_584_n 7.74266e-19 $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.345
cc_31 VNB N_A_570_47#_c_585_n 0.00336493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_570_47#_c_586_n 0.00189785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_570_47#_c_587_n 7.4479e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_570_47#_c_588_n 0.0170028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_570_47#_c_589_n 0.0040802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_570_47#_c_590_n 0.0328433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_570_47#_c_591_n 0.00376571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_570_47#_c_592_n 0.0029799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_570_47#_c_593_n 0.0264806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_570_47#_c_594_n 0.00369179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_570_47#_c_595_n 0.00306848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_570_47#_c_596_n 0.00262135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_570_47#_c_597_n 9.82756e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_570_47#_c_598_n 0.00226055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_570_47#_c_599_n 0.0530515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_570_47#_c_600_n 0.0566532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_914_245#_c_823_n 0.00424104f $X=-0.19 $Y=-0.245 $X2=1.905
+ $Y2=0.445
cc_48 VNB N_A_914_245#_c_824_n 0.0358987f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=0.445
cc_49 VNB N_A_914_245#_c_825_n 0.00570298f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=2.2
cc_50 VNB N_A_914_245#_c_826_n 0.0150563f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.925
cc_51 VNB N_A_914_245#_c_827_n 0.00108377f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.15
cc_52 VNB N_A_914_245#_c_828_n 0.0174795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_786_139#_M1038_g 0.0309975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_786_139#_c_926_n 0.0136982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_786_139#_c_927_n 0.00297481f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_56 VNB N_A_786_139#_c_928_n 0.042428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_540_21#_M1025_g 0.0225807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_540_21#_c_1069_n 0.0458704f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.275
cc_59 VNB N_A_540_21#_M1005_g 0.0482494f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.2
cc_60 VNB N_A_540_21#_c_1071_n 0.0160682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_540_21#_c_1072_n 0.0108116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_540_21#_M1026_g 0.0561044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_540_21#_c_1074_n 0.0203704f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.345
cc_64 VNB N_A_540_21#_c_1075_n 0.0241542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_540_21#_c_1076_n 0.00843425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_540_21#_c_1077_n 0.00860914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_540_21#_c_1078_n 0.00126411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_540_21#_c_1079_n 8.45852e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_540_21#_c_1080_n 0.00263872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_540_21#_c_1081_n 0.00729321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_540_21#_c_1082_n 0.00888978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1319_69#_M1020_g 0.0201106f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.275
cc_73 VNB N_A_1319_69#_M1007_g 0.0210191f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=0.445
cc_74 VNB N_A_1319_69#_c_1314_n 0.0155231f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.18
cc_75 VNB N_A_1319_69#_c_1315_n 0.0309008f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.15
cc_76 VNB N_A_1319_69#_M1032_g 0.0285287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1319_69#_c_1317_n 0.0251141f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.18
cc_78 VNB N_A_1319_69#_c_1318_n 0.0120632f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.345
cc_79 VNB N_A_1319_69#_c_1319_n 0.0121646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1319_69#_c_1320_n 0.00307899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1319_69#_c_1321_n 0.00465671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1319_69#_c_1322_n 0.00145347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1319_69#_c_1323_n 0.0207932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1319_69#_c_1324_n 0.0139923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1319_69#_c_1325_n 0.0221316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1493_21#_M1019_g 0.0221392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1493_21#_c_1529_n 0.0112394f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.2
cc_88 VNB N_A_1493_21#_c_1530_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.275
cc_89 VNB N_A_1493_21#_M1006_g 0.0270989f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.18
cc_90 VNB N_A_1493_21#_c_1532_n 0.116729f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=0.445
cc_91 VNB N_A_1493_21#_c_1533_n 0.0394147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1493_21#_c_1534_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=0.59
+ $Y2=0.925
cc_93 VNB N_A_1493_21#_c_1535_n 0.030503f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.15
cc_94 VNB N_A_1493_21#_c_1536_n 0.00544618f $X=-0.19 $Y=-0.245 $X2=2.075
+ $Y2=1.21
cc_95 VNB N_A_1493_21#_c_1537_n 0.0178664f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.15
cc_96 VNB N_A_1493_21#_c_1538_n 0.00307732f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.15
cc_97 VNB N_A_1493_21#_c_1539_n 0.00509066f $X=-0.19 $Y=-0.245 $X2=1.965
+ $Y2=1.345
cc_98 VNB N_A_1493_21#_c_1540_n 0.00541257f $X=-0.19 $Y=-0.245 $X2=2.16
+ $Y2=1.345
cc_99 VNB N_A_1493_21#_c_1541_n 0.00278572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1493_21#_c_1542_n 0.0118341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1493_21#_c_1543_n 0.00580002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1493_21#_c_1544_n 0.00393584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1493_21#_c_1545_n 0.052763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_SLEEP_B_M1010_g 0.0695713f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.275
cc_105 VNB N_SLEEP_B_M1002_g 0.0198397f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_106 VNB N_SLEEP_B_c_1684_n 0.0336704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_SLEEP_B_c_1685_n 0.057206f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.275
cc_108 VNB N_SLEEP_B_c_1686_n 0.0239567f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.705
cc_109 VNB N_SLEEP_B_c_1687_n 0.00385799f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=2.2
cc_110 VNB N_SLEEP_B_c_1688_n 0.0544928f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.15
cc_111 VNB N_SLEEP_B_c_1689_n 0.00429603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_CLK_M1013_g 0.021129f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_113 VNB CLK 0.0146227f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.2
cc_114 VNB N_CLK_c_1750_n 0.034138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2504_57#_M1031_g 0.0273065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2504_57#_M1024_g 5.51802e-19 $X=-0.19 $Y=-0.245 $X2=0.945
+ $Y2=2.705
cc_117 VNB N_A_2504_57#_c_1799_n 0.0134666f $X=-0.19 $Y=-0.245 $X2=1.905
+ $Y2=0.445
cc_118 VNB N_A_2504_57#_c_1800_n 0.00931953f $X=-0.19 $Y=-0.245 $X2=1.88
+ $Y2=1.18
cc_119 VNB N_A_2504_57#_c_1801_n 0.0353509f $X=-0.19 $Y=-0.245 $X2=0.59
+ $Y2=0.925
cc_120 VNB N_A_2504_57#_c_1802_n 0.00424566f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.15
cc_121 VNB N_VPWR_c_1854_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_282_477#_c_1995_n 0.00162906f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=2.2
cc_123 VNB N_A_282_477#_c_1996_n 0.00159669f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=0.925
cc_124 VNB N_A_282_477#_c_1997_n 0.015501f $X=-0.19 $Y=-0.245 $X2=0.755
+ $Y2=0.925
cc_125 VNB N_A_282_477#_c_1998_n 0.00350631f $X=-0.19 $Y=-0.245 $X2=1.88
+ $Y2=1.01
cc_126 VNB N_A_282_477#_c_1999_n 0.00948639f $X=-0.19 $Y=-0.245 $X2=0.59
+ $Y2=0.925
cc_127 VNB N_A_282_477#_c_2000_n 0.00563468f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.15
cc_128 VNB N_A_282_477#_c_2001_n 0.00281813f $X=-0.19 $Y=-0.245 $X2=1.965
+ $Y2=1.18
cc_129 VNB N_A_282_477#_c_2002_n 0.00626963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_Q_c_2283_n 0.0239803f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.18
cc_131 VNB Q 0.00968796f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=0.445
cc_132 VNB N_Q_c_2285_n 0.0301489f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.925
cc_133 VNB N_VGND_c_2305_n 0.00292296f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.2
cc_134 VNB N_VGND_c_2306_n 0.00645063f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.18
cc_135 VNB N_VGND_c_2307_n 0.00509157f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.15
cc_136 VNB N_VGND_c_2308_n 0.0113677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2309_n 0.0291661f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.345
cc_138 VNB N_VGND_c_2310_n 0.0117347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2311_n 0.0658628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2312_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2313_n 0.0950052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2314_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2315_n 0.0169287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2316_n 0.0423732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2317_n 0.0506272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2318_n 0.0215724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2319_n 0.0187292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2320_n 0.69255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2321_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2322_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2323_n 0.00477645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2324_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VPB N_SCE_c_292_n 0.02898f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=2.125
cc_154 VPB N_SCE_c_302_n 0.0192508f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.275
cc_155 VPB N_SCE_c_303_n 0.0193814f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=2.2
cc_156 VPB N_SCE_c_304_n 0.0238031f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.2
cc_157 VPB N_SCE_c_305_n 0.0160737f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.275
cc_158 VPB N_A_31_477#_M1004_g 0.0276108f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.705
cc_159 VPB N_A_31_477#_c_395_n 0.00872581f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=0.445
cc_160 VPB N_A_31_477#_c_401_n 0.0357216f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=2.2
cc_161 VPB N_A_31_477#_c_402_n 0.00384212f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.2
cc_162 VPB N_A_31_477#_c_403_n 0.0131888f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.18
cc_163 VPB N_A_31_477#_c_404_n 0.0370933f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.925
cc_164 VPB N_A_31_477#_c_405_n 0.00725125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_31_477#_c_397_n 0.0032515f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.15
cc_166 VPB N_A_31_477#_c_398_n 0.0243048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_D_M1021_g 0.051181f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.275
cc_168 VPB N_SCD_M1039_g 0.0316118f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.275
cc_169 VPB N_SCD_c_525_n 0.0329217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_SCD_c_526_n 0.00858753f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=2.2
cc_171 VPB N_SCD_c_523_n 0.00809944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_570_47#_c_601_n 0.0382222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_570_47#_c_602_n 0.0193343f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=1.18
cc_174 VPB N_A_570_47#_c_603_n 0.0266616f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.01
cc_175 VPB N_A_570_47#_c_604_n 0.0186626f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.15
cc_176 VPB N_A_570_47#_c_580_n 0.00206664f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_177 VPB N_A_570_47#_c_606_n 0.0077635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_570_47#_c_607_n 0.00686414f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.15
cc_179 VPB N_A_570_47#_c_608_n 0.0036057f $X=-0.19 $Y=1.655 $X2=1.965 $Y2=1.345
cc_180 VPB N_A_570_47#_c_592_n 0.0016339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_570_47#_c_593_n 0.00904295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_570_47#_c_611_n 0.0422456f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_914_245#_M1036_g 0.0252042f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.275
cc_184 VPB N_A_914_245#_c_826_n 0.00804486f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.925
cc_185 VPB N_A_914_245#_c_831_n 0.00787591f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.15
cc_186 VPB N_A_914_245#_c_832_n 0.00718553f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.15
cc_187 VPB N_A_914_245#_c_833_n 0.0307184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_914_245#_c_834_n 0.0015828f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.15
cc_189 VPB N_A_786_139#_c_929_n 0.0187075f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.2
cc_190 VPB N_A_786_139#_c_930_n 0.112253f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.705
cc_191 VPB N_A_786_139#_c_931_n 0.0125556f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=1.18
cc_192 VPB N_A_786_139#_c_926_n 0.00289447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_786_139#_c_933_n 0.00894875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_786_139#_c_934_n 4.51508e-19 $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.2
cc_195 VPB N_A_786_139#_c_935_n 0.00766971f $X=-0.19 $Y=1.655 $X2=0.755
+ $Y2=0.925
cc_196 VPB N_A_786_139#_c_936_n 0.00341444f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.01
cc_197 VPB N_A_786_139#_c_937_n 0.00743144f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.925
cc_198 VPB N_A_786_139#_c_927_n 0.0030345f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_199 VPB N_A_786_139#_c_939_n 0.0280714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_786_139#_c_940_n 0.00227271f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.15
cc_201 VPB N_A_786_139#_c_941_n 0.00203831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_786_139#_c_942_n 0.00232242f $X=-0.19 $Y=1.655 $X2=1.965 $Y2=1.18
cc_203 VPB N_A_786_139#_c_943_n 0.00185984f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.345
cc_204 VPB N_A_786_139#_c_944_n 0.0588424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_540_21#_c_1069_n 0.00736582f $X=-0.19 $Y=1.655 $X2=0.945
+ $Y2=2.275
cc_206 VPB N_A_540_21#_M1027_g 0.0458011f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=1.18
cc_207 VPB N_A_540_21#_c_1085_n 0.0457685f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=0.445
cc_208 VPB N_A_540_21#_M1005_g 0.00717563f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.2
cc_209 VPB N_A_540_21#_c_1087_n 0.061951f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=0.925
cc_210 VPB N_A_540_21#_M1022_g 0.0519588f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.15
cc_211 VPB N_A_540_21#_c_1089_n 0.0437178f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.15
cc_212 VPB N_A_540_21#_c_1071_n 0.0291027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_540_21#_c_1091_n 0.0156452f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_540_21#_c_1072_n 0.00428232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_540_21#_c_1093_n 0.0157831f $X=-0.19 $Y=1.655 $X2=1.965 $Y2=1.345
cc_216 VPB N_A_540_21#_c_1074_n 0.0275136f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.345
cc_217 VPB N_A_540_21#_c_1095_n 0.011188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_540_21#_c_1096_n 0.00819645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_540_21#_c_1097_n 0.0066402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_540_21#_c_1076_n 0.0208168f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_540_21#_c_1077_n 0.00206952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_540_21#_c_1078_n 0.0025524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_540_21#_c_1101_n 0.00942507f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_540_21#_c_1102_n 5.73999e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_540_21#_c_1103_n 0.00379214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_540_21#_c_1080_n 0.00640376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_540_21#_c_1105_n 0.00240085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_540_21#_c_1106_n 0.0156086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_540_21#_c_1107_n 0.00191138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_540_21#_c_1108_n 0.00212087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_540_21#_c_1082_n 0.0470816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_1319_69#_c_1326_n 0.0285043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_1319_69#_c_1327_n 0.0391384f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.2
cc_234 VPB N_A_1319_69#_c_1328_n 0.0143848f $X=-0.19 $Y=1.655 $X2=1.795
+ $Y2=0.925
cc_235 VPB N_A_1319_69#_c_1314_n 0.00867384f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.18
cc_236 VPB N_A_1319_69#_c_1330_n 0.0192854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_1319_69#_c_1318_n 0.0164372f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.345
cc_238 VPB N_A_1319_69#_c_1320_n 0.00304032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_1319_69#_c_1322_n 0.00980781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_1319_69#_c_1334_n 0.0294176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_1319_69#_c_1335_n 0.0109185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_1319_69#_c_1336_n 0.00146649f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1319_69#_c_1337_n 0.0125266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_1319_69#_c_1338_n 0.00245458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_1319_69#_c_1339_n 0.00146721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_1319_69#_c_1340_n 0.00633646f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_1319_69#_c_1341_n 0.0425817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_1319_69#_c_1342_n 0.00304223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_1319_69#_c_1325_n 0.016201f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_1319_69#_c_1344_n 0.0134962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_1319_69#_c_1345_n 0.0498361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_1493_21#_c_1546_n 0.0309102f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.2
cc_253 VPB N_A_1493_21#_c_1535_n 0.0177311f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.15
cc_254 VPB N_A_1493_21#_c_1539_n 0.0039452f $X=-0.19 $Y=1.655 $X2=1.965
+ $Y2=1.345
cc_255 VPB N_A_1493_21#_c_1549_n 0.00822917f $X=-0.19 $Y=1.655 $X2=1.965
+ $Y2=1.345
cc_256 VPB N_A_1493_21#_c_1550_n 0.00375433f $X=-0.19 $Y=1.655 $X2=1.88
+ $Y2=1.345
cc_257 VPB N_SLEEP_B_M1010_g 0.0365723f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.275
cc_258 VPB N_CLK_M1015_g 0.0276406f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.275
cc_259 VPB CLK 0.00719151f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.2
cc_260 VPB N_CLK_c_1750_n 0.0182137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_2504_57#_M1024_g 0.028321f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.705
cc_262 VPB N_A_2504_57#_c_1804_n 0.0103767f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.2
cc_263 VPB N_VPWR_c_1855_n 0.00455795f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=1.18
cc_264 VPB N_VPWR_c_1856_n 0.0071139f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=2.2
cc_265 VPB N_VPWR_c_1857_n 0.0688491f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.2
cc_266 VPB N_VPWR_c_1858_n 0.0142964f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.18
cc_267 VPB N_VPWR_c_1859_n 0.0168929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1860_n 0.0443325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1861_n 0.180517f $X=-0.19 $Y=1.655 $X2=1.965 $Y2=1.345
cc_270 VPB N_VPWR_c_1862_n 0.0185366f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1854_n 0.0759527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1864_n 0.00522307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1865_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1866_n 0.00981695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1867_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_282_477#_c_2003_n 0.00214822f $X=-0.19 $Y=1.655 $X2=1.905
+ $Y2=1.18
cc_277 VPB N_A_282_477#_c_2004_n 0.0133078f $X=-0.19 $Y=1.655 $X2=1.905
+ $Y2=0.445
cc_278 VPB N_A_282_477#_c_2005_n 0.00273691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_282_477#_c_1999_n 0.0136606f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.925
cc_280 VPB N_A_282_477#_c_2007_n 0.0166962f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.15
cc_281 VPB N_A_282_477#_c_2008_n 0.00158776f $X=-0.19 $Y=1.655 $X2=2.075
+ $Y2=1.21
cc_282 VPB N_A_282_477#_c_2000_n 0.00638063f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.15
cc_283 VPB N_A_282_477#_c_2010_n 0.0101995f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_282_477#_c_2011_n 0.00279403f $X=-0.19 $Y=1.655 $X2=0.525
+ $Y2=1.15
cc_285 VPB N_A_282_477#_c_2012_n 0.00758253f $X=-0.19 $Y=1.655 $X2=1.965
+ $Y2=1.345
cc_286 VPB N_A_282_477#_c_2013_n 0.00510526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_287 VPB N_KAPWR_c_2164_n 0.0591554f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=0.445
cc_288 VPB N_Q_c_2286_n 0.0362634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_289 VPB N_Q_c_2287_n 0.00968796f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.705
cc_290 VPB N_Q_c_2283_n 0.00773243f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=1.18
cc_291 N_SCE_c_292_n N_A_31_477#_M1037_g 0.00335311f $X=0.27 $Y=2.125 $X2=0
+ $Y2=0
cc_292 N_SCE_M1040_g N_A_31_477#_M1037_g 0.0224982f $X=0.545 $Y=0.445 $X2=0
+ $Y2=0
cc_293 N_SCE_c_295_n N_A_31_477#_M1037_g 0.0157143f $X=1.795 $Y=0.925 $X2=0
+ $Y2=0
cc_294 N_SCE_c_297_n N_A_31_477#_M1037_g 0.00503559f $X=0.59 $Y=0.925 $X2=0
+ $Y2=0
cc_295 N_SCE_c_299_n N_A_31_477#_M1037_g 0.0196323f $X=0.545 $Y=1.15 $X2=0 $Y2=0
cc_296 N_SCE_c_292_n N_A_31_477#_c_395_n 0.0213672f $X=0.27 $Y=2.125 $X2=0 $Y2=0
cc_297 N_SCE_M1040_g N_A_31_477#_c_395_n 0.00822873f $X=0.545 $Y=0.445 $X2=0
+ $Y2=0
cc_298 N_SCE_c_297_n N_A_31_477#_c_395_n 0.0308074f $X=0.59 $Y=0.925 $X2=0 $Y2=0
cc_299 N_SCE_c_299_n N_A_31_477#_c_395_n 0.0128393f $X=0.545 $Y=1.15 $X2=0 $Y2=0
cc_300 N_SCE_c_292_n N_A_31_477#_c_401_n 0.00131479f $X=0.27 $Y=2.125 $X2=0
+ $Y2=0
cc_301 N_SCE_c_302_n N_A_31_477#_c_401_n 0.00497446f $X=0.515 $Y=2.275 $X2=0
+ $Y2=0
cc_302 N_SCE_c_304_n N_A_31_477#_c_401_n 0.0173908f $X=0.59 $Y=2.2 $X2=0 $Y2=0
cc_303 N_SCE_c_304_n N_A_31_477#_c_402_n 0.00874435f $X=0.59 $Y=2.2 $X2=0 $Y2=0
cc_304 N_SCE_c_297_n N_A_31_477#_c_402_n 0.00466007f $X=0.59 $Y=0.925 $X2=0
+ $Y2=0
cc_305 N_SCE_c_299_n N_A_31_477#_c_402_n 0.00176494f $X=0.545 $Y=1.15 $X2=0
+ $Y2=0
cc_306 N_SCE_c_303_n N_A_31_477#_c_403_n 0.00299361f $X=0.87 $Y=2.2 $X2=0 $Y2=0
cc_307 SCE N_A_31_477#_c_403_n 0.00628791f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_308 N_SCE_c_300_n N_A_31_477#_c_403_n 4.30942e-19 $X=1.965 $Y=1.345 $X2=0
+ $Y2=0
cc_309 SCE N_A_31_477#_c_404_n 8.51686e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_310 N_SCE_c_300_n N_A_31_477#_c_404_n 0.00863897f $X=1.965 $Y=1.345 $X2=0
+ $Y2=0
cc_311 N_SCE_M1040_g N_A_31_477#_c_396_n 7.72299e-19 $X=0.545 $Y=0.445 $X2=0
+ $Y2=0
cc_312 N_SCE_c_299_n N_A_31_477#_c_396_n 0.00626563f $X=0.545 $Y=1.15 $X2=0
+ $Y2=0
cc_313 N_SCE_c_292_n N_A_31_477#_c_405_n 0.0122461f $X=0.27 $Y=2.125 $X2=0 $Y2=0
cc_314 N_SCE_c_299_n N_A_31_477#_c_405_n 0.00114318f $X=0.545 $Y=1.15 $X2=0
+ $Y2=0
cc_315 N_SCE_c_292_n N_A_31_477#_c_397_n 0.00213587f $X=0.27 $Y=2.125 $X2=0
+ $Y2=0
cc_316 N_SCE_c_304_n N_A_31_477#_c_397_n 0.00389783f $X=0.59 $Y=2.2 $X2=0 $Y2=0
cc_317 N_SCE_c_295_n N_A_31_477#_c_397_n 0.00506983f $X=1.795 $Y=0.925 $X2=0
+ $Y2=0
cc_318 N_SCE_c_297_n N_A_31_477#_c_397_n 0.0106222f $X=0.59 $Y=0.925 $X2=0 $Y2=0
cc_319 N_SCE_c_292_n N_A_31_477#_c_398_n 0.0169297f $X=0.27 $Y=2.125 $X2=0 $Y2=0
cc_320 N_SCE_c_304_n N_A_31_477#_c_398_n 0.0233393f $X=0.59 $Y=2.2 $X2=0 $Y2=0
cc_321 N_SCE_c_295_n N_A_31_477#_c_398_n 7.61156e-19 $X=1.795 $Y=0.925 $X2=0
+ $Y2=0
cc_322 N_SCE_c_297_n N_A_31_477#_c_398_n 6.04465e-19 $X=0.59 $Y=0.925 $X2=0
+ $Y2=0
cc_323 N_SCE_c_299_n N_A_31_477#_c_398_n 0.00578856f $X=0.545 $Y=1.15 $X2=0
+ $Y2=0
cc_324 N_SCE_c_303_n N_D_M1021_g 0.0572147f $X=0.87 $Y=2.2 $X2=0 $Y2=0
cc_325 N_SCE_M1018_g N_D_M1003_g 0.0251845f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_326 N_SCE_c_295_n N_D_M1003_g 0.0122719f $X=1.795 $Y=0.925 $X2=0 $Y2=0
cc_327 N_SCE_c_296_n N_D_M1003_g 0.00294382f $X=1.88 $Y=1.18 $X2=0 $Y2=0
cc_328 N_SCE_c_295_n N_D_c_487_n 0.0041539f $X=1.795 $Y=0.925 $X2=0 $Y2=0
cc_329 SCE N_D_c_487_n 0.001218f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_330 N_SCE_c_300_n N_D_c_487_n 0.0214313f $X=1.965 $Y=1.345 $X2=0 $Y2=0
cc_331 N_SCE_c_295_n N_D_c_488_n 0.038115f $X=1.795 $Y=0.925 $X2=0 $Y2=0
cc_332 N_SCE_c_297_n N_D_c_488_n 0.00729781f $X=0.59 $Y=0.925 $X2=0 $Y2=0
cc_333 SCE N_D_c_488_n 0.0241648f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_334 N_SCE_c_300_n N_D_c_488_n 4.0822e-19 $X=1.965 $Y=1.345 $X2=0 $Y2=0
cc_335 N_SCE_M1018_g N_SCD_M1016_g 0.0452059f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_336 SCE N_SCD_c_522_n 3.60445e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_337 SCE N_SCD_c_525_n 0.00292945f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_338 SCE N_SCD_c_526_n 0.0125477f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_339 N_SCE_c_300_n N_SCD_c_526_n 0.00120763f $X=1.965 $Y=1.345 $X2=0 $Y2=0
cc_340 N_SCE_M1018_g N_SCD_c_523_n 0.00609308f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_341 N_SCE_c_296_n N_SCD_c_523_n 6.28027e-19 $X=1.88 $Y=1.18 $X2=0 $Y2=0
cc_342 SCE N_SCD_c_523_n 0.00337699f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_343 N_SCE_c_300_n N_SCD_c_523_n 0.0193196f $X=1.965 $Y=1.345 $X2=0 $Y2=0
cc_344 N_SCE_c_302_n N_VPWR_c_1855_n 0.0121238f $X=0.515 $Y=2.275 $X2=0 $Y2=0
cc_345 N_SCE_c_303_n N_VPWR_c_1855_n 0.00241555f $X=0.87 $Y=2.2 $X2=0 $Y2=0
cc_346 N_SCE_c_305_n N_VPWR_c_1855_n 0.014904f $X=0.945 $Y=2.275 $X2=0 $Y2=0
cc_347 N_SCE_c_302_n N_VPWR_c_1859_n 0.00429645f $X=0.515 $Y=2.275 $X2=0 $Y2=0
cc_348 N_SCE_c_305_n N_VPWR_c_1860_n 0.00429645f $X=0.945 $Y=2.275 $X2=0 $Y2=0
cc_349 N_SCE_c_302_n N_VPWR_c_1854_n 0.00382156f $X=0.515 $Y=2.275 $X2=0 $Y2=0
cc_350 N_SCE_c_305_n N_VPWR_c_1854_n 0.00325954f $X=0.945 $Y=2.275 $X2=0 $Y2=0
cc_351 N_SCE_c_305_n N_A_282_477#_c_2003_n 0.00168748f $X=0.945 $Y=2.275 $X2=0
+ $Y2=0
cc_352 N_SCE_c_305_n N_A_282_477#_c_2005_n 5.73298e-19 $X=0.945 $Y=2.275 $X2=0
+ $Y2=0
cc_353 N_SCE_M1018_g N_A_282_477#_c_1995_n 0.00838471f $X=1.905 $Y=0.445 $X2=0
+ $Y2=0
cc_354 N_SCE_c_295_n N_A_282_477#_c_1995_n 0.00771488f $X=1.795 $Y=0.925 $X2=0
+ $Y2=0
cc_355 SCE N_A_282_477#_c_1995_n 0.00555289f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_356 N_SCE_c_300_n N_A_282_477#_c_1995_n 0.00260007f $X=1.965 $Y=1.345 $X2=0
+ $Y2=0
cc_357 N_SCE_M1018_g N_A_282_477#_c_1996_n 0.00346967f $X=1.905 $Y=0.445 $X2=0
+ $Y2=0
cc_358 N_SCE_M1018_g N_A_282_477#_c_1997_n 4.88897e-19 $X=1.905 $Y=0.445 $X2=0
+ $Y2=0
cc_359 N_SCE_c_296_n N_A_282_477#_c_1997_n 0.00486623f $X=1.88 $Y=1.18 $X2=0
+ $Y2=0
cc_360 N_SCE_M1018_g N_A_282_477#_c_1998_n 0.00105478f $X=1.905 $Y=0.445 $X2=0
+ $Y2=0
cc_361 N_SCE_c_295_n N_A_282_477#_c_1998_n 0.0148412f $X=1.795 $Y=0.925 $X2=0
+ $Y2=0
cc_362 SCE N_A_282_477#_c_1998_n 0.0121074f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_363 SCE N_A_282_477#_c_1999_n 0.0152008f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_364 N_SCE_M1018_g N_A_282_477#_c_2001_n 0.0062834f $X=1.905 $Y=0.445 $X2=0
+ $Y2=0
cc_365 N_SCE_c_295_n N_A_282_477#_c_2001_n 0.0260342f $X=1.795 $Y=0.925 $X2=0
+ $Y2=0
cc_366 N_SCE_c_302_n N_KAPWR_c_2164_n 0.00250617f $X=0.515 $Y=2.275 $X2=0 $Y2=0
cc_367 N_SCE_c_304_n N_KAPWR_c_2164_n 0.00111799f $X=0.59 $Y=2.2 $X2=0 $Y2=0
cc_368 N_SCE_c_305_n N_KAPWR_c_2164_n 0.00432201f $X=0.945 $Y=2.275 $X2=0 $Y2=0
cc_369 N_SCE_M1040_g N_VGND_c_2305_n 0.010828f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_370 N_SCE_c_295_n N_VGND_c_2305_n 0.0137312f $X=1.795 $Y=0.925 $X2=0 $Y2=0
cc_371 N_SCE_c_297_n N_VGND_c_2305_n 0.0139591f $X=0.59 $Y=0.925 $X2=0 $Y2=0
cc_372 N_SCE_c_299_n N_VGND_c_2305_n 3.90443e-19 $X=0.545 $Y=1.15 $X2=0 $Y2=0
cc_373 N_SCE_M1040_g N_VGND_c_2315_n 0.00486043f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_374 N_SCE_M1018_g N_VGND_c_2316_n 0.00397678f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_375 N_SCE_M1040_g N_VGND_c_2320_n 0.00909748f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_376 N_SCE_M1018_g N_VGND_c_2320_n 0.00586794f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_377 N_SCE_c_295_n N_VGND_c_2320_n 0.019992f $X=1.795 $Y=0.925 $X2=0 $Y2=0
cc_378 N_SCE_c_297_n N_VGND_c_2320_n 8.86269e-19 $X=0.59 $Y=0.925 $X2=0 $Y2=0
cc_379 N_A_31_477#_M1004_g N_D_M1021_g 0.0213394f $X=1.765 $Y=2.705 $X2=0 $Y2=0
cc_380 N_A_31_477#_c_403_n N_D_M1021_g 0.018994f $X=1.785 $Y=1.915 $X2=0 $Y2=0
cc_381 N_A_31_477#_c_404_n N_D_M1021_g 0.0213351f $X=1.785 $Y=1.915 $X2=0 $Y2=0
cc_382 N_A_31_477#_c_397_n N_D_M1021_g 0.00162817f $X=0.75 $Y=1.72 $X2=0 $Y2=0
cc_383 N_A_31_477#_c_398_n N_D_M1021_g 0.0220531f $X=0.975 $Y=1.72 $X2=0 $Y2=0
cc_384 N_A_31_477#_M1037_g N_D_M1003_g 0.0579731f $X=0.975 $Y=0.445 $X2=0 $Y2=0
cc_385 N_A_31_477#_M1037_g N_D_c_487_n 0.0220531f $X=0.975 $Y=0.445 $X2=0 $Y2=0
cc_386 N_A_31_477#_c_403_n N_D_c_487_n 0.00403704f $X=1.785 $Y=1.915 $X2=0 $Y2=0
cc_387 N_A_31_477#_M1037_g N_D_c_488_n 0.00702801f $X=0.975 $Y=0.445 $X2=0 $Y2=0
cc_388 N_A_31_477#_c_403_n N_D_c_488_n 0.0310183f $X=1.785 $Y=1.915 $X2=0 $Y2=0
cc_389 N_A_31_477#_M1004_g N_SCD_M1039_g 0.0437163f $X=1.765 $Y=2.705 $X2=0
+ $Y2=0
cc_390 N_A_31_477#_c_403_n N_SCD_c_525_n 3.18329e-19 $X=1.785 $Y=1.915 $X2=0
+ $Y2=0
cc_391 N_A_31_477#_c_404_n N_SCD_c_525_n 0.020513f $X=1.785 $Y=1.915 $X2=0 $Y2=0
cc_392 N_A_31_477#_M1004_g N_SCD_c_526_n 0.00159902f $X=1.765 $Y=2.705 $X2=0
+ $Y2=0
cc_393 N_A_31_477#_c_403_n N_SCD_c_526_n 0.0281419f $X=1.785 $Y=1.915 $X2=0
+ $Y2=0
cc_394 N_A_31_477#_c_404_n N_SCD_c_526_n 0.00209319f $X=1.785 $Y=1.915 $X2=0
+ $Y2=0
cc_395 N_A_31_477#_c_401_n N_VPWR_c_1855_n 0.029037f $X=0.3 $Y=2.53 $X2=0 $Y2=0
cc_396 N_A_31_477#_c_402_n N_VPWR_c_1855_n 9.4611e-19 $X=0.585 $Y=1.995 $X2=0
+ $Y2=0
cc_397 N_A_31_477#_c_397_n N_VPWR_c_1855_n 0.0179645f $X=0.75 $Y=1.72 $X2=0
+ $Y2=0
cc_398 N_A_31_477#_c_398_n N_VPWR_c_1855_n 6.03083e-19 $X=0.975 $Y=1.72 $X2=0
+ $Y2=0
cc_399 N_A_31_477#_c_401_n N_VPWR_c_1859_n 0.0179493f $X=0.3 $Y=2.53 $X2=0 $Y2=0
cc_400 N_A_31_477#_M1004_g N_VPWR_c_1860_n 0.00485697f $X=1.765 $Y=2.705 $X2=0
+ $Y2=0
cc_401 N_A_31_477#_M1004_g N_VPWR_c_1854_n 0.00439301f $X=1.765 $Y=2.705 $X2=0
+ $Y2=0
cc_402 N_A_31_477#_c_401_n N_VPWR_c_1854_n 0.00286516f $X=0.3 $Y=2.53 $X2=0
+ $Y2=0
cc_403 N_A_31_477#_M1004_g N_A_282_477#_c_2003_n 0.0115695f $X=1.765 $Y=2.705
+ $X2=0 $Y2=0
cc_404 N_A_31_477#_M1004_g N_A_282_477#_c_2004_n 0.00808955f $X=1.765 $Y=2.705
+ $X2=0 $Y2=0
cc_405 N_A_31_477#_c_403_n N_A_282_477#_c_2004_n 0.00988418f $X=1.785 $Y=1.915
+ $X2=0 $Y2=0
cc_406 N_A_31_477#_c_404_n N_A_282_477#_c_2004_n 0.00295814f $X=1.785 $Y=1.915
+ $X2=0 $Y2=0
cc_407 N_A_31_477#_M1004_g N_A_282_477#_c_2005_n 0.00157294f $X=1.765 $Y=2.705
+ $X2=0 $Y2=0
cc_408 N_A_31_477#_c_403_n N_A_282_477#_c_2005_n 0.0209631f $X=1.785 $Y=1.915
+ $X2=0 $Y2=0
cc_409 N_A_31_477#_c_404_n N_A_282_477#_c_2005_n 0.00157029f $X=1.785 $Y=1.915
+ $X2=0 $Y2=0
cc_410 N_A_31_477#_M1030_s N_KAPWR_c_2164_n 9.94816e-19 $X=0.155 $Y=2.385 $X2=0
+ $Y2=0
cc_411 N_A_31_477#_M1004_g N_KAPWR_c_2164_n 0.0041732f $X=1.765 $Y=2.705 $X2=0
+ $Y2=0
cc_412 N_A_31_477#_c_401_n N_KAPWR_c_2164_n 0.0306093f $X=0.3 $Y=2.53 $X2=0
+ $Y2=0
cc_413 N_A_31_477#_c_402_n N_KAPWR_c_2164_n 0.0054446f $X=0.585 $Y=1.995 $X2=0
+ $Y2=0
cc_414 N_A_31_477#_c_403_n N_KAPWR_c_2164_n 0.0166524f $X=1.785 $Y=1.915 $X2=0
+ $Y2=0
cc_415 N_A_31_477#_c_397_n N_KAPWR_c_2164_n 0.00210861f $X=0.75 $Y=1.72 $X2=0
+ $Y2=0
cc_416 N_A_31_477#_M1037_g N_VGND_c_2305_n 0.0136233f $X=0.975 $Y=0.445 $X2=0
+ $Y2=0
cc_417 N_A_31_477#_c_396_n N_VGND_c_2305_n 0.0154668f $X=0.33 $Y=0.465 $X2=0
+ $Y2=0
cc_418 N_A_31_477#_c_396_n N_VGND_c_2315_n 0.0223203f $X=0.33 $Y=0.465 $X2=0
+ $Y2=0
cc_419 N_A_31_477#_M1037_g N_VGND_c_2316_n 0.00486043f $X=0.975 $Y=0.445 $X2=0
+ $Y2=0
cc_420 N_A_31_477#_M1040_s N_VGND_c_2320_n 0.00424065f $X=0.185 $Y=0.235 $X2=0
+ $Y2=0
cc_421 N_A_31_477#_M1037_g N_VGND_c_2320_n 0.0045381f $X=0.975 $Y=0.445 $X2=0
+ $Y2=0
cc_422 N_A_31_477#_c_396_n N_VGND_c_2320_n 0.0126561f $X=0.33 $Y=0.465 $X2=0
+ $Y2=0
cc_423 N_D_M1021_g N_VPWR_c_1855_n 0.00280889f $X=1.335 $Y=2.705 $X2=0 $Y2=0
cc_424 N_D_M1021_g N_VPWR_c_1860_n 0.00485697f $X=1.335 $Y=2.705 $X2=0 $Y2=0
cc_425 N_D_M1021_g N_VPWR_c_1854_n 0.00449887f $X=1.335 $Y=2.705 $X2=0 $Y2=0
cc_426 N_D_M1021_g N_A_282_477#_c_2003_n 0.0084677f $X=1.335 $Y=2.705 $X2=0
+ $Y2=0
cc_427 N_D_M1021_g N_A_282_477#_c_2005_n 0.00412937f $X=1.335 $Y=2.705 $X2=0
+ $Y2=0
cc_428 N_D_M1003_g N_A_282_477#_c_2001_n 0.00589513f $X=1.365 $Y=0.445 $X2=0
+ $Y2=0
cc_429 N_D_M1021_g N_KAPWR_c_2164_n 0.00452956f $X=1.335 $Y=2.705 $X2=0 $Y2=0
cc_430 N_D_M1003_g N_VGND_c_2305_n 0.00242344f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_431 N_D_M1003_g N_VGND_c_2316_n 0.00585385f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_432 N_D_M1003_g N_VGND_c_2320_n 0.00674038f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_433 N_SCD_c_522_n N_A_570_47#_c_580_n 3.01975e-19 $X=2.415 $Y=0.895 $X2=0
+ $Y2=0
cc_434 N_SCD_M1016_g N_A_540_21#_M1025_g 0.0119424f $X=2.295 $Y=0.445 $X2=0
+ $Y2=0
cc_435 N_SCD_c_522_n N_A_540_21#_M1025_g 0.00479298f $X=2.415 $Y=0.895 $X2=0
+ $Y2=0
cc_436 N_SCD_c_523_n N_A_540_21#_c_1069_n 0.0102533f $X=2.325 $Y=1.75 $X2=0
+ $Y2=0
cc_437 N_SCD_M1039_g N_A_540_21#_M1027_g 0.0120268f $X=2.235 $Y=2.705 $X2=0
+ $Y2=0
cc_438 N_SCD_c_525_n N_A_540_21#_M1027_g 0.00293352f $X=2.325 $Y=1.915 $X2=0
+ $Y2=0
cc_439 N_SCD_c_523_n N_A_540_21#_c_1075_n 0.00479298f $X=2.325 $Y=1.75 $X2=0
+ $Y2=0
cc_440 N_SCD_c_525_n N_A_540_21#_c_1095_n 0.0102533f $X=2.325 $Y=1.915 $X2=0
+ $Y2=0
cc_441 N_SCD_M1039_g N_VPWR_c_1856_n 0.0124228f $X=2.235 $Y=2.705 $X2=0 $Y2=0
cc_442 N_SCD_M1039_g N_VPWR_c_1860_n 0.0051746f $X=2.235 $Y=2.705 $X2=0 $Y2=0
cc_443 N_SCD_M1039_g N_VPWR_c_1854_n 0.00480591f $X=2.235 $Y=2.705 $X2=0 $Y2=0
cc_444 N_SCD_M1039_g N_A_282_477#_c_2003_n 0.00333745f $X=2.235 $Y=2.705 $X2=0
+ $Y2=0
cc_445 N_SCD_M1039_g N_A_282_477#_c_2004_n 0.0123518f $X=2.235 $Y=2.705 $X2=0
+ $Y2=0
cc_446 N_SCD_c_525_n N_A_282_477#_c_2004_n 0.00104222f $X=2.325 $Y=1.915 $X2=0
+ $Y2=0
cc_447 N_SCD_c_526_n N_A_282_477#_c_2004_n 0.0311061f $X=2.325 $Y=1.915 $X2=0
+ $Y2=0
cc_448 N_SCD_M1016_g N_A_282_477#_c_1995_n 0.00572428f $X=2.295 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_SCD_M1016_g N_A_282_477#_c_1996_n 0.00400262f $X=2.295 $Y=0.445 $X2=0
+ $Y2=0
cc_450 N_SCD_c_522_n N_A_282_477#_c_1996_n 5.24801e-19 $X=2.415 $Y=0.895 $X2=0
+ $Y2=0
cc_451 N_SCD_c_522_n N_A_282_477#_c_1997_n 0.00723338f $X=2.415 $Y=0.895 $X2=0
+ $Y2=0
cc_452 N_SCD_c_523_n N_A_282_477#_c_1997_n 0.0129214f $X=2.325 $Y=1.75 $X2=0
+ $Y2=0
cc_453 N_SCD_c_522_n N_A_282_477#_c_1998_n 0.00290651f $X=2.415 $Y=0.895 $X2=0
+ $Y2=0
cc_454 N_SCD_M1039_g N_A_282_477#_c_1999_n 0.00351506f $X=2.235 $Y=2.705 $X2=0
+ $Y2=0
cc_455 N_SCD_c_525_n N_A_282_477#_c_1999_n 0.00120327f $X=2.325 $Y=1.915 $X2=0
+ $Y2=0
cc_456 N_SCD_c_526_n N_A_282_477#_c_1999_n 0.0308862f $X=2.325 $Y=1.915 $X2=0
+ $Y2=0
cc_457 N_SCD_c_523_n N_A_282_477#_c_1999_n 0.00834093f $X=2.325 $Y=1.75 $X2=0
+ $Y2=0
cc_458 N_SCD_M1039_g N_A_282_477#_c_2053_n 0.0029209f $X=2.235 $Y=2.705 $X2=0
+ $Y2=0
cc_459 N_SCD_M1016_g N_A_282_477#_c_2001_n 8.13465e-19 $X=2.295 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_SCD_M1039_g N_KAPWR_c_2164_n 0.00911148f $X=2.235 $Y=2.705 $X2=0 $Y2=0
cc_461 N_SCD_M1016_g N_VGND_c_2306_n 0.00527125f $X=2.295 $Y=0.445 $X2=0 $Y2=0
cc_462 N_SCD_c_522_n N_VGND_c_2306_n 3.90429e-19 $X=2.415 $Y=0.895 $X2=0 $Y2=0
cc_463 N_SCD_M1016_g N_VGND_c_2316_n 0.00482425f $X=2.295 $Y=0.445 $X2=0 $Y2=0
cc_464 N_SCD_M1016_g N_VGND_c_2320_n 0.00612587f $X=2.295 $Y=0.445 $X2=0 $Y2=0
cc_465 N_SCD_c_522_n N_VGND_c_2320_n 0.00273152f $X=2.415 $Y=0.895 $X2=0 $Y2=0
cc_466 N_A_570_47#_c_585_n N_A_914_245#_M1038_d 0.00896689f $X=5.95 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_467 N_A_570_47#_c_587_n N_A_914_245#_M1038_d 0.00584604f $X=6.035 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_468 N_A_570_47#_M1008_g N_A_914_245#_c_823_n 7.66947e-19 $X=4.285 $Y=0.905
+ $X2=0 $Y2=0
cc_469 N_A_570_47#_M1008_g N_A_914_245#_c_824_n 0.00117874f $X=4.285 $Y=0.905
+ $X2=0 $Y2=0
cc_470 N_A_570_47#_c_583_n N_A_914_245#_c_824_n 4.99549e-19 $X=5.27 $Y=0.7 $X2=0
+ $Y2=0
cc_471 N_A_570_47#_c_583_n N_A_914_245#_c_825_n 0.0356319f $X=5.27 $Y=0.7 $X2=0
+ $Y2=0
cc_472 N_A_570_47#_c_585_n N_A_914_245#_c_825_n 0.00304585f $X=5.95 $Y=0.34
+ $X2=0 $Y2=0
cc_473 N_A_570_47#_M1008_g N_A_914_245#_c_842_n 5.04789e-19 $X=4.285 $Y=0.905
+ $X2=0 $Y2=0
cc_474 N_A_570_47#_c_583_n N_A_914_245#_c_842_n 0.0187975f $X=5.27 $Y=0.7 $X2=0
+ $Y2=0
cc_475 N_A_570_47#_c_578_n N_A_914_245#_c_844_n 9.86411e-19 $X=6.16 $Y=1.095
+ $X2=0 $Y2=0
cc_476 N_A_570_47#_c_585_n N_A_914_245#_c_844_n 0.0127109f $X=5.95 $Y=0.34 $X2=0
+ $Y2=0
cc_477 N_A_570_47#_c_587_n N_A_914_245#_c_844_n 0.0261115f $X=6.035 $Y=1.095
+ $X2=0 $Y2=0
cc_478 N_A_570_47#_c_598_n N_A_914_245#_c_826_n 0.0235879f $X=6.455 $Y=1.26
+ $X2=0 $Y2=0
cc_479 N_A_570_47#_c_600_n N_A_914_245#_c_826_n 0.00103175f $X=6.52 $Y=1.26
+ $X2=0 $Y2=0
cc_480 N_A_570_47#_c_578_n N_A_914_245#_c_827_n 4.75666e-19 $X=6.16 $Y=1.095
+ $X2=0 $Y2=0
cc_481 N_A_570_47#_c_587_n N_A_914_245#_c_827_n 0.0117304f $X=6.035 $Y=1.095
+ $X2=0 $Y2=0
cc_482 N_A_570_47#_c_598_n N_A_914_245#_c_827_n 0.00255925f $X=6.455 $Y=1.26
+ $X2=0 $Y2=0
cc_483 N_A_570_47#_M1008_g N_A_914_245#_c_828_n 0.0330312f $X=4.285 $Y=0.905
+ $X2=0 $Y2=0
cc_484 N_A_570_47#_c_582_n N_A_914_245#_c_828_n 0.00119102f $X=4.49 $Y=0.615
+ $X2=0 $Y2=0
cc_485 N_A_570_47#_c_583_n N_A_914_245#_c_828_n 0.0112455f $X=5.27 $Y=0.7 $X2=0
+ $Y2=0
cc_486 N_A_570_47#_c_633_p N_A_914_245#_c_828_n 7.75791e-19 $X=5.355 $Y=0.615
+ $X2=0 $Y2=0
cc_487 N_A_570_47#_c_578_n N_A_786_139#_M1038_g 0.0120866f $X=6.16 $Y=1.095
+ $X2=0 $Y2=0
cc_488 N_A_570_47#_c_583_n N_A_786_139#_M1038_g 0.00581632f $X=5.27 $Y=0.7 $X2=0
+ $Y2=0
cc_489 N_A_570_47#_c_633_p N_A_786_139#_M1038_g 0.00641166f $X=5.355 $Y=0.615
+ $X2=0 $Y2=0
cc_490 N_A_570_47#_c_585_n N_A_786_139#_M1038_g 0.00842014f $X=5.95 $Y=0.34
+ $X2=0 $Y2=0
cc_491 N_A_570_47#_c_586_n N_A_786_139#_M1038_g 0.00365595f $X=5.44 $Y=0.34
+ $X2=0 $Y2=0
cc_492 N_A_570_47#_c_587_n N_A_786_139#_M1038_g 0.00211016f $X=6.035 $Y=1.095
+ $X2=0 $Y2=0
cc_493 N_A_570_47#_c_600_n N_A_786_139#_M1038_g 0.00859787f $X=6.52 $Y=1.26
+ $X2=0 $Y2=0
cc_494 N_A_570_47#_c_576_n N_A_786_139#_c_926_n 8.29898e-19 $X=4.21 $Y=0.25
+ $X2=0 $Y2=0
cc_495 N_A_570_47#_M1008_g N_A_786_139#_c_926_n 0.010501f $X=4.285 $Y=0.905
+ $X2=0 $Y2=0
cc_496 N_A_570_47#_c_581_n N_A_786_139#_c_926_n 0.0140954f $X=4.405 $Y=0.34
+ $X2=0 $Y2=0
cc_497 N_A_570_47#_c_584_n N_A_786_139#_c_926_n 0.0048601f $X=4.575 $Y=0.7 $X2=0
+ $Y2=0
cc_498 N_A_570_47#_c_601_n N_A_786_139#_c_933_n 0.00121426f $X=4.47 $Y=2.465
+ $X2=0 $Y2=0
cc_499 N_A_570_47#_M1008_g N_A_786_139#_c_933_n 0.00217334f $X=4.285 $Y=0.905
+ $X2=0 $Y2=0
cc_500 N_A_570_47#_c_601_n N_A_786_139#_c_935_n 0.00464682f $X=4.47 $Y=2.465
+ $X2=0 $Y2=0
cc_501 N_A_570_47#_c_602_n N_A_786_139#_c_935_n 0.0018428f $X=4.545 $Y=2.54
+ $X2=0 $Y2=0
cc_502 N_A_570_47#_c_602_n N_A_786_139#_c_941_n 0.00459979f $X=4.545 $Y=2.54
+ $X2=0 $Y2=0
cc_503 N_A_570_47#_c_603_n N_A_786_139#_c_944_n 0.00448633f $X=9.165 $Y=2.09
+ $X2=0 $Y2=0
cc_504 N_A_570_47#_c_580_n N_A_540_21#_M1025_g 0.00523061f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_505 N_A_570_47#_c_594_n N_A_540_21#_M1025_g 0.00610862f $X=3.17 $Y=0.465
+ $X2=0 $Y2=0
cc_506 N_A_570_47#_c_599_n N_A_540_21#_M1025_g 0.00786141f $X=3.405 $Y=0.25
+ $X2=0 $Y2=0
cc_507 N_A_570_47#_c_580_n N_A_540_21#_c_1069_n 0.0228028f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_508 N_A_570_47#_c_580_n N_A_540_21#_M1027_g 0.00240737f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_509 N_A_570_47#_c_606_n N_A_540_21#_M1027_g 0.00960874f $X=3.33 $Y=2.15 $X2=0
+ $Y2=0
cc_510 N_A_570_47#_c_607_n N_A_540_21#_M1027_g 0.00579578f $X=3.33 $Y=2.405
+ $X2=0 $Y2=0
cc_511 N_A_570_47#_c_580_n N_A_540_21#_c_1085_n 0.00453491f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_512 N_A_570_47#_c_606_n N_A_540_21#_c_1085_n 0.0111275f $X=3.33 $Y=2.15 $X2=0
+ $Y2=0
cc_513 N_A_570_47#_c_608_n N_A_540_21#_c_1085_n 0.00402734f $X=3.76 $Y=2.57
+ $X2=0 $Y2=0
cc_514 N_A_570_47#_c_611_n N_A_540_21#_c_1085_n 0.00397534f $X=3.76 $Y=2.465
+ $X2=0 $Y2=0
cc_515 N_A_570_47#_c_576_n N_A_540_21#_M1005_g 0.00830058f $X=4.21 $Y=0.25 $X2=0
+ $Y2=0
cc_516 N_A_570_47#_M1008_g N_A_540_21#_M1005_g 0.0122255f $X=4.285 $Y=0.905
+ $X2=0 $Y2=0
cc_517 N_A_570_47#_c_580_n N_A_540_21#_M1005_g 0.00516323f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_518 N_A_570_47#_c_581_n N_A_540_21#_M1005_g 0.00301984f $X=4.405 $Y=0.34
+ $X2=0 $Y2=0
cc_519 N_A_570_47#_c_594_n N_A_540_21#_M1005_g 0.00210729f $X=3.17 $Y=0.465
+ $X2=0 $Y2=0
cc_520 N_A_570_47#_c_599_n N_A_540_21#_M1005_g 0.00120024f $X=3.405 $Y=0.25
+ $X2=0 $Y2=0
cc_521 N_A_570_47#_c_601_n N_A_540_21#_c_1087_n 0.00964615f $X=4.47 $Y=2.465
+ $X2=0 $Y2=0
cc_522 N_A_570_47#_M1008_g N_A_540_21#_c_1087_n 0.00265814f $X=4.285 $Y=0.905
+ $X2=0 $Y2=0
cc_523 N_A_570_47#_c_601_n N_A_540_21#_M1022_g 0.0196088f $X=4.47 $Y=2.465 $X2=0
+ $Y2=0
cc_524 N_A_570_47#_c_598_n N_A_540_21#_c_1071_n 0.00393343f $X=6.455 $Y=1.26
+ $X2=0 $Y2=0
cc_525 N_A_570_47#_c_600_n N_A_540_21#_c_1071_n 0.0455666f $X=6.52 $Y=1.26 $X2=0
+ $Y2=0
cc_526 N_A_570_47#_c_579_n N_A_540_21#_M1026_g 0.00964816f $X=6.52 $Y=1.095
+ $X2=0 $Y2=0
cc_527 N_A_570_47#_c_588_n N_A_540_21#_M1026_g 0.00556974f $X=7.38 $Y=0.34 $X2=0
+ $Y2=0
cc_528 N_A_570_47#_c_589_n N_A_540_21#_M1026_g 0.00683964f $X=7.58 $Y=1.085
+ $X2=0 $Y2=0
cc_529 N_A_570_47#_c_591_n N_A_540_21#_M1026_g 0.00313848f $X=7.78 $Y=1.17 $X2=0
+ $Y2=0
cc_530 N_A_570_47#_c_598_n N_A_540_21#_M1026_g 3.22319e-19 $X=6.455 $Y=1.26
+ $X2=0 $Y2=0
cc_531 N_A_570_47#_c_600_n N_A_540_21#_M1026_g 0.00768464f $X=6.52 $Y=1.26 $X2=0
+ $Y2=0
cc_532 N_A_570_47#_c_591_n N_A_540_21#_c_1074_n 0.00111805f $X=7.78 $Y=1.17
+ $X2=0 $Y2=0
cc_533 N_A_570_47#_c_580_n N_A_540_21#_c_1075_n 0.00639285f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_534 N_A_570_47#_c_594_n N_A_540_21#_c_1075_n 0.00690374f $X=3.17 $Y=0.465
+ $X2=0 $Y2=0
cc_535 N_A_570_47#_c_580_n N_A_540_21#_c_1095_n 0.00347705f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_536 N_A_570_47#_c_611_n N_A_540_21#_c_1096_n 0.00964615f $X=3.76 $Y=2.465
+ $X2=0 $Y2=0
cc_537 N_A_570_47#_c_592_n N_A_540_21#_c_1101_n 7.48188e-19 $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_538 N_A_570_47#_c_603_n N_A_540_21#_c_1106_n 0.00880362f $X=9.165 $Y=2.09
+ $X2=0 $Y2=0
cc_539 N_A_570_47#_c_604_n N_A_540_21#_c_1106_n 0.00355563f $X=9.165 $Y=1.965
+ $X2=0 $Y2=0
cc_540 N_A_570_47#_c_590_n N_A_540_21#_c_1106_n 0.00610271f $X=9.09 $Y=1.17
+ $X2=0 $Y2=0
cc_541 N_A_570_47#_c_592_n N_A_540_21#_c_1106_n 0.021805f $X=9.255 $Y=1.56 $X2=0
+ $Y2=0
cc_542 N_A_570_47#_c_603_n N_A_540_21#_c_1107_n 0.00724545f $X=9.165 $Y=2.09
+ $X2=0 $Y2=0
cc_543 N_A_570_47#_c_604_n N_A_540_21#_c_1107_n 4.58566e-19 $X=9.165 $Y=1.965
+ $X2=0 $Y2=0
cc_544 N_A_570_47#_c_593_n N_A_540_21#_c_1107_n 9.74097e-19 $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_545 N_A_570_47#_c_603_n N_A_540_21#_c_1082_n 0.00127031f $X=9.165 $Y=2.09
+ $X2=0 $Y2=0
cc_546 N_A_570_47#_c_588_n N_A_1319_69#_M1012_d 0.0113669f $X=7.38 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_547 N_A_570_47#_c_590_n N_A_1319_69#_M1020_g 0.0135801f $X=9.09 $Y=1.17 $X2=0
+ $Y2=0
cc_548 N_A_570_47#_c_590_n N_A_1319_69#_M1007_g 0.0135356f $X=9.09 $Y=1.17 $X2=0
+ $Y2=0
cc_549 N_A_570_47#_c_590_n N_A_1319_69#_c_1317_n 0.00746018f $X=9.09 $Y=1.17
+ $X2=0 $Y2=0
cc_550 N_A_570_47#_c_592_n N_A_1319_69#_c_1317_n 0.00568477f $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_551 N_A_570_47#_c_579_n N_A_1319_69#_c_1321_n 0.00278513f $X=6.52 $Y=1.095
+ $X2=0 $Y2=0
cc_552 N_A_570_47#_c_589_n N_A_1319_69#_c_1321_n 0.0121398f $X=7.58 $Y=1.085
+ $X2=0 $Y2=0
cc_553 N_A_570_47#_c_591_n N_A_1319_69#_c_1321_n 0.0137153f $X=7.78 $Y=1.17
+ $X2=0 $Y2=0
cc_554 N_A_570_47#_c_598_n N_A_1319_69#_c_1321_n 0.0114446f $X=6.455 $Y=1.26
+ $X2=0 $Y2=0
cc_555 N_A_570_47#_c_600_n N_A_1319_69#_c_1321_n 0.00283821f $X=6.52 $Y=1.26
+ $X2=0 $Y2=0
cc_556 N_A_570_47#_c_590_n N_A_1319_69#_c_1323_n 0.0572601f $X=9.09 $Y=1.17
+ $X2=0 $Y2=0
cc_557 N_A_570_47#_c_591_n N_A_1319_69#_c_1323_n 0.0214984f $X=7.78 $Y=1.17
+ $X2=0 $Y2=0
cc_558 N_A_570_47#_c_603_n N_A_1319_69#_c_1358_n 0.0122916f $X=9.165 $Y=2.09
+ $X2=0 $Y2=0
cc_559 N_A_570_47#_c_579_n N_A_1319_69#_c_1359_n 0.00735876f $X=6.52 $Y=1.095
+ $X2=0 $Y2=0
cc_560 N_A_570_47#_c_588_n N_A_1319_69#_c_1359_n 0.0216064f $X=7.38 $Y=0.34
+ $X2=0 $Y2=0
cc_561 N_A_570_47#_c_589_n N_A_1319_69#_c_1359_n 0.0259734f $X=7.58 $Y=1.085
+ $X2=0 $Y2=0
cc_562 N_A_570_47#_c_591_n N_A_1319_69#_c_1324_n 0.0135853f $X=7.78 $Y=1.17
+ $X2=0 $Y2=0
cc_563 N_A_570_47#_c_590_n N_A_1319_69#_c_1342_n 0.023546f $X=9.09 $Y=1.17 $X2=0
+ $Y2=0
cc_564 N_A_570_47#_c_592_n N_A_1319_69#_c_1342_n 0.019012f $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_565 N_A_570_47#_c_593_n N_A_1319_69#_c_1342_n 0.0012425f $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_566 N_A_570_47#_c_592_n N_A_1319_69#_c_1325_n 0.00125609f $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_567 N_A_570_47#_c_593_n N_A_1319_69#_c_1325_n 0.0221793f $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_568 N_A_570_47#_c_603_n N_A_1319_69#_c_1344_n 0.0149378f $X=9.165 $Y=2.09
+ $X2=0 $Y2=0
cc_569 N_A_570_47#_c_588_n N_A_1493_21#_M1019_g 0.00747458f $X=7.38 $Y=0.34
+ $X2=0 $Y2=0
cc_570 N_A_570_47#_c_589_n N_A_1493_21#_M1019_g 0.0158943f $X=7.58 $Y=1.085
+ $X2=0 $Y2=0
cc_571 N_A_570_47#_c_591_n N_A_1493_21#_M1019_g 0.00255533f $X=7.78 $Y=1.17
+ $X2=0 $Y2=0
cc_572 N_A_570_47#_c_588_n N_A_1493_21#_c_1529_n 0.00212752f $X=7.38 $Y=0.34
+ $X2=0 $Y2=0
cc_573 N_A_570_47#_c_588_n N_A_1493_21#_c_1530_n 0.00128489f $X=7.38 $Y=0.34
+ $X2=0 $Y2=0
cc_574 N_A_570_47#_c_588_n N_A_1493_21#_M1006_g 0.00123283f $X=7.38 $Y=0.34
+ $X2=0 $Y2=0
cc_575 N_A_570_47#_c_589_n N_A_1493_21#_M1006_g 0.00504026f $X=7.58 $Y=1.085
+ $X2=0 $Y2=0
cc_576 N_A_570_47#_c_590_n N_A_1493_21#_M1006_g 0.00874669f $X=9.09 $Y=1.17
+ $X2=0 $Y2=0
cc_577 N_A_570_47#_c_603_n N_A_1493_21#_c_1546_n 0.073022f $X=9.165 $Y=2.09
+ $X2=0 $Y2=0
cc_578 N_A_570_47#_c_604_n N_A_1493_21#_c_1535_n 0.00797159f $X=9.165 $Y=1.965
+ $X2=0 $Y2=0
cc_579 N_A_570_47#_c_590_n N_A_1493_21#_c_1535_n 0.00529938f $X=9.09 $Y=1.17
+ $X2=0 $Y2=0
cc_580 N_A_570_47#_c_592_n N_A_1493_21#_c_1535_n 0.00639316f $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_581 N_A_570_47#_c_593_n N_A_1493_21#_c_1535_n 0.0199261f $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_582 N_A_570_47#_c_590_n N_A_1493_21#_c_1540_n 0.027455f $X=9.09 $Y=1.17 $X2=0
+ $Y2=0
cc_583 N_A_570_47#_c_593_n N_A_1493_21#_c_1540_n 7.81894e-19 $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_584 N_A_570_47#_c_590_n N_A_1493_21#_c_1541_n 0.00983917f $X=9.09 $Y=1.17
+ $X2=0 $Y2=0
cc_585 N_A_570_47#_c_593_n N_A_1493_21#_c_1541_n 2.48737e-19 $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_586 N_A_570_47#_c_590_n N_A_1493_21#_c_1542_n 0.00288132f $X=9.09 $Y=1.17
+ $X2=0 $Y2=0
cc_587 N_A_570_47#_c_590_n N_A_1493_21#_c_1545_n 8.73481e-19 $X=9.09 $Y=1.17
+ $X2=0 $Y2=0
cc_588 N_A_570_47#_c_593_n N_A_1493_21#_c_1545_n 0.00145749f $X=9.255 $Y=1.56
+ $X2=0 $Y2=0
cc_589 N_A_570_47#_c_604_n CLK 5.00887e-19 $X=9.165 $Y=1.965 $X2=0 $Y2=0
cc_590 N_A_570_47#_c_592_n CLK 0.0111791f $X=9.255 $Y=1.56 $X2=0 $Y2=0
cc_591 N_A_570_47#_c_593_n CLK 6.75068e-19 $X=9.255 $Y=1.56 $X2=0 $Y2=0
cc_592 N_A_570_47#_c_602_n N_VPWR_c_1857_n 0.00525141f $X=4.545 $Y=2.54 $X2=0
+ $Y2=0
cc_593 N_A_570_47#_c_603_n N_VPWR_c_1861_n 0.00939206f $X=9.165 $Y=2.09 $X2=0
+ $Y2=0
cc_594 N_A_570_47#_c_602_n N_VPWR_c_1854_n 0.00619862f $X=4.545 $Y=2.54 $X2=0
+ $Y2=0
cc_595 N_A_570_47#_c_603_n N_VPWR_c_1854_n 0.00797221f $X=9.165 $Y=2.09 $X2=0
+ $Y2=0
cc_596 N_A_570_47#_c_580_n N_A_282_477#_c_1997_n 0.020843f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_597 N_A_570_47#_c_594_n N_A_282_477#_c_1997_n 2.58353e-19 $X=3.17 $Y=0.465
+ $X2=0 $Y2=0
cc_598 N_A_570_47#_c_580_n N_A_282_477#_c_1999_n 0.0571074f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_599 N_A_570_47#_c_606_n N_A_282_477#_c_1999_n 0.0130061f $X=3.33 $Y=2.15
+ $X2=0 $Y2=0
cc_600 N_A_570_47#_c_607_n N_A_282_477#_c_1999_n 0.00760173f $X=3.33 $Y=2.405
+ $X2=0 $Y2=0
cc_601 N_A_570_47#_c_607_n N_A_282_477#_c_2053_n 0.00172674f $X=3.33 $Y=2.405
+ $X2=0 $Y2=0
cc_602 N_A_570_47#_M1027_d N_A_282_477#_c_2007_n 0.00175724f $X=3.15 $Y=2.385
+ $X2=0 $Y2=0
cc_603 N_A_570_47#_c_601_n N_A_282_477#_c_2007_n 0.00137294f $X=4.47 $Y=2.465
+ $X2=0 $Y2=0
cc_604 N_A_570_47#_c_602_n N_A_282_477#_c_2007_n 0.00326625f $X=4.545 $Y=2.54
+ $X2=0 $Y2=0
cc_605 N_A_570_47#_c_607_n N_A_282_477#_c_2007_n 0.0175416f $X=3.33 $Y=2.405
+ $X2=0 $Y2=0
cc_606 N_A_570_47#_c_608_n N_A_282_477#_c_2007_n 0.0323504f $X=3.76 $Y=2.57
+ $X2=0 $Y2=0
cc_607 N_A_570_47#_c_611_n N_A_282_477#_c_2007_n 0.00548882f $X=3.76 $Y=2.465
+ $X2=0 $Y2=0
cc_608 N_A_570_47#_c_580_n N_A_282_477#_c_2000_n 0.0305716f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_609 N_A_570_47#_c_606_n N_A_282_477#_c_2000_n 0.00655586f $X=3.33 $Y=2.15
+ $X2=0 $Y2=0
cc_610 N_A_570_47#_c_608_n N_A_282_477#_c_2010_n 0.00858889f $X=3.76 $Y=2.57
+ $X2=0 $Y2=0
cc_611 N_A_570_47#_c_611_n N_A_282_477#_c_2010_n 0.00329776f $X=3.76 $Y=2.465
+ $X2=0 $Y2=0
cc_612 N_A_570_47#_c_606_n N_A_282_477#_c_2011_n 0.00733446f $X=3.33 $Y=2.15
+ $X2=0 $Y2=0
cc_613 N_A_570_47#_c_607_n N_A_282_477#_c_2011_n 0.00707996f $X=3.33 $Y=2.405
+ $X2=0 $Y2=0
cc_614 N_A_570_47#_c_608_n N_A_282_477#_c_2011_n 0.0136071f $X=3.76 $Y=2.57
+ $X2=0 $Y2=0
cc_615 N_A_570_47#_c_611_n N_A_282_477#_c_2011_n 0.0016367f $X=3.76 $Y=2.465
+ $X2=0 $Y2=0
cc_616 N_A_570_47#_c_601_n N_A_282_477#_c_2012_n 0.0199658f $X=4.47 $Y=2.465
+ $X2=0 $Y2=0
cc_617 N_A_570_47#_c_602_n N_A_282_477#_c_2012_n 0.00490472f $X=4.545 $Y=2.54
+ $X2=0 $Y2=0
cc_618 N_A_570_47#_c_607_n N_A_282_477#_c_2012_n 0.00540594f $X=3.33 $Y=2.405
+ $X2=0 $Y2=0
cc_619 N_A_570_47#_c_608_n N_A_282_477#_c_2012_n 0.0262119f $X=3.76 $Y=2.57
+ $X2=0 $Y2=0
cc_620 N_A_570_47#_c_611_n N_A_282_477#_c_2012_n 7.823e-19 $X=3.76 $Y=2.465
+ $X2=0 $Y2=0
cc_621 N_A_570_47#_c_607_n N_A_282_477#_c_2013_n 0.00462618f $X=3.33 $Y=2.405
+ $X2=0 $Y2=0
cc_622 N_A_570_47#_c_576_n N_A_282_477#_c_2002_n 5.54456e-19 $X=4.21 $Y=0.25
+ $X2=0 $Y2=0
cc_623 N_A_570_47#_M1008_g N_A_282_477#_c_2002_n 2.12319e-19 $X=4.285 $Y=0.905
+ $X2=0 $Y2=0
cc_624 N_A_570_47#_c_580_n N_A_282_477#_c_2002_n 0.0200899f $X=3.085 $Y=1.98
+ $X2=0 $Y2=0
cc_625 N_A_570_47#_c_581_n N_A_282_477#_c_2002_n 0.00903258f $X=4.405 $Y=0.34
+ $X2=0 $Y2=0
cc_626 N_A_570_47#_c_596_n N_A_282_477#_c_2002_n 0.00718034f $X=3.57 $Y=0.42
+ $X2=0 $Y2=0
cc_627 N_A_570_47#_c_599_n N_A_282_477#_c_2002_n 0.00224756f $X=3.405 $Y=0.25
+ $X2=0 $Y2=0
cc_628 N_A_570_47#_c_603_n N_KAPWR_c_2176_n 0.00122482f $X=9.165 $Y=2.09 $X2=0
+ $Y2=0
cc_629 N_A_570_47#_M1027_d N_KAPWR_c_2164_n 6.82496e-19 $X=3.15 $Y=2.385 $X2=0
+ $Y2=0
cc_630 N_A_570_47#_c_601_n N_KAPWR_c_2164_n 0.00194672f $X=4.47 $Y=2.465 $X2=0
+ $Y2=0
cc_631 N_A_570_47#_c_602_n N_KAPWR_c_2164_n 0.00958502f $X=4.545 $Y=2.54 $X2=0
+ $Y2=0
cc_632 N_A_570_47#_c_603_n N_KAPWR_c_2164_n 0.00650428f $X=9.165 $Y=2.09 $X2=0
+ $Y2=0
cc_633 N_A_570_47#_c_606_n N_KAPWR_c_2164_n 0.00651503f $X=3.33 $Y=2.15 $X2=0
+ $Y2=0
cc_634 N_A_570_47#_c_607_n N_KAPWR_c_2164_n 0.00963984f $X=3.33 $Y=2.405 $X2=0
+ $Y2=0
cc_635 N_A_570_47#_c_608_n N_KAPWR_c_2164_n 0.0216925f $X=3.76 $Y=2.57 $X2=0
+ $Y2=0
cc_636 N_A_570_47#_c_611_n N_KAPWR_c_2164_n 0.00437773f $X=3.76 $Y=2.465 $X2=0
+ $Y2=0
cc_637 N_A_570_47#_c_583_n N_VGND_M1034_d 0.0140063f $X=5.27 $Y=0.7 $X2=0 $Y2=0
cc_638 N_A_570_47#_c_633_p N_VGND_M1034_d 0.00557095f $X=5.355 $Y=0.615 $X2=0
+ $Y2=0
cc_639 N_A_570_47#_c_586_n N_VGND_M1034_d 9.83603e-19 $X=5.44 $Y=0.34 $X2=0
+ $Y2=0
cc_640 N_A_570_47#_c_594_n N_VGND_c_2306_n 0.016826f $X=3.17 $Y=0.465 $X2=0
+ $Y2=0
cc_641 N_A_570_47#_c_576_n N_VGND_c_2307_n 0.00240303f $X=4.21 $Y=0.25 $X2=0
+ $Y2=0
cc_642 N_A_570_47#_c_581_n N_VGND_c_2307_n 0.0119249f $X=4.405 $Y=0.34 $X2=0
+ $Y2=0
cc_643 N_A_570_47#_c_582_n N_VGND_c_2307_n 0.0012256f $X=4.49 $Y=0.615 $X2=0
+ $Y2=0
cc_644 N_A_570_47#_c_583_n N_VGND_c_2307_n 0.018839f $X=5.27 $Y=0.7 $X2=0 $Y2=0
cc_645 N_A_570_47#_c_633_p N_VGND_c_2307_n 0.00122684f $X=5.355 $Y=0.615 $X2=0
+ $Y2=0
cc_646 N_A_570_47#_c_586_n N_VGND_c_2307_n 0.012091f $X=5.44 $Y=0.34 $X2=0 $Y2=0
cc_647 N_A_570_47#_c_588_n N_VGND_c_2308_n 0.0142967f $X=7.38 $Y=0.34 $X2=0
+ $Y2=0
cc_648 N_A_570_47#_c_589_n N_VGND_c_2308_n 0.0242969f $X=7.58 $Y=1.085 $X2=0
+ $Y2=0
cc_649 N_A_570_47#_c_590_n N_VGND_c_2308_n 0.0243655f $X=9.09 $Y=1.17 $X2=0
+ $Y2=0
cc_650 N_A_570_47#_c_578_n N_VGND_c_2311_n 0.00291433f $X=6.16 $Y=1.095 $X2=0
+ $Y2=0
cc_651 N_A_570_47#_c_579_n N_VGND_c_2311_n 0.0029147f $X=6.52 $Y=1.095 $X2=0
+ $Y2=0
cc_652 N_A_570_47#_c_583_n N_VGND_c_2311_n 0.00390843f $X=5.27 $Y=0.7 $X2=0
+ $Y2=0
cc_653 N_A_570_47#_c_585_n N_VGND_c_2311_n 0.0324632f $X=5.95 $Y=0.34 $X2=0
+ $Y2=0
cc_654 N_A_570_47#_c_586_n N_VGND_c_2311_n 0.0118414f $X=5.44 $Y=0.34 $X2=0
+ $Y2=0
cc_655 N_A_570_47#_c_588_n N_VGND_c_2311_n 0.107875f $X=7.38 $Y=0.34 $X2=0 $Y2=0
cc_656 N_A_570_47#_c_597_n N_VGND_c_2311_n 0.0120637f $X=6.035 $Y=0.34 $X2=0
+ $Y2=0
cc_657 N_A_570_47#_c_581_n N_VGND_c_2317_n 0.0119604f $X=4.405 $Y=0.34 $X2=0
+ $Y2=0
cc_658 N_A_570_47#_c_583_n N_VGND_c_2317_n 0.00407135f $X=5.27 $Y=0.7 $X2=0
+ $Y2=0
cc_659 N_A_570_47#_c_594_n N_VGND_c_2317_n 0.0987335f $X=3.17 $Y=0.465 $X2=0
+ $Y2=0
cc_660 N_A_570_47#_c_599_n N_VGND_c_2317_n 0.0214756f $X=3.405 $Y=0.25 $X2=0
+ $Y2=0
cc_661 N_A_570_47#_M1025_d N_VGND_c_2320_n 0.00226194f $X=2.85 $Y=0.235 $X2=0
+ $Y2=0
cc_662 N_A_570_47#_c_576_n N_VGND_c_2320_n 0.0204505f $X=4.21 $Y=0.25 $X2=0
+ $Y2=0
cc_663 N_A_570_47#_c_578_n N_VGND_c_2320_n 0.00405957f $X=6.16 $Y=1.095 $X2=0
+ $Y2=0
cc_664 N_A_570_47#_c_579_n N_VGND_c_2320_n 0.00424108f $X=6.52 $Y=1.095 $X2=0
+ $Y2=0
cc_665 N_A_570_47#_c_581_n N_VGND_c_2320_n 0.00656672f $X=4.405 $Y=0.34 $X2=0
+ $Y2=0
cc_666 N_A_570_47#_c_583_n N_VGND_c_2320_n 0.0139809f $X=5.27 $Y=0.7 $X2=0 $Y2=0
cc_667 N_A_570_47#_c_585_n N_VGND_c_2320_n 0.0186441f $X=5.95 $Y=0.34 $X2=0
+ $Y2=0
cc_668 N_A_570_47#_c_586_n N_VGND_c_2320_n 0.00640666f $X=5.44 $Y=0.34 $X2=0
+ $Y2=0
cc_669 N_A_570_47#_c_588_n N_VGND_c_2320_n 0.0602353f $X=7.38 $Y=0.34 $X2=0
+ $Y2=0
cc_670 N_A_570_47#_c_594_n N_VGND_c_2320_n 0.0546037f $X=3.17 $Y=0.465 $X2=0
+ $Y2=0
cc_671 N_A_570_47#_c_597_n N_VGND_c_2320_n 0.00644906f $X=6.035 $Y=0.34 $X2=0
+ $Y2=0
cc_672 N_A_570_47#_c_599_n N_VGND_c_2320_n 0.00855338f $X=3.405 $Y=0.25 $X2=0
+ $Y2=0
cc_673 N_A_570_47#_c_584_n A_872_139# 0.00553173f $X=4.575 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_674 N_A_570_47#_c_588_n A_1247_69# 0.00184804f $X=7.38 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_675 N_A_570_47#_c_589_n A_1451_113# 0.00367027f $X=7.58 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_676 N_A_914_245#_c_823_n N_A_786_139#_M1038_g 0.00197384f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_677 N_A_914_245#_c_824_n N_A_786_139#_M1038_g 9.01905e-19 $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_678 N_A_914_245#_c_825_n N_A_786_139#_M1038_g 0.0137328f $X=5.61 $Y=1.04
+ $X2=0 $Y2=0
cc_679 N_A_914_245#_c_826_n N_A_786_139#_M1038_g 0.0101462f $X=5.695 $Y=2.105
+ $X2=0 $Y2=0
cc_680 N_A_914_245#_c_828_n N_A_786_139#_M1038_g 0.00955619f $X=4.735 $Y=1.225
+ $X2=0 $Y2=0
cc_681 N_A_914_245#_c_826_n N_A_786_139#_c_929_n 0.00289172f $X=5.695 $Y=2.105
+ $X2=0 $Y2=0
cc_682 N_A_914_245#_c_831_n N_A_786_139#_c_929_n 0.0174048f $X=6.335 $Y=2.28
+ $X2=0 $Y2=0
cc_683 N_A_914_245#_c_833_n N_A_786_139#_c_929_n 0.00528385f $X=5.455 $Y=2.325
+ $X2=0 $Y2=0
cc_684 N_A_914_245#_c_834_n N_A_786_139#_c_929_n 0.0129796f $X=6.5 $Y=2.28 $X2=0
+ $Y2=0
cc_685 N_A_914_245#_c_823_n N_A_786_139#_c_926_n 0.0200022f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_686 N_A_914_245#_c_824_n N_A_786_139#_c_926_n 0.00291355f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_687 N_A_914_245#_c_842_n N_A_786_139#_c_926_n 0.00381999f $X=4.9 $Y=1.04
+ $X2=0 $Y2=0
cc_688 N_A_914_245#_c_828_n N_A_786_139#_c_926_n 0.00121037f $X=4.735 $Y=1.225
+ $X2=0 $Y2=0
cc_689 N_A_914_245#_c_823_n N_A_786_139#_c_933_n 0.00186111f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_690 N_A_914_245#_c_832_n N_A_786_139#_c_935_n 0.0152507f $X=5.78 $Y=2.28
+ $X2=0 $Y2=0
cc_691 N_A_914_245#_c_833_n N_A_786_139#_c_935_n 7.43628e-19 $X=5.455 $Y=2.325
+ $X2=0 $Y2=0
cc_692 N_A_914_245#_c_825_n N_A_786_139#_c_936_n 0.00576413f $X=5.61 $Y=1.04
+ $X2=0 $Y2=0
cc_693 N_A_914_245#_c_826_n N_A_786_139#_c_936_n 0.0135709f $X=5.695 $Y=2.105
+ $X2=0 $Y2=0
cc_694 N_A_914_245#_c_832_n N_A_786_139#_c_936_n 0.0106788f $X=5.78 $Y=2.28
+ $X2=0 $Y2=0
cc_695 N_A_914_245#_M1036_g N_A_786_139#_c_937_n 0.0123058f $X=5.365 $Y=2.86
+ $X2=0 $Y2=0
cc_696 N_A_914_245#_c_832_n N_A_786_139#_c_937_n 0.0492413f $X=5.78 $Y=2.28
+ $X2=0 $Y2=0
cc_697 N_A_914_245#_c_833_n N_A_786_139#_c_937_n 0.00420524f $X=5.455 $Y=2.325
+ $X2=0 $Y2=0
cc_698 N_A_914_245#_c_823_n N_A_786_139#_c_927_n 0.0164771f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_699 N_A_914_245#_c_824_n N_A_786_139#_c_927_n 9.05556e-19 $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_700 N_A_914_245#_c_825_n N_A_786_139#_c_927_n 0.0258235f $X=5.61 $Y=1.04
+ $X2=0 $Y2=0
cc_701 N_A_914_245#_c_826_n N_A_786_139#_c_927_n 0.0328298f $X=5.695 $Y=2.105
+ $X2=0 $Y2=0
cc_702 N_A_914_245#_M1023_d N_A_786_139#_c_939_n 0.00113814f $X=6.35 $Y=2.125
+ $X2=0 $Y2=0
cc_703 N_A_914_245#_c_831_n N_A_786_139#_c_939_n 0.00262906f $X=6.335 $Y=2.28
+ $X2=0 $Y2=0
cc_704 N_A_914_245#_c_834_n N_A_786_139#_c_939_n 0.0208796f $X=6.5 $Y=2.28 $X2=0
+ $Y2=0
cc_705 N_A_914_245#_c_823_n N_A_786_139#_c_940_n 0.0268602f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_706 N_A_914_245#_c_824_n N_A_786_139#_c_940_n 0.00117923f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_707 N_A_914_245#_c_825_n N_A_786_139#_c_940_n 8.60188e-19 $X=5.61 $Y=1.04
+ $X2=0 $Y2=0
cc_708 N_A_914_245#_M1036_g N_A_786_139#_c_941_n 0.00215476f $X=5.365 $Y=2.86
+ $X2=0 $Y2=0
cc_709 N_A_914_245#_M1036_g N_A_786_139#_c_942_n 0.00301074f $X=5.365 $Y=2.86
+ $X2=0 $Y2=0
cc_710 N_A_914_245#_c_831_n N_A_786_139#_c_942_n 0.011176f $X=6.335 $Y=2.28
+ $X2=0 $Y2=0
cc_711 N_A_914_245#_c_834_n N_A_786_139#_c_942_n 0.00489182f $X=6.5 $Y=2.28
+ $X2=0 $Y2=0
cc_712 N_A_914_245#_c_823_n N_A_786_139#_c_928_n 0.00121458f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_713 N_A_914_245#_c_824_n N_A_786_139#_c_928_n 0.0186271f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_714 N_A_914_245#_c_825_n N_A_786_139#_c_928_n 0.00690382f $X=5.61 $Y=1.04
+ $X2=0 $Y2=0
cc_715 N_A_914_245#_c_824_n N_A_540_21#_M1005_g 0.0034243f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_716 N_A_914_245#_c_823_n N_A_540_21#_c_1087_n 3.64187e-19 $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_717 N_A_914_245#_c_824_n N_A_540_21#_c_1087_n 0.0176355f $X=4.735 $Y=1.39
+ $X2=0 $Y2=0
cc_718 N_A_914_245#_c_826_n N_A_540_21#_M1022_g 0.00352291f $X=5.695 $Y=2.105
+ $X2=0 $Y2=0
cc_719 N_A_914_245#_c_832_n N_A_540_21#_M1022_g 0.00215061f $X=5.78 $Y=2.28
+ $X2=0 $Y2=0
cc_720 N_A_914_245#_c_833_n N_A_540_21#_M1022_g 0.0561686f $X=5.455 $Y=2.325
+ $X2=0 $Y2=0
cc_721 N_A_914_245#_c_825_n N_A_540_21#_c_1089_n 0.00144381f $X=5.61 $Y=1.04
+ $X2=0 $Y2=0
cc_722 N_A_914_245#_c_826_n N_A_540_21#_c_1089_n 0.0187667f $X=5.695 $Y=2.105
+ $X2=0 $Y2=0
cc_723 N_A_914_245#_c_831_n N_A_540_21#_c_1089_n 0.00672123f $X=6.335 $Y=2.28
+ $X2=0 $Y2=0
cc_724 N_A_914_245#_c_832_n N_A_540_21#_c_1089_n 0.00573529f $X=5.78 $Y=2.28
+ $X2=0 $Y2=0
cc_725 N_A_914_245#_c_833_n N_A_540_21#_c_1089_n 0.0195639f $X=5.455 $Y=2.325
+ $X2=0 $Y2=0
cc_726 N_A_914_245#_c_831_n N_A_540_21#_c_1071_n 0.00880404f $X=6.335 $Y=2.28
+ $X2=0 $Y2=0
cc_727 N_A_914_245#_c_834_n N_A_540_21#_c_1071_n 0.010657f $X=6.5 $Y=2.28 $X2=0
+ $Y2=0
cc_728 N_A_914_245#_c_834_n N_A_540_21#_c_1091_n 0.00353049f $X=6.5 $Y=2.28
+ $X2=0 $Y2=0
cc_729 N_A_914_245#_c_825_n N_A_540_21#_c_1097_n 0.00101558f $X=5.61 $Y=1.04
+ $X2=0 $Y2=0
cc_730 N_A_914_245#_c_826_n N_A_540_21#_c_1076_n 0.00798499f $X=5.695 $Y=2.105
+ $X2=0 $Y2=0
cc_731 N_A_914_245#_c_834_n N_A_1319_69#_c_1335_n 0.00710417f $X=6.5 $Y=2.28
+ $X2=0 $Y2=0
cc_732 N_A_914_245#_c_831_n N_VPWR_M1036_d 0.00319583f $X=6.335 $Y=2.28 $X2=0
+ $Y2=0
cc_733 N_A_914_245#_M1036_g N_VPWR_c_1857_n 0.00390008f $X=5.365 $Y=2.86 $X2=0
+ $Y2=0
cc_734 N_A_914_245#_M1036_g N_VPWR_c_1854_n 0.00564254f $X=5.365 $Y=2.86 $X2=0
+ $Y2=0
cc_735 N_A_914_245#_M1036_g N_VPWR_c_1866_n 0.00654528f $X=5.365 $Y=2.86 $X2=0
+ $Y2=0
cc_736 N_A_914_245#_M1023_d N_KAPWR_c_2164_n 0.001781f $X=6.35 $Y=2.125 $X2=0
+ $Y2=0
cc_737 N_A_914_245#_M1036_g N_KAPWR_c_2164_n 0.00446495f $X=5.365 $Y=2.86 $X2=0
+ $Y2=0
cc_738 N_A_914_245#_c_831_n N_KAPWR_c_2164_n 0.00584325f $X=6.335 $Y=2.28 $X2=0
+ $Y2=0
cc_739 N_A_914_245#_c_832_n N_KAPWR_c_2164_n 0.00478771f $X=5.78 $Y=2.28 $X2=0
+ $Y2=0
cc_740 N_A_914_245#_c_834_n N_KAPWR_c_2164_n 0.025744f $X=6.5 $Y=2.28 $X2=0
+ $Y2=0
cc_741 N_A_914_245#_c_825_n N_VGND_M1034_d 0.00598865f $X=5.61 $Y=1.04 $X2=0
+ $Y2=0
cc_742 N_A_914_245#_c_842_n N_VGND_M1034_d 0.00101671f $X=4.9 $Y=1.04 $X2=0
+ $Y2=0
cc_743 N_A_914_245#_c_828_n N_VGND_c_2317_n 0.00294293f $X=4.735 $Y=1.225 $X2=0
+ $Y2=0
cc_744 N_A_914_245#_c_828_n N_VGND_c_2320_n 0.0045051f $X=4.735 $Y=1.225 $X2=0
+ $Y2=0
cc_745 N_A_786_139#_c_926_n N_A_540_21#_M1005_g 0.00893747f $X=4.07 $Y=0.905
+ $X2=0 $Y2=0
cc_746 N_A_786_139#_c_934_n N_A_540_21#_M1005_g 0.00201289f $X=4.235 $Y=1.81
+ $X2=0 $Y2=0
cc_747 N_A_786_139#_c_933_n N_A_540_21#_c_1087_n 0.0116565f $X=4.595 $Y=1.81
+ $X2=0 $Y2=0
cc_748 N_A_786_139#_c_934_n N_A_540_21#_c_1087_n 0.0110739f $X=4.235 $Y=1.81
+ $X2=0 $Y2=0
cc_749 N_A_786_139#_c_935_n N_A_540_21#_c_1087_n 0.0112313f $X=4.76 $Y=2.625
+ $X2=0 $Y2=0
cc_750 N_A_786_139#_c_940_n N_A_540_21#_c_1087_n 0.00409344f $X=4.76 $Y=1.81
+ $X2=0 $Y2=0
cc_751 N_A_786_139#_c_935_n N_A_540_21#_M1022_g 0.0264164f $X=4.76 $Y=2.625
+ $X2=0 $Y2=0
cc_752 N_A_786_139#_c_937_n N_A_540_21#_M1022_g 0.0113296f $X=5.995 $Y=2.71
+ $X2=0 $Y2=0
cc_753 N_A_786_139#_c_941_n N_A_540_21#_M1022_g 0.00692209f $X=4.76 $Y=2.71
+ $X2=0 $Y2=0
cc_754 N_A_786_139#_c_936_n N_A_540_21#_c_1089_n 0.0195936f $X=5.11 $Y=1.81
+ $X2=0 $Y2=0
cc_755 N_A_786_139#_c_937_n N_A_540_21#_c_1089_n 0.00487452f $X=5.995 $Y=2.71
+ $X2=0 $Y2=0
cc_756 N_A_786_139#_c_928_n N_A_540_21#_c_1089_n 0.0292966f $X=5.48 $Y=1.425
+ $X2=0 $Y2=0
cc_757 N_A_786_139#_c_929_n N_A_540_21#_c_1071_n 0.0100137f $X=6.275 $Y=3.075
+ $X2=0 $Y2=0
cc_758 N_A_786_139#_c_929_n N_A_540_21#_c_1091_n 0.0212536f $X=6.275 $Y=3.075
+ $X2=0 $Y2=0
cc_759 N_A_786_139#_c_930_n N_A_540_21#_c_1091_n 0.00933385f $X=8.01 $Y=3.15
+ $X2=0 $Y2=0
cc_760 N_A_786_139#_c_939_n N_A_540_21#_c_1091_n 0.00310404f $X=8.01 $Y=2.99
+ $X2=0 $Y2=0
cc_761 N_A_786_139#_c_930_n N_A_540_21#_c_1093_n 0.00933385f $X=8.01 $Y=3.15
+ $X2=0 $Y2=0
cc_762 N_A_786_139#_c_939_n N_A_540_21#_c_1093_n 0.00273636f $X=8.01 $Y=2.99
+ $X2=0 $Y2=0
cc_763 N_A_786_139#_c_935_n N_A_540_21#_c_1097_n 0.00270075f $X=4.76 $Y=2.625
+ $X2=0 $Y2=0
cc_764 N_A_786_139#_c_936_n N_A_540_21#_c_1097_n 0.00851924f $X=5.11 $Y=1.81
+ $X2=0 $Y2=0
cc_765 N_A_786_139#_c_940_n N_A_540_21#_c_1097_n 6.14813e-19 $X=4.76 $Y=1.81
+ $X2=0 $Y2=0
cc_766 N_A_786_139#_c_944_n N_A_540_21#_c_1082_n 0.00383676f $X=8.175 $Y=2.91
+ $X2=0 $Y2=0
cc_767 N_A_786_139#_c_939_n N_A_1319_69#_c_1334_n 0.0102584f $X=8.01 $Y=2.99
+ $X2=0 $Y2=0
cc_768 N_A_786_139#_c_943_n N_A_1319_69#_c_1334_n 0.0105366f $X=8.175 $Y=2.91
+ $X2=0 $Y2=0
cc_769 N_A_786_139#_c_944_n N_A_1319_69#_c_1334_n 0.00133836f $X=8.175 $Y=2.91
+ $X2=0 $Y2=0
cc_770 N_A_786_139#_c_939_n N_A_1319_69#_c_1335_n 0.0224621f $X=8.01 $Y=2.99
+ $X2=0 $Y2=0
cc_771 N_A_786_139#_c_943_n N_A_1319_69#_c_1344_n 0.0108679f $X=8.175 $Y=2.91
+ $X2=0 $Y2=0
cc_772 N_A_786_139#_c_944_n N_A_1319_69#_c_1344_n 0.00239429f $X=8.175 $Y=2.91
+ $X2=0 $Y2=0
cc_773 N_A_786_139#_c_937_n N_VPWR_M1036_d 0.00698915f $X=5.995 $Y=2.71 $X2=0
+ $Y2=0
cc_774 N_A_786_139#_c_942_n N_VPWR_M1036_d 0.00571808f $X=6.08 $Y=2.71 $X2=0
+ $Y2=0
cc_775 N_A_786_139#_c_937_n N_VPWR_c_1857_n 0.0123942f $X=5.995 $Y=2.71 $X2=0
+ $Y2=0
cc_776 N_A_786_139#_c_941_n N_VPWR_c_1857_n 0.0233446f $X=4.76 $Y=2.71 $X2=0
+ $Y2=0
cc_777 N_A_786_139#_c_931_n N_VPWR_c_1861_n 0.0451836f $X=6.35 $Y=3.15 $X2=0
+ $Y2=0
cc_778 N_A_786_139#_c_937_n N_VPWR_c_1861_n 0.00412764f $X=5.995 $Y=2.71 $X2=0
+ $Y2=0
cc_779 N_A_786_139#_c_939_n N_VPWR_c_1861_n 0.118383f $X=8.01 $Y=2.99 $X2=0
+ $Y2=0
cc_780 N_A_786_139#_c_942_n N_VPWR_c_1861_n 0.0116773f $X=6.08 $Y=2.71 $X2=0
+ $Y2=0
cc_781 N_A_786_139#_c_943_n N_VPWR_c_1861_n 0.0212434f $X=8.175 $Y=2.91 $X2=0
+ $Y2=0
cc_782 N_A_786_139#_c_930_n N_VPWR_c_1854_n 0.0299428f $X=8.01 $Y=3.15 $X2=0
+ $Y2=0
cc_783 N_A_786_139#_c_931_n N_VPWR_c_1854_n 0.00544415f $X=6.35 $Y=3.15 $X2=0
+ $Y2=0
cc_784 N_A_786_139#_c_937_n N_VPWR_c_1854_n 0.00307306f $X=5.995 $Y=2.71 $X2=0
+ $Y2=0
cc_785 N_A_786_139#_c_939_n N_VPWR_c_1854_n 0.0140507f $X=8.01 $Y=2.99 $X2=0
+ $Y2=0
cc_786 N_A_786_139#_c_941_n N_VPWR_c_1854_n 0.00303042f $X=4.76 $Y=2.71 $X2=0
+ $Y2=0
cc_787 N_A_786_139#_c_942_n N_VPWR_c_1854_n 0.00151024f $X=6.08 $Y=2.71 $X2=0
+ $Y2=0
cc_788 N_A_786_139#_c_943_n N_VPWR_c_1854_n 0.00250438f $X=8.175 $Y=2.91 $X2=0
+ $Y2=0
cc_789 N_A_786_139#_c_944_n N_VPWR_c_1854_n 0.008512f $X=8.175 $Y=2.91 $X2=0
+ $Y2=0
cc_790 N_A_786_139#_c_931_n N_VPWR_c_1866_n 0.00339574f $X=6.35 $Y=3.15 $X2=0
+ $Y2=0
cc_791 N_A_786_139#_c_937_n N_VPWR_c_1866_n 0.0220718f $X=5.995 $Y=2.71 $X2=0
+ $Y2=0
cc_792 N_A_786_139#_c_941_n N_VPWR_c_1866_n 0.00159381f $X=4.76 $Y=2.71 $X2=0
+ $Y2=0
cc_793 N_A_786_139#_c_942_n N_VPWR_c_1866_n 0.00855308f $X=6.08 $Y=2.71 $X2=0
+ $Y2=0
cc_794 N_A_786_139#_c_941_n N_A_282_477#_c_2007_n 0.00714249f $X=4.76 $Y=2.71
+ $X2=0 $Y2=0
cc_795 N_A_786_139#_c_934_n N_A_282_477#_c_2000_n 0.0126741f $X=4.235 $Y=1.81
+ $X2=0 $Y2=0
cc_796 N_A_786_139#_c_933_n N_A_282_477#_c_2010_n 0.0152946f $X=4.595 $Y=1.81
+ $X2=0 $Y2=0
cc_797 N_A_786_139#_c_934_n N_A_282_477#_c_2010_n 0.0212331f $X=4.235 $Y=1.81
+ $X2=0 $Y2=0
cc_798 N_A_786_139#_c_935_n N_A_282_477#_c_2010_n 0.0150383f $X=4.76 $Y=2.625
+ $X2=0 $Y2=0
cc_799 N_A_786_139#_c_935_n N_A_282_477#_c_2012_n 0.045275f $X=4.76 $Y=2.625
+ $X2=0 $Y2=0
cc_800 N_A_786_139#_c_926_n N_A_282_477#_c_2002_n 0.0559818f $X=4.07 $Y=0.905
+ $X2=0 $Y2=0
cc_801 N_A_786_139#_c_937_n A_1010_530# 0.00133423f $X=5.995 $Y=2.71 $X2=-0.19
+ $Y2=-0.245
cc_802 N_A_786_139#_c_929_n N_KAPWR_c_2164_n 0.00666989f $X=6.275 $Y=3.075 $X2=0
+ $Y2=0
cc_803 N_A_786_139#_c_937_n N_KAPWR_c_2164_n 0.0509743f $X=5.995 $Y=2.71 $X2=0
+ $Y2=0
cc_804 N_A_786_139#_c_939_n N_KAPWR_c_2164_n 0.0548122f $X=8.01 $Y=2.99 $X2=0
+ $Y2=0
cc_805 N_A_786_139#_c_941_n N_KAPWR_c_2164_n 0.0376714f $X=4.76 $Y=2.71 $X2=0
+ $Y2=0
cc_806 N_A_786_139#_c_942_n N_KAPWR_c_2164_n 0.0194881f $X=6.08 $Y=2.71 $X2=0
+ $Y2=0
cc_807 N_A_786_139#_c_943_n N_KAPWR_c_2164_n 0.020347f $X=8.175 $Y=2.91 $X2=0
+ $Y2=0
cc_808 N_A_786_139#_c_944_n N_KAPWR_c_2164_n 0.00650736f $X=8.175 $Y=2.91 $X2=0
+ $Y2=0
cc_809 N_A_786_139#_M1038_g N_VGND_c_2307_n 0.00190212f $X=5.48 $Y=0.665 $X2=0
+ $Y2=0
cc_810 N_A_786_139#_M1038_g N_VGND_c_2311_n 0.00291433f $X=5.48 $Y=0.665 $X2=0
+ $Y2=0
cc_811 N_A_786_139#_M1038_g N_VGND_c_2320_n 0.00440467f $X=5.48 $Y=0.665 $X2=0
+ $Y2=0
cc_812 N_A_540_21#_c_1103_n N_A_1319_69#_c_1326_n 0.00168271f $X=11.18 $Y=2.085
+ $X2=0 $Y2=0
cc_813 N_A_540_21#_c_1080_n N_A_1319_69#_c_1328_n 0.00170526f $X=11.265 $Y=2
+ $X2=0 $Y2=0
cc_814 N_A_540_21#_M1026_g N_A_1319_69#_c_1321_n 0.0178538f $X=7.18 $Y=0.775
+ $X2=0 $Y2=0
cc_815 N_A_540_21#_c_1091_n N_A_1319_69#_c_1322_n 0.00205152f $X=6.785 $Y=1.785
+ $X2=0 $Y2=0
cc_816 N_A_540_21#_c_1093_n N_A_1319_69#_c_1322_n 0.0110102f $X=7.145 $Y=1.785
+ $X2=0 $Y2=0
cc_817 N_A_540_21#_M1026_g N_A_1319_69#_c_1322_n 0.00250392f $X=7.18 $Y=0.775
+ $X2=0 $Y2=0
cc_818 N_A_540_21#_c_1074_n N_A_1319_69#_c_1322_n 0.0203111f $X=8.01 $Y=1.71
+ $X2=0 $Y2=0
cc_819 N_A_540_21#_c_1078_n N_A_1319_69#_c_1322_n 0.00799646f $X=7.162 $Y=1.71
+ $X2=0 $Y2=0
cc_820 N_A_540_21#_c_1105_n N_A_1319_69#_c_1322_n 0.0118413f $X=8.175 $Y=1.93
+ $X2=0 $Y2=0
cc_821 N_A_540_21#_c_1082_n N_A_1319_69#_c_1322_n 0.0056463f $X=8.175 $Y=1.71
+ $X2=0 $Y2=0
cc_822 N_A_540_21#_c_1074_n N_A_1319_69#_c_1323_n 0.0206024f $X=8.01 $Y=1.71
+ $X2=0 $Y2=0
cc_823 N_A_540_21#_c_1105_n N_A_1319_69#_c_1323_n 0.0247693f $X=8.175 $Y=1.93
+ $X2=0 $Y2=0
cc_824 N_A_540_21#_c_1106_n N_A_1319_69#_c_1323_n 0.00999161f $X=9.235 $Y=2.047
+ $X2=0 $Y2=0
cc_825 N_A_540_21#_c_1074_n N_A_1319_69#_c_1334_n 0.00646389f $X=8.01 $Y=1.71
+ $X2=0 $Y2=0
cc_826 N_A_540_21#_c_1105_n N_A_1319_69#_c_1334_n 0.02413f $X=8.175 $Y=1.93
+ $X2=0 $Y2=0
cc_827 N_A_540_21#_c_1106_n N_A_1319_69#_c_1334_n 0.0289233f $X=9.235 $Y=2.047
+ $X2=0 $Y2=0
cc_828 N_A_540_21#_c_1082_n N_A_1319_69#_c_1334_n 0.00134938f $X=8.175 $Y=1.71
+ $X2=0 $Y2=0
cc_829 N_A_540_21#_c_1091_n N_A_1319_69#_c_1335_n 0.00136768f $X=6.785 $Y=1.785
+ $X2=0 $Y2=0
cc_830 N_A_540_21#_c_1093_n N_A_1319_69#_c_1335_n 0.0105791f $X=7.145 $Y=1.785
+ $X2=0 $Y2=0
cc_831 N_A_540_21#_c_1101_n N_A_1319_69#_c_1358_n 0.0110768f $X=10.515 $Y=2.085
+ $X2=0 $Y2=0
cc_832 N_A_540_21#_c_1106_n N_A_1319_69#_c_1358_n 0.0080038f $X=9.235 $Y=2.047
+ $X2=0 $Y2=0
cc_833 N_A_540_21#_c_1107_n N_A_1319_69#_c_1358_n 0.0486656f $X=9.405 $Y=2.047
+ $X2=0 $Y2=0
cc_834 N_A_540_21#_c_1102_n N_A_1319_69#_c_1336_n 0.0091171f $X=10.6 $Y=2.405
+ $X2=0 $Y2=0
cc_835 N_A_540_21#_c_1102_n N_A_1319_69#_c_1337_n 0.0119316f $X=10.6 $Y=2.405
+ $X2=0 $Y2=0
cc_836 N_A_540_21#_c_1102_n N_A_1319_69#_c_1339_n 0.0091171f $X=10.6 $Y=2.405
+ $X2=0 $Y2=0
cc_837 N_A_540_21#_c_1103_n N_A_1319_69#_c_1401_n 0.0201438f $X=11.18 $Y=2.085
+ $X2=0 $Y2=0
cc_838 N_A_540_21#_c_1103_n N_A_1319_69#_c_1402_n 0.0110768f $X=11.18 $Y=2.085
+ $X2=0 $Y2=0
cc_839 N_A_540_21#_M1026_g N_A_1319_69#_c_1359_n 0.00632057f $X=7.18 $Y=0.775
+ $X2=0 $Y2=0
cc_840 N_A_540_21#_c_1072_n N_A_1319_69#_c_1324_n 0.00356788f $X=7.07 $Y=1.71
+ $X2=0 $Y2=0
cc_841 N_A_540_21#_M1026_g N_A_1319_69#_c_1324_n 0.0161155f $X=7.18 $Y=0.775
+ $X2=0 $Y2=0
cc_842 N_A_540_21#_c_1106_n N_A_1319_69#_c_1342_n 0.0247729f $X=9.235 $Y=2.047
+ $X2=0 $Y2=0
cc_843 N_A_540_21#_c_1082_n N_A_1319_69#_c_1342_n 9.22812e-19 $X=8.175 $Y=1.71
+ $X2=0 $Y2=0
cc_844 N_A_540_21#_c_1106_n N_A_1319_69#_c_1325_n 0.00228259f $X=9.235 $Y=2.047
+ $X2=0 $Y2=0
cc_845 N_A_540_21#_c_1082_n N_A_1319_69#_c_1325_n 0.00857262f $X=8.175 $Y=1.71
+ $X2=0 $Y2=0
cc_846 N_A_540_21#_c_1106_n N_A_1319_69#_c_1344_n 0.023919f $X=9.235 $Y=2.047
+ $X2=0 $Y2=0
cc_847 N_A_540_21#_M1026_g N_A_1493_21#_M1019_g 0.0397972f $X=7.18 $Y=0.775
+ $X2=0 $Y2=0
cc_848 N_A_540_21#_c_1074_n N_A_1493_21#_M1019_g 0.00250476f $X=8.01 $Y=1.71
+ $X2=0 $Y2=0
cc_849 N_A_540_21#_c_1074_n N_A_1493_21#_M1006_g 0.0024696f $X=8.01 $Y=1.71
+ $X2=0 $Y2=0
cc_850 N_A_540_21#_c_1101_n N_A_1493_21#_c_1546_n 0.0201733f $X=10.515 $Y=2.085
+ $X2=0 $Y2=0
cc_851 N_A_540_21#_c_1107_n N_A_1493_21#_c_1546_n 0.00101436f $X=9.405 $Y=2.047
+ $X2=0 $Y2=0
cc_852 N_A_540_21#_c_1107_n N_A_1493_21#_c_1535_n 0.00104244f $X=9.405 $Y=2.047
+ $X2=0 $Y2=0
cc_853 N_A_540_21#_c_1079_n N_A_1493_21#_c_1537_n 0.00528701f $X=11.18 $Y=1.245
+ $X2=0 $Y2=0
cc_854 N_A_540_21#_c_1081_n N_A_1493_21#_c_1537_n 0.0260128f $X=10.81 $Y=1.13
+ $X2=0 $Y2=0
cc_855 N_A_540_21#_c_1079_n N_A_1493_21#_c_1538_n 0.00284755f $X=11.18 $Y=1.245
+ $X2=0 $Y2=0
cc_856 N_A_540_21#_c_1079_n N_A_1493_21#_c_1539_n 0.0128122f $X=11.18 $Y=1.245
+ $X2=0 $Y2=0
cc_857 N_A_540_21#_c_1080_n N_A_1493_21#_c_1539_n 0.0492667f $X=11.265 $Y=2
+ $X2=0 $Y2=0
cc_858 N_A_540_21#_c_1081_n N_A_1493_21#_c_1539_n 0.00508536f $X=10.81 $Y=1.13
+ $X2=0 $Y2=0
cc_859 N_A_540_21#_c_1103_n N_A_1493_21#_c_1583_n 0.014897f $X=11.18 $Y=2.085
+ $X2=0 $Y2=0
cc_860 N_A_540_21#_c_1079_n N_A_1493_21#_c_1544_n 0.00892776f $X=11.18 $Y=1.245
+ $X2=0 $Y2=0
cc_861 N_A_540_21#_c_1081_n N_A_1493_21#_c_1544_n 0.00406959f $X=10.81 $Y=1.13
+ $X2=0 $Y2=0
cc_862 N_A_540_21#_c_1101_n N_SLEEP_B_M1010_g 0.0121053f $X=10.515 $Y=2.085
+ $X2=0 $Y2=0
cc_863 N_A_540_21#_c_1102_n N_SLEEP_B_M1010_g 0.00528139f $X=10.6 $Y=2.405 $X2=0
+ $Y2=0
cc_864 N_A_540_21#_c_1081_n N_SLEEP_B_M1010_g 0.0124866f $X=10.81 $Y=1.13 $X2=0
+ $Y2=0
cc_865 N_A_540_21#_c_1079_n N_SLEEP_B_M1002_g 0.00107413f $X=11.18 $Y=1.245
+ $X2=0 $Y2=0
cc_866 N_A_540_21#_c_1080_n N_SLEEP_B_M1002_g 6.36922e-19 $X=11.265 $Y=2 $X2=0
+ $Y2=0
cc_867 N_A_540_21#_c_1081_n N_SLEEP_B_M1002_g 2.85458e-19 $X=10.81 $Y=1.13 $X2=0
+ $Y2=0
cc_868 N_A_540_21#_c_1102_n N_CLK_M1015_g 0.00528139f $X=10.6 $Y=2.405 $X2=0
+ $Y2=0
cc_869 N_A_540_21#_c_1103_n N_CLK_M1015_g 0.0119501f $X=11.18 $Y=2.085 $X2=0
+ $Y2=0
cc_870 N_A_540_21#_c_1079_n N_CLK_M1013_g 0.0113745f $X=11.18 $Y=1.245 $X2=0
+ $Y2=0
cc_871 N_A_540_21#_c_1080_n N_CLK_M1013_g 0.00531226f $X=11.265 $Y=2 $X2=0 $Y2=0
cc_872 N_A_540_21#_c_1081_n N_CLK_M1013_g 0.00691782f $X=10.81 $Y=1.13 $X2=0
+ $Y2=0
cc_873 N_A_540_21#_c_1101_n CLK 0.0609839f $X=10.515 $Y=2.085 $X2=0 $Y2=0
cc_874 N_A_540_21#_c_1103_n CLK 0.0238828f $X=11.18 $Y=2.085 $X2=0 $Y2=0
cc_875 N_A_540_21#_c_1079_n CLK 0.00263029f $X=11.18 $Y=1.245 $X2=0 $Y2=0
cc_876 N_A_540_21#_c_1080_n CLK 0.0258604f $X=11.265 $Y=2 $X2=0 $Y2=0
cc_877 N_A_540_21#_c_1108_n CLK 0.0150178f $X=10.6 $Y=2.085 $X2=0 $Y2=0
cc_878 N_A_540_21#_c_1081_n CLK 0.0266002f $X=10.81 $Y=1.13 $X2=0 $Y2=0
cc_879 N_A_540_21#_c_1103_n N_CLK_c_1750_n 0.00781714f $X=11.18 $Y=2.085 $X2=0
+ $Y2=0
cc_880 N_A_540_21#_c_1079_n N_CLK_c_1750_n 0.00251917f $X=11.18 $Y=1.245 $X2=0
+ $Y2=0
cc_881 N_A_540_21#_c_1080_n N_CLK_c_1750_n 0.0160034f $X=11.265 $Y=2 $X2=0 $Y2=0
cc_882 N_A_540_21#_c_1081_n N_CLK_c_1750_n 0.00775699f $X=10.81 $Y=1.13 $X2=0
+ $Y2=0
cc_883 N_A_540_21#_M1027_g N_VPWR_c_1856_n 0.00194333f $X=3.075 $Y=2.705 $X2=0
+ $Y2=0
cc_884 N_A_540_21#_M1027_g N_VPWR_c_1857_n 0.00313972f $X=3.075 $Y=2.705 $X2=0
+ $Y2=0
cc_885 N_A_540_21#_M1022_g N_VPWR_c_1857_n 0.00383348f $X=4.975 $Y=2.86 $X2=0
+ $Y2=0
cc_886 N_A_540_21#_M1027_g N_VPWR_c_1854_n 0.00513578f $X=3.075 $Y=2.705 $X2=0
+ $Y2=0
cc_887 N_A_540_21#_M1022_g N_VPWR_c_1854_n 0.00460802f $X=4.975 $Y=2.86 $X2=0
+ $Y2=0
cc_888 N_A_540_21#_M1025_g N_A_282_477#_c_1996_n 8.90508e-19 $X=2.775 $Y=0.445
+ $X2=0 $Y2=0
cc_889 N_A_540_21#_c_1069_n N_A_282_477#_c_1997_n 0.00180231f $X=2.975 $Y=1.765
+ $X2=0 $Y2=0
cc_890 N_A_540_21#_c_1075_n N_A_282_477#_c_1997_n 0.00865889f $X=2.975 $Y=0.9
+ $X2=0 $Y2=0
cc_891 N_A_540_21#_c_1069_n N_A_282_477#_c_1999_n 0.00649709f $X=2.975 $Y=1.765
+ $X2=0 $Y2=0
cc_892 N_A_540_21#_M1027_g N_A_282_477#_c_1999_n 0.00317906f $X=3.075 $Y=2.705
+ $X2=0 $Y2=0
cc_893 N_A_540_21#_M1027_g N_A_282_477#_c_2053_n 0.00534066f $X=3.075 $Y=2.705
+ $X2=0 $Y2=0
cc_894 N_A_540_21#_M1027_g N_A_282_477#_c_2007_n 0.0134823f $X=3.075 $Y=2.705
+ $X2=0 $Y2=0
cc_895 N_A_540_21#_c_1069_n N_A_282_477#_c_2000_n 0.00289628f $X=2.975 $Y=1.765
+ $X2=0 $Y2=0
cc_896 N_A_540_21#_M1027_g N_A_282_477#_c_2000_n 6.02528e-19 $X=3.075 $Y=2.705
+ $X2=0 $Y2=0
cc_897 N_A_540_21#_c_1085_n N_A_282_477#_c_2000_n 0.0089591f $X=3.78 $Y=1.84
+ $X2=0 $Y2=0
cc_898 N_A_540_21#_M1005_g N_A_282_477#_c_2000_n 0.0176702f $X=3.855 $Y=0.905
+ $X2=0 $Y2=0
cc_899 N_A_540_21#_c_1096_n N_A_282_477#_c_2000_n 0.00527111f $X=3.855 $Y=1.857
+ $X2=0 $Y2=0
cc_900 N_A_540_21#_c_1087_n N_A_282_477#_c_2010_n 0.0029378f $X=4.9 $Y=1.875
+ $X2=0 $Y2=0
cc_901 N_A_540_21#_M1022_g N_A_282_477#_c_2010_n 7.07726e-19 $X=4.975 $Y=2.86
+ $X2=0 $Y2=0
cc_902 N_A_540_21#_c_1096_n N_A_282_477#_c_2010_n 0.0054437f $X=3.855 $Y=1.857
+ $X2=0 $Y2=0
cc_903 N_A_540_21#_M1027_g N_A_282_477#_c_2011_n 5.32675e-19 $X=3.075 $Y=2.705
+ $X2=0 $Y2=0
cc_904 N_A_540_21#_M1022_g N_A_282_477#_c_2012_n 6.92234e-19 $X=4.975 $Y=2.86
+ $X2=0 $Y2=0
cc_905 N_A_540_21#_M1027_g N_A_282_477#_c_2013_n 0.00193912f $X=3.075 $Y=2.705
+ $X2=0 $Y2=0
cc_906 N_A_540_21#_c_1095_n N_A_282_477#_c_2013_n 0.00291312f $X=3.025 $Y=1.84
+ $X2=0 $Y2=0
cc_907 N_A_540_21#_c_1085_n N_A_282_477#_c_2002_n 0.0037361f $X=3.78 $Y=1.84
+ $X2=0 $Y2=0
cc_908 N_A_540_21#_M1005_g N_A_282_477#_c_2002_n 0.00460697f $X=3.855 $Y=0.905
+ $X2=0 $Y2=0
cc_909 N_A_540_21#_c_1075_n N_A_282_477#_c_2002_n 0.00165565f $X=2.975 $Y=0.9
+ $X2=0 $Y2=0
cc_910 N_A_540_21#_c_1101_n A_1858_419# 6.98275e-19 $X=10.515 $Y=2.085 $X2=-0.19
+ $Y2=-0.245
cc_911 N_A_540_21#_c_1107_n A_1858_419# 6.11325e-19 $X=9.405 $Y=2.047 $X2=-0.19
+ $Y2=-0.245
cc_912 N_A_540_21#_c_1101_n N_KAPWR_M1017_d 0.00307194f $X=10.515 $Y=2.085
+ $X2=-0.19 $Y2=-0.245
cc_913 N_A_540_21#_c_1103_n N_KAPWR_M1015_d 0.00400127f $X=11.18 $Y=2.085 $X2=0
+ $Y2=0
cc_914 N_A_540_21#_M1010_d N_KAPWR_c_2164_n 0.00425678f $X=10.325 $Y=2.095 $X2=0
+ $Y2=0
cc_915 N_A_540_21#_M1027_g N_KAPWR_c_2164_n 0.00717829f $X=3.075 $Y=2.705 $X2=0
+ $Y2=0
cc_916 N_A_540_21#_M1022_g N_KAPWR_c_2164_n 0.00163688f $X=4.975 $Y=2.86 $X2=0
+ $Y2=0
cc_917 N_A_540_21#_c_1091_n N_KAPWR_c_2164_n 0.00945542f $X=6.785 $Y=1.785 $X2=0
+ $Y2=0
cc_918 N_A_540_21#_c_1093_n N_KAPWR_c_2164_n 0.00856204f $X=7.145 $Y=1.785 $X2=0
+ $Y2=0
cc_919 N_A_540_21#_c_1101_n N_KAPWR_c_2164_n 0.00652937f $X=10.515 $Y=2.085
+ $X2=0 $Y2=0
cc_920 N_A_540_21#_c_1102_n N_KAPWR_c_2164_n 0.0133164f $X=10.6 $Y=2.405 $X2=0
+ $Y2=0
cc_921 N_A_540_21#_c_1103_n N_KAPWR_c_2164_n 0.00652937f $X=11.18 $Y=2.085 $X2=0
+ $Y2=0
cc_922 N_A_540_21#_c_1106_n N_KAPWR_c_2164_n 0.0019668f $X=9.235 $Y=2.047 $X2=0
+ $Y2=0
cc_923 N_A_540_21#_M1025_g N_VGND_c_2306_n 0.00304304f $X=2.775 $Y=0.445 $X2=0
+ $Y2=0
cc_924 N_A_540_21#_M1025_g N_VGND_c_2317_n 0.00547467f $X=2.775 $Y=0.445 $X2=0
+ $Y2=0
cc_925 N_A_540_21#_M1025_g N_VGND_c_2320_n 0.0108841f $X=2.775 $Y=0.445 $X2=0
+ $Y2=0
cc_926 N_A_540_21#_c_1079_n A_2243_178# 0.00210406f $X=11.18 $Y=1.245 $X2=-0.19
+ $Y2=-0.245
cc_927 N_A_1319_69#_c_1340_n N_A_1493_21#_M1029_d 0.0107826f $X=12.43 $Y=2.91
+ $X2=0 $Y2=0
cc_928 N_A_1319_69#_c_1323_n N_A_1493_21#_M1019_g 2.367e-19 $X=8.55 $Y=1.51
+ $X2=0 $Y2=0
cc_929 N_A_1319_69#_c_1359_n N_A_1493_21#_M1019_g 3.25444e-19 $X=7.125 $Y=0.76
+ $X2=0 $Y2=0
cc_930 N_A_1319_69#_M1020_g N_A_1493_21#_M1006_g 0.011623f $X=8.445 $Y=0.835
+ $X2=0 $Y2=0
cc_931 N_A_1319_69#_c_1323_n N_A_1493_21#_M1006_g 3.98653e-19 $X=8.55 $Y=1.51
+ $X2=0 $Y2=0
cc_932 N_A_1319_69#_M1020_g N_A_1493_21#_c_1532_n 0.00907339f $X=8.445 $Y=0.835
+ $X2=0 $Y2=0
cc_933 N_A_1319_69#_M1007_g N_A_1493_21#_c_1532_n 0.00907339f $X=8.805 $Y=0.835
+ $X2=0 $Y2=0
cc_934 N_A_1319_69#_M1007_g N_A_1493_21#_c_1533_n 0.00934585f $X=8.805 $Y=0.835
+ $X2=0 $Y2=0
cc_935 N_A_1319_69#_c_1358_n N_A_1493_21#_c_1546_n 0.0154247f $X=10.175 $Y=2.425
+ $X2=0 $Y2=0
cc_936 N_A_1319_69#_c_1336_n N_A_1493_21#_c_1546_n 0.00106365f $X=10.26 $Y=2.905
+ $X2=0 $Y2=0
cc_937 N_A_1319_69#_c_1338_n N_A_1493_21#_c_1546_n 3.12331e-19 $X=10.345 $Y=2.99
+ $X2=0 $Y2=0
cc_938 N_A_1319_69#_c_1344_n N_A_1493_21#_c_1546_n 0.00222472f $X=8.9 $Y=2.43
+ $X2=0 $Y2=0
cc_939 N_A_1319_69#_c_1326_n N_A_1493_21#_c_1539_n 3.96587e-19 $X=11.545
+ $Y=1.985 $X2=0 $Y2=0
cc_940 N_A_1319_69#_c_1327_n N_A_1493_21#_c_1539_n 0.00734115f $X=12.265 $Y=1.91
+ $X2=0 $Y2=0
cc_941 N_A_1319_69#_c_1328_n N_A_1493_21#_c_1539_n 0.00616348f $X=11.67 $Y=1.91
+ $X2=0 $Y2=0
cc_942 N_A_1319_69#_c_1318_n N_A_1493_21#_c_1539_n 0.00603977f $X=12.34 $Y=1.65
+ $X2=0 $Y2=0
cc_943 N_A_1319_69#_c_1345_n N_A_1493_21#_c_1539_n 2.03474e-19 $X=12.43 $Y=2.745
+ $X2=0 $Y2=0
cc_944 N_A_1319_69#_c_1327_n N_A_1493_21#_c_1549_n 0.0149438f $X=12.265 $Y=1.91
+ $X2=0 $Y2=0
cc_945 N_A_1319_69#_c_1340_n N_A_1493_21#_c_1549_n 0.00244802f $X=12.43 $Y=2.91
+ $X2=0 $Y2=0
cc_946 N_A_1319_69#_c_1345_n N_A_1493_21#_c_1549_n 0.00221043f $X=12.43 $Y=2.745
+ $X2=0 $Y2=0
cc_947 N_A_1319_69#_c_1326_n N_A_1493_21#_c_1583_n 0.00878936f $X=11.545
+ $Y=1.985 $X2=0 $Y2=0
cc_948 N_A_1319_69#_c_1401_n N_A_1493_21#_c_1583_n 0.0120334f $X=11.535 $Y=2.425
+ $X2=0 $Y2=0
cc_949 N_A_1319_69#_c_1326_n N_A_1493_21#_c_1550_n 0.00511894f $X=11.545
+ $Y=1.985 $X2=0 $Y2=0
cc_950 N_A_1319_69#_c_1340_n N_A_1493_21#_c_1550_n 0.0173211f $X=12.43 $Y=2.91
+ $X2=0 $Y2=0
cc_951 N_A_1319_69#_c_1345_n N_A_1493_21#_c_1550_n 0.00593971f $X=12.43 $Y=2.745
+ $X2=0 $Y2=0
cc_952 N_A_1319_69#_M1007_g N_A_1493_21#_c_1540_n 0.00929831f $X=8.805 $Y=0.835
+ $X2=0 $Y2=0
cc_953 N_A_1319_69#_M1007_g N_A_1493_21#_c_1545_n 0.00257227f $X=8.805 $Y=0.835
+ $X2=0 $Y2=0
cc_954 N_A_1319_69#_c_1358_n N_SLEEP_B_M1010_g 0.00859173f $X=10.175 $Y=2.425
+ $X2=0 $Y2=0
cc_955 N_A_1319_69#_c_1336_n N_SLEEP_B_M1010_g 0.0131929f $X=10.26 $Y=2.905
+ $X2=0 $Y2=0
cc_956 N_A_1319_69#_c_1339_n N_SLEEP_B_M1010_g 3.40635e-19 $X=10.94 $Y=2.905
+ $X2=0 $Y2=0
cc_957 N_A_1319_69#_c_1328_n N_SLEEP_B_M1002_g 0.00551877f $X=11.67 $Y=1.91
+ $X2=0 $Y2=0
cc_958 N_A_1319_69#_c_1327_n N_SLEEP_B_c_1684_n 0.00906292f $X=12.265 $Y=1.91
+ $X2=0 $Y2=0
cc_959 N_A_1319_69#_c_1318_n N_SLEEP_B_c_1684_n 8.93998e-19 $X=12.34 $Y=1.65
+ $X2=0 $Y2=0
cc_960 N_A_1319_69#_c_1328_n N_CLK_M1015_g 0.0274148f $X=11.67 $Y=1.91 $X2=0
+ $Y2=0
cc_961 N_A_1319_69#_c_1336_n N_CLK_M1015_g 3.40635e-19 $X=10.26 $Y=2.905 $X2=0
+ $Y2=0
cc_962 N_A_1319_69#_c_1339_n N_CLK_M1015_g 0.0127487f $X=10.94 $Y=2.905 $X2=0
+ $Y2=0
cc_963 N_A_1319_69#_c_1402_n N_CLK_M1015_g 0.00856139f $X=11.025 $Y=2.425 $X2=0
+ $Y2=0
cc_964 N_A_1319_69#_c_1448_p N_CLK_M1015_g 5.47824e-19 $X=11.62 $Y=2.745 $X2=0
+ $Y2=0
cc_965 N_A_1319_69#_c_1315_n N_A_2504_57#_M1031_g 0.00585127f $X=12.85 $Y=1.575
+ $X2=0 $Y2=0
cc_966 N_A_1319_69#_M1032_g N_A_2504_57#_M1031_g 0.0139382f $X=12.88 $Y=0.495
+ $X2=0 $Y2=0
cc_967 N_A_1319_69#_c_1320_n N_A_2504_57#_M1024_g 0.0153393f $X=12.865 $Y=1.65
+ $X2=0 $Y2=0
cc_968 N_A_1319_69#_c_1315_n N_A_2504_57#_c_1799_n 0.0094645f $X=12.85 $Y=1.575
+ $X2=0 $Y2=0
cc_969 N_A_1319_69#_M1032_g N_A_2504_57#_c_1799_n 0.0131268f $X=12.88 $Y=0.495
+ $X2=0 $Y2=0
cc_970 N_A_1319_69#_c_1319_n N_A_2504_57#_c_1799_n 0.00580594f $X=12.865
+ $Y=1.075 $X2=0 $Y2=0
cc_971 N_A_1319_69#_c_1314_n N_A_2504_57#_c_1804_n 0.0104477f $X=12.775 $Y=1.65
+ $X2=0 $Y2=0
cc_972 N_A_1319_69#_c_1330_n N_A_2504_57#_c_1804_n 0.0115158f $X=12.88 $Y=1.725
+ $X2=0 $Y2=0
cc_973 N_A_1319_69#_c_1318_n N_A_2504_57#_c_1804_n 0.013513f $X=12.34 $Y=1.65
+ $X2=0 $Y2=0
cc_974 N_A_1319_69#_c_1320_n N_A_2504_57#_c_1804_n 0.0018089f $X=12.865 $Y=1.65
+ $X2=0 $Y2=0
cc_975 N_A_1319_69#_c_1340_n N_A_2504_57#_c_1804_n 0.00428806f $X=12.43 $Y=2.91
+ $X2=0 $Y2=0
cc_976 N_A_1319_69#_c_1341_n N_A_2504_57#_c_1804_n 0.00156195f $X=12.43 $Y=2.91
+ $X2=0 $Y2=0
cc_977 N_A_1319_69#_c_1315_n N_A_2504_57#_c_1800_n 0.00939885f $X=12.85 $Y=1.575
+ $X2=0 $Y2=0
cc_978 N_A_1319_69#_c_1319_n N_A_2504_57#_c_1800_n 7.69146e-19 $X=12.865
+ $Y=1.075 $X2=0 $Y2=0
cc_979 N_A_1319_69#_c_1320_n N_A_2504_57#_c_1800_n 0.00777516f $X=12.865 $Y=1.65
+ $X2=0 $Y2=0
cc_980 N_A_1319_69#_c_1315_n N_A_2504_57#_c_1801_n 0.0142245f $X=12.85 $Y=1.575
+ $X2=0 $Y2=0
cc_981 N_A_1319_69#_c_1320_n N_A_2504_57#_c_1801_n 0.00457333f $X=12.865 $Y=1.65
+ $X2=0 $Y2=0
cc_982 N_A_1319_69#_c_1314_n N_A_2504_57#_c_1802_n 0.0111895f $X=12.775 $Y=1.65
+ $X2=0 $Y2=0
cc_983 N_A_1319_69#_c_1315_n N_A_2504_57#_c_1802_n 0.00645076f $X=12.85 $Y=1.575
+ $X2=0 $Y2=0
cc_984 N_A_1319_69#_c_1320_n N_A_2504_57#_c_1802_n 3.62533e-19 $X=12.865 $Y=1.65
+ $X2=0 $Y2=0
cc_985 N_A_1319_69#_c_1330_n N_VPWR_c_1858_n 0.00881619f $X=12.88 $Y=1.725 $X2=0
+ $Y2=0
cc_986 N_A_1319_69#_c_1340_n N_VPWR_c_1858_n 0.009564f $X=12.43 $Y=2.91 $X2=0
+ $Y2=0
cc_987 N_A_1319_69#_c_1341_n N_VPWR_c_1858_n 0.00168289f $X=12.43 $Y=2.91 $X2=0
+ $Y2=0
cc_988 N_A_1319_69#_c_1345_n N_VPWR_c_1858_n 0.0026375f $X=12.43 $Y=2.745 $X2=0
+ $Y2=0
cc_989 N_A_1319_69#_c_1326_n N_VPWR_c_1861_n 0.00770696f $X=11.545 $Y=1.985
+ $X2=0 $Y2=0
cc_990 N_A_1319_69#_c_1330_n N_VPWR_c_1861_n 0.00312414f $X=12.88 $Y=1.725 $X2=0
+ $Y2=0
cc_991 N_A_1319_69#_c_1337_n N_VPWR_c_1861_n 0.0449818f $X=10.855 $Y=2.99 $X2=0
+ $Y2=0
cc_992 N_A_1319_69#_c_1338_n N_VPWR_c_1861_n 0.0121867f $X=10.345 $Y=2.99 $X2=0
+ $Y2=0
cc_993 N_A_1319_69#_c_1477_p N_VPWR_c_1861_n 0.0104451f $X=11.705 $Y=2.91 $X2=0
+ $Y2=0
cc_994 N_A_1319_69#_c_1340_n N_VPWR_c_1861_n 0.0578702f $X=12.43 $Y=2.91 $X2=0
+ $Y2=0
cc_995 N_A_1319_69#_c_1341_n N_VPWR_c_1861_n 0.00783549f $X=12.43 $Y=2.91 $X2=0
+ $Y2=0
cc_996 N_A_1319_69#_c_1344_n N_VPWR_c_1861_n 0.0210192f $X=8.9 $Y=2.43 $X2=0
+ $Y2=0
cc_997 N_A_1319_69#_M1001_s N_VPWR_c_1854_n 0.00119401f $X=8.755 $Y=2.095 $X2=0
+ $Y2=0
cc_998 N_A_1319_69#_c_1326_n N_VPWR_c_1854_n 0.00998876f $X=11.545 $Y=1.985
+ $X2=0 $Y2=0
cc_999 N_A_1319_69#_c_1337_n N_VPWR_c_1854_n 0.00574275f $X=10.855 $Y=2.99 $X2=0
+ $Y2=0
cc_1000 N_A_1319_69#_c_1338_n N_VPWR_c_1854_n 0.0015975f $X=10.345 $Y=2.99 $X2=0
+ $Y2=0
cc_1001 N_A_1319_69#_c_1477_p N_VPWR_c_1854_n 0.00145179f $X=11.705 $Y=2.91
+ $X2=0 $Y2=0
cc_1002 N_A_1319_69#_c_1340_n N_VPWR_c_1854_n 0.00755029f $X=12.43 $Y=2.91 $X2=0
+ $Y2=0
cc_1003 N_A_1319_69#_c_1341_n N_VPWR_c_1854_n 0.00625434f $X=12.43 $Y=2.91 $X2=0
+ $Y2=0
cc_1004 N_A_1319_69#_c_1344_n N_VPWR_c_1854_n 0.00303861f $X=8.9 $Y=2.43 $X2=0
+ $Y2=0
cc_1005 N_A_1319_69#_c_1358_n A_1858_419# 0.00290533f $X=10.175 $Y=2.425
+ $X2=-0.19 $Y2=-0.245
cc_1006 N_A_1319_69#_c_1358_n N_KAPWR_M1017_d 0.00640065f $X=10.175 $Y=2.425
+ $X2=-0.19 $Y2=-0.245
cc_1007 N_A_1319_69#_c_1401_n N_KAPWR_M1015_d 0.00675338f $X=11.535 $Y=2.425
+ $X2=0 $Y2=0
cc_1008 N_A_1319_69#_c_1358_n N_KAPWR_c_2176_n 0.0151698f $X=10.175 $Y=2.425
+ $X2=0 $Y2=0
cc_1009 N_A_1319_69#_c_1336_n N_KAPWR_c_2176_n 0.0152291f $X=10.26 $Y=2.905
+ $X2=0 $Y2=0
cc_1010 N_A_1319_69#_c_1338_n N_KAPWR_c_2176_n 0.0140409f $X=10.345 $Y=2.99
+ $X2=0 $Y2=0
cc_1011 N_A_1319_69#_c_1344_n N_KAPWR_c_2176_n 0.00537831f $X=8.9 $Y=2.43 $X2=0
+ $Y2=0
cc_1012 N_A_1319_69#_c_1326_n N_KAPWR_c_2214_n 4.19303e-19 $X=11.545 $Y=1.985
+ $X2=0 $Y2=0
cc_1013 N_A_1319_69#_c_1337_n N_KAPWR_c_2214_n 0.0136755f $X=10.855 $Y=2.99
+ $X2=0 $Y2=0
cc_1014 N_A_1319_69#_c_1339_n N_KAPWR_c_2214_n 0.0151292f $X=10.94 $Y=2.905
+ $X2=0 $Y2=0
cc_1015 N_A_1319_69#_c_1401_n N_KAPWR_c_2214_n 0.0108529f $X=11.535 $Y=2.425
+ $X2=0 $Y2=0
cc_1016 N_A_1319_69#_c_1448_p N_KAPWR_c_2214_n 0.00322291f $X=11.62 $Y=2.745
+ $X2=0 $Y2=0
cc_1017 N_A_1319_69#_c_1477_p N_KAPWR_c_2214_n 0.0156321f $X=11.705 $Y=2.91
+ $X2=0 $Y2=0
cc_1018 N_A_1319_69#_c_1326_n N_KAPWR_c_2164_n 0.0018092f $X=11.545 $Y=1.985
+ $X2=0 $Y2=0
cc_1019 N_A_1319_69#_c_1330_n N_KAPWR_c_2164_n 0.00480838f $X=12.88 $Y=1.725
+ $X2=0 $Y2=0
cc_1020 N_A_1319_69#_c_1334_n N_KAPWR_c_2164_n 0.0416403f $X=8.735 $Y=2.35 $X2=0
+ $Y2=0
cc_1021 N_A_1319_69#_c_1335_n N_KAPWR_c_2164_n 0.0272675f $X=7.525 $Y=2.35 $X2=0
+ $Y2=0
cc_1022 N_A_1319_69#_c_1358_n N_KAPWR_c_2164_n 0.0448732f $X=10.175 $Y=2.425
+ $X2=0 $Y2=0
cc_1023 N_A_1319_69#_c_1336_n N_KAPWR_c_2164_n 0.014022f $X=10.26 $Y=2.905 $X2=0
+ $Y2=0
cc_1024 N_A_1319_69#_c_1337_n N_KAPWR_c_2164_n 0.0203156f $X=10.855 $Y=2.99
+ $X2=0 $Y2=0
cc_1025 N_A_1319_69#_c_1338_n N_KAPWR_c_2164_n 0.00253087f $X=10.345 $Y=2.99
+ $X2=0 $Y2=0
cc_1026 N_A_1319_69#_c_1339_n N_KAPWR_c_2164_n 0.0139877f $X=10.94 $Y=2.905
+ $X2=0 $Y2=0
cc_1027 N_A_1319_69#_c_1401_n N_KAPWR_c_2164_n 0.0204638f $X=11.535 $Y=2.425
+ $X2=0 $Y2=0
cc_1028 N_A_1319_69#_c_1448_p N_KAPWR_c_2164_n 0.00743295f $X=11.62 $Y=2.745
+ $X2=0 $Y2=0
cc_1029 N_A_1319_69#_c_1477_p N_KAPWR_c_2164_n 0.00705435f $X=11.705 $Y=2.91
+ $X2=0 $Y2=0
cc_1030 N_A_1319_69#_c_1340_n N_KAPWR_c_2164_n 0.0410287f $X=12.43 $Y=2.91 $X2=0
+ $Y2=0
cc_1031 N_A_1319_69#_c_1341_n N_KAPWR_c_2164_n 0.00491829f $X=12.43 $Y=2.91
+ $X2=0 $Y2=0
cc_1032 N_A_1319_69#_c_1344_n N_KAPWR_c_2164_n 0.0318014f $X=8.9 $Y=2.43 $X2=0
+ $Y2=0
cc_1033 N_A_1319_69#_c_1345_n N_KAPWR_c_2164_n 0.00841226f $X=12.43 $Y=2.745
+ $X2=0 $Y2=0
cc_1034 N_A_1319_69#_M1020_g N_VGND_c_2308_n 0.0114696f $X=8.445 $Y=0.835 $X2=0
+ $Y2=0
cc_1035 N_A_1319_69#_c_1327_n N_VGND_c_2309_n 0.00631373f $X=12.265 $Y=1.91
+ $X2=0 $Y2=0
cc_1036 N_A_1319_69#_M1032_g N_VGND_c_2309_n 0.00346692f $X=12.88 $Y=0.495 $X2=0
+ $Y2=0
cc_1037 N_A_1319_69#_c_1319_n N_VGND_c_2309_n 0.00163265f $X=12.865 $Y=1.075
+ $X2=0 $Y2=0
cc_1038 N_A_1319_69#_c_1315_n N_VGND_c_2310_n 5.94772e-19 $X=12.85 $Y=1.575
+ $X2=0 $Y2=0
cc_1039 N_A_1319_69#_M1032_g N_VGND_c_2310_n 0.00953123f $X=12.88 $Y=0.495 $X2=0
+ $Y2=0
cc_1040 N_A_1319_69#_M1032_g N_VGND_c_2318_n 0.00502664f $X=12.88 $Y=0.495 $X2=0
+ $Y2=0
cc_1041 N_A_1319_69#_M1020_g N_VGND_c_2320_n 9.49986e-19 $X=8.445 $Y=0.835 $X2=0
+ $Y2=0
cc_1042 N_A_1319_69#_M1007_g N_VGND_c_2320_n 9.49986e-19 $X=8.805 $Y=0.835 $X2=0
+ $Y2=0
cc_1043 N_A_1319_69#_M1032_g N_VGND_c_2320_n 0.0106059f $X=12.88 $Y=0.495 $X2=0
+ $Y2=0
cc_1044 N_A_1493_21#_c_1533_n N_SLEEP_B_M1010_g 0.00421284f $X=9.43 $Y=0.79
+ $X2=0 $Y2=0
cc_1045 N_A_1493_21#_c_1535_n N_SLEEP_B_M1010_g 0.0546137f $X=9.655 $Y=1.965
+ $X2=0 $Y2=0
cc_1046 N_A_1493_21#_c_1536_n N_SLEEP_B_M1010_g 0.0107943f $X=10.305 $Y=0.83
+ $X2=0 $Y2=0
cc_1047 N_A_1493_21#_c_1537_n N_SLEEP_B_M1010_g 9.02832e-19 $X=11.145 $Y=0.68
+ $X2=0 $Y2=0
cc_1048 N_A_1493_21#_c_1542_n N_SLEEP_B_M1010_g 0.00130768f $X=9.92 $Y=0.932
+ $X2=0 $Y2=0
cc_1049 N_A_1493_21#_c_1543_n N_SLEEP_B_M1010_g 0.0131683f $X=10.39 $Y=0.68
+ $X2=0 $Y2=0
cc_1050 N_A_1493_21#_c_1545_n N_SLEEP_B_M1010_g 0.0159881f $X=9.705 $Y=0.955
+ $X2=0 $Y2=0
cc_1051 N_A_1493_21#_c_1538_n N_SLEEP_B_M1002_g 0.00931478f $X=11.52 $Y=0.905
+ $X2=0 $Y2=0
cc_1052 N_A_1493_21#_c_1539_n N_SLEEP_B_M1002_g 0.0106555f $X=11.605 $Y=2 $X2=0
+ $Y2=0
cc_1053 N_A_1493_21#_c_1538_n N_SLEEP_B_c_1684_n 0.00136906f $X=11.52 $Y=0.905
+ $X2=0 $Y2=0
cc_1054 N_A_1493_21#_c_1539_n N_SLEEP_B_c_1684_n 0.008638f $X=11.605 $Y=2 $X2=0
+ $Y2=0
cc_1055 N_A_1493_21#_c_1544_n N_SLEEP_B_c_1684_n 2.4946e-19 $X=11.23 $Y=0.68
+ $X2=0 $Y2=0
cc_1056 N_A_1493_21#_c_1532_n N_SLEEP_B_c_1685_n 0.0128286f $X=9.355 $Y=0.18
+ $X2=0 $Y2=0
cc_1057 N_A_1493_21#_c_1542_n N_SLEEP_B_c_1685_n 0.00645963f $X=9.92 $Y=0.932
+ $X2=0 $Y2=0
cc_1058 N_A_1493_21#_c_1545_n N_SLEEP_B_c_1685_n 0.00718371f $X=9.705 $Y=0.955
+ $X2=0 $Y2=0
cc_1059 N_A_1493_21#_c_1536_n N_SLEEP_B_c_1686_n 0.00617561f $X=10.305 $Y=0.83
+ $X2=0 $Y2=0
cc_1060 N_A_1493_21#_c_1537_n N_SLEEP_B_c_1686_n 0.0474754f $X=11.145 $Y=0.68
+ $X2=0 $Y2=0
cc_1061 N_A_1493_21#_c_1538_n N_SLEEP_B_c_1686_n 0.00696688f $X=11.52 $Y=0.905
+ $X2=0 $Y2=0
cc_1062 N_A_1493_21#_c_1543_n N_SLEEP_B_c_1686_n 0.0123916f $X=10.39 $Y=0.68
+ $X2=0 $Y2=0
cc_1063 N_A_1493_21#_c_1544_n N_SLEEP_B_c_1686_n 0.0127302f $X=11.23 $Y=0.68
+ $X2=0 $Y2=0
cc_1064 N_A_1493_21#_c_1533_n N_SLEEP_B_c_1687_n 0.0019553f $X=9.43 $Y=0.79
+ $X2=0 $Y2=0
cc_1065 N_A_1493_21#_c_1542_n N_SLEEP_B_c_1687_n 0.0243417f $X=9.92 $Y=0.932
+ $X2=0 $Y2=0
cc_1066 N_A_1493_21#_c_1544_n N_SLEEP_B_c_1688_n 0.0065751f $X=11.23 $Y=0.68
+ $X2=0 $Y2=0
cc_1067 N_A_1493_21#_c_1538_n N_SLEEP_B_c_1689_n 0.0137308f $X=11.52 $Y=0.905
+ $X2=0 $Y2=0
cc_1068 N_A_1493_21#_c_1544_n N_SLEEP_B_c_1689_n 0.00359117f $X=11.23 $Y=0.68
+ $X2=0 $Y2=0
cc_1069 N_A_1493_21#_c_1537_n N_CLK_M1013_g 0.00318151f $X=11.145 $Y=0.68 $X2=0
+ $Y2=0
cc_1070 N_A_1493_21#_c_1538_n N_CLK_M1013_g 2.09135e-19 $X=11.52 $Y=0.905 $X2=0
+ $Y2=0
cc_1071 N_A_1493_21#_c_1539_n N_CLK_M1013_g 0.00125649f $X=11.605 $Y=2 $X2=0
+ $Y2=0
cc_1072 N_A_1493_21#_c_1543_n N_CLK_M1013_g 0.00217799f $X=10.39 $Y=0.68 $X2=0
+ $Y2=0
cc_1073 N_A_1493_21#_c_1544_n N_CLK_M1013_g 0.00887359f $X=11.23 $Y=0.68 $X2=0
+ $Y2=0
cc_1074 N_A_1493_21#_c_1535_n CLK 0.0128156f $X=9.655 $Y=1.965 $X2=0 $Y2=0
cc_1075 N_A_1493_21#_c_1536_n CLK 0.0119014f $X=10.305 $Y=0.83 $X2=0 $Y2=0
cc_1076 N_A_1493_21#_c_1542_n CLK 0.00832895f $X=9.92 $Y=0.932 $X2=0 $Y2=0
cc_1077 N_A_1493_21#_c_1543_n CLK 0.00576953f $X=10.39 $Y=0.68 $X2=0 $Y2=0
cc_1078 N_A_1493_21#_c_1545_n CLK 0.00276564f $X=9.705 $Y=0.955 $X2=0 $Y2=0
cc_1079 N_A_1493_21#_c_1537_n N_CLK_c_1750_n 4.57092e-19 $X=11.145 $Y=0.68 $X2=0
+ $Y2=0
cc_1080 N_A_1493_21#_c_1549_n N_A_2504_57#_c_1804_n 0.00856903f $X=11.875
+ $Y=2.085 $X2=0 $Y2=0
cc_1081 N_A_1493_21#_c_1550_n N_A_2504_57#_c_1804_n 0.0152551f $X=11.96 $Y=2.325
+ $X2=0 $Y2=0
cc_1082 N_A_1493_21#_c_1546_n N_VPWR_c_1861_n 0.00892222f $X=9.655 $Y=2.09 $X2=0
+ $Y2=0
cc_1083 N_A_1493_21#_M1029_d N_VPWR_c_1854_n 0.00186062f $X=11.67 $Y=2.095 $X2=0
+ $Y2=0
cc_1084 N_A_1493_21#_c_1546_n N_VPWR_c_1854_n 0.00865691f $X=9.655 $Y=2.09 $X2=0
+ $Y2=0
cc_1085 N_A_1493_21#_c_1546_n N_KAPWR_c_2176_n 0.00900644f $X=9.655 $Y=2.09
+ $X2=0 $Y2=0
cc_1086 N_A_1493_21#_M1029_d N_KAPWR_c_2164_n 0.00393414f $X=11.67 $Y=2.095
+ $X2=0 $Y2=0
cc_1087 N_A_1493_21#_c_1546_n N_KAPWR_c_2164_n 0.00618057f $X=9.655 $Y=2.09
+ $X2=0 $Y2=0
cc_1088 N_A_1493_21#_c_1549_n N_KAPWR_c_2164_n 0.00398295f $X=11.875 $Y=2.085
+ $X2=0 $Y2=0
cc_1089 N_A_1493_21#_c_1583_n N_KAPWR_c_2164_n 6.47155e-19 $X=11.69 $Y=2.085
+ $X2=0 $Y2=0
cc_1090 N_A_1493_21#_c_1550_n N_KAPWR_c_2164_n 0.00780915f $X=11.96 $Y=2.325
+ $X2=0 $Y2=0
cc_1091 N_A_1493_21#_M1019_g N_VGND_c_2308_n 5.0787e-19 $X=7.54 $Y=0.775 $X2=0
+ $Y2=0
cc_1092 N_A_1493_21#_M1006_g N_VGND_c_2308_n 0.0126459f $X=7.9 $Y=0.775 $X2=0
+ $Y2=0
cc_1093 N_A_1493_21#_c_1532_n N_VGND_c_2308_n 0.0186723f $X=9.355 $Y=0.18 $X2=0
+ $Y2=0
cc_1094 N_A_1493_21#_c_1534_n N_VGND_c_2308_n 0.00442488f $X=7.9 $Y=0.18 $X2=0
+ $Y2=0
cc_1095 N_A_1493_21#_c_1538_n N_VGND_c_2309_n 0.0061366f $X=11.52 $Y=0.905 $X2=0
+ $Y2=0
cc_1096 N_A_1493_21#_c_1539_n N_VGND_c_2309_n 0.00806148f $X=11.605 $Y=2 $X2=0
+ $Y2=0
cc_1097 N_A_1493_21#_c_1549_n N_VGND_c_2309_n 0.00362475f $X=11.875 $Y=2.085
+ $X2=0 $Y2=0
cc_1098 N_A_1493_21#_c_1530_n N_VGND_c_2311_n 0.0139733f $X=7.615 $Y=0.18 $X2=0
+ $Y2=0
cc_1099 N_A_1493_21#_c_1532_n N_VGND_c_2313_n 0.0384433f $X=9.355 $Y=0.18 $X2=0
+ $Y2=0
cc_1100 N_A_1493_21#_c_1540_n N_VGND_c_2313_n 0.00700261f $X=9.135 $Y=0.75 $X2=0
+ $Y2=0
cc_1101 N_A_1493_21#_c_1541_n N_VGND_c_2313_n 0.00730889f $X=9.59 $Y=0.932 $X2=0
+ $Y2=0
cc_1102 N_A_1493_21#_c_1529_n N_VGND_c_2320_n 0.00673026f $X=7.825 $Y=0.18 $X2=0
+ $Y2=0
cc_1103 N_A_1493_21#_c_1530_n N_VGND_c_2320_n 0.00604505f $X=7.615 $Y=0.18 $X2=0
+ $Y2=0
cc_1104 N_A_1493_21#_c_1532_n N_VGND_c_2320_n 0.0481416f $X=9.355 $Y=0.18 $X2=0
+ $Y2=0
cc_1105 N_A_1493_21#_c_1534_n N_VGND_c_2320_n 0.00749832f $X=7.9 $Y=0.18 $X2=0
+ $Y2=0
cc_1106 N_A_1493_21#_c_1538_n N_VGND_c_2320_n 3.25845e-19 $X=11.52 $Y=0.905
+ $X2=0 $Y2=0
cc_1107 N_A_1493_21#_c_1540_n N_VGND_c_2320_n 0.00870923f $X=9.135 $Y=0.75 $X2=0
+ $Y2=0
cc_1108 N_A_1493_21#_c_1541_n N_VGND_c_2320_n 0.0134555f $X=9.59 $Y=0.932 $X2=0
+ $Y2=0
cc_1109 N_A_1493_21#_c_1538_n A_2243_178# 0.00243848f $X=11.52 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_1110 N_A_1493_21#_c_1544_n A_2243_178# 6.94404e-19 $X=11.23 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_1111 N_A_1493_21#_c_1538_n A_2321_178# 0.00109775f $X=11.52 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_1112 N_A_1493_21#_c_1539_n A_2321_178# 0.0034525f $X=11.605 $Y=2 $X2=-0.19
+ $Y2=-0.245
cc_1113 N_SLEEP_B_M1010_g N_CLK_M1015_g 0.0180733f $X=10.25 $Y=2.415 $X2=0 $Y2=0
cc_1114 N_SLEEP_B_M1002_g N_CLK_M1013_g 0.0343257f $X=11.53 $Y=1.1 $X2=0 $Y2=0
cc_1115 N_SLEEP_B_c_1684_n N_CLK_M1013_g 0.00189667f $X=11.89 $Y=0.65 $X2=0
+ $Y2=0
cc_1116 N_SLEEP_B_c_1686_n N_CLK_M1013_g 6.95937e-19 $X=11.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1117 N_SLEEP_B_M1010_g CLK 0.0204751f $X=10.25 $Y=2.415 $X2=0 $Y2=0
cc_1118 N_SLEEP_B_M1010_g N_CLK_c_1750_n 0.0134213f $X=10.25 $Y=2.415 $X2=0
+ $Y2=0
cc_1119 N_SLEEP_B_c_1684_n N_A_2504_57#_c_1802_n 0.00698754f $X=11.89 $Y=0.65
+ $X2=0 $Y2=0
cc_1120 N_SLEEP_B_M1010_g N_VPWR_c_1861_n 5.65238e-19 $X=10.25 $Y=2.415 $X2=0
+ $Y2=0
cc_1121 N_SLEEP_B_M1010_g N_KAPWR_c_2176_n 0.00100017f $X=10.25 $Y=2.415 $X2=0
+ $Y2=0
cc_1122 N_SLEEP_B_M1010_g N_KAPWR_c_2164_n 0.00156815f $X=10.25 $Y=2.415 $X2=0
+ $Y2=0
cc_1123 N_SLEEP_B_c_1688_n N_VGND_c_2309_n 0.0190276f $X=11.89 $Y=0.485 $X2=0
+ $Y2=0
cc_1124 N_SLEEP_B_c_1689_n N_VGND_c_2309_n 0.0308482f $X=11.685 $Y=0.34 $X2=0
+ $Y2=0
cc_1125 N_SLEEP_B_c_1685_n N_VGND_c_2313_n 0.0120585f $X=10.175 $Y=0.415 $X2=0
+ $Y2=0
cc_1126 N_SLEEP_B_c_1687_n N_VGND_c_2313_n 0.109794f $X=10.135 $Y=0.415 $X2=0
+ $Y2=0
cc_1127 N_SLEEP_B_c_1688_n N_VGND_c_2313_n 0.00613609f $X=11.89 $Y=0.485 $X2=0
+ $Y2=0
cc_1128 N_SLEEP_B_c_1689_n N_VGND_c_2313_n 0.0225819f $X=11.685 $Y=0.34 $X2=0
+ $Y2=0
cc_1129 N_SLEEP_B_c_1685_n N_VGND_c_2320_n 0.0172795f $X=10.175 $Y=0.415 $X2=0
+ $Y2=0
cc_1130 N_SLEEP_B_c_1687_n N_VGND_c_2320_n 0.0643497f $X=10.135 $Y=0.415 $X2=0
+ $Y2=0
cc_1131 N_SLEEP_B_c_1688_n N_VGND_c_2320_n 0.00406047f $X=11.89 $Y=0.485 $X2=0
+ $Y2=0
cc_1132 N_SLEEP_B_c_1689_n N_VGND_c_2320_n 0.0125782f $X=11.685 $Y=0.34 $X2=0
+ $Y2=0
cc_1133 N_CLK_M1015_g N_VPWR_c_1861_n 5.65238e-19 $X=10.95 $Y=2.415 $X2=0 $Y2=0
cc_1134 N_CLK_M1015_g N_KAPWR_c_2214_n 9.84121e-19 $X=10.95 $Y=2.415 $X2=0 $Y2=0
cc_1135 N_CLK_M1015_g N_KAPWR_c_2164_n 0.00156815f $X=10.95 $Y=2.415 $X2=0 $Y2=0
cc_1136 N_A_2504_57#_M1024_g N_VPWR_c_1858_n 0.0071691f $X=13.425 $Y=2.465 $X2=0
+ $Y2=0
cc_1137 N_A_2504_57#_c_1804_n N_VPWR_c_1858_n 0.0431951f $X=12.665 $Y=1.98 $X2=0
+ $Y2=0
cc_1138 N_A_2504_57#_c_1800_n N_VPWR_c_1858_n 0.0214059f $X=13.33 $Y=1.48 $X2=0
+ $Y2=0
cc_1139 N_A_2504_57#_c_1801_n N_VPWR_c_1858_n 0.00300514f $X=13.33 $Y=1.48 $X2=0
+ $Y2=0
cc_1140 N_A_2504_57#_M1024_g N_VPWR_c_1862_n 0.0054895f $X=13.425 $Y=2.465 $X2=0
+ $Y2=0
cc_1141 N_A_2504_57#_M1024_g N_VPWR_c_1854_n 0.0072954f $X=13.425 $Y=2.465 $X2=0
+ $Y2=0
cc_1142 N_A_2504_57#_M1024_g N_KAPWR_c_2164_n 0.00753768f $X=13.425 $Y=2.465
+ $X2=0 $Y2=0
cc_1143 N_A_2504_57#_c_1804_n N_KAPWR_c_2164_n 0.0156751f $X=12.665 $Y=1.98
+ $X2=0 $Y2=0
cc_1144 N_A_2504_57#_M1024_g N_Q_c_2286_n 0.0137945f $X=13.425 $Y=2.465 $X2=0
+ $Y2=0
cc_1145 N_A_2504_57#_M1024_g N_Q_c_2287_n 0.00270474f $X=13.425 $Y=2.465 $X2=0
+ $Y2=0
cc_1146 N_A_2504_57#_c_1800_n N_Q_c_2287_n 0.00151667f $X=13.33 $Y=1.48 $X2=0
+ $Y2=0
cc_1147 N_A_2504_57#_M1031_g N_Q_c_2283_n 0.0157191f $X=13.425 $Y=0.705 $X2=0
+ $Y2=0
cc_1148 N_A_2504_57#_c_1800_n N_Q_c_2283_n 0.0262122f $X=13.33 $Y=1.48 $X2=0
+ $Y2=0
cc_1149 N_A_2504_57#_M1031_g Q 0.00270753f $X=13.425 $Y=0.705 $X2=0 $Y2=0
cc_1150 N_A_2504_57#_c_1800_n Q 0.00151667f $X=13.33 $Y=1.48 $X2=0 $Y2=0
cc_1151 N_A_2504_57#_M1031_g N_Q_c_2285_n 0.0112513f $X=13.425 $Y=0.705 $X2=0
+ $Y2=0
cc_1152 N_A_2504_57#_c_1799_n N_VGND_c_2309_n 0.0692985f $X=12.665 $Y=0.495
+ $X2=0 $Y2=0
cc_1153 N_A_2504_57#_c_1802_n N_VGND_c_2309_n 0.0010522f $X=12.665 $Y=1.48 $X2=0
+ $Y2=0
cc_1154 N_A_2504_57#_M1031_g N_VGND_c_2310_n 0.00381831f $X=13.425 $Y=0.705
+ $X2=0 $Y2=0
cc_1155 N_A_2504_57#_c_1799_n N_VGND_c_2310_n 0.0564479f $X=12.665 $Y=0.495
+ $X2=0 $Y2=0
cc_1156 N_A_2504_57#_c_1800_n N_VGND_c_2310_n 0.0214059f $X=13.33 $Y=1.48 $X2=0
+ $Y2=0
cc_1157 N_A_2504_57#_c_1801_n N_VGND_c_2310_n 0.00300514f $X=13.33 $Y=1.48 $X2=0
+ $Y2=0
cc_1158 N_A_2504_57#_c_1799_n N_VGND_c_2318_n 0.0220321f $X=12.665 $Y=0.495
+ $X2=0 $Y2=0
cc_1159 N_A_2504_57#_M1031_g N_VGND_c_2319_n 0.00502664f $X=13.425 $Y=0.705
+ $X2=0 $Y2=0
cc_1160 N_A_2504_57#_M1031_g N_VGND_c_2320_n 0.0102688f $X=13.425 $Y=0.705 $X2=0
+ $Y2=0
cc_1161 N_A_2504_57#_c_1799_n N_VGND_c_2320_n 0.0125808f $X=12.665 $Y=0.495
+ $X2=0 $Y2=0
cc_1162 N_VPWR_c_1855_n N_A_282_477#_c_2003_n 0.0133692f $X=0.73 $Y=2.53 $X2=0
+ $Y2=0
cc_1163 N_VPWR_c_1860_n N_A_282_477#_c_2003_n 0.0195955f $X=2.4 $Y=3.33 $X2=0
+ $Y2=0
cc_1164 N_VPWR_c_1854_n N_A_282_477#_c_2003_n 0.00309878f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1165 N_VPWR_M1039_d N_A_282_477#_c_2004_n 0.00395567f $X=2.31 $Y=2.385 $X2=0
+ $Y2=0
cc_1166 N_VPWR_c_1856_n N_A_282_477#_c_2004_n 0.0185325f $X=2.565 $Y=2.85 $X2=0
+ $Y2=0
cc_1167 N_VPWR_c_1855_n N_A_282_477#_c_2005_n 0.00419988f $X=0.73 $Y=2.53 $X2=0
+ $Y2=0
cc_1168 N_VPWR_M1039_d N_A_282_477#_c_2053_n 0.00581526f $X=2.31 $Y=2.385 $X2=0
+ $Y2=0
cc_1169 N_VPWR_c_1856_n N_A_282_477#_c_2053_n 0.0169891f $X=2.565 $Y=2.85 $X2=0
+ $Y2=0
cc_1170 N_VPWR_c_1857_n N_A_282_477#_c_2007_n 0.0943177f $X=5.495 $Y=3.33 $X2=0
+ $Y2=0
cc_1171 N_VPWR_c_1854_n N_A_282_477#_c_2007_n 0.0119304f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1172 N_VPWR_M1039_d N_A_282_477#_c_2008_n 9.80244e-19 $X=2.31 $Y=2.385 $X2=0
+ $Y2=0
cc_1173 N_VPWR_c_1856_n N_A_282_477#_c_2008_n 0.0138368f $X=2.565 $Y=2.85 $X2=0
+ $Y2=0
cc_1174 N_VPWR_c_1857_n N_A_282_477#_c_2008_n 0.0120507f $X=5.495 $Y=3.33 $X2=0
+ $Y2=0
cc_1175 N_VPWR_c_1854_n N_A_282_477#_c_2008_n 0.0015719f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1176 N_VPWR_M1039_d N_A_282_477#_c_2013_n 0.00407303f $X=2.31 $Y=2.385 $X2=0
+ $Y2=0
cc_1177 N_VPWR_c_1854_n N_A_282_477#_c_2013_n 2.59564e-19 $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1178 N_VPWR_c_1854_n A_1858_419# 0.00145452f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1179 N_VPWR_c_1854_n N_KAPWR_M1017_d 0.00131698f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1180 N_VPWR_c_1854_n N_KAPWR_M1015_d 0.00142981f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1181 N_VPWR_c_1861_n N_KAPWR_c_2176_n 0.0168759f $X=13.045 $Y=3.33 $X2=0
+ $Y2=0
cc_1182 N_VPWR_c_1854_n N_KAPWR_c_2176_n 0.00242436f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1183 N_VPWR_c_1861_n N_KAPWR_c_2214_n 0.0113274f $X=13.045 $Y=3.33 $X2=0
+ $Y2=0
cc_1184 N_VPWR_c_1854_n N_KAPWR_c_2214_n 0.00148498f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1185 N_VPWR_M1039_d N_KAPWR_c_2164_n 0.00388447f $X=2.31 $Y=2.385 $X2=0 $Y2=0
cc_1186 N_VPWR_M1036_d N_KAPWR_c_2164_n 0.00321696f $X=5.44 $Y=2.65 $X2=0 $Y2=0
cc_1187 N_VPWR_M1011_d N_KAPWR_c_2164_n 0.00244555f $X=12.955 $Y=1.835 $X2=0
+ $Y2=0
cc_1188 N_VPWR_c_1855_n N_KAPWR_c_2164_n 0.0290096f $X=0.73 $Y=2.53 $X2=0 $Y2=0
cc_1189 N_VPWR_c_1856_n N_KAPWR_c_2164_n 0.0245903f $X=2.565 $Y=2.85 $X2=0 $Y2=0
cc_1190 N_VPWR_c_1857_n N_KAPWR_c_2164_n 0.00467425f $X=5.495 $Y=3.33 $X2=0
+ $Y2=0
cc_1191 N_VPWR_c_1858_n N_KAPWR_c_2164_n 0.0341776f $X=13.21 $Y=1.98 $X2=0 $Y2=0
cc_1192 N_VPWR_c_1859_n N_KAPWR_c_2164_n 0.00122026f $X=0.565 $Y=3.33 $X2=0
+ $Y2=0
cc_1193 N_VPWR_c_1860_n N_KAPWR_c_2164_n 0.00637057f $X=2.4 $Y=3.33 $X2=0 $Y2=0
cc_1194 N_VPWR_c_1861_n N_KAPWR_c_2164_n 0.0145253f $X=13.045 $Y=3.33 $X2=0
+ $Y2=0
cc_1195 N_VPWR_c_1862_n N_KAPWR_c_2164_n 0.00124399f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1854_n N_KAPWR_c_2164_n 1.44221f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1197 N_VPWR_c_1866_n N_KAPWR_c_2164_n 0.00273721f $X=5.66 $Y=3.05 $X2=0 $Y2=0
cc_1198 N_VPWR_c_1854_n N_Q_M1024_d 0.00119401f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1199 N_VPWR_c_1862_n N_Q_c_2286_n 0.0231698f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1200 N_VPWR_c_1854_n N_Q_c_2286_n 0.00332052f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1201 N_VPWR_c_1858_n N_Q_c_2287_n 0.0494754f $X=13.21 $Y=1.98 $X2=0 $Y2=0
cc_1202 A_204_477# N_KAPWR_c_2164_n 0.00450483f $X=1.02 $Y=2.385 $X2=11.28
+ $Y2=2.82
cc_1203 N_A_282_477#_c_2004_n A_368_477# 0.00270984f $X=2.66 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_1204 N_A_282_477#_M1035_s N_KAPWR_c_2164_n 0.00199666f $X=4.115 $Y=2.65 $X2=0
+ $Y2=0
cc_1205 N_A_282_477#_c_2003_n N_KAPWR_c_2164_n 0.0317182f $X=1.55 $Y=2.53 $X2=0
+ $Y2=0
cc_1206 N_A_282_477#_c_2004_n N_KAPWR_c_2164_n 0.0406236f $X=2.66 $Y=2.405 $X2=0
+ $Y2=0
cc_1207 N_A_282_477#_c_2053_n N_KAPWR_c_2164_n 0.0150085f $X=2.905 $Y=2.905
+ $X2=0 $Y2=0
cc_1208 N_A_282_477#_c_2007_n N_KAPWR_c_2164_n 0.0329459f $X=4.095 $Y=2.99 $X2=0
+ $Y2=0
cc_1209 N_A_282_477#_c_2008_n N_KAPWR_c_2164_n 0.00250961f $X=2.99 $Y=2.99 $X2=0
+ $Y2=0
cc_1210 N_A_282_477#_c_2010_n N_KAPWR_c_2164_n 0.00485026f $X=4.095 $Y=2.15
+ $X2=0 $Y2=0
cc_1211 N_A_282_477#_c_2011_n N_KAPWR_c_2164_n 8.07963e-19 $X=3.805 $Y=2.15
+ $X2=0 $Y2=0
cc_1212 N_A_282_477#_c_2012_n N_KAPWR_c_2164_n 0.0275397f $X=4.26 $Y=2.85 $X2=0
+ $Y2=0
cc_1213 N_A_282_477#_c_2013_n N_KAPWR_c_2164_n 7.49401e-19 $X=2.905 $Y=2.405
+ $X2=0 $Y2=0
cc_1214 N_A_282_477#_c_2001_n N_VGND_c_2305_n 0.0119341f $X=1.69 $Y=0.46 $X2=0
+ $Y2=0
cc_1215 N_A_282_477#_c_1995_n N_VGND_c_2306_n 0.0129505f $X=2.135 $Y=0.585 $X2=0
+ $Y2=0
cc_1216 N_A_282_477#_c_1997_n N_VGND_c_2306_n 0.0144963f $X=2.485 $Y=0.925 $X2=0
+ $Y2=0
cc_1217 N_A_282_477#_c_2001_n N_VGND_c_2306_n 0.00650943f $X=1.69 $Y=0.46 $X2=0
+ $Y2=0
cc_1218 N_A_282_477#_c_1995_n N_VGND_c_2316_n 0.00968009f $X=2.135 $Y=0.585
+ $X2=0 $Y2=0
cc_1219 N_A_282_477#_c_2001_n N_VGND_c_2316_n 0.0203614f $X=1.69 $Y=0.46 $X2=0
+ $Y2=0
cc_1220 N_A_282_477#_M1003_d N_VGND_c_2320_n 0.00371678f $X=1.44 $Y=0.235 $X2=0
+ $Y2=0
cc_1221 N_A_282_477#_c_1995_n N_VGND_c_2320_n 0.0134428f $X=2.135 $Y=0.585 $X2=0
+ $Y2=0
cc_1222 N_A_282_477#_c_1997_n N_VGND_c_2320_n 0.00597146f $X=2.485 $Y=0.925
+ $X2=0 $Y2=0
cc_1223 N_A_282_477#_c_2001_n N_VGND_c_2320_n 0.0124836f $X=1.69 $Y=0.46 $X2=0
+ $Y2=0
cc_1224 N_A_282_477#_c_1995_n A_396_47# 0.0018379f $X=2.135 $Y=0.585 $X2=-0.19
+ $Y2=-0.245
cc_1225 A_368_477# N_KAPWR_c_2164_n 0.00430099f $X=1.84 $Y=2.385 $X2=2.66
+ $Y2=2.405
cc_1226 A_1010_530# N_KAPWR_c_2164_n 0.00117632f $X=5.05 $Y=2.65 $X2=4.11
+ $Y2=0.905
cc_1227 A_1372_379# N_KAPWR_c_2164_n 0.00850025f $X=6.86 $Y=1.895 $X2=11.28
+ $Y2=2.82
cc_1228 A_1858_419# N_KAPWR_c_2164_n 0.00318255f $X=9.29 $Y=2.095 $X2=3.78
+ $Y2=1.84
cc_1229 N_KAPWR_c_2164_n N_Q_c_2286_n 0.041515f $X=11.28 $Y=2.82 $X2=0 $Y2=0
cc_1230 N_Q_c_2285_n N_VGND_c_2310_n 0.0333828f $X=13.64 $Y=0.43 $X2=0 $Y2=0
cc_1231 N_Q_c_2285_n N_VGND_c_2319_n 0.0240548f $X=13.64 $Y=0.43 $X2=0 $Y2=0
cc_1232 N_Q_c_2285_n N_VGND_c_2320_n 0.0137416f $X=13.64 $Y=0.43 $X2=0 $Y2=0
cc_1233 N_VGND_c_2320_n A_210_47# 0.00352191f $X=13.68 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1234 N_VGND_c_2320_n A_396_47# 0.00235397f $X=13.68 $Y=0 $X2=-0.19 $Y2=-0.245
