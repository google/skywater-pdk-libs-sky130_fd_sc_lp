# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dfxbp_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.525000 1.315000 1.855000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.402600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.225000 0.905000 9.925000 1.075000 ;
        RECT 9.225000 1.075000 9.555000 2.890000 ;
        RECT 9.595000 0.615000 9.925000 0.905000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.515000 0.265000 12.845000 3.065000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.600000 0.440000 0.930000 1.285000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.110000  0.405000  0.420000 1.995000 ;
      RECT  0.110000  1.995000  0.440000 2.425000 ;
      RECT  0.110000  2.425000  1.320000 2.595000 ;
      RECT  0.110000  2.595000  0.440000 3.035000 ;
      RECT  0.640000  2.775000  0.970000 3.245000 ;
      RECT  1.110000  0.085000  1.360000 0.865000 ;
      RECT  1.150000  2.595000  1.320000 2.775000 ;
      RECT  1.150000  2.775000  2.315000 3.065000 ;
      RECT  1.170000  2.035000  3.110000 2.205000 ;
      RECT  1.170000  2.205000  1.500000 2.245000 ;
      RECT  1.720000  2.385000  2.050000 2.425000 ;
      RECT  1.720000  2.425000  3.665000 2.595000 ;
      RECT  1.820000  0.405000  2.150000 0.865000 ;
      RECT  1.820000  0.865000  1.990000 2.035000 ;
      RECT  2.250000  1.595000  2.660000 1.635000 ;
      RECT  2.250000  1.635000  4.215000 1.805000 ;
      RECT  2.250000  1.805000  2.580000 1.855000 ;
      RECT  2.330000  0.405000  2.660000 1.595000 ;
      RECT  2.780000  1.985000  3.110000 2.035000 ;
      RECT  2.780000  2.205000  3.110000 2.245000 ;
      RECT  3.075000  0.965000  4.780000 1.135000 ;
      RECT  3.075000  1.135000  3.405000 1.455000 ;
      RECT  3.280000  0.085000  3.610000 0.785000 ;
      RECT  3.335000  1.985000  3.665000 2.425000 ;
      RECT  3.335000  2.595000  3.665000 2.755000 ;
      RECT  3.865000  1.985000  4.195000 3.245000 ;
      RECT  4.045000  1.315000  4.430000 1.575000 ;
      RECT  4.045000  1.575000  4.215000 1.635000 ;
      RECT  4.150000  0.265000  5.480000 0.435000 ;
      RECT  4.150000  0.435000  4.480000 0.965000 ;
      RECT  4.395000  1.755000  4.780000 2.115000 ;
      RECT  4.395000  2.115000  6.470000 2.285000 ;
      RECT  4.395000  2.285000  4.780000 2.755000 ;
      RECT  4.610000  1.135000  4.780000 1.755000 ;
      RECT  4.710000  0.615000  5.130000 0.785000 ;
      RECT  4.960000  0.785000  5.130000 1.685000 ;
      RECT  4.960000  1.685000  7.265000 1.855000 ;
      RECT  4.960000  1.855000  5.290000 1.935000 ;
      RECT  5.310000  0.435000  5.480000 1.335000 ;
      RECT  5.310000  1.335000  6.740000 1.505000 ;
      RECT  5.490000  2.465000  5.820000 3.245000 ;
      RECT  5.660000  0.085000  5.910000 1.065000 ;
      RECT  6.140000  0.265000  8.155000 0.435000 ;
      RECT  6.140000  0.435000  6.390000 1.155000 ;
      RECT  6.140000  2.075000  6.470000 2.115000 ;
      RECT  6.140000  2.285000  6.470000 3.065000 ;
      RECT  6.570000  0.615000  7.600000 0.785000 ;
      RECT  6.570000  0.785000  6.740000 1.335000 ;
      RECT  6.670000  2.115000  7.615000 2.285000 ;
      RECT  6.670000  2.285000  7.000000 3.065000 ;
      RECT  6.920000  0.965000  7.090000 1.265000 ;
      RECT  6.920000  1.265000  8.695000 1.435000 ;
      RECT  6.935000  1.615000  7.265000 1.685000 ;
      RECT  6.935000  1.855000  7.265000 1.935000 ;
      RECT  7.270000  0.785000  7.600000 1.085000 ;
      RECT  7.445000  1.435000  7.615000 2.115000 ;
      RECT  7.795000  1.615000  8.125000 2.020000 ;
      RECT  7.795000  2.020000  9.045000 2.190000 ;
      RECT  7.795000  2.370000  8.125000 3.245000 ;
      RECT  7.825000  0.435000  8.155000 0.725000 ;
      RECT  8.335000  0.085000  8.585000 0.725000 ;
      RECT  8.365000  1.170000  8.695000 1.265000 ;
      RECT  8.365000  1.435000  8.695000 1.840000 ;
      RECT  8.590000  2.190000  9.045000 3.065000 ;
      RECT  8.875000  0.265000 10.275000 0.435000 ;
      RECT  8.875000  0.435000  9.375000 0.725000 ;
      RECT  8.875000  0.725000  9.045000 2.020000 ;
      RECT  9.735000  1.255000 11.765000 1.585000 ;
      RECT  9.755000  1.815000 10.085000 3.245000 ;
      RECT 10.105000  0.435000 10.275000 1.255000 ;
      RECT 10.285000  1.765000 12.335000 1.935000 ;
      RECT 10.285000  1.935000 10.615000 2.855000 ;
      RECT 10.465000  0.085000 10.715000 1.075000 ;
      RECT 11.175000  0.615000 11.505000 0.905000 ;
      RECT 11.175000  0.905000 12.175000 1.075000 ;
      RECT 11.725000  0.085000 12.055000 0.725000 ;
      RECT 11.985000  2.115000 12.315000 3.245000 ;
      RECT 12.005000  1.075000 12.175000 1.215000 ;
      RECT 12.005000  1.215000 12.335000 1.765000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
  END
END sky130_fd_sc_lp__dfxbp_lp
