* File: sky130_fd_sc_lp__maj3_1.pxi.spice
* Created: Fri Aug 28 10:42:53 2020
* 
x_PM_SKY130_FD_SC_LP__MAJ3_1%A N_A_M1002_g N_A_M1003_g N_A_M1013_g N_A_M1006_g A
+ A N_A_c_71_n PM_SKY130_FD_SC_LP__MAJ3_1%A
x_PM_SKY130_FD_SC_LP__MAJ3_1%B N_B_c_112_n N_B_M1000_g N_B_M1007_g N_B_c_107_n
+ N_B_M1001_g N_B_M1008_g N_B_c_115_n B B N_B_c_111_n
+ PM_SKY130_FD_SC_LP__MAJ3_1%B
x_PM_SKY130_FD_SC_LP__MAJ3_1%C N_C_M1004_g N_C_M1005_g N_C_c_156_n N_C_c_157_n
+ N_C_M1012_g N_C_M1009_g C C C N_C_c_160_n PM_SKY130_FD_SC_LP__MAJ3_1%C
x_PM_SKY130_FD_SC_LP__MAJ3_1%A_30_57# N_A_30_57#_M1004_s N_A_30_57#_M1007_d
+ N_A_30_57#_M1005_s N_A_30_57#_M1000_d N_A_30_57#_M1011_g N_A_30_57#_M1010_g
+ N_A_30_57#_c_207_n N_A_30_57#_c_217_n N_A_30_57#_c_208_n N_A_30_57#_c_218_n
+ N_A_30_57#_c_209_n N_A_30_57#_c_210_n N_A_30_57#_c_219_n N_A_30_57#_c_211_n
+ N_A_30_57#_c_221_n N_A_30_57#_c_212_n N_A_30_57#_c_213_n N_A_30_57#_c_214_n
+ N_A_30_57#_c_215_n PM_SKY130_FD_SC_LP__MAJ3_1%A_30_57#
x_PM_SKY130_FD_SC_LP__MAJ3_1%VPWR N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_c_297_n
+ N_VPWR_c_298_n VPWR N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n
+ N_VPWR_c_296_n N_VPWR_c_303_n N_VPWR_c_304_n PM_SKY130_FD_SC_LP__MAJ3_1%VPWR
x_PM_SKY130_FD_SC_LP__MAJ3_1%X N_X_M1011_d N_X_M1010_d X X X X X X X N_X_c_335_n
+ X PM_SKY130_FD_SC_LP__MAJ3_1%X
x_PM_SKY130_FD_SC_LP__MAJ3_1%VGND N_VGND_M1003_d N_VGND_M1012_d N_VGND_c_357_n
+ N_VGND_c_358_n N_VGND_c_359_n N_VGND_c_360_n VGND N_VGND_c_361_n
+ N_VGND_c_362_n N_VGND_c_363_n N_VGND_c_364_n PM_SKY130_FD_SC_LP__MAJ3_1%VGND
cc_1 VNB N_A_M1002_g 0.0098958f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.165
cc_2 VNB N_A_M1003_g 0.0337023f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.495
cc_3 VNB N_A_M1013_g 0.0115241f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.165
cc_4 VNB N_A_M1006_g 0.0315833f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=0.495
cc_5 VNB A 0.0140932f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_6 VNB N_A_c_71_n 0.0527773f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.29
cc_7 VNB N_B_M1007_g 0.0328822f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.495
cc_8 VNB N_B_c_107_n 0.0083577f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.455
cc_9 VNB N_B_M1001_g 0.031479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_M1008_g 0.00713519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB B 0.00758657f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.29
cc_12 VNB N_B_c_111_n 0.0366747f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.29
cc_13 VNB N_C_M1004_g 0.0686582f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.165
cc_14 VNB N_C_M1012_g 0.0551446f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.165
cc_15 VNB N_A_30_57#_M1011_g 0.0271637f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=0.495
cc_16 VNB N_A_30_57#_c_207_n 0.0217276f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.29
cc_17 VNB N_A_30_57#_c_208_n 0.00340376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_30_57#_c_209_n 0.0123431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_30_57#_c_210_n 0.0109271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_30_57#_c_211_n 0.0344089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_30_57#_c_212_n 0.0230986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_30_57#_c_213_n 0.00915735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_30_57#_c_214_n 0.00266963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_30_57#_c_215_n 0.0361206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_296_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB X 0.0101713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0261165f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.455
cc_28 VNB N_X_c_335_n 0.0303701f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.29
cc_29 VNB A_117_57# 0.00242931f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.455
cc_30 VNB N_VGND_c_357_n 0.00421131f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.455
cc_31 VNB N_VGND_c_358_n 0.0130575f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=1.125
cc_32 VNB N_VGND_c_359_n 0.0396119f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_33 VNB N_VGND_c_360_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_361_n 0.0301612f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.29
cc_35 VNB N_VGND_c_362_n 0.0199099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_363_n 0.230394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_364_n 0.00548753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_M1002_g 0.0326858f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=2.165
cc_39 VPB N_A_M1013_g 0.0246279f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.165
cc_40 VPB N_B_c_112_n 0.0310526f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.455
cc_41 VPB N_B_c_107_n 0.00226355f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=1.455
cc_42 VPB N_B_M1008_g 0.026099f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_B_c_115_n 0.0248112f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_C_M1004_g 0.0607767f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=2.165
cc_45 VPB N_C_c_156_n 0.125675f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=0.495
cc_46 VPB N_C_c_157_n 0.0146273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_C_M1012_g 0.0423658f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.165
cc_48 VPB C 0.02106f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_49 VPB N_C_c_160_n 0.0369217f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=1.29
cc_50 VPB N_A_30_57#_M1010_g 0.0265186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_30_57#_c_217_n 0.00326015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_30_57#_c_218_n 0.00243716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_30_57#_c_219_n 0.0349498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_30_57#_c_211_n 0.013647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_30_57#_c_221_n 0.00733693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_30_57#_c_215_n 0.00746577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_297_n 0.0171925f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=1.455
cc_58 VPB N_VPWR_c_298_n 0.0125909f $X=-0.19 $Y=1.655 $X2=1.5 $Y2=1.125
cc_59 VPB N_VPWR_c_299_n 0.0314195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_300_n 0.043554f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=1.29
cc_61 VPB N_VPWR_c_301_n 0.0161515f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.29
cc_62 VPB N_VPWR_c_296_n 0.0913406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_303_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_304_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB X 0.0551511f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=1.455
cc_66 N_A_M1002_g N_B_c_112_n 0.00196173f $X=0.87 $Y=2.165 $X2=-0.19 $Y2=-0.245
cc_67 N_A_M1006_g N_B_M1007_g 0.0303016f $X=1.5 $Y=0.495 $X2=0 $Y2=0
cc_68 A N_B_M1007_g 2.33261e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_M1013_g N_B_c_107_n 0.00586864f $X=1.3 $Y=2.165 $X2=0 $Y2=0
cc_70 N_A_M1013_g N_B_c_115_n 0.0498116f $X=1.3 $Y=2.165 $X2=0 $Y2=0
cc_71 A B 0.0220126f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_c_71_n B 0.00523388f $X=1.3 $Y=1.29 $X2=0 $Y2=0
cc_73 A N_B_c_111_n 2.16395e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_c_71_n N_B_c_111_n 0.0361703f $X=1.3 $Y=1.29 $X2=0 $Y2=0
cc_75 N_A_M1003_g N_C_M1004_g 0.0314383f $X=1.02 $Y=0.495 $X2=0 $Y2=0
cc_76 A N_C_M1004_g 0.0038312f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_71_n N_C_M1004_g 0.0821168f $X=1.3 $Y=1.29 $X2=0 $Y2=0
cc_78 N_A_M1002_g N_C_c_156_n 0.00917051f $X=0.87 $Y=2.165 $X2=0 $Y2=0
cc_79 N_A_M1013_g N_C_c_156_n 0.00536039f $X=1.3 $Y=2.165 $X2=0 $Y2=0
cc_80 N_A_M1002_g N_A_30_57#_c_219_n 0.00125204f $X=0.87 $Y=2.165 $X2=0 $Y2=0
cc_81 A N_A_30_57#_c_211_n 0.018391f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_M1003_g N_A_30_57#_c_212_n 0.0122644f $X=1.02 $Y=0.495 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_A_30_57#_c_212_n 0.0154714f $X=1.5 $Y=0.495 $X2=0 $Y2=0
cc_84 A N_A_30_57#_c_212_n 0.056283f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A_c_71_n N_A_30_57#_c_212_n 0.00460521f $X=1.3 $Y=1.29 $X2=0 $Y2=0
cc_86 N_A_M1006_g N_A_30_57#_c_213_n 0.00183449f $X=1.5 $Y=0.495 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_VPWR_c_297_n 0.0179957f $X=0.87 $Y=2.165 $X2=0 $Y2=0
cc_88 N_A_M1013_g N_VPWR_c_297_n 0.0132446f $X=1.3 $Y=2.165 $X2=0 $Y2=0
cc_89 A N_VPWR_c_297_n 0.0125214f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A_c_71_n N_VPWR_c_297_n 0.00218712f $X=1.3 $Y=1.29 $X2=0 $Y2=0
cc_91 N_A_M1003_g A_117_57# 0.00179116f $X=1.02 $Y=0.495 $X2=-0.19 $Y2=-0.245
cc_92 N_A_M1003_g N_VGND_c_357_n 0.00808391f $X=1.02 $Y=0.495 $X2=0 $Y2=0
cc_93 N_A_M1006_g N_VGND_c_357_n 0.00299959f $X=1.5 $Y=0.495 $X2=0 $Y2=0
cc_94 N_A_M1006_g N_VGND_c_359_n 0.0053602f $X=1.5 $Y=0.495 $X2=0 $Y2=0
cc_95 N_A_M1003_g N_VGND_c_361_n 0.00445056f $X=1.02 $Y=0.495 $X2=0 $Y2=0
cc_96 N_A_M1003_g N_VGND_c_363_n 0.00436882f $X=1.02 $Y=0.495 $X2=0 $Y2=0
cc_97 N_A_M1006_g N_VGND_c_363_n 0.00564987f $X=1.5 $Y=0.495 $X2=0 $Y2=0
cc_98 N_B_c_112_n N_C_c_156_n 0.00825049f $X=1.66 $Y=1.845 $X2=0 $Y2=0
cc_99 N_B_M1008_g N_C_c_156_n 0.00380464f $X=2.32 $Y=2.155 $X2=0 $Y2=0
cc_100 N_B_M1001_g N_C_M1012_g 0.145405f $X=2.32 $Y=0.495 $X2=0 $Y2=0
cc_101 B N_C_M1012_g 2.61234e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B_c_112_n C 0.00956853f $X=1.66 $Y=1.845 $X2=0 $Y2=0
cc_103 N_B_M1008_g C 0.00218263f $X=2.32 $Y=2.155 $X2=0 $Y2=0
cc_104 N_B_M1008_g N_A_30_57#_c_217_n 0.014988f $X=2.32 $Y=2.155 $X2=0 $Y2=0
cc_105 B N_A_30_57#_c_217_n 0.0045153f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B_M1001_g N_A_30_57#_c_208_n 0.00641404f $X=2.32 $Y=0.495 $X2=0 $Y2=0
cc_107 B N_A_30_57#_c_208_n 0.0110184f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_108 N_B_M1008_g N_A_30_57#_c_218_n 0.00610804f $X=2.32 $Y=2.155 $X2=0 $Y2=0
cc_109 N_B_c_112_n N_A_30_57#_c_221_n 0.00721757f $X=1.66 $Y=1.845 $X2=0 $Y2=0
cc_110 N_B_M1008_g N_A_30_57#_c_221_n 0.00900888f $X=2.32 $Y=2.155 $X2=0 $Y2=0
cc_111 N_B_c_115_n N_A_30_57#_c_221_n 0.00472421f $X=1.89 $Y=1.77 $X2=0 $Y2=0
cc_112 B N_A_30_57#_c_221_n 0.0137742f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B_c_111_n N_A_30_57#_c_221_n 0.00193648f $X=2.32 $Y=1.345 $X2=0 $Y2=0
cc_114 N_B_M1007_g N_A_30_57#_c_212_n 0.00840192f $X=1.89 $Y=0.495 $X2=0 $Y2=0
cc_115 B N_A_30_57#_c_212_n 0.0444499f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_116 N_B_M1007_g N_A_30_57#_c_213_n 0.0136704f $X=1.89 $Y=0.495 $X2=0 $Y2=0
cc_117 N_B_M1001_g N_A_30_57#_c_213_n 0.026982f $X=2.32 $Y=0.495 $X2=0 $Y2=0
cc_118 N_B_c_111_n N_A_30_57#_c_213_n 0.00224358f $X=2.32 $Y=1.345 $X2=0 $Y2=0
cc_119 B N_A_30_57#_c_214_n 0.0157531f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B_c_111_n N_A_30_57#_c_214_n 0.00599578f $X=2.32 $Y=1.345 $X2=0 $Y2=0
cc_121 N_B_c_112_n N_VPWR_c_297_n 0.00536519f $X=1.66 $Y=1.845 $X2=0 $Y2=0
cc_122 N_B_M1007_g N_VGND_c_359_n 0.00501304f $X=1.89 $Y=0.495 $X2=0 $Y2=0
cc_123 N_B_M1001_g N_VGND_c_359_n 0.00327726f $X=2.32 $Y=0.495 $X2=0 $Y2=0
cc_124 N_B_M1007_g N_VGND_c_363_n 0.00560802f $X=1.89 $Y=0.495 $X2=0 $Y2=0
cc_125 N_B_M1001_g N_VGND_c_363_n 0.00476272f $X=2.32 $Y=0.495 $X2=0 $Y2=0
cc_126 N_C_M1012_g N_A_30_57#_M1011_g 0.0213049f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_127 N_C_M1012_g N_A_30_57#_M1010_g 0.0155191f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_128 N_C_M1004_g N_A_30_57#_c_207_n 0.00382024f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_129 N_C_M1012_g N_A_30_57#_c_217_n 0.00447293f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_130 C N_A_30_57#_c_217_n 0.0130564f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_131 N_C_c_160_n N_A_30_57#_c_217_n 6.35942e-19 $X=2.59 $Y=2.9 $X2=0 $Y2=0
cc_132 N_C_M1012_g N_A_30_57#_c_208_n 0.00794704f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_133 N_C_M1012_g N_A_30_57#_c_218_n 0.00636649f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_134 N_C_M1012_g N_A_30_57#_c_209_n 0.0192428f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_135 N_C_M1004_g N_A_30_57#_c_219_n 0.0110828f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_136 N_C_M1004_g N_A_30_57#_c_211_n 0.0305642f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_137 N_C_c_156_n N_A_30_57#_c_221_n 0.00145861f $X=2.425 $Y=2.99 $X2=0 $Y2=0
cc_138 C N_A_30_57#_c_221_n 0.0209841f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_139 N_C_M1004_g N_A_30_57#_c_212_n 0.0178835f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_140 N_C_M1012_g N_A_30_57#_c_213_n 0.0140123f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_141 N_C_M1012_g N_A_30_57#_c_214_n 0.00248261f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_142 N_C_M1012_g N_A_30_57#_c_215_n 0.021376f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_143 N_C_M1004_g N_VPWR_c_297_n 0.0101104f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_144 N_C_c_156_n N_VPWR_c_297_n 0.0284974f $X=2.425 $Y=2.99 $X2=0 $Y2=0
cc_145 C N_VPWR_c_297_n 0.0218728f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_146 N_C_M1012_g N_VPWR_c_298_n 0.0181165f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_147 C N_VPWR_c_298_n 0.028797f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_148 N_C_c_157_n N_VPWR_c_299_n 0.0156578f $X=0.585 $Y=2.99 $X2=0 $Y2=0
cc_149 N_C_c_156_n N_VPWR_c_300_n 0.03313f $X=2.425 $Y=2.99 $X2=0 $Y2=0
cc_150 C N_VPWR_c_300_n 0.0728629f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_151 N_C_c_157_n N_VPWR_c_296_n 0.0596458f $X=0.585 $Y=2.99 $X2=0 $Y2=0
cc_152 C N_VPWR_c_296_n 0.0446602f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_153 N_C_M1004_g A_117_57# 0.00435548f $X=0.51 $Y=0.495 $X2=-0.19 $Y2=-0.245
cc_154 N_C_M1004_g N_VGND_c_357_n 8.06754e-19 $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_155 N_C_M1012_g N_VGND_c_358_n 0.0113398f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_156 N_C_M1012_g N_VGND_c_359_n 0.00508247f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_157 N_C_M1004_g N_VGND_c_361_n 0.00502664f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_158 N_C_M1004_g N_VGND_c_363_n 0.00647671f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_159 N_C_M1012_g N_VGND_c_363_n 0.00984795f $X=2.68 $Y=0.495 $X2=0 $Y2=0
cc_160 N_A_30_57#_c_219_n N_VPWR_c_297_n 0.0153904f $X=0.295 $Y=2.165 $X2=0
+ $Y2=0
cc_161 N_A_30_57#_c_221_n N_VPWR_c_297_n 0.0137622f $X=1.99 $Y=2.01 $X2=0 $Y2=0
cc_162 N_A_30_57#_M1010_g N_VPWR_c_298_n 0.0229076f $X=3.345 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_30_57#_c_217_n N_VPWR_c_298_n 0.00801352f $X=2.455 $Y=2.01 $X2=0
+ $Y2=0
cc_164 N_A_30_57#_c_218_n N_VPWR_c_298_n 0.00404551f $X=2.54 $Y=1.925 $X2=0
+ $Y2=0
cc_165 N_A_30_57#_c_209_n N_VPWR_c_298_n 0.0233889f $X=3.13 $Y=1.49 $X2=0 $Y2=0
cc_166 N_A_30_57#_c_215_n N_VPWR_c_298_n 0.00702351f $X=3.345 $Y=1.49 $X2=0
+ $Y2=0
cc_167 N_A_30_57#_M1010_g N_VPWR_c_301_n 0.00486043f $X=3.345 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_30_57#_M1010_g N_VPWR_c_296_n 0.00919827f $X=3.345 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_30_57#_c_217_n A_479_389# 0.00165069f $X=2.455 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A_30_57#_M1011_g X 0.00360697f $X=3.305 $Y=0.705 $X2=0 $Y2=0
cc_171 N_A_30_57#_c_215_n X 0.00191463f $X=3.345 $Y=1.49 $X2=0 $Y2=0
cc_172 N_A_30_57#_M1011_g X 0.00696188f $X=3.305 $Y=0.705 $X2=0 $Y2=0
cc_173 N_A_30_57#_c_209_n X 0.0258106f $X=3.13 $Y=1.49 $X2=0 $Y2=0
cc_174 N_A_30_57#_c_215_n X 0.0195681f $X=3.345 $Y=1.49 $X2=0 $Y2=0
cc_175 N_A_30_57#_M1011_g N_X_c_335_n 0.0112926f $X=3.305 $Y=0.705 $X2=0 $Y2=0
cc_176 N_A_30_57#_c_207_n A_117_57# 0.0125556f $X=0.295 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_177 N_A_30_57#_c_212_n A_117_57# 0.0212895f $X=1.94 $Y=0.605 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A_30_57#_c_212_n N_VGND_c_357_n 0.0211715f $X=1.94 $Y=0.605 $X2=0 $Y2=0
cc_179 N_A_30_57#_c_213_n N_VGND_c_357_n 0.00569139f $X=2.54 $Y=0.605 $X2=0
+ $Y2=0
cc_180 N_A_30_57#_M1011_g N_VGND_c_358_n 0.00865202f $X=3.305 $Y=0.705 $X2=0
+ $Y2=0
cc_181 N_A_30_57#_c_208_n N_VGND_c_358_n 0.0124602f $X=2.54 $Y=1.325 $X2=0 $Y2=0
cc_182 N_A_30_57#_c_209_n N_VGND_c_358_n 0.0269919f $X=3.13 $Y=1.49 $X2=0 $Y2=0
cc_183 N_A_30_57#_c_213_n N_VGND_c_358_n 0.0461867f $X=2.54 $Y=0.605 $X2=0 $Y2=0
cc_184 N_A_30_57#_c_215_n N_VGND_c_358_n 0.00484479f $X=3.345 $Y=1.49 $X2=0
+ $Y2=0
cc_185 N_A_30_57#_c_213_n N_VGND_c_359_n 0.0452281f $X=2.54 $Y=0.605 $X2=0 $Y2=0
cc_186 N_A_30_57#_c_207_n N_VGND_c_361_n 0.0167213f $X=0.295 $Y=0.495 $X2=0
+ $Y2=0
cc_187 N_A_30_57#_M1011_g N_VGND_c_362_n 0.00502664f $X=3.305 $Y=0.705 $X2=0
+ $Y2=0
cc_188 N_A_30_57#_M1011_g N_VGND_c_363_n 0.0103937f $X=3.305 $Y=0.705 $X2=0
+ $Y2=0
cc_189 N_A_30_57#_c_207_n N_VGND_c_363_n 0.0095959f $X=0.295 $Y=0.495 $X2=0
+ $Y2=0
cc_190 N_A_30_57#_c_212_n N_VGND_c_363_n 0.0309328f $X=1.94 $Y=0.605 $X2=0 $Y2=0
cc_191 N_A_30_57#_c_213_n N_VGND_c_363_n 0.025591f $X=2.54 $Y=0.605 $X2=0 $Y2=0
cc_192 N_VPWR_c_296_n N_X_M1010_d 0.0042346f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_301_n X 0.0163773f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_c_296_n X 0.00959046f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_195 N_X_c_335_n N_VGND_c_358_n 0.0335795f $X=3.52 $Y=0.43 $X2=0 $Y2=0
cc_196 N_X_c_335_n N_VGND_c_362_n 0.0247291f $X=3.52 $Y=0.43 $X2=0 $Y2=0
cc_197 N_X_c_335_n N_VGND_c_363_n 0.0141285f $X=3.52 $Y=0.43 $X2=0 $Y2=0
cc_198 A_117_57# N_VGND_c_357_n 0.0125869f $X=0.585 $Y=0.285 $X2=0 $Y2=0
cc_199 A_117_57# N_VGND_c_361_n 0.0208937f $X=0.585 $Y=0.285 $X2=0 $Y2=0
cc_200 A_117_57# N_VGND_c_363_n 0.0123466f $X=0.585 $Y=0.285 $X2=0 $Y2=0
