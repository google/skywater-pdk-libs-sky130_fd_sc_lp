* File: sky130_fd_sc_lp__dfbbn_1.spice
* Created: Wed Sep  2 09:42:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfbbn_1.pex.spice"
.subckt sky130_fd_sc_lp__dfbbn_1  VNB VPB CLK_N D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK_N	CLK_N
* VPB	VPB
* VNB	VNB
MM1029 N_A_113_67#_M1029_d N_CLK_N_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_113_67#_M1009_g N_A_223_119#_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.15645 AS=0.1155 PD=1.165 PS=1.39 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1022 N_A_460_449#_M1022_d N_D_M1022_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.15645 PD=0.7 PS=1.165 NRD=0 NRS=109.992 M=1 R=2.8 SA=75001.1
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1023 N_A_546_449#_M1023_d N_A_223_119#_M1023_g N_A_460_449#_M1022_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.110475 AS=0.0588 PD=0.96 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1038 A_702_110# N_A_113_67#_M1038_g N_A_546_449#_M1023_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.110475 PD=0.84 PS=0.96 NRD=44.28 NRS=38.568 M=1 R=2.8
+ SA=75002 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_A_755_398#_M1031_g A_702_110# VNB NSHORT L=0.15 W=0.42
+ AD=0.201283 AS=0.0882 PD=1.16887 PS=0.84 NRD=37.14 NRS=44.28 M=1 R=2.8
+ SA=75002.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1024 N_A_1013_66#_M1024_d N_SET_B_M1024_g N_VGND_M1031_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0912 AS=0.306717 PD=0.925 PS=1.78113 NRD=0 NRS=80.616 M=1
+ R=4.26667 SA=75002.5 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_755_398#_M1017_d N_A_546_449#_M1017_g N_A_1013_66#_M1024_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1803 AS=0.0912 PD=1.375 PS=0.925 NRD=42.504 NRS=0.936 M=1
+ R=4.26667 SA=75003 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1012 N_A_1013_66#_M1012_d N_A_1186_21#_M1012_g N_A_755_398#_M1017_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1803 PD=1.85 PS=1.375 NRD=0 NRS=42.504 M=1
+ R=4.26667 SA=75003.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 A_1442_119# N_A_755_398#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1152 AS=0.1824 PD=1 PS=1.85 NRD=23.436 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1025 N_A_1531_428#_M1025_d N_A_113_67#_M1025_g A_1442_119# VNB NSHORT L=0.15
+ W=0.64 AD=0.219955 AS=0.1152 PD=1.49132 PS=1 NRD=44.052 NRS=23.436 M=1
+ R=4.26667 SA=75000.7 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1018 A_1693_163# N_A_223_119#_M1018_g N_A_1531_428#_M1025_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.144345 PD=0.66 PS=0.978679 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.5 SB=75002 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_1741_137#_M1006_g A_1693_163# VNB NSHORT L=0.15 W=0.42
+ AD=0.110864 AS=0.0504 PD=0.883585 PS=0.66 NRD=34.284 NRS=18.564 M=1 R=2.8
+ SA=75001.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1026 N_A_1896_119#_M1026_d N_SET_B_M1026_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1088 AS=0.168936 PD=0.98 PS=1.34642 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75001.7 SB=75001 A=0.096 P=1.58 MULT=1
MM1001 N_A_1741_137#_M1001_d N_A_1531_428#_M1001_g N_A_1896_119#_M1026_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.122375 AS=0.1088 PD=1.175 PS=0.98 NRD=3.744
+ NRS=11.244 M=1 R=4.26667 SA=75002.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1014 N_A_1896_119#_M1014_d N_A_1186_21#_M1014_g N_A_1741_137#_M1001_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.2176 AS=0.122375 PD=1.96 PS=1.175 NRD=10.308
+ NRS=4.68 M=1 R=4.26667 SA=75001.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1002_d N_RESET_B_M1002_g N_A_1186_21#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1030 N_Q_N_M1030_d N_A_1741_137#_M1030_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1806 PD=2.25 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1034 N_VGND_M1034_d N_A_1741_137#_M1034_g N_A_2511_137#_M1034_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1035 N_Q_M1035_d N_A_2511_137#_M1035_g N_VGND_M1034_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1806 PD=2.25 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1027 N_A_113_67#_M1027_d N_CLK_N_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2336 AS=0.1824 PD=2.01 PS=1.85 NRD=24.6053 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1032 N_VPWR_M1032_d N_A_113_67#_M1032_g N_A_223_119#_M1032_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.17274 AS=0.1824 PD=1.36453 PS=1.85 NRD=24.6053 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75004.7 A=0.096 P=1.58 MULT=1
MM1008 N_A_460_449#_M1008_d N_D_M1008_g N_VPWR_M1032_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.11336 PD=0.7 PS=0.895472 NRD=0 NRS=62.1338 M=1 R=2.8 SA=75000.8
+ SB=75006.3 A=0.063 P=1.14 MULT=1
MM1036 N_A_546_449#_M1036_d N_A_113_67#_M1036_g N_A_460_449#_M1008_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.13755 AS=0.0588 PD=1.075 PS=0.7 NRD=175.882 NRS=0 M=1 R=2.8
+ SA=75001.3 SB=75005.9 A=0.063 P=1.14 MULT=1
MM1033 A_707_449# N_A_223_119#_M1033_g N_A_546_449#_M1036_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.13755 PD=0.66 PS=1.075 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75005.1 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_755_398#_M1010_g A_707_449# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.222917 AS=0.0504 PD=1.42667 PS=0.66 NRD=223.142 NRS=30.4759 M=1 R=2.8
+ SA=75002.5 SB=75004.7 A=0.063 P=1.14 MULT=1
MM1037 N_A_755_398#_M1037_d N_SET_B_M1037_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.357 AS=0.445833 PD=1.69 PS=2.85333 NRD=133.665 NRS=111.561 M=1
+ R=5.6 SA=75002 SB=75003.2 A=0.126 P=1.98 MULT=1
MM1003 A_1228_379# N_A_546_449#_M1003_g N_A_755_398#_M1037_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1008 AS=0.357 PD=1.08 PS=1.69 NRD=15.2281 NRS=0 M=1 R=5.6 SA=75003
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1020 N_VPWR_M1020_d N_A_1186_21#_M1020_g A_1228_379# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.21 AS=0.1008 PD=1.34 PS=1.08 NRD=51.5943 NRS=15.2281 M=1 R=5.6 SA=75003.4
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1004 A_1436_379# N_A_755_398#_M1004_g N_VPWR_M1020_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.157937 AS=0.21 PD=1.41 PS=1.34 NRD=31.1851 NRS=0 M=1 R=5.6 SA=75004
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1021 N_A_1531_428#_M1021_d N_A_223_119#_M1021_g A_1436_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2254 AS=0.157937 PD=1.70667 PS=1.41 NRD=18.7544 NRS=31.1851 M=1
+ R=5.6 SA=75003.7 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1039 A_1649_512# N_A_113_67#_M1039_g N_A_1531_428#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.13545 AS=0.1127 PD=1.065 PS=0.853333 NRD=125.469 NRS=100.056 M=1
+ R=2.8 SA=75002.7 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_1741_137#_M1000_g A_1649_512# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.117808 AS=0.13545 PD=0.933333 PS=1.065 NRD=93.7917 NRS=125.469 M=1
+ R=2.8 SA=75003.5 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1015 N_A_1741_137#_M1015_d N_SET_B_M1015_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1176 AS=0.235617 PD=1.12 PS=1.86667 NRD=0 NRS=18.7544 M=1 R=5.6
+ SA=75002.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1028 A_2036_451# N_A_1531_428#_M1028_g N_A_1741_137#_M1015_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.0882 AS=0.1176 PD=1.05 PS=1.12 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75002.6 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_A_1186_21#_M1013_g A_2036_451# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2352 AS=0.0882 PD=2.24 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75003
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_RESET_B_M1007_g N_A_1186_21#_M1007_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.135006 AS=0.176 PD=1.088 PS=1.83 NRD=47.9892 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1011 N_Q_N_M1011_d N_A_1741_137#_M1011_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3465 AS=0.265794 PD=3.07 PS=2.142 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1019_d N_A_1741_137#_M1019_g N_A_2511_137#_M1019_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.137128 AS=0.176 PD=1.09137 PS=1.83 NRD=25.3933 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1016 N_Q_M1016_d N_A_2511_137#_M1016_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.269972 PD=3.09 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=26.8573 P=32.57
c_148 VNB 0 2.36507e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dfbbn_1.pxi.spice"
*
.ends
*
*
