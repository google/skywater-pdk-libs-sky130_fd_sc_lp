* File: sky130_fd_sc_lp__o31a_lp.pxi.spice
* Created: Wed Sep  2 10:24:51 2020
* 
x_PM_SKY130_FD_SC_LP__O31A_LP%B1 N_B1_M1010_g N_B1_M1009_g N_B1_c_78_n
+ N_B1_c_79_n B1 B1 N_B1_c_80_n N_B1_c_81_n PM_SKY130_FD_SC_LP__O31A_LP%B1
x_PM_SKY130_FD_SC_LP__O31A_LP%A3 N_A3_M1004_g N_A3_M1006_g N_A3_c_116_n
+ N_A3_c_117_n A3 A3 N_A3_c_119_n PM_SKY130_FD_SC_LP__O31A_LP%A3
x_PM_SKY130_FD_SC_LP__O31A_LP%A2 N_A2_M1002_g N_A2_M1005_g N_A2_c_163_n
+ N_A2_c_168_n A2 A2 N_A2_c_165_n PM_SKY130_FD_SC_LP__O31A_LP%A2
x_PM_SKY130_FD_SC_LP__O31A_LP%A1 N_A1_M1008_g N_A1_M1007_g N_A1_c_206_n
+ N_A1_c_207_n N_A1_c_208_n N_A1_c_209_n N_A1_c_214_n A1 A1 N_A1_c_211_n
+ PM_SKY130_FD_SC_LP__O31A_LP%A1
x_PM_SKY130_FD_SC_LP__O31A_LP%A_37_57# N_A_37_57#_M1009_s N_A_37_57#_M1010_d
+ N_A_37_57#_c_255_n N_A_37_57#_M1000_g N_A_37_57#_M1003_g N_A_37_57#_M1001_g
+ N_A_37_57#_c_257_n N_A_37_57#_c_258_n N_A_37_57#_c_259_n N_A_37_57#_c_267_n
+ N_A_37_57#_c_268_n N_A_37_57#_c_269_n N_A_37_57#_c_270_n N_A_37_57#_c_260_n
+ N_A_37_57#_c_261_n N_A_37_57#_c_262_n N_A_37_57#_c_263_n N_A_37_57#_c_272_n
+ N_A_37_57#_c_264_n PM_SKY130_FD_SC_LP__O31A_LP%A_37_57#
x_PM_SKY130_FD_SC_LP__O31A_LP%VPWR N_VPWR_M1010_s N_VPWR_M1007_d N_VPWR_c_349_n
+ N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n VPWR
+ N_VPWR_c_354_n N_VPWR_c_348_n PM_SKY130_FD_SC_LP__O31A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O31A_LP%X N_X_M1001_d N_X_M1003_d N_X_c_385_n X X X
+ N_X_c_386_n X PM_SKY130_FD_SC_LP__O31A_LP%X
x_PM_SKY130_FD_SC_LP__O31A_LP%A_140_57# N_A_140_57#_M1009_d N_A_140_57#_M1005_d
+ N_A_140_57#_c_404_n N_A_140_57#_c_405_n N_A_140_57#_c_406_n
+ N_A_140_57#_c_407_n PM_SKY130_FD_SC_LP__O31A_LP%A_140_57#
x_PM_SKY130_FD_SC_LP__O31A_LP%VGND N_VGND_M1004_d N_VGND_M1008_d N_VGND_c_439_n
+ N_VGND_c_440_n N_VGND_c_441_n VGND N_VGND_c_442_n N_VGND_c_443_n
+ N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_446_n PM_SKY130_FD_SC_LP__O31A_LP%VGND
cc_1 VNB N_B1_M1009_g 0.0374413f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.495
cc_2 VNB N_B1_c_78_n 0.0234927f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.63
cc_3 VNB N_B1_c_79_n 0.00173762f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.795
cc_4 VNB N_B1_c_80_n 0.0165772f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.29
cc_5 VNB N_B1_c_81_n 0.00724108f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.29
cc_6 VNB N_A3_M1004_g 0.0349725f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.55
cc_7 VNB N_A3_c_116_n 0.0208807f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.63
cc_8 VNB N_A3_c_117_n 0.00154443f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.795
cc_9 VNB A3 0.00534248f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_A3_c_119_n 0.01542f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.29
cc_11 VNB N_A2_M1005_g 0.0367745f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.495
cc_12 VNB N_A2_c_163_n 0.0217596f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.63
cc_13 VNB A2 0.00184734f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_14 VNB N_A2_c_165_n 0.0163353f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.29
cc_15 VNB N_A1_c_206_n 0.0145128f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.125
cc_16 VNB N_A1_c_207_n 0.0131584f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.63
cc_17 VNB N_A1_c_208_n 0.0143108f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_18 VNB N_A1_c_209_n 0.019754f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_19 VNB A1 0.00579675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_211_n 0.0153029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_37_57#_c_255_n 0.0319623f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.495
cc_22 VNB N_A_37_57#_M1003_g 0.00335186f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.795
cc_23 VNB N_A_37_57#_c_257_n 0.0243688f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.29
cc_24 VNB N_A_37_57#_c_258_n 0.0147236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_37_57#_c_259_n 0.0452662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_37_57#_c_260_n 0.00455898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_37_57#_c_261_n 0.0367122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_37_57#_c_262_n 3.35121e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_37_57#_c_263_n 0.0308105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_37_57#_c_264_n 0.00307274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_348_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_385_n 0.0268447f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.125
cc_33 VNB N_X_c_386_n 0.0438671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_140_57#_c_404_n 0.00312002f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.29
cc_35 VNB N_A_140_57#_c_405_n 0.0197287f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.63
cc_36 VNB N_A_140_57#_c_406_n 0.008113f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.795
cc_37 VNB N_A_140_57#_c_407_n 0.00249624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_439_n 0.00645068f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.29
cc_39 VNB N_VGND_c_440_n 0.0163422f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.63
cc_40 VNB N_VGND_c_441_n 0.00548867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_442_n 0.0330936f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.29
cc_42 VNB N_VGND_c_443_n 0.0269679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_444_n 0.209831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_445_n 0.00632158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_446_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_B1_M1010_g 0.0350283f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.55
cc_47 VPB N_B1_c_79_n 0.0119856f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.795
cc_48 VPB N_B1_c_81_n 0.00194981f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.29
cc_49 VPB N_A3_M1006_g 0.0315535f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.495
cc_50 VPB N_A3_c_117_n 0.0109177f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.795
cc_51 VPB A3 0.00164914f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_52 VPB N_A2_M1002_g 0.0291847f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.55
cc_53 VPB N_A2_c_163_n 0.00129603f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.63
cc_54 VPB N_A2_c_168_n 0.0135443f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.795
cc_55 VPB A2 7.46703e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_56 VPB N_A1_M1007_g 0.0288441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A1_c_209_n 0.00118947f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_58 VPB N_A1_c_214_n 0.0125844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB A1 0.00207774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_37_57#_M1003_g 0.0439947f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.795
cc_61 VPB N_A_37_57#_c_259_n 0.0156122f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_37_57#_c_267_n 0.00670675f $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.665
cc_63 VPB N_A_37_57#_c_268_n 0.0122924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_37_57#_c_269_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_37_57#_c_270_n 0.0215294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_37_57#_c_262_n 0.00295236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_37_57#_c_272_n 0.00796264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_349_n 0.0138708f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.495
cc_69 VPB N_VPWR_c_350_n 0.0327755f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.29
cc_70 VPB N_VPWR_c_351_n 0.00164766f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_71 VPB N_VPWR_c_352_n 0.0523707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_353_n 0.00491794f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.29
cc_73 VPB N_VPWR_c_354_n 0.0209811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_348_n 0.0769451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB X 0.0590168f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_76 VPB N_X_c_386_n 0.0127377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 N_B1_M1009_g N_A3_M1004_g 0.0240663f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_78 N_B1_M1010_g N_A3_M1006_g 0.0197584f $X=0.625 $Y=2.55 $X2=0 $Y2=0
cc_79 N_B1_c_78_n N_A3_c_116_n 0.0139302f $X=0.605 $Y=1.63 $X2=0 $Y2=0
cc_80 N_B1_c_79_n N_A3_c_117_n 0.0139302f $X=0.605 $Y=1.795 $X2=0 $Y2=0
cc_81 N_B1_c_80_n A3 7.74725e-19 $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_82 N_B1_c_81_n A3 0.0511345f $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_83 N_B1_c_80_n N_A3_c_119_n 0.0139302f $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_84 N_B1_c_81_n N_A3_c_119_n 0.00386561f $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_85 N_B1_M1010_g N_A_37_57#_c_259_n 0.00603123f $X=0.625 $Y=2.55 $X2=0 $Y2=0
cc_86 N_B1_M1009_g N_A_37_57#_c_259_n 0.00952738f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_87 N_B1_c_80_n N_A_37_57#_c_259_n 0.0148853f $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_88 N_B1_c_81_n N_A_37_57#_c_259_n 0.0485328f $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_89 N_B1_M1010_g N_A_37_57#_c_267_n 0.0195058f $X=0.625 $Y=2.55 $X2=0 $Y2=0
cc_90 N_B1_c_79_n N_A_37_57#_c_267_n 4.05894e-19 $X=0.605 $Y=1.795 $X2=0 $Y2=0
cc_91 N_B1_c_81_n N_A_37_57#_c_267_n 0.0208232f $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_92 N_B1_M1010_g N_A_37_57#_c_269_n 0.0192808f $X=0.625 $Y=2.55 $X2=0 $Y2=0
cc_93 N_B1_M1009_g N_A_37_57#_c_263_n 0.00891111f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_94 N_B1_c_80_n N_A_37_57#_c_263_n 3.54928e-19 $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_95 N_B1_c_81_n N_A_37_57#_c_263_n 0.00244611f $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_96 N_B1_M1010_g N_A_37_57#_c_272_n 0.00381008f $X=0.625 $Y=2.55 $X2=0 $Y2=0
cc_97 N_B1_c_81_n N_A_37_57#_c_272_n 0.00677849f $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_98 N_B1_M1010_g N_VPWR_c_350_n 0.0188987f $X=0.625 $Y=2.55 $X2=0 $Y2=0
cc_99 N_B1_M1010_g N_VPWR_c_352_n 0.0077588f $X=0.625 $Y=2.55 $X2=0 $Y2=0
cc_100 N_B1_M1010_g N_VPWR_c_348_n 0.0134709f $X=0.625 $Y=2.55 $X2=0 $Y2=0
cc_101 N_B1_M1009_g N_A_140_57#_c_404_n 0.0073428f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_102 N_B1_M1009_g N_A_140_57#_c_406_n 0.00540509f $X=0.625 $Y=0.495 $X2=0
+ $Y2=0
cc_103 N_B1_c_80_n N_A_140_57#_c_406_n 5.40842e-19 $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_104 N_B1_c_81_n N_A_140_57#_c_406_n 0.0110421f $X=0.605 $Y=1.29 $X2=0 $Y2=0
cc_105 N_B1_M1009_g N_VGND_c_442_n 0.00502664f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_106 N_B1_M1009_g N_VGND_c_444_n 0.0103301f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_107 N_A3_M1006_g N_A2_M1002_g 0.0698785f $X=1.155 $Y=2.55 $X2=0 $Y2=0
cc_108 N_A3_M1004_g N_A2_M1005_g 0.0220632f $X=1.085 $Y=0.495 $X2=0 $Y2=0
cc_109 A3 N_A2_M1005_g 9.46497e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A3_c_119_n N_A2_M1005_g 0.00203482f $X=1.145 $Y=1.29 $X2=0 $Y2=0
cc_111 N_A3_c_116_n N_A2_c_163_n 0.0130541f $X=1.145 $Y=1.63 $X2=0 $Y2=0
cc_112 N_A3_M1006_g N_A2_c_168_n 0.00257269f $X=1.155 $Y=2.55 $X2=0 $Y2=0
cc_113 N_A3_c_117_n N_A2_c_168_n 0.0130541f $X=1.145 $Y=1.795 $X2=0 $Y2=0
cc_114 N_A3_M1006_g A2 3.02847e-19 $X=1.155 $Y=2.55 $X2=0 $Y2=0
cc_115 A3 A2 0.0429319f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A3_c_119_n A2 7.8e-19 $X=1.145 $Y=1.29 $X2=0 $Y2=0
cc_117 A3 N_A2_c_165_n 0.0035618f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_118 N_A3_c_119_n N_A2_c_165_n 0.0130541f $X=1.145 $Y=1.29 $X2=0 $Y2=0
cc_119 N_A3_M1006_g N_A_37_57#_c_269_n 0.0179394f $X=1.155 $Y=2.55 $X2=0 $Y2=0
cc_120 N_A3_M1006_g N_A_37_57#_c_270_n 0.0189134f $X=1.155 $Y=2.55 $X2=0 $Y2=0
cc_121 A3 N_A_37_57#_c_270_n 0.0158531f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A3_M1006_g N_A_37_57#_c_272_n 0.00261321f $X=1.155 $Y=2.55 $X2=0 $Y2=0
cc_123 N_A3_c_117_n N_A_37_57#_c_272_n 6.26696e-19 $X=1.145 $Y=1.795 $X2=0 $Y2=0
cc_124 A3 N_A_37_57#_c_272_n 0.00577003f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A3_M1006_g N_VPWR_c_350_n 8.9247e-19 $X=1.155 $Y=2.55 $X2=0 $Y2=0
cc_126 N_A3_M1006_g N_VPWR_c_352_n 0.00867649f $X=1.155 $Y=2.55 $X2=0 $Y2=0
cc_127 N_A3_M1006_g N_VPWR_c_348_n 0.015834f $X=1.155 $Y=2.55 $X2=0 $Y2=0
cc_128 N_A3_M1004_g N_A_140_57#_c_404_n 0.00233034f $X=1.085 $Y=0.495 $X2=0
+ $Y2=0
cc_129 N_A3_M1004_g N_A_140_57#_c_405_n 0.0125094f $X=1.085 $Y=0.495 $X2=0 $Y2=0
cc_130 A3 N_A_140_57#_c_405_n 0.0230313f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_131 N_A3_c_119_n N_A_140_57#_c_405_n 0.00106308f $X=1.145 $Y=1.29 $X2=0 $Y2=0
cc_132 A3 N_A_140_57#_c_406_n 0.00162016f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_133 N_A3_c_119_n N_A_140_57#_c_406_n 4.2995e-19 $X=1.145 $Y=1.29 $X2=0 $Y2=0
cc_134 N_A3_M1004_g N_A_140_57#_c_407_n 8.24409e-19 $X=1.085 $Y=0.495 $X2=0
+ $Y2=0
cc_135 N_A3_M1004_g N_VGND_c_439_n 0.00300153f $X=1.085 $Y=0.495 $X2=0 $Y2=0
cc_136 N_A3_M1004_g N_VGND_c_442_n 0.0053602f $X=1.085 $Y=0.495 $X2=0 $Y2=0
cc_137 N_A3_M1004_g N_VGND_c_444_n 0.00589472f $X=1.085 $Y=0.495 $X2=0 $Y2=0
cc_138 N_A2_M1002_g N_A1_M1007_g 0.0658237f $X=1.675 $Y=2.55 $X2=0 $Y2=0
cc_139 N_A2_M1005_g N_A1_c_206_n 0.01647f $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_140 N_A2_M1005_g N_A1_c_208_n 0.00999702f $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_141 N_A2_c_163_n N_A1_c_209_n 0.0139741f $X=1.685 $Y=1.675 $X2=0 $Y2=0
cc_142 N_A2_c_168_n N_A1_c_214_n 0.0139741f $X=1.685 $Y=1.84 $X2=0 $Y2=0
cc_143 A2 A1 0.0479466f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A2_c_165_n A1 0.00382624f $X=1.685 $Y=1.335 $X2=0 $Y2=0
cc_145 A2 N_A1_c_211_n 8.17732e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A2_c_165_n N_A1_c_211_n 0.0139741f $X=1.685 $Y=1.335 $X2=0 $Y2=0
cc_147 N_A2_M1002_g N_A_37_57#_c_269_n 0.00376793f $X=1.675 $Y=2.55 $X2=0 $Y2=0
cc_148 N_A2_M1002_g N_A_37_57#_c_270_n 0.0224765f $X=1.675 $Y=2.55 $X2=0 $Y2=0
cc_149 N_A2_c_168_n N_A_37_57#_c_270_n 5.36606e-19 $X=1.685 $Y=1.84 $X2=0 $Y2=0
cc_150 A2 N_A_37_57#_c_270_n 0.0241241f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_151 N_A2_M1002_g N_VPWR_c_351_n 0.00367597f $X=1.675 $Y=2.55 $X2=0 $Y2=0
cc_152 N_A2_M1002_g N_VPWR_c_352_n 0.00901271f $X=1.675 $Y=2.55 $X2=0 $Y2=0
cc_153 N_A2_M1002_g N_VPWR_c_348_n 0.0167409f $X=1.675 $Y=2.55 $X2=0 $Y2=0
cc_154 N_A2_M1005_g N_A_140_57#_c_405_n 0.0116186f $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_155 A2 N_A_140_57#_c_405_n 0.0217131f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A2_c_165_n N_A_140_57#_c_405_n 0.00129241f $X=1.685 $Y=1.335 $X2=0
+ $Y2=0
cc_157 N_A2_M1005_g N_A_140_57#_c_407_n 0.00826863f $X=1.645 $Y=0.495 $X2=0
+ $Y2=0
cc_158 N_A2_M1005_g N_VGND_c_439_n 0.00343383f $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_159 N_A2_M1005_g N_VGND_c_440_n 0.00502664f $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_160 N_A2_M1005_g N_VGND_c_441_n 5.43415e-19 $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_161 N_A2_M1005_g N_VGND_c_444_n 0.00576058f $X=1.645 $Y=0.495 $X2=0 $Y2=0
cc_162 N_A1_c_206_n N_A_37_57#_c_255_n 0.0106065f $X=2.105 $Y=0.78 $X2=0 $Y2=0
cc_163 N_A1_M1007_g N_A_37_57#_M1003_g 0.028901f $X=2.215 $Y=2.55 $X2=0 $Y2=0
cc_164 N_A1_c_209_n N_A_37_57#_M1003_g 0.0133154f $X=2.225 $Y=1.675 $X2=0 $Y2=0
cc_165 A1 N_A_37_57#_M1003_g 2.78512e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_166 N_A1_c_207_n N_A_37_57#_c_257_n 0.0100718f $X=2.105 $Y=0.93 $X2=0 $Y2=0
cc_167 N_A1_c_209_n N_A_37_57#_c_258_n 0.0134404f $X=2.225 $Y=1.675 $X2=0 $Y2=0
cc_168 N_A1_M1007_g N_A_37_57#_c_270_n 0.0218129f $X=2.215 $Y=2.55 $X2=0 $Y2=0
cc_169 N_A1_c_214_n N_A_37_57#_c_270_n 5.43235e-19 $X=2.225 $Y=1.84 $X2=0 $Y2=0
cc_170 A1 N_A_37_57#_c_270_n 0.0253346f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A1_c_208_n N_A_37_57#_c_260_n 0.00455969f $X=2.225 $Y=1.17 $X2=0 $Y2=0
cc_172 A1 N_A_37_57#_c_260_n 0.0489912f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A1_c_211_n N_A_37_57#_c_260_n 0.00125722f $X=2.225 $Y=1.335 $X2=0 $Y2=0
cc_174 N_A1_c_208_n N_A_37_57#_c_261_n 0.00643306f $X=2.225 $Y=1.17 $X2=0 $Y2=0
cc_175 A1 N_A_37_57#_c_261_n 5.17119e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_176 N_A1_c_211_n N_A_37_57#_c_261_n 0.0134404f $X=2.225 $Y=1.335 $X2=0 $Y2=0
cc_177 N_A1_M1007_g N_A_37_57#_c_262_n 0.00348712f $X=2.215 $Y=2.55 $X2=0 $Y2=0
cc_178 N_A1_c_214_n N_A_37_57#_c_262_n 0.00125722f $X=2.225 $Y=1.84 $X2=0 $Y2=0
cc_179 N_A1_c_209_n N_A_37_57#_c_264_n 0.00125722f $X=2.225 $Y=1.675 $X2=0 $Y2=0
cc_180 N_A1_M1007_g N_VPWR_c_351_n 0.0191131f $X=2.215 $Y=2.55 $X2=0 $Y2=0
cc_181 N_A1_M1007_g N_VPWR_c_352_n 0.00809503f $X=2.215 $Y=2.55 $X2=0 $Y2=0
cc_182 N_A1_M1007_g N_VPWR_c_348_n 0.0143777f $X=2.215 $Y=2.55 $X2=0 $Y2=0
cc_183 N_A1_c_206_n N_A_140_57#_c_405_n 0.004951f $X=2.105 $Y=0.78 $X2=0 $Y2=0
cc_184 N_A1_c_208_n N_A_140_57#_c_405_n 2.19279e-19 $X=2.225 $Y=1.17 $X2=0 $Y2=0
cc_185 N_A1_c_206_n N_A_140_57#_c_407_n 0.00167928f $X=2.105 $Y=0.78 $X2=0 $Y2=0
cc_186 N_A1_c_206_n N_VGND_c_440_n 0.00445056f $X=2.105 $Y=0.78 $X2=0 $Y2=0
cc_187 N_A1_c_206_n N_VGND_c_441_n 0.00957284f $X=2.105 $Y=0.78 $X2=0 $Y2=0
cc_188 N_A1_c_207_n N_VGND_c_441_n 0.00218225f $X=2.105 $Y=0.93 $X2=0 $Y2=0
cc_189 A1 N_VGND_c_441_n 0.0112443f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A1_c_211_n N_VGND_c_441_n 0.00122446f $X=2.225 $Y=1.335 $X2=0 $Y2=0
cc_191 N_A1_c_206_n N_VGND_c_444_n 0.0081158f $X=2.105 $Y=0.78 $X2=0 $Y2=0
cc_192 N_A_37_57#_c_267_n N_VPWR_M1010_s 0.00228864f $X=0.725 $Y=2.06 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_37_57#_c_268_n N_VPWR_M1010_s 7.4681e-19 $X=0.26 $Y=2.06 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_37_57#_c_270_n N_VPWR_M1007_d 0.00180746f $X=2.575 $Y=2.105 $X2=0
+ $Y2=0
cc_195 N_A_37_57#_c_267_n N_VPWR_c_350_n 0.0159361f $X=0.725 $Y=2.06 $X2=0 $Y2=0
cc_196 N_A_37_57#_c_268_n N_VPWR_c_350_n 0.00559555f $X=0.26 $Y=2.06 $X2=0 $Y2=0
cc_197 N_A_37_57#_c_269_n N_VPWR_c_350_n 0.0487591f $X=0.89 $Y=2.195 $X2=0 $Y2=0
cc_198 N_A_37_57#_M1003_g N_VPWR_c_351_n 0.0163608f $X=2.745 $Y=2.55 $X2=0 $Y2=0
cc_199 N_A_37_57#_c_270_n N_VPWR_c_351_n 0.016545f $X=2.575 $Y=2.105 $X2=0 $Y2=0
cc_200 N_A_37_57#_c_269_n N_VPWR_c_352_n 0.021949f $X=0.89 $Y=2.195 $X2=0 $Y2=0
cc_201 N_A_37_57#_M1003_g N_VPWR_c_354_n 0.00809503f $X=2.745 $Y=2.55 $X2=0
+ $Y2=0
cc_202 N_A_37_57#_M1003_g N_VPWR_c_348_n 0.0150743f $X=2.745 $Y=2.55 $X2=0 $Y2=0
cc_203 N_A_37_57#_c_269_n N_VPWR_c_348_n 0.0124703f $X=0.89 $Y=2.195 $X2=0 $Y2=0
cc_204 N_A_37_57#_c_270_n A_256_410# 0.00595227f $X=2.575 $Y=2.105 $X2=-0.19
+ $Y2=-0.245
cc_205 N_A_37_57#_c_270_n A_360_410# 0.00671538f $X=2.575 $Y=2.105 $X2=-0.19
+ $Y2=-0.245
cc_206 N_A_37_57#_c_255_n N_X_c_385_n 0.0113995f $X=2.505 $Y=0.78 $X2=0 $Y2=0
cc_207 N_A_37_57#_M1003_g X 0.00363627f $X=2.745 $Y=2.55 $X2=0 $Y2=0
cc_208 N_A_37_57#_c_258_n X 5.77237e-19 $X=2.77 $Y=1.6 $X2=0 $Y2=0
cc_209 N_A_37_57#_c_270_n X 0.00800963f $X=2.575 $Y=2.105 $X2=0 $Y2=0
cc_210 N_A_37_57#_c_262_n X 0.00722769f $X=2.66 $Y=2.02 $X2=0 $Y2=0
cc_211 N_A_37_57#_c_255_n N_X_c_386_n 0.0215046f $X=2.505 $Y=0.78 $X2=0 $Y2=0
cc_212 N_A_37_57#_M1003_g N_X_c_386_n 0.0058106f $X=2.745 $Y=2.55 $X2=0 $Y2=0
cc_213 N_A_37_57#_c_260_n N_X_c_386_n 0.0482504f $X=2.765 $Y=1.095 $X2=0 $Y2=0
cc_214 N_A_37_57#_c_262_n N_X_c_386_n 0.0111464f $X=2.66 $Y=2.02 $X2=0 $Y2=0
cc_215 N_A_37_57#_c_259_n N_A_140_57#_c_404_n 0.00190863f $X=0.175 $Y=1.975
+ $X2=0 $Y2=0
cc_216 N_A_37_57#_c_263_n N_A_140_57#_c_404_n 0.0179795f $X=0.33 $Y=0.495 $X2=0
+ $Y2=0
cc_217 N_A_37_57#_c_260_n N_A_140_57#_c_405_n 5.26873e-19 $X=2.765 $Y=1.095
+ $X2=0 $Y2=0
cc_218 N_A_37_57#_c_259_n N_A_140_57#_c_406_n 0.00692851f $X=0.175 $Y=1.975
+ $X2=0 $Y2=0
cc_219 N_A_37_57#_c_255_n N_VGND_c_441_n 0.015388f $X=2.505 $Y=0.78 $X2=0 $Y2=0
cc_220 N_A_37_57#_c_263_n N_VGND_c_442_n 0.0263576f $X=0.33 $Y=0.495 $X2=0 $Y2=0
cc_221 N_A_37_57#_c_255_n N_VGND_c_443_n 0.00947719f $X=2.505 $Y=0.78 $X2=0
+ $Y2=0
cc_222 N_A_37_57#_c_257_n N_VGND_c_443_n 5.84996e-19 $X=2.685 $Y=0.93 $X2=0
+ $Y2=0
cc_223 N_A_37_57#_c_255_n N_VGND_c_444_n 0.0180243f $X=2.505 $Y=0.78 $X2=0 $Y2=0
cc_224 N_A_37_57#_c_257_n N_VGND_c_444_n 7.94744e-19 $X=2.685 $Y=0.93 $X2=0
+ $Y2=0
cc_225 N_A_37_57#_c_263_n N_VGND_c_444_n 0.0154994f $X=0.33 $Y=0.495 $X2=0 $Y2=0
cc_226 N_VPWR_c_351_n X 0.0179162f $X=2.48 $Y=2.535 $X2=0 $Y2=0
cc_227 N_VPWR_c_354_n X 0.0231266f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_228 N_VPWR_c_348_n X 0.0132718f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_229 N_X_c_385_n N_VGND_c_441_n 0.0154769f $X=3.08 $Y=0.495 $X2=0 $Y2=0
cc_230 N_X_c_385_n N_VGND_c_443_n 0.0233657f $X=3.08 $Y=0.495 $X2=0 $Y2=0
cc_231 N_X_c_385_n N_VGND_c_444_n 0.0134749f $X=3.08 $Y=0.495 $X2=0 $Y2=0
cc_232 N_A_140_57#_c_404_n N_VGND_c_439_n 0.00151838f $X=0.84 $Y=0.495 $X2=0
+ $Y2=0
cc_233 N_A_140_57#_c_405_n N_VGND_c_439_n 0.0237709f $X=1.695 $Y=0.86 $X2=0
+ $Y2=0
cc_234 N_A_140_57#_c_407_n N_VGND_c_439_n 0.0120942f $X=1.86 $Y=0.495 $X2=0
+ $Y2=0
cc_235 N_A_140_57#_c_407_n N_VGND_c_440_n 0.0166382f $X=1.86 $Y=0.495 $X2=0
+ $Y2=0
cc_236 N_A_140_57#_c_407_n N_VGND_c_441_n 0.0179429f $X=1.86 $Y=0.495 $X2=0
+ $Y2=0
cc_237 N_A_140_57#_c_404_n N_VGND_c_442_n 0.0220321f $X=0.84 $Y=0.495 $X2=0
+ $Y2=0
cc_238 N_A_140_57#_c_404_n N_VGND_c_444_n 0.0125808f $X=0.84 $Y=0.495 $X2=0
+ $Y2=0
cc_239 N_A_140_57#_c_405_n N_VGND_c_444_n 0.0124074f $X=1.695 $Y=0.86 $X2=0
+ $Y2=0
cc_240 N_A_140_57#_c_407_n N_VGND_c_444_n 0.00948536f $X=1.86 $Y=0.495 $X2=0
+ $Y2=0
