* File: sky130_fd_sc_lp__decap_3.pxi.spice
* Created: Wed Sep  2 09:41:53 2020
* 
x_PM_SKY130_FD_SC_LP__DECAP_3%VGND N_VGND_M1001_s N_VGND_c_21_n N_VGND_M1000_g
+ N_VGND_c_22_n N_VGND_c_23_n N_VGND_c_24_n N_VGND_c_25_n N_VGND_c_26_n VGND
+ N_VGND_c_27_n N_VGND_c_28_n PM_SKY130_FD_SC_LP__DECAP_3%VGND
x_PM_SKY130_FD_SC_LP__DECAP_3%VPWR N_VPWR_M1000_s N_VPWR_c_48_n N_VPWR_M1001_g
+ N_VPWR_c_52_n N_VPWR_c_53_n N_VPWR_c_54_n N_VPWR_c_49_n N_VPWR_c_50_n VPWR
+ N_VPWR_c_56_n N_VPWR_c_51_n PM_SKY130_FD_SC_LP__DECAP_3%VPWR
cc_1 VNB N_VGND_c_21_n 0.012024f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.135
cc_2 VNB N_VGND_c_22_n 0.012758f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.085
cc_3 VNB N_VGND_c_23_n 0.0667513f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.48
cc_4 VNB N_VGND_c_24_n 0.0124146f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.085
cc_5 VNB N_VGND_c_25_n 0.018083f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.46
cc_6 VNB N_VGND_c_26_n 0.0043934f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.77
cc_7 VNB N_VGND_c_27_n 0.0121627f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=0
cc_8 VNB N_VGND_c_28_n 0.113154f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0
cc_9 VNB N_VPWR_c_48_n 0.0882018f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.135
cc_10 VNB N_VPWR_c_49_n 0.0258712f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.77
cc_11 VNB N_VPWR_c_50_n 0.0186797f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=0
cc_12 VNB N_VPWR_c_51_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0
cc_13 VPB N_VGND_c_21_n 0.0833936f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.135
cc_14 VPB N_VGND_c_26_n 0.0138032f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.77
cc_15 VPB N_VPWR_c_52_n 0.0103989f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.085
cc_16 VPB N_VPWR_c_53_n 0.0424658f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.48
cc_17 VPB N_VPWR_c_54_n 0.0144866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_18 VPB N_VPWR_c_49_n 0.0607744f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.77
cc_19 VPB N_VPWR_c_56_n 0.0124809f $X=-0.19 $Y=1.655 $X2=0.25 $Y2=0
cc_20 VPB N_VPWR_c_51_n 0.0485751f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=0
cc_21 N_VGND_c_21_n N_VPWR_c_48_n 0.0107128f $X=0.66 $Y=2.135 $X2=0 $Y2=0
cc_22 N_VGND_c_23_n N_VPWR_c_48_n 0.0411391f $X=0.335 $Y=0.48 $X2=0 $Y2=0
cc_23 N_VGND_c_25_n N_VPWR_c_48_n 0.0160601f $X=1.115 $Y=0.46 $X2=0 $Y2=0
cc_24 N_VGND_c_26_n N_VPWR_c_48_n 0.00102763f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_25 N_VGND_c_27_n N_VPWR_c_48_n 0.017526f $X=0.95 $Y=0 $X2=0 $Y2=0
cc_26 N_VGND_c_28_n N_VPWR_c_48_n 0.019115f $X=1.2 $Y=0 $X2=0 $Y2=0
cc_27 N_VGND_c_21_n N_VPWR_c_53_n 0.0290763f $X=0.66 $Y=2.135 $X2=0 $Y2=0
cc_28 N_VGND_c_26_n N_VPWR_c_53_n 0.0205444f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_29 N_VGND_c_21_n N_VPWR_c_49_n 0.0505388f $X=0.66 $Y=2.135 $X2=0 $Y2=0
cc_30 N_VGND_c_23_n N_VPWR_c_49_n 0.017965f $X=0.335 $Y=0.48 $X2=0 $Y2=0
cc_31 N_VGND_c_26_n N_VPWR_c_49_n 0.0215873f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_32 N_VGND_c_21_n N_VPWR_c_50_n 0.00139445f $X=0.66 $Y=2.135 $X2=0 $Y2=0
cc_33 N_VGND_c_23_n N_VPWR_c_50_n 0.0297314f $X=0.335 $Y=0.48 $X2=0 $Y2=0
cc_34 N_VGND_c_25_n N_VPWR_c_50_n 0.0151419f $X=1.115 $Y=0.46 $X2=0 $Y2=0
cc_35 N_VGND_c_28_n N_VPWR_c_50_n 0.00916521f $X=1.2 $Y=0 $X2=0 $Y2=0
cc_36 N_VGND_c_21_n N_VPWR_c_56_n 0.0179162f $X=0.66 $Y=2.135 $X2=0 $Y2=0
cc_37 N_VGND_c_21_n N_VPWR_c_51_n 0.0279709f $X=0.66 $Y=2.135 $X2=0 $Y2=0
