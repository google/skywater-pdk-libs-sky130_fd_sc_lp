* NGSPICE file created from sky130_fd_sc_lp__dlrbp_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlrbp_lp D GATE RESET_B VGND VNB VPB VPWR Q Q_N
M1000 a_272_419# GATE a_272_112# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1001 VGND a_1028_23# a_1701_74# VNB nshort w=420000u l=150000u
+  ad=6.258e+11p pd=7.18e+06u as=8.82e+10p ps=1.26e+06u
M1002 VPWR a_1028_23# a_955_367# VPB phighvt w=1e+06u l=250000u
+  ad=1.553e+12p pd=1.337e+07u as=3.65e+11p ps=2.73e+06u
M1003 Q a_1028_23# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1004 VPWR a_1028_23# a_1614_74# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1005 a_1431_49# a_1028_23# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1006 VGND D a_114_112# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 a_778_49# a_272_419# a_692_367# VPB phighvt w=1e+06u l=250000u
+  ad=5.75e+11p pd=3.15e+06u as=2.4e+11p ps=2.48e+06u
M1008 a_272_112# GATE VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_955_367# a_455_49# a_778_49# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_272_419# a_542_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1011 VPWR a_272_419# a_455_49# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1012 Q_N a_1614_74# a_1859_74# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1013 a_272_419# GATE VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1014 a_114_112# D a_27_112# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1015 VPWR RESET_B a_1028_23# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=4.69e+11p ps=3.08e+06u
M1016 a_542_49# a_272_419# a_455_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1017 a_1859_74# a_1614_74# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_700_49# a_27_112# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1019 a_944_49# a_272_419# a_778_49# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=2.856e+11p ps=2.2e+06u
M1020 a_1273_49# a_778_49# a_1028_23# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1021 a_1028_23# a_778_49# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q_N a_1614_74# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1023 VGND RESET_B a_1273_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Q a_1028_23# a_1431_49# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1025 a_692_367# a_27_112# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_778_49# a_455_49# a_700_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR D a_27_112# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1028 VGND a_1028_23# a_944_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1701_74# a_1028_23# a_1614_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends

