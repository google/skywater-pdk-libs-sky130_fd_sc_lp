* File: sky130_fd_sc_lp__a2bb2oi_2.pxi.spice
* Created: Fri Aug 28 09:56:45 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%B1 N_B1_M1015_g N_B1_M1002_g N_B1_M1018_g
+ N_B1_M1011_g N_B1_c_108_n N_B1_c_109_n N_B1_c_114_n N_B1_c_115_n N_B1_c_110_n
+ N_B1_c_111_n B1 B1 B1 PM_SKY130_FD_SC_LP__A2BB2OI_2%B1
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%B2 N_B2_M1004_g N_B2_M1005_g N_B2_M1008_g
+ N_B2_M1012_g B2 N_B2_c_196_n N_B2_c_193_n PM_SKY130_FD_SC_LP__A2BB2OI_2%B2
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%A_459_39# N_A_459_39#_M1010_s
+ N_A_459_39#_M1000_s N_A_459_39#_M1006_d N_A_459_39#_M1003_g
+ N_A_459_39#_M1007_g N_A_459_39#_c_243_n N_A_459_39#_c_244_n
+ N_A_459_39#_M1009_g N_A_459_39#_M1016_g N_A_459_39#_c_246_n
+ N_A_459_39#_c_247_n N_A_459_39#_c_248_n N_A_459_39#_c_249_n
+ N_A_459_39#_c_250_n N_A_459_39#_c_251_n N_A_459_39#_c_252_n
+ N_A_459_39#_c_253_n N_A_459_39#_c_254_n N_A_459_39#_c_255_n
+ N_A_459_39#_c_260_n N_A_459_39#_c_261_n N_A_459_39#_c_336_p
+ N_A_459_39#_c_256_n N_A_459_39#_c_257_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_2%A_459_39#
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%A1_N N_A1_N_M1010_g N_A1_N_M1001_g
+ N_A1_N_M1019_g N_A1_N_M1013_g A1_N N_A1_N_c_361_n N_A1_N_c_362_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_2%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%A2_N N_A2_N_c_417_n N_A2_N_M1000_g
+ N_A2_N_M1006_g N_A2_N_c_419_n N_A2_N_M1017_g N_A2_N_M1014_g N_A2_N_c_421_n
+ A2_N A2_N N_A2_N_c_423_n PM_SKY130_FD_SC_LP__A2BB2OI_2%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%A_30_367# N_A_30_367#_M1002_d
+ N_A_30_367#_M1005_d N_A_30_367#_M1011_d N_A_30_367#_M1016_d
+ N_A_30_367#_c_463_n N_A_30_367#_c_464_n N_A_30_367#_c_474_n
+ N_A_30_367#_c_478_n N_A_30_367#_c_465_n N_A_30_367#_c_489_n
+ N_A_30_367#_c_504_p N_A_30_367#_c_466_n N_A_30_367#_c_467_n
+ N_A_30_367#_c_468_n N_A_30_367#_c_485_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_2%A_30_367#
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%VPWR N_VPWR_M1002_s N_VPWR_M1012_s
+ N_VPWR_M1001_d N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n VPWR
+ N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_524_n
+ N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%Y N_Y_M1004_d N_Y_M1003_d N_Y_M1007_s
+ N_Y_c_607_n N_Y_c_601_n N_Y_c_602_n N_Y_c_605_n N_Y_c_628_n N_Y_c_603_n
+ N_Y_c_638_n Y Y N_Y_c_604_n PM_SKY130_FD_SC_LP__A2BB2OI_2%Y
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%A_699_367# N_A_699_367#_M1001_s
+ N_A_699_367#_M1013_s N_A_699_367#_M1014_s N_A_699_367#_c_659_n
+ N_A_699_367#_c_660_n N_A_699_367#_c_664_n N_A_699_367#_c_666_n
+ N_A_699_367#_c_693_n N_A_699_367#_c_667_n N_A_699_367#_c_661_n
+ N_A_699_367#_c_662_n PM_SKY130_FD_SC_LP__A2BB2OI_2%A_699_367#
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%VGND N_VGND_M1015_d N_VGND_M1018_d
+ N_VGND_M1009_s N_VGND_M1019_d N_VGND_M1017_d N_VGND_c_699_n N_VGND_c_700_n
+ N_VGND_c_701_n N_VGND_c_702_n N_VGND_c_703_n N_VGND_c_704_n VGND
+ N_VGND_c_705_n N_VGND_c_706_n N_VGND_c_707_n N_VGND_c_708_n N_VGND_c_709_n
+ N_VGND_c_710_n N_VGND_c_711_n PM_SKY130_FD_SC_LP__A2BB2OI_2%VGND
x_PM_SKY130_FD_SC_LP__A2BB2OI_2%A_113_65# N_A_113_65#_M1015_s
+ N_A_113_65#_M1008_s N_A_113_65#_c_777_n N_A_113_65#_c_778_n
+ N_A_113_65#_c_779_n N_A_113_65#_c_784_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_2%A_113_65#
cc_1 VNB N_B1_M1015_g 0.022827f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.745
cc_2 VNB N_B1_M1002_g 0.00221461f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_3 VNB N_B1_M1018_g 0.0217405f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.745
cc_4 VNB N_B1_c_108_n 0.0133945f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.5
cc_5 VNB N_B1_c_109_n 0.0369181f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.46
cc_6 VNB N_B1_c_110_n 0.00225608f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.51
cc_7 VNB N_B1_c_111_n 0.0256594f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.51
cc_8 VNB N_B2_M1004_g 0.0198827f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.745
cc_9 VNB N_B2_M1008_g 0.0203074f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.745
cc_10 VNB N_B2_c_193_n 0.0333769f $X=-0.19 $Y=-0.245 $X2=1.737 $Y2=1.655
cc_11 VNB N_A_459_39#_M1003_g 0.0243953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_459_39#_M1007_g 0.00411396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_459_39#_c_243_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.5
cc_14 VNB N_A_459_39#_c_244_n 0.0180861f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.46
cc_15 VNB N_A_459_39#_M1016_g 0.00425929f $X=-0.19 $Y=-0.245 $X2=1.737 $Y2=1.92
cc_16 VNB N_A_459_39#_c_246_n 0.0160355f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.51
cc_17 VNB N_A_459_39#_c_247_n 0.00535129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_459_39#_c_248_n 0.00891687f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.655
cc_19 VNB N_A_459_39#_c_249_n 0.00766626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_459_39#_c_250_n 0.00627546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_459_39#_c_251_n 6.24889e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_459_39#_c_252_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.625
cc_23 VNB N_A_459_39#_c_253_n 0.00115399f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.675
cc_24 VNB N_A_459_39#_c_254_n 0.00634013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_459_39#_c_255_n 0.0038594f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=2.02
cc_26 VNB N_A_459_39#_c_256_n 0.00168223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_459_39#_c_257_n 0.0402148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_N_M1010_g 0.0228515f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.745
cc_29 VNB N_A1_N_M1019_g 0.0189298f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.745
cc_30 VNB N_A1_N_c_361_n 0.00304874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A1_N_c_362_n 0.0397838f $X=-0.19 $Y=-0.245 $X2=1.737 $Y2=1.655
cc_32 VNB N_A2_N_c_417_n 0.0156569f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.295
cc_33 VNB N_A2_N_M1006_g 0.0119872f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_34 VNB N_A2_N_c_419_n 0.0475088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_N_M1014_g 0.00303933f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=2.465
cc_36 VNB N_A2_N_c_421_n 0.00537411f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.5
cc_37 VNB A2_N 0.028155f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.5
cc_38 VNB N_A2_N_c_423_n 0.0203221f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.92
cc_39 VNB N_VPWR_c_524_n 0.243291f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.02
cc_40 VNB N_Y_c_601_n 0.0112625f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=2.465
cc_41 VNB N_Y_c_602_n 0.00232524f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=2.465
cc_42 VNB N_Y_c_603_n 0.00238193f $X=-0.19 $Y=-0.245 $X2=1.737 $Y2=1.655
cc_43 VNB N_Y_c_604_n 0.00209028f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_44 VNB N_VGND_c_699_n 0.0113841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_700_n 0.0464301f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.5
cc_46 VNB N_VGND_c_701_n 0.00455363f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.625
cc_47 VNB N_VGND_c_702_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.51
cc_48 VNB N_VGND_c_703_n 0.0161518f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.51
cc_49 VNB N_VGND_c_704_n 0.0350549f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.655
cc_50 VNB N_VGND_c_705_n 0.0389003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_706_n 0.0410254f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.51
cc_52 VNB N_VGND_c_707_n 0.0143188f $X=-0.19 $Y=-0.245 $X2=0.767 $Y2=2.02
cc_53 VNB N_VGND_c_708_n 0.0144602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_709_n 0.00581671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_710_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_711_n 0.31983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_113_65#_c_777_n 0.00468699f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.345
cc_58 VNB N_A_113_65#_c_778_n 0.00499024f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.745
cc_59 VNB N_A_113_65#_c_779_n 0.00221252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VPB N_B1_M1002_g 0.026333f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_61 VPB N_B1_M1011_g 0.0200063f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=2.465
cc_62 VPB N_B1_c_114_n 0.00136397f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.92
cc_63 VPB N_B1_c_115_n 0.00143908f $X=-0.19 $Y=1.655 $X2=1.737 $Y2=1.92
cc_64 VPB N_B1_c_111_n 0.00647089f $X=-0.19 $Y=1.655 $X2=1.85 $Y2=1.51
cc_65 VPB N_B2_M1005_g 0.0184684f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_66 VPB N_B2_M1012_g 0.0202431f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=2.465
cc_67 VPB N_B2_c_196_n 0.00259635f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.92
cc_68 VPB N_B2_c_193_n 0.00485967f $X=-0.19 $Y=1.655 $X2=1.737 $Y2=1.655
cc_69 VPB N_A_459_39#_M1007_g 0.0199701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_459_39#_M1016_g 0.0239746f $X=-0.19 $Y=1.655 $X2=1.737 $Y2=1.92
cc_71 VPB N_A_459_39#_c_260_n 0.00739529f $X=-0.19 $Y=1.655 $X2=0.767 $Y2=2.02
cc_72 VPB N_A_459_39#_c_261_n 8.26403e-19 $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.02
cc_73 VPB N_A1_N_M1001_g 0.0222503f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_74 VPB N_A1_N_M1013_g 0.0174026f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=2.465
cc_75 VPB N_A1_N_c_361_n 0.00385574f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A1_N_c_362_n 0.00913024f $X=-0.19 $Y=1.655 $X2=1.737 $Y2=1.655
cc_77 VPB N_A2_N_M1006_g 0.0188143f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_78 VPB N_A2_N_M1014_g 0.026001f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=2.465
cc_79 VPB A2_N 0.0135375f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.5
cc_80 VPB N_A_30_367#_c_463_n 0.0211977f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=2.465
cc_81 VPB N_A_30_367#_c_464_n 0.0233935f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.46
cc_82 VPB N_A_30_367#_c_465_n 0.0033084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A_30_367#_c_466_n 0.00206973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_30_367#_c_467_n 0.0151077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A_30_367#_c_468_n 0.00717518f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.46
cc_86 VPB N_VPWR_c_525_n 4.14e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_526_n 0.00504096f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_527_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.46
cc_89 VPB N_VPWR_c_528_n 0.0158532f $X=-0.19 $Y=1.655 $X2=1.737 $Y2=1.655
cc_90 VPB N_VPWR_c_529_n 0.0167565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_530_n 0.0512789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_531_n 0.0394434f $X=-0.19 $Y=1.655 $X2=0.767 $Y2=2.02
cc_93 VPB N_VPWR_c_524_n 0.064663f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.02
cc_94 VPB N_VPWR_c_533_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.02
cc_95 VPB N_VPWR_c_534_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_535_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_Y_c_605_n 7.44467e-19 $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.5
cc_98 VPB N_Y_c_603_n 0.00138773f $X=-0.19 $Y=1.655 $X2=1.737 $Y2=1.655
cc_99 VPB N_A_699_367#_c_659_n 0.00340764f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=0.745
cc_100 VPB N_A_699_367#_c_660_n 0.00909614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_699_367#_c_661_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.46
cc_102 VPB N_A_699_367#_c_662_n 0.0384572f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.625
cc_103 N_B1_M1015_g N_B2_M1004_g 0.0286544f $X=0.49 $Y=0.745 $X2=0 $Y2=0
cc_104 N_B1_M1002_g N_B2_M1005_g 0.0286544f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_105 B1 N_B2_M1005_g 0.0136686f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_106 N_B1_M1018_g N_B2_M1008_g 0.0262771f $X=1.86 $Y=0.745 $X2=0 $Y2=0
cc_107 N_B1_M1011_g N_B2_M1012_g 0.0353167f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_108 N_B1_c_115_n N_B2_M1012_g 0.00321181f $X=1.737 $Y=1.92 $X2=0 $Y2=0
cc_109 B1 N_B2_M1012_g 0.012487f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_110 N_B1_c_108_n N_B2_c_196_n 0.0162461f $X=0.55 $Y=1.5 $X2=0 $Y2=0
cc_111 N_B1_c_109_n N_B2_c_196_n 2.84562e-19 $X=0.4 $Y=1.46 $X2=0 $Y2=0
cc_112 N_B1_c_114_n N_B2_c_196_n 0.00927785f $X=0.64 $Y=1.92 $X2=0 $Y2=0
cc_113 N_B1_c_110_n N_B2_c_196_n 0.026767f $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_114 N_B1_c_111_n N_B2_c_196_n 2.70823e-19 $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_115 B1 N_B2_c_196_n 0.0348015f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_116 N_B1_c_108_n N_B2_c_193_n 0.00311053f $X=0.55 $Y=1.5 $X2=0 $Y2=0
cc_117 N_B1_c_109_n N_B2_c_193_n 0.0286544f $X=0.4 $Y=1.46 $X2=0 $Y2=0
cc_118 N_B1_c_114_n N_B2_c_193_n 0.0046388f $X=0.64 $Y=1.92 $X2=0 $Y2=0
cc_119 N_B1_c_110_n N_B2_c_193_n 0.00321181f $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_120 N_B1_c_111_n N_B2_c_193_n 0.0174855f $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_121 B1 N_B2_c_193_n 5.84466e-19 $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_122 N_B1_M1018_g N_A_459_39#_M1003_g 0.0245792f $X=1.86 $Y=0.745 $X2=0 $Y2=0
cc_123 N_B1_c_111_n N_A_459_39#_M1003_g 0.0165666f $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_124 N_B1_c_115_n N_A_459_39#_M1007_g 5.31474e-19 $X=1.737 $Y=1.92 $X2=0 $Y2=0
cc_125 N_B1_M1011_g N_A_459_39#_c_247_n 0.0165666f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B1_c_110_n N_A_459_39#_c_247_n 0.00100492f $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_127 B1 N_A_30_367#_M1005_d 0.00334146f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_128 N_B1_M1002_g N_A_30_367#_c_463_n 0.00241112f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_129 N_B1_c_108_n N_A_30_367#_c_463_n 0.0109602f $X=0.55 $Y=1.5 $X2=0 $Y2=0
cc_130 N_B1_c_109_n N_A_30_367#_c_463_n 0.00332032f $X=0.4 $Y=1.46 $X2=0 $Y2=0
cc_131 N_B1_c_114_n N_A_30_367#_c_463_n 0.00432257f $X=0.64 $Y=1.92 $X2=0 $Y2=0
cc_132 N_B1_M1002_g N_A_30_367#_c_474_n 0.0142333f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_133 N_B1_c_108_n N_A_30_367#_c_474_n 0.00339833f $X=0.55 $Y=1.5 $X2=0 $Y2=0
cc_134 N_B1_c_114_n N_A_30_367#_c_474_n 0.00988447f $X=0.64 $Y=1.92 $X2=0 $Y2=0
cc_135 B1 N_A_30_367#_c_474_n 0.0144893f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_136 N_B1_M1011_g N_A_30_367#_c_478_n 0.0156363f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_137 N_B1_c_115_n N_A_30_367#_c_478_n 0.0184178f $X=1.737 $Y=1.92 $X2=0 $Y2=0
cc_138 N_B1_c_110_n N_A_30_367#_c_478_n 0.00311532f $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_139 N_B1_c_111_n N_A_30_367#_c_478_n 4.56216e-19 $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_140 B1 N_A_30_367#_c_478_n 0.0184648f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_141 N_B1_M1011_g N_A_30_367#_c_465_n 3.34222e-19 $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_142 N_B1_c_115_n N_A_30_367#_c_465_n 0.00379586f $X=1.737 $Y=1.92 $X2=0 $Y2=0
cc_143 B1 N_A_30_367#_c_485_n 0.0136549f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_144 N_B1_c_114_n N_VPWR_M1002_s 0.00213723f $X=0.64 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_145 B1 N_VPWR_M1002_s 0.00282854f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_146 N_B1_c_115_n N_VPWR_M1012_s 0.00455943f $X=1.737 $Y=1.92 $X2=0 $Y2=0
cc_147 B1 N_VPWR_M1012_s 0.00358643f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_148 N_B1_M1002_g N_VPWR_c_525_n 0.011946f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_149 N_B1_M1011_g N_VPWR_c_526_n 0.00611917f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_150 N_B1_M1002_g N_VPWR_c_528_n 0.00486043f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_151 N_B1_M1011_g N_VPWR_c_530_n 0.00585385f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_152 N_B1_M1002_g N_VPWR_c_524_n 0.00919377f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_153 N_B1_M1011_g N_VPWR_c_524_n 0.0111412f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_154 N_B1_M1018_g N_Y_c_607_n 6.08169e-19 $X=1.86 $Y=0.745 $X2=0 $Y2=0
cc_155 N_B1_M1018_g N_Y_c_601_n 0.0148518f $X=1.86 $Y=0.745 $X2=0 $Y2=0
cc_156 N_B1_c_110_n N_Y_c_601_n 0.0310439f $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_157 N_B1_c_111_n N_Y_c_601_n 0.00476197f $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_158 B1 N_Y_c_601_n 0.00392693f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_159 N_B1_M1015_g N_Y_c_602_n 3.20368e-19 $X=0.49 $Y=0.745 $X2=0 $Y2=0
cc_160 N_B1_c_115_n N_Y_c_605_n 5.75163e-19 $X=1.737 $Y=1.92 $X2=0 $Y2=0
cc_161 N_B1_c_115_n N_Y_c_603_n 0.0042283f $X=1.737 $Y=1.92 $X2=0 $Y2=0
cc_162 N_B1_c_110_n N_Y_c_603_n 0.00764285f $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_163 N_B1_c_111_n N_Y_c_603_n 4.27505e-19 $X=1.85 $Y=1.51 $X2=0 $Y2=0
cc_164 N_B1_M1015_g N_VGND_c_700_n 0.00783332f $X=0.49 $Y=0.745 $X2=0 $Y2=0
cc_165 N_B1_c_108_n N_VGND_c_700_n 0.0128647f $X=0.55 $Y=1.5 $X2=0 $Y2=0
cc_166 N_B1_c_109_n N_VGND_c_700_n 0.00429667f $X=0.4 $Y=1.46 $X2=0 $Y2=0
cc_167 N_B1_M1018_g N_VGND_c_701_n 0.00518042f $X=1.86 $Y=0.745 $X2=0 $Y2=0
cc_168 N_B1_M1015_g N_VGND_c_705_n 0.00499542f $X=0.49 $Y=0.745 $X2=0 $Y2=0
cc_169 N_B1_M1018_g N_VGND_c_705_n 0.00453911f $X=1.86 $Y=0.745 $X2=0 $Y2=0
cc_170 N_B1_M1015_g N_VGND_c_711_n 0.01008f $X=0.49 $Y=0.745 $X2=0 $Y2=0
cc_171 N_B1_M1018_g N_VGND_c_711_n 0.00866891f $X=1.86 $Y=0.745 $X2=0 $Y2=0
cc_172 N_B1_M1015_g N_A_113_65#_c_777_n 8.9451e-19 $X=0.49 $Y=0.745 $X2=0 $Y2=0
cc_173 N_B1_c_108_n N_A_113_65#_c_777_n 0.013331f $X=0.55 $Y=1.5 $X2=0 $Y2=0
cc_174 N_B1_M1018_g N_A_113_65#_c_778_n 0.00293805f $X=1.86 $Y=0.745 $X2=0 $Y2=0
cc_175 N_B1_M1015_g N_A_113_65#_c_779_n 5.28944e-19 $X=0.49 $Y=0.745 $X2=0 $Y2=0
cc_176 N_B1_M1018_g N_A_113_65#_c_784_n 0.00569398f $X=1.86 $Y=0.745 $X2=0 $Y2=0
cc_177 N_B2_M1005_g N_A_30_367#_c_474_n 0.0122129f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_178 N_B2_M1012_g N_A_30_367#_c_478_n 0.013664f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_179 N_B2_M1005_g N_VPWR_c_525_n 0.0104601f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_180 N_B2_M1012_g N_VPWR_c_525_n 6.11746e-19 $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B2_M1012_g N_VPWR_c_526_n 0.00662445f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B2_M1005_g N_VPWR_c_529_n 0.00486043f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B2_M1012_g N_VPWR_c_529_n 0.00585385f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_184 N_B2_M1005_g N_VPWR_c_524_n 0.00824727f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_185 N_B2_M1012_g N_VPWR_c_524_n 0.0111705f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B2_M1004_g N_Y_c_607_n 0.00506691f $X=0.92 $Y=0.745 $X2=0 $Y2=0
cc_187 N_B2_M1008_g N_Y_c_607_n 0.00668486f $X=1.35 $Y=0.745 $X2=0 $Y2=0
cc_188 N_B2_M1008_g N_Y_c_601_n 0.00957731f $X=1.35 $Y=0.745 $X2=0 $Y2=0
cc_189 N_B2_c_196_n N_Y_c_601_n 0.00845751f $X=1.075 $Y=1.51 $X2=0 $Y2=0
cc_190 N_B2_M1004_g N_Y_c_602_n 0.00361035f $X=0.92 $Y=0.745 $X2=0 $Y2=0
cc_191 N_B2_M1008_g N_Y_c_602_n 0.0016917f $X=1.35 $Y=0.745 $X2=0 $Y2=0
cc_192 N_B2_c_196_n N_Y_c_602_n 0.0263959f $X=1.075 $Y=1.51 $X2=0 $Y2=0
cc_193 N_B2_c_193_n N_Y_c_602_n 0.00254355f $X=1.35 $Y=1.51 $X2=0 $Y2=0
cc_194 N_B2_M1004_g N_VGND_c_705_n 0.0030414f $X=0.92 $Y=0.745 $X2=0 $Y2=0
cc_195 N_B2_M1008_g N_VGND_c_705_n 0.0030414f $X=1.35 $Y=0.745 $X2=0 $Y2=0
cc_196 N_B2_M1004_g N_VGND_c_711_n 0.00435814f $X=0.92 $Y=0.745 $X2=0 $Y2=0
cc_197 N_B2_M1008_g N_VGND_c_711_n 0.0044277f $X=1.35 $Y=0.745 $X2=0 $Y2=0
cc_198 N_B2_M1004_g N_A_113_65#_c_777_n 8.30663e-19 $X=0.92 $Y=0.745 $X2=0 $Y2=0
cc_199 N_B2_M1004_g N_A_113_65#_c_778_n 0.0118256f $X=0.92 $Y=0.745 $X2=0 $Y2=0
cc_200 N_B2_M1008_g N_A_113_65#_c_778_n 0.0116012f $X=1.35 $Y=0.745 $X2=0 $Y2=0
cc_201 N_A_459_39#_c_249_n N_A1_N_M1010_g 0.00116512f $X=3.25 $Y=1.44 $X2=0
+ $Y2=0
cc_202 N_A_459_39#_c_250_n N_A1_N_M1010_g 0.0151939f $X=3.955 $Y=1.16 $X2=0
+ $Y2=0
cc_203 N_A_459_39#_c_252_n N_A1_N_M1010_g 8.28776e-19 $X=4.05 $Y=0.47 $X2=0
+ $Y2=0
cc_204 N_A_459_39#_c_253_n N_A1_N_M1010_g 0.00193172f $X=4.22 $Y=1.705 $X2=0
+ $Y2=0
cc_205 N_A_459_39#_c_257_n N_A1_N_M1010_g 0.00291799f $X=3.25 $Y=1.35 $X2=0
+ $Y2=0
cc_206 N_A_459_39#_c_261_n N_A1_N_M1001_g 5.04096e-19 $X=4.305 $Y=1.79 $X2=0
+ $Y2=0
cc_207 N_A_459_39#_c_252_n N_A1_N_M1019_g 8.28776e-19 $X=4.05 $Y=0.47 $X2=0
+ $Y2=0
cc_208 N_A_459_39#_c_253_n N_A1_N_M1019_g 0.00320692f $X=4.22 $Y=1.705 $X2=0
+ $Y2=0
cc_209 N_A_459_39#_c_254_n N_A1_N_M1019_g 0.00405091f $X=4.825 $Y=1.16 $X2=0
+ $Y2=0
cc_210 N_A_459_39#_c_255_n N_A1_N_M1019_g 0.00814406f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_211 N_A_459_39#_c_253_n N_A1_N_M1013_g 8.0536e-19 $X=4.22 $Y=1.705 $X2=0
+ $Y2=0
cc_212 N_A_459_39#_c_260_n N_A1_N_M1013_g 0.00373666f $X=4.785 $Y=1.79 $X2=0
+ $Y2=0
cc_213 N_A_459_39#_c_261_n N_A1_N_M1013_g 0.00428833f $X=4.305 $Y=1.79 $X2=0
+ $Y2=0
cc_214 N_A_459_39#_M1016_g N_A1_N_c_361_n 0.00538914f $X=2.8 $Y=2.465 $X2=0
+ $Y2=0
cc_215 N_A_459_39#_c_249_n N_A1_N_c_361_n 0.0151101f $X=3.25 $Y=1.44 $X2=0 $Y2=0
cc_216 N_A_459_39#_c_250_n N_A1_N_c_361_n 0.034619f $X=3.955 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_459_39#_c_253_n N_A1_N_c_361_n 0.0205211f $X=4.22 $Y=1.705 $X2=0
+ $Y2=0
cc_218 N_A_459_39#_c_261_n N_A1_N_c_361_n 0.0112511f $X=4.305 $Y=1.79 $X2=0
+ $Y2=0
cc_219 N_A_459_39#_c_257_n N_A1_N_c_361_n 0.00130038f $X=3.25 $Y=1.35 $X2=0
+ $Y2=0
cc_220 N_A_459_39#_c_249_n N_A1_N_c_362_n 6.18944e-19 $X=3.25 $Y=1.44 $X2=0
+ $Y2=0
cc_221 N_A_459_39#_c_250_n N_A1_N_c_362_n 0.00328782f $X=3.955 $Y=1.16 $X2=0
+ $Y2=0
cc_222 N_A_459_39#_c_253_n N_A1_N_c_362_n 0.0162294f $X=4.22 $Y=1.705 $X2=0
+ $Y2=0
cc_223 N_A_459_39#_c_255_n N_A1_N_c_362_n 0.00405355f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_224 N_A_459_39#_c_257_n N_A1_N_c_362_n 0.0172304f $X=3.25 $Y=1.35 $X2=0 $Y2=0
cc_225 N_A_459_39#_c_253_n N_A2_N_c_417_n 0.00285052f $X=4.22 $Y=1.705 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A_459_39#_c_254_n N_A2_N_c_417_n 0.0143103f $X=4.825 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_459_39#_c_256_n N_A2_N_c_417_n 8.13177e-19 $X=4.91 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_228 N_A_459_39#_c_260_n N_A2_N_M1006_g 0.0155177f $X=4.785 $Y=1.79 $X2=0
+ $Y2=0
cc_229 N_A_459_39#_c_254_n N_A2_N_c_419_n 0.00293735f $X=4.825 $Y=1.16 $X2=0
+ $Y2=0
cc_230 N_A_459_39#_c_260_n N_A2_N_c_419_n 0.00210337f $X=4.785 $Y=1.79 $X2=0
+ $Y2=0
cc_231 N_A_459_39#_c_260_n N_A2_N_M1014_g 0.00306651f $X=4.785 $Y=1.79 $X2=0
+ $Y2=0
cc_232 N_A_459_39#_c_254_n A2_N 0.00290947f $X=4.825 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A_459_39#_c_260_n A2_N 0.00390572f $X=4.785 $Y=1.79 $X2=0 $Y2=0
cc_234 N_A_459_39#_c_254_n N_A2_N_c_423_n 0.00168652f $X=4.825 $Y=1.16 $X2=0
+ $Y2=0
cc_235 N_A_459_39#_c_256_n N_A2_N_c_423_n 8.13177e-19 $X=4.91 $Y=0.47 $X2=0
+ $Y2=0
cc_236 N_A_459_39#_M1007_g N_A_30_367#_c_465_n 3.27305e-19 $X=2.37 $Y=2.465
+ $X2=0 $Y2=0
cc_237 N_A_459_39#_M1007_g N_A_30_367#_c_489_n 0.0115031f $X=2.37 $Y=2.465 $X2=0
+ $Y2=0
cc_238 N_A_459_39#_M1016_g N_A_30_367#_c_489_n 0.0114565f $X=2.8 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A_459_39#_M1016_g N_A_30_367#_c_467_n 0.00293325f $X=2.8 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_A_459_39#_c_246_n N_A_30_367#_c_467_n 0.00527123f $X=3.085 $Y=1.35
+ $X2=0 $Y2=0
cc_241 N_A_459_39#_c_249_n N_A_30_367#_c_467_n 0.00670541f $X=3.25 $Y=1.44 $X2=0
+ $Y2=0
cc_242 N_A_459_39#_c_257_n N_A_30_367#_c_467_n 7.12986e-19 $X=3.25 $Y=1.35 $X2=0
+ $Y2=0
cc_243 N_A_459_39#_M1007_g N_VPWR_c_530_n 0.00357877f $X=2.37 $Y=2.465 $X2=0
+ $Y2=0
cc_244 N_A_459_39#_M1016_g N_VPWR_c_530_n 0.00357877f $X=2.8 $Y=2.465 $X2=0
+ $Y2=0
cc_245 N_A_459_39#_M1006_d N_VPWR_c_524_n 0.00225186f $X=4.77 $Y=1.835 $X2=0
+ $Y2=0
cc_246 N_A_459_39#_M1007_g N_VPWR_c_524_n 0.00537654f $X=2.37 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_A_459_39#_M1016_g N_VPWR_c_524_n 0.00665089f $X=2.8 $Y=2.465 $X2=0
+ $Y2=0
cc_248 N_A_459_39#_M1003_g N_Y_c_601_n 0.0177379f $X=2.37 $Y=0.745 $X2=0 $Y2=0
cc_249 N_A_459_39#_M1007_g N_Y_c_605_n 0.00278152f $X=2.37 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A_459_39#_M1016_g N_Y_c_605_n 0.00276064f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A_459_39#_M1007_g N_Y_c_628_n 0.00802865f $X=2.37 $Y=2.465 $X2=0 $Y2=0
cc_252 N_A_459_39#_M1016_g N_Y_c_628_n 0.00846694f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_253 N_A_459_39#_M1003_g N_Y_c_603_n 0.00459881f $X=2.37 $Y=0.745 $X2=0 $Y2=0
cc_254 N_A_459_39#_M1007_g N_Y_c_603_n 0.00292236f $X=2.37 $Y=2.465 $X2=0 $Y2=0
cc_255 N_A_459_39#_c_243_n N_Y_c_603_n 0.0104412f $X=2.725 $Y=1.5 $X2=0 $Y2=0
cc_256 N_A_459_39#_c_244_n N_Y_c_603_n 6.73763e-19 $X=2.8 $Y=1.275 $X2=0 $Y2=0
cc_257 N_A_459_39#_M1016_g N_Y_c_603_n 0.0108421f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A_459_39#_c_248_n N_Y_c_603_n 0.00676826f $X=2.8 $Y=1.35 $X2=0 $Y2=0
cc_259 N_A_459_39#_c_249_n N_Y_c_603_n 0.0150678f $X=3.25 $Y=1.44 $X2=0 $Y2=0
cc_260 N_A_459_39#_c_257_n N_Y_c_603_n 5.20269e-19 $X=3.25 $Y=1.35 $X2=0 $Y2=0
cc_261 N_A_459_39#_c_244_n N_Y_c_638_n 0.00348978f $X=2.8 $Y=1.275 $X2=0 $Y2=0
cc_262 N_A_459_39#_c_251_n N_Y_c_638_n 0.00894079f $X=3.335 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_459_39#_M1003_g N_Y_c_604_n 8.74036e-19 $X=2.37 $Y=0.745 $X2=0 $Y2=0
cc_264 N_A_459_39#_c_244_n N_Y_c_604_n 0.0158663f $X=2.8 $Y=1.275 $X2=0 $Y2=0
cc_265 N_A_459_39#_c_260_n N_A_699_367#_M1013_s 0.00176461f $X=4.785 $Y=1.79
+ $X2=0 $Y2=0
cc_266 N_A_459_39#_c_260_n N_A_699_367#_c_664_n 0.00230453f $X=4.785 $Y=1.79
+ $X2=0 $Y2=0
cc_267 N_A_459_39#_c_261_n N_A_699_367#_c_664_n 0.00866254f $X=4.305 $Y=1.79
+ $X2=0 $Y2=0
cc_268 N_A_459_39#_c_260_n N_A_699_367#_c_666_n 0.0135055f $X=4.785 $Y=1.79
+ $X2=0 $Y2=0
cc_269 N_A_459_39#_M1006_d N_A_699_367#_c_667_n 0.00332344f $X=4.77 $Y=1.835
+ $X2=0 $Y2=0
cc_270 N_A_459_39#_c_336_p N_A_699_367#_c_667_n 0.0126348f $X=4.91 $Y=1.98 $X2=0
+ $Y2=0
cc_271 N_A_459_39#_c_250_n N_VGND_M1009_s 0.00450833f $X=3.955 $Y=1.16 $X2=0
+ $Y2=0
cc_272 N_A_459_39#_c_251_n N_VGND_M1009_s 0.00410939f $X=3.335 $Y=1.16 $X2=0
+ $Y2=0
cc_273 N_A_459_39#_c_254_n N_VGND_M1019_d 0.00180746f $X=4.825 $Y=1.16 $X2=0
+ $Y2=0
cc_274 N_A_459_39#_M1003_g N_VGND_c_701_n 0.0100135f $X=2.37 $Y=0.745 $X2=0
+ $Y2=0
cc_275 N_A_459_39#_c_244_n N_VGND_c_701_n 5.46016e-19 $X=2.8 $Y=1.275 $X2=0
+ $Y2=0
cc_276 N_A_459_39#_c_252_n N_VGND_c_702_n 0.0228652f $X=4.05 $Y=0.47 $X2=0 $Y2=0
cc_277 N_A_459_39#_c_254_n N_VGND_c_702_n 0.0163515f $X=4.825 $Y=1.16 $X2=0
+ $Y2=0
cc_278 N_A_459_39#_c_256_n N_VGND_c_702_n 0.0218329f $X=4.91 $Y=0.47 $X2=0 $Y2=0
cc_279 N_A_459_39#_c_256_n N_VGND_c_704_n 0.0270299f $X=4.91 $Y=0.47 $X2=0 $Y2=0
cc_280 N_A_459_39#_M1003_g N_VGND_c_706_n 0.00414769f $X=2.37 $Y=0.745 $X2=0
+ $Y2=0
cc_281 N_A_459_39#_c_244_n N_VGND_c_706_n 0.019155f $X=2.8 $Y=1.275 $X2=0 $Y2=0
cc_282 N_A_459_39#_c_246_n N_VGND_c_706_n 0.00518719f $X=3.085 $Y=1.35 $X2=0
+ $Y2=0
cc_283 N_A_459_39#_c_250_n N_VGND_c_706_n 0.0303575f $X=3.955 $Y=1.16 $X2=0
+ $Y2=0
cc_284 N_A_459_39#_c_251_n N_VGND_c_706_n 0.0212027f $X=3.335 $Y=1.16 $X2=0
+ $Y2=0
cc_285 N_A_459_39#_c_252_n N_VGND_c_706_n 0.0254628f $X=4.05 $Y=0.47 $X2=0 $Y2=0
cc_286 N_A_459_39#_c_257_n N_VGND_c_706_n 0.00143271f $X=3.25 $Y=1.35 $X2=0
+ $Y2=0
cc_287 N_A_459_39#_c_252_n N_VGND_c_707_n 0.0102275f $X=4.05 $Y=0.47 $X2=0 $Y2=0
cc_288 N_A_459_39#_c_256_n N_VGND_c_708_n 0.00913949f $X=4.91 $Y=0.47 $X2=0
+ $Y2=0
cc_289 N_A_459_39#_M1003_g N_VGND_c_711_n 0.00787505f $X=2.37 $Y=0.745 $X2=0
+ $Y2=0
cc_290 N_A_459_39#_c_244_n N_VGND_c_711_n 0.00939634f $X=2.8 $Y=1.275 $X2=0
+ $Y2=0
cc_291 N_A_459_39#_c_252_n N_VGND_c_711_n 0.00712543f $X=4.05 $Y=0.47 $X2=0
+ $Y2=0
cc_292 N_A_459_39#_c_256_n N_VGND_c_711_n 0.0063674f $X=4.91 $Y=0.47 $X2=0 $Y2=0
cc_293 N_A1_N_M1019_g N_A2_N_c_417_n 0.0204753f $X=4.265 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_294 N_A1_N_M1013_g N_A2_N_M1006_g 0.0204753f $X=4.265 $Y=2.465 $X2=0 $Y2=0
cc_295 N_A1_N_c_362_n N_A2_N_c_421_n 0.0204753f $X=4.265 $Y=1.51 $X2=0 $Y2=0
cc_296 N_A1_N_M1001_g N_A_30_367#_c_467_n 0.00389357f $X=3.835 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_A1_N_c_361_n N_A_30_367#_c_467_n 0.00255884f $X=3.79 $Y=1.51 $X2=0
+ $Y2=0
cc_298 N_A1_N_M1001_g N_VPWR_c_527_n 0.0139526f $X=3.835 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A1_N_M1013_g N_VPWR_c_527_n 0.0133041f $X=4.265 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A1_N_M1001_g N_VPWR_c_530_n 0.00486043f $X=3.835 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A1_N_M1013_g N_VPWR_c_531_n 0.00486043f $X=4.265 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A1_N_M1001_g N_VPWR_c_524_n 0.00954696f $X=3.835 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A1_N_M1013_g N_VPWR_c_524_n 0.0082726f $X=4.265 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A1_N_c_361_n N_A_699_367#_M1001_s 0.0027721f $X=3.79 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_305 N_A1_N_c_361_n N_A_699_367#_c_659_n 0.0172673f $X=3.79 $Y=1.51 $X2=0
+ $Y2=0
cc_306 N_A1_N_c_362_n N_A_699_367#_c_659_n 4.25149e-19 $X=4.265 $Y=1.51 $X2=0
+ $Y2=0
cc_307 N_A1_N_M1001_g N_A_699_367#_c_664_n 0.0122129f $X=3.835 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A1_N_M1013_g N_A_699_367#_c_664_n 0.0122411f $X=4.265 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A1_N_c_361_n N_A_699_367#_c_664_n 0.0109713f $X=3.79 $Y=1.51 $X2=0
+ $Y2=0
cc_310 N_A1_N_c_362_n N_A_699_367#_c_664_n 0.00303798f $X=4.265 $Y=1.51 $X2=0
+ $Y2=0
cc_311 N_A1_N_M1010_g N_VGND_c_702_n 5.06642e-19 $X=3.835 $Y=0.745 $X2=0 $Y2=0
cc_312 N_A1_N_M1019_g N_VGND_c_702_n 0.00999441f $X=4.265 $Y=0.745 $X2=0 $Y2=0
cc_313 N_A1_N_M1010_g N_VGND_c_706_n 0.011597f $X=3.835 $Y=0.745 $X2=0 $Y2=0
cc_314 N_A1_N_M1019_g N_VGND_c_706_n 5.09255e-19 $X=4.265 $Y=0.745 $X2=0 $Y2=0
cc_315 N_A1_N_M1010_g N_VGND_c_707_n 0.00416285f $X=3.835 $Y=0.745 $X2=0 $Y2=0
cc_316 N_A1_N_M1019_g N_VGND_c_707_n 0.00414769f $X=4.265 $Y=0.745 $X2=0 $Y2=0
cc_317 N_A1_N_M1010_g N_VGND_c_711_n 0.00787505f $X=3.835 $Y=0.745 $X2=0 $Y2=0
cc_318 N_A1_N_M1019_g N_VGND_c_711_n 0.00787505f $X=4.265 $Y=0.745 $X2=0 $Y2=0
cc_319 N_A2_N_M1006_g N_VPWR_c_527_n 0.00109252f $X=4.695 $Y=2.465 $X2=0 $Y2=0
cc_320 N_A2_N_M1006_g N_VPWR_c_531_n 0.00357877f $X=4.695 $Y=2.465 $X2=0 $Y2=0
cc_321 N_A2_N_M1014_g N_VPWR_c_531_n 0.00357842f $X=5.125 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A2_N_M1006_g N_VPWR_c_524_n 0.00537654f $X=4.695 $Y=2.465 $X2=0 $Y2=0
cc_323 N_A2_N_M1014_g N_VPWR_c_524_n 0.00640398f $X=5.125 $Y=2.465 $X2=0 $Y2=0
cc_324 N_A2_N_M1006_g N_A_699_367#_c_667_n 0.012237f $X=4.695 $Y=2.465 $X2=0
+ $Y2=0
cc_325 N_A2_N_M1014_g N_A_699_367#_c_667_n 0.010474f $X=5.125 $Y=2.465 $X2=0
+ $Y2=0
cc_326 N_A2_N_M1014_g N_A_699_367#_c_661_n 5.81207e-19 $X=5.125 $Y=2.465 $X2=0
+ $Y2=0
cc_327 N_A2_N_M1006_g N_A_699_367#_c_662_n 6.71626e-19 $X=4.695 $Y=2.465 $X2=0
+ $Y2=0
cc_328 N_A2_N_c_419_n N_A_699_367#_c_662_n 0.00112434f $X=5.05 $Y=1.35 $X2=0
+ $Y2=0
cc_329 N_A2_N_M1014_g N_A_699_367#_c_662_n 0.0125112f $X=5.125 $Y=2.465 $X2=0
+ $Y2=0
cc_330 A2_N N_A_699_367#_c_662_n 0.026915f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_331 N_A2_N_c_417_n N_VGND_c_702_n 0.01013f $X=4.695 $Y=1.275 $X2=0 $Y2=0
cc_332 N_A2_N_c_423_n N_VGND_c_702_n 5.15793e-19 $X=5.237 $Y=1.275 $X2=0 $Y2=0
cc_333 N_A2_N_c_417_n N_VGND_c_704_n 5.59064e-19 $X=4.695 $Y=1.275 $X2=0 $Y2=0
cc_334 N_A2_N_c_419_n N_VGND_c_704_n 0.00134937f $X=5.05 $Y=1.35 $X2=0 $Y2=0
cc_335 A2_N N_VGND_c_704_n 0.0269149f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_336 N_A2_N_c_423_n N_VGND_c_704_n 0.0146435f $X=5.237 $Y=1.275 $X2=0 $Y2=0
cc_337 N_A2_N_c_417_n N_VGND_c_708_n 0.00414769f $X=4.695 $Y=1.275 $X2=0 $Y2=0
cc_338 N_A2_N_c_423_n N_VGND_c_708_n 0.00414769f $X=5.237 $Y=1.275 $X2=0 $Y2=0
cc_339 N_A2_N_c_417_n N_VGND_c_711_n 0.00787505f $X=4.695 $Y=1.275 $X2=0 $Y2=0
cc_340 N_A2_N_c_423_n N_VGND_c_711_n 0.00787505f $X=5.237 $Y=1.275 $X2=0 $Y2=0
cc_341 N_A_30_367#_c_474_n N_VPWR_M1002_s 0.0035201f $X=1.04 $Y=2.375 $X2=-0.19
+ $Y2=1.655
cc_342 N_A_30_367#_c_478_n N_VPWR_M1012_s 0.00780749f $X=2.05 $Y=2.375 $X2=0
+ $Y2=0
cc_343 N_A_30_367#_c_474_n N_VPWR_c_525_n 0.0170777f $X=1.04 $Y=2.375 $X2=0
+ $Y2=0
cc_344 N_A_30_367#_c_478_n N_VPWR_c_526_n 0.0257907f $X=2.05 $Y=2.375 $X2=0
+ $Y2=0
cc_345 N_A_30_367#_c_464_n N_VPWR_c_528_n 0.0178111f $X=0.275 $Y=2.47 $X2=0
+ $Y2=0
cc_346 N_A_30_367#_c_485_n N_VPWR_c_529_n 0.0128073f $X=1.135 $Y=2.455 $X2=0
+ $Y2=0
cc_347 N_A_30_367#_c_489_n N_VPWR_c_530_n 0.0361172f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_348 N_A_30_367#_c_504_p N_VPWR_c_530_n 0.0128782f $X=2.25 $Y=2.99 $X2=0 $Y2=0
cc_349 N_A_30_367#_c_466_n N_VPWR_c_530_n 0.0179183f $X=3.05 $Y=2.905 $X2=0
+ $Y2=0
cc_350 N_A_30_367#_M1002_d N_VPWR_c_524_n 0.00371702f $X=0.15 $Y=1.835 $X2=0
+ $Y2=0
cc_351 N_A_30_367#_M1005_d N_VPWR_c_524_n 0.00501859f $X=0.995 $Y=1.835 $X2=0
+ $Y2=0
cc_352 N_A_30_367#_M1011_d N_VPWR_c_524_n 0.00341839f $X=2.015 $Y=1.835 $X2=0
+ $Y2=0
cc_353 N_A_30_367#_M1016_d N_VPWR_c_524_n 0.00215161f $X=2.875 $Y=1.835 $X2=0
+ $Y2=0
cc_354 N_A_30_367#_c_464_n N_VPWR_c_524_n 0.0100304f $X=0.275 $Y=2.47 $X2=0
+ $Y2=0
cc_355 N_A_30_367#_c_489_n N_VPWR_c_524_n 0.023676f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_356 N_A_30_367#_c_504_p N_VPWR_c_524_n 0.00776497f $X=2.25 $Y=2.99 $X2=0
+ $Y2=0
cc_357 N_A_30_367#_c_466_n N_VPWR_c_524_n 0.0101029f $X=3.05 $Y=2.905 $X2=0
+ $Y2=0
cc_358 N_A_30_367#_c_485_n N_VPWR_c_524_n 0.00769778f $X=1.135 $Y=2.455 $X2=0
+ $Y2=0
cc_359 N_A_30_367#_c_489_n N_Y_M1007_s 0.00332344f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_360 N_A_30_367#_c_465_n N_Y_c_601_n 0.00711126f $X=2.155 $Y=1.99 $X2=0 $Y2=0
cc_361 N_A_30_367#_c_465_n N_Y_c_605_n 0.0177575f $X=2.155 $Y=1.99 $X2=0 $Y2=0
cc_362 N_A_30_367#_c_467_n N_Y_c_605_n 0.034469f $X=3.015 $Y=1.99 $X2=0 $Y2=0
cc_363 N_A_30_367#_c_489_n N_Y_c_628_n 0.0159805f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_364 N_A_30_367#_c_467_n N_A_699_367#_c_659_n 0.0105682f $X=3.015 $Y=1.99
+ $X2=0 $Y2=0
cc_365 N_A_30_367#_c_466_n N_A_699_367#_c_660_n 0.0105682f $X=3.05 $Y=2.905
+ $X2=0 $Y2=0
cc_366 N_A_30_367#_c_467_n N_A_699_367#_c_660_n 0.0396179f $X=3.015 $Y=1.99
+ $X2=0 $Y2=0
cc_367 N_A_30_367#_c_463_n N_VGND_c_700_n 0.00463729f $X=0.275 $Y=1.98 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_524_n N_Y_M1007_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_369 N_VPWR_c_524_n N_A_699_367#_M1001_s 0.00371702f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_370 N_VPWR_c_524_n N_A_699_367#_M1013_s 0.00373407f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_524_n N_A_699_367#_M1014_s 0.00215158f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_372 N_VPWR_c_530_n N_A_699_367#_c_660_n 0.0178111f $X=3.885 $Y=3.33 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_524_n N_A_699_367#_c_660_n 0.0100304f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_374 N_VPWR_M1001_d N_A_699_367#_c_664_n 0.00565274f $X=3.91 $Y=1.835 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_527_n N_A_699_367#_c_664_n 0.0170777f $X=4.05 $Y=2.49 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_531_n N_A_699_367#_c_693_n 0.0139427f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_524_n N_A_699_367#_c_693_n 0.00894187f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_531_n N_A_699_367#_c_667_n 0.0315814f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_524_n N_A_699_367#_c_667_n 0.0197252f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_531_n N_A_699_367#_c_661_n 0.0211538f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_524_n N_A_699_367#_c_661_n 0.0126374f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_382 N_Y_c_601_n N_VGND_M1018_d 0.00267852f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_383 N_Y_c_601_n N_VGND_c_701_n 0.0208822f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_384 N_Y_c_604_n N_VGND_c_701_n 0.0244537f $X=2.585 $Y=0.45 $X2=0 $Y2=0
cc_385 N_Y_c_604_n N_VGND_c_706_n 0.0393378f $X=2.585 $Y=0.45 $X2=0 $Y2=0
cc_386 N_Y_c_604_n N_VGND_c_711_n 0.00977127f $X=2.585 $Y=0.45 $X2=0 $Y2=0
cc_387 N_Y_c_601_n N_A_113_65#_M1008_s 0.00261503f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_388 N_Y_c_602_n N_A_113_65#_c_777_n 0.00538273f $X=1.3 $Y=1.16 $X2=0 $Y2=0
cc_389 N_Y_M1004_d N_A_113_65#_c_778_n 0.00176461f $X=0.995 $Y=0.325 $X2=0 $Y2=0
cc_390 N_Y_c_607_n N_A_113_65#_c_778_n 0.0159398f $X=1.135 $Y=0.7 $X2=0 $Y2=0
cc_391 N_Y_c_601_n N_A_113_65#_c_778_n 0.00280043f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_392 N_Y_c_601_n N_A_113_65#_c_784_n 0.0224504f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_393 N_VGND_c_700_n N_A_113_65#_c_777_n 0.0015231f $X=0.275 $Y=0.47 $X2=0
+ $Y2=0
cc_394 N_VGND_c_701_n N_A_113_65#_c_778_n 0.00962613f $X=2.155 $Y=0.45 $X2=0
+ $Y2=0
cc_395 N_VGND_c_705_n N_A_113_65#_c_778_n 0.0630824f $X=1.99 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_c_711_n N_A_113_65#_c_778_n 0.0370174f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_c_700_n N_A_113_65#_c_779_n 0.00517394f $X=0.275 $Y=0.47 $X2=0
+ $Y2=0
cc_398 N_VGND_c_705_n N_A_113_65#_c_779_n 0.0151705f $X=1.99 $Y=0 $X2=0 $Y2=0
cc_399 N_VGND_c_711_n N_A_113_65#_c_779_n 0.00870596f $X=5.52 $Y=0 $X2=0 $Y2=0
