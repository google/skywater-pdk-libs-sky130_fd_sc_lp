* File: sky130_fd_sc_lp__o211ai_1.pxi.spice
* Created: Wed Sep  2 10:14:29 2020
* 
x_PM_SKY130_FD_SC_LP__O211AI_1%A1 N_A1_M1001_g N_A1_M1007_g A1 A1 N_A1_c_50_n
+ PM_SKY130_FD_SC_LP__O211AI_1%A1
x_PM_SKY130_FD_SC_LP__O211AI_1%A2 N_A2_M1006_g N_A2_M1002_g A2 A2 A2 A2 A2
+ N_A2_c_77_n N_A2_c_78_n N_A2_c_79_n PM_SKY130_FD_SC_LP__O211AI_1%A2
x_PM_SKY130_FD_SC_LP__O211AI_1%B1 N_B1_M1000_g N_B1_M1004_g B1 B1 B1 B1
+ N_B1_c_124_n N_B1_c_127_n B1 PM_SKY130_FD_SC_LP__O211AI_1%B1
x_PM_SKY130_FD_SC_LP__O211AI_1%C1 N_C1_M1005_g N_C1_M1003_g C1 N_C1_c_169_n
+ N_C1_c_170_n PM_SKY130_FD_SC_LP__O211AI_1%C1
x_PM_SKY130_FD_SC_LP__O211AI_1%VPWR N_VPWR_M1007_s N_VPWR_M1000_d N_VPWR_c_199_n
+ N_VPWR_c_200_n N_VPWR_c_201_n VPWR N_VPWR_c_202_n N_VPWR_c_203_n
+ N_VPWR_c_198_n N_VPWR_c_205_n PM_SKY130_FD_SC_LP__O211AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O211AI_1%Y N_Y_M1005_d N_Y_M1006_d N_Y_M1003_d N_Y_c_239_n
+ N_Y_c_243_n N_Y_c_245_n Y Y Y Y Y Y Y N_Y_c_235_n
+ PM_SKY130_FD_SC_LP__O211AI_1%Y
x_PM_SKY130_FD_SC_LP__O211AI_1%A_27_47# N_A_27_47#_M1001_s N_A_27_47#_M1002_d
+ N_A_27_47#_c_278_n N_A_27_47#_c_281_n N_A_27_47#_c_279_n N_A_27_47#_c_293_n
+ PM_SKY130_FD_SC_LP__O211AI_1%A_27_47#
x_PM_SKY130_FD_SC_LP__O211AI_1%VGND N_VGND_M1001_d N_VGND_c_305_n VGND
+ N_VGND_c_306_n N_VGND_c_307_n N_VGND_c_308_n N_VGND_c_309_n
+ PM_SKY130_FD_SC_LP__O211AI_1%VGND
cc_1 VNB N_A1_M1001_g 0.0247879f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A1_M1007_g 0.00692203f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB A1 0.0208507f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_50_n 0.0473626f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.375
cc_5 VNB N_A2_M1006_g 0.00681205f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_6 VNB A2 0.00125489f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_A2_c_77_n 0.0320549f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.295
cc_8 VNB N_A2_c_78_n 0.00653914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A2_c_79_n 0.0185512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_M1004_g 0.024081f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_11 VNB B1 0.00230031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB B1 0.00610792f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_B1_c_124_n 0.0252154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_C1_M1005_g 0.0270421f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_15 VNB N_C1_M1003_g 0.0017608f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_16 VNB N_C1_c_169_n 0.0455283f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.375
cc_17 VNB N_C1_c_170_n 0.00639456f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.375
cc_18 VNB N_VPWR_c_198_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB Y 0.0313003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_235_n 0.050682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_278_n 0.0230847f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_A_27_47#_c_279_n 0.00745492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_305_n 0.0055721f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_24 VNB N_VGND_c_306_n 0.0178675f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_25 VNB N_VGND_c_307_n 0.0524005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_308_n 0.170422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_309_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A1_M1007_g 0.0246048f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_29 VPB A1 0.00695305f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_30 VPB N_A2_M1006_g 0.0197056f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_31 VPB A2 0.00134908f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_32 VPB B1 0.00395756f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_33 VPB N_B1_c_124_n 0.00991804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_B1_c_127_n 0.0182358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_C1_M1003_g 0.0254867f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_36 VPB N_C1_c_170_n 0.00404109f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.375
cc_37 VPB N_VPWR_c_199_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_38 VPB N_VPWR_c_200_n 0.0483776f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_39 VPB N_VPWR_c_201_n 0.0055721f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.375
cc_40 VPB N_VPWR_c_202_n 0.0285189f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.295
cc_41 VPB N_VPWR_c_203_n 0.0285663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_198_n 0.0459344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_205_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB Y 0.0155252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB Y 0.0080869f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.665
cc_46 VPB Y 0.0466859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 N_A1_c_50_n N_A2_M1006_g 0.0608796f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_48 A1 A2 0.0181767f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_49 N_A1_c_50_n A2 0.0068886f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_50 N_A1_M1001_g N_A2_c_77_n 0.0608796f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_51 A1 N_A2_c_77_n 2.55898e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_52 N_A1_M1001_g N_A2_c_78_n 0.0025016f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_53 A1 N_A2_c_78_n 0.0269735f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_A1_M1001_g N_A2_c_79_n 0.0256249f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_55 N_A1_M1007_g N_VPWR_c_200_n 0.0233639f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_56 A1 N_VPWR_c_200_n 0.0270156f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_A1_c_50_n N_VPWR_c_200_n 0.00132775f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_58 N_A1_M1007_g N_VPWR_c_202_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A1_M1007_g N_VPWR_c_198_n 0.00818711f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_60 N_A1_M1001_g N_A_27_47#_c_278_n 0.0111213f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_61 N_A1_M1001_g N_A_27_47#_c_281_n 0.0127239f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_62 A1 N_A_27_47#_c_281_n 6.40987e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A1_M1001_g N_A_27_47#_c_279_n 7.3104e-19 $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_64 A1 N_A_27_47#_c_279_n 0.0271908f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A1_c_50_n N_A_27_47#_c_279_n 0.00201405f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_66 N_A1_M1001_g N_VGND_c_305_n 0.00563167f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_67 N_A1_M1001_g N_VGND_c_306_n 0.0054895f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_68 N_A1_M1001_g N_VGND_c_308_n 0.00735185f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_69 N_A2_c_78_n N_B1_M1004_g 5.90752e-19 $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_70 N_A2_c_79_n N_B1_M1004_g 0.0232272f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_71 N_A2_c_78_n B1 0.00513415f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_72 N_A2_c_79_n B1 0.00107993f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_73 N_A2_M1006_g B1 9.75472e-19 $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_74 A2 B1 0.0089903f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_75 N_A2_c_77_n B1 2.12376e-19 $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_76 N_A2_c_78_n B1 0.0114245f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_77 N_A2_M1006_g N_B1_c_124_n 0.0294577f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_78 A2 N_B1_c_124_n 0.00177376f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_79 N_A2_c_77_n N_B1_c_124_n 0.0107049f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_80 N_A2_c_78_n N_B1_c_124_n 5.88442e-19 $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_81 N_A2_M1006_g N_VPWR_c_200_n 0.00259911f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A2_M1006_g N_VPWR_c_202_n 0.00480784f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_83 A2 N_VPWR_c_202_n 0.00597736f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A2_M1006_g N_VPWR_c_198_n 0.00812063f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_85 A2 N_VPWR_c_198_n 0.00770133f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_86 A2 A_110_367# 0.00139886f $X=0.635 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_87 N_A2_M1006_g N_Y_c_239_n 0.0014537f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_88 A2 N_Y_c_239_n 0.0137332f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A2_c_77_n N_Y_c_239_n 0.00169907f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A2_c_78_n N_Y_c_239_n 0.00299772f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_91 N_A2_M1006_g N_Y_c_243_n 0.00862145f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_92 A2 N_Y_c_243_n 0.0551246f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_93 N_A2_c_79_n N_A_27_47#_c_278_n 7.0638e-19 $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_94 N_A2_c_77_n N_A_27_47#_c_281_n 0.00450164f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_95 N_A2_c_78_n N_A_27_47#_c_281_n 0.0339425f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_96 N_A2_c_79_n N_A_27_47#_c_281_n 0.0127398f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_97 N_A2_c_79_n N_VGND_c_305_n 0.00403719f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_98 N_A2_c_79_n N_VGND_c_307_n 0.00585385f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_99 N_A2_c_79_n N_VGND_c_308_n 0.00689251f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_100 N_B1_M1004_g N_C1_M1005_g 0.0486209f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_101 B1 N_C1_M1005_g 0.00466307f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_102 N_B1_c_127_n N_C1_M1003_g 0.0228447f $X=1.465 $Y=1.725 $X2=0 $Y2=0
cc_103 B1 N_C1_c_169_n 0.00466307f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B1_c_124_n N_C1_c_169_n 0.0486209f $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B1_M1004_g N_C1_c_170_n 3.26672e-19 $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_106 B1 N_C1_c_170_n 0.0393682f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_107 N_B1_c_127_n N_VPWR_c_201_n 0.00422051f $X=1.465 $Y=1.725 $X2=0 $Y2=0
cc_108 N_B1_c_127_n N_VPWR_c_202_n 0.00585385f $X=1.465 $Y=1.725 $X2=0 $Y2=0
cc_109 N_B1_c_127_n N_VPWR_c_198_n 0.0111121f $X=1.465 $Y=1.725 $X2=0 $Y2=0
cc_110 B1 N_Y_c_245_n 0.0366899f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B1_c_124_n N_Y_c_245_n 9.67719e-19 $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_112 N_B1_c_127_n N_Y_c_245_n 0.0135074f $X=1.465 $Y=1.725 $X2=0 $Y2=0
cc_113 B1 Y 0.00455092f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_114 N_B1_c_127_n Y 6.9385e-19 $X=1.465 $Y=1.725 $X2=0 $Y2=0
cc_115 N_B1_M1004_g N_Y_c_235_n 9.23438e-19 $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_116 B1 N_Y_c_235_n 0.0303031f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_117 B1 N_A_27_47#_c_281_n 0.013673f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_118 B1 N_A_27_47#_c_281_n 0.00501954f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_119 N_B1_c_124_n N_A_27_47#_c_281_n 7.14813e-19 $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_120 N_B1_M1004_g N_A_27_47#_c_293_n 0.00266525f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_121 B1 N_A_27_47#_c_293_n 0.0338166f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_122 N_B1_M1004_g N_VGND_c_307_n 0.00506294f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_123 B1 N_VGND_c_307_n 0.00703416f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_124 N_B1_M1004_g N_VGND_c_308_n 0.00882722f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_125 B1 N_VGND_c_308_n 0.00774524f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_126 B1 A_326_47# 0.00122477f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_127 N_C1_M1003_g N_VPWR_c_201_n 0.00422051f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_128 N_C1_M1003_g N_VPWR_c_203_n 0.00571722f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_129 N_C1_M1003_g N_VPWR_c_198_n 0.0118478f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_130 N_C1_M1003_g N_Y_c_245_n 0.0166238f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_131 N_C1_c_170_n N_Y_c_245_n 0.00100284f $X=2.1 $Y=1.46 $X2=0 $Y2=0
cc_132 N_C1_M1005_g Y 0.00254121f $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_133 N_C1_M1003_g Y 0.00304773f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_134 N_C1_c_169_n Y 0.00220283f $X=2.1 $Y=1.46 $X2=0 $Y2=0
cc_135 N_C1_c_170_n Y 0.040237f $X=2.1 $Y=1.46 $X2=0 $Y2=0
cc_136 N_C1_M1003_g Y 2.7414e-19 $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_137 N_C1_c_169_n Y 0.00137401f $X=2.1 $Y=1.46 $X2=0 $Y2=0
cc_138 N_C1_c_170_n Y 0.0259024f $X=2.1 $Y=1.46 $X2=0 $Y2=0
cc_139 N_C1_M1003_g Y 0.0130693f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_140 N_C1_M1005_g N_Y_c_235_n 0.0143157f $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_141 N_C1_c_169_n N_Y_c_235_n 0.00213231f $X=2.1 $Y=1.46 $X2=0 $Y2=0
cc_142 N_C1_c_170_n N_Y_c_235_n 0.0256707f $X=2.1 $Y=1.46 $X2=0 $Y2=0
cc_143 N_C1_M1005_g N_VGND_c_307_n 0.0054895f $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_144 N_C1_M1005_g N_VGND_c_308_n 0.0111524f $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_145 N_VPWR_c_198_n A_110_367# 0.00385363f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_146 N_VPWR_c_198_n N_Y_M1006_d 0.00752153f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_147 N_VPWR_c_198_n N_Y_M1003_d 0.00500006f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_148 N_VPWR_c_200_n N_Y_c_243_n 0.00615351f $X=0.26 $Y=2.005 $X2=0 $Y2=0
cc_149 N_VPWR_c_202_n N_Y_c_243_n 0.0172383f $X=1.48 $Y=3.33 $X2=0 $Y2=0
cc_150 N_VPWR_c_198_n N_Y_c_243_n 0.0102248f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_151 N_VPWR_M1000_d N_Y_c_245_n 0.00588714f $X=1.45 $Y=1.835 $X2=0 $Y2=0
cc_152 N_VPWR_c_201_n N_Y_c_245_n 0.022455f $X=1.645 $Y=2.39 $X2=0 $Y2=0
cc_153 N_VPWR_c_203_n Y 0.0543249f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_154 N_VPWR_c_198_n Y 0.03091f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_155 N_Y_c_235_n N_A_27_47#_c_293_n 0.00424342f $X=2.47 $Y=0.38 $X2=0 $Y2=0
cc_156 N_Y_c_235_n N_VGND_c_307_n 0.0553475f $X=2.47 $Y=0.38 $X2=0 $Y2=0
cc_157 N_Y_M1005_d N_VGND_c_308_n 0.00500006f $X=1.99 $Y=0.235 $X2=0 $Y2=0
cc_158 N_Y_c_235_n N_VGND_c_308_n 0.0314246f $X=2.47 $Y=0.38 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_281_n N_VGND_M1001_d 0.0058207f $X=1.125 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_27_47#_c_281_n N_VGND_c_305_n 0.0219723f $X=1.125 $Y=0.93 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_278_n N_VGND_c_306_n 0.0210467f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_293_n N_VGND_c_307_n 0.0184639f $X=1.29 $Y=0.42 $X2=0 $Y2=0
cc_163 N_A_27_47#_M1001_s N_VGND_c_308_n 0.00215158f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_M1002_d N_VGND_c_308_n 0.00614803f $X=1.09 $Y=0.235 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_278_n N_VGND_c_308_n 0.0125689f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_281_n N_VGND_c_308_n 0.0117712f $X=1.125 $Y=0.93 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_293_n N_VGND_c_308_n 0.0106136f $X=1.29 $Y=0.42 $X2=0 $Y2=0
cc_168 N_VGND_c_308_n A_326_47# 0.00339089f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
