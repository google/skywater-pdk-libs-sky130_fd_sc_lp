* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_89_367# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_89_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR A2 a_89_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_63_65# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_867_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND B2 a_63_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR A1 a_89_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 Y B1 a_89_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_63_65# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VGND B2 a_63_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_63_65# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 Y A1 a_867_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_867_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_89_367# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VGND A2 a_867_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_89_367# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 Y B2 a_89_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 Y A1 a_867_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 Y B1 a_63_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_63_65# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_89_367# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 Y B1 a_89_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 Y B1 a_63_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_867_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_867_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 VPWR A2 a_89_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 VGND A2 a_867_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 VPWR A1 a_89_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 a_89_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_89_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_89_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 Y B2 a_89_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
