* File: sky130_fd_sc_lp__o311a_0.pxi.spice
* Created: Wed Sep  2 10:22:46 2020
* 
x_PM_SKY130_FD_SC_LP__O311A_0%A_96_161# N_A_96_161#_M1010_d N_A_96_161#_M1007_d
+ N_A_96_161#_M1001_d N_A_96_161#_c_92_n N_A_96_161#_c_93_n N_A_96_161#_M1000_g
+ N_A_96_161#_c_94_n N_A_96_161#_M1002_g N_A_96_161#_c_95_n N_A_96_161#_c_101_n
+ N_A_96_161#_c_102_n N_A_96_161#_c_96_n N_A_96_161#_c_97_n N_A_96_161#_c_105_n
+ N_A_96_161#_c_106_n N_A_96_161#_c_107_n N_A_96_161#_c_108_n N_A_96_161#_c_98_n
+ N_A_96_161#_c_110_n N_A_96_161#_c_111_n N_A_96_161#_c_99_n N_A_96_161#_c_112_n
+ PM_SKY130_FD_SC_LP__O311A_0%A_96_161#
x_PM_SKY130_FD_SC_LP__O311A_0%A1 N_A1_M1003_g N_A1_c_198_n N_A1_M1011_g
+ N_A1_c_199_n N_A1_c_200_n N_A1_c_207_n N_A1_c_201_n A1 A1 A1 N_A1_c_203_n
+ N_A1_c_204_n PM_SKY130_FD_SC_LP__O311A_0%A1
x_PM_SKY130_FD_SC_LP__O311A_0%A2 N_A2_c_259_n N_A2_M1006_g N_A2_M1005_g
+ N_A2_c_256_n A2 A2 N_A2_c_258_n PM_SKY130_FD_SC_LP__O311A_0%A2
x_PM_SKY130_FD_SC_LP__O311A_0%A3 N_A3_M1007_g N_A3_M1004_g N_A3_c_302_n
+ N_A3_c_303_n A3 A3 N_A3_c_304_n N_A3_c_305_n PM_SKY130_FD_SC_LP__O311A_0%A3
x_PM_SKY130_FD_SC_LP__O311A_0%B1 N_B1_M1009_g N_B1_M1008_g N_B1_c_346_n B1 B1
+ N_B1_c_348_n PM_SKY130_FD_SC_LP__O311A_0%B1
x_PM_SKY130_FD_SC_LP__O311A_0%C1 N_C1_c_391_n N_C1_M1010_g N_C1_M1001_g
+ N_C1_c_392_n N_C1_c_393_n N_C1_c_399_n N_C1_c_400_n N_C1_c_394_n N_C1_c_395_n
+ C1 C1 C1 N_C1_c_397_n PM_SKY130_FD_SC_LP__O311A_0%C1
x_PM_SKY130_FD_SC_LP__O311A_0%X N_X_M1002_s N_X_M1000_s N_X_c_439_n X X X X X X
+ X N_X_c_436_n X PM_SKY130_FD_SC_LP__O311A_0%X
x_PM_SKY130_FD_SC_LP__O311A_0%VPWR N_VPWR_M1000_d N_VPWR_M1009_d N_VPWR_c_458_n
+ N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n N_VPWR_c_463_n
+ VPWR N_VPWR_c_464_n N_VPWR_c_457_n PM_SKY130_FD_SC_LP__O311A_0%VPWR
x_PM_SKY130_FD_SC_LP__O311A_0%VGND N_VGND_M1002_d N_VGND_M1005_d N_VGND_c_495_n
+ N_VGND_c_496_n VGND N_VGND_c_497_n N_VGND_c_498_n N_VGND_c_499_n
+ N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n PM_SKY130_FD_SC_LP__O311A_0%VGND
x_PM_SKY130_FD_SC_LP__O311A_0%A_292_55# N_A_292_55#_M1011_d N_A_292_55#_M1004_d
+ N_A_292_55#_c_542_n N_A_292_55#_c_543_n N_A_292_55#_c_544_n
+ N_A_292_55#_c_546_n PM_SKY130_FD_SC_LP__O311A_0%A_292_55#
cc_1 VNB N_A_96_161#_c_92_n 0.0270634f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.88
cc_2 VNB N_A_96_161#_c_93_n 0.00994638f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.88
cc_3 VNB N_A_96_161#_c_94_n 0.0206899f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.805
cc_4 VNB N_A_96_161#_c_95_n 0.0366948f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.545
cc_5 VNB N_A_96_161#_c_96_n 0.0043422f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.71
cc_6 VNB N_A_96_161#_c_97_n 0.0115152f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.71
cc_7 VNB N_A_96_161#_c_98_n 0.0170045f $X=-0.19 $Y=-0.245 $X2=3.197 $Y2=2.045
cc_8 VNB N_A_96_161#_c_99_n 0.0136503f $X=-0.19 $Y=-0.245 $X2=3.32 $Y2=0.485
cc_9 VNB N_A1_c_198_n 0.0169204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_199_n 0.0132826f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.545
cc_11 VNB N_A1_c_200_n 0.019452f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.88
cc_12 VNB N_A1_c_201_n 0.0174054f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.725
cc_13 VNB A1 0.003449f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.485
cc_14 VNB N_A1_c_203_n 0.0165202f $X=-0.19 $Y=-0.245 $X2=0.702 $Y2=2.045
cc_15 VNB N_A1_c_204_n 0.00720152f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.71
cc_16 VNB N_A2_M1005_g 0.0376256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_256_n 0.0181551f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.545
cc_18 VNB A2 0.00519626f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.88
cc_19 VNB N_A2_c_258_n 0.0153265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A3_M1004_g 0.0309607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A3_c_302_n 0.0212748f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.545
cc_22 VNB N_A3_c_303_n 0.00440602f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.88
cc_23 VNB N_A3_c_304_n 0.0154282f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.805
cc_24 VNB N_A3_c_305_n 0.0059353f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.485
cc_25 VNB N_B1_M1008_g 0.0363403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B1_c_346_n 0.0205972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB B1 0.00929886f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.88
cc_28 VNB N_B1_c_348_n 0.0188296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_C1_c_391_n 0.0201336f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=0.275
cc_30 VNB N_C1_c_392_n 0.0400352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C1_c_393_n 0.0108563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_C1_c_394_n 0.00971496f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.88
cc_33 VNB N_C1_c_395_n 0.0195023f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.725
cc_34 VNB C1 0.03088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C1_c_397_n 0.0323749f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.215
cc_36 VNB X 0.0566872f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.88
cc_37 VNB N_X_c_436_n 0.0164934f $X=-0.19 $Y=-0.245 $X2=0.702 $Y2=1.71
cc_38 VNB N_VPWR_c_457_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_495_n 0.00125039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_496_n 0.00364944f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.88
cc_41 VNB N_VGND_c_497_n 0.026705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_498_n 0.0136923f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.545
cc_43 VNB N_VGND_c_499_n 0.0478807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_500_n 0.234109f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=2.13
cc_45 VNB N_VGND_c_501_n 0.0048828f $X=-0.19 $Y=-0.245 $X2=2.405 $Y2=2.55
cc_46 VNB N_VGND_c_502_n 0.00541044f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=2.13
cc_47 VNB N_A_292_55#_c_542_n 8.37384e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_292_55#_c_543_n 0.0158542f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.545
cc_49 VNB N_A_292_55#_c_544_n 0.00408748f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.88
cc_50 VPB N_A_96_161#_M1000_g 0.0261503f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.725
cc_51 VPB N_A_96_161#_c_101_n 0.0243921f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.05
cc_52 VPB N_A_96_161#_c_102_n 0.017452f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.215
cc_53 VPB N_A_96_161#_c_96_n 0.0034089f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.71
cc_54 VPB N_A_96_161#_c_97_n 0.00377125f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.71
cc_55 VPB N_A_96_161#_c_105_n 0.0442846f $X=-0.19 $Y=1.655 $X2=2.24 $Y2=2.13
cc_56 VPB N_A_96_161#_c_106_n 0.00240336f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.13
cc_57 VPB N_A_96_161#_c_107_n 0.0022968f $X=-0.19 $Y=1.655 $X2=2.405 $Y2=2.55
cc_58 VPB N_A_96_161#_c_108_n 0.0084939f $X=-0.19 $Y=1.655 $X2=3.09 $Y2=2.13
cc_59 VPB N_A_96_161#_c_98_n 0.00865455f $X=-0.19 $Y=1.655 $X2=3.197 $Y2=2.045
cc_60 VPB N_A_96_161#_c_110_n 0.0339812f $X=-0.19 $Y=1.655 $X2=3.35 $Y2=2.55
cc_61 VPB N_A_96_161#_c_111_n 0.00579008f $X=-0.19 $Y=1.655 $X2=2.405 $Y2=2.13
cc_62 VPB N_A_96_161#_c_112_n 0.00407275f $X=-0.19 $Y=1.655 $X2=3.302 $Y2=2.13
cc_63 VPB N_A1_M1003_g 0.0415206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A1_c_200_n 0.00271795f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=0.88
cc_65 VPB N_A1_c_207_n 0.0153157f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.88
cc_66 VPB A1 0.00304703f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.485
cc_67 VPB N_A2_c_259_n 0.0152409f $X=-0.19 $Y=1.655 $X2=3.18 $Y2=0.275
cc_68 VPB N_A2_M1006_g 0.0394795f $X=-0.19 $Y=1.655 $X2=3.21 $Y2=2.405
cc_69 VPB N_A2_c_256_n 0.00271709f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.545
cc_70 VPB A2 0.00288963f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=0.88
cc_71 VPB N_A3_M1007_g 0.0444266f $X=-0.19 $Y=1.655 $X2=3.21 $Y2=2.405
cc_72 VPB N_A3_c_303_n 0.0111009f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=0.88
cc_73 VPB N_A3_c_305_n 0.0034354f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.485
cc_74 VPB N_B1_M1009_g 0.024821f $X=-0.19 $Y=1.655 $X2=3.21 $Y2=2.405
cc_75 VPB N_B1_c_346_n 0.0449815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB B1 0.00342416f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=0.88
cc_77 VPB N_C1_M1001_g 0.0222366f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_C1_c_399_n 0.0304247f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.955
cc_79 VPB N_C1_c_400_n 0.00912178f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.545
cc_80 VPB N_C1_c_394_n 0.034149f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.88
cc_81 VPB C1 0.015712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB X 0.0396636f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=0.88
cc_83 VPB X 0.0448256f $X=-0.19 $Y=1.655 $X2=3.377 $Y2=2.215
cc_84 VPB N_VPWR_c_458_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_459_n 0.00675677f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.88
cc_86 VPB N_VPWR_c_460_n 0.0234952f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.725
cc_87 VPB N_VPWR_c_461_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_462_n 0.0468709f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.485
cc_89 VPB N_VPWR_c_463_n 0.00554856f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.485
cc_90 VPB N_VPWR_c_464_n 0.02341f $X=-0.19 $Y=1.655 $X2=2.405 $Y2=2.55
cc_91 VPB N_VPWR_c_457_n 0.0909202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 N_A_96_161#_c_101_n N_A1_M1003_g 0.0204786f $X=0.645 $Y=2.05 $X2=0 $Y2=0
cc_93 N_A_96_161#_c_96_n N_A1_M1003_g 0.00352602f $X=0.645 $Y=1.71 $X2=0 $Y2=0
cc_94 N_A_96_161#_c_105_n N_A1_M1003_g 0.015718f $X=2.24 $Y=2.13 $X2=0 $Y2=0
cc_95 N_A_96_161#_c_94_n N_A1_c_198_n 0.0104989f $X=0.915 $Y=0.805 $X2=0 $Y2=0
cc_96 N_A_96_161#_c_95_n N_A1_c_199_n 0.00349479f $X=0.645 $Y=1.545 $X2=0 $Y2=0
cc_97 N_A_96_161#_c_96_n N_A1_c_200_n 0.00180329f $X=0.645 $Y=1.71 $X2=0 $Y2=0
cc_98 N_A_96_161#_c_97_n N_A1_c_200_n 0.00996349f $X=0.645 $Y=1.71 $X2=0 $Y2=0
cc_99 N_A_96_161#_c_101_n N_A1_c_207_n 0.00996349f $X=0.645 $Y=2.05 $X2=0 $Y2=0
cc_100 N_A_96_161#_c_105_n N_A1_c_207_n 0.00144107f $X=2.24 $Y=2.13 $X2=0 $Y2=0
cc_101 N_A_96_161#_c_92_n N_A1_c_201_n 0.0098294f $X=0.84 $Y=0.88 $X2=0 $Y2=0
cc_102 N_A_96_161#_c_95_n A1 0.00162431f $X=0.645 $Y=1.545 $X2=0 $Y2=0
cc_103 N_A_96_161#_c_96_n A1 0.0251567f $X=0.645 $Y=1.71 $X2=0 $Y2=0
cc_104 N_A_96_161#_c_97_n A1 3.61015e-19 $X=0.645 $Y=1.71 $X2=0 $Y2=0
cc_105 N_A_96_161#_c_105_n A1 0.024955f $X=2.24 $Y=2.13 $X2=0 $Y2=0
cc_106 N_A_96_161#_c_95_n N_A1_c_203_n 0.0101706f $X=0.645 $Y=1.545 $X2=0 $Y2=0
cc_107 N_A_96_161#_c_92_n N_A1_c_204_n 0.00169658f $X=0.84 $Y=0.88 $X2=0 $Y2=0
cc_108 N_A_96_161#_c_95_n N_A1_c_204_n 0.00201796f $X=0.645 $Y=1.545 $X2=0 $Y2=0
cc_109 N_A_96_161#_c_105_n N_A2_c_259_n 0.00263933f $X=2.24 $Y=2.13 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_96_161#_c_105_n N_A2_M1006_g 0.0152669f $X=2.24 $Y=2.13 $X2=0 $Y2=0
cc_111 N_A_96_161#_c_107_n N_A2_M1006_g 0.00399634f $X=2.405 $Y=2.55 $X2=0 $Y2=0
cc_112 N_A_96_161#_c_105_n A2 0.02387f $X=2.24 $Y=2.13 $X2=0 $Y2=0
cc_113 N_A_96_161#_c_105_n N_A3_M1007_g 0.0125426f $X=2.24 $Y=2.13 $X2=0 $Y2=0
cc_114 N_A_96_161#_c_107_n N_A3_M1007_g 0.0175276f $X=2.405 $Y=2.55 $X2=0 $Y2=0
cc_115 N_A_96_161#_c_111_n N_A3_M1007_g 0.00247816f $X=2.405 $Y=2.13 $X2=0 $Y2=0
cc_116 N_A_96_161#_c_111_n N_A3_c_303_n 0.00403626f $X=2.405 $Y=2.13 $X2=0 $Y2=0
cc_117 N_A_96_161#_c_105_n N_A3_c_305_n 0.0147182f $X=2.24 $Y=2.13 $X2=0 $Y2=0
cc_118 N_A_96_161#_c_111_n N_A3_c_305_n 0.00869822f $X=2.405 $Y=2.13 $X2=0 $Y2=0
cc_119 N_A_96_161#_c_107_n N_B1_M1009_g 0.0122634f $X=2.405 $Y=2.55 $X2=0 $Y2=0
cc_120 N_A_96_161#_c_108_n N_B1_M1009_g 0.00811981f $X=3.09 $Y=2.13 $X2=0 $Y2=0
cc_121 N_A_96_161#_c_111_n N_B1_M1009_g 0.00100835f $X=2.405 $Y=2.13 $X2=0 $Y2=0
cc_122 N_A_96_161#_c_98_n N_B1_M1008_g 0.0056631f $X=3.197 $Y=2.045 $X2=0 $Y2=0
cc_123 N_A_96_161#_c_99_n N_B1_M1008_g 9.91949e-19 $X=3.32 $Y=0.485 $X2=0 $Y2=0
cc_124 N_A_96_161#_c_108_n N_B1_c_346_n 0.0124789f $X=3.09 $Y=2.13 $X2=0 $Y2=0
cc_125 N_A_96_161#_c_98_n N_B1_c_346_n 0.00425691f $X=3.197 $Y=2.045 $X2=0 $Y2=0
cc_126 N_A_96_161#_c_111_n N_B1_c_346_n 0.00137218f $X=2.405 $Y=2.13 $X2=0 $Y2=0
cc_127 N_A_96_161#_c_108_n B1 0.0261827f $X=3.09 $Y=2.13 $X2=0 $Y2=0
cc_128 N_A_96_161#_c_98_n B1 0.0584892f $X=3.197 $Y=2.045 $X2=0 $Y2=0
cc_129 N_A_96_161#_c_111_n B1 0.00436171f $X=2.405 $Y=2.13 $X2=0 $Y2=0
cc_130 N_A_96_161#_c_98_n N_B1_c_348_n 0.00613237f $X=3.197 $Y=2.045 $X2=0 $Y2=0
cc_131 N_A_96_161#_c_98_n N_C1_c_391_n 0.0055724f $X=3.197 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A_96_161#_c_99_n N_C1_c_391_n 0.00750098f $X=3.32 $Y=0.485 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_96_161#_c_110_n N_C1_M1001_g 0.00486636f $X=3.35 $Y=2.55 $X2=0 $Y2=0
cc_134 N_A_96_161#_c_98_n N_C1_c_392_n 0.00935096f $X=3.197 $Y=2.045 $X2=0 $Y2=0
cc_135 N_A_96_161#_c_99_n N_C1_c_392_n 0.00788201f $X=3.32 $Y=0.485 $X2=0 $Y2=0
cc_136 N_A_96_161#_c_98_n N_C1_c_393_n 0.005224f $X=3.197 $Y=2.045 $X2=0 $Y2=0
cc_137 N_A_96_161#_c_110_n N_C1_c_399_n 0.00994145f $X=3.35 $Y=2.55 $X2=0 $Y2=0
cc_138 N_A_96_161#_c_112_n N_C1_c_399_n 0.0129722f $X=3.302 $Y=2.13 $X2=0 $Y2=0
cc_139 N_A_96_161#_c_107_n N_C1_c_400_n 5.7515e-19 $X=2.405 $Y=2.55 $X2=0 $Y2=0
cc_140 N_A_96_161#_c_108_n N_C1_c_400_n 0.00316416f $X=3.09 $Y=2.13 $X2=0 $Y2=0
cc_141 N_A_96_161#_c_112_n N_C1_c_400_n 0.0104893f $X=3.302 $Y=2.13 $X2=0 $Y2=0
cc_142 N_A_96_161#_c_112_n N_C1_c_394_n 0.00745704f $X=3.302 $Y=2.13 $X2=0 $Y2=0
cc_143 N_A_96_161#_c_98_n C1 0.0779791f $X=3.197 $Y=2.045 $X2=0 $Y2=0
cc_144 N_A_96_161#_c_99_n C1 7.35155e-19 $X=3.32 $Y=0.485 $X2=0 $Y2=0
cc_145 N_A_96_161#_c_112_n C1 0.00308258f $X=3.302 $Y=2.13 $X2=0 $Y2=0
cc_146 N_A_96_161#_c_98_n N_C1_c_397_n 0.0114326f $X=3.197 $Y=2.045 $X2=0 $Y2=0
cc_147 N_A_96_161#_c_93_n N_X_c_439_n 0.0129787f $X=0.63 $Y=0.88 $X2=0 $Y2=0
cc_148 N_A_96_161#_c_93_n X 0.0378791f $X=0.63 $Y=0.88 $X2=0 $Y2=0
cc_149 N_A_96_161#_M1000_g X 0.00549575f $X=0.735 $Y=2.725 $X2=0 $Y2=0
cc_150 N_A_96_161#_c_94_n X 0.00377806f $X=0.915 $Y=0.805 $X2=0 $Y2=0
cc_151 N_A_96_161#_c_96_n X 0.0389168f $X=0.645 $Y=1.71 $X2=0 $Y2=0
cc_152 N_A_96_161#_c_106_n X 0.0141027f $X=0.855 $Y=2.13 $X2=0 $Y2=0
cc_153 N_A_96_161#_M1000_g X 0.0073672f $X=0.735 $Y=2.725 $X2=0 $Y2=0
cc_154 N_A_96_161#_c_102_n X 0.00422121f $X=0.645 $Y=2.215 $X2=0 $Y2=0
cc_155 N_A_96_161#_c_106_n X 0.0105576f $X=0.855 $Y=2.13 $X2=0 $Y2=0
cc_156 N_A_96_161#_M1000_g N_VPWR_c_458_n 0.00312359f $X=0.735 $Y=2.725 $X2=0
+ $Y2=0
cc_157 N_A_96_161#_c_105_n N_VPWR_c_458_n 0.0264827f $X=2.24 $Y=2.13 $X2=0 $Y2=0
cc_158 N_A_96_161#_c_106_n N_VPWR_c_458_n 0.00126356f $X=0.855 $Y=2.13 $X2=0
+ $Y2=0
cc_159 N_A_96_161#_c_107_n N_VPWR_c_459_n 0.0263049f $X=2.405 $Y=2.55 $X2=0
+ $Y2=0
cc_160 N_A_96_161#_c_108_n N_VPWR_c_459_n 0.0265262f $X=3.09 $Y=2.13 $X2=0 $Y2=0
cc_161 N_A_96_161#_c_110_n N_VPWR_c_459_n 0.0262732f $X=3.35 $Y=2.55 $X2=0 $Y2=0
cc_162 N_A_96_161#_M1000_g N_VPWR_c_460_n 0.00523511f $X=0.735 $Y=2.725 $X2=0
+ $Y2=0
cc_163 N_A_96_161#_c_107_n N_VPWR_c_462_n 0.0220529f $X=2.405 $Y=2.55 $X2=0
+ $Y2=0
cc_164 N_A_96_161#_c_110_n N_VPWR_c_464_n 0.0184069f $X=3.35 $Y=2.55 $X2=0 $Y2=0
cc_165 N_A_96_161#_M1000_g N_VPWR_c_457_n 0.0108546f $X=0.735 $Y=2.725 $X2=0
+ $Y2=0
cc_166 N_A_96_161#_c_107_n N_VPWR_c_457_n 0.0126084f $X=2.405 $Y=2.55 $X2=0
+ $Y2=0
cc_167 N_A_96_161#_c_110_n N_VPWR_c_457_n 0.0105632f $X=3.35 $Y=2.55 $X2=0 $Y2=0
cc_168 N_A_96_161#_c_94_n N_VGND_c_495_n 0.0101345f $X=0.915 $Y=0.805 $X2=0
+ $Y2=0
cc_169 N_A_96_161#_c_94_n N_VGND_c_497_n 0.00525707f $X=0.915 $Y=0.805 $X2=0
+ $Y2=0
cc_170 N_A_96_161#_c_99_n N_VGND_c_499_n 0.0171532f $X=3.32 $Y=0.485 $X2=0 $Y2=0
cc_171 N_A_96_161#_c_92_n N_VGND_c_500_n 6.15481e-19 $X=0.84 $Y=0.88 $X2=0 $Y2=0
cc_172 N_A_96_161#_c_94_n N_VGND_c_500_n 0.010392f $X=0.915 $Y=0.805 $X2=0 $Y2=0
cc_173 N_A_96_161#_c_99_n N_VGND_c_500_n 0.0140776f $X=3.32 $Y=0.485 $X2=0 $Y2=0
cc_174 N_A_96_161#_c_98_n N_A_292_55#_c_543_n 0.00663892f $X=3.197 $Y=2.045
+ $X2=0 $Y2=0
cc_175 N_A_96_161#_c_98_n N_A_292_55#_c_546_n 0.00329679f $X=3.197 $Y=2.045
+ $X2=0 $Y2=0
cc_176 N_A_96_161#_c_99_n N_A_292_55#_c_546_n 0.0126869f $X=3.32 $Y=0.485 $X2=0
+ $Y2=0
cc_177 N_A1_c_207_n N_A2_c_259_n 0.014448f $X=1.185 $Y=1.865 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A1_M1003_g N_A2_M1006_g 0.0579734f $X=1.275 $Y=2.725 $X2=0 $Y2=0
cc_179 N_A1_c_198_n N_A2_M1005_g 0.0180403f $X=1.385 $Y=0.805 $X2=0 $Y2=0
cc_180 N_A1_c_199_n N_A2_M1005_g 0.00663444f $X=1.185 $Y=1.195 $X2=0 $Y2=0
cc_181 A1 N_A2_M1005_g 2.35678e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A1_c_204_n N_A2_M1005_g 0.00282942f $X=1.192 $Y=1.167 $X2=0 $Y2=0
cc_183 N_A1_c_200_n N_A2_c_256_n 0.014448f $X=1.185 $Y=1.7 $X2=0 $Y2=0
cc_184 A1 A2 0.0557038f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A1_c_203_n A2 0.00214114f $X=1.185 $Y=1.36 $X2=0 $Y2=0
cc_186 A1 N_A2_c_258_n 0.00205669f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_187 N_A1_c_203_n N_A2_c_258_n 0.014448f $X=1.185 $Y=1.36 $X2=0 $Y2=0
cc_188 A1 N_A3_c_305_n 8.78701e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A1_c_204_n N_A3_c_305_n 0.00278474f $X=1.192 $Y=1.167 $X2=0 $Y2=0
cc_190 A1 X 0.0107558f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_191 N_A1_c_204_n X 0.0105032f $X=1.192 $Y=1.167 $X2=0 $Y2=0
cc_192 N_A1_M1003_g N_VPWR_c_458_n 0.00388829f $X=1.275 $Y=2.725 $X2=0 $Y2=0
cc_193 N_A1_M1003_g N_VPWR_c_462_n 0.0053602f $X=1.275 $Y=2.725 $X2=0 $Y2=0
cc_194 N_A1_M1003_g N_VPWR_c_457_n 0.010475f $X=1.275 $Y=2.725 $X2=0 $Y2=0
cc_195 N_A1_c_198_n N_VGND_c_495_n 0.00734999f $X=1.385 $Y=0.805 $X2=0 $Y2=0
cc_196 N_A1_c_201_n N_VGND_c_495_n 0.00288829f $X=1.385 $Y=0.88 $X2=0 $Y2=0
cc_197 N_A1_c_203_n N_VGND_c_495_n 6.20658e-19 $X=1.185 $Y=1.36 $X2=0 $Y2=0
cc_198 N_A1_c_204_n N_VGND_c_495_n 0.0198472f $X=1.192 $Y=1.167 $X2=0 $Y2=0
cc_199 N_A1_c_198_n N_VGND_c_496_n 5.60389e-19 $X=1.385 $Y=0.805 $X2=0 $Y2=0
cc_200 N_A1_c_198_n N_VGND_c_498_n 0.00525707f $X=1.385 $Y=0.805 $X2=0 $Y2=0
cc_201 N_A1_c_198_n N_VGND_c_500_n 0.00878876f $X=1.385 $Y=0.805 $X2=0 $Y2=0
cc_202 N_A1_c_204_n N_VGND_c_500_n 0.00173248f $X=1.192 $Y=1.167 $X2=0 $Y2=0
cc_203 N_A1_c_198_n N_A_292_55#_c_542_n 0.00113463f $X=1.385 $Y=0.805 $X2=0
+ $Y2=0
cc_204 N_A1_c_198_n N_A_292_55#_c_544_n 0.00383564f $X=1.385 $Y=0.805 $X2=0
+ $Y2=0
cc_205 N_A1_c_204_n N_A_292_55#_c_544_n 0.0059061f $X=1.192 $Y=1.167 $X2=0 $Y2=0
cc_206 N_A2_c_259_n N_A3_M1007_g 0.0120534f $X=1.725 $Y=1.865 $X2=0 $Y2=0
cc_207 N_A2_M1006_g N_A3_M1007_g 0.056981f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_208 N_A2_M1005_g N_A3_M1004_g 0.0249578f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_209 N_A2_c_258_n N_A3_c_302_n 0.0120534f $X=1.725 $Y=1.36 $X2=0 $Y2=0
cc_210 N_A2_c_256_n N_A3_c_303_n 0.0120534f $X=1.725 $Y=1.7 $X2=0 $Y2=0
cc_211 N_A2_M1005_g N_A3_c_304_n 0.0120534f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_212 A2 N_A3_c_304_n 6.37093e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_213 N_A2_M1005_g N_A3_c_305_n 0.00523253f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_214 A2 N_A3_c_305_n 0.0504588f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_215 A2 B1 8.42414e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_216 N_A2_M1006_g N_VPWR_c_462_n 0.0053602f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_217 N_A2_M1006_g N_VPWR_c_457_n 0.010529f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_218 N_A2_M1005_g N_VGND_c_495_n 5.65458e-19 $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_219 N_A2_M1005_g N_VGND_c_496_n 0.00753755f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_220 N_A2_M1005_g N_VGND_c_498_n 0.00337855f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_221 N_A2_M1005_g N_VGND_c_500_n 0.00422396f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_222 N_A2_M1005_g N_A_292_55#_c_542_n 6.54411e-19 $X=1.815 $Y=0.485 $X2=0
+ $Y2=0
cc_223 N_A2_M1005_g N_A_292_55#_c_543_n 0.0135583f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_224 A2 N_A_292_55#_c_543_n 0.00788499f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_225 N_A2_c_258_n N_A_292_55#_c_543_n 2.78643e-19 $X=1.725 $Y=1.36 $X2=0 $Y2=0
cc_226 A2 N_A_292_55#_c_544_n 0.00993463f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_227 N_A2_c_258_n N_A_292_55#_c_544_n 9.71289e-19 $X=1.725 $Y=1.36 $X2=0 $Y2=0
cc_228 N_A2_M1005_g N_A_292_55#_c_546_n 3.22122e-19 $X=1.815 $Y=0.485 $X2=0
+ $Y2=0
cc_229 N_A3_M1004_g N_B1_M1008_g 0.0260851f $X=2.315 $Y=0.485 $X2=0 $Y2=0
cc_230 N_A3_c_304_n N_B1_M1008_g 0.0116081f $X=2.265 $Y=1.245 $X2=0 $Y2=0
cc_231 N_A3_c_305_n N_B1_M1008_g 7.3009e-19 $X=2.265 $Y=1.245 $X2=0 $Y2=0
cc_232 N_A3_M1007_g N_B1_c_346_n 0.0298208f $X=2.175 $Y=2.725 $X2=0 $Y2=0
cc_233 N_A3_c_303_n N_B1_c_346_n 0.0116081f $X=2.265 $Y=1.75 $X2=0 $Y2=0
cc_234 N_A3_c_305_n N_B1_c_346_n 2.31787e-19 $X=2.265 $Y=1.245 $X2=0 $Y2=0
cc_235 N_A3_M1007_g B1 6.0385e-19 $X=2.175 $Y=2.725 $X2=0 $Y2=0
cc_236 N_A3_c_304_n B1 0.0045821f $X=2.265 $Y=1.245 $X2=0 $Y2=0
cc_237 N_A3_c_305_n B1 0.058134f $X=2.265 $Y=1.245 $X2=0 $Y2=0
cc_238 N_A3_c_302_n N_B1_c_348_n 0.0116081f $X=2.265 $Y=1.585 $X2=0 $Y2=0
cc_239 N_A3_M1007_g N_VPWR_c_462_n 0.00523511f $X=2.175 $Y=2.725 $X2=0 $Y2=0
cc_240 N_A3_M1007_g N_VPWR_c_457_n 0.0102117f $X=2.175 $Y=2.725 $X2=0 $Y2=0
cc_241 N_A3_M1004_g N_VGND_c_496_n 0.00466345f $X=2.315 $Y=0.485 $X2=0 $Y2=0
cc_242 N_A3_M1004_g N_VGND_c_499_n 0.0039722f $X=2.315 $Y=0.485 $X2=0 $Y2=0
cc_243 N_A3_M1004_g N_VGND_c_500_n 0.00570792f $X=2.315 $Y=0.485 $X2=0 $Y2=0
cc_244 N_A3_M1004_g N_A_292_55#_c_543_n 0.013218f $X=2.315 $Y=0.485 $X2=0 $Y2=0
cc_245 N_A3_c_304_n N_A_292_55#_c_543_n 0.00285043f $X=2.265 $Y=1.245 $X2=0
+ $Y2=0
cc_246 N_A3_c_305_n N_A_292_55#_c_543_n 0.0261637f $X=2.265 $Y=1.245 $X2=0 $Y2=0
cc_247 N_A3_M1004_g N_A_292_55#_c_546_n 0.00686876f $X=2.315 $Y=0.485 $X2=0
+ $Y2=0
cc_248 N_B1_M1008_g N_C1_c_391_n 0.0487548f $X=2.745 $Y=0.485 $X2=-0.19
+ $Y2=-0.245
cc_249 N_B1_M1009_g N_C1_c_400_n 0.0130671f $X=2.635 $Y=2.725 $X2=0 $Y2=0
cc_250 N_B1_c_346_n N_C1_c_400_n 0.0019268f $X=2.835 $Y=1.7 $X2=0 $Y2=0
cc_251 N_B1_c_346_n N_C1_c_394_n 0.00178227f $X=2.835 $Y=1.7 $X2=0 $Y2=0
cc_252 N_B1_c_346_n N_C1_c_395_n 0.00741861f $X=2.835 $Y=1.7 $X2=0 $Y2=0
cc_253 N_B1_M1008_g N_C1_c_397_n 0.0019432f $X=2.745 $Y=0.485 $X2=0 $Y2=0
cc_254 N_B1_c_348_n N_C1_c_397_n 0.00741861f $X=2.835 $Y=1.36 $X2=0 $Y2=0
cc_255 N_B1_M1009_g N_VPWR_c_459_n 0.00296463f $X=2.635 $Y=2.725 $X2=0 $Y2=0
cc_256 N_B1_c_346_n N_VPWR_c_459_n 5.09294e-19 $X=2.835 $Y=1.7 $X2=0 $Y2=0
cc_257 N_B1_M1009_g N_VPWR_c_462_n 0.00523511f $X=2.635 $Y=2.725 $X2=0 $Y2=0
cc_258 N_B1_M1009_g N_VPWR_c_457_n 0.0101005f $X=2.635 $Y=2.725 $X2=0 $Y2=0
cc_259 N_B1_M1008_g N_VGND_c_499_n 0.00513261f $X=2.745 $Y=0.485 $X2=0 $Y2=0
cc_260 N_B1_M1008_g N_VGND_c_500_n 0.00955386f $X=2.745 $Y=0.485 $X2=0 $Y2=0
cc_261 N_B1_M1008_g N_A_292_55#_c_543_n 0.00489368f $X=2.745 $Y=0.485 $X2=0
+ $Y2=0
cc_262 B1 N_A_292_55#_c_543_n 0.0138955f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_263 N_B1_M1008_g N_A_292_55#_c_546_n 0.00708203f $X=2.745 $Y=0.485 $X2=0
+ $Y2=0
cc_264 N_C1_M1001_g N_VPWR_c_459_n 0.0111201f $X=3.135 $Y=2.725 $X2=0 $Y2=0
cc_265 N_C1_M1001_g N_VPWR_c_464_n 0.00498658f $X=3.135 $Y=2.725 $X2=0 $Y2=0
cc_266 N_C1_M1001_g N_VPWR_c_457_n 0.0097852f $X=3.135 $Y=2.725 $X2=0 $Y2=0
cc_267 N_C1_c_391_n N_VGND_c_499_n 0.00424578f $X=3.105 $Y=0.805 $X2=0 $Y2=0
cc_268 N_C1_c_391_n N_VGND_c_500_n 0.0079407f $X=3.105 $Y=0.805 $X2=0 $Y2=0
cc_269 N_C1_c_392_n N_VGND_c_500_n 0.00651136f $X=3.405 $Y=0.88 $X2=0 $Y2=0
cc_270 C1 N_VGND_c_500_n 0.00982604f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_271 N_C1_c_391_n N_A_292_55#_c_543_n 5.2519e-19 $X=3.105 $Y=0.805 $X2=0 $Y2=0
cc_272 N_C1_c_391_n N_A_292_55#_c_546_n 0.00110333f $X=3.105 $Y=0.805 $X2=0
+ $Y2=0
cc_273 X N_VPWR_c_458_n 0.0294301f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_274 X N_VPWR_c_460_n 0.0392773f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_275 X N_VPWR_c_457_n 0.0225167f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_276 N_X_c_439_n N_VGND_c_497_n 0.0195375f $X=0.7 $Y=0.485 $X2=0 $Y2=0
cc_277 N_X_c_436_n N_VGND_c_497_n 0.0147766f $X=0.232 $Y=0.65 $X2=0 $Y2=0
cc_278 N_X_c_439_n N_VGND_c_500_n 0.0157946f $X=0.7 $Y=0.485 $X2=0 $Y2=0
cc_279 N_X_c_436_n N_VGND_c_500_n 0.0110879f $X=0.232 $Y=0.65 $X2=0 $Y2=0
cc_280 N_VGND_c_498_n N_A_292_55#_c_542_n 0.00869451f $X=1.865 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_500_n N_A_292_55#_c_542_n 0.00703445f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_496_n N_A_292_55#_c_543_n 0.0229339f $X=2.03 $Y=0.465 $X2=0
+ $Y2=0
cc_283 N_VGND_c_498_n N_A_292_55#_c_543_n 0.00226785f $X=1.865 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_499_n N_A_292_55#_c_543_n 0.00226968f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_500_n N_A_292_55#_c_543_n 0.00898392f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_499_n N_A_292_55#_c_546_n 0.013285f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_c_500_n N_A_292_55#_c_546_n 0.0120222f $X=3.6 $Y=0 $X2=0 $Y2=0
