# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfxbp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfxbp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.84000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 1.215000 2.275000 1.885000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.396300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.125000 1.125000 12.760000 1.295000 ;
        RECT 12.125000 1.295000 12.295000 1.985000 ;
        RECT 12.125000 1.985000 12.835000 3.025000 ;
        RECT 12.510000 0.615000 12.760000 1.125000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.398400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.715000 1.920000 15.740000 3.065000 ;
        RECT 15.410000 0.265000 15.740000 1.920000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.955000 1.245000 3.285000 1.915000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 1.515000 0.860000 1.845000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.180000 4.195000 1.510000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.840000 0.085000 ;
        RECT  1.150000  0.085000  1.480000 0.985000 ;
        RECT  2.950000  0.085000  3.280000 1.065000 ;
        RECT  4.280000  0.085000  4.610000 0.650000 ;
        RECT  7.850000  0.085000  8.180000 0.715000 ;
        RECT 11.280000  0.085000 11.530000 0.595000 ;
        RECT 13.300000  0.085000 13.630000 1.075000 ;
        RECT 14.620000  0.085000 14.950000 0.725000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 15.840000 3.415000 ;
        RECT  0.630000 2.025000  0.960000 3.245000 ;
        RECT  2.690000 2.855000  3.020000 3.245000 ;
        RECT  4.320000 2.505000  4.650000 3.245000 ;
        RECT  7.875000 2.015000  8.205000 3.245000 ;
        RECT 10.750000 2.130000 11.080000 3.245000 ;
        RECT 13.015000 1.985000 13.345000 3.245000 ;
        RECT 14.185000 2.335000 14.515000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 15.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.100000 0.605000  0.580000 1.165000 ;
      RECT  0.100000 1.165000  1.685000 1.335000 ;
      RECT  0.100000 1.335000  0.350000 3.065000 ;
      RECT  1.160000 2.065000  1.490000 2.505000 ;
      RECT  1.160000 2.505000  3.550000 2.675000 ;
      RECT  1.160000 2.675000  1.490000 3.065000 ;
      RECT  1.355000 1.335000  1.685000 1.835000 ;
      RECT  1.690000 2.065000  2.625000 2.155000 ;
      RECT  1.690000 2.155000  6.655000 2.325000 ;
      RECT  2.160000 0.605000  2.625000 1.035000 ;
      RECT  2.455000 1.035000  2.625000 2.065000 ;
      RECT  3.220000 2.675000  3.550000 3.065000 ;
      RECT  3.490000 0.310000  3.820000 0.830000 ;
      RECT  3.490000 0.830000  4.910000 1.000000 ;
      RECT  3.790000 1.715000  4.545000 1.975000 ;
      RECT  4.375000 1.000000  4.910000 1.530000 ;
      RECT  4.375000 1.530000  4.545000 1.715000 ;
      RECT  4.850000 1.715000  5.660000 1.975000 ;
      RECT  5.070000 0.310000  5.400000 0.650000 ;
      RECT  5.230000 0.650000  5.400000 1.305000 ;
      RECT  5.230000 1.305000  5.660000 1.715000 ;
      RECT  5.595000 0.265000  7.605000 0.435000 ;
      RECT  5.595000 0.435000  5.845000 1.125000 ;
      RECT  6.025000 0.615000  7.135000 0.785000 ;
      RECT  6.025000 0.785000  6.195000 1.745000 ;
      RECT  6.025000 1.745000  6.655000 2.155000 ;
      RECT  6.025000 2.325000  6.655000 2.755000 ;
      RECT  6.375000 0.965000  6.705000 1.395000 ;
      RECT  6.375000 1.395000  7.185000 1.565000 ;
      RECT  6.855000 1.565000  7.185000 1.665000 ;
      RECT  6.855000 1.665000  8.550000 1.835000 ;
      RECT  6.855000 1.835000  7.185000 2.755000 ;
      RECT  6.885000 0.785000  7.135000 1.215000 ;
      RECT  7.355000 0.435000  7.605000 0.975000 ;
      RECT  7.650000 1.155000  7.980000 1.485000 ;
      RECT  7.810000 0.895000  9.075000 1.065000 ;
      RECT  7.810000 1.065000  7.980000 1.155000 ;
      RECT  8.220000 1.245000  8.550000 1.665000 ;
      RECT  8.705000 0.265000 10.575000 0.435000 ;
      RECT  8.705000 0.435000  9.075000 0.895000 ;
      RECT  8.745000 1.065000  9.075000 2.755000 ;
      RECT  9.255000 0.615000 11.100000 0.785000 ;
      RECT  9.255000 0.785000  9.505000 1.215000 ;
      RECT  9.565000 1.715000 10.080000 1.780000 ;
      RECT  9.565000 1.780000 11.550000 1.950000 ;
      RECT  9.565000 1.950000  9.895000 2.780000 ;
      RECT  9.750000 0.965000 10.080000 1.715000 ;
      RECT 10.565000 0.965000 11.900000 1.135000 ;
      RECT 10.565000 1.135000 10.895000 1.600000 ;
      RECT 10.770000 0.265000 11.100000 0.615000 ;
      RECT 11.220000 1.315000 11.550000 1.780000 ;
      RECT 11.360000 2.130000 11.900000 2.300000 ;
      RECT 11.360000 2.300000 11.690000 2.825000 ;
      RECT 11.730000 0.775000 12.320000 0.945000 ;
      RECT 11.730000 0.945000 11.900000 0.965000 ;
      RECT 11.730000 1.135000 11.900000 2.130000 ;
      RECT 11.990000 0.265000 13.110000 0.435000 ;
      RECT 11.990000 0.435000 12.320000 0.775000 ;
      RECT 12.475000 1.475000 14.165000 1.805000 ;
      RECT 12.940000 0.435000 13.110000 1.475000 ;
      RECT 13.545000 1.985000 14.515000 2.155000 ;
      RECT 13.545000 2.155000 13.875000 3.025000 ;
      RECT 14.090000 0.615000 14.420000 0.905000 ;
      RECT 14.090000 0.905000 14.825000 1.075000 ;
      RECT 14.345000 1.075000 14.825000 1.575000 ;
      RECT 14.345000 1.575000 14.515000 1.985000 ;
  END
END sky130_fd_sc_lp__sdfxbp_lp
