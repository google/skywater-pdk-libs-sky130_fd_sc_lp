# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__a21bo_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a21bo_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.900000 1.345000 5.265000 1.770000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.280000 1.335000 4.645000 1.625000 ;
        RECT 4.475000 1.625000 4.645000 1.940000 ;
        RECT 4.475000 1.940000 5.665000 2.120000 ;
        RECT 5.435000 1.340000 6.010000 1.645000 ;
        RECT 5.435000 1.645000 5.665000 1.940000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.200000 0.805000 1.760000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  1.184400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.930000 2.725000 2.200000 ;
        RECT 0.995000 1.005000 2.480000 1.175000 ;
        RECT 0.995000 1.175000 1.165000 1.800000 ;
        RECT 0.995000 1.800000 2.725000 1.930000 ;
        RECT 1.440000 0.255000 1.630000 1.005000 ;
        RECT 2.300000 0.255000 2.480000 1.005000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 6.240000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 6.430000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.090000  0.255000 0.430000 1.030000 ;
      RECT 0.090000  1.030000 0.270000 1.930000 ;
      RECT 0.090000  1.930000 0.455000 2.370000 ;
      RECT 0.090000  2.370000 3.075000 2.540000 ;
      RECT 0.090000  2.540000 0.455000 3.075000 ;
      RECT 0.600000  0.085000 1.270000 0.835000 ;
      RECT 0.635000  2.710000 0.965000 3.245000 ;
      RECT 1.345000  1.355000 2.820000 1.535000 ;
      RECT 1.495000  2.710000 1.825000 3.245000 ;
      RECT 1.800000  0.085000 2.130000 0.825000 ;
      RECT 2.355000  2.710000 2.685000 3.245000 ;
      RECT 2.650000  0.995000 5.215000 1.165000 ;
      RECT 2.650000  1.165000 2.820000 1.355000 ;
      RECT 2.670000  0.085000 3.475000 0.825000 ;
      RECT 2.905000  1.705000 3.320000 1.875000 ;
      RECT 2.905000  1.875000 3.075000 2.370000 ;
      RECT 2.990000  1.345000 3.320000 1.705000 ;
      RECT 3.245000  2.045000 3.445000 2.905000 ;
      RECT 3.245000  2.905000 4.305000 3.075000 ;
      RECT 3.615000  1.165000 3.945000 2.735000 ;
      RECT 3.645000  0.255000 3.835000 0.995000 ;
      RECT 4.005000  0.085000 4.335000 0.825000 ;
      RECT 4.115000  1.795000 4.305000 2.290000 ;
      RECT 4.115000  2.290000 6.135000 2.460000 ;
      RECT 4.115000  2.460000 4.305000 2.905000 ;
      RECT 4.475000  2.630000 4.805000 3.245000 ;
      RECT 4.515000  0.255000 5.685000 0.425000 ;
      RECT 4.515000  0.425000 4.845000 0.825000 ;
      RECT 4.975000  2.460000 5.205000 3.075000 ;
      RECT 5.015000  0.595000 5.215000 0.995000 ;
      RECT 5.375000  2.630000 5.705000 3.245000 ;
      RECT 5.435000  0.425000 5.685000 1.095000 ;
      RECT 5.835000  1.815000 6.135000 2.290000 ;
      RECT 5.855000  0.085000 6.135000 1.095000 ;
      RECT 5.875000  2.460000 6.135000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__a21bo_4
END LIBRARY
