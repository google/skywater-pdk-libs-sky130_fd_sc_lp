* File: sky130_fd_sc_lp__and4b_4.pxi.spice
* Created: Wed Sep  2 09:33:40 2020
* 
x_PM_SKY130_FD_SC_LP__AND4B_4%A_N N_A_N_M1017_g N_A_N_M1010_g A_N A_N A_N A_N
+ A_N N_A_N_c_90_n N_A_N_c_91_n PM_SKY130_FD_SC_LP__AND4B_4%A_N
x_PM_SKY130_FD_SC_LP__AND4B_4%A_242_23# N_A_242_23#_M1004_d N_A_242_23#_M1001_d
+ N_A_242_23#_M1015_d N_A_242_23#_M1002_g N_A_242_23#_M1000_g
+ N_A_242_23#_M1003_g N_A_242_23#_M1007_g N_A_242_23#_M1008_g
+ N_A_242_23#_M1014_g N_A_242_23#_M1013_g N_A_242_23#_M1016_g
+ N_A_242_23#_c_202_p N_A_242_23#_c_121_n N_A_242_23#_c_131_n
+ N_A_242_23#_c_210_p N_A_242_23#_c_175_p N_A_242_23#_c_140_p
+ N_A_242_23#_c_122_n N_A_242_23#_c_123_n N_A_242_23#_c_124_n
+ N_A_242_23#_c_125_n N_A_242_23#_c_126_n PM_SKY130_FD_SC_LP__AND4B_4%A_242_23#
x_PM_SKY130_FD_SC_LP__AND4B_4%D N_D_M1001_g N_D_M1012_g D N_D_c_246_n
+ N_D_c_247_n PM_SKY130_FD_SC_LP__AND4B_4%D
x_PM_SKY130_FD_SC_LP__AND4B_4%C N_C_M1005_g N_C_M1006_g C N_C_c_284_n
+ N_C_c_285_n PM_SKY130_FD_SC_LP__AND4B_4%C
x_PM_SKY130_FD_SC_LP__AND4B_4%B N_B_M1011_g N_B_M1015_g B B N_B_c_318_n
+ PM_SKY130_FD_SC_LP__AND4B_4%B
x_PM_SKY130_FD_SC_LP__AND4B_4%A_49_133# N_A_49_133#_M1017_s N_A_49_133#_M1010_s
+ N_A_49_133#_M1004_g N_A_49_133#_M1009_g N_A_49_133#_c_352_n
+ N_A_49_133#_c_353_n N_A_49_133#_c_358_n N_A_49_133#_c_359_n
+ N_A_49_133#_c_354_n N_A_49_133#_c_355_n PM_SKY130_FD_SC_LP__AND4B_4%A_49_133#
x_PM_SKY130_FD_SC_LP__AND4B_4%VPWR N_VPWR_M1010_d N_VPWR_M1007_s N_VPWR_M1016_s
+ N_VPWR_M1006_d N_VPWR_M1009_d N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n
+ N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_425_n
+ N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n N_VPWR_c_429_n N_VPWR_c_430_n
+ VPWR N_VPWR_c_431_n N_VPWR_c_417_n N_VPWR_c_433_n N_VPWR_c_434_n
+ PM_SKY130_FD_SC_LP__AND4B_4%VPWR
x_PM_SKY130_FD_SC_LP__AND4B_4%X N_X_M1002_d N_X_M1008_d N_X_M1000_d N_X_M1014_d
+ N_X_c_496_n N_X_c_497_n N_X_c_498_n N_X_c_539_p N_X_c_499_n N_X_c_540_p
+ N_X_c_500_n X X X X N_X_c_521_n PM_SKY130_FD_SC_LP__AND4B_4%X
x_PM_SKY130_FD_SC_LP__AND4B_4%VGND N_VGND_M1017_d N_VGND_M1003_s N_VGND_M1013_s
+ N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n N_VGND_c_548_n N_VGND_c_549_n
+ N_VGND_c_550_n N_VGND_c_551_n N_VGND_c_552_n N_VGND_c_553_n VGND
+ N_VGND_c_554_n N_VGND_c_555_n PM_SKY130_FD_SC_LP__AND4B_4%VGND
cc_1 VNB N_A_N_M1010_g 0.00750648f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.045
cc_2 VNB A_N 0.010532f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_3 VNB N_A_N_c_90_n 0.0419534f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_4 VNB N_A_N_c_91_n 0.0218424f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.195
cc_5 VNB N_A_242_23#_M1002_g 0.026297f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_6 VNB N_A_242_23#_M1003_g 0.0222407f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_7 VNB N_A_242_23#_M1008_g 0.0222554f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.295
cc_8 VNB N_A_242_23#_M1013_g 0.0246709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_242_23#_c_121_n 0.00227867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_242_23#_c_122_n 0.00673785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_242_23#_c_123_n 0.0521254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_242_23#_c_124_n 0.00143519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_242_23#_c_125_n 0.00634034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_242_23#_c_126_n 0.0670688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_D_M1012_g 0.0245716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_D_c_246_n 0.023977f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_17 VNB N_D_c_247_n 0.00328537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C_M1005_g 0.024226f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.875
cc_19 VNB N_C_c_284_n 0.0242961f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_20 VNB N_C_c_285_n 0.0036209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_M1011_g 0.0268186f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.875
cc_22 VNB B 0.00599377f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_23 VNB N_B_c_318_n 0.0223059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_49_133#_M1004_g 0.0298927f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_25 VNB N_A_49_133#_M1009_g 0.00140042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_49_133#_c_352_n 0.00923992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_49_133#_c_353_n 0.0443193f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_28 VNB N_A_49_133#_c_354_n 0.0013024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_49_133#_c_355_n 0.0693276f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.295
cc_30 VNB N_VPWR_c_417_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_496_n 0.00701696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_497_n 6.30069e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_498_n 0.00123683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_499_n 0.00567406f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.195
cc_35 VNB N_X_c_500_n 0.00181876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_545_n 0.00460397f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_37 VNB N_VGND_c_546_n 5.01583e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_547_n 0.00535193f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_39 VNB N_VGND_c_548_n 0.0311972f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.555
cc_40 VNB N_VGND_c_549_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_550_n 0.014949f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.925
cc_42 VNB N_VGND_c_551_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_552_n 0.0164391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_553_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.665
cc_45 VNB N_VGND_c_554_n 0.0575633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_555_n 0.29662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VPB N_A_N_M1010_g 0.0225859f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.045
cc_48 VPB A_N 0.00122212f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_49 VPB N_A_242_23#_M1000_g 0.0218972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_242_23#_M1007_g 0.0185418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_242_23#_M1014_g 0.0185375f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.035
cc_52 VPB N_A_242_23#_M1016_g 0.0186923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_242_23#_c_131_n 0.00129303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_242_23#_c_126_n 0.0121738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_D_M1001_g 0.0193048f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.875
cc_56 VPB N_D_c_246_n 0.00616041f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_57 VPB N_D_c_247_n 0.00246605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_C_M1006_g 0.0206966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_C_c_284_n 0.00638147f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_60 VPB N_C_c_285_n 0.00235431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_B_M1015_g 0.0206033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB B 0.00567615f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_63 VPB N_B_c_318_n 0.00624794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_49_133#_M1009_g 0.022194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_49_133#_c_353_n 0.0356313f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.36
cc_66 VPB N_A_49_133#_c_358_n 0.0315299f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.555
cc_67 VPB N_A_49_133#_c_359_n 0.0126274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_49_133#_c_354_n 0.0355983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_418_n 0.0150717f $X=-0.19 $Y=1.655 $X2=0.707 $Y2=1.36
cc_70 VPB N_VPWR_c_419_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.707 $Y2=1.525
cc_71 VPB N_VPWR_c_420_n 0.0127282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_421_n 0.00213954f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.295
cc_73 VPB N_VPWR_c_422_n 0.0158804f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.665
cc_74 VPB N_VPWR_c_423_n 0.00276847f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_424_n 0.015161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_425_n 0.0283007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_426_n 0.00510611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_427_n 0.0127282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_428_n 0.00436638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_429_n 0.0199508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_430_n 0.00510611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_431_n 0.0113076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_417_n 0.0608418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_433_n 0.00510611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_434_n 0.00510611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_X_c_496_n 0.00309762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 A_N N_A_242_23#_M1002_g 0.00247319f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_88 N_A_N_c_90_n N_A_242_23#_M1002_g 0.0108616f $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_89 N_A_N_c_91_n N_A_242_23#_M1002_g 0.00793174f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_90 A_N N_A_242_23#_M1000_g 0.00124056f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_91 N_A_N_M1010_g N_A_242_23#_c_126_n 0.0157137f $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_92 A_N N_A_49_133#_c_353_n 0.104965f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_93 N_A_N_c_91_n N_A_49_133#_c_353_n 0.0264883f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_94 N_A_N_M1010_g N_A_49_133#_c_358_n 0.00646164f $X=0.605 $Y=2.045 $X2=0
+ $Y2=0
cc_95 A_N N_A_49_133#_c_358_n 0.00940954f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_96 A_N N_VPWR_M1010_d 0.00422784f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_97 N_A_N_M1010_g N_X_c_496_n 0.0028198f $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_98 A_N N_X_c_496_n 0.0724963f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_99 N_A_N_c_90_n N_X_c_496_n 0.00220591f $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_100 A_N N_X_c_498_n 0.0141915f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_101 N_A_N_c_90_n N_X_c_498_n 4.42419e-19 $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_102 N_A_N_c_91_n N_X_c_498_n 4.07562e-19 $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_103 A_N N_VGND_M1017_d 0.00492489f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_104 A_N N_VGND_c_545_n 0.0385531f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_105 N_A_N_c_91_n N_VGND_c_545_n 0.00101849f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_106 A_N N_VGND_c_548_n 0.00708719f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_107 N_A_N_c_91_n N_VGND_c_548_n 0.00295909f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_108 A_N N_VGND_c_555_n 0.00645391f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_109 N_A_N_c_91_n N_VGND_c_555_n 0.00324018f $X=0.707 $Y=1.195 $X2=0 $Y2=0
cc_110 N_A_242_23#_M1016_g N_D_M1001_g 0.0455281f $X=2.575 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_242_23#_c_131_n N_D_M1001_g 0.00388564f $X=2.71 $Y=1.93 $X2=0 $Y2=0
cc_112 N_A_242_23#_c_140_p N_D_M1001_g 0.013472f $X=4.375 $Y=2.095 $X2=0 $Y2=0
cc_113 N_A_242_23#_M1013_g N_D_M1012_g 0.0276321f $X=2.575 $Y=0.665 $X2=0 $Y2=0
cc_114 N_A_242_23#_c_121_n N_D_M1012_g 0.0034595f $X=2.71 $Y=1.415 $X2=0 $Y2=0
cc_115 N_A_242_23#_c_122_n N_D_M1012_g 0.0100999f $X=3.75 $Y=0.71 $X2=0 $Y2=0
cc_116 N_A_242_23#_c_125_n N_D_M1012_g 0.015296f $X=3.295 $Y=0.71 $X2=0 $Y2=0
cc_117 N_A_242_23#_c_121_n N_D_c_246_n 4.22693e-19 $X=2.71 $Y=1.415 $X2=0 $Y2=0
cc_118 N_A_242_23#_c_140_p N_D_c_246_n 0.00257775f $X=4.375 $Y=2.095 $X2=0 $Y2=0
cc_119 N_A_242_23#_c_124_n N_D_c_246_n 0.00183709f $X=2.71 $Y=1.545 $X2=0 $Y2=0
cc_120 N_A_242_23#_c_125_n N_D_c_246_n 0.00339108f $X=3.295 $Y=0.71 $X2=0 $Y2=0
cc_121 N_A_242_23#_c_126_n N_D_c_246_n 0.0205334f $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_122 N_A_242_23#_c_121_n N_D_c_247_n 0.0051848f $X=2.71 $Y=1.415 $X2=0 $Y2=0
cc_123 N_A_242_23#_c_131_n N_D_c_247_n 0.00586273f $X=2.71 $Y=1.93 $X2=0 $Y2=0
cc_124 N_A_242_23#_c_140_p N_D_c_247_n 0.0190809f $X=4.375 $Y=2.095 $X2=0 $Y2=0
cc_125 N_A_242_23#_c_124_n N_D_c_247_n 0.0217824f $X=2.71 $Y=1.545 $X2=0 $Y2=0
cc_126 N_A_242_23#_c_125_n N_D_c_247_n 0.0214937f $X=3.295 $Y=0.71 $X2=0 $Y2=0
cc_127 N_A_242_23#_c_126_n N_D_c_247_n 2.96798e-19 $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_128 N_A_242_23#_c_122_n N_C_M1005_g 0.0354751f $X=3.75 $Y=0.71 $X2=0 $Y2=0
cc_129 N_A_242_23#_c_140_p N_C_M1006_g 0.01462f $X=4.375 $Y=2.095 $X2=0 $Y2=0
cc_130 N_A_242_23#_c_140_p N_C_c_284_n 9.61193e-19 $X=4.375 $Y=2.095 $X2=0 $Y2=0
cc_131 N_A_242_23#_c_122_n N_C_c_284_n 0.00140991f $X=3.75 $Y=0.71 $X2=0 $Y2=0
cc_132 N_A_242_23#_c_140_p N_C_c_285_n 0.0234302f $X=4.375 $Y=2.095 $X2=0 $Y2=0
cc_133 N_A_242_23#_c_122_n N_C_c_285_n 0.0265848f $X=3.75 $Y=0.71 $X2=0 $Y2=0
cc_134 N_A_242_23#_c_123_n N_B_M1011_g 0.0435753f $X=4.805 $Y=0.42 $X2=0 $Y2=0
cc_135 N_A_242_23#_c_140_p N_B_M1015_g 0.0146262f $X=4.375 $Y=2.095 $X2=0 $Y2=0
cc_136 N_A_242_23#_c_140_p B 0.0368176f $X=4.375 $Y=2.095 $X2=0 $Y2=0
cc_137 N_A_242_23#_c_123_n B 0.0606804f $X=4.805 $Y=0.42 $X2=0 $Y2=0
cc_138 N_A_242_23#_c_140_p N_B_c_318_n 8.24464e-19 $X=4.375 $Y=2.095 $X2=0 $Y2=0
cc_139 N_A_242_23#_c_123_n N_B_c_318_n 0.00137675f $X=4.805 $Y=0.42 $X2=0 $Y2=0
cc_140 N_A_242_23#_c_123_n N_A_49_133#_M1004_g 0.034795f $X=4.805 $Y=0.42 $X2=0
+ $Y2=0
cc_141 N_A_242_23#_M1001_d N_A_49_133#_c_358_n 0.00494544f $X=3.155 $Y=1.835
+ $X2=0 $Y2=0
cc_142 N_A_242_23#_M1015_d N_A_49_133#_c_358_n 0.00494544f $X=4.235 $Y=1.835
+ $X2=0 $Y2=0
cc_143 N_A_242_23#_M1000_g N_A_49_133#_c_358_n 0.0144624f $X=1.285 $Y=2.465
+ $X2=0 $Y2=0
cc_144 N_A_242_23#_M1007_g N_A_49_133#_c_358_n 0.0123004f $X=1.715 $Y=2.465
+ $X2=0 $Y2=0
cc_145 N_A_242_23#_M1014_g N_A_49_133#_c_358_n 0.0123004f $X=2.145 $Y=2.465
+ $X2=0 $Y2=0
cc_146 N_A_242_23#_M1016_g N_A_49_133#_c_358_n 0.0165142f $X=2.575 $Y=2.465
+ $X2=0 $Y2=0
cc_147 N_A_242_23#_c_175_p N_A_49_133#_c_358_n 0.0090121f $X=2.795 $Y=2.095
+ $X2=0 $Y2=0
cc_148 N_A_242_23#_c_140_p N_A_49_133#_c_358_n 0.0989194f $X=4.375 $Y=2.095
+ $X2=0 $Y2=0
cc_149 N_A_242_23#_c_123_n N_A_49_133#_c_354_n 0.0127803f $X=4.805 $Y=0.42 $X2=0
+ $Y2=0
cc_150 N_A_242_23#_c_123_n N_A_49_133#_c_355_n 0.0109593f $X=4.805 $Y=0.42 $X2=0
+ $Y2=0
cc_151 N_A_242_23#_c_131_n N_VPWR_M1016_s 0.00112177f $X=2.71 $Y=1.93 $X2=0
+ $Y2=0
cc_152 N_A_242_23#_c_175_p N_VPWR_M1016_s 9.65132e-19 $X=2.795 $Y=2.095 $X2=0
+ $Y2=0
cc_153 N_A_242_23#_c_140_p N_VPWR_M1016_s 0.00645603f $X=4.375 $Y=2.095 $X2=0
+ $Y2=0
cc_154 N_A_242_23#_c_140_p N_VPWR_M1006_d 0.0157822f $X=4.375 $Y=2.095 $X2=0
+ $Y2=0
cc_155 N_A_242_23#_M1000_g N_VPWR_c_418_n 0.0105259f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_242_23#_M1007_g N_VPWR_c_418_n 0.00135454f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_242_23#_M1000_g N_VPWR_c_419_n 0.00135454f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A_242_23#_M1007_g N_VPWR_c_419_n 0.0094624f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A_242_23#_M1014_g N_VPWR_c_419_n 0.0094624f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_242_23#_M1016_g N_VPWR_c_419_n 0.00135454f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_242_23#_M1014_g N_VPWR_c_420_n 0.0036352f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_242_23#_M1016_g N_VPWR_c_420_n 0.0036352f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_242_23#_M1014_g N_VPWR_c_421_n 0.00135454f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_242_23#_M1016_g N_VPWR_c_421_n 0.00948316f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_242_23#_M1000_g N_VPWR_c_427_n 0.0036352f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_242_23#_M1007_g N_VPWR_c_427_n 0.0036352f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_242_23#_M1001_d N_VPWR_c_417_n 0.00360572f $X=3.155 $Y=1.835 $X2=0
+ $Y2=0
cc_168 N_A_242_23#_M1015_d N_VPWR_c_417_n 0.00360572f $X=4.235 $Y=1.835 $X2=0
+ $Y2=0
cc_169 N_A_242_23#_M1000_g N_VPWR_c_417_n 0.00436741f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_242_23#_M1007_g N_VPWR_c_417_n 0.00436741f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_242_23#_M1014_g N_VPWR_c_417_n 0.00436741f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_242_23#_M1016_g N_VPWR_c_417_n 0.00436741f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_242_23#_M1002_g N_X_c_496_n 0.0120086f $X=1.285 $Y=0.665 $X2=0 $Y2=0
cc_174 N_A_242_23#_c_202_p N_X_c_496_n 0.0207007f $X=2.625 $Y=1.545 $X2=0 $Y2=0
cc_175 N_A_242_23#_M1002_g N_X_c_497_n 0.0166776f $X=1.285 $Y=0.665 $X2=0 $Y2=0
cc_176 N_A_242_23#_c_202_p N_X_c_497_n 0.00208315f $X=2.625 $Y=1.545 $X2=0 $Y2=0
cc_177 N_A_242_23#_M1003_g N_X_c_499_n 0.0140849f $X=1.715 $Y=0.665 $X2=0 $Y2=0
cc_178 N_A_242_23#_M1008_g N_X_c_499_n 0.0137525f $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_179 N_A_242_23#_M1013_g N_X_c_499_n 0.00131418f $X=2.575 $Y=0.665 $X2=0 $Y2=0
cc_180 N_A_242_23#_c_202_p N_X_c_499_n 0.0640257f $X=2.625 $Y=1.545 $X2=0 $Y2=0
cc_181 N_A_242_23#_c_121_n N_X_c_499_n 0.00641961f $X=2.71 $Y=1.415 $X2=0 $Y2=0
cc_182 N_A_242_23#_c_210_p N_X_c_499_n 0.00750776f $X=2.795 $Y=1.08 $X2=0 $Y2=0
cc_183 N_A_242_23#_c_126_n N_X_c_499_n 0.00497162f $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_184 N_A_242_23#_c_202_p N_X_c_500_n 0.0190874f $X=2.625 $Y=1.545 $X2=0 $Y2=0
cc_185 N_A_242_23#_c_126_n N_X_c_500_n 0.00253619f $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A_242_23#_M1000_g N_X_c_521_n 0.0175301f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A_242_23#_M1007_g N_X_c_521_n 0.0151877f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_242_23#_M1014_g N_X_c_521_n 0.0151938f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_242_23#_c_202_p N_X_c_521_n 0.0704561f $X=2.625 $Y=1.545 $X2=0 $Y2=0
cc_190 N_A_242_23#_c_126_n N_X_c_521_n 0.00683322f $X=2.575 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A_242_23#_c_210_p N_VGND_M1013_s 9.73829e-19 $X=2.795 $Y=1.08 $X2=0
+ $Y2=0
cc_192 N_A_242_23#_c_125_n N_VGND_M1013_s 0.0026801f $X=3.295 $Y=0.71 $X2=0
+ $Y2=0
cc_193 N_A_242_23#_M1002_g N_VGND_c_545_n 0.00327945f $X=1.285 $Y=0.665 $X2=0
+ $Y2=0
cc_194 N_A_242_23#_M1002_g N_VGND_c_546_n 6.30876e-19 $X=1.285 $Y=0.665 $X2=0
+ $Y2=0
cc_195 N_A_242_23#_M1003_g N_VGND_c_546_n 0.0113264f $X=1.715 $Y=0.665 $X2=0
+ $Y2=0
cc_196 N_A_242_23#_M1008_g N_VGND_c_546_n 0.0113984f $X=2.145 $Y=0.665 $X2=0
+ $Y2=0
cc_197 N_A_242_23#_M1013_g N_VGND_c_546_n 6.43775e-19 $X=2.575 $Y=0.665 $X2=0
+ $Y2=0
cc_198 N_A_242_23#_M1013_g N_VGND_c_547_n 0.00519269f $X=2.575 $Y=0.665 $X2=0
+ $Y2=0
cc_199 N_A_242_23#_c_210_p N_VGND_c_547_n 0.00793424f $X=2.795 $Y=1.08 $X2=0
+ $Y2=0
cc_200 N_A_242_23#_c_125_n N_VGND_c_547_n 0.0181065f $X=3.295 $Y=0.71 $X2=0
+ $Y2=0
cc_201 N_A_242_23#_M1002_g N_VGND_c_550_n 0.00575161f $X=1.285 $Y=0.665 $X2=0
+ $Y2=0
cc_202 N_A_242_23#_M1003_g N_VGND_c_550_n 0.00477554f $X=1.715 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_242_23#_M1008_g N_VGND_c_552_n 0.00477554f $X=2.145 $Y=0.665 $X2=0
+ $Y2=0
cc_204 N_A_242_23#_M1013_g N_VGND_c_552_n 0.00575161f $X=2.575 $Y=0.665 $X2=0
+ $Y2=0
cc_205 N_A_242_23#_c_122_n N_VGND_c_554_n 0.104218f $X=3.75 $Y=0.71 $X2=0 $Y2=0
cc_206 N_A_242_23#_M1004_d N_VGND_c_555_n 0.00212318f $X=4.665 $Y=0.245 $X2=0
+ $Y2=0
cc_207 N_A_242_23#_M1002_g N_VGND_c_555_n 0.0118487f $X=1.285 $Y=0.665 $X2=0
+ $Y2=0
cc_208 N_A_242_23#_M1003_g N_VGND_c_555_n 0.00825815f $X=1.715 $Y=0.665 $X2=0
+ $Y2=0
cc_209 N_A_242_23#_M1008_g N_VGND_c_555_n 0.00825815f $X=2.145 $Y=0.665 $X2=0
+ $Y2=0
cc_210 N_A_242_23#_M1013_g N_VGND_c_555_n 0.0110258f $X=2.575 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_242_23#_c_122_n N_VGND_c_555_n 0.0629508f $X=3.75 $Y=0.71 $X2=0 $Y2=0
cc_212 N_A_242_23#_c_122_n A_645_49# 0.00880535f $X=3.75 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_242_23#_c_125_n A_645_49# 4.57867e-19 $X=3.295 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_214 N_A_242_23#_c_122_n A_717_49# 0.00105839f $X=3.75 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A_242_23#_c_123_n A_717_49# 0.00301315f $X=4.805 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A_242_23#_c_123_n A_825_49# 0.00408134f $X=4.805 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_217 N_D_M1012_g N_C_M1005_g 0.0478602f $X=3.15 $Y=0.665 $X2=0 $Y2=0
cc_218 N_D_M1001_g N_C_M1006_g 0.0535965f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_219 N_D_c_246_n N_C_c_284_n 0.0478602f $X=3.06 $Y=1.51 $X2=0 $Y2=0
cc_220 N_D_c_247_n N_C_c_284_n 0.00227595f $X=3.06 $Y=1.51 $X2=0 $Y2=0
cc_221 N_D_c_246_n N_C_c_285_n 3.80616e-19 $X=3.06 $Y=1.51 $X2=0 $Y2=0
cc_222 N_D_c_247_n N_C_c_285_n 0.0318075f $X=3.06 $Y=1.51 $X2=0 $Y2=0
cc_223 N_D_M1001_g N_A_49_133#_c_358_n 0.0129331f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_224 N_D_M1001_g N_VPWR_c_421_n 0.00325225f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_225 N_D_M1001_g N_VPWR_c_422_n 0.00437171f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_226 N_D_M1001_g N_VPWR_c_423_n 0.00141133f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_227 N_D_M1001_g N_VPWR_c_417_n 0.00633763f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_228 N_D_M1012_g N_VGND_c_547_n 0.00663855f $X=3.15 $Y=0.665 $X2=0 $Y2=0
cc_229 N_D_M1012_g N_VGND_c_554_n 0.00575161f $X=3.15 $Y=0.665 $X2=0 $Y2=0
cc_230 N_D_M1012_g N_VGND_c_555_n 0.0109023f $X=3.15 $Y=0.665 $X2=0 $Y2=0
cc_231 N_C_M1005_g N_B_M1011_g 0.0376705f $X=3.51 $Y=0.665 $X2=0 $Y2=0
cc_232 N_C_M1006_g N_B_M1015_g 0.0310548f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_233 N_C_c_285_n N_B_M1015_g 2.13899e-19 $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_234 N_C_M1005_g B 2.03444e-19 $X=3.51 $Y=0.665 $X2=0 $Y2=0
cc_235 N_C_M1006_g B 2.21216e-19 $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_236 N_C_c_284_n B 0.00123119f $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_237 N_C_c_285_n B 0.0358678f $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_238 N_C_c_284_n N_B_c_318_n 0.0214125f $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_239 N_C_c_285_n N_B_c_318_n 9.97393e-19 $X=3.6 $Y=1.51 $X2=0 $Y2=0
cc_240 N_C_M1006_g N_A_49_133#_c_358_n 0.0132134f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_241 N_C_M1006_g N_VPWR_c_422_n 0.0036352f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_242 N_C_M1006_g N_VPWR_c_423_n 0.0103197f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_243 N_C_M1006_g N_VPWR_c_417_n 0.00439469f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_244 N_C_M1005_g N_VGND_c_554_n 0.00351226f $X=3.51 $Y=0.665 $X2=0 $Y2=0
cc_245 N_C_M1005_g N_VGND_c_555_n 0.00542362f $X=3.51 $Y=0.665 $X2=0 $Y2=0
cc_246 N_B_M1011_g N_A_49_133#_M1004_g 0.0378729f $X=4.05 $Y=0.665 $X2=0 $Y2=0
cc_247 N_B_M1015_g N_A_49_133#_M1009_g 0.0537565f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_248 B N_A_49_133#_M1009_g 0.00987555f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_249 B N_A_49_133#_c_352_n 0.0124137f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_250 N_B_c_318_n N_A_49_133#_c_352_n 0.0214293f $X=4.14 $Y=1.51 $X2=0 $Y2=0
cc_251 N_B_M1015_g N_A_49_133#_c_358_n 0.0135561f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_252 B N_A_49_133#_c_354_n 0.0320446f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_253 N_B_M1015_g N_VPWR_c_423_n 0.0101551f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_254 N_B_M1015_g N_VPWR_c_424_n 0.00256693f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_255 N_B_M1015_g N_VPWR_c_429_n 0.00437171f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_256 N_B_M1015_g N_VPWR_c_417_n 0.0067625f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_257 N_B_M1011_g N_VGND_c_554_n 0.00351226f $X=4.05 $Y=0.665 $X2=0 $Y2=0
cc_258 N_B_M1011_g N_VGND_c_555_n 0.00584707f $X=4.05 $Y=0.665 $X2=0 $Y2=0
cc_259 N_A_49_133#_c_358_n N_VPWR_M1010_d 0.00631102f $X=4.825 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_49_133#_c_358_n N_VPWR_M1007_s 0.00349458f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_261 N_A_49_133#_c_358_n N_VPWR_M1016_s 0.00506052f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_262 N_A_49_133#_c_358_n N_VPWR_M1006_d 0.010701f $X=4.825 $Y=2.52 $X2=0 $Y2=0
cc_263 N_A_49_133#_c_358_n N_VPWR_M1009_d 0.00694561f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_264 N_A_49_133#_c_354_n N_VPWR_M1009_d 0.0102885f $X=4.99 $Y=1.46 $X2=0 $Y2=0
cc_265 N_A_49_133#_c_358_n N_VPWR_c_418_n 0.021205f $X=4.825 $Y=2.52 $X2=0 $Y2=0
cc_266 N_A_49_133#_c_358_n N_VPWR_c_419_n 0.0164573f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_267 N_A_49_133#_c_358_n N_VPWR_c_420_n 0.00670101f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_268 N_A_49_133#_c_358_n N_VPWR_c_421_n 0.0206179f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_269 N_A_49_133#_c_358_n N_VPWR_c_422_n 0.00742693f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_270 N_A_49_133#_c_358_n N_VPWR_c_423_n 0.0210884f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_271 N_A_49_133#_M1009_g N_VPWR_c_424_n 0.011903f $X=4.59 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A_49_133#_c_358_n N_VPWR_c_424_n 0.0222812f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_273 N_A_49_133#_c_358_n N_VPWR_c_425_n 0.00692254f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_274 N_A_49_133#_c_359_n N_VPWR_c_425_n 0.00426603f $X=0.455 $Y=2.52 $X2=0
+ $Y2=0
cc_275 N_A_49_133#_c_358_n N_VPWR_c_427_n 0.00670101f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_276 N_A_49_133#_M1009_g N_VPWR_c_429_n 0.0036352f $X=4.59 $Y=2.465 $X2=0
+ $Y2=0
cc_277 N_A_49_133#_c_358_n N_VPWR_c_429_n 0.00950964f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_278 N_A_49_133#_c_358_n N_VPWR_c_431_n 0.00315343f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_279 N_A_49_133#_M1009_g N_VPWR_c_417_n 0.00439469f $X=4.59 $Y=2.465 $X2=0
+ $Y2=0
cc_280 N_A_49_133#_c_358_n N_VPWR_c_417_n 0.0835084f $X=4.825 $Y=2.52 $X2=0
+ $Y2=0
cc_281 N_A_49_133#_c_359_n N_VPWR_c_417_n 0.00710942f $X=0.455 $Y=2.52 $X2=0
+ $Y2=0
cc_282 N_A_49_133#_c_358_n N_X_M1000_d 0.00494544f $X=4.825 $Y=2.52 $X2=0 $Y2=0
cc_283 N_A_49_133#_c_358_n N_X_M1014_d 0.00494544f $X=4.825 $Y=2.52 $X2=0 $Y2=0
cc_284 N_A_49_133#_c_353_n N_X_c_496_n 0.00250461f $X=0.37 $Y=0.87 $X2=0 $Y2=0
cc_285 N_A_49_133#_c_358_n N_X_c_496_n 0.0136761f $X=4.825 $Y=2.52 $X2=0 $Y2=0
cc_286 N_A_49_133#_c_358_n N_X_c_521_n 0.071525f $X=4.825 $Y=2.52 $X2=0 $Y2=0
cc_287 N_A_49_133#_c_353_n N_VGND_c_548_n 0.00425501f $X=0.37 $Y=0.87 $X2=0
+ $Y2=0
cc_288 N_A_49_133#_M1004_g N_VGND_c_554_n 0.00351226f $X=4.59 $Y=0.665 $X2=0
+ $Y2=0
cc_289 N_A_49_133#_M1004_g N_VGND_c_555_n 0.00665279f $X=4.59 $Y=0.665 $X2=0
+ $Y2=0
cc_290 N_A_49_133#_c_353_n N_VGND_c_555_n 0.00719928f $X=0.37 $Y=0.87 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_417_n N_X_M1000_d 0.00360572f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_292 N_VPWR_c_417_n N_X_M1014_d 0.00360572f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_293 N_VPWR_M1010_d N_X_c_496_n 0.00719849f $X=0.68 $Y=1.835 $X2=0 $Y2=0
cc_294 N_VPWR_M1007_s N_X_c_521_n 0.00343809f $X=1.79 $Y=1.835 $X2=0 $Y2=0
cc_295 N_X_c_498_n N_VGND_M1017_d 0.00200503f $X=1.165 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_296 N_X_c_499_n N_VGND_M1003_s 0.00176461f $X=2.265 $Y=1.16 $X2=0 $Y2=0
cc_297 N_X_c_498_n N_VGND_c_545_n 0.014423f $X=1.165 $Y=1.16 $X2=0 $Y2=0
cc_298 N_X_c_499_n N_VGND_c_546_n 0.0170777f $X=2.265 $Y=1.16 $X2=0 $Y2=0
cc_299 N_X_c_539_p N_VGND_c_550_n 0.0138717f $X=1.5 $Y=0.42 $X2=0 $Y2=0
cc_300 N_X_c_540_p N_VGND_c_552_n 0.0124525f $X=2.36 $Y=0.42 $X2=0 $Y2=0
cc_301 N_X_M1002_d N_VGND_c_555_n 0.00397496f $X=1.36 $Y=0.245 $X2=0 $Y2=0
cc_302 N_X_M1008_d N_VGND_c_555_n 0.00536646f $X=2.22 $Y=0.245 $X2=0 $Y2=0
cc_303 N_X_c_539_p N_VGND_c_555_n 0.00886411f $X=1.5 $Y=0.42 $X2=0 $Y2=0
cc_304 N_X_c_540_p N_VGND_c_555_n 0.00730901f $X=2.36 $Y=0.42 $X2=0 $Y2=0
cc_305 N_VGND_c_555_n A_645_49# 0.00412397f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
cc_306 N_VGND_c_555_n A_717_49# 0.00313651f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
cc_307 N_VGND_c_555_n A_825_49# 0.00313651f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
