* File: sky130_fd_sc_lp__decap_4.pex.spice
* Created: Wed Sep  2 09:42:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAP_4%VGND 1 7 9 11 14 17 19 26 29 32 42
r27 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r28 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 36 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r30 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r31 33 38 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.25
+ $Y2=0
r32 33 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=1.2 $Y2=0
r33 32 41 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.685
+ $Y2=0
r34 32 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.2
+ $Y2=0
r35 29 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r36 29 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r37 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.77 $X2=0.575 $Y2=1.77
r38 23 26 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.335 $Y=1.77
+ $X2=0.575 $Y2=1.77
r39 19 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.615 $Y=0.36
+ $X2=1.615 $Y2=1.04
r40 17 41 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.685 $Y2=0
r41 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0.36
r42 14 16 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.335 $Y=0.38
+ $X2=0.335 $Y2=1.06
r43 12 23 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.335 $Y=1.605
+ $X2=0.335 $Y2=1.77
r44 12 16 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.335 $Y=1.605
+ $X2=0.335 $Y2=1.06
r45 11 38 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.25 $Y2=0
r46 11 14 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.38
r47 7 27 22.6591 $w=1e-06 $l=4.09268e-07 $layer=POLY_cond $X=0.91 $Y=1.935
+ $X2=0.575 $Y2=1.77
r48 7 9 33.9353 $w=1e-06 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.935 $X2=0.91
+ $Y2=2.595
r49 1 21 121.333 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=1.615 $Y2=1.04
r50 1 19 121.333 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=1.615 $Y2=0.36
r51 1 16 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=0.335 $Y2=1.06
r52 1 14 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=0.335 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DECAP_4%VPWR 1 7 9 14 16 23 25 28 30 40
r27 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r28 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 34 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r30 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r31 31 36 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r32 31 33 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 30 39 4.56733 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.652 $Y2=3.33
r34 30 33 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.2 $Y2=3.33
r35 25 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r36 25 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 21 28 44.365 $w=8.68e-07 $l=9.34987e-07 $layer=POLY_cond $X=1.345 $Y=1.51
+ $X2=0.992 $Y2=0.735
r38 20 23 7.05226 $w=3.33e-07 $l=2.05e-07 $layer=LI1_cond $X=1.345 $Y=1.507
+ $X2=1.55 $Y2=1.507
r39 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.345
+ $Y=1.51 $X2=1.345 $Y2=1.51
r40 16 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.29
+ $X2=1.55 $Y2=2.97
r41 14 39 3.19884 $w=3.3e-07 $l=1.38109e-07 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.652 $Y2=3.33
r42 14 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.55 $Y2=2.97
r43 13 23 0.808037 $w=3.3e-07 $l=1.68e-07 $layer=LI1_cond $X=1.55 $Y=1.675
+ $X2=1.55 $Y2=1.507
r44 13 16 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.55 $Y=1.675
+ $X2=1.55 $Y2=2.29
r45 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.27 $X2=0.26
+ $Y2=2.95
r46 7 36 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r47 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r48 1 18 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.095 $X2=1.55 $Y2=2.97
r49 1 16 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.095 $X2=1.55 $Y2=2.29
r50 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.095 $X2=0.26 $Y2=2.95
r51 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.095 $X2=0.26 $Y2=2.27
.ends

