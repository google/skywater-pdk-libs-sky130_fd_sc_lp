* File: sky130_fd_sc_lp__dlrtp_1.pxi.spice
* Created: Fri Aug 28 10:26:57 2020
* 
x_PM_SKY130_FD_SC_LP__DLRTP_1%D N_D_c_145_n N_D_M1015_g N_D_M1000_g N_D_c_147_n
+ D D D N_D_c_149_n N_D_c_150_n PM_SKY130_FD_SC_LP__DLRTP_1%D
x_PM_SKY130_FD_SC_LP__DLRTP_1%GATE N_GATE_M1013_g N_GATE_c_180_n N_GATE_M1014_g
+ N_GATE_c_182_n GATE GATE GATE N_GATE_c_184_n N_GATE_c_185_n
+ PM_SKY130_FD_SC_LP__DLRTP_1%GATE
x_PM_SKY130_FD_SC_LP__DLRTP_1%A_249_70# N_A_249_70#_M1013_d N_A_249_70#_M1014_d
+ N_A_249_70#_c_222_n N_A_249_70#_M1001_g N_A_249_70#_c_223_n
+ N_A_249_70#_M1012_g N_A_249_70#_M1007_g N_A_249_70#_c_224_n
+ N_A_249_70#_c_225_n N_A_249_70#_M1009_g N_A_249_70#_c_241_n
+ N_A_249_70#_c_242_n N_A_249_70#_c_227_n N_A_249_70#_c_228_n
+ N_A_249_70#_c_229_n N_A_249_70#_c_230_n N_A_249_70#_c_231_n
+ N_A_249_70#_c_244_n N_A_249_70#_c_232_n N_A_249_70#_c_233_n
+ N_A_249_70#_c_234_n N_A_249_70#_c_235_n PM_SKY130_FD_SC_LP__DLRTP_1%A_249_70#
x_PM_SKY130_FD_SC_LP__DLRTP_1%A_41_464# N_A_41_464#_M1000_s N_A_41_464#_M1015_s
+ N_A_41_464#_M1003_g N_A_41_464#_M1002_g N_A_41_464#_c_372_n
+ N_A_41_464#_c_373_n N_A_41_464#_c_368_n N_A_41_464#_c_375_n
+ N_A_41_464#_c_376_n N_A_41_464#_c_377_n N_A_41_464#_c_378_n
+ N_A_41_464#_c_379_n N_A_41_464#_c_380_n N_A_41_464#_c_381_n
+ N_A_41_464#_c_369_n N_A_41_464#_c_370_n PM_SKY130_FD_SC_LP__DLRTP_1%A_41_464#
x_PM_SKY130_FD_SC_LP__DLRTP_1%A_371_473# N_A_371_473#_M1012_s
+ N_A_371_473#_M1001_s N_A_371_473#_M1005_g N_A_371_473#_M1017_g
+ N_A_371_473#_c_466_n N_A_371_473#_c_467_n N_A_371_473#_c_468_n
+ N_A_371_473#_c_469_n N_A_371_473#_c_477_n N_A_371_473#_c_478_n
+ N_A_371_473#_c_479_n N_A_371_473#_c_470_n N_A_371_473#_c_471_n
+ N_A_371_473#_c_472_n N_A_371_473#_c_473_n N_A_371_473#_c_480_n
+ N_A_371_473#_c_481_n PM_SKY130_FD_SC_LP__DLRTP_1%A_371_473#
x_PM_SKY130_FD_SC_LP__DLRTP_1%A_809_21# N_A_809_21#_M1006_s N_A_809_21#_M1004_d
+ N_A_809_21#_c_581_n N_A_809_21#_M1010_g N_A_809_21#_M1008_g
+ N_A_809_21#_M1011_g N_A_809_21#_M1018_g N_A_809_21#_c_583_n
+ N_A_809_21#_c_591_n N_A_809_21#_c_592_n N_A_809_21#_c_584_n
+ N_A_809_21#_c_585_n N_A_809_21#_c_614_p N_A_809_21#_c_615_p
+ N_A_809_21#_c_645_p N_A_809_21#_c_594_n N_A_809_21#_c_611_p
+ N_A_809_21#_c_586_n N_A_809_21#_c_587_n N_A_809_21#_c_588_n
+ PM_SKY130_FD_SC_LP__DLRTP_1%A_809_21#
x_PM_SKY130_FD_SC_LP__DLRTP_1%A_659_47# N_A_659_47#_M1005_d N_A_659_47#_M1007_d
+ N_A_659_47#_M1006_g N_A_659_47#_M1004_g N_A_659_47#_c_705_n
+ N_A_659_47#_c_706_n N_A_659_47#_c_716_n N_A_659_47#_c_720_n
+ N_A_659_47#_c_707_n N_A_659_47#_c_726_n N_A_659_47#_c_708_n
+ N_A_659_47#_c_709_n N_A_659_47#_c_710_n N_A_659_47#_c_736_n
+ N_A_659_47#_c_711_n N_A_659_47#_c_712_n PM_SKY130_FD_SC_LP__DLRTP_1%A_659_47#
x_PM_SKY130_FD_SC_LP__DLRTP_1%RESET_B N_RESET_B_M1019_g N_RESET_B_M1016_g
+ RESET_B RESET_B RESET_B RESET_B RESET_B N_RESET_B_c_813_n N_RESET_B_c_814_n
+ RESET_B PM_SKY130_FD_SC_LP__DLRTP_1%RESET_B
x_PM_SKY130_FD_SC_LP__DLRTP_1%VPWR N_VPWR_M1015_d N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_M1016_d N_VPWR_c_859_n N_VPWR_c_860_n N_VPWR_c_861_n N_VPWR_c_862_n
+ N_VPWR_c_863_n VPWR N_VPWR_c_864_n N_VPWR_c_865_n N_VPWR_c_866_n
+ N_VPWR_c_858_n N_VPWR_c_868_n N_VPWR_c_869_n N_VPWR_c_870_n
+ PM_SKY130_FD_SC_LP__DLRTP_1%VPWR
x_PM_SKY130_FD_SC_LP__DLRTP_1%Q N_Q_M1011_d N_Q_M1018_d N_Q_c_941_n N_Q_c_942_n
+ Q Q Q Q N_Q_c_943_n PM_SKY130_FD_SC_LP__DLRTP_1%Q
x_PM_SKY130_FD_SC_LP__DLRTP_1%VGND N_VGND_M1000_d N_VGND_M1012_d N_VGND_M1010_d
+ N_VGND_M1019_d N_VGND_c_963_n N_VGND_c_964_n N_VGND_c_965_n N_VGND_c_966_n
+ N_VGND_c_967_n N_VGND_c_968_n VGND N_VGND_c_969_n N_VGND_c_970_n
+ N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n N_VGND_c_974_n N_VGND_c_975_n
+ PM_SKY130_FD_SC_LP__DLRTP_1%VGND
cc_1 VNB N_D_c_145_n 0.0213841f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.343
cc_2 VNB N_D_M1015_g 0.0064277f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.64
cc_3 VNB N_D_c_147_n 0.0250537f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.55
cc_4 VNB D 0.00397283f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_5 VNB N_D_c_149_n 0.0255231f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_6 VNB N_D_c_150_n 0.0224261f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.88
cc_7 VNB N_GATE_c_180_n 0.0250155f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.64
cc_8 VNB N_GATE_M1014_g 0.00667554f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.56
cc_9 VNB N_GATE_c_182_n 0.0199943f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.55
cc_10 VNB GATE 0.00865102f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_11 VNB N_GATE_c_184_n 0.0182715f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_12 VNB N_GATE_c_185_n 0.0213431f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.88
cc_13 VNB N_A_249_70#_c_222_n 0.0353204f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.56
cc_14 VNB N_A_249_70#_c_223_n 0.0196964f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_15 VNB N_A_249_70#_c_224_n 0.0162136f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.88
cc_16 VNB N_A_249_70#_c_225_n 0.00807223f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.925
cc_17 VNB N_A_249_70#_M1009_g 0.0372302f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.045
cc_18 VNB N_A_249_70#_c_227_n 0.0135321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_249_70#_c_228_n 0.020087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_249_70#_c_229_n 0.016862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_249_70#_c_230_n 0.00265019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_249_70#_c_231_n 0.0111371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_249_70#_c_232_n 0.00232174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_249_70#_c_233_n 0.00503425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_249_70#_c_234_n 0.0160071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_249_70#_c_235_n 0.0459606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_41_464#_M1003_g 0.0555522f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_28 VNB N_A_41_464#_c_368_n 0.0628147f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.925
cc_29 VNB N_A_41_464#_c_369_n 0.00412769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_41_464#_c_370_n 0.0175432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_371_473#_M1005_g 0.0264986f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.56
cc_32 VNB N_A_371_473#_c_466_n 0.0125511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_371_473#_c_467_n 0.00531428f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_34 VNB N_A_371_473#_c_468_n 0.0113757f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.925
cc_35 VNB N_A_371_473#_c_469_n 0.0059897f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.045
cc_36 VNB N_A_371_473#_c_470_n 0.00636425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_371_473#_c_471_n 0.00157813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_371_473#_c_472_n 0.0126825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_371_473#_c_473_n 0.0300411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_809_21#_c_581_n 0.0191232f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.88
cc_41 VNB N_A_809_21#_M1011_g 0.0243733f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_42 VNB N_A_809_21#_c_583_n 0.0231338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_809_21#_c_584_n 0.00240204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_809_21#_c_585_n 0.00163828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_809_21#_c_586_n 0.0040335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_809_21#_c_587_n 0.0259394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_809_21#_c_588_n 0.0404406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_659_47#_M1006_g 0.0207961f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.56
cc_49 VNB N_A_659_47#_c_705_n 0.0325311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_659_47#_c_706_n 0.010488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_659_47#_c_707_n 0.0092328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_659_47#_c_708_n 5.86216e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_659_47#_c_709_n 0.0132658f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.665
cc_54 VNB N_A_659_47#_c_710_n 0.00233604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_659_47#_c_711_n 0.00975489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_659_47#_c_712_n 0.00892717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_M1019_g 0.018795f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.55
cc_58 VNB RESET_B 0.00149042f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.56
cc_59 VNB RESET_B 0.00497525f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_60 VNB N_RESET_B_c_813_n 0.0249092f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.925
cc_61 VNB N_RESET_B_c_814_n 9.13189e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VPWR_c_858_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_Q_c_941_n 0.0308122f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.56
cc_64 VNB N_Q_c_942_n 0.0108163f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_65 VNB N_Q_c_943_n 0.0231323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_963_n 0.00924355f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.045
cc_67 VNB N_VGND_c_964_n 0.00250426f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.925
cc_68 VNB N_VGND_c_965_n 0.00933245f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.295
cc_69 VNB N_VGND_c_966_n 0.00828611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_967_n 0.0326946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_968_n 0.00413547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_969_n 0.0379644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_970_n 0.038269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_971_n 0.0216814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_972_n 0.37535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_973_n 0.0291634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_974_n 0.00414071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_975_n 0.00478125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VPB N_D_M1015_g 0.0576313f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.64
cc_80 VPB D 0.00432776f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_81 VPB N_GATE_M1014_g 0.0525326f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.56
cc_82 VPB GATE 0.0075402f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_83 VPB N_A_249_70#_c_222_n 0.00823582f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.56
cc_84 VPB N_A_249_70#_M1001_g 0.0262946f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_85 VPB N_A_249_70#_M1007_g 0.0497057f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.045
cc_86 VPB N_A_249_70#_c_224_n 0.0100472f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=0.88
cc_87 VPB N_A_249_70#_c_225_n 3.95165e-19 $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.925
cc_88 VPB N_A_249_70#_c_241_n 0.0762637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_249_70#_c_242_n 0.00860329f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.665
cc_90 VPB N_A_249_70#_c_228_n 0.00632426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_249_70#_c_244_n 0.00581445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_41_464#_M1002_g 0.0212166f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_41_464#_c_372_n 0.0237526f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=1.045
cc_94 VPB N_A_41_464#_c_373_n 0.0385219f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.045
cc_95 VPB N_A_41_464#_c_368_n 0.0157013f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.925
cc_96 VPB N_A_41_464#_c_375_n 0.0372332f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.295
cc_97 VPB N_A_41_464#_c_376_n 0.0182604f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.665
cc_98 VPB N_A_41_464#_c_377_n 0.00171253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_41_464#_c_378_n 0.0163816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_41_464#_c_379_n 0.00137942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_41_464#_c_380_n 0.00202821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_41_464#_c_381_n 0.00770964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_41_464#_c_369_n 0.00242568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_41_464#_c_370_n 0.00873377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_371_473#_M1017_g 0.0185645f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_106 VPB N_A_371_473#_c_467_n 0.0052655f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.045
cc_107 VPB N_A_371_473#_c_469_n 0.00803827f $X=-0.19 $Y=1.655 $X2=0.745
+ $Y2=1.045
cc_108 VPB N_A_371_473#_c_477_n 0.0110867f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.295
cc_109 VPB N_A_371_473#_c_478_n 3.20306e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_371_473#_c_479_n 0.00251057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_371_473#_c_480_n 0.0332719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_371_473#_c_481_n 0.00358839f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_809_21#_M1008_g 0.0227682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_809_21#_M1018_g 0.023547f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_809_21#_c_591_n 0.00803573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_809_21#_c_592_n 0.0319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_809_21#_c_585_n 0.00302819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_809_21#_c_594_n 0.00133778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_809_21#_c_586_n 3.95463e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_809_21#_c_587_n 0.00676868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_809_21#_c_588_n 0.0193871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_659_47#_M1004_g 0.0239246f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_123 VPB N_A_659_47#_c_705_n 0.0134213f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_659_47#_c_706_n 3.27749e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_659_47#_c_716_n 0.00704323f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.045
cc_126 VPB N_A_659_47#_c_707_n 0.0121832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_659_47#_c_711_n 0.0043672f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_RESET_B_M1016_g 0.0183094f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.88
cc_129 VPB N_RESET_B_c_813_n 0.00674372f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.925
cc_130 VPB N_RESET_B_c_814_n 0.00214788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_859_n 0.0100469f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=1.045
cc_132 VPB N_VPWR_c_860_n 0.00885927f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.925
cc_133 VPB N_VPWR_c_861_n 0.00505115f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.295
cc_134 VPB N_VPWR_c_862_n 0.0173748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_863_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_864_n 0.0419316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_865_n 0.0388713f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_866_n 0.0198429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_858_n 0.0969181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_868_n 0.0243656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_869_n 0.0043944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_870_n 0.0269064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB Q 0.0540904f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_Q_c_943_n 0.00934303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 N_D_c_145_n N_GATE_c_180_n 0.0141165f $X=0.677 $Y=1.343 $X2=0 $Y2=0
cc_146 N_D_M1015_g N_GATE_M1014_g 0.0253859f $X=0.545 $Y=2.64 $X2=0 $Y2=0
cc_147 D N_GATE_M1014_g 8.0025e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_148 N_D_c_147_n N_GATE_c_182_n 0.0141165f $X=0.677 $Y=1.55 $X2=0 $Y2=0
cc_149 D GATE 0.0746948f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_150 N_D_c_149_n GATE 0.00404989f $X=0.72 $Y=1.045 $X2=0 $Y2=0
cc_151 D N_GATE_c_184_n 7.17666e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_152 N_D_c_149_n N_GATE_c_184_n 0.0141165f $X=0.72 $Y=1.045 $X2=0 $Y2=0
cc_153 N_D_c_150_n N_GATE_c_185_n 0.0143642f $X=0.677 $Y=0.88 $X2=0 $Y2=0
cc_154 D N_A_41_464#_c_368_n 0.0735381f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_155 N_D_c_149_n N_A_41_464#_c_368_n 0.0320974f $X=0.72 $Y=1.045 $X2=0 $Y2=0
cc_156 N_D_c_150_n N_A_41_464#_c_368_n 0.00413045f $X=0.677 $Y=0.88 $X2=0 $Y2=0
cc_157 N_D_M1015_g N_A_41_464#_c_375_n 0.00594899f $X=0.545 $Y=2.64 $X2=0 $Y2=0
cc_158 N_D_M1015_g N_A_41_464#_c_376_n 0.0219015f $X=0.545 $Y=2.64 $X2=0 $Y2=0
cc_159 N_D_c_147_n N_A_41_464#_c_376_n 0.00182204f $X=0.677 $Y=1.55 $X2=0 $Y2=0
cc_160 D N_A_41_464#_c_376_n 0.0201012f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_161 N_D_M1015_g N_A_41_464#_c_377_n 0.00216509f $X=0.545 $Y=2.64 $X2=0 $Y2=0
cc_162 N_D_M1015_g N_VPWR_c_859_n 0.00340641f $X=0.545 $Y=2.64 $X2=0 $Y2=0
cc_163 N_D_M1015_g N_VPWR_c_858_n 0.00913333f $X=0.545 $Y=2.64 $X2=0 $Y2=0
cc_164 N_D_M1015_g N_VPWR_c_868_n 0.00461464f $X=0.545 $Y=2.64 $X2=0 $Y2=0
cc_165 D N_VGND_c_963_n 0.0132262f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_166 N_D_c_149_n N_VGND_c_963_n 0.00200223f $X=0.72 $Y=1.045 $X2=0 $Y2=0
cc_167 N_D_c_150_n N_VGND_c_963_n 0.00557049f $X=0.677 $Y=0.88 $X2=0 $Y2=0
cc_168 D N_VGND_c_972_n 0.00382542f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_169 N_D_c_149_n N_VGND_c_972_n 0.00100004f $X=0.72 $Y=1.045 $X2=0 $Y2=0
cc_170 N_D_c_150_n N_VGND_c_972_n 0.00866141f $X=0.677 $Y=0.88 $X2=0 $Y2=0
cc_171 N_D_c_150_n N_VGND_c_973_n 0.00478016f $X=0.677 $Y=0.88 $X2=0 $Y2=0
cc_172 N_GATE_c_180_n N_A_249_70#_c_222_n 0.00317452f $X=1.265 $Y=1.38 $X2=0
+ $Y2=0
cc_173 N_GATE_M1014_g N_A_249_70#_c_241_n 0.0205338f $X=1.17 $Y=2.64 $X2=0 $Y2=0
cc_174 N_GATE_M1014_g N_A_249_70#_c_228_n 0.00773225f $X=1.17 $Y=2.64 $X2=0
+ $Y2=0
cc_175 GATE N_A_249_70#_c_228_n 0.072954f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_176 N_GATE_c_184_n N_A_249_70#_c_228_n 0.00800895f $X=1.27 $Y=1.045 $X2=0
+ $Y2=0
cc_177 N_GATE_c_185_n N_A_249_70#_c_228_n 0.00486249f $X=1.265 $Y=0.88 $X2=0
+ $Y2=0
cc_178 GATE N_A_249_70#_c_231_n 0.0105465f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_179 N_GATE_c_184_n N_A_249_70#_c_231_n 0.00329097f $X=1.27 $Y=1.045 $X2=0
+ $Y2=0
cc_180 N_GATE_c_185_n N_A_249_70#_c_231_n 0.00452475f $X=1.265 $Y=0.88 $X2=0
+ $Y2=0
cc_181 GATE N_A_249_70#_c_244_n 6.52566e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_182 N_GATE_c_184_n N_A_249_70#_c_235_n 0.00317452f $X=1.27 $Y=1.045 $X2=0
+ $Y2=0
cc_183 N_GATE_M1014_g N_A_41_464#_c_376_n 0.00735805f $X=1.17 $Y=2.64 $X2=0
+ $Y2=0
cc_184 GATE N_A_41_464#_c_376_n 0.0131467f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_185 N_GATE_M1014_g N_A_41_464#_c_377_n 0.0252916f $X=1.17 $Y=2.64 $X2=0 $Y2=0
cc_186 N_GATE_M1014_g N_A_41_464#_c_378_n 0.00788427f $X=1.17 $Y=2.64 $X2=0
+ $Y2=0
cc_187 N_GATE_M1014_g N_A_41_464#_c_379_n 0.00346309f $X=1.17 $Y=2.64 $X2=0
+ $Y2=0
cc_188 N_GATE_c_185_n N_A_371_473#_c_470_n 0.00204328f $X=1.265 $Y=0.88 $X2=0
+ $Y2=0
cc_189 N_GATE_M1014_g N_VPWR_c_859_n 0.00266777f $X=1.17 $Y=2.64 $X2=0 $Y2=0
cc_190 N_GATE_M1014_g N_VPWR_c_864_n 0.00278184f $X=1.17 $Y=2.64 $X2=0 $Y2=0
cc_191 N_GATE_M1014_g N_VPWR_c_858_n 0.00360052f $X=1.17 $Y=2.64 $X2=0 $Y2=0
cc_192 GATE N_VGND_c_963_n 4.4689e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_193 N_GATE_c_185_n N_VGND_c_963_n 0.00526137f $X=1.265 $Y=0.88 $X2=0 $Y2=0
cc_194 N_GATE_c_185_n N_VGND_c_969_n 0.00448345f $X=1.265 $Y=0.88 $X2=0 $Y2=0
cc_195 GATE N_VGND_c_972_n 0.00628107f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_196 N_GATE_c_185_n N_VGND_c_972_n 0.0050896f $X=1.265 $Y=0.88 $X2=0 $Y2=0
cc_197 N_A_249_70#_c_222_n N_A_41_464#_M1003_g 0.0109574f $X=2.195 $Y=1.83 $X2=0
+ $Y2=0
cc_198 N_A_249_70#_c_223_n N_A_41_464#_M1003_g 0.0159908f $X=2.43 $Y=0.765 $X2=0
+ $Y2=0
cc_199 N_A_249_70#_c_225_n N_A_41_464#_M1003_g 0.00657043f $X=3.475 $Y=1.59
+ $X2=0 $Y2=0
cc_200 N_A_249_70#_c_229_n N_A_41_464#_M1003_g 0.0116933f $X=3.655 $Y=0.79 $X2=0
+ $Y2=0
cc_201 N_A_249_70#_c_232_n N_A_41_464#_M1003_g 0.00112723f $X=2.41 $Y=0.79 $X2=0
+ $Y2=0
cc_202 N_A_249_70#_c_235_n N_A_41_464#_M1003_g 0.0219164f $X=2.43 $Y=0.93 $X2=0
+ $Y2=0
cc_203 N_A_249_70#_M1001_g N_A_41_464#_M1002_g 0.00900704f $X=2.195 $Y=2.685
+ $X2=0 $Y2=0
cc_204 N_A_249_70#_c_242_n N_A_41_464#_c_372_n 0.014474f $X=2.195 $Y=1.995 $X2=0
+ $Y2=0
cc_205 N_A_249_70#_M1001_g N_A_41_464#_c_373_n 0.014474f $X=2.195 $Y=2.685 $X2=0
+ $Y2=0
cc_206 N_A_249_70#_M1007_g N_A_41_464#_c_373_n 0.0650737f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_207 N_A_249_70#_c_241_n N_A_41_464#_c_376_n 6.63789e-19 $X=2.12 $Y=1.995
+ $X2=0 $Y2=0
cc_208 N_A_249_70#_c_228_n N_A_41_464#_c_376_n 0.00710042f $X=1.63 $Y=1.995
+ $X2=0 $Y2=0
cc_209 N_A_249_70#_c_228_n N_A_41_464#_c_377_n 0.0110514f $X=1.63 $Y=1.995 $X2=0
+ $Y2=0
cc_210 N_A_249_70#_c_244_n N_A_41_464#_c_377_n 0.0246186f $X=1.635 $Y=2.57 $X2=0
+ $Y2=0
cc_211 N_A_249_70#_M1014_d N_A_41_464#_c_378_n 0.00467848f $X=1.245 $Y=2.32
+ $X2=0 $Y2=0
cc_212 N_A_249_70#_M1001_g N_A_41_464#_c_378_n 0.0154258f $X=2.195 $Y=2.685
+ $X2=0 $Y2=0
cc_213 N_A_249_70#_c_244_n N_A_41_464#_c_378_n 0.0269181f $X=1.635 $Y=2.57 $X2=0
+ $Y2=0
cc_214 N_A_249_70#_M1001_g N_A_41_464#_c_380_n 0.0224701f $X=2.195 $Y=2.685
+ $X2=0 $Y2=0
cc_215 N_A_249_70#_c_222_n N_A_41_464#_c_369_n 0.00596736f $X=2.195 $Y=1.83
+ $X2=0 $Y2=0
cc_216 N_A_249_70#_M1001_g N_A_41_464#_c_369_n 2.71045e-19 $X=2.195 $Y=2.685
+ $X2=0 $Y2=0
cc_217 N_A_249_70#_c_242_n N_A_41_464#_c_369_n 0.00837673f $X=2.195 $Y=1.995
+ $X2=0 $Y2=0
cc_218 N_A_249_70#_c_222_n N_A_41_464#_c_370_n 0.014474f $X=2.195 $Y=1.83 $X2=0
+ $Y2=0
cc_219 N_A_249_70#_M1007_g N_A_41_464#_c_370_n 0.00657043f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_220 N_A_249_70#_c_235_n N_A_41_464#_c_370_n 0.00213794f $X=2.43 $Y=0.93 $X2=0
+ $Y2=0
cc_221 N_A_249_70#_M1009_g N_A_371_473#_M1005_g 0.0208141f $X=3.76 $Y=0.445
+ $X2=0 $Y2=0
cc_222 N_A_249_70#_c_229_n N_A_371_473#_M1005_g 0.0121724f $X=3.655 $Y=0.79
+ $X2=0 $Y2=0
cc_223 N_A_249_70#_c_230_n N_A_371_473#_M1005_g 0.00171438f $X=3.74 $Y=1.175
+ $X2=0 $Y2=0
cc_224 N_A_249_70#_M1007_g N_A_371_473#_M1017_g 0.0139144f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_225 N_A_249_70#_c_223_n N_A_371_473#_c_466_n 0.00432882f $X=2.43 $Y=0.765
+ $X2=0 $Y2=0
cc_226 N_A_249_70#_c_228_n N_A_371_473#_c_466_n 0.039839f $X=1.63 $Y=1.995 $X2=0
+ $Y2=0
cc_227 N_A_249_70#_c_231_n N_A_371_473#_c_466_n 0.0110884f $X=1.635 $Y=0.5 $X2=0
+ $Y2=0
cc_228 N_A_249_70#_c_232_n N_A_371_473#_c_466_n 0.0243998f $X=2.41 $Y=0.79 $X2=0
+ $Y2=0
cc_229 N_A_249_70#_c_235_n N_A_371_473#_c_466_n 0.0103593f $X=2.43 $Y=0.93 $X2=0
+ $Y2=0
cc_230 N_A_249_70#_c_222_n N_A_371_473#_c_467_n 0.0113993f $X=2.195 $Y=1.83
+ $X2=0 $Y2=0
cc_231 N_A_249_70#_M1001_g N_A_371_473#_c_467_n 0.00476424f $X=2.195 $Y=2.685
+ $X2=0 $Y2=0
cc_232 N_A_249_70#_c_241_n N_A_371_473#_c_467_n 0.023067f $X=2.12 $Y=1.995 $X2=0
+ $Y2=0
cc_233 N_A_249_70#_c_228_n N_A_371_473#_c_467_n 0.0765617f $X=1.63 $Y=1.995
+ $X2=0 $Y2=0
cc_234 N_A_249_70#_c_244_n N_A_371_473#_c_467_n 0.0260803f $X=1.635 $Y=2.57
+ $X2=0 $Y2=0
cc_235 N_A_249_70#_c_222_n N_A_371_473#_c_468_n 0.0175079f $X=2.195 $Y=1.83
+ $X2=0 $Y2=0
cc_236 N_A_249_70#_c_241_n N_A_371_473#_c_468_n 0.00107415f $X=2.12 $Y=1.995
+ $X2=0 $Y2=0
cc_237 N_A_249_70#_c_229_n N_A_371_473#_c_468_n 0.0189809f $X=3.655 $Y=0.79
+ $X2=0 $Y2=0
cc_238 N_A_249_70#_c_232_n N_A_371_473#_c_468_n 0.0246232f $X=2.41 $Y=0.79 $X2=0
+ $Y2=0
cc_239 N_A_249_70#_c_235_n N_A_371_473#_c_468_n 0.00656366f $X=2.43 $Y=0.93
+ $X2=0 $Y2=0
cc_240 N_A_249_70#_c_225_n N_A_371_473#_c_469_n 0.0082585f $X=3.475 $Y=1.59
+ $X2=0 $Y2=0
cc_241 N_A_249_70#_c_227_n N_A_371_473#_c_469_n 0.00244022f $X=3.85 $Y=1.515
+ $X2=0 $Y2=0
cc_242 N_A_249_70#_c_233_n N_A_371_473#_c_469_n 0.00261617f $X=3.85 $Y=1.34
+ $X2=0 $Y2=0
cc_243 N_A_249_70#_M1007_g N_A_371_473#_c_477_n 0.0111299f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_244 N_A_249_70#_M1007_g N_A_371_473#_c_479_n 0.00107963f $X=3.4 $Y=2.685
+ $X2=0 $Y2=0
cc_245 N_A_249_70#_c_223_n N_A_371_473#_c_470_n 0.00243824f $X=2.43 $Y=0.765
+ $X2=0 $Y2=0
cc_246 N_A_249_70#_c_231_n N_A_371_473#_c_470_n 0.0180763f $X=1.635 $Y=0.5 $X2=0
+ $Y2=0
cc_247 N_A_249_70#_c_232_n N_A_371_473#_c_470_n 0.00653721f $X=2.41 $Y=0.79
+ $X2=0 $Y2=0
cc_248 N_A_249_70#_c_235_n N_A_371_473#_c_470_n 0.00430008f $X=2.43 $Y=0.93
+ $X2=0 $Y2=0
cc_249 N_A_249_70#_c_228_n N_A_371_473#_c_471_n 0.0144138f $X=1.63 $Y=1.995
+ $X2=0 $Y2=0
cc_250 N_A_249_70#_c_225_n N_A_371_473#_c_472_n 0.00136982f $X=3.475 $Y=1.59
+ $X2=0 $Y2=0
cc_251 N_A_249_70#_c_229_n N_A_371_473#_c_472_n 0.0328032f $X=3.655 $Y=0.79
+ $X2=0 $Y2=0
cc_252 N_A_249_70#_c_230_n N_A_371_473#_c_472_n 0.00940213f $X=3.74 $Y=1.175
+ $X2=0 $Y2=0
cc_253 N_A_249_70#_c_233_n N_A_371_473#_c_472_n 0.015553f $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_254 N_A_249_70#_c_234_n N_A_371_473#_c_472_n 5.8211e-19 $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_255 N_A_249_70#_c_225_n N_A_371_473#_c_473_n 0.00990992f $X=3.475 $Y=1.59
+ $X2=0 $Y2=0
cc_256 N_A_249_70#_M1009_g N_A_371_473#_c_473_n 0.0211732f $X=3.76 $Y=0.445
+ $X2=0 $Y2=0
cc_257 N_A_249_70#_c_229_n N_A_371_473#_c_473_n 0.0043813f $X=3.655 $Y=0.79
+ $X2=0 $Y2=0
cc_258 N_A_249_70#_c_230_n N_A_371_473#_c_473_n 0.00179762f $X=3.74 $Y=1.175
+ $X2=0 $Y2=0
cc_259 N_A_249_70#_c_233_n N_A_371_473#_c_473_n 4.37106e-19 $X=3.85 $Y=1.34
+ $X2=0 $Y2=0
cc_260 N_A_249_70#_M1007_g N_A_371_473#_c_480_n 0.0205563f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_261 N_A_249_70#_c_224_n N_A_371_473#_c_480_n 0.0207526f $X=3.685 $Y=1.59
+ $X2=0 $Y2=0
cc_262 N_A_249_70#_M1007_g N_A_371_473#_c_481_n 3.06081e-19 $X=3.4 $Y=2.685
+ $X2=0 $Y2=0
cc_263 N_A_249_70#_c_224_n N_A_371_473#_c_481_n 2.91744e-19 $X=3.685 $Y=1.59
+ $X2=0 $Y2=0
cc_264 N_A_249_70#_M1009_g N_A_809_21#_c_581_n 0.0507147f $X=3.76 $Y=0.445 $X2=0
+ $Y2=0
cc_265 N_A_249_70#_M1009_g N_A_809_21#_c_588_n 0.00807357f $X=3.76 $Y=0.445
+ $X2=0 $Y2=0
cc_266 N_A_249_70#_c_230_n N_A_809_21#_c_588_n 0.00147717f $X=3.74 $Y=1.175
+ $X2=0 $Y2=0
cc_267 N_A_249_70#_c_233_n N_A_809_21#_c_588_n 9.7532e-19 $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_268 N_A_249_70#_c_234_n N_A_809_21#_c_588_n 0.0302003f $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_269 N_A_249_70#_M1007_g N_A_659_47#_c_716_n 0.0147958f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_270 N_A_249_70#_M1009_g N_A_659_47#_c_720_n 0.00889484f $X=3.76 $Y=0.445
+ $X2=0 $Y2=0
cc_271 N_A_249_70#_c_229_n N_A_659_47#_c_720_n 0.0301062f $X=3.655 $Y=0.79 $X2=0
+ $Y2=0
cc_272 N_A_249_70#_c_233_n N_A_659_47#_c_720_n 0.00364504f $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_273 N_A_249_70#_c_234_n N_A_659_47#_c_720_n 0.00263277f $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_274 N_A_249_70#_c_224_n N_A_659_47#_c_707_n 0.0179222f $X=3.685 $Y=1.59 $X2=0
+ $Y2=0
cc_275 N_A_249_70#_c_233_n N_A_659_47#_c_707_n 0.0253088f $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_276 N_A_249_70#_M1007_g N_A_659_47#_c_726_n 0.0045686f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_277 N_A_249_70#_c_224_n N_A_659_47#_c_726_n 0.00251808f $X=3.685 $Y=1.59
+ $X2=0 $Y2=0
cc_278 N_A_249_70#_c_225_n N_A_659_47#_c_726_n 0.00220002f $X=3.475 $Y=1.59
+ $X2=0 $Y2=0
cc_279 N_A_249_70#_M1009_g N_A_659_47#_c_708_n 0.00138212f $X=3.76 $Y=0.445
+ $X2=0 $Y2=0
cc_280 N_A_249_70#_c_229_n N_A_659_47#_c_708_n 0.00149399f $X=3.655 $Y=0.79
+ $X2=0 $Y2=0
cc_281 N_A_249_70#_M1009_g N_A_659_47#_c_710_n 9.78418e-19 $X=3.76 $Y=0.445
+ $X2=0 $Y2=0
cc_282 N_A_249_70#_c_229_n N_A_659_47#_c_710_n 0.0128337f $X=3.655 $Y=0.79 $X2=0
+ $Y2=0
cc_283 N_A_249_70#_c_230_n N_A_659_47#_c_710_n 0.00151728f $X=3.74 $Y=1.175
+ $X2=0 $Y2=0
cc_284 N_A_249_70#_c_233_n N_A_659_47#_c_710_n 5.64806e-19 $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_285 N_A_249_70#_c_234_n N_A_659_47#_c_710_n 2.34038e-19 $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_286 N_A_249_70#_M1007_g N_A_659_47#_c_736_n 0.00801981f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_287 N_A_249_70#_c_233_n N_A_659_47#_c_712_n 0.00857094f $X=3.85 $Y=1.34 $X2=0
+ $Y2=0
cc_288 N_A_249_70#_M1001_g N_VPWR_c_860_n 0.00315744f $X=2.195 $Y=2.685 $X2=0
+ $Y2=0
cc_289 N_A_249_70#_M1001_g N_VPWR_c_864_n 0.00302479f $X=2.195 $Y=2.685 $X2=0
+ $Y2=0
cc_290 N_A_249_70#_M1007_g N_VPWR_c_865_n 0.00302501f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_291 N_A_249_70#_M1001_g N_VPWR_c_858_n 0.00512844f $X=2.195 $Y=2.685 $X2=0
+ $Y2=0
cc_292 N_A_249_70#_M1007_g N_VPWR_c_858_n 0.00478661f $X=3.4 $Y=2.685 $X2=0
+ $Y2=0
cc_293 N_A_249_70#_c_231_n N_VGND_c_963_n 0.0140296f $X=1.635 $Y=0.5 $X2=0 $Y2=0
cc_294 N_A_249_70#_c_223_n N_VGND_c_964_n 0.00303181f $X=2.43 $Y=0.765 $X2=0
+ $Y2=0
cc_295 N_A_249_70#_c_229_n N_VGND_c_964_n 0.0157811f $X=3.655 $Y=0.79 $X2=0
+ $Y2=0
cc_296 N_A_249_70#_c_232_n N_VGND_c_964_n 0.00218915f $X=2.41 $Y=0.79 $X2=0
+ $Y2=0
cc_297 N_A_249_70#_c_235_n N_VGND_c_964_n 2.05862e-19 $X=2.43 $Y=0.93 $X2=0
+ $Y2=0
cc_298 N_A_249_70#_c_223_n N_VGND_c_969_n 0.004324f $X=2.43 $Y=0.765 $X2=0 $Y2=0
cc_299 N_A_249_70#_c_231_n N_VGND_c_969_n 0.0231285f $X=1.635 $Y=0.5 $X2=0 $Y2=0
cc_300 N_A_249_70#_c_232_n N_VGND_c_969_n 0.00252135f $X=2.41 $Y=0.79 $X2=0
+ $Y2=0
cc_301 N_A_249_70#_M1009_g N_VGND_c_970_n 0.00370116f $X=3.76 $Y=0.445 $X2=0
+ $Y2=0
cc_302 N_A_249_70#_c_229_n N_VGND_c_970_n 0.00849173f $X=3.655 $Y=0.79 $X2=0
+ $Y2=0
cc_303 N_A_249_70#_c_223_n N_VGND_c_972_n 0.00710831f $X=2.43 $Y=0.765 $X2=0
+ $Y2=0
cc_304 N_A_249_70#_M1009_g N_VGND_c_972_n 0.00547618f $X=3.76 $Y=0.445 $X2=0
+ $Y2=0
cc_305 N_A_249_70#_c_229_n N_VGND_c_972_n 0.0154797f $X=3.655 $Y=0.79 $X2=0
+ $Y2=0
cc_306 N_A_249_70#_c_231_n N_VGND_c_972_n 0.0183373f $X=1.635 $Y=0.5 $X2=0 $Y2=0
cc_307 N_A_249_70#_c_232_n N_VGND_c_972_n 0.00435665f $X=2.41 $Y=0.79 $X2=0
+ $Y2=0
cc_308 N_A_41_464#_c_378_n N_A_371_473#_M1001_s 0.00380539f $X=2.25 $Y=2.99
+ $X2=0 $Y2=0
cc_309 N_A_41_464#_M1003_g N_A_371_473#_M1005_g 0.0759412f $X=2.86 $Y=0.445
+ $X2=0 $Y2=0
cc_310 N_A_41_464#_c_372_n N_A_371_473#_c_467_n 2.08622e-19 $X=2.797 $Y=2.055
+ $X2=0 $Y2=0
cc_311 N_A_41_464#_c_378_n N_A_371_473#_c_467_n 0.0127109f $X=2.25 $Y=2.99 $X2=0
+ $Y2=0
cc_312 N_A_41_464#_c_369_n N_A_371_473#_c_467_n 0.0752472f $X=2.645 $Y=1.7 $X2=0
+ $Y2=0
cc_313 N_A_41_464#_M1003_g N_A_371_473#_c_468_n 0.0164944f $X=2.86 $Y=0.445
+ $X2=0 $Y2=0
cc_314 N_A_41_464#_c_373_n N_A_371_473#_c_468_n 0.00119948f $X=2.797 $Y=2.205
+ $X2=0 $Y2=0
cc_315 N_A_41_464#_c_369_n N_A_371_473#_c_468_n 0.0452336f $X=2.645 $Y=1.7 $X2=0
+ $Y2=0
cc_316 N_A_41_464#_c_370_n N_A_371_473#_c_468_n 0.0018026f $X=2.645 $Y=1.7 $X2=0
+ $Y2=0
cc_317 N_A_41_464#_M1003_g N_A_371_473#_c_469_n 0.011558f $X=2.86 $Y=0.445 $X2=0
+ $Y2=0
cc_318 N_A_41_464#_M1002_g N_A_371_473#_c_469_n 0.0152599f $X=3.04 $Y=2.685
+ $X2=0 $Y2=0
cc_319 N_A_41_464#_c_373_n N_A_371_473#_c_469_n 0.00767537f $X=2.797 $Y=2.205
+ $X2=0 $Y2=0
cc_320 N_A_41_464#_c_380_n N_A_371_473#_c_469_n 0.00485367f $X=2.335 $Y=2.905
+ $X2=0 $Y2=0
cc_321 N_A_41_464#_c_369_n N_A_371_473#_c_469_n 0.0474674f $X=2.645 $Y=1.7 $X2=0
+ $Y2=0
cc_322 N_A_41_464#_M1002_g N_A_371_473#_c_478_n 0.00524418f $X=3.04 $Y=2.685
+ $X2=0 $Y2=0
cc_323 N_A_41_464#_M1003_g N_A_371_473#_c_472_n 0.00100252f $X=2.86 $Y=0.445
+ $X2=0 $Y2=0
cc_324 N_A_41_464#_c_373_n N_A_659_47#_c_716_n 3.94505e-19 $X=2.797 $Y=2.205
+ $X2=0 $Y2=0
cc_325 N_A_41_464#_M1002_g N_A_659_47#_c_736_n 3.70502e-19 $X=3.04 $Y=2.685
+ $X2=0 $Y2=0
cc_326 N_A_41_464#_c_377_n N_VPWR_M1015_d 0.00533256f $X=1.1 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_327 N_A_41_464#_c_379_n N_VPWR_M1015_d 5.22721e-19 $X=1.185 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_328 N_A_41_464#_c_378_n N_VPWR_M1001_d 9.99249e-19 $X=2.25 $Y=2.99 $X2=0
+ $Y2=0
cc_329 N_A_41_464#_c_380_n N_VPWR_M1001_d 0.00517437f $X=2.335 $Y=2.905 $X2=0
+ $Y2=0
cc_330 N_A_41_464#_c_375_n N_VPWR_c_859_n 0.00267962f $X=0.33 $Y=2.465 $X2=0
+ $Y2=0
cc_331 N_A_41_464#_c_376_n N_VPWR_c_859_n 0.0158786f $X=1.015 $Y=2.045 $X2=0
+ $Y2=0
cc_332 N_A_41_464#_c_377_n N_VPWR_c_859_n 0.0443297f $X=1.1 $Y=2.905 $X2=0 $Y2=0
cc_333 N_A_41_464#_c_379_n N_VPWR_c_859_n 0.0142942f $X=1.185 $Y=2.99 $X2=0
+ $Y2=0
cc_334 N_A_41_464#_M1002_g N_VPWR_c_860_n 0.0085467f $X=3.04 $Y=2.685 $X2=0
+ $Y2=0
cc_335 N_A_41_464#_c_373_n N_VPWR_c_860_n 0.00657084f $X=2.797 $Y=2.205 $X2=0
+ $Y2=0
cc_336 N_A_41_464#_c_378_n N_VPWR_c_860_n 0.014341f $X=2.25 $Y=2.99 $X2=0 $Y2=0
cc_337 N_A_41_464#_c_380_n N_VPWR_c_860_n 0.0416354f $X=2.335 $Y=2.905 $X2=0
+ $Y2=0
cc_338 N_A_41_464#_c_369_n N_VPWR_c_860_n 0.0193502f $X=2.645 $Y=1.7 $X2=0 $Y2=0
cc_339 N_A_41_464#_c_378_n N_VPWR_c_864_n 0.0800837f $X=2.25 $Y=2.99 $X2=0 $Y2=0
cc_340 N_A_41_464#_c_379_n N_VPWR_c_864_n 0.0118704f $X=1.185 $Y=2.99 $X2=0
+ $Y2=0
cc_341 N_A_41_464#_M1002_g N_VPWR_c_865_n 0.00335204f $X=3.04 $Y=2.685 $X2=0
+ $Y2=0
cc_342 N_A_41_464#_M1002_g N_VPWR_c_858_n 0.00549498f $X=3.04 $Y=2.685 $X2=0
+ $Y2=0
cc_343 N_A_41_464#_c_375_n N_VPWR_c_858_n 0.0106368f $X=0.33 $Y=2.465 $X2=0
+ $Y2=0
cc_344 N_A_41_464#_c_378_n N_VPWR_c_858_n 0.0456831f $X=2.25 $Y=2.99 $X2=0 $Y2=0
cc_345 N_A_41_464#_c_379_n N_VPWR_c_858_n 0.0061974f $X=1.185 $Y=2.99 $X2=0
+ $Y2=0
cc_346 N_A_41_464#_c_375_n N_VPWR_c_868_n 0.0128508f $X=0.33 $Y=2.465 $X2=0
+ $Y2=0
cc_347 N_A_41_464#_M1003_g N_VGND_c_964_n 0.0100885f $X=2.86 $Y=0.445 $X2=0
+ $Y2=0
cc_348 N_A_41_464#_M1003_g N_VGND_c_970_n 0.00361815f $X=2.86 $Y=0.445 $X2=0
+ $Y2=0
cc_349 N_A_41_464#_M1003_g N_VGND_c_972_n 0.00416812f $X=2.86 $Y=0.445 $X2=0
+ $Y2=0
cc_350 N_A_41_464#_c_368_n N_VGND_c_972_n 0.0103695f $X=0.37 $Y=0.555 $X2=0
+ $Y2=0
cc_351 N_A_41_464#_c_368_n N_VGND_c_973_n 0.0108128f $X=0.37 $Y=0.555 $X2=0
+ $Y2=0
cc_352 N_A_371_473#_M1017_g N_A_809_21#_M1008_g 0.0353053f $X=3.925 $Y=2.575
+ $X2=0 $Y2=0
cc_353 N_A_371_473#_c_479_n N_A_809_21#_M1008_g 0.0050849f $X=3.965 $Y=2.905
+ $X2=0 $Y2=0
cc_354 N_A_371_473#_c_480_n N_A_809_21#_c_591_n 3.01893e-19 $X=3.855 $Y=2.04
+ $X2=0 $Y2=0
cc_355 N_A_371_473#_c_481_n N_A_809_21#_c_591_n 0.0209658f $X=3.965 $Y=2.075
+ $X2=0 $Y2=0
cc_356 N_A_371_473#_c_480_n N_A_809_21#_c_592_n 0.0220907f $X=3.855 $Y=2.04
+ $X2=0 $Y2=0
cc_357 N_A_371_473#_c_481_n N_A_809_21#_c_592_n 8.74212e-19 $X=3.965 $Y=2.075
+ $X2=0 $Y2=0
cc_358 N_A_371_473#_c_477_n N_A_659_47#_M1007_d 0.00339864f $X=3.88 $Y=2.99
+ $X2=0 $Y2=0
cc_359 N_A_371_473#_M1017_g N_A_659_47#_c_716_n 0.00113749f $X=3.925 $Y=2.575
+ $X2=0 $Y2=0
cc_360 N_A_371_473#_c_469_n N_A_659_47#_c_716_n 0.0416516f $X=3.075 $Y=2.905
+ $X2=0 $Y2=0
cc_361 N_A_371_473#_c_479_n N_A_659_47#_c_716_n 0.00710387f $X=3.965 $Y=2.905
+ $X2=0 $Y2=0
cc_362 N_A_371_473#_c_480_n N_A_659_47#_c_716_n 0.00220609f $X=3.855 $Y=2.04
+ $X2=0 $Y2=0
cc_363 N_A_371_473#_c_481_n N_A_659_47#_c_716_n 0.0187835f $X=3.965 $Y=2.075
+ $X2=0 $Y2=0
cc_364 N_A_371_473#_M1005_g N_A_659_47#_c_720_n 0.00339307f $X=3.22 $Y=0.445
+ $X2=0 $Y2=0
cc_365 N_A_371_473#_c_480_n N_A_659_47#_c_707_n 0.00219961f $X=3.855 $Y=2.04
+ $X2=0 $Y2=0
cc_366 N_A_371_473#_c_481_n N_A_659_47#_c_707_n 0.0266895f $X=3.965 $Y=2.075
+ $X2=0 $Y2=0
cc_367 N_A_371_473#_c_469_n N_A_659_47#_c_726_n 0.0129671f $X=3.075 $Y=2.905
+ $X2=0 $Y2=0
cc_368 N_A_371_473#_c_472_n N_A_659_47#_c_726_n 0.00874882f $X=3.075 $Y=1.205
+ $X2=0 $Y2=0
cc_369 N_A_371_473#_M1017_g N_A_659_47#_c_736_n 0.00241057f $X=3.925 $Y=2.575
+ $X2=0 $Y2=0
cc_370 N_A_371_473#_c_477_n N_A_659_47#_c_736_n 0.021054f $X=3.88 $Y=2.99 $X2=0
+ $Y2=0
cc_371 N_A_371_473#_c_479_n N_A_659_47#_c_736_n 0.0235002f $X=3.965 $Y=2.905
+ $X2=0 $Y2=0
cc_372 N_A_371_473#_c_480_n N_A_659_47#_c_736_n 2.23801e-19 $X=3.855 $Y=2.04
+ $X2=0 $Y2=0
cc_373 N_A_371_473#_c_481_n N_A_659_47#_c_736_n 6.73161e-19 $X=3.965 $Y=2.075
+ $X2=0 $Y2=0
cc_374 N_A_371_473#_c_469_n N_VPWR_c_860_n 0.0402512f $X=3.075 $Y=2.905 $X2=0
+ $Y2=0
cc_375 N_A_371_473#_c_478_n N_VPWR_c_860_n 0.0137471f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_376 N_A_371_473#_M1017_g N_VPWR_c_865_n 6.53345e-19 $X=3.925 $Y=2.575 $X2=0
+ $Y2=0
cc_377 N_A_371_473#_c_477_n N_VPWR_c_865_n 0.058073f $X=3.88 $Y=2.99 $X2=0 $Y2=0
cc_378 N_A_371_473#_c_478_n N_VPWR_c_865_n 0.0116785f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_379 N_A_371_473#_c_477_n N_VPWR_c_858_n 0.032989f $X=3.88 $Y=2.99 $X2=0 $Y2=0
cc_380 N_A_371_473#_c_478_n N_VPWR_c_858_n 0.00602728f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_381 N_A_371_473#_M1017_g N_VPWR_c_870_n 5.10473e-19 $X=3.925 $Y=2.575 $X2=0
+ $Y2=0
cc_382 N_A_371_473#_c_477_n N_VPWR_c_870_n 0.0103458f $X=3.88 $Y=2.99 $X2=0
+ $Y2=0
cc_383 N_A_371_473#_c_479_n N_VPWR_c_870_n 0.01572f $X=3.965 $Y=2.905 $X2=0
+ $Y2=0
cc_384 N_A_371_473#_c_477_n A_623_473# 0.00366293f $X=3.88 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_385 N_A_371_473#_M1005_g N_VGND_c_964_n 0.0021589f $X=3.22 $Y=0.445 $X2=0
+ $Y2=0
cc_386 N_A_371_473#_c_470_n N_VGND_c_969_n 0.0289237f $X=2.195 $Y=0.42 $X2=0
+ $Y2=0
cc_387 N_A_371_473#_M1005_g N_VGND_c_970_n 0.00435108f $X=3.22 $Y=0.445 $X2=0
+ $Y2=0
cc_388 N_A_371_473#_M1012_s N_VGND_c_972_n 0.00228716f $X=2.07 $Y=0.235 $X2=0
+ $Y2=0
cc_389 N_A_371_473#_M1005_g N_VGND_c_972_n 0.00631645f $X=3.22 $Y=0.445 $X2=0
+ $Y2=0
cc_390 N_A_371_473#_c_470_n N_VGND_c_972_n 0.0175819f $X=2.195 $Y=0.42 $X2=0
+ $Y2=0
cc_391 N_A_809_21#_c_584_n N_A_659_47#_M1006_g 0.0139692f $X=4.99 $Y=0.51 $X2=0
+ $Y2=0
cc_392 N_A_809_21#_c_585_n N_A_659_47#_M1006_g 0.00485053f $X=5.17 $Y=1.945
+ $X2=0 $Y2=0
cc_393 N_A_809_21#_c_611_p N_A_659_47#_M1006_g 0.00315522f $X=5.065 $Y=1.165
+ $X2=0 $Y2=0
cc_394 N_A_809_21#_c_592_n N_A_659_47#_M1004_g 0.0050896f $X=4.395 $Y=2.04 $X2=0
+ $Y2=0
cc_395 N_A_809_21#_c_585_n N_A_659_47#_M1004_g 0.00839993f $X=5.17 $Y=1.945
+ $X2=0 $Y2=0
cc_396 N_A_809_21#_c_614_p N_A_659_47#_M1004_g 0.0236002f $X=5.405 $Y=2.47 $X2=0
+ $Y2=0
cc_397 N_A_809_21#_c_615_p N_A_659_47#_M1004_g 0.00871612f $X=5.42 $Y=2.91 $X2=0
+ $Y2=0
cc_398 N_A_809_21#_c_591_n N_A_659_47#_c_705_n 0.00714735f $X=5.085 $Y=2.075
+ $X2=0 $Y2=0
cc_399 N_A_809_21#_c_585_n N_A_659_47#_c_705_n 0.00796982f $X=5.17 $Y=1.945
+ $X2=0 $Y2=0
cc_400 N_A_809_21#_c_611_p N_A_659_47#_c_705_n 0.00760991f $X=5.065 $Y=1.165
+ $X2=0 $Y2=0
cc_401 N_A_809_21#_c_588_n N_A_659_47#_c_705_n 0.0134163f $X=4.395 $Y=1.875
+ $X2=0 $Y2=0
cc_402 N_A_809_21#_c_585_n N_A_659_47#_c_706_n 0.0055112f $X=5.17 $Y=1.945 $X2=0
+ $Y2=0
cc_403 N_A_809_21#_c_581_n N_A_659_47#_c_720_n 0.00728916f $X=4.12 $Y=0.765
+ $X2=0 $Y2=0
cc_404 N_A_809_21#_c_583_n N_A_659_47#_c_707_n 0.00434948f $X=4.305 $Y=0.84
+ $X2=0 $Y2=0
cc_405 N_A_809_21#_c_591_n N_A_659_47#_c_707_n 0.0219496f $X=5.085 $Y=2.075
+ $X2=0 $Y2=0
cc_406 N_A_809_21#_c_592_n N_A_659_47#_c_707_n 0.00381742f $X=4.395 $Y=2.04
+ $X2=0 $Y2=0
cc_407 N_A_809_21#_c_588_n N_A_659_47#_c_707_n 0.0165834f $X=4.395 $Y=1.875
+ $X2=0 $Y2=0
cc_408 N_A_809_21#_c_581_n N_A_659_47#_c_708_n 0.00905385f $X=4.12 $Y=0.765
+ $X2=0 $Y2=0
cc_409 N_A_809_21#_c_581_n N_A_659_47#_c_709_n 0.00140825f $X=4.12 $Y=0.765
+ $X2=0 $Y2=0
cc_410 N_A_809_21#_c_583_n N_A_659_47#_c_709_n 0.0164534f $X=4.305 $Y=0.84 $X2=0
+ $Y2=0
cc_411 N_A_809_21#_c_584_n N_A_659_47#_c_709_n 0.0149588f $X=4.99 $Y=0.51 $X2=0
+ $Y2=0
cc_412 N_A_809_21#_c_581_n N_A_659_47#_c_710_n 5.74535e-19 $X=4.12 $Y=0.765
+ $X2=0 $Y2=0
cc_413 N_A_809_21#_c_583_n N_A_659_47#_c_710_n 0.00743428f $X=4.305 $Y=0.84
+ $X2=0 $Y2=0
cc_414 N_A_809_21#_c_591_n N_A_659_47#_c_711_n 0.0320916f $X=5.085 $Y=2.075
+ $X2=0 $Y2=0
cc_415 N_A_809_21#_c_592_n N_A_659_47#_c_711_n 6.08687e-19 $X=4.395 $Y=2.04
+ $X2=0 $Y2=0
cc_416 N_A_809_21#_c_585_n N_A_659_47#_c_711_n 0.0326551f $X=5.17 $Y=1.945 $X2=0
+ $Y2=0
cc_417 N_A_809_21#_c_611_p N_A_659_47#_c_711_n 0.00321828f $X=5.065 $Y=1.165
+ $X2=0 $Y2=0
cc_418 N_A_809_21#_c_588_n N_A_659_47#_c_711_n 0.0100356f $X=4.395 $Y=1.875
+ $X2=0 $Y2=0
cc_419 N_A_809_21#_c_583_n N_A_659_47#_c_712_n 0.0093992f $X=4.305 $Y=0.84 $X2=0
+ $Y2=0
cc_420 N_A_809_21#_c_584_n N_A_659_47#_c_712_n 0.0211453f $X=4.99 $Y=0.51 $X2=0
+ $Y2=0
cc_421 N_A_809_21#_c_585_n N_A_659_47#_c_712_n 0.00643373f $X=5.17 $Y=1.945
+ $X2=0 $Y2=0
cc_422 N_A_809_21#_M1011_g N_RESET_B_M1019_g 0.0180006f $X=6.105 $Y=0.785 $X2=0
+ $Y2=0
cc_423 N_A_809_21#_c_584_n N_RESET_B_M1019_g 7.06311e-19 $X=4.99 $Y=0.51 $X2=0
+ $Y2=0
cc_424 N_A_809_21#_M1018_g N_RESET_B_M1016_g 0.0371176f $X=6.14 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_809_21#_c_585_n N_RESET_B_M1016_g 2.66039e-19 $X=5.17 $Y=1.945 $X2=0
+ $Y2=0
cc_426 N_A_809_21#_c_614_p N_RESET_B_M1016_g 5.48082e-19 $X=5.405 $Y=2.47 $X2=0
+ $Y2=0
cc_427 N_A_809_21#_c_645_p N_RESET_B_M1016_g 0.0103985f $X=5.92 $Y=2.385 $X2=0
+ $Y2=0
cc_428 N_A_809_21#_c_594_n N_RESET_B_M1016_g 0.00319994f $X=6.005 $Y=2.3 $X2=0
+ $Y2=0
cc_429 N_A_809_21#_M1011_g RESET_B 0.00107235f $X=6.105 $Y=0.785 $X2=0 $Y2=0
cc_430 N_A_809_21#_c_584_n RESET_B 0.0396969f $X=4.99 $Y=0.51 $X2=0 $Y2=0
cc_431 N_A_809_21#_c_611_p RESET_B 0.0396969f $X=5.065 $Y=1.165 $X2=0 $Y2=0
cc_432 N_A_809_21#_c_586_n RESET_B 0.0247282f $X=6.195 $Y=1.505 $X2=0 $Y2=0
cc_433 N_A_809_21#_c_587_n RESET_B 2.89063e-19 $X=6.195 $Y=1.505 $X2=0 $Y2=0
cc_434 N_A_809_21#_M1018_g N_RESET_B_c_813_n 2.26231e-19 $X=6.14 $Y=2.465 $X2=0
+ $Y2=0
cc_435 N_A_809_21#_c_645_p N_RESET_B_c_813_n 0.00159663f $X=5.92 $Y=2.385 $X2=0
+ $Y2=0
cc_436 N_A_809_21#_c_611_p N_RESET_B_c_813_n 7.06311e-19 $X=5.065 $Y=1.165 $X2=0
+ $Y2=0
cc_437 N_A_809_21#_c_586_n N_RESET_B_c_813_n 0.00217544f $X=6.195 $Y=1.505 $X2=0
+ $Y2=0
cc_438 N_A_809_21#_c_587_n N_RESET_B_c_813_n 0.0201445f $X=6.195 $Y=1.505 $X2=0
+ $Y2=0
cc_439 N_A_809_21#_M1004_d N_RESET_B_c_814_n 0.00334483f $X=5.28 $Y=1.835 $X2=0
+ $Y2=0
cc_440 N_A_809_21#_M1018_g N_RESET_B_c_814_n 6.39063e-19 $X=6.14 $Y=2.465 $X2=0
+ $Y2=0
cc_441 N_A_809_21#_c_585_n N_RESET_B_c_814_n 0.0396969f $X=5.17 $Y=1.945 $X2=0
+ $Y2=0
cc_442 N_A_809_21#_c_614_p N_RESET_B_c_814_n 0.0221356f $X=5.405 $Y=2.47 $X2=0
+ $Y2=0
cc_443 N_A_809_21#_c_645_p N_RESET_B_c_814_n 0.0113922f $X=5.92 $Y=2.385 $X2=0
+ $Y2=0
cc_444 N_A_809_21#_c_594_n N_RESET_B_c_814_n 0.0227231f $X=6.005 $Y=2.3 $X2=0
+ $Y2=0
cc_445 N_A_809_21#_c_591_n N_VPWR_M1008_d 0.00701689f $X=5.085 $Y=2.075 $X2=0
+ $Y2=0
cc_446 N_A_809_21#_c_645_p N_VPWR_M1016_d 0.00723121f $X=5.92 $Y=2.385 $X2=0
+ $Y2=0
cc_447 N_A_809_21#_c_594_n N_VPWR_M1016_d 0.00496116f $X=6.005 $Y=2.3 $X2=0
+ $Y2=0
cc_448 N_A_809_21#_M1018_g N_VPWR_c_861_n 0.00408238f $X=6.14 $Y=2.465 $X2=0
+ $Y2=0
cc_449 N_A_809_21#_c_645_p N_VPWR_c_861_n 0.0198746f $X=5.92 $Y=2.385 $X2=0
+ $Y2=0
cc_450 N_A_809_21#_c_615_p N_VPWR_c_862_n 0.0171073f $X=5.42 $Y=2.91 $X2=0 $Y2=0
cc_451 N_A_809_21#_M1008_g N_VPWR_c_865_n 0.00382362f $X=4.315 $Y=2.575 $X2=0
+ $Y2=0
cc_452 N_A_809_21#_M1018_g N_VPWR_c_866_n 0.00585385f $X=6.14 $Y=2.465 $X2=0
+ $Y2=0
cc_453 N_A_809_21#_M1004_d N_VPWR_c_858_n 0.00219538f $X=5.28 $Y=1.835 $X2=0
+ $Y2=0
cc_454 N_A_809_21#_M1008_g N_VPWR_c_858_n 0.00410091f $X=4.315 $Y=2.575 $X2=0
+ $Y2=0
cc_455 N_A_809_21#_M1018_g N_VPWR_c_858_n 0.011125f $X=6.14 $Y=2.465 $X2=0 $Y2=0
cc_456 N_A_809_21#_c_614_p N_VPWR_c_858_n 0.00557334f $X=5.405 $Y=2.47 $X2=0
+ $Y2=0
cc_457 N_A_809_21#_c_615_p N_VPWR_c_858_n 0.0114026f $X=5.42 $Y=2.91 $X2=0 $Y2=0
cc_458 N_A_809_21#_c_645_p N_VPWR_c_858_n 0.00684813f $X=5.92 $Y=2.385 $X2=0
+ $Y2=0
cc_459 N_A_809_21#_M1008_g N_VPWR_c_870_n 0.0114814f $X=4.315 $Y=2.575 $X2=0
+ $Y2=0
cc_460 N_A_809_21#_c_591_n N_VPWR_c_870_n 0.0457322f $X=5.085 $Y=2.075 $X2=0
+ $Y2=0
cc_461 N_A_809_21#_c_592_n N_VPWR_c_870_n 0.00372277f $X=4.395 $Y=2.04 $X2=0
+ $Y2=0
cc_462 N_A_809_21#_c_615_p N_VPWR_c_870_n 0.00802427f $X=5.42 $Y=2.91 $X2=0
+ $Y2=0
cc_463 N_A_809_21#_M1011_g N_Q_c_941_n 0.00877915f $X=6.105 $Y=0.785 $X2=0 $Y2=0
cc_464 N_A_809_21#_M1011_g N_Q_c_942_n 0.00259502f $X=6.105 $Y=0.785 $X2=0 $Y2=0
cc_465 N_A_809_21#_c_586_n N_Q_c_942_n 0.00717444f $X=6.195 $Y=1.505 $X2=0 $Y2=0
cc_466 N_A_809_21#_c_587_n N_Q_c_942_n 0.00471609f $X=6.195 $Y=1.505 $X2=0 $Y2=0
cc_467 N_A_809_21#_c_586_n Q 0.00102804f $X=6.195 $Y=1.505 $X2=0 $Y2=0
cc_468 N_A_809_21#_c_587_n Q 0.00279611f $X=6.195 $Y=1.505 $X2=0 $Y2=0
cc_469 N_A_809_21#_M1011_g N_Q_c_943_n 0.00370067f $X=6.105 $Y=0.785 $X2=0 $Y2=0
cc_470 N_A_809_21#_M1018_g N_Q_c_943_n 0.00253293f $X=6.14 $Y=2.465 $X2=0 $Y2=0
cc_471 N_A_809_21#_c_594_n N_Q_c_943_n 0.00532674f $X=6.005 $Y=2.3 $X2=0 $Y2=0
cc_472 N_A_809_21#_c_586_n N_Q_c_943_n 0.0250436f $X=6.195 $Y=1.505 $X2=0 $Y2=0
cc_473 N_A_809_21#_c_587_n N_Q_c_943_n 0.00817336f $X=6.195 $Y=1.505 $X2=0 $Y2=0
cc_474 N_A_809_21#_c_581_n N_VGND_c_965_n 0.0113315f $X=4.12 $Y=0.765 $X2=0
+ $Y2=0
cc_475 N_A_809_21#_c_583_n N_VGND_c_965_n 2.3658e-19 $X=4.305 $Y=0.84 $X2=0
+ $Y2=0
cc_476 N_A_809_21#_c_584_n N_VGND_c_965_n 0.0119203f $X=4.99 $Y=0.51 $X2=0 $Y2=0
cc_477 N_A_809_21#_M1011_g N_VGND_c_966_n 0.00369209f $X=6.105 $Y=0.785 $X2=0
+ $Y2=0
cc_478 N_A_809_21#_c_586_n N_VGND_c_966_n 0.00526356f $X=6.195 $Y=1.505 $X2=0
+ $Y2=0
cc_479 N_A_809_21#_c_584_n N_VGND_c_967_n 0.0168381f $X=4.99 $Y=0.51 $X2=0 $Y2=0
cc_480 N_A_809_21#_c_581_n N_VGND_c_970_n 0.00378975f $X=4.12 $Y=0.765 $X2=0
+ $Y2=0
cc_481 N_A_809_21#_c_583_n N_VGND_c_970_n 4.89446e-19 $X=4.305 $Y=0.84 $X2=0
+ $Y2=0
cc_482 N_A_809_21#_M1011_g N_VGND_c_971_n 0.00443766f $X=6.105 $Y=0.785 $X2=0
+ $Y2=0
cc_483 N_A_809_21#_c_581_n N_VGND_c_972_n 0.0067851f $X=4.12 $Y=0.765 $X2=0
+ $Y2=0
cc_484 N_A_809_21#_M1011_g N_VGND_c_972_n 0.00856022f $X=6.105 $Y=0.785 $X2=0
+ $Y2=0
cc_485 N_A_809_21#_c_584_n N_VGND_c_972_n 0.0134058f $X=4.99 $Y=0.51 $X2=0 $Y2=0
cc_486 N_A_659_47#_M1006_g N_RESET_B_M1019_g 0.0435445f $X=5.205 $Y=0.785 $X2=0
+ $Y2=0
cc_487 N_A_659_47#_M1004_g N_RESET_B_M1016_g 0.0327799f $X=5.205 $Y=2.465 $X2=0
+ $Y2=0
cc_488 N_A_659_47#_M1006_g RESET_B 0.00331404f $X=5.205 $Y=0.785 $X2=0 $Y2=0
cc_489 N_A_659_47#_c_706_n RESET_B 0.00331404f $X=5.205 $Y=1.5 $X2=0 $Y2=0
cc_490 N_A_659_47#_c_706_n N_RESET_B_c_813_n 0.0435445f $X=5.205 $Y=1.5 $X2=0
+ $Y2=0
cc_491 N_A_659_47#_M1004_g N_RESET_B_c_814_n 0.00331404f $X=5.205 $Y=2.465 $X2=0
+ $Y2=0
cc_492 N_A_659_47#_M1004_g N_VPWR_c_862_n 0.0054895f $X=5.205 $Y=2.465 $X2=0
+ $Y2=0
cc_493 N_A_659_47#_M1004_g N_VPWR_c_858_n 0.00758249f $X=5.205 $Y=2.465 $X2=0
+ $Y2=0
cc_494 N_A_659_47#_M1004_g N_VPWR_c_870_n 0.00877502f $X=5.205 $Y=2.465 $X2=0
+ $Y2=0
cc_495 N_A_659_47#_c_720_n N_VGND_c_964_n 0.00687891f $X=4.005 $Y=0.425 $X2=0
+ $Y2=0
cc_496 N_A_659_47#_M1006_g N_VGND_c_965_n 0.00304769f $X=5.205 $Y=0.785 $X2=0
+ $Y2=0
cc_497 N_A_659_47#_c_720_n N_VGND_c_965_n 0.017769f $X=4.005 $Y=0.425 $X2=0
+ $Y2=0
cc_498 N_A_659_47#_c_708_n N_VGND_c_965_n 0.0014134f $X=4.09 $Y=0.725 $X2=0
+ $Y2=0
cc_499 N_A_659_47#_c_709_n N_VGND_c_965_n 0.0202455f $X=4.535 $Y=0.81 $X2=0
+ $Y2=0
cc_500 N_A_659_47#_M1006_g N_VGND_c_967_n 0.00323392f $X=5.205 $Y=0.785 $X2=0
+ $Y2=0
cc_501 N_A_659_47#_c_709_n N_VGND_c_967_n 0.00185996f $X=4.535 $Y=0.81 $X2=0
+ $Y2=0
cc_502 N_A_659_47#_c_720_n N_VGND_c_970_n 0.0335141f $X=4.005 $Y=0.425 $X2=0
+ $Y2=0
cc_503 N_A_659_47#_c_709_n N_VGND_c_970_n 0.00253464f $X=4.535 $Y=0.81 $X2=0
+ $Y2=0
cc_504 N_A_659_47#_M1005_d N_VGND_c_972_n 0.00357675f $X=3.295 $Y=0.235 $X2=0
+ $Y2=0
cc_505 N_A_659_47#_M1006_g N_VGND_c_972_n 0.0047183f $X=5.205 $Y=0.785 $X2=0
+ $Y2=0
cc_506 N_A_659_47#_c_720_n N_VGND_c_972_n 0.0277614f $X=4.005 $Y=0.425 $X2=0
+ $Y2=0
cc_507 N_A_659_47#_c_709_n N_VGND_c_972_n 0.00860976f $X=4.535 $Y=0.81 $X2=0
+ $Y2=0
cc_508 N_A_659_47#_c_720_n A_767_47# 0.00276484f $X=4.005 $Y=0.425 $X2=-0.19
+ $Y2=-0.245
cc_509 N_RESET_B_M1016_g N_VPWR_c_861_n 0.00259664f $X=5.635 $Y=2.465 $X2=0
+ $Y2=0
cc_510 N_RESET_B_M1016_g N_VPWR_c_862_n 0.00585385f $X=5.635 $Y=2.465 $X2=0
+ $Y2=0
cc_511 N_RESET_B_M1016_g N_VPWR_c_858_n 0.00651119f $X=5.635 $Y=2.465 $X2=0
+ $Y2=0
cc_512 N_RESET_B_M1019_g N_VGND_c_966_n 0.00855674f $X=5.565 $Y=0.785 $X2=0
+ $Y2=0
cc_513 RESET_B N_VGND_c_966_n 0.0592671f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_514 N_RESET_B_c_813_n N_VGND_c_966_n 0.00194488f $X=5.655 $Y=1.51 $X2=0 $Y2=0
cc_515 N_RESET_B_M1019_g N_VGND_c_967_n 0.00334856f $X=5.565 $Y=0.785 $X2=0
+ $Y2=0
cc_516 RESET_B N_VGND_c_967_n 0.00776145f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_517 N_RESET_B_M1019_g N_VGND_c_972_n 0.00500611f $X=5.565 $Y=0.785 $X2=0
+ $Y2=0
cc_518 RESET_B N_VGND_c_972_n 0.00604519f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_519 RESET_B A_1056_73# 0.00698634f $X=5.435 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_520 N_VPWR_c_858_n N_Q_M1018_d 0.00371702f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_521 N_VPWR_c_866_n Q 0.0256966f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_522 N_VPWR_c_858_n Q 0.014307f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_523 N_Q_c_941_n N_VGND_c_966_n 0.0333777f $X=6.32 $Y=0.51 $X2=0 $Y2=0
cc_524 N_Q_c_941_n N_VGND_c_971_n 0.0212526f $X=6.32 $Y=0.51 $X2=0 $Y2=0
cc_525 N_Q_c_941_n N_VGND_c_972_n 0.0172451f $X=6.32 $Y=0.51 $X2=0 $Y2=0
cc_526 N_VGND_c_972_n A_587_47# 0.00265743f $X=6.48 $Y=0 $X2=-0.19 $Y2=-0.245
cc_527 N_VGND_c_972_n A_767_47# 0.00172061f $X=6.48 $Y=0 $X2=-0.19 $Y2=-0.245
