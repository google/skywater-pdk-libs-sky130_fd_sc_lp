* NGSPICE file created from sky130_fd_sc_lp__o2111ai_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o2111ai_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 VPWR C1 Y VPB phighvt w=640000u l=150000u
+  ad=9.536e+11p pd=6.82e+06u as=3.904e+11p ps=3.78e+06u
M1001 VGND A2 a_339_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=3.717e+11p ps=3.45e+06u
M1002 Y B1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y D1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_339_47# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_520_465# A2 Y VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1006 a_195_47# D1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.541e+11p ps=2.05e+06u
M1007 a_267_47# C1 a_195_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 VPWR A1 a_520_465# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_339_47# B1 a_267_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

