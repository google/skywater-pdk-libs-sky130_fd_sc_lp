* File: sky130_fd_sc_lp__a21o_0.pxi.spice
* Created: Fri Aug 28 09:50:36 2020
* 
x_PM_SKY130_FD_SC_LP__A21O_0%A_80_275# N_A_80_275#_M1002_d N_A_80_275#_M1000_s
+ N_A_80_275#_M1003_g N_A_80_275#_c_68_n N_A_80_275#_c_69_n N_A_80_275#_M1007_g
+ N_A_80_275#_c_71_n N_A_80_275#_c_72_n N_A_80_275#_c_73_n N_A_80_275#_c_80_n
+ N_A_80_275#_c_74_n N_A_80_275#_c_75_n N_A_80_275#_c_76_n N_A_80_275#_c_77_n
+ N_A_80_275#_c_78_n N_A_80_275#_c_82_n PM_SKY130_FD_SC_LP__A21O_0%A_80_275#
x_PM_SKY130_FD_SC_LP__A21O_0%B1 N_B1_M1002_g N_B1_M1000_g N_B1_c_134_n
+ N_B1_c_135_n B1 B1 N_B1_c_136_n N_B1_c_137_n PM_SKY130_FD_SC_LP__A21O_0%B1
x_PM_SKY130_FD_SC_LP__A21O_0%A1 N_A1_M1004_g N_A1_M1006_g N_A1_c_179_n
+ N_A1_c_183_n A1 A1 A1 A1 N_A1_c_181_n A1 PM_SKY130_FD_SC_LP__A21O_0%A1
x_PM_SKY130_FD_SC_LP__A21O_0%A2 N_A2_c_227_n N_A2_M1005_g N_A2_M1001_g
+ N_A2_c_228_n N_A2_c_229_n N_A2_c_235_n N_A2_c_230_n A2 A2 A2 N_A2_c_232_n
+ PM_SKY130_FD_SC_LP__A21O_0%A2
x_PM_SKY130_FD_SC_LP__A21O_0%X N_X_M1007_s N_X_M1003_s N_X_c_270_n X X X X X X X
+ N_X_c_272_n PM_SKY130_FD_SC_LP__A21O_0%X
x_PM_SKY130_FD_SC_LP__A21O_0%VPWR N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_c_291_n
+ N_VPWR_c_292_n VPWR N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_295_n
+ N_VPWR_c_290_n N_VPWR_c_297_n N_VPWR_c_298_n PM_SKY130_FD_SC_LP__A21O_0%VPWR
x_PM_SKY130_FD_SC_LP__A21O_0%A_319_473# N_A_319_473#_M1000_d
+ N_A_319_473#_M1001_d N_A_319_473#_c_324_n N_A_319_473#_c_325_n
+ N_A_319_473#_c_326_n N_A_319_473#_c_327_n
+ PM_SKY130_FD_SC_LP__A21O_0%A_319_473#
x_PM_SKY130_FD_SC_LP__A21O_0%VGND N_VGND_M1007_d N_VGND_M1005_d N_VGND_c_352_n
+ N_VGND_c_353_n N_VGND_c_354_n VGND N_VGND_c_355_n N_VGND_c_356_n
+ N_VGND_c_357_n N_VGND_c_358_n PM_SKY130_FD_SC_LP__A21O_0%VGND
cc_1 VNB N_A_80_275#_M1003_g 0.00838526f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_2 VNB N_A_80_275#_c_68_n 0.0339399f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.45
cc_3 VNB N_A_80_275#_c_69_n 0.0143573f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.45
cc_4 VNB N_A_80_275#_M1007_g 0.0260553f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.445
cc_5 VNB N_A_80_275#_c_71_n 0.0264246f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.375
cc_6 VNB N_A_80_275#_c_72_n 0.00304983f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.02
cc_7 VNB N_A_80_275#_c_73_n 0.017984f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.02
cc_8 VNB N_A_80_275#_c_74_n 0.00929619f $X=-0.19 $Y=-0.245 $X2=1.55 $Y2=0.825
cc_9 VNB N_A_80_275#_c_75_n 0.00473557f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.825
cc_10 VNB N_A_80_275#_c_76_n 0.00147743f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.445
cc_11 VNB N_A_80_275#_c_77_n 0.0146932f $X=-0.19 $Y=-0.245 $X2=0.957 $Y2=1.525
cc_12 VNB N_A_80_275#_c_78_n 0.00228447f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.055
cc_13 VNB N_B1_M1002_g 0.0342131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_134_n 0.022359f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.45
cc_15 VNB N_B1_c_135_n 0.00489944f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.45
cc_16 VNB N_B1_c_136_n 0.0157002f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=0.855
cc_17 VNB N_B1_c_137_n 0.00578518f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.375
cc_18 VNB N_A1_M1004_g 0.0364437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_179_n 0.0214986f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.45
cc_20 VNB A1 0.00443152f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.445
cc_21 VNB N_A1_c_181_n 0.0157584f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.02
cc_22 VNB N_A2_c_227_n 0.0212662f $X=-0.19 $Y=-0.245 $X2=1.53 $Y2=0.235
cc_23 VNB N_A2_c_228_n 0.00891899f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_24 VNB N_A2_c_229_n 0.0333851f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.855
cc_25 VNB N_A2_c_230_n 0.0185653f $X=-0.19 $Y=-0.245 $X2=0.957 $Y2=0.91
cc_26 VNB A2 0.0327919f $X=-0.19 $Y=-0.245 $X2=0.957 $Y2=1.278
cc_27 VNB N_A2_c_232_n 0.0363074f $X=-0.19 $Y=-0.245 $X2=1.282 $Y2=2.51
cc_28 VNB N_X_c_270_n 0.0130354f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_29 VNB X 0.0599398f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.45
cc_30 VNB N_X_c_272_n 0.0195816f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.055
cc_31 VNB N_VPWR_c_290_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_352_n 0.00561404f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_33 VNB N_VGND_c_353_n 0.0120881f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.45
cc_34 VNB N_VGND_c_354_n 0.0188195f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.855
cc_35 VNB N_VGND_c_355_n 0.0283918f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.02
cc_36 VNB N_VGND_c_356_n 0.0293867f $X=-0.19 $Y=-0.245 $X2=0.957 $Y2=1.02
cc_37 VNB N_VGND_c_357_n 0.00632031f $X=-0.19 $Y=-0.245 $X2=1.282 $Y2=2.51
cc_38 VNB N_VGND_c_358_n 0.172325f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.825
cc_39 VPB N_A_80_275#_M1003_g 0.0650741f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_40 VPB N_A_80_275#_c_80_n 0.0139249f $X=-0.19 $Y=1.655 $X2=1.305 $Y2=2.51
cc_41 VPB N_A_80_275#_c_78_n 0.0101019f $X=-0.19 $Y=1.655 $X2=1.23 $Y2=2.055
cc_42 VPB N_A_80_275#_c_82_n 0.0150746f $X=-0.19 $Y=1.655 $X2=1.23 $Y2=2.225
cc_43 VPB N_B1_M1000_g 0.0473582f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.525
cc_44 VPB N_B1_c_135_n 0.0117805f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.45
cc_45 VPB N_B1_c_137_n 0.00483496f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.375
cc_46 VPB N_A1_M1006_g 0.0397156f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.525
cc_47 VPB N_A1_c_183_n 0.0158728f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.45
cc_48 VPB A1 0.00376771f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=0.445
cc_49 VPB N_A2_M1001_g 0.0226699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A2_c_228_n 0.0298101f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_51 VPB N_A2_c_235_n 0.0193948f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.02
cc_52 VPB A2 0.00952973f $X=-0.19 $Y=1.655 $X2=0.957 $Y2=1.278
cc_53 VPB X 0.0720449f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.45
cc_54 VPB N_VPWR_c_291_n 0.0258536f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_55 VPB N_VPWR_c_292_n 0.010042f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=0.855
cc_56 VPB N_VPWR_c_293_n 0.0172252f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.02
cc_57 VPB N_VPWR_c_294_n 0.0328891f $X=-0.19 $Y=1.655 $X2=0.957 $Y2=1.02
cc_58 VPB N_VPWR_c_295_n 0.0182082f $X=-0.19 $Y=1.655 $X2=1.305 $Y2=2.51
cc_59 VPB N_VPWR_c_290_n 0.0683785f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_297_n 0.00555219f $X=-0.19 $Y=1.655 $X2=1.667 $Y2=0.74
cc_61 VPB N_VPWR_c_298_n 0.00487897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_319_473#_c_324_n 0.00590952f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_63 VPB N_A_319_473#_c_325_n 0.0180949f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.45
cc_64 VPB N_A_319_473#_c_326_n 0.00578121f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.45
cc_65 VPB N_A_319_473#_c_327_n 0.0358998f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=0.445
cc_66 N_A_80_275#_M1007_g N_B1_M1002_g 0.0208042f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_67 N_A_80_275#_c_72_n N_B1_M1002_g 0.00438952f $X=0.875 $Y=1.02 $X2=0 $Y2=0
cc_68 N_A_80_275#_c_74_n N_B1_M1002_g 0.012608f $X=1.55 $Y=0.825 $X2=0 $Y2=0
cc_69 N_A_80_275#_c_76_n N_B1_M1002_g 0.00236935f $X=1.68 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_80_275#_c_78_n N_B1_M1000_g 0.00701711f $X=1.23 $Y=2.055 $X2=0 $Y2=0
cc_71 N_A_80_275#_c_82_n N_B1_M1000_g 0.00771356f $X=1.23 $Y=2.225 $X2=0 $Y2=0
cc_72 N_A_80_275#_c_68_n N_B1_c_134_n 0.0101822f $X=0.71 $Y=1.45 $X2=0 $Y2=0
cc_73 N_A_80_275#_c_77_n N_B1_c_134_n 0.00298031f $X=0.957 $Y=1.525 $X2=0 $Y2=0
cc_74 N_A_80_275#_c_78_n N_B1_c_135_n 0.00298031f $X=1.23 $Y=2.055 $X2=0 $Y2=0
cc_75 N_A_80_275#_c_82_n N_B1_c_135_n 0.0036079f $X=1.23 $Y=2.225 $X2=0 $Y2=0
cc_76 N_A_80_275#_c_71_n N_B1_c_136_n 0.0101822f $X=0.875 $Y=1.375 $X2=0 $Y2=0
cc_77 N_A_80_275#_c_72_n N_B1_c_136_n 0.00298031f $X=0.875 $Y=1.02 $X2=0 $Y2=0
cc_78 N_A_80_275#_c_74_n N_B1_c_136_n 0.0038778f $X=1.55 $Y=0.825 $X2=0 $Y2=0
cc_79 N_A_80_275#_c_71_n N_B1_c_137_n 3.79227e-19 $X=0.875 $Y=1.375 $X2=0 $Y2=0
cc_80 N_A_80_275#_c_72_n N_B1_c_137_n 0.057803f $X=0.875 $Y=1.02 $X2=0 $Y2=0
cc_81 N_A_80_275#_c_74_n N_B1_c_137_n 0.0339442f $X=1.55 $Y=0.825 $X2=0 $Y2=0
cc_82 N_A_80_275#_c_82_n N_B1_c_137_n 0.00292015f $X=1.23 $Y=2.225 $X2=0 $Y2=0
cc_83 N_A_80_275#_c_74_n N_A1_M1004_g 0.0014103f $X=1.55 $Y=0.825 $X2=0 $Y2=0
cc_84 N_A_80_275#_c_76_n N_A1_M1004_g 0.00350679f $X=1.68 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_80_275#_c_74_n A1 0.0143625f $X=1.55 $Y=0.825 $X2=0 $Y2=0
cc_86 N_A_80_275#_c_76_n A1 0.027403f $X=1.68 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_80_275#_c_73_n N_X_c_270_n 9.19401e-19 $X=0.875 $Y=1.02 $X2=0 $Y2=0
cc_88 N_A_80_275#_c_75_n N_X_c_270_n 0.0123978f $X=1.205 $Y=0.825 $X2=0 $Y2=0
cc_89 N_A_80_275#_c_69_n X 0.0352903f $X=0.55 $Y=1.45 $X2=0 $Y2=0
cc_90 N_A_80_275#_M1007_g X 0.00404473f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_80_275#_c_72_n X 0.0314129f $X=0.875 $Y=1.02 $X2=0 $Y2=0
cc_92 N_A_80_275#_c_73_n X 0.00994234f $X=0.875 $Y=1.02 $X2=0 $Y2=0
cc_93 N_A_80_275#_c_75_n X 0.00840406f $X=1.205 $Y=0.825 $X2=0 $Y2=0
cc_94 N_A_80_275#_c_78_n X 0.0219735f $X=1.23 $Y=2.055 $X2=0 $Y2=0
cc_95 N_A_80_275#_M1003_g N_VPWR_c_291_n 0.00504732f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_96 N_A_80_275#_c_80_n N_VPWR_c_291_n 0.0358911f $X=1.305 $Y=2.51 $X2=0 $Y2=0
cc_97 N_A_80_275#_M1003_g N_VPWR_c_293_n 0.00545548f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_98 N_A_80_275#_c_80_n N_VPWR_c_294_n 0.0153957f $X=1.305 $Y=2.51 $X2=0 $Y2=0
cc_99 N_A_80_275#_M1003_g N_VPWR_c_290_n 0.0120267f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_100 N_A_80_275#_c_80_n N_VPWR_c_290_n 0.010726f $X=1.305 $Y=2.51 $X2=0 $Y2=0
cc_101 N_A_80_275#_c_82_n N_A_319_473#_c_324_n 0.0428014f $X=1.23 $Y=2.225 $X2=0
+ $Y2=0
cc_102 N_A_80_275#_c_78_n N_A_319_473#_c_326_n 0.00211536f $X=1.23 $Y=2.055
+ $X2=0 $Y2=0
cc_103 N_A_80_275#_c_82_n N_A_319_473#_c_326_n 0.0101966f $X=1.23 $Y=2.225 $X2=0
+ $Y2=0
cc_104 N_A_80_275#_M1007_g N_VGND_c_352_n 0.0033471f $X=0.965 $Y=0.445 $X2=0
+ $Y2=0
cc_105 N_A_80_275#_c_74_n N_VGND_c_352_n 0.0113433f $X=1.55 $Y=0.825 $X2=0 $Y2=0
cc_106 N_A_80_275#_c_75_n N_VGND_c_352_n 0.0115505f $X=1.205 $Y=0.825 $X2=0
+ $Y2=0
cc_107 N_A_80_275#_M1007_g N_VGND_c_355_n 0.0058053f $X=0.965 $Y=0.445 $X2=0
+ $Y2=0
cc_108 N_A_80_275#_c_75_n N_VGND_c_355_n 2.29031e-19 $X=1.205 $Y=0.825 $X2=0
+ $Y2=0
cc_109 N_A_80_275#_c_74_n N_VGND_c_356_n 0.00222198f $X=1.55 $Y=0.825 $X2=0
+ $Y2=0
cc_110 N_A_80_275#_c_76_n N_VGND_c_356_n 0.0129772f $X=1.68 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_80_275#_M1002_d N_VGND_c_358_n 0.00604286f $X=1.53 $Y=0.235 $X2=0
+ $Y2=0
cc_112 N_A_80_275#_M1007_g N_VGND_c_358_n 0.00771011f $X=0.965 $Y=0.445 $X2=0
+ $Y2=0
cc_113 N_A_80_275#_c_74_n N_VGND_c_358_n 0.00438922f $X=1.55 $Y=0.825 $X2=0
+ $Y2=0
cc_114 N_A_80_275#_c_75_n N_VGND_c_358_n 0.00670992f $X=1.205 $Y=0.825 $X2=0
+ $Y2=0
cc_115 N_A_80_275#_c_76_n N_VGND_c_358_n 0.00892897f $X=1.68 $Y=0.445 $X2=0
+ $Y2=0
cc_116 N_B1_M1002_g N_A1_M1004_g 0.0190003f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_117 N_B1_c_136_n N_A1_M1004_g 0.0115258f $X=1.47 $Y=1.245 $X2=0 $Y2=0
cc_118 N_B1_c_137_n N_A1_M1004_g 0.00540004f $X=1.47 $Y=1.245 $X2=0 $Y2=0
cc_119 N_B1_c_135_n N_A1_c_179_n 0.0115258f $X=1.47 $Y=1.75 $X2=0 $Y2=0
cc_120 N_B1_M1000_g N_A1_c_183_n 0.0318751f $X=1.52 $Y=2.685 $X2=0 $Y2=0
cc_121 N_B1_M1002_g A1 2.31087e-19 $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_122 N_B1_M1002_g A1 8.69456e-19 $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B1_c_136_n A1 5.68885e-19 $X=1.47 $Y=1.245 $X2=0 $Y2=0
cc_124 N_B1_c_137_n A1 0.0604337f $X=1.47 $Y=1.245 $X2=0 $Y2=0
cc_125 N_B1_c_134_n N_A1_c_181_n 0.0115258f $X=1.47 $Y=1.585 $X2=0 $Y2=0
cc_126 N_B1_M1000_g N_VPWR_c_291_n 0.00326526f $X=1.52 $Y=2.685 $X2=0 $Y2=0
cc_127 N_B1_M1000_g N_VPWR_c_294_n 0.00499542f $X=1.52 $Y=2.685 $X2=0 $Y2=0
cc_128 N_B1_M1000_g N_VPWR_c_290_n 0.0104152f $X=1.52 $Y=2.685 $X2=0 $Y2=0
cc_129 N_B1_M1000_g N_A_319_473#_c_324_n 0.001706f $X=1.52 $Y=2.685 $X2=0 $Y2=0
cc_130 N_B1_M1000_g N_A_319_473#_c_326_n 0.00177623f $X=1.52 $Y=2.685 $X2=0
+ $Y2=0
cc_131 N_B1_c_135_n N_A_319_473#_c_326_n 2.54754e-19 $X=1.47 $Y=1.75 $X2=0 $Y2=0
cc_132 N_B1_c_137_n N_A_319_473#_c_326_n 0.0173454f $X=1.47 $Y=1.245 $X2=0 $Y2=0
cc_133 N_B1_M1002_g N_VGND_c_352_n 0.00341356f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_134 N_B1_M1002_g N_VGND_c_356_n 0.00439071f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_135 N_B1_M1002_g N_VGND_c_358_n 0.00637652f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_136 N_A1_M1004_g N_A2_c_227_n 0.0444996f $X=1.95 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_137 A1 N_A2_c_227_n 0.0138583f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_138 N_A1_M1006_g N_A2_c_228_n 0.00772999f $X=1.95 $Y=2.685 $X2=0 $Y2=0
cc_139 N_A1_c_183_n N_A2_c_228_n 0.0113746f $X=2.04 $Y=1.825 $X2=0 $Y2=0
cc_140 A1 N_A2_c_229_n 8.20289e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_141 A1 N_A2_c_229_n 0.00520644f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_142 N_A1_M1006_g N_A2_c_235_n 0.0180168f $X=1.95 $Y=2.685 $X2=0 $Y2=0
cc_143 N_A1_c_179_n N_A2_c_230_n 0.0113746f $X=2.04 $Y=1.66 $X2=0 $Y2=0
cc_144 A1 N_A2_c_230_n 0.00322951f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_145 N_A1_M1004_g A2 2.78937e-19 $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_146 A1 A2 0.0825863f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_147 N_A1_c_181_n A2 6.56752e-19 $X=2.04 $Y=1.32 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_A2_c_232_n 0.00569061f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_149 A1 N_A2_c_232_n 0.00322951f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_150 N_A1_c_181_n N_A2_c_232_n 0.0113746f $X=2.04 $Y=1.32 $X2=0 $Y2=0
cc_151 N_A1_M1006_g N_VPWR_c_292_n 0.00308207f $X=1.95 $Y=2.685 $X2=0 $Y2=0
cc_152 N_A1_M1006_g N_VPWR_c_294_n 0.00499542f $X=1.95 $Y=2.685 $X2=0 $Y2=0
cc_153 N_A1_M1006_g N_VPWR_c_290_n 0.00973692f $X=1.95 $Y=2.685 $X2=0 $Y2=0
cc_154 N_A1_M1006_g N_A_319_473#_c_324_n 0.0027941f $X=1.95 $Y=2.685 $X2=0 $Y2=0
cc_155 N_A1_M1006_g N_A_319_473#_c_325_n 0.0176957f $X=1.95 $Y=2.685 $X2=0 $Y2=0
cc_156 N_A1_c_183_n N_A_319_473#_c_325_n 0.00121735f $X=2.04 $Y=1.825 $X2=0
+ $Y2=0
cc_157 A1 N_A_319_473#_c_325_n 0.0292401f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_158 N_A1_M1004_g N_VGND_c_356_n 0.00492032f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_159 A1 N_VGND_c_356_n 0.011025f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_160 N_A1_M1004_g N_VGND_c_358_n 0.00857209f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_161 A1 N_VGND_c_358_n 0.0119334f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_162 A1 N_VGND_c_358_n 3.04069e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_163 A1 A_405_47# 0.00157923f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_164 N_A2_M1001_g N_VPWR_c_292_n 0.003107f $X=2.38 $Y=2.685 $X2=0 $Y2=0
cc_165 N_A2_M1001_g N_VPWR_c_295_n 0.00499542f $X=2.38 $Y=2.685 $X2=0 $Y2=0
cc_166 N_A2_M1001_g N_VPWR_c_290_n 0.0100834f $X=2.38 $Y=2.685 $X2=0 $Y2=0
cc_167 N_A2_c_228_n N_A_319_473#_c_325_n 0.0061292f $X=2.52 $Y=2.065 $X2=0 $Y2=0
cc_168 N_A2_c_235_n N_A_319_473#_c_325_n 0.015311f $X=2.52 $Y=2.14 $X2=0 $Y2=0
cc_169 N_A2_c_230_n N_A_319_473#_c_325_n 6.54377e-19 $X=2.61 $Y=1.51 $X2=0 $Y2=0
cc_170 A2 N_A_319_473#_c_325_n 0.0245687f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_171 N_A2_M1001_g N_A_319_473#_c_327_n 0.00483547f $X=2.38 $Y=2.685 $X2=0
+ $Y2=0
cc_172 N_A2_c_235_n N_A_319_473#_c_327_n 0.00507638f $X=2.52 $Y=2.14 $X2=0 $Y2=0
cc_173 N_A2_c_229_n N_VGND_c_353_n 0.00109359f $X=2.61 $Y=0.915 $X2=0 $Y2=0
cc_174 N_A2_c_227_n N_VGND_c_354_n 0.00476035f $X=2.34 $Y=0.765 $X2=0 $Y2=0
cc_175 N_A2_c_229_n N_VGND_c_354_n 0.00705477f $X=2.61 $Y=0.915 $X2=0 $Y2=0
cc_176 A2 N_VGND_c_354_n 0.0202609f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_177 N_A2_c_227_n N_VGND_c_356_n 0.00539385f $X=2.34 $Y=0.765 $X2=0 $Y2=0
cc_178 N_A2_c_229_n N_VGND_c_356_n 9.57268e-19 $X=2.61 $Y=0.915 $X2=0 $Y2=0
cc_179 N_A2_c_227_n N_VGND_c_358_n 0.0102824f $X=2.34 $Y=0.765 $X2=0 $Y2=0
cc_180 N_A2_c_229_n N_VGND_c_358_n 0.00280483f $X=2.61 $Y=0.915 $X2=0 $Y2=0
cc_181 A2 N_VGND_c_358_n 0.00375713f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_182 X N_VPWR_c_291_n 0.00311641f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_183 X N_VPWR_c_293_n 0.0220795f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_184 X N_VPWR_c_290_n 0.0119743f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_185 N_X_c_270_n N_VGND_c_355_n 0.0267391f $X=0.75 $Y=0.445 $X2=0 $Y2=0
cc_186 N_X_c_272_n N_VGND_c_355_n 0.0191846f $X=0.24 $Y=0.61 $X2=0 $Y2=0
cc_187 N_X_M1007_s N_VGND_c_358_n 0.00222632f $X=0.625 $Y=0.235 $X2=0 $Y2=0
cc_188 N_X_c_270_n N_VGND_c_358_n 0.018247f $X=0.75 $Y=0.445 $X2=0 $Y2=0
cc_189 N_X_c_272_n N_VGND_c_358_n 0.0119057f $X=0.24 $Y=0.61 $X2=0 $Y2=0
cc_190 N_VPWR_c_292_n N_A_319_473#_c_324_n 0.00305835f $X=2.165 $Y=2.51 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_294_n N_A_319_473#_c_324_n 0.0148517f $X=2.04 $Y=3.33 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_290_n N_A_319_473#_c_324_n 0.010347f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_292_n N_A_319_473#_c_325_n 0.0213684f $X=2.165 $Y=2.51 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_292_n N_A_319_473#_c_327_n 0.00307479f $X=2.165 $Y=2.51 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_295_n N_A_319_473#_c_327_n 0.0159397f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_290_n N_A_319_473#_c_327_n 0.0111051f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_197 N_VGND_c_358_n A_405_47# 0.00206003f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
