* File: sky130_fd_sc_lp__a221oi_0.spice
* Created: Wed Sep  2 09:21:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a221oi_0.pex.spice"
.subckt sky130_fd_sc_lp__a221oi_0  VNB VPB C1 B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_C1_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.08715 AS=0.1113 PD=0.835 PS=1.37 NRD=8.568 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1000 A_228_47# N_B2_M1000_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.08715 PD=0.66 PS=0.835 NRD=18.564 NRS=30 M=1 R=2.8 SA=75000.8 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g A_228_47# VNB NSHORT L=0.15 W=0.42 AD=0.0756
+ AS=0.0504 PD=0.78 PS=0.66 NRD=12.852 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 A_408_47# N_A1_M1006_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=9.996 M=1 R=2.8 SA=75001.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_408_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_156_487#_M1007_d N_C1_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_242_487#_M1002_d N_B2_M1002_g N_A_156_487#_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1312 AS=0.0896 PD=1.05 PS=0.92 NRD=40.0107 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_242_487#_M1002_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.112 AS=0.1312 PD=0.99 PS=1.05 NRD=21.5321 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1004 N_A_242_487#_M1004_d N_A2_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.112 AS=0.112 PD=0.99 PS=0.99 NRD=21.5321 NRS=0 M=1 R=4.26667
+ SA=75001.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1008 N_A_156_487#_M1008_d N_B1_M1008_g N_A_242_487#_M1004_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2144 AS=0.112 PD=1.95 PS=0.99 NRD=21.5321 NRS=0 M=1 R=4.26667
+ SA=75002.2 SB=75000.3 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a221oi_0.pxi.spice"
*
.ends
*
*
