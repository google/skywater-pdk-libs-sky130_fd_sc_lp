* File: sky130_fd_sc_lp__nor2_lp2.pex.spice
* Created: Fri Aug 28 10:53:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2_LP2%A 3 7 9 13 15 17 23
r33 26 28 31.9995 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=1.51
r34 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=1.345 $X2=0.485 $Y2=1.345
r35 23 26 14.8382 $w=3.5e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=1.255
+ $X2=0.495 $Y2=1.345
r36 23 24 31.5932 $w=3.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.255
+ $X2=0.495 $Y2=1.18
r37 17 27 4.68464 $w=5.98e-07 $l=2.35e-07 $layer=LI1_cond $X=0.72 $Y=1.48
+ $X2=0.485 $Y2=1.48
r38 15 27 4.88399 $w=5.98e-07 $l=2.45e-07 $layer=LI1_cond $X=0.24 $Y=1.48
+ $X2=0.485 $Y2=1.48
r39 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.965 $Y=1.18
+ $X2=0.965 $Y2=0.77
r40 10 23 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.67 $Y=1.255
+ $X2=0.495 $Y2=1.255
r41 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.89 $Y=1.255
+ $X2=0.965 $Y2=1.18
r42 9 10 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.89 $Y=1.255
+ $X2=0.67 $Y2=1.255
r43 7 24 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.575 $Y=0.77
+ $X2=0.575 $Y2=1.18
r44 3 28 213.67 $w=2.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.545 $Y=2.37
+ $X2=0.545 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_LP2%B 1 3 4 5 8 10 14 16 17 18 19 20 21 38
c41 16 0 1.59193e-19 $X=1.395 $Y=1.72
r42 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.875
+ $Y=1.345 $X2=1.875 $Y2=1.345
r43 20 21 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.405
+ $X2=1.92 $Y2=2.775
r44 19 20 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=1.92 $Y2=2.405
r45 18 19 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=1.665
+ $X2=1.92 $Y2=2.035
r46 18 39 5.39078 $w=7.08e-07 $l=3.2e-07 $layer=LI1_cond $X=1.92 $Y=1.665
+ $X2=1.92 $Y2=1.345
r47 17 39 0.842309 $w=7.08e-07 $l=5e-08 $layer=LI1_cond $X=1.92 $Y=1.295
+ $X2=1.92 $Y2=1.345
r48 12 38 39.6178 $w=2.46e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.785 $Y=1.18
+ $X2=1.875 $Y2=1.345
r49 12 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.785 $Y=1.18
+ $X2=1.785 $Y2=0.77
r50 11 16 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.47 $Y=1.72
+ $X2=1.395 $Y2=1.72
r51 10 38 73.4756 $w=2.46e-07 $l=4.5e-07 $layer=POLY_cond $X=1.71 $Y=1.72
+ $X2=1.875 $Y2=1.345
r52 10 11 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.71 $Y=1.72
+ $X2=1.47 $Y2=1.72
r53 6 16 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=1.645
+ $X2=1.395 $Y2=1.72
r54 6 8 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.395 $Y=1.645
+ $X2=1.395 $Y2=0.77
r55 4 16 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.32 $Y=1.72
+ $X2=1.395 $Y2=1.72
r56 4 5 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.32 $Y=1.72 $X2=1.13
+ $Y2=1.72
r57 1 5 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=1.005 $Y=1.795
+ $X2=1.13 $Y2=1.72
r58 1 3 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.005 $Y=1.795
+ $X2=1.005 $Y2=2.37
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_LP2%VPWR 1 4 6 10 17 18
r18 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r19 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r20 15 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r21 14 17 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r22 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r23 12 21 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r24 12 14 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 10 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r26 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 6 9 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=2.065 $X2=0.28
+ $Y2=2.745
r28 4 21 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r29 4 9 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.28 $Y=3.245 $X2=0.28
+ $Y2=2.745
r30 1 9 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.87 $X2=0.28 $Y2=2.745
r31 1 6 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.87 $X2=0.28 $Y2=2.065
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_LP2%Y 1 2 7 8 9 10 11 12 13
r23 12 13 9.70478 $w=3.78e-07 $l=3.2e-07 $layer=LI1_cond $X=1.205 $Y=2.405
+ $X2=1.205 $Y2=2.725
r24 11 12 11.8277 $w=3.78e-07 $l=3.9e-07 $layer=LI1_cond $X=1.205 $Y=2.015
+ $X2=1.205 $Y2=2.405
r25 10 11 10.6146 $w=3.78e-07 $l=3.5e-07 $layer=LI1_cond $X=1.205 $Y=1.665
+ $X2=1.205 $Y2=2.015
r26 9 10 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=1.295
+ $X2=1.205 $Y2=1.665
r27 8 9 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=0.925
+ $X2=1.205 $Y2=1.295
r28 8 25 4.70075 $w=3.78e-07 $l=1.55e-07 $layer=LI1_cond $X=1.205 $Y=0.925
+ $X2=1.205 $Y2=0.77
r29 7 25 6.5204 $w=3.78e-07 $l=2.15e-07 $layer=LI1_cond $X=1.205 $Y=0.555
+ $X2=1.205 $Y2=0.77
r30 2 13 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.87 $X2=1.27 $Y2=2.725
r31 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.87 $X2=1.27 $Y2=2.015
r32 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.56 $X2=1.18 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_LP2%VGND 1 2 7 9 11 13 15 17 30
r26 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r29 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r30 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r31 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r32 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r33 18 26 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.262
+ $Y2=0
r34 18 20 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.72
+ $Y2=0
r35 17 29 4.52492 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2.117
+ $Y2=0
r36 17 23 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.68
+ $Y2=0
r37 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r38 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r39 11 29 3.24126 $w=3.3e-07 $l=1.53734e-07 $layer=LI1_cond $X=2 $Y=0.085
+ $X2=2.117 $Y2=0
r40 11 13 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0.77
r41 7 26 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.262 $Y2=0
r42 7 9 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.36 $Y2=0.77
r43 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.56 $X2=2 $Y2=0.77
r44 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.56 $X2=0.36 $Y2=0.77
.ends

