* File: sky130_fd_sc_lp__o2111a_1.pex.spice
* Created: Wed Sep  2 10:12:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111A_1%A_80_21# 1 2 3 12 15 17 20 23 24 25 28 32
+ 34 36 38 40 43 47
c68 43 0 1.26666e-19 $X=1.755 $Y=2.015
c69 20 0 7.70883e-20 $X=0.63 $Y=1.35
r70 36 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=2.1 $X2=3.095
+ $Y2=2.015
r71 36 38 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.095 $Y=2.1 $X2=3.095
+ $Y2=2.5
r72 35 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.85 $Y=2.015
+ $X2=1.755 $Y2=2.015
r73 34 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=2.015
+ $X2=3.095 $Y2=2.015
r74 34 35 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=2.93 $Y=2.015
+ $X2=1.85 $Y2=2.015
r75 30 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=2.1
+ $X2=1.755 $Y2=2.015
r76 30 32 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.755 $Y=2.1
+ $X2=1.755 $Y2=2.47
r77 26 40 16.4798 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.395 $Y=1.245
+ $X2=1.06 $Y2=1.245
r78 26 28 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.395 $Y=1.075
+ $X2=1.395 $Y2=0.42
r79 24 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.66 $Y=2.015
+ $X2=1.755 $Y2=2.015
r80 24 25 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.66 $Y=2.015
+ $X2=1.145 $Y2=2.015
r81 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=1.93
+ $X2=1.145 $Y2=2.015
r82 22 40 2.94836 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=1.06 $Y=1.515
+ $X2=1.06 $Y2=1.245
r83 22 23 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.06 $Y=1.515
+ $X2=1.06 $Y2=1.93
r84 20 48 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.35
+ $X2=0.597 $Y2=1.515
r85 20 47 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.35
+ $X2=0.597 $Y2=1.185
r86 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.35 $X2=0.63 $Y2=1.35
r87 17 40 3.92342 $w=3.3e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.975 $Y=1.35
+ $X2=1.06 $Y2=1.245
r88 17 19 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.975 $Y=1.35
+ $X2=0.63 $Y2=1.35
r89 15 48 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.515
r90 12 47 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.655
+ $X2=0.475 $Y2=1.185
r91 3 45 600 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_PDIFF $count=1 $X=2.885
+ $Y=1.835 $X2=3.095 $Y2=2.015
r92 3 38 300 $w=1.7e-07 $l=7.62807e-07 $layer=licon1_PDIFF $count=2 $X=2.885
+ $Y=1.835 $X2=3.095 $Y2=2.5
r93 2 43 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=1.615
+ $Y=1.835 $X2=1.755 $Y2=2.015
r94 2 32 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=1.615
+ $Y=1.835 $X2=1.755 $Y2=2.47
r95 1 28 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=1.27
+ $Y=0.245 $X2=1.395 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_1%D1 3 7 9 12
c34 12 0 1.26666e-19 $X=1.49 $Y=1.51
c35 9 0 7.70883e-20 $X=1.68 $Y=1.665
c36 3 0 6.94505e-20 $X=1.54 $Y=2.465
r37 12 15 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.51
+ $X2=1.505 $Y2=1.675
r38 12 14 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.51
+ $X2=1.505 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.51 $X2=1.49 $Y2=1.51
r40 9 13 6.34679 $w=3.43e-07 $l=1.9e-07 $layer=LI1_cond $X=1.68 $Y=1.587
+ $X2=1.49 $Y2=1.587
r41 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.61 $Y=0.665
+ $X2=1.61 $Y2=1.345
r42 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.54 $Y=2.465
+ $X2=1.54 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_1%C1 3 6 8 9 10 11 17 19
c41 19 0 1.30966e-19 $X=2.06 $Y=1.195
c42 17 0 1.79609e-19 $X=2.06 $Y=1.36
c43 8 0 6.94505e-20 $X=2.16 $Y=0.555
r44 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.36
+ $X2=2.06 $Y2=1.525
r45 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.36
+ $X2=2.06 $Y2=1.195
r46 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=1.36 $X2=2.06 $Y2=1.36
r47 11 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=1.36
r48 10 18 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=2.14 $Y=1.295
+ $X2=2.14 $Y2=1.36
r49 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.14 $Y=0.925
+ $X2=2.14 $Y2=1.295
r50 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.14 $Y=0.555 $X2=2.14
+ $Y2=0.925
r51 6 20 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.97 $Y=2.465 $X2=1.97
+ $Y2=1.525
r52 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.97 $Y=0.665
+ $X2=1.97 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_1%B1 3 7 9 15 16
c32 15 0 2.41518e-19 $X=2.64 $Y=1.51
c33 3 0 9.66986e-20 $X=2.51 $Y=0.665
r34 14 16 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.64 $Y=1.51
+ $X2=2.81 $Y2=1.51
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.64
+ $Y=1.51 $X2=2.64 $Y2=1.51
r36 11 14 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.51 $Y=1.51 $X2=2.64
+ $Y2=1.51
r37 9 15 5.49627 $w=3.23e-07 $l=1.55e-07 $layer=LI1_cond $X=2.637 $Y=1.665
+ $X2=2.637 $Y2=1.51
r38 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.675
+ $X2=2.81 $Y2=1.51
r39 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.81 $Y=1.675 $X2=2.81
+ $Y2=2.465
r40 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.345
+ $X2=2.51 $Y2=1.51
r41 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.51 $Y=1.345 $X2=2.51
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_1%A2 3 7 9 10 14
c33 14 0 1.58704e-19 $X=3.26 $Y=1.51
c34 10 0 9.66986e-20 $X=3.6 $Y=1.665
c35 7 0 6.19094e-20 $X=3.35 $Y=2.465
c36 3 0 4.7142e-21 $X=3.28 $Y=0.665
r37 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.51
+ $X2=3.26 $Y2=1.675
r38 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.51
+ $X2=3.26 $Y2=1.345
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.26
+ $Y=1.51 $X2=3.26 $Y2=1.51
r40 10 15 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=3.6 $Y=1.547
+ $X2=3.26 $Y2=1.547
r41 9 15 3.79628 $w=4.23e-07 $l=1.4e-07 $layer=LI1_cond $X=3.12 $Y=1.547
+ $X2=3.26 $Y2=1.547
r42 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.35 $Y=2.465
+ $X2=3.35 $Y2=1.675
r43 3 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.28 $Y=0.665
+ $X2=3.28 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_1%A1 3 7 9 14 15
c23 15 0 1.63418e-19 $X=4.03 $Y=1.46
r24 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.46 $X2=4.03 $Y2=1.46
r25 11 14 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=3.71 $Y=1.46
+ $X2=4.03 $Y2=1.46
r26 9 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.05 $Y=1.665
+ $X2=4.05 $Y2=1.46
r27 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.625
+ $X2=3.71 $Y2=1.46
r28 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.71 $Y=1.625 $X2=3.71
+ $Y2=2.465
r29 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.295
+ $X2=3.71 $Y2=1.46
r30 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.71 $Y=1.295 $X2=3.71
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_1%X 1 2 7 8 9 10 11 12 13 22
r13 13 40 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.23 $Y=2.775
+ $X2=0.23 $Y2=2.91
r14 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=2.405
+ $X2=0.23 $Y2=2.775
r15 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.23 $Y=1.98
+ $X2=0.23 $Y2=2.405
r16 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.23 $Y=1.665
+ $X2=0.23 $Y2=1.98
r17 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.665
r18 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=0.925 $X2=0.23
+ $Y2=1.295
r19 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=0.555 $X2=0.23
+ $Y2=0.925
r20 7 22 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.23 $Y=0.555
+ $X2=0.23 $Y2=0.42
r21 2 40 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r22 2 11 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
r23 1 22 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_1%VPWR 1 2 3 12 17 20 22 24 29 31 33 38 43 49
+ 52 56
r61 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r64 47 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 47 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r67 44 52 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=2.76 $Y=3.33 $X2=2.39
+ $Y2=3.33
r68 44 46 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.76 $Y=3.33 $X2=3.6
+ $Y2=3.33
r69 43 55 4.78145 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.73 $Y=3.33
+ $X2=4.025 $Y2=3.33
r70 43 46 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.73 $Y=3.33 $X2=3.6
+ $Y2=3.33
r71 42 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r72 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 39 49 15.9462 $w=1.7e-07 $l=4.78e-07 $layer=LI1_cond $X=1.49 $Y=3.33
+ $X2=1.012 $Y2=3.33
r74 39 41 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.49 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 38 52 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=2.02 $Y=3.33 $X2=2.39
+ $Y2=3.33
r76 38 41 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.02 $Y=3.33
+ $X2=1.68 $Y2=3.33
r77 36 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r78 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r79 33 49 15.9462 $w=1.7e-07 $l=4.77e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=1.012 $Y2=3.33
r80 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 31 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 29 30 8.10591 $w=9.53e-07 $l=8.5e-08 $layer=LI1_cond $X=1.012 $Y=2.355
+ $X2=1.012 $Y2=2.27
r84 24 27 29.9315 $w=3.58e-07 $l=9.35e-07 $layer=LI1_cond $X=3.91 $Y=2.015
+ $X2=3.91 $Y2=2.95
r85 22 55 3.24166 $w=3.6e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.91 $Y=3.245
+ $X2=4.025 $Y2=3.33
r86 22 27 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.91 $Y=3.245
+ $X2=3.91 $Y2=2.95
r87 18 52 2.97738 $w=7.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=3.245
+ $X2=2.39 $Y2=3.33
r88 18 20 13.9812 $w=7.38e-07 $l=8.65e-07 $layer=LI1_cond $X=2.39 $Y=3.245
+ $X2=2.39 $Y2=2.38
r89 15 49 3.45294 $w=9.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.012 $Y=3.245
+ $X2=1.012 $Y2=3.33
r90 15 17 3.76859 $w=9.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.012 $Y=3.245
+ $X2=1.012 $Y2=2.95
r91 14 29 5.00775 $w=9.53e-07 $l=3.92e-07 $layer=LI1_cond $X=1.012 $Y=2.747
+ $X2=1.012 $Y2=2.355
r92 14 17 2.5933 $w=9.53e-07 $l=2.03e-07 $layer=LI1_cond $X=1.012 $Y=2.747
+ $X2=1.012 $Y2=2.95
r93 12 30 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.67 $Y=1.98
+ $X2=0.67 $Y2=2.27
r94 3 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.785
+ $Y=1.835 $X2=3.925 $Y2=2.95
r95 3 24 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=3.785
+ $Y=1.835 $X2=3.925 $Y2=2.015
r96 2 20 150 $w=1.7e-07 $l=7.76048e-07 $layer=licon1_PDIFF $count=4 $X=2.045
+ $Y=1.835 $X2=2.595 $Y2=2.38
r97 1 29 480 $w=1.7e-07 $l=1.00181e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=1.325 $Y2=2.355
r98 1 17 480 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.95
r99 1 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_1%VGND 1 2 10 13 17 18 19 21 34 35 38
r45 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r47 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r48 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 29 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r50 28 31 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r51 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 26 38 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.695
+ $Y2=0
r53 26 28 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r54 24 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r55 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r56 21 38 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.695
+ $Y2=0
r57 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r58 19 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r59 19 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r60 17 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.12
+ $Y2=0
r61 17 18 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.495
+ $Y2=0
r62 16 34 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.66 $Y=0 $X2=4.08
+ $Y2=0
r63 16 18 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.66 $Y=0 $X2=3.495
+ $Y2=0
r64 11 18 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=0.085
+ $X2=3.495 $Y2=0
r65 11 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.495 $Y=0.085
+ $X2=3.495 $Y2=0.37
r66 7 38 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0
r67 7 10 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0.38
r68 2 13 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.355
+ $Y=0.245 $X2=3.495 $Y2=0.37
r69 1 10 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_1%A_517_49# 1 2 9 11 12 15
c26 12 0 1.30966e-19 $X=3.16 $Y=1.08
r27 13 15 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=3.96 $Y=0.995
+ $X2=3.96 $Y2=0.42
r28 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.83 $Y=1.08
+ $X2=3.96 $Y2=0.995
r29 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.83 $Y=1.08
+ $X2=3.16 $Y2=1.08
r30 7 12 10.0451 $w=1.7e-07 $l=3.39853e-07 $layer=LI1_cond $X=2.86 $Y=0.995
+ $X2=3.16 $Y2=1.08
r31 7 9 11.4624 $w=5.98e-07 $l=5.75e-07 $layer=LI1_cond $X=2.86 $Y=0.995
+ $X2=2.86 $Y2=0.42
r32 2 15 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.785
+ $Y=0.245 $X2=3.925 $Y2=0.42
r33 1 9 45.5 $w=1.7e-07 $l=5.60714e-07 $layer=licon1_NDIFF $count=4 $X=2.585
+ $Y=0.245 $X2=3.065 $Y2=0.42
.ends

