# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__o311ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o311ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.185000 0.945000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 1.185000 1.900000 1.435000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.070000 1.185000 3.205000 1.435000 ;
        RECT 2.340000 1.435000 3.205000 1.525000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.470000 1.185000 4.285000 1.515000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.295000 1.210000 5.675000 1.545000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.818600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.695000 5.125000 1.715000 ;
        RECT 2.375000 1.715000 5.665000 1.865000 ;
        RECT 2.375000 1.865000 2.635000 2.735000 ;
        RECT 3.305000 1.865000 3.495000 3.075000 ;
        RECT 4.455000 0.595000 4.805000 0.870000 ;
        RECT 4.455000 0.870000 5.665000 1.040000 ;
        RECT 4.455000 1.040000 5.125000 1.695000 ;
        RECT 4.545000 1.865000 5.665000 1.885000 ;
        RECT 4.545000 1.885000 4.735000 3.075000 ;
        RECT 5.395000 0.335000 5.665000 0.870000 ;
        RECT 5.405000 1.885000 5.665000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 5.760000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 5.950000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.135000  0.255000 0.395000 0.845000 ;
      RECT 0.135000  0.845000 4.285000 1.015000 ;
      RECT 0.135000  1.605000 2.185000 1.775000 ;
      RECT 0.135000  1.775000 0.395000 3.075000 ;
      RECT 0.565000  0.085000 0.895000 0.675000 ;
      RECT 0.565000  1.945000 0.895000 3.245000 ;
      RECT 1.065000  0.255000 1.255000 0.845000 ;
      RECT 1.065000  1.775000 1.255000 3.075000 ;
      RECT 1.425000  0.085000 1.755000 0.675000 ;
      RECT 1.425000  1.945000 1.755000 2.905000 ;
      RECT 1.425000  2.905000 3.135000 3.075000 ;
      RECT 1.925000  0.255000 2.155000 0.845000 ;
      RECT 1.925000  1.775000 2.185000 2.735000 ;
      RECT 2.325000  0.085000 3.000000 0.675000 ;
      RECT 2.805000  2.035000 3.135000 2.905000 ;
      RECT 3.170000  0.255000 3.355000 0.845000 ;
      RECT 3.525000  0.255000 5.225000 0.425000 ;
      RECT 3.525000  0.425000 3.855000 0.675000 ;
      RECT 3.665000  2.035000 4.375000 3.245000 ;
      RECT 4.025000  0.595000 4.285000 0.845000 ;
      RECT 4.905000  2.055000 5.235000 3.245000 ;
      RECT 4.975000  0.425000 5.225000 0.700000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__o311ai_2
END LIBRARY
