* File: sky130_fd_sc_lp__inv_16.pex.spice
* Created: Fri Aug 28 10:37:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INV_16%A 3 5 7 10 12 14 17 19 21 24 26 28 31 33 35
+ 38 40 42 45 47 49 52 54 56 59 61 63 66 68 70 73 75 77 80 82 84 87 89 91 94 96
+ 98 101 103 105 108 110 112 113 120 125 130 135 140 145 150 152 187
r273 182 187 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=5.495 $Y=1.665
+ $X2=6.355 $Y2=1.665
r274 177 182 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=4.635 $Y=1.665
+ $X2=5.495 $Y2=1.665
r275 162 167 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=2.055 $Y=1.665
+ $X2=2.915 $Y2=1.665
r276 157 162 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=1.195 $Y=1.665
+ $X2=2.055 $Y2=1.665
r277 151 152 61.3195 $w=3.9e-07 $l=4.3e-07 $layer=POLY_cond $X=6.57 $Y=1.53
+ $X2=7 $Y2=1.53
r278 150 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.355 $Y=1.665
+ $X2=6.355 $Y2=1.665
r279 149 151 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=6.355 $Y=1.53
+ $X2=6.57 $Y2=1.53
r280 149 150 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.355
+ $Y=1.5 $X2=6.355 $Y2=1.5
r281 147 149 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=6.14 $Y=1.53
+ $X2=6.355 $Y2=1.53
r282 146 147 61.3195 $w=3.9e-07 $l=4.3e-07 $layer=POLY_cond $X=5.71 $Y=1.53
+ $X2=6.14 $Y2=1.53
r283 145 182 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.495 $Y=1.665
+ $X2=5.495 $Y2=1.665
r284 144 146 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=5.495 $Y=1.53
+ $X2=5.71 $Y2=1.53
r285 144 145 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.495
+ $Y=1.5 $X2=5.495 $Y2=1.5
r286 142 144 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=5.28 $Y=1.53
+ $X2=5.495 $Y2=1.53
r287 141 142 61.3195 $w=3.9e-07 $l=4.3e-07 $layer=POLY_cond $X=4.85 $Y=1.53
+ $X2=5.28 $Y2=1.53
r288 140 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.665
+ $X2=4.635 $Y2=1.665
r289 139 141 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=4.635 $Y=1.53
+ $X2=4.85 $Y2=1.53
r290 139 140 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.635
+ $Y=1.5 $X2=4.635 $Y2=1.5
r291 137 139 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=4.42 $Y=1.53
+ $X2=4.635 $Y2=1.53
r292 136 137 61.3195 $w=3.9e-07 $l=4.3e-07 $layer=POLY_cond $X=3.99 $Y=1.53
+ $X2=4.42 $Y2=1.53
r293 134 136 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=3.775 $Y=1.53
+ $X2=3.99 $Y2=1.53
r294 134 135 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=1.5 $X2=3.775 $Y2=1.5
r295 132 134 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=3.56 $Y=1.53
+ $X2=3.775 $Y2=1.53
r296 131 132 61.3195 $w=3.9e-07 $l=4.3e-07 $layer=POLY_cond $X=3.13 $Y=1.53
+ $X2=3.56 $Y2=1.53
r297 130 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.915 $Y=1.665
+ $X2=2.915 $Y2=1.665
r298 129 131 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=2.915 $Y=1.53
+ $X2=3.13 $Y2=1.53
r299 129 130 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.5 $X2=2.915 $Y2=1.5
r300 127 129 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=2.7 $Y=1.53
+ $X2=2.915 $Y2=1.53
r301 126 127 61.3195 $w=3.9e-07 $l=4.3e-07 $layer=POLY_cond $X=2.27 $Y=1.53
+ $X2=2.7 $Y2=1.53
r302 125 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.055 $Y=1.665
+ $X2=2.055 $Y2=1.665
r303 124 126 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=2.055 $Y=1.53
+ $X2=2.27 $Y2=1.53
r304 124 125 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=1.5 $X2=2.055 $Y2=1.5
r305 122 124 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=1.84 $Y=1.53
+ $X2=2.055 $Y2=1.53
r306 121 122 61.3195 $w=3.9e-07 $l=4.3e-07 $layer=POLY_cond $X=1.41 $Y=1.53
+ $X2=1.84 $Y2=1.53
r307 120 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.195 $Y=1.665
+ $X2=1.195 $Y2=1.665
r308 119 121 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=1.195 $Y=1.53
+ $X2=1.41 $Y2=1.53
r309 119 120 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.5 $X2=1.195 $Y2=1.5
r310 117 119 30.6598 $w=3.9e-07 $l=2.15e-07 $layer=POLY_cond $X=0.98 $Y=1.53
+ $X2=1.195 $Y2=1.53
r311 115 117 61.3195 $w=3.9e-07 $l=4.3e-07 $layer=POLY_cond $X=0.55 $Y=1.53
+ $X2=0.98 $Y2=1.53
r312 113 177 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=3.775 $Y=1.665
+ $X2=4.635 $Y2=1.665
r313 113 167 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=3.775 $Y=1.665
+ $X2=2.915 $Y2=1.665
r314 113 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.775 $Y=1.665
+ $X2=3.775 $Y2=1.665
r315 110 152 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=7 $Y=1.725 $X2=7
+ $Y2=1.53
r316 110 112 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7 $Y=1.725 $X2=7
+ $Y2=2.465
r317 106 152 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=7 $Y=1.335 $X2=7
+ $Y2=1.53
r318 106 108 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7 $Y=1.335 $X2=7
+ $Y2=0.655
r319 103 151 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=6.57 $Y=1.725
+ $X2=6.57 $Y2=1.53
r320 103 105 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.57 $Y=1.725
+ $X2=6.57 $Y2=2.465
r321 99 151 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=6.57 $Y=1.335
+ $X2=6.57 $Y2=1.53
r322 99 101 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.57 $Y=1.335
+ $X2=6.57 $Y2=0.655
r323 96 147 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=6.14 $Y=1.725
+ $X2=6.14 $Y2=1.53
r324 96 98 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.14 $Y=1.725
+ $X2=6.14 $Y2=2.465
r325 92 147 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=6.14 $Y=1.335
+ $X2=6.14 $Y2=1.53
r326 92 94 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.14 $Y=1.335
+ $X2=6.14 $Y2=0.655
r327 89 146 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=5.71 $Y=1.725
+ $X2=5.71 $Y2=1.53
r328 89 91 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.71 $Y=1.725
+ $X2=5.71 $Y2=2.465
r329 85 146 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=5.71 $Y=1.335
+ $X2=5.71 $Y2=1.53
r330 85 87 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.71 $Y=1.335
+ $X2=5.71 $Y2=0.655
r331 82 142 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=5.28 $Y=1.725
+ $X2=5.28 $Y2=1.53
r332 82 84 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.28 $Y=1.725
+ $X2=5.28 $Y2=2.465
r333 78 142 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=5.28 $Y=1.335
+ $X2=5.28 $Y2=1.53
r334 78 80 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.28 $Y=1.335
+ $X2=5.28 $Y2=0.655
r335 75 141 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.85 $Y=1.725
+ $X2=4.85 $Y2=1.53
r336 75 77 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.85 $Y=1.725
+ $X2=4.85 $Y2=2.465
r337 71 141 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.85 $Y=1.335
+ $X2=4.85 $Y2=1.53
r338 71 73 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.85 $Y=1.335
+ $X2=4.85 $Y2=0.655
r339 68 137 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.42 $Y=1.725
+ $X2=4.42 $Y2=1.53
r340 68 70 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.42 $Y=1.725
+ $X2=4.42 $Y2=2.465
r341 64 137 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.42 $Y=1.335
+ $X2=4.42 $Y2=1.53
r342 64 66 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.42 $Y=1.335
+ $X2=4.42 $Y2=0.655
r343 61 136 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.99 $Y=1.725
+ $X2=3.99 $Y2=1.53
r344 61 63 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.99 $Y=1.725
+ $X2=3.99 $Y2=2.465
r345 57 136 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.99 $Y=1.335
+ $X2=3.99 $Y2=1.53
r346 57 59 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.99 $Y=1.335
+ $X2=3.99 $Y2=0.655
r347 54 132 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.56 $Y=1.725
+ $X2=3.56 $Y2=1.53
r348 54 56 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.56 $Y=1.725
+ $X2=3.56 $Y2=2.465
r349 50 132 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.56 $Y=1.335
+ $X2=3.56 $Y2=1.53
r350 50 52 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.56 $Y=1.335
+ $X2=3.56 $Y2=0.655
r351 47 131 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.13 $Y=1.725
+ $X2=3.13 $Y2=1.53
r352 47 49 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.13 $Y=1.725
+ $X2=3.13 $Y2=2.465
r353 43 131 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.13 $Y=1.335
+ $X2=3.13 $Y2=1.53
r354 43 45 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.13 $Y=1.335
+ $X2=3.13 $Y2=0.655
r355 40 127 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.7 $Y=1.725
+ $X2=2.7 $Y2=1.53
r356 40 42 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.7 $Y=1.725
+ $X2=2.7 $Y2=2.465
r357 36 127 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.7 $Y=1.335
+ $X2=2.7 $Y2=1.53
r358 36 38 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.7 $Y=1.335
+ $X2=2.7 $Y2=0.655
r359 33 126 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.27 $Y=1.725
+ $X2=2.27 $Y2=1.53
r360 33 35 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.27 $Y=1.725
+ $X2=2.27 $Y2=2.465
r361 29 126 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.27 $Y=1.335
+ $X2=2.27 $Y2=1.53
r362 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.27 $Y=1.335
+ $X2=2.27 $Y2=0.655
r363 26 122 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.84 $Y=1.725
+ $X2=1.84 $Y2=1.53
r364 26 28 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.84 $Y=1.725
+ $X2=1.84 $Y2=2.465
r365 22 122 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.84 $Y=1.335
+ $X2=1.84 $Y2=1.53
r366 22 24 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.84 $Y=1.335
+ $X2=1.84 $Y2=0.655
r367 19 121 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.41 $Y=1.725
+ $X2=1.41 $Y2=1.53
r368 19 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.41 $Y=1.725
+ $X2=1.41 $Y2=2.465
r369 15 121 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.41 $Y=1.335
+ $X2=1.41 $Y2=1.53
r370 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.41 $Y=1.335
+ $X2=1.41 $Y2=0.655
r371 12 117 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.98 $Y=1.725
+ $X2=0.98 $Y2=1.53
r372 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.98 $Y=1.725
+ $X2=0.98 $Y2=2.465
r373 8 117 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.98 $Y=1.335
+ $X2=0.98 $Y2=1.53
r374 8 10 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.98 $Y=1.335
+ $X2=0.98 $Y2=0.655
r375 5 115 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.55 $Y=1.725
+ $X2=0.55 $Y2=1.53
r376 5 7 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.55 $Y=1.725
+ $X2=0.55 $Y2=2.465
r377 1 115 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.55 $Y=1.335
+ $X2=0.55 $Y2=1.53
r378 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.55 $Y=1.335
+ $X2=0.55 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__INV_16%VPB 1 2 3 4 5 6 7 8 9 28 30 36 42 48 54 58 62
+ 68 74 80 85 86 88 89 90 91 93 94 95 96 97 98 100 115 129 134 137 140
r152 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r153 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r155 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r156 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r157 126 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r158 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r159 123 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r160 123 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r161 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r162 120 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.625 $Y=3.33
+ $X2=5.495 $Y2=3.33
r163 120 122 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.625 $Y=3.33
+ $X2=6 $Y2=3.33
r164 119 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r165 119 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r166 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r167 116 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.765 $Y=3.33
+ $X2=4.635 $Y2=3.33
r168 116 118 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.765 $Y=3.33
+ $X2=5.04 $Y2=3.33
r169 115 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.365 $Y=3.33
+ $X2=5.495 $Y2=3.33
r170 115 118 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.365 $Y=3.33
+ $X2=5.04 $Y2=3.33
r171 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r172 111 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r173 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r174 108 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r175 108 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r176 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r177 105 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.195 $Y2=3.33
r178 105 107 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.68 $Y2=3.33
r179 104 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r180 104 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r181 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r182 101 131 4.32323 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r183 101 103 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.72 $Y2=3.33
r184 100 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.195 $Y2=3.33
r185 100 103 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r186 98 138 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r187 98 114 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r188 96 125 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.085 $Y=3.33
+ $X2=6.96 $Y2=3.33
r189 96 97 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.085 $Y=3.33
+ $X2=7.232 $Y2=3.33
r190 95 128 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=7.38 $Y=3.33 $X2=7.44
+ $Y2=3.33
r191 95 97 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.38 $Y=3.33
+ $X2=7.232 $Y2=3.33
r192 93 122 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.225 $Y=3.33
+ $X2=6 $Y2=3.33
r193 93 94 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.225 $Y=3.33
+ $X2=6.355 $Y2=3.33
r194 92 125 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=6.485 $Y=3.33
+ $X2=6.96 $Y2=3.33
r195 92 94 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.485 $Y=3.33
+ $X2=6.355 $Y2=3.33
r196 90 113 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.6 $Y2=3.33
r197 90 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.775 $Y2=3.33
r198 88 110 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.785 $Y=3.33
+ $X2=2.64 $Y2=3.33
r199 88 89 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.785 $Y=3.33
+ $X2=2.915 $Y2=3.33
r200 87 113 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.045 $Y=3.33
+ $X2=3.6 $Y2=3.33
r201 87 89 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.045 $Y=3.33
+ $X2=2.915 $Y2=3.33
r202 85 107 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.925 $Y=3.33
+ $X2=1.68 $Y2=3.33
r203 85 86 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.925 $Y=3.33
+ $X2=2.055 $Y2=3.33
r204 84 110 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=2.64 $Y2=3.33
r205 84 86 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=2.055 $Y2=3.33
r206 80 83 31.6434 $w=2.93e-07 $l=8.1e-07 $layer=LI1_cond $X=7.232 $Y=2.085
+ $X2=7.232 $Y2=2.895
r207 78 97 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.232 $Y=3.245
+ $X2=7.232 $Y2=3.33
r208 78 83 13.6731 $w=2.93e-07 $l=3.5e-07 $layer=LI1_cond $X=7.232 $Y=3.245
+ $X2=7.232 $Y2=2.895
r209 74 77 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=6.355 $Y=2.085
+ $X2=6.355 $Y2=2.895
r210 72 94 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.355 $Y=3.245
+ $X2=6.355 $Y2=3.33
r211 72 77 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=6.355 $Y=3.245
+ $X2=6.355 $Y2=2.895
r212 68 71 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=5.495 $Y=2.085
+ $X2=5.495 $Y2=2.895
r213 66 140 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=3.245
+ $X2=5.495 $Y2=3.33
r214 66 71 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=5.495 $Y=3.245
+ $X2=5.495 $Y2=2.895
r215 62 65 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=4.635 $Y=2.085
+ $X2=4.635 $Y2=2.895
r216 60 137 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.635 $Y=3.245
+ $X2=4.635 $Y2=3.33
r217 60 65 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=4.635 $Y=3.245
+ $X2=4.635 $Y2=2.895
r218 59 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.775 $Y2=3.33
r219 58 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.505 $Y=3.33
+ $X2=4.635 $Y2=3.33
r220 58 59 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.505 $Y=3.33
+ $X2=3.905 $Y2=3.33
r221 54 57 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=3.775 $Y=2.085
+ $X2=3.775 $Y2=2.895
r222 52 91 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=3.245
+ $X2=3.775 $Y2=3.33
r223 52 57 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=3.775 $Y=3.245
+ $X2=3.775 $Y2=2.895
r224 48 51 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=2.915 $Y=2.085
+ $X2=2.915 $Y2=2.895
r225 46 89 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=3.33
r226 46 51 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=2.895
r227 42 45 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=2.055 $Y=2.085
+ $X2=2.055 $Y2=2.895
r228 40 86 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=3.33
r229 40 45 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=2.895
r230 36 39 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=1.195 $Y=2.085
+ $X2=1.195 $Y2=2.895
r231 34 134 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.195 $Y2=3.33
r232 34 39 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.195 $Y2=2.895
r233 30 33 31.6434 $w=2.93e-07 $l=8.1e-07 $layer=LI1_cond $X=0.317 $Y=2.085
+ $X2=0.317 $Y2=2.895
r234 28 131 3.15429 $w=2.95e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.317 $Y=3.245
+ $X2=0.232 $Y2=3.33
r235 28 33 13.6731 $w=2.93e-07 $l=3.5e-07 $layer=LI1_cond $X=0.317 $Y=3.245
+ $X2=0.317 $Y2=2.895
r236 9 83 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=7.075
+ $Y=1.835 $X2=7.215 $Y2=2.895
r237 9 80 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=7.075
+ $Y=1.835 $X2=7.215 $Y2=2.085
r238 8 77 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=1.835 $X2=6.355 $Y2=2.895
r239 8 74 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=1.835 $X2=6.355 $Y2=2.085
r240 7 71 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.835 $X2=5.495 $Y2=2.895
r241 7 68 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.835 $X2=5.495 $Y2=2.085
r242 6 65 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=4.495
+ $Y=1.835 $X2=4.635 $Y2=2.895
r243 6 62 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=4.495
+ $Y=1.835 $X2=4.635 $Y2=2.085
r244 5 57 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.835 $X2=3.775 $Y2=2.895
r245 5 54 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.835 $X2=3.775 $Y2=2.085
r246 4 51 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.915 $Y2=2.895
r247 4 48 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.915 $Y2=2.085
r248 3 45 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.895
r249 3 42 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.085
r250 2 39 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.835 $X2=1.195 $Y2=2.895
r251 2 36 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.835 $X2=1.195 $Y2=2.085
r252 1 33 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=1.835 $X2=0.335 $Y2=2.895
r253 1 30 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=1.835 $X2=0.335 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__INV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 49
+ 52 62 72 82 92 102 112 122 126
r180 125 129 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=6.785 $Y=2.035
+ $X2=6.785 $Y2=2.885
r181 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.785 $Y=2.035
+ $X2=6.785 $Y2=2.035
r182 122 125 69.3682 $w=2.58e-07 $l=1.565e-06 $layer=LI1_cond $X=6.785 $Y=0.47
+ $X2=6.785 $Y2=2.035
r183 116 126 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=5.925 $Y=2.035
+ $X2=6.785 $Y2=2.035
r184 115 119 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=5.925 $Y=2.035
+ $X2=5.925 $Y2=2.885
r185 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.925 $Y=2.035
+ $X2=5.925 $Y2=2.035
r186 112 115 69.3682 $w=2.58e-07 $l=1.565e-06 $layer=LI1_cond $X=5.925 $Y=0.47
+ $X2=5.925 $Y2=2.035
r187 106 116 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=5.065 $Y=2.035
+ $X2=5.925 $Y2=2.035
r188 105 109 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=5.065 $Y=2.035
+ $X2=5.065 $Y2=2.885
r189 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.065 $Y=2.035
+ $X2=5.065 $Y2=2.035
r190 102 105 69.3682 $w=2.58e-07 $l=1.565e-06 $layer=LI1_cond $X=5.065 $Y=0.47
+ $X2=5.065 $Y2=2.035
r191 96 106 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=4.205 $Y=2.035
+ $X2=5.065 $Y2=2.035
r192 95 99 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=4.205 $Y=2.035
+ $X2=4.205 $Y2=2.885
r193 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.205 $Y=2.035
+ $X2=4.205 $Y2=2.035
r194 92 95 69.3682 $w=2.58e-07 $l=1.565e-06 $layer=LI1_cond $X=4.205 $Y=0.47
+ $X2=4.205 $Y2=2.035
r195 85 89 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=3.345 $Y=2.035
+ $X2=3.345 $Y2=2.885
r196 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.345 $Y=2.035
+ $X2=3.345 $Y2=2.035
r197 82 85 69.3682 $w=2.58e-07 $l=1.565e-06 $layer=LI1_cond $X=3.345 $Y=0.47
+ $X2=3.345 $Y2=2.035
r198 76 86 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=2.485 $Y=2.035
+ $X2=3.345 $Y2=2.035
r199 75 79 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=2.485 $Y=2.035
+ $X2=2.485 $Y2=2.885
r200 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.485 $Y=2.035
+ $X2=2.485 $Y2=2.035
r201 72 75 69.3682 $w=2.58e-07 $l=1.565e-06 $layer=LI1_cond $X=2.485 $Y=0.47
+ $X2=2.485 $Y2=2.035
r202 66 76 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=1.625 $Y=2.035
+ $X2=2.485 $Y2=2.035
r203 65 69 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=1.625 $Y=2.035
+ $X2=1.625 $Y2=2.885
r204 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.625 $Y=2.035
+ $X2=1.625 $Y2=2.035
r205 62 65 69.3682 $w=2.58e-07 $l=1.565e-06 $layer=LI1_cond $X=1.625 $Y=0.47
+ $X2=1.625 $Y2=2.035
r206 56 66 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=0.765 $Y=2.035
+ $X2=1.625 $Y2=2.035
r207 55 59 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=0.765 $Y=2.035
+ $X2=0.765 $Y2=2.885
r208 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.765 $Y=2.035
+ $X2=0.765 $Y2=2.035
r209 52 55 69.3682 $w=2.58e-07 $l=1.565e-06 $layer=LI1_cond $X=0.765 $Y=0.47
+ $X2=0.765 $Y2=2.035
r210 49 96 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=3.775 $Y=2.035
+ $X2=4.205 $Y2=2.035
r211 49 86 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=3.775 $Y=2.035
+ $X2=3.345 $Y2=2.035
r212 16 129 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=6.645
+ $Y=1.835 $X2=6.785 $Y2=2.885
r213 16 125 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.645
+ $Y=1.835 $X2=6.785 $Y2=2.045
r214 15 119 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.835 $X2=5.925 $Y2=2.885
r215 15 115 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.835 $X2=5.925 $Y2=2.045
r216 14 109 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.835 $X2=5.065 $Y2=2.885
r217 14 105 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.835 $X2=5.065 $Y2=2.045
r218 13 99 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.835 $X2=4.205 $Y2=2.885
r219 13 95 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.835 $X2=4.205 $Y2=2.045
r220 12 89 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.835 $X2=3.345 $Y2=2.885
r221 12 85 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.835 $X2=3.345 $Y2=2.045
r222 11 79 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.835 $X2=2.485 $Y2=2.885
r223 11 75 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.835 $X2=2.485 $Y2=2.045
r224 10 69 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=2.885
r225 10 65 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=2.045
r226 9 59 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.835 $X2=0.765 $Y2=2.885
r227 9 55 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.835 $X2=0.765 $Y2=2.045
r228 8 122 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=6.645
+ $Y=0.235 $X2=6.785 $Y2=0.47
r229 7 112 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.785
+ $Y=0.235 $X2=5.925 $Y2=0.47
r230 6 102 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.925
+ $Y=0.235 $X2=5.065 $Y2=0.47
r231 5 92 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.065
+ $Y=0.235 $X2=4.205 $Y2=0.47
r232 4 82 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=3.205
+ $Y=0.235 $X2=3.345 $Y2=0.47
r233 3 72 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=2.345
+ $Y=0.235 $X2=2.485 $Y2=0.47
r234 2 62 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.235 $X2=1.625 $Y2=0.47
r235 1 52 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=0.625
+ $Y=0.235 $X2=0.765 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__INV_16%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 48
+ 52 56 60 64 67 68 70 71 72 73 75 76 77 78 79 80 82 97 111 116 119 122
r121 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r122 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r123 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r124 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r125 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r126 108 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r127 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r128 105 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r129 105 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r130 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r131 102 122 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.625 $Y=0
+ $X2=5.495 $Y2=0
r132 102 104 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.625 $Y=0 $X2=6
+ $Y2=0
r133 101 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r134 101 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r135 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r136 98 119 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=4.635 $Y2=0
r137 98 100 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=5.04 $Y2=0
r138 97 122 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.365 $Y=0
+ $X2=5.495 $Y2=0
r139 97 100 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.365 $Y=0
+ $X2=5.04 $Y2=0
r140 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r141 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r142 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r143 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r144 90 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r145 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r146 87 116 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.325 $Y=0
+ $X2=1.195 $Y2=0
r147 87 89 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.325 $Y=0
+ $X2=1.68 $Y2=0
r148 86 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r149 86 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r150 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r151 83 113 4.32323 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=0
+ $X2=0.232 $Y2=0
r152 83 85 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.465 $Y=0
+ $X2=0.72 $Y2=0
r153 82 116 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.065 $Y=0
+ $X2=1.195 $Y2=0
r154 82 85 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r155 80 120 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.56 $Y2=0
r156 80 96 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r157 78 107 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=6.96 $Y2=0
r158 78 79 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=7.232 $Y2=0
r159 77 110 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=7.38 $Y=0 $X2=7.44
+ $Y2=0
r160 77 79 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.38 $Y=0 $X2=7.232
+ $Y2=0
r161 75 104 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6
+ $Y2=0
r162 75 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.355
+ $Y2=0
r163 74 107 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=6.485 $Y=0
+ $X2=6.96 $Y2=0
r164 74 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.485 $Y=0 $X2=6.355
+ $Y2=0
r165 72 95 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.6
+ $Y2=0
r166 72 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.775
+ $Y2=0
r167 70 92 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.785 $Y=0
+ $X2=2.64 $Y2=0
r168 70 71 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.785 $Y=0 $X2=2.915
+ $Y2=0
r169 69 95 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.6
+ $Y2=0
r170 69 71 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=2.915
+ $Y2=0
r171 67 89 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=1.68
+ $Y2=0
r172 67 68 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=2.055
+ $Y2=0
r173 66 92 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=2.64 $Y2=0
r174 66 68 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.055
+ $Y2=0
r175 62 79 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.232 $Y=0.085
+ $X2=7.232 $Y2=0
r176 62 64 15.0404 $w=2.93e-07 $l=3.85e-07 $layer=LI1_cond $X=7.232 $Y=0.085
+ $X2=7.232 $Y2=0.47
r177 58 76 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.355 $Y=0.085
+ $X2=6.355 $Y2=0
r178 58 60 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=6.355 $Y=0.085
+ $X2=6.355 $Y2=0.47
r179 54 122 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=0.085
+ $X2=5.495 $Y2=0
r180 54 56 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=5.495 $Y=0.085
+ $X2=5.495 $Y2=0.47
r181 50 119 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.635 $Y=0.085
+ $X2=4.635 $Y2=0
r182 50 52 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=4.635 $Y=0.085
+ $X2=4.635 $Y2=0.47
r183 49 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.905 $Y=0 $X2=3.775
+ $Y2=0
r184 48 119 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.505 $Y=0
+ $X2=4.635 $Y2=0
r185 48 49 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.505 $Y=0 $X2=3.905
+ $Y2=0
r186 44 73 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=0.085
+ $X2=3.775 $Y2=0
r187 44 46 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=3.775 $Y=0.085
+ $X2=3.775 $Y2=0.47
r188 40 71 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0
r189 40 42 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.47
r190 36 68 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0
r191 36 38 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0.47
r192 32 116 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0
r193 32 34 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0.47
r194 28 113 3.15429 $w=2.95e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.317 $Y=0.085
+ $X2=0.232 $Y2=0
r195 28 30 15.0404 $w=2.93e-07 $l=3.85e-07 $layer=LI1_cond $X=0.317 $Y=0.085
+ $X2=0.317 $Y2=0.47
r196 9 64 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=7.075
+ $Y=0.235 $X2=7.215 $Y2=0.47
r197 8 60 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=6.215
+ $Y=0.235 $X2=6.355 $Y2=0.47
r198 7 56 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.355
+ $Y=0.235 $X2=5.495 $Y2=0.47
r199 6 52 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.495
+ $Y=0.235 $X2=4.635 $Y2=0.47
r200 5 46 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=3.635
+ $Y=0.235 $X2=3.775 $Y2=0.47
r201 4 42 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=2.775
+ $Y=0.235 $X2=2.915 $Y2=0.47
r202 3 38 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=1.915
+ $Y=0.235 $X2=2.055 $Y2=0.47
r203 2 34 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=1.055
+ $Y=0.235 $X2=1.195 $Y2=0.47
r204 1 30 91 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.235 $X2=0.335 $Y2=0.47
.ends

