* File: sky130_fd_sc_lp__o22a_0.pex.spice
* Created: Fri Aug 28 11:09:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22A_0%A_80_313# 1 2 8 11 15 17 20 21 24 25 26 27 31
+ 34 35 36 38 41 44 49
c125 36 0 6.30536e-20 $X=3.075 $Y=1.67
c126 27 0 9.6968e-20 $X=2.905 $Y=1.12
c127 26 0 1.12607e-19 $X=0.765 $Y=2.52
c128 17 0 1.77161e-19 $X=0.572 $Y=2.235
c129 15 0 4.9202e-21 $X=0.575 $Y=0.835
r130 44 46 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.02 $Y=0.89
+ $X2=2.02 $Y2=1.12
r131 39 41 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.58 $Y=2.15 $X2=0.68
+ $Y2=2.15
r132 37 38 36.7894 $w=2.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.642 $Y=1.755
+ $X2=3.642 $Y2=2.435
r133 35 37 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=3.54 $Y=1.67
+ $X2=3.642 $Y2=1.755
r134 35 36 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.54 $Y=1.67
+ $X2=3.075 $Y2=1.67
r135 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=1.585
+ $X2=3.075 $Y2=1.67
r136 33 34 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.99 $Y=1.205
+ $X2=2.99 $Y2=1.585
r137 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.555 $Y=2.52
+ $X2=2.39 $Y2=2.52
r138 31 38 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=3.54 $Y=2.52
+ $X2=3.642 $Y2=2.435
r139 31 32 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=3.54 $Y=2.52
+ $X2=2.555 $Y2=2.52
r140 28 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=1.12
+ $X2=2.02 $Y2=1.12
r141 27 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=1.12
+ $X2=2.99 $Y2=1.205
r142 27 28 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.905 $Y=1.12
+ $X2=2.185 $Y2=1.12
r143 25 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=2.52
+ $X2=2.39 $Y2=2.52
r144 25 26 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.225 $Y=2.52
+ $X2=0.765 $Y2=2.52
r145 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=2.435
+ $X2=0.765 $Y2=2.52
r146 23 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.235
+ $X2=0.68 $Y2=2.15
r147 23 24 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.68 $Y=2.235
+ $X2=0.68 $Y2=2.435
r148 21 51 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.572 $Y=1.73
+ $X2=0.572 $Y2=1.565
r149 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.73 $X2=0.58 $Y2=1.73
r150 18 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.58 $Y=2.065
+ $X2=0.58 $Y2=2.15
r151 18 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.58 $Y=2.065
+ $X2=0.58 $Y2=1.73
r152 15 51 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.575 $Y=0.835
+ $X2=0.575 $Y2=1.565
r153 11 17 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=2.765
+ $X2=0.475 $Y2=2.235
r154 8 17 47.5363 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=0.572 $Y=2.063
+ $X2=0.572 $Y2=2.235
r155 7 21 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=0.572 $Y=1.737
+ $X2=0.572 $Y2=1.73
r156 7 8 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=0.572 $Y=1.737
+ $X2=0.572 $Y2=2.063
r157 2 49 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.25
+ $Y=2.445 $X2=2.39 $Y2=2.59
r158 1 44 182 $w=1.7e-07 $l=3.35596e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.625 $X2=2.02 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_0%A1 1 3 6 8 11 12 13 15 16 20 21 22 31 36 37
+ 39
c85 36 0 8.73193e-21 $X=1.205 $Y=0.5
c86 16 0 6.30536e-20 $X=3.225 $Y=2.1
c87 15 0 9.29322e-20 $X=3.225 $Y=2.1
c88 1 0 1.51092e-19 $X=1.355 $Y=0.515
r89 36 39 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=1.205 $Y=0.5
+ $X2=1.205 $Y2=0.555
r90 28 31 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.16 $Y=0.35
+ $X2=1.355 $Y2=0.35
r91 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=0.35 $X2=1.16 $Y2=0.35
r92 22 37 3.39854 $w=1.8e-07 $l=1.4e-07 $layer=LI1_cond $X=1.142 $Y=1.282
+ $X2=1.205 $Y2=1.17
r93 21 37 15.096 $w=1.78e-07 $l=2.45e-07 $layer=LI1_cond $X=1.205 $Y=0.925
+ $X2=1.205 $Y2=1.17
r94 20 36 2.9051 $w=3.21e-07 $l=5.19615e-08 $layer=LI1_cond $X=1.16 $Y=0.485
+ $X2=1.205 $Y2=0.5
r95 20 29 5.13084 $w=3.21e-07 $l=1.35e-07 $layer=LI1_cond $X=1.16 $Y=0.485
+ $X2=1.16 $Y2=0.35
r96 20 21 21.8737 $w=1.78e-07 $l=3.55e-07 $layer=LI1_cond $X=1.205 $Y=0.57
+ $X2=1.205 $Y2=0.925
r97 20 39 0.924242 $w=1.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.205 $Y=0.57
+ $X2=1.205 $Y2=0.555
r98 16 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=2.1
+ $X2=3.225 $Y2=2.265
r99 15 18 2.97405 $w=3.08e-07 $l=8e-08 $layer=LI1_cond $X=3.215 $Y=2.1 $X2=3.215
+ $Y2=2.18
r100 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=2.1 $X2=3.225 $Y2=2.1
r101 12 18 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.06 $Y=2.18
+ $X2=3.215 $Y2=2.18
r102 12 13 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=3.06 $Y=2.18
+ $X2=1.685 $Y2=2.18
r103 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=2.095
+ $X2=1.685 $Y2=2.18
r104 10 11 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.6 $Y=1.395 $X2=1.6
+ $Y2=2.095
r105 9 22 3.41796 $w=1.8e-07 $l=1.64098e-07 $layer=LI1_cond $X=1.295 $Y=1.305
+ $X2=1.142 $Y2=1.282
r106 8 10 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.515 $Y=1.305
+ $X2=1.6 $Y2=1.395
r107 8 9 13.5556 $w=1.78e-07 $l=2.2e-07 $layer=LI1_cond $X=1.515 $Y=1.305
+ $X2=1.295 $Y2=1.305
r108 6 35 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.135 $Y=2.765
+ $X2=3.135 $Y2=2.265
r109 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=0.515
+ $X2=1.355 $Y2=0.35
r110 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.355 $Y=0.515
+ $X2=1.355 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_0%B1 3 7 9 10 11 12
c48 11 0 1.90671e-19 $X=1.2 $Y=1.665
c49 3 0 1.0078e-19 $X=1.785 $Y=0.835
r50 11 12 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.2
+ $Y2=2.035
r51 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.24
+ $Y=1.73 $X2=1.24 $Y2=1.73
r52 9 16 37.5319 $w=6.7e-07 $l=4.7e-07 $layer=POLY_cond $X=1.71 $Y=1.9 $X2=1.24
+ $Y2=1.9
r53 9 10 11.9686 $w=6.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.71 $Y=1.9 $X2=1.785
+ $Y2=1.9
r54 5 10 56.3093 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.785 $Y=2.235
+ $X2=1.785 $Y2=1.9
r55 5 7 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.785 $Y=2.235
+ $X2=1.785 $Y2=2.765
r56 1 10 56.3093 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.785 $Y=1.565
+ $X2=1.785 $Y2=1.9
r57 1 3 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.785 $Y=1.565
+ $X2=1.785 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_0%B2 3 7 11 12 13 14 18
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.265
+ $Y=1.47 $X2=2.265 $Y2=1.47
r47 14 19 8.3061 $w=5.38e-07 $l=3.75e-07 $layer=LI1_cond $X=2.64 $Y=1.655
+ $X2=2.265 $Y2=1.655
r48 13 19 2.32571 $w=5.38e-07 $l=1.05e-07 $layer=LI1_cond $X=2.16 $Y=1.655
+ $X2=2.265 $Y2=1.655
r49 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.265 $Y=1.81
+ $X2=2.265 $Y2=1.47
r50 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.81
+ $X2=2.265 $Y2=1.975
r51 10 18 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.305
+ $X2=2.265 $Y2=1.47
r52 7 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.235 $Y=0.835 $X2=2.235
+ $Y2=1.305
r53 3 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.175 $Y=2.765
+ $X2=2.175 $Y2=1.975
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_0%A2 1 3 4 6 8 11 14 15 18
c46 18 0 9.29322e-20 $X=3.42 $Y=1.32
c47 4 0 9.20945e-20 $X=2.745 $Y=1.155
r48 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.32 $X2=3.42 $Y2=1.32
r49 15 19 6.91466 $w=2.98e-07 $l=1.8e-07 $layer=LI1_cond $X=3.6 $Y=1.265
+ $X2=3.42 $Y2=1.265
r50 13 18 104.917 $w=3.3e-07 $l=6e-07 $layer=POLY_cond $X=2.82 $Y=1.32 $X2=3.42
+ $Y2=1.32
r51 13 14 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.82 $Y=1.32
+ $X2=2.745 $Y2=1.32
r52 9 11 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.605 $Y=2.26
+ $X2=2.745 $Y2=2.26
r53 8 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.745 $Y=2.185
+ $X2=2.745 $Y2=2.26
r54 7 14 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.485
+ $X2=2.745 $Y2=1.32
r55 7 8 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=2.745 $Y=1.485 $X2=2.745
+ $Y2=2.185
r56 4 14 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.155
+ $X2=2.745 $Y2=1.32
r57 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.745 $Y=1.155
+ $X2=2.745 $Y2=0.835
r58 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.605 $Y=2.335
+ $X2=2.605 $Y2=2.26
r59 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.605 $Y=2.335
+ $X2=2.605 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_0%X 1 2 7 8 9 10 11 12 32 42
r24 33 47 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=0.255 $Y=2.595
+ $X2=0.255 $Y2=2.59
r25 32 45 0.960369 $w=2.38e-07 $l=2e-08 $layer=LI1_cond $X=0.205 $Y=2.405
+ $X2=0.205 $Y2=2.425
r26 21 37 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.205 $Y=0.935
+ $X2=0.205 $Y2=0.77
r27 12 33 6.10117 $w=3.38e-07 $l=1.8e-07 $layer=LI1_cond $X=0.255 $Y=2.775
+ $X2=0.255 $Y2=2.595
r28 11 47 4.50809 $w=3.38e-07 $l=1.33e-07 $layer=LI1_cond $X=0.255 $Y=2.457
+ $X2=0.255 $Y2=2.59
r29 11 45 2.0963 $w=3.38e-07 $l=3.2e-08 $layer=LI1_cond $X=0.255 $Y=2.457
+ $X2=0.255 $Y2=2.425
r30 11 32 1.58461 $w=2.38e-07 $l=3.3e-08 $layer=LI1_cond $X=0.205 $Y=2.372
+ $X2=0.205 $Y2=2.405
r31 10 11 16.1822 $w=2.38e-07 $l=3.37e-07 $layer=LI1_cond $X=0.205 $Y=2.035
+ $X2=0.205 $Y2=2.372
r32 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.205 $Y=1.665
+ $X2=0.205 $Y2=2.035
r33 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.205 $Y=1.295
+ $X2=0.205 $Y2=1.665
r34 7 42 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.24 $Y=0.77 $X2=0.36
+ $Y2=0.77
r35 7 37 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=0.77
+ $X2=0.205 $Y2=0.77
r36 7 8 15.51 $w=2.38e-07 $l=3.23e-07 $layer=LI1_cond $X=0.205 $Y=0.972
+ $X2=0.205 $Y2=1.295
r37 7 21 1.77668 $w=2.38e-07 $l=3.7e-08 $layer=LI1_cond $X=0.205 $Y=0.972
+ $X2=0.205 $Y2=0.935
r38 2 47 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.445 $X2=0.26 $Y2=2.59
r39 1 42 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.625 $X2=0.36 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_0%VPWR 1 2 9 11 15 17 18 19 25 34 35 42
r48 40 42 8.3611 $w=6.38e-07 $l=5.5e-08 $layer=LI1_cond $X=1.68 $Y=3.095
+ $X2=1.735 $Y2=3.095
r49 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 38 40 2.05576 $w=6.38e-07 $l=1.1e-07 $layer=LI1_cond $X=1.57 $Y=3.095
+ $X2=1.68 $Y2=3.095
r51 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r53 31 42 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=1.735 $Y2=3.33
r54 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 25 38 2.89675 $w=6.38e-07 $l=1.55e-07 $layer=LI1_cond $X=1.415 $Y=3.095
+ $X2=1.57 $Y2=3.095
r58 25 27 4.01808 $w=6.38e-07 $l=2.15e-07 $layer=LI1_cond $X=1.415 $Y=3.095
+ $X2=1.2 $Y2=3.095
r59 23 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 19 32 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 19 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 17 31 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.12 $Y2=3.33
r64 17 18 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.35 $Y2=3.33
r65 16 34 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.6 $Y2=3.33
r66 16 18 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.35 $Y2=3.33
r67 15 22 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.24 $Y2=3.33
r68 14 15 9.10865 $w=6.38e-07 $l=9.5e-08 $layer=LI1_cond $X=0.69 $Y=3.095
+ $X2=0.595 $Y2=3.095
r69 11 27 5.32629 $w=6.38e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=3.095
+ $X2=1.2 $Y2=3.095
r70 11 14 4.20496 $w=6.38e-07 $l=2.25e-07 $layer=LI1_cond $X=0.915 $Y=3.095
+ $X2=0.69 $Y2=3.095
r71 7 18 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=3.245 $X2=3.35
+ $Y2=3.33
r72 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.35 $Y=3.245
+ $X2=3.35 $Y2=2.89
r73 2 9 600 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=2.445 $X2=3.35 $Y2=2.89
r74 1 38 400 $w=1.7e-07 $l=1.2431e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.445 $X2=1.57 $Y2=2.94
r75 1 14 400 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.445 $X2=0.69 $Y2=2.94
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_0%VGND 1 2 10 13 18 20 22 32 33 36 39
r43 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r46 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r47 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.04
+ $Y2=0
r48 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.6
+ $Y2=0
r49 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r50 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r51 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r53 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 23 36 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.735
+ $Y2=0
r55 23 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.825 $Y=0 $X2=1.2
+ $Y2=0
r56 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=3.04
+ $Y2=0
r57 22 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.64
+ $Y2=0
r58 20 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r59 20 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r60 15 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.735 $Y=0.835
+ $X2=0.825 $Y2=0.835
r61 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0
r62 11 13 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0.77
r63 10 15 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=0.67
+ $X2=0.735 $Y2=0.835
r64 9 36 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0
r65 9 10 36.0455 $w=1.78e-07 $l=5.85e-07 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0.67
r66 2 13 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.625 $X2=3.04 $Y2=0.77
r67 1 18 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.625 $X2=0.825 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_0%A_286_125# 1 2 9 11 12 13
c24 12 0 1.37581e-19 $X=1.685 $Y=0.53
c25 11 0 9.20945e-20 $X=2.365 $Y=0.53
r26 13 16 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.53 $Y=0.53
+ $X2=2.53 $Y2=0.76
r27 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0.53
+ $X2=2.53 $Y2=0.53
r28 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.365 $Y=0.53
+ $X2=1.685 $Y2=0.53
r29 7 12 5.96496 $w=2.27e-07 $l=2.43875e-07 $layer=LI1_cond $X=1.575 $Y=0.725
+ $X2=1.685 $Y2=0.53
r30 7 9 5.76222 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=1.575 $Y=0.725
+ $X2=1.575 $Y2=0.835
r31 2 16 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.625 $X2=2.53 $Y2=0.76
r32 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.625 $X2=1.57 $Y2=0.835
.ends

