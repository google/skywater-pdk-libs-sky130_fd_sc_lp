* File: sky130_fd_sc_lp__decapkapwr_6.spice
* Created: Wed Sep  2 09:42:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__decapkapwr_6.pex.spice"
.subckt sky130_fd_sc_lp__decapkapwr_6  VNB VPB VGND KAPWR VPWR
* 
* KAPWR	KAPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_s N_KAPWR_M1001_g N_VGND_M1001_s VNB NSHORT L=2 W=1 AD=0.265
+ AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=0.5 SA=999999 SB=999999 A=2 P=6
+ MULT=1
MM1000 N_KAPWR_M1000_s N_VGND_M1000_g N_KAPWR_M1000_s VPB PHIGHVT L=2 W=1
+ AD=0.285 AS=0.275 PD=2.57 PS=2.55 NRD=0 NRS=1.9503 M=1 R=0.5 SA=999999
+ SB=999999 A=2 P=6 MULT=1
DX2_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__decapkapwr_6.pxi.spice"
*
.ends
*
*
