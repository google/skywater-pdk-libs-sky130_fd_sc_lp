* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_0 A0 A1 S VGND VNB VPB VPWR X
X0 a_89_200# A0 a_467_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_89_200# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_89_200# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 VPWR S a_509_99# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND S a_257_94# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_89_200# A1 a_423_515# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_423_515# a_509_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_257_94# A1 a_89_200# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_467_125# a_509_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR S a_227_491# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_227_491# A0 a_89_200# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND S a_509_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
