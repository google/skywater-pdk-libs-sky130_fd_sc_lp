* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__isobufsrc_2 A SLEEP VGND VNB VPB VPWR X
M1000 VGND SLEEP X VNB nshort w=840000u l=150000u
+  ad=1.0038e+12p pd=7.52e+06u as=4.704e+11p ps=4.48e+06u
M1001 VGND A a_40_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1002 a_283_367# a_40_131# X VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=3.528e+11p ps=3.08e+06u
M1003 VPWR A a_40_131# VPB phighvt w=420000u l=150000u
+  ad=7.14e+11p pd=6.32e+06u as=1.113e+11p ps=1.37e+06u
M1004 VGND a_40_131# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_40_131# a_283_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_40_131# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X SLEEP VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR SLEEP a_283_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_283_367# SLEEP VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
