# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a22oi_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a22oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 1.180000 1.845000 1.750000 ;
        RECT 1.585000 0.365000 1.810000 1.100000 ;
        RECT 1.585000 1.100000 1.845000 1.180000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015000 1.210000 2.795000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.210000 1.350000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.535000 1.750000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.693000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.705000 0.860000 1.415000 1.040000 ;
        RECT 0.705000 1.040000 0.875000 1.920000 ;
        RECT 0.705000 1.920000 2.245000 2.130000 ;
        RECT 0.705000 2.130000 1.045000 2.735000 ;
        RECT 1.205000 0.325000 1.415000 0.860000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.880000 0.085000 ;
        RECT 0.285000  0.085000 0.535000 1.040000 ;
        RECT 2.170000  0.085000 2.500000 0.995000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 2.880000 3.415000 ;
        RECT 1.630000 2.640000 2.300000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.285000 1.920000 0.535000 2.905000 ;
      RECT 0.285000 2.905000 1.460000 3.075000 ;
      RECT 1.215000 2.300000 2.730000 2.470000 ;
      RECT 1.215000 2.470000 1.460000 2.905000 ;
      RECT 2.415000 1.920000 2.730000 2.300000 ;
      RECT 2.470000 2.470000 2.730000 3.075000 ;
  END
END sky130_fd_sc_lp__a22oi_1
