* File: sky130_fd_sc_lp__or4b_1.pxi.spice
* Created: Fri Aug 28 11:25:38 2020
* 
x_PM_SKY130_FD_SC_LP__OR4B_1%D_N N_D_N_M1006_g N_D_N_M1005_g D_N D_N
+ N_D_N_c_72_n PM_SKY130_FD_SC_LP__OR4B_1%D_N
x_PM_SKY130_FD_SC_LP__OR4B_1%A_64_131# N_A_64_131#_M1006_s N_A_64_131#_M1005_s
+ N_A_64_131#_M1002_g N_A_64_131#_c_97_n N_A_64_131#_M1009_g N_A_64_131#_c_98_n
+ N_A_64_131#_c_102_n N_A_64_131#_c_99_n N_A_64_131#_c_100_n
+ PM_SKY130_FD_SC_LP__OR4B_1%A_64_131#
x_PM_SKY130_FD_SC_LP__OR4B_1%C N_C_c_145_n N_C_M1010_g N_C_c_146_n N_C_c_147_n
+ N_C_M1007_g C C C C N_C_c_152_n PM_SKY130_FD_SC_LP__OR4B_1%C
x_PM_SKY130_FD_SC_LP__OR4B_1%B N_B_M1011_g N_B_M1003_g N_B_c_197_n B B
+ N_B_c_199_n PM_SKY130_FD_SC_LP__OR4B_1%B
x_PM_SKY130_FD_SC_LP__OR4B_1%A N_A_M1000_g N_A_M1004_g A A A N_A_c_237_n
+ PM_SKY130_FD_SC_LP__OR4B_1%A
x_PM_SKY130_FD_SC_LP__OR4B_1%A_220_367# N_A_220_367#_M1002_d
+ N_A_220_367#_M1011_d N_A_220_367#_M1009_s N_A_220_367#_c_270_n
+ N_A_220_367#_M1001_g N_A_220_367#_M1008_g N_A_220_367#_c_272_n
+ N_A_220_367#_c_273_n N_A_220_367#_c_274_n N_A_220_367#_c_304_n
+ N_A_220_367#_c_275_n N_A_220_367#_c_280_n N_A_220_367#_c_291_n
+ N_A_220_367#_c_276_n N_A_220_367#_c_277_n
+ PM_SKY130_FD_SC_LP__OR4B_1%A_220_367#
x_PM_SKY130_FD_SC_LP__OR4B_1%VPWR N_VPWR_M1005_d N_VPWR_M1004_d N_VPWR_c_348_n
+ N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n
+ VPWR N_VPWR_c_354_n N_VPWR_c_347_n PM_SKY130_FD_SC_LP__OR4B_1%VPWR
x_PM_SKY130_FD_SC_LP__OR4B_1%X N_X_M1008_d N_X_M1001_d X X X X X X X N_X_c_387_n
+ X X N_X_c_391_n PM_SKY130_FD_SC_LP__OR4B_1%X
x_PM_SKY130_FD_SC_LP__OR4B_1%VGND N_VGND_M1006_d N_VGND_M1010_d N_VGND_M1000_d
+ N_VGND_c_404_n N_VGND_c_405_n N_VGND_c_406_n N_VGND_c_407_n N_VGND_c_408_n
+ N_VGND_c_409_n N_VGND_c_410_n VGND N_VGND_c_411_n N_VGND_c_412_n
+ N_VGND_c_413_n N_VGND_c_414_n PM_SKY130_FD_SC_LP__OR4B_1%VGND
cc_1 VNB N_D_N_M1006_g 0.0469463f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.865
cc_2 VNB D_N 0.0136354f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_3 VNB N_D_N_c_72_n 0.0192016f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.73
cc_4 VNB N_A_64_131#_M1002_g 0.0196427f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_5 VNB N_A_64_131#_c_97_n 0.0474312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_64_131#_c_98_n 0.020893f $X=-0.19 $Y=-0.245 $X2=0.477 $Y2=1.565
cc_7 VNB N_A_64_131#_c_99_n 9.84849e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_64_131#_c_100_n 0.0230472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C_c_145_n 0.0189395f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.565
cc_10 VNB N_C_c_146_n 0.0254851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_c_147_n 0.00771144f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.235
cc_12 VNB N_C_M1007_g 0.016693f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB C 0.00314404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_M1011_g 0.0283541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_197_n 0.00697213f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_16 VNB B 0.0119697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_c_199_n 0.0464063f $X=-0.19 $Y=-0.245 $X2=0.477 $Y2=1.565
cc_18 VNB N_A_M1000_g 0.0397827f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.865
cc_19 VNB N_A_220_367#_c_270_n 0.0413896f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_20 VNB N_A_220_367#_M1008_g 0.0283553f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.73
cc_21 VNB N_A_220_367#_c_272_n 0.00147461f $X=-0.19 $Y=-0.245 $X2=0.282
+ $Y2=1.665
cc_22 VNB N_A_220_367#_c_273_n 0.00332048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_220_367#_c_274_n 0.0137087f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.73
cc_24 VNB N_A_220_367#_c_275_n 0.0169902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_220_367#_c_276_n 0.00101194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_220_367#_c_277_n 0.00528547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_347_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB X 0.0296845f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_X_c_387_n 0.0290325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB X 0.0109066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_404_n 0.031188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_405_n 0.0217376f $X=-0.19 $Y=-0.245 $X2=0.477 $Y2=1.565
cc_33 VNB N_VGND_c_406_n 0.00681128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_407_n 0.0256816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_408_n 0.00442399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_409_n 0.020667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_410_n 0.00384695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_411_n 0.0257961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_412_n 0.0170749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_413_n 0.252231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_414_n 0.00532666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_D_N_M1005_g 0.0497309f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.865
cc_43 VPB D_N 0.0318572f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_44 VPB N_D_N_c_72_n 0.071146f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.73
cc_45 VPB N_A_64_131#_c_97_n 0.0347411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_64_131#_c_102_n 0.0193198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_64_131#_c_99_n 0.0272543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_C_M1007_g 0.0154125f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_49 VPB C 0.0123202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_C_c_152_n 0.0818792f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=1.73
cc_51 VPB N_B_M1003_g 0.0182705f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.865
cc_52 VPB N_B_c_197_n 0.00450165f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_53 VPB N_A_M1000_g 0.0303882f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=0.865
cc_54 VPB A 0.00473766f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.865
cc_55 VPB N_A_c_237_n 0.0462589f $X=-0.19 $Y=1.655 $X2=0.477 $Y2=2.235
cc_56 VPB N_A_220_367#_c_270_n 0.029193f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_57 VPB N_A_220_367#_c_273_n 0.00116565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_220_367#_c_280_n 0.00448485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_348_n 0.0135216f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_60 VPB N_VPWR_c_349_n 0.00474522f $X=-0.19 $Y=1.655 $X2=0.477 $Y2=1.73
cc_61 VPB N_VPWR_c_350_n 0.0227191f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=1.665
cc_62 VPB N_VPWR_c_351_n 0.00564791f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_352_n 0.0516856f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=1.73
cc_64 VPB N_VPWR_c_353_n 0.00382116f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=2.035
cc_65 VPB N_VPWR_c_354_n 0.0186439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_347_n 0.0990708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB X 0.00890576f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_68 VPB X 0.0489747f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_X_c_391_n 0.0141306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 N_D_N_M1006_g N_A_64_131#_M1002_g 0.00973518f $X=0.66 $Y=0.865 $X2=0 $Y2=0
cc_71 N_D_N_M1006_g N_A_64_131#_c_97_n 0.0262667f $X=0.66 $Y=0.865 $X2=0 $Y2=0
cc_72 N_D_N_c_72_n N_A_64_131#_c_97_n 0.00579945f $X=0.385 $Y=1.73 $X2=0 $Y2=0
cc_73 N_D_N_M1006_g N_A_64_131#_c_98_n 0.0103794f $X=0.66 $Y=0.865 $X2=0 $Y2=0
cc_74 N_D_N_M1005_g N_A_64_131#_c_102_n 0.00376522f $X=0.66 $Y=2.865 $X2=0 $Y2=0
cc_75 N_D_N_M1006_g N_A_64_131#_c_99_n 7.30551e-19 $X=0.66 $Y=0.865 $X2=0 $Y2=0
cc_76 N_D_N_M1005_g N_A_64_131#_c_99_n 0.0262926f $X=0.66 $Y=2.865 $X2=0 $Y2=0
cc_77 D_N N_A_64_131#_c_99_n 0.0664361f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_78 N_D_N_c_72_n N_A_64_131#_c_99_n 0.028728f $X=0.385 $Y=1.73 $X2=0 $Y2=0
cc_79 N_D_N_M1006_g N_A_64_131#_c_100_n 0.0261273f $X=0.66 $Y=0.865 $X2=0 $Y2=0
cc_80 D_N N_A_64_131#_c_100_n 0.0186524f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_81 N_D_N_c_72_n N_A_64_131#_c_100_n 0.00651155f $X=0.385 $Y=1.73 $X2=0 $Y2=0
cc_82 N_D_N_c_72_n N_A_220_367#_c_273_n 2.50228e-19 $X=0.385 $Y=1.73 $X2=0 $Y2=0
cc_83 N_D_N_c_72_n N_A_220_367#_c_280_n 0.00104278f $X=0.385 $Y=1.73 $X2=0 $Y2=0
cc_84 N_D_N_M1005_g N_VPWR_c_348_n 0.00487711f $X=0.66 $Y=2.865 $X2=0 $Y2=0
cc_85 N_D_N_M1005_g N_VPWR_c_350_n 0.00424641f $X=0.66 $Y=2.865 $X2=0 $Y2=0
cc_86 N_D_N_M1005_g N_VPWR_c_347_n 0.00804212f $X=0.66 $Y=2.865 $X2=0 $Y2=0
cc_87 N_D_N_M1006_g N_VGND_c_404_n 0.00344874f $X=0.66 $Y=0.865 $X2=0 $Y2=0
cc_88 N_D_N_M1006_g N_VGND_c_407_n 0.00385987f $X=0.66 $Y=0.865 $X2=0 $Y2=0
cc_89 N_D_N_M1006_g N_VGND_c_413_n 0.0046122f $X=0.66 $Y=0.865 $X2=0 $Y2=0
cc_90 N_A_64_131#_M1002_g N_C_c_145_n 0.0123309f $X=1.13 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A_64_131#_c_97_n N_C_c_147_n 0.0091082f $X=1.44 $Y=1.725 $X2=0 $Y2=0
cc_92 N_A_64_131#_c_97_n N_C_M1007_g 0.0333112f $X=1.44 $Y=1.725 $X2=0 $Y2=0
cc_93 N_A_64_131#_c_97_n C 0.00684869f $X=1.44 $Y=1.725 $X2=0 $Y2=0
cc_94 N_A_64_131#_M1002_g N_A_220_367#_c_272_n 0.0037672f $X=1.13 $Y=0.865 $X2=0
+ $Y2=0
cc_95 N_A_64_131#_c_100_n N_A_220_367#_c_272_n 0.00195992f $X=0.77 $Y=1.38 $X2=0
+ $Y2=0
cc_96 N_A_64_131#_c_97_n N_A_220_367#_c_273_n 0.0156412f $X=1.44 $Y=1.725 $X2=0
+ $Y2=0
cc_97 N_A_64_131#_c_99_n N_A_220_367#_c_273_n 0.011672f $X=0.77 $Y=2.405 $X2=0
+ $Y2=0
cc_98 N_A_64_131#_c_100_n N_A_220_367#_c_273_n 0.0106057f $X=0.77 $Y=1.38 $X2=0
+ $Y2=0
cc_99 N_A_64_131#_c_97_n N_A_220_367#_c_280_n 0.0210515f $X=1.44 $Y=1.725 $X2=0
+ $Y2=0
cc_100 N_A_64_131#_c_99_n N_A_220_367#_c_280_n 0.0276097f $X=0.77 $Y=2.405 $X2=0
+ $Y2=0
cc_101 N_A_64_131#_c_100_n N_A_220_367#_c_280_n 0.00631233f $X=0.77 $Y=1.38
+ $X2=0 $Y2=0
cc_102 N_A_64_131#_M1002_g N_A_220_367#_c_291_n 0.0044676f $X=1.13 $Y=0.865
+ $X2=0 $Y2=0
cc_103 N_A_64_131#_c_97_n N_A_220_367#_c_291_n 0.00433885f $X=1.44 $Y=1.725
+ $X2=0 $Y2=0
cc_104 N_A_64_131#_c_100_n N_A_220_367#_c_291_n 0.00105697f $X=0.77 $Y=1.38
+ $X2=0 $Y2=0
cc_105 N_A_64_131#_c_97_n N_A_220_367#_c_276_n 0.00158073f $X=1.44 $Y=1.725
+ $X2=0 $Y2=0
cc_106 N_A_64_131#_c_100_n N_A_220_367#_c_276_n 0.0151196f $X=0.77 $Y=1.38 $X2=0
+ $Y2=0
cc_107 N_A_64_131#_c_99_n N_VPWR_c_348_n 0.009432f $X=0.77 $Y=2.405 $X2=0 $Y2=0
cc_108 N_A_64_131#_c_102_n N_VPWR_c_350_n 0.0144155f $X=0.445 $Y=2.865 $X2=0
+ $Y2=0
cc_109 N_A_64_131#_c_99_n N_VPWR_c_350_n 0.00218971f $X=0.77 $Y=2.405 $X2=0
+ $Y2=0
cc_110 N_A_64_131#_c_102_n N_VPWR_c_347_n 0.0110041f $X=0.445 $Y=2.865 $X2=0
+ $Y2=0
cc_111 N_A_64_131#_c_99_n N_VPWR_c_347_n 0.00429416f $X=0.77 $Y=2.405 $X2=0
+ $Y2=0
cc_112 N_A_64_131#_M1002_g N_VGND_c_404_n 0.00344874f $X=1.13 $Y=0.865 $X2=0
+ $Y2=0
cc_113 N_A_64_131#_c_97_n N_VGND_c_404_n 4.6602e-19 $X=1.44 $Y=1.725 $X2=0 $Y2=0
cc_114 N_A_64_131#_c_100_n N_VGND_c_404_n 0.0179643f $X=0.77 $Y=1.38 $X2=0 $Y2=0
cc_115 N_A_64_131#_c_98_n N_VGND_c_407_n 0.00503613f $X=0.445 $Y=0.865 $X2=0
+ $Y2=0
cc_116 N_A_64_131#_M1002_g N_VGND_c_409_n 0.00385418f $X=1.13 $Y=0.865 $X2=0
+ $Y2=0
cc_117 N_A_64_131#_M1002_g N_VGND_c_413_n 0.0046122f $X=1.13 $Y=0.865 $X2=0
+ $Y2=0
cc_118 N_A_64_131#_c_98_n N_VGND_c_413_n 0.0094461f $X=0.445 $Y=0.865 $X2=0
+ $Y2=0
cc_119 N_C_c_145_n N_B_M1011_g 0.00659796f $X=1.56 $Y=1.185 $X2=0 $Y2=0
cc_120 N_C_c_146_n N_B_M1011_g 0.0167384f $X=1.835 $Y=1.26 $X2=0 $Y2=0
cc_121 N_C_M1007_g N_B_M1003_g 0.0305896f $X=1.91 $Y=2.045 $X2=0 $Y2=0
cc_122 C N_B_M1003_g 0.0175875f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_123 N_C_M1007_g N_B_c_197_n 0.0167384f $X=1.91 $Y=2.045 $X2=0 $Y2=0
cc_124 C N_B_c_197_n 0.00775303f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_125 N_C_c_145_n N_B_c_199_n 4.17479e-19 $X=1.56 $Y=1.185 $X2=0 $Y2=0
cc_126 N_C_M1007_g N_A_M1000_g 3.48548e-19 $X=1.91 $Y=2.045 $X2=0 $Y2=0
cc_127 C N_A_M1000_g 0.0024253f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_128 N_C_c_152_n N_A_M1000_g 0.003155f $X=1.89 $Y=2.58 $X2=0 $Y2=0
cc_129 N_C_M1007_g A 2.5745e-19 $X=1.91 $Y=2.045 $X2=0 $Y2=0
cc_130 C A 0.0901796f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_131 N_C_c_152_n A 7.4294e-19 $X=1.89 $Y=2.58 $X2=0 $Y2=0
cc_132 C N_A_c_237_n 0.00302284f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_133 N_C_c_152_n N_A_c_237_n 0.0108392f $X=1.89 $Y=2.58 $X2=0 $Y2=0
cc_134 N_C_c_145_n N_A_220_367#_c_272_n 0.00464206f $X=1.56 $Y=1.185 $X2=0 $Y2=0
cc_135 N_C_c_147_n N_A_220_367#_c_272_n 0.00164626f $X=1.635 $Y=1.26 $X2=0 $Y2=0
cc_136 N_C_M1007_g N_A_220_367#_c_273_n 0.00411196f $X=1.91 $Y=2.045 $X2=0 $Y2=0
cc_137 C N_A_220_367#_c_273_n 0.0222455f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_138 N_C_c_146_n N_A_220_367#_c_274_n 0.0141367f $X=1.835 $Y=1.26 $X2=0 $Y2=0
cc_139 N_C_c_147_n N_A_220_367#_c_274_n 0.00611461f $X=1.635 $Y=1.26 $X2=0 $Y2=0
cc_140 N_C_M1007_g N_A_220_367#_c_274_n 0.00500946f $X=1.91 $Y=2.045 $X2=0 $Y2=0
cc_141 C N_A_220_367#_c_274_n 0.046671f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_142 N_C_c_145_n N_A_220_367#_c_304_n 6.4293e-19 $X=1.56 $Y=1.185 $X2=0 $Y2=0
cc_143 N_C_c_146_n N_A_220_367#_c_304_n 3.05389e-19 $X=1.835 $Y=1.26 $X2=0 $Y2=0
cc_144 C N_A_220_367#_c_275_n 0.00132427f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_145 N_C_c_145_n N_A_220_367#_c_291_n 0.00509922f $X=1.56 $Y=1.185 $X2=0 $Y2=0
cc_146 N_C_c_147_n N_A_220_367#_c_276_n 0.00244238f $X=1.635 $Y=1.26 $X2=0 $Y2=0
cc_147 N_C_c_152_n N_VPWR_c_348_n 0.00798875f $X=1.89 $Y=2.58 $X2=0 $Y2=0
cc_148 C N_VPWR_c_349_n 0.00513087f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_149 C N_VPWR_c_352_n 0.0402787f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_C_c_152_n N_VPWR_c_352_n 0.00604818f $X=1.89 $Y=2.58 $X2=0 $Y2=0
cc_151 C N_VPWR_c_347_n 0.0209659f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_152 N_C_c_152_n N_VPWR_c_347_n 0.0118983f $X=1.89 $Y=2.58 $X2=0 $Y2=0
cc_153 C A_303_367# 0.00399078f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_154 N_C_c_145_n N_VGND_c_405_n 0.00549449f $X=1.56 $Y=1.185 $X2=0 $Y2=0
cc_155 N_C_c_146_n N_VGND_c_405_n 0.0046525f $X=1.835 $Y=1.26 $X2=0 $Y2=0
cc_156 N_C_c_145_n N_VGND_c_409_n 0.00370979f $X=1.56 $Y=1.185 $X2=0 $Y2=0
cc_157 N_C_c_145_n N_VGND_c_413_n 0.0046122f $X=1.56 $Y=1.185 $X2=0 $Y2=0
cc_158 N_B_M1011_g N_A_M1000_g 0.0306263f $X=2.27 $Y=0.865 $X2=0 $Y2=0
cc_159 N_B_c_197_n N_A_M1000_g 0.049237f $X=2.305 $Y=1.705 $X2=0 $Y2=0
cc_160 B N_A_M1000_g 0.00777305f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_161 N_B_c_199_n N_A_M1000_g 0.00121998f $X=2.24 $Y=0.38 $X2=0 $Y2=0
cc_162 N_B_M1003_g A 0.00334391f $X=2.34 $Y=2.045 $X2=0 $Y2=0
cc_163 N_B_M1003_g N_A_c_237_n 0.00139852f $X=2.34 $Y=2.045 $X2=0 $Y2=0
cc_164 N_B_M1011_g N_A_220_367#_c_272_n 8.37321e-19 $X=2.27 $Y=0.865 $X2=0 $Y2=0
cc_165 N_B_M1011_g N_A_220_367#_c_274_n 0.00895723f $X=2.27 $Y=0.865 $X2=0 $Y2=0
cc_166 B N_A_220_367#_c_274_n 0.0072898f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_167 N_B_c_199_n N_A_220_367#_c_274_n 5.18627e-19 $X=2.24 $Y=0.38 $X2=0 $Y2=0
cc_168 N_B_M1011_g N_A_220_367#_c_304_n 0.0099921f $X=2.27 $Y=0.865 $X2=0 $Y2=0
cc_169 B N_A_220_367#_c_304_n 0.0223985f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_170 N_B_c_199_n N_A_220_367#_c_304_n 2.21056e-19 $X=2.24 $Y=0.38 $X2=0 $Y2=0
cc_171 B N_A_220_367#_c_275_n 0.00193308f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_172 N_B_M1011_g N_A_220_367#_c_277_n 0.00358489f $X=2.27 $Y=0.865 $X2=0 $Y2=0
cc_173 N_B_c_197_n N_A_220_367#_c_277_n 0.00339944f $X=2.305 $Y=1.705 $X2=0
+ $Y2=0
cc_174 N_B_M1011_g N_VGND_c_405_n 0.00567419f $X=2.27 $Y=0.865 $X2=0 $Y2=0
cc_175 B N_VGND_c_405_n 0.0293367f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_176 N_B_c_199_n N_VGND_c_405_n 0.0045193f $X=2.24 $Y=0.38 $X2=0 $Y2=0
cc_177 B N_VGND_c_406_n 0.03104f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_178 N_B_c_199_n N_VGND_c_406_n 0.00284648f $X=2.24 $Y=0.38 $X2=0 $Y2=0
cc_179 B N_VGND_c_411_n 0.0342932f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_180 N_B_c_199_n N_VGND_c_411_n 0.00625935f $X=2.24 $Y=0.38 $X2=0 $Y2=0
cc_181 B N_VGND_c_413_n 0.0227615f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_182 N_B_c_199_n N_VGND_c_413_n 0.00876757f $X=2.24 $Y=0.38 $X2=0 $Y2=0
cc_183 N_A_M1000_g N_A_220_367#_c_270_n 0.0446874f $X=2.7 $Y=0.865 $X2=0 $Y2=0
cc_184 A N_A_220_367#_c_270_n 4.15161e-19 $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_185 N_A_M1000_g N_A_220_367#_M1008_g 0.0171592f $X=2.7 $Y=0.865 $X2=0 $Y2=0
cc_186 N_A_M1000_g N_A_220_367#_c_304_n 0.00869913f $X=2.7 $Y=0.865 $X2=0 $Y2=0
cc_187 N_A_M1000_g N_A_220_367#_c_275_n 0.015757f $X=2.7 $Y=0.865 $X2=0 $Y2=0
cc_188 A N_A_220_367#_c_275_n 0.00293993f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_189 N_A_M1000_g N_A_220_367#_c_277_n 0.00296801f $X=2.7 $Y=0.865 $X2=0 $Y2=0
cc_190 A N_A_220_367#_c_277_n 0.00652936f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_191 N_A_M1000_g N_VPWR_c_349_n 0.00884515f $X=2.7 $Y=0.865 $X2=0 $Y2=0
cc_192 A N_VPWR_c_349_n 0.0827025f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_193 A N_VPWR_c_352_n 0.00971876f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_194 N_A_c_237_n N_VPWR_c_352_n 0.00507663f $X=2.7 $Y=2.79 $X2=0 $Y2=0
cc_195 A N_VPWR_c_347_n 0.00916124f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_196 N_A_c_237_n N_VPWR_c_347_n 0.0037897f $X=2.7 $Y=2.79 $X2=0 $Y2=0
cc_197 A A_483_367# 0.00496341f $X=2.555 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_198 N_A_M1000_g N_VGND_c_406_n 0.00794577f $X=2.7 $Y=0.865 $X2=0 $Y2=0
cc_199 N_A_M1000_g N_VGND_c_411_n 0.00168672f $X=2.7 $Y=0.865 $X2=0 $Y2=0
cc_200 N_A_M1000_g N_VGND_c_413_n 0.0015374f $X=2.7 $Y=0.865 $X2=0 $Y2=0
cc_201 N_A_220_367#_c_270_n N_VPWR_c_349_n 0.0225231f $X=3.225 $Y=1.76 $X2=0
+ $Y2=0
cc_202 N_A_220_367#_c_275_n N_VPWR_c_349_n 0.0185189f $X=2.96 $Y=1.325 $X2=0
+ $Y2=0
cc_203 N_A_220_367#_c_270_n N_VPWR_c_354_n 0.00525069f $X=3.225 $Y=1.76 $X2=0
+ $Y2=0
cc_204 N_A_220_367#_c_270_n N_VPWR_c_347_n 0.00990586f $X=3.225 $Y=1.76 $X2=0
+ $Y2=0
cc_205 N_A_220_367#_c_270_n X 0.0158422f $X=3.225 $Y=1.76 $X2=0 $Y2=0
cc_206 N_A_220_367#_M1008_g X 0.00659419f $X=3.285 $Y=0.655 $X2=0 $Y2=0
cc_207 N_A_220_367#_c_275_n X 0.0301108f $X=2.96 $Y=1.325 $X2=0 $Y2=0
cc_208 N_A_220_367#_M1008_g X 0.00315726f $X=3.285 $Y=0.655 $X2=0 $Y2=0
cc_209 N_A_220_367#_c_270_n N_X_c_391_n 0.00623546f $X=3.225 $Y=1.76 $X2=0 $Y2=0
cc_210 N_A_220_367#_c_274_n N_VGND_c_405_n 0.0132523f $X=2.32 $Y=1.325 $X2=0
+ $Y2=0
cc_211 N_A_220_367#_c_304_n N_VGND_c_405_n 0.00769385f $X=2.485 $Y=0.93 $X2=0
+ $Y2=0
cc_212 N_A_220_367#_c_291_n N_VGND_c_405_n 0.0247741f $X=1.45 $Y=0.865 $X2=0
+ $Y2=0
cc_213 N_A_220_367#_c_270_n N_VGND_c_406_n 0.00137872f $X=3.225 $Y=1.76 $X2=0
+ $Y2=0
cc_214 N_A_220_367#_M1008_g N_VGND_c_406_n 0.0223834f $X=3.285 $Y=0.655 $X2=0
+ $Y2=0
cc_215 N_A_220_367#_c_304_n N_VGND_c_406_n 0.0144016f $X=2.485 $Y=0.93 $X2=0
+ $Y2=0
cc_216 N_A_220_367#_c_275_n N_VGND_c_406_n 0.026604f $X=2.96 $Y=1.325 $X2=0
+ $Y2=0
cc_217 N_A_220_367#_c_291_n N_VGND_c_409_n 0.00467815f $X=1.45 $Y=0.865 $X2=0
+ $Y2=0
cc_218 N_A_220_367#_M1008_g N_VGND_c_412_n 0.00486043f $X=3.285 $Y=0.655 $X2=0
+ $Y2=0
cc_219 N_A_220_367#_M1008_g N_VGND_c_413_n 0.00924722f $X=3.285 $Y=0.655 $X2=0
+ $Y2=0
cc_220 N_A_220_367#_c_291_n N_VGND_c_413_n 0.00980632f $X=1.45 $Y=0.865 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_347_n N_X_M1001_d 0.00336915f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_354_n X 0.0289189f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_c_347_n X 0.0162509f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_224 N_VPWR_c_349_n N_X_c_391_n 0.0464021f $X=3.01 $Y=1.98 $X2=0 $Y2=0
cc_225 N_X_c_387_n N_VGND_c_412_n 0.0242629f $X=3.5 $Y=0.42 $X2=0 $Y2=0
cc_226 N_X_M1008_d N_VGND_c_413_n 0.00371702f $X=3.36 $Y=0.235 $X2=0 $Y2=0
cc_227 N_X_c_387_n N_VGND_c_413_n 0.0135294f $X=3.5 $Y=0.42 $X2=0 $Y2=0
