* File: sky130_fd_sc_lp__o21a_2.pex.spice
* Created: Wed Sep  2 10:15:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21A_2%A_86_21# 1 2 7 9 12 16 18 21 23 25 26 28 29
+ 32 34 36 38 42 47
c73 21 0 1.03991e-20 $X=0.935 $Y=2.465
r74 46 47 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.935 $Y=1.35
+ $X2=0.86 $Y2=1.35
r75 42 46 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.15 $Y=1.35
+ $X2=0.935 $Y2=1.35
r76 41 43 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.15 $Y=1.35
+ $X2=1.15 $Y2=1.52
r77 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.35 $X2=1.15 $Y2=1.35
r78 38 41 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.15 $Y2=1.35
r79 34 45 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=2.09
+ $X2=2.135 $Y2=2.005
r80 34 36 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=2.135 $Y=2.09
+ $X2=2.135 $Y2=2.45
r81 30 32 25.5881 $w=2.93e-07 $l=6.55e-07 $layer=LI1_cond $X=1.652 $Y=1.075
+ $X2=1.652 $Y2=0.42
r82 28 45 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.005 $Y=2.005
+ $X2=2.135 $Y2=2.005
r83 28 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.005 $Y=2.005
+ $X2=1.315 $Y2=2.005
r84 27 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=1.16
+ $X2=1.15 $Y2=1.16
r85 26 30 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=1.505 $Y=1.16
+ $X2=1.652 $Y2=1.075
r86 26 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.505 $Y=1.16
+ $X2=1.315 $Y2=1.16
r87 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=1.92
+ $X2=1.315 $Y2=2.005
r88 25 43 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.23 $Y=1.92 $X2=1.23
+ $Y2=1.52
r89 19 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.515
+ $X2=0.935 $Y2=1.35
r90 19 21 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.935 $Y=1.515
+ $X2=0.935 $Y2=2.465
r91 16 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.185
+ $X2=0.935 $Y2=1.35
r92 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.935 $Y=1.185
+ $X2=0.935 $Y2=0.655
r93 15 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.58 $Y=1.26
+ $X2=0.505 $Y2=1.26
r94 15 47 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.58 $Y=1.26
+ $X2=0.86 $Y2=1.26
r95 10 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.505 $Y=1.335
+ $X2=0.505 $Y2=1.26
r96 10 12 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=0.505 $Y=1.335
+ $X2=0.505 $Y2=2.465
r97 7 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.505 $Y=1.185
+ $X2=0.505 $Y2=1.26
r98 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.505 $Y=1.185
+ $X2=0.505 $Y2=0.655
r99 2 45 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.835 $X2=2.1 $Y2=2.005
r100 2 36 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=1.835 $X2=2.1 $Y2=2.45
r101 1 32 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.545
+ $Y=0.255 $X2=1.67 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_2%B1 3 7 9 12 13
c34 13 0 7.37516e-20 $X=1.73 $Y=1.51
r35 12 15 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.762 $Y=1.51
+ $X2=1.762 $Y2=1.675
r36 12 14 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.762 $Y=1.51
+ $X2=1.762 $Y2=1.345
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.51 $X2=1.73 $Y2=1.51
r38 9 13 4.3568 $w=4.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.69 $Y=1.665
+ $X2=1.69 $Y2=1.51
r39 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.885 $Y=2.465
+ $X2=1.885 $Y2=1.675
r40 3 14 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.885 $Y=0.675
+ $X2=1.885 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_2%A2 3 7 9 10 14
c34 14 0 1.54831e-19 $X=2.335 $Y=1.51
c35 7 0 6.33525e-20 $X=2.315 $Y=2.465
r36 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.51
+ $X2=2.335 $Y2=1.675
r37 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.51
+ $X2=2.335 $Y2=1.345
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.335
+ $Y=1.51 $X2=2.335 $Y2=1.51
r39 10 15 9.3732 $w=3.73e-07 $l=3.05e-07 $layer=LI1_cond $X=2.64 $Y=1.562
+ $X2=2.335 $Y2=1.562
r40 9 15 5.37807 $w=3.73e-07 $l=1.75e-07 $layer=LI1_cond $X=2.16 $Y=1.562
+ $X2=2.335 $Y2=1.562
r41 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.315 $Y=2.465
+ $X2=2.315 $Y2=1.675
r42 3 16 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.315 $Y=0.675
+ $X2=2.315 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_2%A1 3 7 9 14 15
c25 15 0 1.54831e-19 $X=3.07 $Y=1.46
r26 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.46 $X2=3.07 $Y2=1.46
r27 11 14 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.785 $Y=1.46
+ $X2=3.07 $Y2=1.46
r28 9 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.46
r29 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.625
+ $X2=2.785 $Y2=1.46
r30 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.785 $Y=1.625
+ $X2=2.785 $Y2=2.465
r31 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.295
+ $X2=2.785 $Y2=1.46
r32 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.785 $Y=1.295
+ $X2=2.785 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_2%VPWR 1 2 3 10 12 18 20 22 26 28 33 42 46
r44 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 37 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 34 42 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.41 $Y2=3.33
r49 34 36 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 33 45 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.097 $Y2=3.33
r51 33 36 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 32 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 29 39 4.1687 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.197 $Y2=3.33
r55 29 31 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 28 42 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.41 $Y2=3.33
r57 28 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 26 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 26 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 26 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 22 25 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=3 $Y=2.005 $X2=3
+ $Y2=2.95
r62 20 45 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=3 $Y=3.245
+ $X2=3.097 $Y2=3.33
r63 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.95
r64 16 42 3.24638 $w=8.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=3.245
+ $X2=1.41 $Y2=3.33
r65 16 18 12.2718 $w=8.48e-07 $l=8.55e-07 $layer=LI1_cond $X=1.41 $Y=3.245
+ $X2=1.41 $Y2=2.39
r66 12 15 41.4026 $w=2.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.26 $Y=1.98
+ $X2=0.26 $Y2=2.95
r67 10 39 3.116 $w=2.7e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.197 $Y2=3.33
r68 10 15 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r69 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.835 $X2=3 $Y2=2.95
r70 3 22 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.835 $X2=3 $Y2=2.005
r71 2 18 150 $w=1.7e-07 $l=8.95489e-07 $layer=licon1_PDIFF $count=4 $X=1.01
+ $Y=1.835 $X2=1.67 $Y2=2.39
r72 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.95
r73 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_2%X 1 2 7 8 9 10 11 12 13 22
r18 13 40 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.69 $Y=2.775
+ $X2=0.69 $Y2=2.91
r19 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=2.405
+ $X2=0.69 $Y2=2.775
r20 11 12 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=0.69 $Y=1.98
+ $X2=0.69 $Y2=2.405
r21 10 11 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=1.665
+ $X2=0.69 $Y2=1.98
r22 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=1.295
+ $X2=0.69 $Y2=1.665
r23 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=0.925 $X2=0.69
+ $Y2=1.295
r24 7 8 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=0.555 $X2=0.69
+ $Y2=0.925
r25 7 22 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.69 $Y=0.555
+ $X2=0.69 $Y2=0.42
r26 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.91
r27 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=1.98
r28 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.58
+ $Y=0.235 $X2=0.72 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_2%VGND 1 2 3 10 12 16 20 23 24 25 27 37 38 44
r43 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r45 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r47 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=1.15
+ $Y2=0
r49 32 34 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=2.16
+ $Y2=0
r50 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r51 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r52 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 28 41 4.1687 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r54 28 30 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.72
+ $Y2=0
r55 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.15
+ $Y2=0
r56 27 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r57 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r58 25 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 23 34 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.16
+ $Y2=0
r60 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.55
+ $Y2=0
r61 22 37 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=3.12
+ $Y2=0
r62 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.55
+ $Y2=0
r63 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=0.085
+ $X2=2.55 $Y2=0
r64 18 20 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.55 $Y=0.085
+ $X2=2.55 $Y2=0.4
r65 14 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0
r66 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.38
r67 10 41 3.116 $w=2.7e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.197 $Y2=0
r68 10 12 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r69 3 20 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=2.39
+ $Y=0.255 $X2=2.55 $Y2=0.4
r70 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.01
+ $Y=0.235 $X2=1.15 $Y2=0.38
r71 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_2%A_392_51# 1 2 9 11 12 15
r20 13 15 25.3126 $w=2.78e-07 $l=6.15e-07 $layer=LI1_cond $X=3.025 $Y=1.035
+ $X2=3.025 $Y2=0.42
r21 11 13 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.885 $Y=1.12
+ $X2=3.025 $Y2=1.035
r22 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.885 $Y=1.12
+ $X2=2.215 $Y2=1.12
r23 7 12 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=2.092 $Y=1.035
+ $X2=2.215 $Y2=1.12
r24 7 9 28.9287 $w=2.43e-07 $l=6.15e-07 $layer=LI1_cond $X=2.092 $Y=1.035
+ $X2=2.092 $Y2=0.42
r25 2 15 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.86
+ $Y=0.255 $X2=3 $Y2=0.42
r26 1 9 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.96
+ $Y=0.255 $X2=2.1 $Y2=0.42
.ends

