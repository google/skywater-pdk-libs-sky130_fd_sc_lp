# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__or3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__or3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.910000 1.425000 2.305000 2.120000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 1.125000 2.815000 2.120000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.405000 0.580000 1.750000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.100000 0.255000 1.360000 1.010000 ;
        RECT 1.100000 1.010000 1.270000 1.815000 ;
        RECT 1.100000 1.815000 1.575000 2.120000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.125000  0.700000 0.385000 1.065000 ;
      RECT 0.125000  1.065000 0.930000 1.235000 ;
      RECT 0.290000  1.920000 0.930000 2.290000 ;
      RECT 0.290000  2.290000 2.815000 2.460000 ;
      RECT 0.555000  0.085000 0.930000 0.895000 ;
      RECT 0.750000  1.235000 0.930000 1.920000 ;
      RECT 0.815000  2.640000 1.145000 3.245000 ;
      RECT 1.440000  1.190000 2.305000 1.235000 ;
      RECT 1.440000  1.235000 1.720000 1.520000 ;
      RECT 1.530000  0.085000 1.930000 0.895000 ;
      RECT 1.550000  1.065000 2.305000 1.190000 ;
      RECT 1.675000  2.640000 2.005000 3.245000 ;
      RECT 2.100000  0.280000 2.315000 0.785000 ;
      RECT 2.100000  0.785000 3.265000 0.955000 ;
      RECT 2.100000  0.955000 2.305000 1.065000 ;
      RECT 2.485000  0.085000 2.815000 0.615000 ;
      RECT 2.485000  2.460000 2.815000 2.965000 ;
      RECT 2.985000  0.280000 3.265000 0.785000 ;
      RECT 2.985000  0.955000 3.265000 2.300000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__or3b_2
END LIBRARY
