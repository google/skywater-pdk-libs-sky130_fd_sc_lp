* File: sky130_fd_sc_lp__a311o_lp.pxi.spice
* Created: Wed Sep  2 09:25:20 2020
* 
x_PM_SKY130_FD_SC_LP__A311O_LP%A_85_21# N_A_85_21#_M1002_d N_A_85_21#_M1013_d
+ N_A_85_21#_M1009_d N_A_85_21#_M1014_g N_A_85_21#_c_107_n N_A_85_21#_M1006_g
+ N_A_85_21#_M1007_g N_A_85_21#_c_96_n N_A_85_21#_c_97_n N_A_85_21#_c_98_n
+ N_A_85_21#_c_99_n N_A_85_21#_c_133_p N_A_85_21#_c_100_n N_A_85_21#_c_110_n
+ N_A_85_21#_c_101_n N_A_85_21#_c_102_n N_A_85_21#_c_103_n N_A_85_21#_c_104_n
+ N_A_85_21#_c_111_n N_A_85_21#_c_105_n N_A_85_21#_c_106_n
+ PM_SKY130_FD_SC_LP__A311O_LP%A_85_21#
x_PM_SKY130_FD_SC_LP__A311O_LP%A3 N_A3_c_215_n N_A3_M1003_g N_A3_c_209_n
+ N_A3_M1004_g N_A3_c_210_n N_A3_c_211_n N_A3_c_212_n A3 N_A3_c_213_n
+ N_A3_c_214_n PM_SKY130_FD_SC_LP__A311O_LP%A3
x_PM_SKY130_FD_SC_LP__A311O_LP%A2 N_A2_M1008_g N_A2_M1001_g N_A2_c_263_n
+ N_A2_c_268_n A2 N_A2_c_264_n N_A2_c_265_n PM_SKY130_FD_SC_LP__A311O_LP%A2
x_PM_SKY130_FD_SC_LP__A311O_LP%A1 N_A1_M1002_g N_A1_c_307_n N_A1_M1000_g
+ N_A1_c_308_n N_A1_c_309_n N_A1_c_315_n A1 A1 N_A1_c_311_n N_A1_c_312_n
+ PM_SKY130_FD_SC_LP__A311O_LP%A1
x_PM_SKY130_FD_SC_LP__A311O_LP%B1 N_B1_c_361_n N_B1_M1010_g N_B1_M1011_g
+ N_B1_c_362_n N_B1_M1005_g N_B1_c_363_n B1 B1 B1 B1 N_B1_c_364_n N_B1_c_365_n
+ N_B1_c_366_n PM_SKY130_FD_SC_LP__A311O_LP%B1
x_PM_SKY130_FD_SC_LP__A311O_LP%C1 N_C1_c_419_n N_C1_M1012_g N_C1_M1009_g
+ N_C1_c_420_n N_C1_M1013_g N_C1_c_421_n N_C1_c_422_n N_C1_c_423_n N_C1_c_428_n
+ C1 N_C1_c_424_n N_C1_c_425_n PM_SKY130_FD_SC_LP__A311O_LP%C1
x_PM_SKY130_FD_SC_LP__A311O_LP%X N_X_M1014_s N_X_M1006_s N_X_c_467_n N_X_c_470_n
+ N_X_c_471_n N_X_c_468_n X X PM_SKY130_FD_SC_LP__A311O_LP%X
x_PM_SKY130_FD_SC_LP__A311O_LP%VPWR N_VPWR_M1006_d N_VPWR_M1008_d N_VPWR_c_497_n
+ N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n
+ VPWR N_VPWR_c_503_n N_VPWR_c_496_n PM_SKY130_FD_SC_LP__A311O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A311O_LP%A_257_414# N_A_257_414#_M1003_d
+ N_A_257_414#_M1000_d N_A_257_414#_c_544_n N_A_257_414#_c_550_n
+ N_A_257_414#_c_545_n N_A_257_414#_c_546_n N_A_257_414#_c_558_n
+ PM_SKY130_FD_SC_LP__A311O_LP%A_257_414#
x_PM_SKY130_FD_SC_LP__A311O_LP%VGND N_VGND_M1007_d N_VGND_M1005_d N_VGND_c_583_n
+ N_VGND_c_584_n VGND N_VGND_c_585_n N_VGND_c_586_n N_VGND_c_587_n
+ N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n PM_SKY130_FD_SC_LP__A311O_LP%VGND
cc_1 VNB N_A_85_21#_M1014_g 0.0209274f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_2 VNB N_A_85_21#_M1007_g 0.0184814f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.445
cc_3 VNB N_A_85_21#_c_96_n 0.0189012f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.96
cc_4 VNB N_A_85_21#_c_97_n 0.0186396f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.52
cc_5 VNB N_A_85_21#_c_98_n 0.00807508f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.76
cc_6 VNB N_A_85_21#_c_99_n 0.0345744f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.935
cc_7 VNB N_A_85_21#_c_100_n 0.0155823f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=0.935
cc_8 VNB N_A_85_21#_c_101_n 0.0230694f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=0.47
cc_9 VNB N_A_85_21#_c_102_n 0.00233856f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.015
cc_10 VNB N_A_85_21#_c_103_n 0.0311545f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.015
cc_11 VNB N_A_85_21#_c_104_n 0.00222923f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.935
cc_12 VNB N_A_85_21#_c_105_n 0.0302905f $X=-0.19 $Y=-0.245 $X2=3.957 $Y2=2.05
cc_13 VNB N_A_85_21#_c_106_n 0.0166071f $X=-0.19 $Y=-0.245 $X2=3.995 $Y2=0.935
cc_14 VNB N_A3_c_209_n 0.0148488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_c_210_n 0.0175882f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_16 VNB N_A3_c_211_n 0.0204286f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_17 VNB N_A3_c_212_n 0.0174729f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.76
cc_18 VNB N_A3_c_213_n 0.0163656f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.81
cc_19 VNB N_A3_c_214_n 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.445
cc_20 VNB N_A2_M1001_g 0.0378953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_c_263_n 0.0200641f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_22 VNB N_A2_c_264_n 0.0164034f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.885
cc_23 VNB N_A2_c_265_n 0.00166572f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.57
cc_24 VNB N_A1_c_307_n 0.0173545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_c_308_n 0.0140052f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.445
cc_26 VNB N_A1_c_309_n 0.00718099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A1 0.00553354f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.885
cc_28 VNB N_A1_c_311_n 0.0156903f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.81
cc_29 VNB N_A1_c_312_n 0.0172406f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.445
cc_30 VNB N_B1_c_361_n 0.0135257f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.235
cc_31 VNB N_B1_c_362_n 0.0136222f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.81
cc_32 VNB N_B1_c_363_n 0.0222409f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.885
cc_33 VNB N_B1_c_364_n 0.0458148f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.34
cc_34 VNB N_B1_c_365_n 0.00307656f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.52
cc_35 VNB N_B1_c_366_n 0.0232525f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.76
cc_36 VNB N_C1_c_419_n 0.0136222f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.235
cc_37 VNB N_C1_c_420_n 0.0172357f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.81
cc_38 VNB N_C1_c_421_n 0.024124f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.885
cc_39 VNB N_C1_c_422_n 0.0231934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_C1_c_423_n 0.0204984f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.81
cc_41 VNB N_C1_c_424_n 0.0147484f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.81
cc_42 VNB N_C1_c_425_n 0.00473252f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.96
cc_43 VNB N_X_c_467_n 0.0173365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_X_c_468_n 0.0468363f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.76
cc_45 VNB X 0.00758559f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.57
cc_46 VNB N_VPWR_c_496_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_583_n 0.00507466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_584_n 0.0027509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_585_n 0.027718f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.57
cc_50 VNB N_VGND_c_586_n 0.0479595f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.445
cc_51 VNB N_VGND_c_587_n 0.0290969f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.935
cc_52 VNB N_VGND_c_588_n 0.230975f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.935
cc_53 VNB N_VGND_c_589_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.47
cc_54 VNB N_VGND_c_590_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=0.935
cc_55 VPB N_A_85_21#_c_107_n 0.0101691f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.885
cc_56 VPB N_A_85_21#_M1006_g 0.0310091f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.57
cc_57 VPB N_A_85_21#_c_98_n 0.00626723f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.76
cc_58 VPB N_A_85_21#_c_110_n 0.0357647f $X=-0.19 $Y=1.655 $X2=3.895 $Y2=2.9
cc_59 VPB N_A_85_21#_c_111_n 0.0179524f $X=-0.19 $Y=1.655 $X2=3.895 $Y2=2.215
cc_60 VPB N_A_85_21#_c_105_n 0.0189541f $X=-0.19 $Y=1.655 $X2=3.957 $Y2=2.05
cc_61 VPB N_A3_c_215_n 0.0139268f $X=-0.19 $Y=1.655 $X2=2.25 $Y2=0.235
cc_62 VPB N_A3_M1003_g 0.0281322f $X=-0.19 $Y=1.655 $X2=3.755 $Y2=2.07
cc_63 VPB N_A3_c_211_n 0.00360137f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_64 VPB N_A3_c_214_n 7.45264e-19 $X=-0.19 $Y=1.655 $X2=0.86 $Y2=0.445
cc_65 VPB N_A2_M1008_g 0.0293588f $X=-0.19 $Y=1.655 $X2=3.755 $Y2=2.07
cc_66 VPB N_A2_c_263_n 0.00340188f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_67 VPB N_A2_c_268_n 0.0135495f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_68 VPB N_A2_c_265_n 7.46168e-19 $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.57
cc_69 VPB N_A1_c_307_n 0.00258471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A1_M1000_g 0.0296766f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.81
cc_71 VPB N_A1_c_315_n 0.0130609f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.52
cc_72 VPB A1 0.00459983f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.885
cc_73 VPB N_B1_M1011_g 0.0271805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_B1_c_364_n 0.0308659f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.34
cc_75 VPB N_B1_c_365_n 0.00171813f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.52
cc_76 VPB N_C1_M1009_g 0.0359841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_C1_c_423_n 0.00347552f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=0.81
cc_78 VPB N_C1_c_428_n 0.0139582f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=0.445
cc_79 VPB N_C1_c_425_n 0.00298138f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.96
cc_80 VPB N_X_c_470_n 0.0350556f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_81 VPB N_X_c_471_n 0.0162763f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.52
cc_82 VPB N_X_c_468_n 0.0199387f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.76
cc_83 VPB N_VPWR_c_497_n 0.0103441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_498_n 0.00356003f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.76
cc_85 VPB N_VPWR_c_499_n 0.0205887f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.57
cc_86 VPB N_VPWR_c_500_n 0.00467382f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_501_n 0.018376f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=0.445
cc_88 VPB N_VPWR_c_502_n 0.00529797f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=0.445
cc_89 VPB N_VPWR_c_503_n 0.0627992f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=0.47
cc_90 VPB N_VPWR_c_496_n 0.0718784f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_257_414#_c_544_n 0.00906025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_257_414#_c_545_n 0.00768109f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.445
cc_93 VPB N_A_257_414#_c_546_n 0.00268116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 N_A_85_21#_c_107_n N_A3_c_215_n 0.00634947f $X=0.63 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A_85_21#_c_107_n N_A3_M1003_g 0.0166121f $X=0.63 $Y=1.885 $X2=0 $Y2=0
cc_96 N_A_85_21#_M1007_g N_A3_c_209_n 0.0119319f $X=0.86 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_85_21#_c_96_n N_A3_c_210_n 0.00681265f $X=0.68 $Y=0.96 $X2=0 $Y2=0
cc_98 N_A_85_21#_c_99_n N_A3_c_210_n 0.0077922f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_99 N_A_85_21#_c_102_n N_A3_c_210_n 0.00103519f $X=0.62 $Y=1.015 $X2=0 $Y2=0
cc_100 N_A_85_21#_c_103_n N_A3_c_210_n 0.00785859f $X=0.62 $Y=1.015 $X2=0 $Y2=0
cc_101 N_A_85_21#_c_97_n N_A3_c_211_n 0.0097844f $X=0.605 $Y=1.52 $X2=0 $Y2=0
cc_102 N_A_85_21#_c_98_n N_A3_c_211_n 0.00930496f $X=0.63 $Y=1.76 $X2=0 $Y2=0
cc_103 N_A_85_21#_M1007_g N_A3_c_212_n 0.00681265f $X=0.86 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_85_21#_c_99_n N_A3_c_212_n 0.00852073f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_105 N_A_85_21#_c_99_n N_A3_c_213_n 0.00123028f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_106 N_A_85_21#_c_102_n N_A3_c_213_n 0.00111105f $X=0.62 $Y=1.015 $X2=0 $Y2=0
cc_107 N_A_85_21#_c_103_n N_A3_c_213_n 0.0097844f $X=0.62 $Y=1.015 $X2=0 $Y2=0
cc_108 N_A_85_21#_c_107_n N_A3_c_214_n 7.47265e-19 $X=0.63 $Y=1.885 $X2=0 $Y2=0
cc_109 N_A_85_21#_c_98_n N_A3_c_214_n 0.00142919f $X=0.63 $Y=1.76 $X2=0 $Y2=0
cc_110 N_A_85_21#_c_99_n N_A3_c_214_n 0.0245051f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_111 N_A_85_21#_c_102_n N_A3_c_214_n 0.0202161f $X=0.62 $Y=1.015 $X2=0 $Y2=0
cc_112 N_A_85_21#_c_103_n N_A3_c_214_n 0.00112926f $X=0.62 $Y=1.015 $X2=0 $Y2=0
cc_113 N_A_85_21#_c_99_n N_A2_M1001_g 0.0122247f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_114 N_A_85_21#_c_133_p N_A2_M1001_g 0.00289391f $X=2.39 $Y=0.47 $X2=0 $Y2=0
cc_115 N_A_85_21#_c_99_n N_A2_c_264_n 0.00119584f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_116 N_A_85_21#_c_99_n N_A2_c_265_n 0.0245014f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_117 N_A_85_21#_c_133_p N_A1_c_308_n 0.00940601f $X=2.39 $Y=0.47 $X2=0 $Y2=0
cc_118 N_A_85_21#_c_99_n N_A1_c_309_n 0.00372778f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_119 N_A_85_21#_c_133_p N_A1_c_309_n 0.00365256f $X=2.39 $Y=0.47 $X2=0 $Y2=0
cc_120 N_A_85_21#_c_104_n N_A1_c_309_n 4.29605e-19 $X=2.39 $Y=0.935 $X2=0 $Y2=0
cc_121 N_A_85_21#_c_99_n A1 0.013485f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_122 N_A_85_21#_c_100_n A1 0.0158875f $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_123 N_A_85_21#_c_104_n A1 0.0283601f $X=2.39 $Y=0.935 $X2=0 $Y2=0
cc_124 N_A_85_21#_c_104_n N_A1_c_311_n 0.00528112f $X=2.39 $Y=0.935 $X2=0 $Y2=0
cc_125 N_A_85_21#_c_99_n N_A1_c_312_n 0.00465552f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_126 N_A_85_21#_c_104_n N_A1_c_312_n 0.00321152f $X=2.39 $Y=0.935 $X2=0 $Y2=0
cc_127 N_A_85_21#_c_133_p N_B1_c_361_n 0.00866012f $X=2.39 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_85_21#_c_133_p N_B1_c_362_n 0.00139826f $X=2.39 $Y=0.47 $X2=0 $Y2=0
cc_129 N_A_85_21#_c_133_p N_B1_c_363_n 0.0070021f $X=2.39 $Y=0.47 $X2=0 $Y2=0
cc_130 N_A_85_21#_c_100_n N_B1_c_363_n 0.0174595f $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_131 N_A_85_21#_c_104_n N_B1_c_363_n 8.50662e-19 $X=2.39 $Y=0.935 $X2=0 $Y2=0
cc_132 N_A_85_21#_c_100_n N_B1_c_364_n 0.00306381f $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_133 N_A_85_21#_c_100_n N_B1_c_365_n 0.0215685f $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_134 N_A_85_21#_c_111_n N_B1_c_365_n 0.0306368f $X=3.895 $Y=2.215 $X2=0 $Y2=0
cc_135 N_A_85_21#_c_100_n N_B1_c_366_n 0.0129007f $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_136 N_A_85_21#_c_101_n N_C1_c_419_n 0.00139826f $X=3.97 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_85_21#_c_110_n N_C1_M1009_g 0.020649f $X=3.895 $Y=2.9 $X2=0 $Y2=0
cc_138 N_A_85_21#_c_111_n N_C1_M1009_g 0.00536428f $X=3.895 $Y=2.215 $X2=0 $Y2=0
cc_139 N_A_85_21#_c_105_n N_C1_M1009_g 0.00427061f $X=3.957 $Y=2.05 $X2=0 $Y2=0
cc_140 N_A_85_21#_c_101_n N_C1_c_420_n 0.00936739f $X=3.97 $Y=0.47 $X2=0 $Y2=0
cc_141 N_A_85_21#_c_100_n N_C1_c_421_n 0.0174273f $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_142 N_A_85_21#_c_101_n N_C1_c_421_n 0.00801072f $X=3.97 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A_85_21#_c_106_n N_C1_c_421_n 9.00015e-19 $X=3.995 $Y=0.935 $X2=0 $Y2=0
cc_144 N_A_85_21#_c_100_n N_C1_c_422_n 0.00991684f $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_145 N_A_85_21#_c_105_n N_C1_c_422_n 0.00362326f $X=3.957 $Y=2.05 $X2=0 $Y2=0
cc_146 N_A_85_21#_c_111_n N_C1_c_428_n 6.14058e-19 $X=3.895 $Y=2.215 $X2=0 $Y2=0
cc_147 N_A_85_21#_c_100_n N_C1_c_424_n 4.88897e-19 $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_148 N_A_85_21#_c_105_n N_C1_c_424_n 0.0148853f $X=3.957 $Y=2.05 $X2=0 $Y2=0
cc_149 N_A_85_21#_c_100_n N_C1_c_425_n 0.0238642f $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_150 N_A_85_21#_c_111_n N_C1_c_425_n 0.00867382f $X=3.895 $Y=2.215 $X2=0 $Y2=0
cc_151 N_A_85_21#_c_105_n N_C1_c_425_n 0.0483772f $X=3.957 $Y=2.05 $X2=0 $Y2=0
cc_152 N_A_85_21#_c_106_n N_C1_c_425_n 0.00247288f $X=3.995 $Y=0.935 $X2=0 $Y2=0
cc_153 N_A_85_21#_M1006_g N_X_c_470_n 0.0137539f $X=0.63 $Y=2.57 $X2=0 $Y2=0
cc_154 N_A_85_21#_M1006_g N_X_c_471_n 0.00464668f $X=0.63 $Y=2.57 $X2=0 $Y2=0
cc_155 N_A_85_21#_c_97_n N_X_c_471_n 0.0013496f $X=0.605 $Y=1.52 $X2=0 $Y2=0
cc_156 N_A_85_21#_c_102_n N_X_c_471_n 0.00264316f $X=0.62 $Y=1.015 $X2=0 $Y2=0
cc_157 N_A_85_21#_M1014_g N_X_c_468_n 0.0223711f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_85_21#_c_98_n N_X_c_468_n 0.017514f $X=0.63 $Y=1.76 $X2=0 $Y2=0
cc_159 N_A_85_21#_c_102_n N_X_c_468_n 0.0488877f $X=0.62 $Y=1.015 $X2=0 $Y2=0
cc_160 N_A_85_21#_M1014_g X 0.0141751f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_85_21#_M1007_g X 0.00976617f $X=0.86 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_85_21#_c_96_n X 8.36052e-19 $X=0.68 $Y=0.96 $X2=0 $Y2=0
cc_163 N_A_85_21#_c_99_n X 0.00334559f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_164 N_A_85_21#_c_102_n X 0.0256578f $X=0.62 $Y=1.015 $X2=0 $Y2=0
cc_165 N_A_85_21#_M1006_g N_VPWR_c_497_n 0.0239485f $X=0.63 $Y=2.57 $X2=0 $Y2=0
cc_166 N_A_85_21#_c_97_n N_VPWR_c_497_n 2.0969e-19 $X=0.605 $Y=1.52 $X2=0 $Y2=0
cc_167 N_A_85_21#_c_102_n N_VPWR_c_497_n 0.00188819f $X=0.62 $Y=1.015 $X2=0
+ $Y2=0
cc_168 N_A_85_21#_M1006_g N_VPWR_c_499_n 0.00803832f $X=0.63 $Y=2.57 $X2=0 $Y2=0
cc_169 N_A_85_21#_c_110_n N_VPWR_c_503_n 0.0281861f $X=3.895 $Y=2.9 $X2=0 $Y2=0
cc_170 N_A_85_21#_M1006_g N_VPWR_c_496_n 0.0144375f $X=0.63 $Y=2.57 $X2=0 $Y2=0
cc_171 N_A_85_21#_c_110_n N_VPWR_c_496_n 0.0174072f $X=3.895 $Y=2.9 $X2=0 $Y2=0
cc_172 N_A_85_21#_M1007_g N_VGND_c_583_n 0.00707908f $X=0.86 $Y=0.445 $X2=0
+ $Y2=0
cc_173 N_A_85_21#_c_99_n N_VGND_c_583_n 0.0252198f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_174 N_A_85_21#_c_133_p N_VGND_c_584_n 0.0135502f $X=2.39 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A_85_21#_c_100_n N_VGND_c_584_n 0.025548f $X=3.805 $Y=0.935 $X2=0 $Y2=0
cc_176 N_A_85_21#_c_101_n N_VGND_c_584_n 0.0135502f $X=3.97 $Y=0.47 $X2=0 $Y2=0
cc_177 N_A_85_21#_M1014_g N_VGND_c_585_n 0.00359964f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A_85_21#_M1007_g N_VGND_c_585_n 0.00510244f $X=0.86 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_A_85_21#_c_133_p N_VGND_c_586_n 0.0178561f $X=2.39 $Y=0.47 $X2=0 $Y2=0
cc_180 N_A_85_21#_c_101_n N_VGND_c_587_n 0.0197885f $X=3.97 $Y=0.47 $X2=0 $Y2=0
cc_181 N_A_85_21#_M1002_d N_VGND_c_588_n 0.0022543f $X=2.25 $Y=0.235 $X2=0 $Y2=0
cc_182 N_A_85_21#_M1013_d N_VGND_c_588_n 0.00232985f $X=3.83 $Y=0.235 $X2=0
+ $Y2=0
cc_183 N_A_85_21#_M1014_g N_VGND_c_588_n 0.00624174f $X=0.5 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_85_21#_M1007_g N_VGND_c_588_n 0.0061947f $X=0.86 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A_85_21#_c_99_n N_VGND_c_588_n 0.0338503f $X=2.225 $Y=0.935 $X2=0 $Y2=0
cc_186 N_A_85_21#_c_133_p N_VGND_c_588_n 0.0124703f $X=2.39 $Y=0.47 $X2=0 $Y2=0
cc_187 N_A_85_21#_c_100_n N_VGND_c_588_n 0.0276035f $X=3.805 $Y=0.935 $X2=0
+ $Y2=0
cc_188 N_A_85_21#_c_101_n N_VGND_c_588_n 0.0125808f $X=3.97 $Y=0.47 $X2=0 $Y2=0
cc_189 N_A_85_21#_c_106_n N_VGND_c_588_n 0.00195436f $X=3.995 $Y=0.935 $X2=0
+ $Y2=0
cc_190 N_A3_M1003_g N_A2_M1008_g 0.0172924f $X=1.16 $Y=2.57 $X2=0 $Y2=0
cc_191 N_A3_c_209_n N_A2_M1001_g 0.0435687f $X=1.395 $Y=0.73 $X2=0 $Y2=0
cc_192 N_A3_c_210_n N_A2_M1001_g 0.0109094f $X=1.16 $Y=1.2 $X2=0 $Y2=0
cc_193 N_A3_c_211_n N_A2_c_263_n 0.0135694f $X=1.16 $Y=1.705 $X2=0 $Y2=0
cc_194 N_A3_c_215_n N_A2_c_268_n 0.0135694f $X=1.16 $Y=1.87 $X2=0 $Y2=0
cc_195 N_A3_c_213_n N_A2_c_264_n 0.0135694f $X=1.16 $Y=1.365 $X2=0 $Y2=0
cc_196 N_A3_c_214_n N_A2_c_264_n 0.00232658f $X=1.16 $Y=1.365 $X2=0 $Y2=0
cc_197 N_A3_c_213_n N_A2_c_265_n 0.00232658f $X=1.16 $Y=1.365 $X2=0 $Y2=0
cc_198 N_A3_c_214_n N_A2_c_265_n 0.0423335f $X=1.16 $Y=1.365 $X2=0 $Y2=0
cc_199 N_A3_M1003_g N_X_c_471_n 2.63752e-19 $X=1.16 $Y=2.57 $X2=0 $Y2=0
cc_200 N_A3_c_215_n N_VPWR_c_497_n 3.03142e-19 $X=1.16 $Y=1.87 $X2=0 $Y2=0
cc_201 N_A3_M1003_g N_VPWR_c_497_n 0.0225921f $X=1.16 $Y=2.57 $X2=0 $Y2=0
cc_202 N_A3_c_214_n N_VPWR_c_497_n 0.00526295f $X=1.16 $Y=1.365 $X2=0 $Y2=0
cc_203 N_A3_M1003_g N_VPWR_c_498_n 8.17405e-19 $X=1.16 $Y=2.57 $X2=0 $Y2=0
cc_204 N_A3_M1003_g N_VPWR_c_501_n 0.00803832f $X=1.16 $Y=2.57 $X2=0 $Y2=0
cc_205 N_A3_M1003_g N_VPWR_c_496_n 0.0135635f $X=1.16 $Y=2.57 $X2=0 $Y2=0
cc_206 N_A3_c_215_n N_A_257_414#_c_544_n 3.02817e-19 $X=1.16 $Y=1.87 $X2=0 $Y2=0
cc_207 N_A3_M1003_g N_A_257_414#_c_544_n 0.00353295f $X=1.16 $Y=2.57 $X2=0 $Y2=0
cc_208 N_A3_c_214_n N_A_257_414#_c_544_n 0.00534367f $X=1.16 $Y=1.365 $X2=0
+ $Y2=0
cc_209 N_A3_M1003_g N_A_257_414#_c_550_n 0.0143275f $X=1.16 $Y=2.57 $X2=0 $Y2=0
cc_210 N_A3_c_209_n N_VGND_c_583_n 0.0134854f $X=1.395 $Y=0.73 $X2=0 $Y2=0
cc_211 N_A3_c_212_n N_VGND_c_583_n 0.00453864f $X=1.395 $Y=0.805 $X2=0 $Y2=0
cc_212 N_A3_c_209_n N_VGND_c_586_n 0.00486043f $X=1.395 $Y=0.73 $X2=0 $Y2=0
cc_213 N_A3_c_209_n N_VGND_c_588_n 0.00455901f $X=1.395 $Y=0.73 $X2=0 $Y2=0
cc_214 N_A2_c_263_n N_A1_c_307_n 0.0117619f $X=1.7 $Y=1.705 $X2=0 $Y2=0
cc_215 N_A2_M1008_g N_A1_M1000_g 0.0296596f $X=1.69 $Y=2.57 $X2=0 $Y2=0
cc_216 N_A2_M1001_g N_A1_c_308_n 0.0424044f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_217 N_A2_c_268_n N_A1_c_315_n 0.0117619f $X=1.7 $Y=1.87 $X2=0 $Y2=0
cc_218 N_A2_c_264_n A1 0.00437388f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_219 N_A2_c_265_n A1 0.0540841f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_220 N_A2_c_264_n N_A1_c_311_n 0.0117619f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_221 N_A2_c_265_n N_A1_c_311_n 7.52017e-19 $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_222 N_A2_M1001_g N_A1_c_312_n 0.0176854f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_223 N_A2_M1008_g N_VPWR_c_497_n 0.00108285f $X=1.69 $Y=2.57 $X2=0 $Y2=0
cc_224 N_A2_M1008_g N_VPWR_c_498_n 0.0166179f $X=1.69 $Y=2.57 $X2=0 $Y2=0
cc_225 N_A2_M1008_g N_VPWR_c_501_n 0.00803832f $X=1.69 $Y=2.57 $X2=0 $Y2=0
cc_226 N_A2_M1008_g N_VPWR_c_496_n 0.0135635f $X=1.69 $Y=2.57 $X2=0 $Y2=0
cc_227 N_A2_M1008_g N_A_257_414#_c_544_n 9.81754e-19 $X=1.69 $Y=2.57 $X2=0 $Y2=0
cc_228 N_A2_c_268_n N_A_257_414#_c_544_n 2.25414e-19 $X=1.7 $Y=1.87 $X2=0 $Y2=0
cc_229 N_A2_c_265_n N_A_257_414#_c_544_n 0.00449095f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_230 N_A2_M1008_g N_A_257_414#_c_550_n 0.0154098f $X=1.69 $Y=2.57 $X2=0 $Y2=0
cc_231 N_A2_M1008_g N_A_257_414#_c_545_n 0.0184003f $X=1.69 $Y=2.57 $X2=0 $Y2=0
cc_232 N_A2_c_268_n N_A_257_414#_c_545_n 3.36724e-19 $X=1.7 $Y=1.87 $X2=0 $Y2=0
cc_233 N_A2_c_265_n N_A_257_414#_c_545_n 0.020059f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_234 N_A2_M1008_g N_A_257_414#_c_558_n 6.84026e-19 $X=1.69 $Y=2.57 $X2=0 $Y2=0
cc_235 N_A2_M1001_g N_VGND_c_583_n 0.00324405f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_236 N_A2_M1001_g N_VGND_c_586_n 0.00585385f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_237 N_A2_M1001_g N_VGND_c_588_n 0.00639597f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_238 N_A1_c_308_n N_B1_c_361_n 0.0118425f $X=2.177 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_239 N_A1_c_315_n N_B1_M1011_g 0.0156928f $X=2.277 $Y=1.87 $X2=0 $Y2=0
cc_240 N_A1_c_309_n N_B1_c_363_n 0.00696367f $X=2.177 $Y=0.88 $X2=0 $Y2=0
cc_241 A1 N_B1_c_363_n 0.00112807f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_242 N_A1_c_307_n N_B1_c_364_n 0.0156928f $X=2.277 $Y=1.698 $X2=0 $Y2=0
cc_243 A1 N_B1_c_364_n 0.0187503f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_244 N_A1_M1000_g N_B1_c_365_n 2.10892e-19 $X=2.325 $Y=2.57 $X2=0 $Y2=0
cc_245 N_A1_c_315_n N_B1_c_365_n 8.01853e-19 $X=2.277 $Y=1.87 $X2=0 $Y2=0
cc_246 A1 N_B1_c_365_n 0.0481139f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_247 N_A1_c_311_n N_B1_c_365_n 3.78927e-19 $X=2.27 $Y=1.365 $X2=0 $Y2=0
cc_248 A1 N_B1_c_366_n 0.00261851f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_249 N_A1_c_311_n N_B1_c_366_n 0.0156928f $X=2.27 $Y=1.365 $X2=0 $Y2=0
cc_250 N_A1_c_312_n N_B1_c_366_n 0.00856413f $X=2.277 $Y=1.2 $X2=0 $Y2=0
cc_251 N_A1_M1000_g N_VPWR_c_498_n 0.0104853f $X=2.325 $Y=2.57 $X2=0 $Y2=0
cc_252 N_A1_M1000_g N_VPWR_c_503_n 0.00898892f $X=2.325 $Y=2.57 $X2=0 $Y2=0
cc_253 N_A1_M1000_g N_VPWR_c_496_n 0.0162227f $X=2.325 $Y=2.57 $X2=0 $Y2=0
cc_254 N_A1_M1000_g N_A_257_414#_c_550_n 8.85586e-19 $X=2.325 $Y=2.57 $X2=0
+ $Y2=0
cc_255 N_A1_M1000_g N_A_257_414#_c_545_n 0.0191335f $X=2.325 $Y=2.57 $X2=0 $Y2=0
cc_256 N_A1_c_315_n N_A_257_414#_c_545_n 0.00248655f $X=2.277 $Y=1.87 $X2=0
+ $Y2=0
cc_257 A1 N_A_257_414#_c_545_n 0.0283057f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_258 N_A1_M1000_g N_A_257_414#_c_546_n 9.82838e-19 $X=2.325 $Y=2.57 $X2=0
+ $Y2=0
cc_259 A1 N_A_257_414#_c_546_n 0.0290713f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_260 N_A1_M1000_g N_A_257_414#_c_558_n 0.0146152f $X=2.325 $Y=2.57 $X2=0 $Y2=0
cc_261 N_A1_c_308_n N_VGND_c_586_n 0.00549284f $X=2.177 $Y=0.73 $X2=0 $Y2=0
cc_262 N_A1_c_308_n N_VGND_c_588_n 0.00630621f $X=2.177 $Y=0.73 $X2=0 $Y2=0
cc_263 N_B1_c_362_n N_C1_c_419_n 0.00979708f $X=2.965 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_264 N_B1_M1011_g N_C1_M1009_g 0.0251001f $X=2.855 $Y=2.57 $X2=0 $Y2=0
cc_265 N_B1_c_365_n N_C1_M1009_g 0.0130022f $X=3.1 $Y=1.405 $X2=0 $Y2=0
cc_266 N_B1_c_363_n N_C1_c_421_n 0.00979708f $X=2.965 $Y=0.805 $X2=0 $Y2=0
cc_267 N_B1_c_366_n N_C1_c_422_n 0.00662178f $X=2.997 $Y=1.24 $X2=0 $Y2=0
cc_268 N_B1_c_364_n N_C1_c_424_n 0.0370542f $X=3.1 $Y=1.405 $X2=0 $Y2=0
cc_269 N_B1_c_365_n N_C1_c_424_n 7.75152e-19 $X=3.1 $Y=1.405 $X2=0 $Y2=0
cc_270 N_B1_c_364_n N_C1_c_425_n 0.00409483f $X=3.1 $Y=1.405 $X2=0 $Y2=0
cc_271 N_B1_c_365_n N_C1_c_425_n 0.0413195f $X=3.1 $Y=1.405 $X2=0 $Y2=0
cc_272 N_B1_c_366_n N_C1_c_425_n 6.43907e-19 $X=2.997 $Y=1.24 $X2=0 $Y2=0
cc_273 N_B1_M1011_g N_VPWR_c_503_n 0.00844498f $X=2.855 $Y=2.57 $X2=0 $Y2=0
cc_274 N_B1_c_365_n N_VPWR_c_503_n 0.00946574f $X=3.1 $Y=1.405 $X2=0 $Y2=0
cc_275 N_B1_M1011_g N_VPWR_c_496_n 0.0149187f $X=2.855 $Y=2.57 $X2=0 $Y2=0
cc_276 N_B1_c_365_n N_VPWR_c_496_n 0.011217f $X=3.1 $Y=1.405 $X2=0 $Y2=0
cc_277 N_B1_M1011_g N_A_257_414#_c_546_n 0.00352132f $X=2.855 $Y=2.57 $X2=0
+ $Y2=0
cc_278 N_B1_c_365_n N_A_257_414#_c_546_n 0.0129587f $X=3.1 $Y=1.405 $X2=0 $Y2=0
cc_279 N_B1_M1011_g N_A_257_414#_c_558_n 0.0191487f $X=2.855 $Y=2.57 $X2=0 $Y2=0
cc_280 N_B1_c_365_n N_A_257_414#_c_558_n 0.0479915f $X=3.1 $Y=1.405 $X2=0 $Y2=0
cc_281 N_B1_c_365_n A_596_414# 0.0187652f $X=3.1 $Y=1.405 $X2=-0.19 $Y2=-0.245
cc_282 N_B1_c_361_n N_VGND_c_584_n 0.00238433f $X=2.605 $Y=0.73 $X2=0 $Y2=0
cc_283 N_B1_c_362_n N_VGND_c_584_n 0.0126359f $X=2.965 $Y=0.73 $X2=0 $Y2=0
cc_284 N_B1_c_361_n N_VGND_c_586_n 0.00549284f $X=2.605 $Y=0.73 $X2=0 $Y2=0
cc_285 N_B1_c_362_n N_VGND_c_586_n 0.00486043f $X=2.965 $Y=0.73 $X2=0 $Y2=0
cc_286 N_B1_c_363_n N_VGND_c_586_n 6.21075e-19 $X=2.965 $Y=0.805 $X2=0 $Y2=0
cc_287 N_B1_c_361_n N_VGND_c_588_n 0.00617664f $X=2.605 $Y=0.73 $X2=0 $Y2=0
cc_288 N_B1_c_362_n N_VGND_c_588_n 0.00442943f $X=2.965 $Y=0.73 $X2=0 $Y2=0
cc_289 N_B1_c_363_n N_VGND_c_588_n 8.18184e-19 $X=2.965 $Y=0.805 $X2=0 $Y2=0
cc_290 N_C1_M1009_g N_VPWR_c_503_n 0.00898892f $X=3.63 $Y=2.57 $X2=0 $Y2=0
cc_291 N_C1_M1009_g N_VPWR_c_496_n 0.0174031f $X=3.63 $Y=2.57 $X2=0 $Y2=0
cc_292 N_C1_c_419_n N_VGND_c_584_n 0.0126494f $X=3.395 $Y=0.73 $X2=0 $Y2=0
cc_293 N_C1_c_420_n N_VGND_c_584_n 0.00238433f $X=3.755 $Y=0.73 $X2=0 $Y2=0
cc_294 N_C1_c_419_n N_VGND_c_587_n 0.00486043f $X=3.395 $Y=0.73 $X2=0 $Y2=0
cc_295 N_C1_c_420_n N_VGND_c_587_n 0.00549284f $X=3.755 $Y=0.73 $X2=0 $Y2=0
cc_296 N_C1_c_421_n N_VGND_c_587_n 6.21075e-19 $X=3.755 $Y=0.805 $X2=0 $Y2=0
cc_297 N_C1_c_419_n N_VGND_c_588_n 0.00442943f $X=3.395 $Y=0.73 $X2=0 $Y2=0
cc_298 N_C1_c_420_n N_VGND_c_588_n 0.00723412f $X=3.755 $Y=0.73 $X2=0 $Y2=0
cc_299 N_C1_c_421_n N_VGND_c_588_n 8.18184e-19 $X=3.755 $Y=0.805 $X2=0 $Y2=0
cc_300 N_X_c_471_n N_VPWR_c_497_n 0.0681645f $X=0.365 $Y=2.215 $X2=0 $Y2=0
cc_301 N_X_c_470_n N_VPWR_c_499_n 0.0261633f $X=0.365 $Y=2.9 $X2=0 $Y2=0
cc_302 N_X_c_470_n N_VPWR_c_496_n 0.0162464f $X=0.365 $Y=2.9 $X2=0 $Y2=0
cc_303 X A_115_47# 9.46545e-19 $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_304 X N_VGND_c_583_n 0.0317852f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_305 N_X_c_467_n N_VGND_c_585_n 0.0112786f $X=0.19 $Y=0.67 $X2=0 $Y2=0
cc_306 X N_VGND_c_585_n 0.0298725f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_307 N_X_M1014_s N_VGND_c_588_n 0.00233004f $X=0.14 $Y=0.235 $X2=0 $Y2=0
cc_308 N_X_c_467_n N_VGND_c_588_n 0.00657784f $X=0.19 $Y=0.67 $X2=0 $Y2=0
cc_309 X N_VGND_c_588_n 0.0204363f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_310 N_VPWR_c_497_n N_A_257_414#_c_544_n 0.0119061f $X=0.895 $Y=2.215 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_497_n N_A_257_414#_c_550_n 0.0556447f $X=0.895 $Y=2.215 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_498_n N_A_257_414#_c_550_n 0.0438173f $X=1.955 $Y=2.565 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_501_n N_A_257_414#_c_550_n 0.0177952f $X=1.79 $Y=3.33 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_496_n N_A_257_414#_c_550_n 0.0124497f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_315 N_VPWR_M1008_d N_A_257_414#_c_545_n 0.00381132f $X=1.815 $Y=2.07 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_498_n N_A_257_414#_c_545_n 0.0209601f $X=1.955 $Y=2.565 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_498_n N_A_257_414#_c_558_n 0.032976f $X=1.955 $Y=2.565 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_503_n N_A_257_414#_c_558_n 0.0177952f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_496_n N_A_257_414#_c_558_n 0.0124497f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_320 A_115_47# N_VGND_c_588_n 0.00169099f $X=0.575 $Y=0.235 $X2=0 $Y2=0
cc_321 N_VGND_c_588_n A_294_47# 0.00355777f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_322 N_VGND_c_588_n A_372_47# 0.00355777f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_323 N_VGND_c_588_n A_536_47# 0.00311305f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_324 N_VGND_c_588_n A_694_47# 0.00311305f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
