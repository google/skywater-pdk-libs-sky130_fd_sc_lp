* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor3_1 A B C VGND VNB VPB VPWR X
X0 a_1263_295# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_425_117# a_474_313# a_86_305# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 a_86_305# B a_402_411# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 a_474_313# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_1263_295# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_402_411# a_1263_295# a_1363_127# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 VPWR A a_86_305# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND a_1363_127# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_42_411# a_86_305# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_86_305# B a_425_117# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 a_42_411# a_86_305# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_402_411# a_474_313# a_42_411# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_1363_127# C a_402_411# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_425_117# a_1263_295# a_1363_127# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 VGND A a_86_305# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_402_411# a_474_313# a_86_305# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 a_42_411# B a_425_117# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_425_117# a_474_313# a_42_411# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_1363_127# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_474_313# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_42_411# B a_402_411# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_1363_127# C a_425_117# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
