* File: sky130_fd_sc_lp__o211a_0.spice
* Created: Wed Sep  2 10:13:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o211a_0.pex.spice"
.subckt sky130_fd_sc_lp__o211a_0  VNB VPB A1 A2 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A1_M1007_g N_A_257_47#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0609 AS=0.1113 PD=0.71 PS=1.37 NRD=2.856 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_A_257_47#_M1001_d N_A2_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.0609 PD=0.73 PS=0.71 NRD=8.568 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 A_520_47# N_B1_M1004_g N_A_257_47#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0651 PD=0.63 PS=0.73 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_80_21#_M1008_d N_C1_M1008_g A_520_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_80_21#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1152 AS=0.3872 PD=1 PS=2.49 NRD=24.6053 NRS=0 M=1 R=4.26667 SA=75000.5
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1002 A_340_485# N_A1_M1002_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1152 PD=0.85 PS=1 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1000 N_A_80_21#_M1000_d N_A2_M1000_g A_340_485# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1024 AS=0.0672 PD=0.96 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.4
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_B1_M1009_g N_A_80_21#_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=12.2928 M=1 R=4.26667 SA=75001.9
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_80_21#_M1006_d N_C1_M1006_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_483 A_520_47# 0 1.99675e-19 $X=2.6 $Y=0.235
*
.include "sky130_fd_sc_lp__o211a_0.pxi.spice"
*
.ends
*
*
