* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__clkbuf_0 A VGND VNB VPB VPWR X
M1000 a_70_157# A VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.428e+11p ps=1.52e+06u
M1001 VPWR a_70_157# X VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=1.696e+11p ps=1.81e+06u
M1002 VGND a_70_157# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 a_70_157# A VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
.ends
