* File: sky130_fd_sc_lp__sdfsbp_2.spice
* Created: Wed Sep  2 10:35:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfsbp_2.pex.spice"
.subckt sky130_fd_sc_lp__sdfsbp_2  VNB VPB SCE D SCD CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_SCE_M1004_g N_A_27_467#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1027 A_268_47# N_A_27_467#_M1027_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=15.708 M=1 R=2.8 SA=75000.7
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1016 N_A_268_467#_M1016_d N_D_M1016_g A_268_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.10605 AS=0.0441 PD=0.925 PS=0.63 NRD=61.428 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1011 A_471_47# N_SCE_M1011_g N_A_268_467#_M1016_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.10605 PD=0.63 PS=0.925 NRD=14.28 NRS=2.856 M=1 R=2.8 SA=75001.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_SCD_M1012_g A_471_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1023 N_A_629_47#_M1023_d N_CLK_M1023_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1033 N_A_920_73#_M1033_d N_A_629_47#_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1039 N_A_1163_119#_M1039_d N_A_629_47#_M1039_g N_A_268_467#_M1039_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1019 A_1249_119# N_A_920_73#_M1019_g N_A_1163_119#_M1039_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_1291_93#_M1035_g A_1249_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1036 A_1530_119# N_A_1163_119#_M1036_g N_A_1291_93#_M1036_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_SET_B_M1024_g A_1530_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.132458 AS=0.0441 PD=1.0183 PS=0.63 NRD=45.708 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1017 A_1735_119# N_A_1163_119#_M1017_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0944 AS=0.201842 PD=0.935 PS=1.5517 NRD=17.34 NRS=15.936 M=1 R=4.26667
+ SA=75000.9 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1041 N_A_1799_408#_M1041_d N_A_920_73#_M1041_g A_1735_119# VNB NSHORT L=0.15
+ W=0.64 AD=0.130294 AS=0.0944 PD=1.22566 PS=0.935 NRD=7.488 NRS=17.34 M=1
+ R=4.26667 SA=75001.3 SB=75001 A=0.096 P=1.58 MULT=1
MM1032 A_1929_119# N_A_629_47#_M1032_g N_A_1799_408#_M1041_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0855057 PD=0.63 PS=0.80434 NRD=14.28 NRS=15.708 M=1
+ R=2.8 SA=75002.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1038 A_2001_119# N_A_1946_369#_M1038_g A_1929_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75002.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1045 N_VGND_M1045_d N_SET_B_M1045_g A_2001_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_A_1799_408#_M1028_g N_A_1946_369#_M1028_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1078 AS=0.1113 PD=0.853333 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1018 N_Q_N_M1018_d N_A_1799_408#_M1018_g N_VGND_M1028_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2156 PD=1.12 PS=1.70667 NRD=0 NRS=11.424 M=1 R=5.6
+ SA=75000.5 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1037 N_Q_N_M1018_d N_A_1799_408#_M1037_g N_VGND_M1037_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=6.78 M=1 R=5.6 SA=75000.9
+ SB=75000.5 A=0.126 P=1.98 MULT=1
MM1042 N_A_2624_49#_M1042_d N_A_1799_408#_M1042_g N_VGND_M1037_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0896 PD=1.37 PS=0.81 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_2624_49#_M1007_g N_Q_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.273 PD=2.21 PS=1.49 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75001
+ A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_A_2624_49#_M1015_g N_Q_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.273 PD=2.21 PS=1.49 NRD=0 NRS=0 M=1 R=5.6 SA=75001 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1029 N_VPWR_M1029_d N_SCE_M1029_g N_A_27_467#_M1029_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003 A=0.096 P=1.58 MULT=1
MM1005 A_196_467# N_SCE_M1005_g N_VPWR_M1029_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_268_467#_M1008_d N_D_M1008_g A_196_467# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=33.8446 NRS=15.3857 M=1 R=4.26667
+ SA=75001 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1020 A_376_467# N_A_27_467#_M1020_g N_A_268_467#_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1152 AS=0.1248 PD=1 PS=1.03 NRD=38.4741 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1021 N_VPWR_M1021_d N_SCD_M1021_g A_376_467# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2927 AS=0.1152 PD=1.675 PS=1 NRD=123.834 NRS=38.4741 M=1 R=4.26667
+ SA=75002 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1025 N_A_629_47#_M1025_d N_CLK_M1025_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.2927 PD=1.85 PS=1.675 NRD=0 NRS=123.834 M=1 R=4.26667
+ SA=75003 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_920_73#_M1006_d N_A_629_47#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.3691 PD=1.85 PS=2.86 NRD=0 NRS=160.575 M=1 R=4.26667
+ SA=75000.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_1163_119#_M1001_d N_A_920_73#_M1001_g N_A_268_467#_M1001_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1026 A_1275_463# N_A_629_47#_M1026_g N_A_1163_119#_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1034 N_VPWR_M1034_d N_A_1291_93#_M1034_g A_1275_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.110525 AS=0.0441 PD=0.985 PS=0.63 NRD=39.8531 NRS=23.443 M=1 R=2.8
+ SA=75001 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1003 N_A_1291_93#_M1003_d N_A_1163_119#_M1003_g N_VPWR_M1034_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.110525 PD=0.7 PS=0.985 NRD=0 NRS=39.8531 M=1
+ R=2.8 SA=75001.6 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1030 N_VPWR_M1030_d N_SET_B_M1030_g N_A_1291_93#_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.128283 AS=0.0588 PD=1.03 PS=0.7 NRD=105.533 NRS=0 M=1 R=2.8
+ SA=75002 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1013 A_1697_379# N_A_1163_119#_M1013_g N_VPWR_M1030_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.16135 AS=0.256567 PD=1.345 PS=2.06 NRD=32.1307 NRS=19.9167 M=1
+ R=5.6 SA=75001.5 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1031 N_A_1799_408#_M1031_d N_A_629_47#_M1031_g A_1697_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1792 AS=0.16135 PD=1.62 PS=1.345 NRD=0 NRS=32.1307 M=1 R=5.6
+ SA=75001.9 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1043 A_1904_492# N_A_920_73#_M1043_g N_A_1799_408#_M1031_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0896 PD=0.63 PS=0.81 NRD=23.443 NRS=44.5417 M=1 R=2.8
+ SA=75002.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_1946_369#_M1002_g A_1904_492# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.113425 AS=0.0441 PD=1.005 PS=0.63 NRD=37.5088 NRS=23.443 M=1 R=2.8
+ SA=75003.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1000 N_A_1799_408#_M1000_d N_SET_B_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.113425 PD=1.41 PS=1.005 NRD=0 NRS=37.5088 M=1 R=2.8
+ SA=75003.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_1799_408#_M1010_g N_A_1946_369#_M1010_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=80.3169 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1010_d N_A_1799_408#_M1022_g N_Q_N_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.4 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1040 N_VPWR_M1040_d N_A_1799_408#_M1040_g N_Q_N_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.268115 AS=0.1764 PD=2.16853 PS=1.54 NRD=2.3443 NRS=0 M=1 R=8.4
+ SA=75000.8 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1009 N_A_2624_49#_M1009_d N_A_1799_408#_M1009_g N_VPWR_M1040_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.136185 PD=1.81 PS=1.10147 NRD=0 NRS=23.0687 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_Q_M1014_d N_A_2624_49#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1044 N_Q_M1014_d N_A_2624_49#_M1044_g N_VPWR_M1044_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX46_noxref VNB VPB NWDIODE A=29.3551 P=35.21
c_160 VNB 0 1.29912e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__sdfsbp_2.pxi.spice"
*
.ends
*
*
