* File: sky130_fd_sc_lp__nor3_2.pex.spice
* Created: Wed Sep  2 10:09:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3_2%A 3 5 7 8 10 13 15 16 24 25
r47 23 25 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.075 $Y=1.35
+ $X2=1.295 $Y2=1.35
r48 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.075
+ $Y=1.35 $X2=1.075 $Y2=1.35
r49 21 23 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.845 $Y=1.35
+ $X2=1.075 $Y2=1.35
r50 19 21 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=0.52 $Y=1.35
+ $X2=0.845 $Y2=1.35
r51 16 24 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.72 $Y=1.35
+ $X2=1.075 $Y2=1.35
r52 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.35
+ $X2=0.72 $Y2=1.35
r53 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.295 $Y=1.515
+ $X2=1.295 $Y2=1.35
r54 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.295 $Y=1.515
+ $X2=1.295 $Y2=2.465
r55 8 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.295 $Y=1.185
+ $X2=1.295 $Y2=1.35
r56 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.295 $Y=1.185
+ $X2=1.295 $Y2=0.655
r57 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.845 $Y=1.185
+ $X2=0.845 $Y2=1.35
r58 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.845 $Y=1.185
+ $X2=0.845 $Y2=0.655
r59 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.515
+ $X2=0.52 $Y2=1.35
r60 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.52 $Y=1.515 $X2=0.52
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_2%B 3 7 9 11 14 19 20 24 25 36 39 46 48
r78 39 48 1.67451 $w=4.98e-07 $l=7e-08 $layer=LI1_cond $X=3.19 $Y=1.535 $X2=3.12
+ $Y2=1.535
r79 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.45 $X2=3.57 $Y2=1.45
r80 34 36 26.5143 $w=4.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.365 $Y=1.4
+ $X2=3.57 $Y2=1.4
r81 32 34 38.8014 $w=4.3e-07 $l=3e-07 $layer=POLY_cond $X=3.065 $Y=1.4 $X2=3.365
+ $Y2=1.4
r82 25 37 0.717647 $w=4.98e-07 $l=3e-08 $layer=LI1_cond $X=3.6 $Y=1.535 $X2=3.57
+ $Y2=1.535
r83 24 48 0.191373 $w=4.98e-07 $l=8e-09 $layer=LI1_cond $X=3.112 $Y=1.535
+ $X2=3.12 $Y2=1.535
r84 24 46 9.28579 $w=4.98e-07 $l=1.72e-07 $layer=LI1_cond $X=3.112 $Y=1.535
+ $X2=2.94 $Y2=1.535
r85 24 37 8.92274 $w=4.98e-07 $l=3.73e-07 $layer=LI1_cond $X=3.197 $Y=1.535
+ $X2=3.57 $Y2=1.535
r86 24 39 0.167451 $w=4.98e-07 $l=7e-09 $layer=LI1_cond $X=3.197 $Y=1.535
+ $X2=3.19 $Y2=1.535
r87 20 31 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.51
+ $X2=1.75 $Y2=1.675
r88 20 30 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.51
+ $X2=1.75 $Y2=1.345
r89 19 22 10.2591 $w=1.98e-07 $l=1.85e-07 $layer=LI1_cond $X=1.77 $Y=1.51
+ $X2=1.77 $Y2=1.695
r90 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.755
+ $Y=1.51 $X2=1.755 $Y2=1.51
r91 17 22 1.35108 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=1.87 $Y=1.695 $X2=1.77
+ $Y2=1.695
r92 17 46 65.9293 $w=1.78e-07 $l=1.07e-06 $layer=LI1_cond $X=1.87 $Y=1.695
+ $X2=2.94 $Y2=1.695
r93 12 34 27.6395 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.365 $Y=1.615
+ $X2=3.365 $Y2=1.4
r94 12 14 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=3.365 $Y=1.615
+ $X2=3.365 $Y2=2.465
r95 9 32 27.6395 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.065 $Y=1.185
+ $X2=3.065 $Y2=1.4
r96 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.065 $Y=1.185
+ $X2=3.065 $Y2=0.655
r97 7 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.725 $Y=2.465
+ $X2=1.725 $Y2=1.675
r98 3 30 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.725 $Y=0.655
+ $X2=1.725 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_2%C 1 3 4 6 7 9 10 12 13 14 22
r51 20 22 24.2745 $w=5.4e-07 $l=2.45e-07 $layer=POLY_cond $X=2.39 $Y=1.455
+ $X2=2.635 $Y2=1.455
r52 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.39
+ $Y=1.35 $X2=2.39 $Y2=1.35
r53 17 20 18.3297 $w=5.4e-07 $l=1.85e-07 $layer=POLY_cond $X=2.205 $Y=1.455
+ $X2=2.39 $Y2=1.455
r54 14 21 12.8049 $w=2.23e-07 $l=2.5e-07 $layer=LI1_cond $X=2.64 $Y=1.322
+ $X2=2.39 $Y2=1.322
r55 13 21 11.7805 $w=2.23e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=1.322
+ $X2=2.39 $Y2=1.322
r56 10 22 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.635 $Y=1.725
+ $X2=2.635 $Y2=1.455
r57 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.635 $Y=1.725
+ $X2=2.635 $Y2=2.465
r58 7 22 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.635 $Y=1.185
+ $X2=2.635 $Y2=1.455
r59 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.635 $Y=1.185
+ $X2=2.635 $Y2=0.655
r60 4 17 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.205 $Y=1.725
+ $X2=2.205 $Y2=1.455
r61 4 6 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.205 $Y=1.725
+ $X2=2.205 $Y2=2.465
r62 1 17 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.205 $Y=1.185
+ $X2=2.205 $Y2=1.455
r63 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.205 $Y=1.185
+ $X2=2.205 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_2%A_36_367# 1 2 3 12 16 17 19 20 21 24 26 29 30
+ 31 32 34 37
r68 32 39 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=2.125
+ $X2=3.615 $Y2=2.04
r69 32 34 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.615 $Y=2.125
+ $X2=3.615 $Y2=2.495
r70 30 39 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.485 $Y=2.04
+ $X2=3.615 $Y2=2.04
r71 30 31 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.485 $Y=2.04
+ $X2=2.845 $Y2=2.04
r72 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.76 $Y=2.125
+ $X2=2.845 $Y2=2.04
r73 28 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.76 $Y=2.125
+ $X2=2.76 $Y2=2.465
r74 27 37 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.605 $Y=2.555
+ $X2=1.51 $Y2=2.555
r75 26 29 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.675 $Y=2.555
+ $X2=2.76 $Y2=2.465
r76 26 27 65.9293 $w=1.78e-07 $l=1.07e-06 $layer=LI1_cond $X=2.675 $Y=2.555
+ $X2=1.605 $Y2=2.555
r77 22 37 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=1.51 $Y=2.645 $X2=1.51
+ $Y2=2.555
r78 22 24 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=1.51 $Y=2.645
+ $X2=1.51 $Y2=2.91
r79 20 37 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.415 $Y=2.555
+ $X2=1.51 $Y2=2.555
r80 20 21 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=1.415 $Y=2.555
+ $X2=1.16 $Y2=2.555
r81 19 21 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.075 $Y=2.465
+ $X2=1.16 $Y2=2.555
r82 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.075 $Y=1.855
+ $X2=1.075 $Y2=2.465
r83 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.99 $Y=1.77
+ $X2=1.075 $Y2=1.855
r84 16 17 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=0.99 $Y=1.77
+ $X2=0.41 $Y2=1.77
r85 12 14 39.6953 $w=2.68e-07 $l=9.3e-07 $layer=LI1_cond $X=0.275 $Y=1.98
+ $X2=0.275 $Y2=2.91
r86 10 17 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.275 $Y=1.855
+ $X2=0.41 $Y2=1.77
r87 10 12 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.275 $Y=1.855
+ $X2=0.275 $Y2=1.98
r88 3 39 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.835 $X2=3.58 $Y2=2.04
r89 3 34 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=3.44
+ $Y=1.835 $X2=3.58 $Y2=2.495
r90 2 37 600 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_PDIFF $count=1 $X=1.37
+ $Y=1.835 $X2=1.51 $Y2=2.55
r91 2 24 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.37
+ $Y=1.835 $X2=1.51 $Y2=2.91
r92 1 14 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.835 $X2=0.305 $Y2=2.91
r93 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.835 $X2=0.305 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_2%VPWR 1 6 8 17 18 21 32
r49 30 32 7.76391 $w=5.98e-07 $l=4.5e-08 $layer=LI1_cond $X=1.2 $Y=3.115
+ $X2=1.245 $Y2=3.115
r50 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 28 30 2.39216 $w=5.98e-07 $l=1.2e-07 $layer=LI1_cond $X=1.08 $Y=3.115
+ $X2=1.2 $Y2=3.115
r52 26 28 6.87745 $w=5.98e-07 $l=3.45e-07 $layer=LI1_cond $X=0.735 $Y=3.115
+ $X2=1.08 $Y2=3.115
r53 24 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 23 26 0.29902 $w=5.98e-07 $l=1.5e-08 $layer=LI1_cond $X=0.72 $Y=3.115
+ $X2=0.735 $Y2=3.115
r55 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 20 23 0.398693 $w=5.98e-07 $l=2e-08 $layer=LI1_cond $X=0.7 $Y=3.115 $X2=0.72
+ $Y2=3.115
r57 20 21 9.25901 $w=5.98e-07 $l=1.2e-07 $layer=LI1_cond $X=0.7 $Y=3.115
+ $X2=0.58 $Y2=3.115
r58 17 32 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=1.245 $Y2=3.33
r59 17 18 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 13 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 12 21 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=0.58 $Y2=3.33
r62 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 8 18 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.6 $Y2=3.33
r64 8 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33 $X2=1.2
+ $Y2=3.33
r65 4 20 6.14847 $w=2.4e-07 $l=3e-07 $layer=LI1_cond $X=0.7 $Y=2.815 $X2=0.7
+ $Y2=3.115
r66 4 6 30.0115 $w=2.38e-07 $l=6.25e-07 $layer=LI1_cond $X=0.7 $Y=2.815 $X2=0.7
+ $Y2=2.19
r67 1 28 600 $w=1.7e-07 $l=1.33566e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.835 $X2=1.08 $Y2=2.95
r68 1 26 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.835 $X2=0.735 $Y2=2.95
r69 1 6 300 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.835 $X2=0.735 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_2%A_360_367# 1 2 7 15
r21 13 15 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=3.165 $Y=2.815
+ $X2=3.165 $Y2=2.46
r22 9 12 40.3355 $w=2.58e-07 $l=9.1e-07 $layer=LI1_cond $X=1.94 $Y=2.945
+ $X2=2.85 $Y2=2.945
r23 7 13 6.86182 $w=2.6e-07 $l=2.04939e-07 $layer=LI1_cond $X=3.015 $Y=2.945
+ $X2=3.165 $Y2=2.815
r24 7 12 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=2.945
+ $X2=2.85 $Y2=2.945
r25 2 15 600 $w=1.7e-07 $l=8.15858e-07 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.835 $X2=3.15 $Y2=2.46
r26 2 12 600 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.835 $X2=2.85 $Y2=2.94
r27 1 9 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.8
+ $Y=1.835 $X2=1.94 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_2%Y 1 2 3 4 14 15 17 21 23 24 25 26 33 34 39 43
+ 48
r67 37 39 4.15909 $w=1.98e-07 $l=7.5e-08 $layer=LI1_cond $X=2.085 $Y=0.94
+ $X2=2.16 $Y2=0.94
r68 34 54 5.30787 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=0.94 $X2=1.415
+ $Y2=0.94
r69 26 33 5.99569 $w=2e-07 $l=1.2e-07 $layer=LI1_cond $X=1.965 $Y=0.94 $X2=1.845
+ $Y2=0.94
r70 26 37 5.99569 $w=2e-07 $l=1.2e-07 $layer=LI1_cond $X=1.965 $Y=0.94 $X2=2.085
+ $Y2=0.94
r71 26 48 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=1.965 $Y=0.84
+ $X2=1.965 $Y2=0.42
r72 26 39 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=2.165 $Y=0.94
+ $X2=2.16 $Y2=0.94
r73 25 33 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=0.94 $X2=1.845
+ $Y2=0.94
r74 25 34 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=0.94 $X2=1.5
+ $Y2=0.94
r75 24 54 14.4121 $w=1.82e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=0.94
+ $X2=1.415 $Y2=0.94
r76 24 43 18.5268 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.07 $Y=0.84
+ $X2=1.07 $Y2=0.42
r77 23 26 32.7182 $w=1.98e-07 $l=5.9e-07 $layer=LI1_cond $X=2.755 $Y=0.94
+ $X2=2.165 $Y2=0.94
r78 19 23 6.84722 $w=2e-07 $l=1.54091e-07 $layer=LI1_cond $X=2.867 $Y=0.84
+ $X2=2.755 $Y2=0.94
r79 19 21 21.5123 $w=2.23e-07 $l=4.2e-07 $layer=LI1_cond $X=2.867 $Y=0.84
+ $X2=2.867 $Y2=0.42
r80 15 17 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=1.5 $Y=2.13 $X2=2.42
+ $Y2=2.13
r81 14 15 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.415 $Y=1.965
+ $X2=1.5 $Y2=2.13
r82 13 54 1.129 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.415 $Y=1.04 $X2=1.415
+ $Y2=0.94
r83 13 14 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.415 $Y=1.04
+ $X2=1.415 $Y2=1.965
r84 4 17 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=2.13
r85 3 21 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.71
+ $Y=0.235 $X2=2.85 $Y2=0.42
r86 2 26 182 $w=1.7e-07 $l=7.68082e-07 $layer=licon1_NDIFF $count=1 $X=1.8
+ $Y=0.235 $X2=1.965 $Y2=0.925
r87 2 48 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.8
+ $Y=0.235 $X2=1.965 $Y2=0.42
r88 1 43 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.92
+ $Y=0.235 $X2=1.06 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_2%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37 39
+ 40 41 57 58
r60 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r61 55 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r62 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r63 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r64 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r65 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r66 45 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r67 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r68 41 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r69 41 49 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r70 39 54 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.15 $Y=0 $X2=3.12
+ $Y2=0
r71 39 40 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=3.15 $Y=0 $X2=3.297
+ $Y2=0
r72 38 57 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.6
+ $Y2=0
r73 38 40 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.297
+ $Y2=0
r74 36 51 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.16
+ $Y2=0
r75 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.42
+ $Y2=0
r76 35 54 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.585 $Y=0 $X2=3.12
+ $Y2=0
r77 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.42
+ $Y2=0
r78 33 48 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.2
+ $Y2=0
r79 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.51
+ $Y2=0
r80 32 51 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=2.16
+ $Y2=0
r81 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.51
+ $Y2=0
r82 30 44 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.24
+ $Y2=0
r83 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.63
+ $Y2=0
r84 29 48 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.2
+ $Y2=0
r85 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.63
+ $Y2=0
r86 25 40 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.297 $Y=0.085
+ $X2=3.297 $Y2=0
r87 25 27 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=3.297 $Y=0.085
+ $X2=3.297 $Y2=0.38
r88 21 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=0.085
+ $X2=2.42 $Y2=0
r89 21 23 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.42 $Y=0.085
+ $X2=2.42 $Y2=0.545
r90 17 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=0.085
+ $X2=1.51 $Y2=0
r91 17 19 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.51 $Y=0.085
+ $X2=1.51 $Y2=0.545
r92 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.085
+ $X2=0.63 $Y2=0
r93 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.63 $Y=0.085
+ $X2=0.63 $Y2=0.38
r94 4 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.14
+ $Y=0.235 $X2=3.28 $Y2=0.38
r95 3 23 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.235 $X2=2.42 $Y2=0.545
r96 2 19 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=1.37
+ $Y=0.235 $X2=1.51 $Y2=0.545
r97 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.505
+ $Y=0.235 $X2=0.63 $Y2=0.38
.ends

