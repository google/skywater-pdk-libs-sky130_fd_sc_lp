* File: sky130_fd_sc_lp__o2bb2a_m.pex.spice
* Created: Wed Sep  2 10:21:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%A_85_187# 1 2 9 13 17 18 21 22 24 25 28 31
+ 32 36
c73 36 0 9.13536e-20 $X=2.505 $Y=2.835
c74 32 0 1.8647e-19 $X=2.207 $Y=1.66
r75 33 36 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.29 $Y=2.835
+ $X2=2.505 $Y2=2.835
r76 31 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=2.67
+ $X2=2.29 $Y2=2.835
r77 30 32 4.70473 $w=1.9e-07 $l=1.19499e-07 $layer=LI1_cond $X=2.29 $Y=1.745
+ $X2=2.207 $Y2=1.66
r78 30 31 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.29 $Y=1.745
+ $X2=2.29 $Y2=2.67
r79 26 32 4.70473 $w=1.9e-07 $l=1.11781e-07 $layer=LI1_cond $X=2.145 $Y=1.575
+ $X2=2.207 $Y2=1.66
r80 26 28 24.5584 $w=2.08e-07 $l=4.65e-07 $layer=LI1_cond $X=2.145 $Y=1.575
+ $X2=2.145 $Y2=1.11
r81 24 32 1.74598 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.04 $Y=1.66
+ $X2=2.207 $Y2=1.66
r82 24 25 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=2.04 $Y=1.66
+ $X2=0.675 $Y2=1.66
r83 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59 $Y=1.1
+ $X2=0.59 $Y2=1.1
r84 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.59 $Y=1.575
+ $X2=0.675 $Y2=1.66
r85 19 21 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.59 $Y=1.575
+ $X2=0.59 $Y2=1.1
r86 17 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.59 $Y=1.44
+ $X2=0.59 $Y2=1.1
r87 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.44
+ $X2=0.59 $Y2=1.605
r88 16 22 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=0.935
+ $X2=0.59 $Y2=1.1
r89 13 16 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.61 $Y=0.445
+ $X2=0.61 $Y2=0.935
r90 9 18 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=0.5 $Y=2.885 $X2=0.5
+ $Y2=1.605
r91 2 36 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=2.675 $X2=2.505 $Y2=2.835
r92 1 28 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.835 $X2=2.145 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%A1_N 3 7 11 12 13 14 18 19
c45 3 0 9.25659e-20 $X=0.97 $Y=2.885
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.95
+ $Y=2.01 $X2=0.95 $Y2=2.01
r47 13 14 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.875 $Y=2.035
+ $X2=0.875 $Y2=2.405
r48 13 19 0.622958 $w=4.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.875 $Y=2.035
+ $X2=0.875 $Y2=2.01
r49 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.95 $Y=2.35
+ $X2=0.95 $Y2=2.01
r50 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.35
+ $X2=0.95 $Y2=2.515
r51 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.845
+ $X2=0.95 $Y2=2.01
r52 7 10 717.872 $w=1.5e-07 $l=1.4e-06 $layer=POLY_cond $X=1.04 $Y=0.445
+ $X2=1.04 $Y2=1.845
r53 3 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.97 $Y=2.885
+ $X2=0.97 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%A2_N 3 7 11 12 13 14 15 20
c43 20 0 2.60315e-20 $X=1.49 $Y=0.955
r44 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.49
+ $Y=0.955 $X2=1.49 $Y2=0.955
r45 15 21 7.53086 $w=5.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.385 $Y=1.295
+ $X2=1.385 $Y2=0.955
r46 14 21 0.664488 $w=5.38e-07 $l=3e-08 $layer=LI1_cond $X=1.385 $Y=0.925
+ $X2=1.385 $Y2=0.955
r47 13 14 8.19535 $w=5.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.385 $Y=0.555
+ $X2=1.385 $Y2=0.925
r48 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.49 $Y=1.295
+ $X2=1.49 $Y2=0.955
r49 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.295
+ $X2=1.49 $Y2=1.46
r50 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=0.79
+ $X2=1.49 $Y2=0.955
r51 7 12 730.691 $w=1.5e-07 $l=1.425e-06 $layer=POLY_cond $X=1.4 $Y=2.885
+ $X2=1.4 $Y2=1.46
r52 3 10 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.4 $Y=0.445 $X2=1.4
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%A_209_535# 1 2 7 9 14 16 17 18 21 28 29 34
c71 34 0 9.25659e-20 $X=1.43 $Y=2.835
r72 32 34 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.185 $Y=2.835
+ $X2=1.43 $Y2=2.835
r73 29 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=0.44
+ $X2=2.34 $Y2=0.605
r74 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.34
+ $Y=0.44 $X2=2.34 $Y2=0.44
r75 25 28 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.92 $Y=0.44
+ $X2=2.34 $Y2=0.44
r76 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.86
+ $Y=2.01 $X2=1.86 $Y2=2.01
r77 19 21 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.86 $Y=2.265
+ $X2=1.86 $Y2=2.01
r78 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.695 $Y=2.35
+ $X2=1.86 $Y2=2.265
r79 17 18 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.695 $Y=2.35
+ $X2=1.515 $Y2=2.35
r80 16 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.43 $Y=2.67
+ $X2=1.43 $Y2=2.835
r81 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.43 $Y=2.435
+ $X2=1.515 $Y2=2.35
r82 15 16 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.43 $Y=2.435
+ $X2=1.43 $Y2=2.67
r83 14 39 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.36 $Y=1.045
+ $X2=2.36 $Y2=0.605
r84 12 22 46.8536 $w=6.85e-07 $l=3.68375e-07 $layer=POLY_cond $X=2.36 $Y=1.845
+ $X2=2.065 $Y2=2.01
r85 12 14 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.36 $Y=1.845 $X2=2.36
+ $Y2=1.045
r86 7 22 70.7777 $w=6.85e-07 $l=6.07166e-07 $layer=POLY_cond $X=2.29 $Y=2.515
+ $X2=2.065 $Y2=2.01
r87 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.29 $Y=2.515 $X2=2.29
+ $Y2=2.885
r88 2 32 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=2.675 $X2=1.185 $Y2=2.835
r89 1 25 182 $w=1.7e-07 $l=5.3782e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=1.92 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%B2 3 7 11 12 13 14 15 20
c41 20 0 1.8647e-19 $X=2.81 $Y=1.665
c42 3 0 9.13536e-20 $X=2.72 $Y=2.885
r43 14 15 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.765 $Y=2.035
+ $X2=2.765 $Y2=2.405
r44 13 14 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.765 $Y=1.665
+ $X2=2.765 $Y2=2.035
r45 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.81
+ $Y=1.665 $X2=2.81 $Y2=1.665
r46 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.81 $Y=2.005
+ $X2=2.81 $Y2=1.665
r47 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=2.005
+ $X2=2.81 $Y2=2.17
r48 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.5
+ $X2=2.81 $Y2=1.665
r49 7 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.79 $Y=1.045
+ $X2=2.79 $Y2=1.5
r50 3 12 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=2.72 $Y=2.885
+ $X2=2.72 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%B1 1 3 6 11 15 16 17 22
r31 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.35
+ $Y=1.865 $X2=3.35 $Y2=1.865
r32 16 17 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.475 $Y=2.035
+ $X2=3.475 $Y2=2.405
r33 16 23 4.66465 $w=4.18e-07 $l=1.7e-07 $layer=LI1_cond $X=3.475 $Y=2.035
+ $X2=3.475 $Y2=1.865
r34 15 23 5.48782 $w=4.18e-07 $l=2e-07 $layer=LI1_cond $X=3.475 $Y=1.665
+ $X2=3.475 $Y2=1.865
r35 14 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=1.7
+ $X2=3.35 $Y2=1.865
r36 11 22 95.2994 $w=3.3e-07 $l=5.45e-07 $layer=POLY_cond $X=3.35 $Y=2.41
+ $X2=3.35 $Y2=1.865
r37 8 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.08 $Y=2.485
+ $X2=3.35 $Y2=2.485
r38 6 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=3.26 $Y=1.045
+ $X2=3.26 $Y2=1.7
r39 1 8 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.08 $Y=2.56 $X2=3.08
+ $Y2=2.485
r40 1 3 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.08 $Y=2.56 $X2=3.08
+ $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%X 1 2 9 12 13 14 15 16 17 36
r19 16 17 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.405
r20 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r21 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r22 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.295
r23 13 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=0.675
r24 12 40 6.97622 $w=3.43e-07 $l=1.2e-07 $layer=LI1_cond $X=0.327 $Y=0.555
+ $X2=0.327 $Y2=0.675
r25 12 36 1.50319 $w=3.43e-07 $l=4.5e-08 $layer=LI1_cond $X=0.327 $Y=0.555
+ $X2=0.327 $Y2=0.51
r26 10 17 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.24 $Y=2.655
+ $X2=0.24 $Y2=2.405
r27 9 10 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=2.82
+ $X2=0.272 $Y2=2.655
r28 2 9 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.675 $X2=0.285 $Y2=2.82
r29 1 36 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.235 $X2=0.395 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%VPWR 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r54 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r57 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 40 43 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r60 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 38 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=0.735 $Y2=3.33
r64 35 37 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=1.68
+ $Y2=3.33
r65 33 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r67 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.735 $Y2=3.33
r68 30 32 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 28 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 28 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 26 43 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.13 $Y=3.33 $X2=3.12
+ $Y2=3.33
r72 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=3.33
+ $X2=3.295 $Y2=3.33
r73 25 46 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.46 $Y=3.33 $X2=3.6
+ $Y2=3.33
r74 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=3.33
+ $X2=3.295 $Y2=3.33
r75 23 37 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.86 $Y2=3.33
r77 22 40 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.86 $Y2=3.33
r79 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=3.245
+ $X2=3.295 $Y2=3.33
r80 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.295 $Y=3.245
+ $X2=3.295 $Y2=2.95
r81 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=3.245
+ $X2=1.86 $Y2=3.33
r82 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.86 $Y=3.245
+ $X2=1.86 $Y2=2.95
r83 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r84 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.95
r85 3 20 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=2.675 $X2=3.295 $Y2=2.95
r86 2 16 600 $w=1.7e-07 $l=5.04083e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=2.675 $X2=1.86 $Y2=2.95
r87 1 12 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.675 $X2=0.735 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%VGND 1 2 11 15 18 19 20 30 31 34
c38 31 0 2.60315e-20 $X=3.6 $Y=0
r39 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r41 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r42 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r44 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r45 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 22 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=0.825
+ $Y2=0
r47 22 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=1.2
+ $Y2=0
r48 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r49 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r50 18 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.64
+ $Y2=0
r51 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=3.025
+ $Y2=0
r52 17 30 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.6
+ $Y2=0
r53 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.025
+ $Y2=0
r54 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.025 $Y=0.085
+ $X2=3.025 $Y2=0
r55 13 15 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=3.025 $Y=0.085
+ $X2=3.025 $Y2=0.96
r56 9 34 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r57 9 11 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.38
r58 2 15 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.835 $X2=3.025 $Y2=0.96
r59 1 11 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.685
+ $Y=0.235 $X2=0.825 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_M%A_487_167# 1 2 9 11 12
r15 13 15 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=3.475 $Y=1.225
+ $X2=3.475 $Y2=1.11
r16 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.37 $Y=1.31
+ $X2=3.475 $Y2=1.225
r17 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.37 $Y=1.31 $X2=2.68
+ $Y2=1.31
r18 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.575 $Y=1.225
+ $X2=2.68 $Y2=1.31
r19 7 9 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.575 $Y=1.225
+ $X2=2.575 $Y2=1.11
r20 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.835 $X2=3.475 $Y2=1.11
r21 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.835 $X2=2.575 $Y2=1.11
.ends

