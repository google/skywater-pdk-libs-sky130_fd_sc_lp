# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__a211o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.310000 1.425000 5.640000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.770000 1.425000 5.100000 1.820000 ;
        RECT 4.900000 1.820000 5.100000 1.950000 ;
        RECT 4.900000 1.950000 6.125000 2.120000 ;
        RECT 5.915000 1.345000 6.500000 1.645000 ;
        RECT 5.915000 1.645000 6.125000 1.950000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 1.345000 3.205000 1.695000 ;
        RECT 2.815000 1.695000 4.450000 1.865000 ;
        RECT 4.120000 1.415000 4.450000 1.695000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 1.185000 3.710000 1.515000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.188600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.390000 0.405000 1.055000 ;
        RECT 0.090000 1.055000 2.305000 1.225000 ;
        RECT 0.090000 1.225000 0.345000 1.755000 ;
        RECT 0.090000 1.755000 1.760000 1.925000 ;
        RECT 0.710000 1.925000 0.900000 3.075000 ;
        RECT 1.265000 0.255000 1.455000 1.045000 ;
        RECT 1.265000 1.045000 2.305000 1.055000 ;
        RECT 1.570000 1.925000 1.760000 3.075000 ;
        RECT 2.125000 0.255000 2.305000 1.045000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.210000  2.095000 0.540000 3.245000 ;
      RECT 0.515000  1.395000 2.645000 1.585000 ;
      RECT 0.765000  0.085000 1.095000 0.885000 ;
      RECT 1.070000  2.105000 1.400000 3.245000 ;
      RECT 1.625000  0.085000 1.955000 0.875000 ;
      RECT 1.930000  1.815000 2.260000 3.245000 ;
      RECT 2.475000  0.985000 4.110000 1.015000 ;
      RECT 2.475000  1.015000 3.205000 1.155000 ;
      RECT 2.475000  1.155000 2.645000 1.395000 ;
      RECT 2.475000  1.585000 2.645000 2.035000 ;
      RECT 2.475000  2.035000 3.785000 2.205000 ;
      RECT 2.500000  0.085000 2.830000 0.805000 ;
      RECT 2.595000  2.375000 2.925000 2.425000 ;
      RECT 2.595000  2.425000 6.625000 2.460000 ;
      RECT 2.595000  2.460000 4.725000 2.595000 ;
      RECT 2.595000  2.595000 2.855000 3.075000 ;
      RECT 3.000000  0.255000 3.205000 0.845000 ;
      RECT 3.000000  0.845000 4.110000 0.985000 ;
      RECT 3.025000  2.765000 4.215000 3.055000 ;
      RECT 3.375000  0.085000 3.705000 0.675000 ;
      RECT 3.455000  2.205000 3.785000 2.255000 ;
      RECT 3.875000  0.255000 4.110000 0.845000 ;
      RECT 3.885000  1.015000 4.110000 1.065000 ;
      RECT 3.885000  1.065000 5.695000 1.235000 ;
      RECT 4.280000  0.085000 4.835000 0.885000 ;
      RECT 4.355000  2.035000 4.730000 2.290000 ;
      RECT 4.355000  2.290000 6.625000 2.425000 ;
      RECT 4.385000  2.595000 4.725000 3.075000 ;
      RECT 4.895000  2.630000 5.225000 3.245000 ;
      RECT 5.005000  0.255000 6.195000 0.425000 ;
      RECT 5.005000  0.425000 5.335000 0.895000 ;
      RECT 5.435000  2.460000 5.695000 3.075000 ;
      RECT 5.505000  0.595000 5.695000 1.065000 ;
      RECT 5.865000  0.425000 6.195000 1.095000 ;
      RECT 5.865000  2.630000 6.195000 3.245000 ;
      RECT 6.295000  1.815000 6.625000 2.290000 ;
      RECT 6.365000  0.085000 6.625000 1.095000 ;
      RECT 6.365000  2.460000 6.625000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__a211o_4
END LIBRARY
