* File: sky130_fd_sc_lp__o22a_m.spice
* Created: Fri Aug 28 11:10:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22a_m.pex.spice"
.subckt sky130_fd_sc_lp__o22a_m  VNB VPB A1 B1 B2 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* B2	B2
* B1	B1
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_88_187#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.1197 PD=0.84 PS=1.41 NRD=17.136 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1007 N_A_237_81#_M1007_d N_A1_M1007_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0882 PD=0.78 PS=0.84 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.8
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_88_187#_M1008_d N_B1_M1008_g N_A_237_81#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75001.3 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_237_81#_M1009_d N_B2_M1009_g N_A_88_187#_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75001.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_237_81#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1449 AS=0.0756 PD=1.53 PS=0.78 NRD=22.848 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_88_187#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.20055 AS=0.1197 PD=1.375 PS=1.41 NRD=0 NRS=9.3772 M=1 R=2.8 SA=75000.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1004 A_339_535# N_B1_M1004_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.20055 PD=0.63 PS=1.375 NRD=23.443 NRS=316.599 M=1 R=2.8
+ SA=75001.3 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_A_88_187#_M1001_d N_B2_M1001_g A_339_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 A_519_535# N_A2_M1006_g N_A_88_187#_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=51.5943 M=1 R=2.8
+ SA=75002.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g A_519_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o22a_m.pxi.spice"
*
.ends
*
*
