* NGSPICE file created from sky130_fd_sc_lp__a32oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_58_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.1214e+12p ps=9.34e+06u
M1001 a_326_69# A1 Y VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=3.36e+11p ps=2.48e+06u
M1002 a_58_367# B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A3 a_58_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.1151e+12p pd=6.81e+06u as=0p ps=0u
M1004 Y B1 a_141_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.89e+11p ps=2.13e+06u
M1005 VPWR A1 a_58_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_141_69# B2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.452e+11p ps=4.42e+06u
M1007 a_58_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_434_69# A2 a_326_69# VNB nshort w=840000u l=150000u
+  ad=3.696e+11p pd=2.56e+06u as=0p ps=0u
M1009 VGND A3 a_434_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

