# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nor2_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.210000 1.525000 1.560000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.425000 4.165000 1.760000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.646400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.825000 0.265000 1.015000 0.870000 ;
        RECT 0.825000 0.870000 1.910000 1.040000 ;
        RECT 1.685000 0.265000 1.910000 0.870000 ;
        RECT 1.695000 1.040000 1.910000 1.325000 ;
        RECT 1.695000 1.325000 2.735000 1.560000 ;
        RECT 2.505000 1.560000 2.735000 1.950000 ;
        RECT 2.505000 1.950000 3.635000 2.120000 ;
        RECT 2.505000 2.120000 2.780000 2.735000 ;
        RECT 2.510000 0.265000 2.735000 1.085000 ;
        RECT 2.510000 1.085000 3.625000 1.255000 ;
        RECT 2.510000 1.255000 2.735000 1.325000 ;
        RECT 3.375000 2.120000 3.635000 2.735000 ;
        RECT 3.405000 0.265000 3.625000 1.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
        RECT 0.325000  0.085000 0.655000 1.040000 ;
        RECT 1.185000  0.085000 1.515000 0.700000 ;
        RECT 2.080000  0.085000 2.340000 1.155000 ;
        RECT 2.905000  0.085000 3.235000 0.915000 ;
        RECT 3.795000  0.085000 4.095000 1.140000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.320000 3.415000 ;
        RECT 0.755000 2.095000 1.085000 3.245000 ;
        RECT 1.615000 2.095000 1.945000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.325000 1.730000 2.335000 1.925000 ;
      RECT 0.325000 1.925000 0.585000 3.075000 ;
      RECT 1.255000 1.925000 1.445000 3.075000 ;
      RECT 2.115000 1.925000 2.335000 2.905000 ;
      RECT 2.115000 2.905000 4.095000 3.075000 ;
      RECT 2.950000 2.290000 3.205000 2.905000 ;
      RECT 3.805000 1.930000 4.095000 2.905000 ;
  END
END sky130_fd_sc_lp__nor2_4
