# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nor4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__nor4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.345000 2.135000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.345000 1.210000 4.375000 1.535000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 1.210000 6.085000 1.535000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.305000 1.210000 7.145000 1.355000 ;
        RECT 6.305000 1.355000 7.655000 1.525000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.587200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.255000 1.080000 1.005000 ;
        RECT 0.865000 1.005000 8.070000 1.040000 ;
        RECT 0.865000 1.040000 1.930000 1.175000 ;
        RECT 1.750000 0.255000 1.940000 0.870000 ;
        RECT 1.750000 0.870000 7.550000 1.005000 ;
        RECT 3.055000 0.265000 3.250000 0.870000 ;
        RECT 3.920000 0.265000 4.110000 0.870000 ;
        RECT 4.780000 0.265000 4.970000 0.870000 ;
        RECT 5.640000 0.265000 5.830000 0.870000 ;
        RECT 6.500000 0.265000 6.690000 0.870000 ;
        RECT 6.500000 1.695000 8.070000 1.875000 ;
        RECT 6.500000 1.875000 6.690000 2.735000 ;
        RECT 7.315000 1.040000 8.070000 1.185000 ;
        RECT 7.360000 0.255000 7.550000 0.870000 ;
        RECT 7.360000 1.875000 7.550000 2.735000 ;
        RECT 7.825000 1.185000 8.070000 1.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.320000  1.920000 2.345000 2.090000 ;
      RECT 0.320000  2.090000 0.580000 3.065000 ;
      RECT 0.390000  0.085000 0.695000 1.095000 ;
      RECT 0.750000  2.260000 1.080000 3.245000 ;
      RECT 1.250000  0.085000 1.580000 0.835000 ;
      RECT 1.250000  2.090000 1.440000 3.065000 ;
      RECT 1.610000  2.260000 1.940000 3.245000 ;
      RECT 2.110000  0.085000 2.885000 0.700000 ;
      RECT 2.110000  2.090000 2.345000 2.895000 ;
      RECT 2.110000  2.895000 4.090000 3.065000 ;
      RECT 2.515000  1.705000 5.820000 1.875000 ;
      RECT 2.515000  1.875000 2.730000 2.725000 ;
      RECT 2.900000  2.055000 3.230000 2.895000 ;
      RECT 3.400000  1.875000 3.615000 2.725000 ;
      RECT 3.420000  0.085000 3.750000 0.700000 ;
      RECT 3.785000  2.055000 4.090000 2.895000 ;
      RECT 4.280000  0.085000 4.610000 0.700000 ;
      RECT 4.280000  2.055000 4.610000 2.905000 ;
      RECT 4.280000  2.905000 8.050000 3.075000 ;
      RECT 4.780000  1.875000 4.970000 2.735000 ;
      RECT 5.140000  0.085000 5.470000 0.700000 ;
      RECT 5.140000  2.055000 5.470000 2.905000 ;
      RECT 5.640000  1.875000 5.820000 2.735000 ;
      RECT 6.000000  0.085000 6.330000 0.700000 ;
      RECT 6.000000  2.055000 6.330000 2.905000 ;
      RECT 6.860000  0.085000 7.190000 0.700000 ;
      RECT 6.860000  2.055000 7.190000 2.905000 ;
      RECT 7.720000  0.085000 8.050000 0.835000 ;
      RECT 7.720000  2.055000 8.050000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__nor4_4
END LIBRARY
