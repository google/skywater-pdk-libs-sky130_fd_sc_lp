* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 X a_100_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=2.4885e+12p ps=2.159e+07u
M1001 a_495_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.079e+12p pd=1.842e+07u as=0p ps=0u
M1002 VGND a_100_23# X VNB nshort w=840000u l=150000u
+  ad=1.1508e+12p pd=1.114e+07u as=4.704e+11p ps=4.48e+06u
M1003 a_667_47# A2 a_922_47# VNB nshort w=840000u l=150000u
+  ad=6.804e+11p pd=6.66e+06u as=4.704e+11p ps=4.48e+06u
M1004 VGND a_100_23# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_495_367# A3 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_100_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_100_23# B1 a_495_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1008 VPWR A2 a_495_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1115_47# A4 VGND VNB nshort w=840000u l=150000u
+  ad=6.804e+11p pd=6.66e+06u as=0p ps=0u
M1010 a_495_367# A4 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1115_47# A3 a_922_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A1 a_495_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_100_23# B1 VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1014 VPWR A3 a_495_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_100_23# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_100_23# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_667_47# A1 a_100_23# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_922_47# A2 a_667_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A4 a_1115_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_100_23# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A4 a_495_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B1 a_100_23# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_495_367# B1 a_100_23# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_100_23# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_100_23# A1 a_667_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_922_47# A3 a_1115_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_495_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
