* File: sky130_fd_sc_lp__o21a_1.spice
* Created: Wed Sep  2 10:15:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21a_1.pex.spice"
.subckt sky130_fd_sc_lp__o21a_1  VNB VPB B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_300_51#_M1005_d N_B1_M1005_g N_A_80_21#_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_300_51#_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1596 AS=0.1176 PD=1.22 PS=1.12 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1006 N_A_300_51#_M1006_d N_A1_M1006_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1596 PD=2.21 PS=1.22 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_80_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4221 AS=0.3339 PD=1.93 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_A_80_21#_M1007_d N_B1_M1007_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.4221 PD=1.65 PS=1.93 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75001
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1001 A_420_367# N_A2_M1001_g N_A_80_21#_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.2457 PD=1.47 PS=1.65 NRD=7.8012 NRS=6.2449 M=1 R=8.4 SA=75001.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_420_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__o21a_1.pxi.spice"
*
.ends
*
*
