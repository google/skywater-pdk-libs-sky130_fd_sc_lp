* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_115_367# C1 a_32_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR A2 a_467_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_684_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_467_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_467_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_32_367# C1 a_115_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_32_367# B1 a_467_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 Y D1 a_115_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_115_367# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VGND A2 a_684_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_684_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_467_367# B1 a_32_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VPWR A1 a_467_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 Y A1 a_684_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
