* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 a_96_49# B2 a_287_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3041e+12p pd=7.11e+06u as=3.024e+11p ps=3e+06u
M1001 a_549_367# A2 a_96_49# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1002 a_179_49# C1 a_96_49# VNB nshort w=840000u l=150000u
+  ad=4.914e+11p pd=4.53e+06u as=2.226e+11p ps=2.21e+06u
M1003 VPWR C1 a_96_49# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0269e+12p pd=6.67e+06u as=0p ps=0u
M1004 a_179_49# B2 a_273_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.48e+06u
M1005 X a_96_49# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=4.914e+11p ps=4.53e+06u
M1006 a_287_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_273_49# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_549_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_96_49# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1010 a_273_49# B1 a_179_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A1 a_273_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
