* File: sky130_fd_sc_lp__o2111ai_0.pex.spice
* Created: Wed Sep  2 10:12:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111AI_0%D1 3 7 9 10 12 13 14 15 20
r38 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=0.93 $X2=0.63 $Y2=0.93
r39 14 15 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=1.665
r40 14 21 13.1451 $w=3.18e-07 $l=3.65e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=0.93
r41 13 21 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=0.705 $Y=0.925
+ $X2=0.705 $Y2=0.93
r42 11 20 51.0643 $w=3.65e-07 $l=3.23e-07 $layer=POLY_cond $X=0.612 $Y=1.253
+ $X2=0.612 $Y2=0.93
r43 11 12 49.3547 $w=3.65e-07 $l=1.82e-07 $layer=POLY_cond $X=0.612 $Y=1.253
+ $X2=0.612 $Y2=1.435
r44 10 20 2.37141 $w=3.65e-07 $l=1.5e-08 $layer=POLY_cond $X=0.612 $Y=0.915
+ $X2=0.612 $Y2=0.93
r45 9 10 44.2957 $w=3.65e-07 $l=1.5e-07 $layer=POLY_cond $X=0.702 $Y=0.765
+ $X2=0.702 $Y2=0.915
r46 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.9 $Y=0.445 $X2=0.9
+ $Y2=0.765
r47 3 12 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=0.505 $Y=2.645
+ $X2=0.505 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_0%C1 3 7 12 16 17 18 19 25
r48 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.665
r49 18 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2 $Y=1.32
+ $X2=1.2 $Y2=1.32
r50 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.925 $X2=1.2
+ $Y2=1.295
r51 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.555 $X2=1.2
+ $Y2=0.925
r52 15 25 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.155
+ $X2=1.2 $Y2=1.32
r53 12 25 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=1.2 $Y=1.645
+ $X2=1.2 $Y2=1.32
r54 9 12 103.008 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=0.935 $Y=1.735
+ $X2=1.2 $Y2=1.735
r55 7 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.26 $Y=0.445
+ $X2=1.26 $Y2=1.155
r56 1 9 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.935 $Y=1.825 $X2=0.935
+ $Y2=1.735
r57 1 3 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.935 $Y=1.825
+ $X2=0.935 $Y2=2.645
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_0%B1 3 5 7 8 9 12 14 15 16 21 23 26
c58 21 0 1.34659e-19 $X=1.77 $Y=0.93
r59 26 28 35.7351 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.27
+ $X2=1.755 $Y2=1.435
r60 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.27 $X2=1.77 $Y2=1.27
r61 22 27 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=1.695 $Y=0.93
+ $X2=1.695 $Y2=1.27
r62 21 24 16.1084 $w=3.9e-07 $l=1.1e-07 $layer=POLY_cond $X=1.74 $Y=0.93
+ $X2=1.74 $Y2=1.04
r63 21 23 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=0.93
+ $X2=1.74 $Y2=0.765
r64 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=0.93 $X2=1.77 $Y2=0.93
r65 15 16 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=1.295
+ $X2=1.695 $Y2=1.665
r66 15 27 0.900346 $w=3.18e-07 $l=2.5e-08 $layer=LI1_cond $X=1.695 $Y=1.295
+ $X2=1.695 $Y2=1.27
r67 14 22 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=1.695 $Y=0.925
+ $X2=1.695 $Y2=0.93
r68 10 12 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.045 $Y=2.185
+ $X2=2.045 $Y2=2.645
r69 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.97 $Y=2.11
+ $X2=2.045 $Y2=2.185
r70 8 9 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.97 $Y=2.11 $X2=1.79
+ $Y2=2.11
r71 7 9 28.0566 $w=1.5e-07 $l=1.40584e-07 $layer=POLY_cond $X=1.682 $Y=2.035
+ $X2=1.79 $Y2=2.11
r72 7 28 179.084 $w=2.15e-07 $l=6e-07 $layer=POLY_cond $X=1.682 $Y=2.035
+ $X2=1.682 $Y2=1.435
r73 5 26 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.755 $Y=1.255
+ $X2=1.755 $Y2=1.27
r74 5 24 34.4622 $w=3.6e-07 $l=2.15e-07 $layer=POLY_cond $X=1.755 $Y=1.255
+ $X2=1.755 $Y2=1.04
r75 3 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.62 $Y=0.445
+ $X2=1.62 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_0%A2 3 6 9 11 12 13 14 15 16 24 42
c55 12 0 1.33668e-19 $X=2.64 $Y=1.295
c56 3 0 4.13819e-20 $X=2.39 $Y=0.445
r57 27 42 2.27456 $w=3.78e-07 $l=7.5e-08 $layer=LI1_cond $X=2.575 $Y=1.59
+ $X2=2.575 $Y2=1.665
r58 24 26 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.32
+ $X2=2.515 $Y2=1.155
r59 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.55
+ $Y=1.32 $X2=2.55 $Y2=1.32
r60 15 16 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=2.405
+ $X2=2.645 $Y2=2.775
r61 14 15 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=2.035
+ $X2=2.645 $Y2=2.405
r62 14 44 12.2447 $w=2.38e-07 $l=2.55e-07 $layer=LI1_cond $X=2.645 $Y=2.035
+ $X2=2.645 $Y2=1.78
r63 13 44 4.89314 $w=3.78e-07 $l=1.1e-07 $layer=LI1_cond $X=2.575 $Y=1.67
+ $X2=2.575 $Y2=1.78
r64 13 42 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=2.575 $Y=1.67
+ $X2=2.575 $Y2=1.665
r65 13 27 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=2.575 $Y=1.585
+ $X2=2.575 $Y2=1.59
r66 13 25 8.03677 $w=3.78e-07 $l=2.65e-07 $layer=LI1_cond $X=2.575 $Y=1.585
+ $X2=2.575 $Y2=1.32
r67 12 25 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.575 $Y=1.295
+ $X2=2.575 $Y2=1.32
r68 9 11 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.525 $Y=2.645
+ $X2=2.525 $Y2=1.825
r69 6 11 39.6483 $w=4e-07 $l=2e-07 $layer=POLY_cond $X=2.515 $Y=1.625 $X2=2.515
+ $Y2=1.825
r70 5 24 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=2.515 $Y=1.355
+ $X2=2.515 $Y2=1.32
r71 5 6 37.5404 $w=4e-07 $l=2.7e-07 $layer=POLY_cond $X=2.515 $Y=1.355 $X2=2.515
+ $Y2=1.625
r72 3 26 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.39 $Y=0.445
+ $X2=2.39 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_0%A1 1 3 6 11 14 15 17 18 19 20 25
c38 11 0 1.33668e-19 $X=3.002 $Y=0.84
r39 19 20 17.2866 $w=2.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.14 $Y=1.63
+ $X2=3.14 $Y2=2.035
r40 19 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.63 $X2=3.09 $Y2=1.63
r41 18 19 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.14 $Y=1.295
+ $X2=3.14 $Y2=1.63
r42 17 25 45.1865 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.465
+ $X2=3.09 $Y2=1.63
r43 14 25 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=3.09 $Y=2.065
+ $X2=3.09 $Y2=1.63
r44 14 15 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.032 $Y=2.065
+ $X2=3.032 $Y2=2.215
r45 9 11 93.3234 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=2.82 $Y=0.84
+ $X2=3.002 $Y2=0.84
r46 7 11 2.19748 $w=1.55e-07 $l=7.5e-08 $layer=POLY_cond $X=3.002 $Y=0.915
+ $X2=3.002 $Y2=0.84
r47 7 17 263.127 $w=1.55e-07 $l=5.5e-07 $layer=POLY_cond $X=3.002 $Y=0.915
+ $X2=3.002 $Y2=1.465
r48 6 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.885 $Y=2.645
+ $X2=2.885 $Y2=2.215
r49 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.82 $Y=0.765 $X2=2.82
+ $Y2=0.84
r50 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.82 $Y=0.765 $X2=2.82
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_0%VPWR 1 2 3 10 12 16 19 21 23 25 30 39 43
r41 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 34 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 31 39 15.2533 $w=1.7e-07 $l=4.35e-07 $layer=LI1_cond $X=1.925 $Y=3.33
+ $X2=1.49 $Y2=3.33
r46 31 33 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.925 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 30 42 4.90987 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.935 $Y=3.33
+ $X2=3.147 $Y2=3.33
r48 30 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 26 36 4.25667 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.202 $Y2=3.33
r52 26 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 25 39 15.2533 $w=1.7e-07 $l=4.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.49 $Y2=3.33
r54 25 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 23 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 23 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 23 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 19 42 2.94129 $w=3.4e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.105 $Y=3.245
+ $X2=3.147 $Y2=3.33
r59 19 21 25.93 $w=3.38e-07 $l=7.65e-07 $layer=LI1_cond $X=3.105 $Y=3.245
+ $X2=3.105 $Y2=2.48
r60 14 39 3.28903 $w=8.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=3.245
+ $X2=1.49 $Y2=3.33
r61 14 16 10.8678 $w=8.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.49 $Y=3.245
+ $X2=1.49 $Y2=2.47
r62 10 36 3.10338 $w=2.8e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.265 $Y=3.245
+ $X2=0.202 $Y2=3.33
r63 10 12 31.898 $w=2.78e-07 $l=7.75e-07 $layer=LI1_cond $X=0.265 $Y=3.245
+ $X2=0.265 $Y2=2.47
r64 3 21 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=2.96
+ $Y=2.325 $X2=3.1 $Y2=2.48
r65 2 16 200 $w=1.7e-07 $l=8.8955e-07 $layer=licon1_PDIFF $count=3 $X=1.01
+ $Y=2.325 $X2=1.83 $Y2=2.47
r66 2 16 200 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=3 $X=1.01
+ $Y=2.325 $X2=1.15 $Y2=2.47
r67 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.325 $X2=0.29 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_0%Y 1 2 3 11 12 14 16 17 20 22 23 24 25 26
+ 27
r58 26 27 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=1.68 $Y2=2.035
r59 26 42 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=0.885 $Y2=2.035
r60 24 25 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=2.405
+ $X2=0.73 $Y2=2.775
r61 23 42 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.73 $Y=2.035
+ $X2=0.885 $Y2=2.035
r62 23 24 8.5987 $w=4.78e-07 $l=2.85e-07 $layer=LI1_cond $X=0.73 $Y=2.12
+ $X2=0.73 $Y2=2.405
r63 22 27 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.095 $Y=2.035
+ $X2=1.68 $Y2=2.035
r64 18 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.225 $Y=2.12
+ $X2=2.095 $Y2=2.035
r65 18 20 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=2.225 $Y=2.12
+ $X2=2.225 $Y2=2.47
r66 16 23 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.575 $Y=2.035
+ $X2=0.73 $Y2=2.035
r67 16 17 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.575 $Y=2.035
+ $X2=0.365 $Y2=2.035
r68 12 14 11.7074 $w=3.13e-07 $l=3.2e-07 $layer=LI1_cond $X=0.365 $Y=0.437
+ $X2=0.685 $Y2=0.437
r69 11 17 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.26 $Y=1.95
+ $X2=0.365 $Y2=2.035
r70 10 12 7.17723 $w=3.15e-07 $l=2.03848e-07 $layer=LI1_cond $X=0.26 $Y=0.595
+ $X2=0.365 $Y2=0.437
r71 10 11 71.5628 $w=2.08e-07 $l=1.355e-06 $layer=LI1_cond $X=0.26 $Y=0.595
+ $X2=0.26 $Y2=1.95
r72 3 20 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.12
+ $Y=2.325 $X2=2.26 $Y2=2.47
r73 2 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.325 $X2=0.72 $Y2=2.47
r74 1 14 91 $w=1.7e-07 $l=5.60245e-07 $layer=licon1_NDIFF $count=2 $X=0.22
+ $Y=0.235 $X2=0.685 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_0%A_339_47# 1 2 7 11 12 13 14 17
c33 17 0 4.13819e-20 $X=3.035 $Y=0.445
c34 12 0 1.34659e-19 $X=2.167 $Y=0.78
r35 15 17 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=3.055 $Y=0.78
+ $X2=3.055 $Y2=0.445
r36 13 15 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.91 $Y=0.865
+ $X2=3.055 $Y2=0.78
r37 13 14 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.91 $Y=0.865
+ $X2=2.3 $Y2=0.865
r38 12 14 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=2.167 $Y=0.78
+ $X2=2.3 $Y2=0.865
r39 11 20 3.74982 $w=2.65e-07 $l=1.58e-07 $layer=LI1_cond $X=2.167 $Y=0.595
+ $X2=2.167 $Y2=0.437
r40 11 12 8.04536 $w=2.63e-07 $l=1.85e-07 $layer=LI1_cond $X=2.167 $Y=0.595
+ $X2=2.167 $Y2=0.78
r41 7 20 3.13276 $w=3.15e-07 $l=1.32e-07 $layer=LI1_cond $X=2.035 $Y=0.437
+ $X2=2.167 $Y2=0.437
r42 7 9 7.3171 $w=3.13e-07 $l=2e-07 $layer=LI1_cond $X=2.035 $Y=0.437 $X2=1.835
+ $Y2=0.437
r43 2 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.035 $Y2=0.445
r44 1 20 182 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.235 $X2=2.175 $Y2=0.445
r45 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.235 $X2=1.835 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_0%VGND 1 6 8 10 20 21 24
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r42 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 18 24 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.605
+ $Y2=0
r44 18 20 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=3.12
+ $Y2=0
r45 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r46 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r47 12 16 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r48 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r49 10 24 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.605
+ $Y2=0
r50 10 16 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.16
+ $Y2=0
r51 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r52 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r53 4 24 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0
r54 4 6 15.3659 $w=2.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0.445
r55 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.605 $Y2=0.445
.ends

