* File: sky130_fd_sc_lp__einvp_lp.pxi.spice
* Created: Fri Aug 28 10:34:14 2020
* 
x_PM_SKY130_FD_SC_LP__EINVP_LP%A N_A_c_40_n N_A_M1006_g N_A_M1005_g A A
+ N_A_c_44_n PM_SKY130_FD_SC_LP__EINVP_LP%A
x_PM_SKY130_FD_SC_LP__EINVP_LP%A_182_321# N_A_182_321#_M1000_d
+ N_A_182_321#_M1003_d N_A_182_321#_M1001_g N_A_182_321#_c_64_n
+ N_A_182_321#_c_71_n N_A_182_321#_c_65_n N_A_182_321#_c_66_n
+ N_A_182_321#_c_67_n N_A_182_321#_c_68_n
+ PM_SKY130_FD_SC_LP__EINVP_LP%A_182_321#
x_PM_SKY130_FD_SC_LP__EINVP_LP%TE N_TE_c_106_n N_TE_M1004_g N_TE_c_107_n
+ N_TE_c_108_n N_TE_M1002_g N_TE_M1003_g N_TE_c_110_n N_TE_M1000_g TE TE TE
+ N_TE_c_112_n N_TE_c_113_n PM_SKY130_FD_SC_LP__EINVP_LP%TE
x_PM_SKY130_FD_SC_LP__EINVP_LP%Z N_Z_M1005_s N_Z_M1006_s Z Z Z Z Z N_Z_c_148_n
+ PM_SKY130_FD_SC_LP__EINVP_LP%Z
x_PM_SKY130_FD_SC_LP__EINVP_LP%VPWR N_VPWR_M1001_d N_VPWR_c_165_n N_VPWR_c_166_n
+ N_VPWR_c_167_n VPWR N_VPWR_c_168_n N_VPWR_c_164_n
+ PM_SKY130_FD_SC_LP__EINVP_LP%VPWR
x_PM_SKY130_FD_SC_LP__EINVP_LP%VGND N_VGND_M1004_d N_VGND_c_187_n VGND
+ N_VGND_c_188_n N_VGND_c_189_n N_VGND_c_190_n N_VGND_c_191_n
+ PM_SKY130_FD_SC_LP__EINVP_LP%VGND
cc_1 VNB N_A_c_40_n 0.0120744f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.36
cc_2 VNB N_A_M1006_g 0.0291831f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_3 VNB N_A_M1005_g 0.0129471f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.915
cc_4 VNB A 0.0361031f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB N_A_c_44_n 0.0440916f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.43
cc_6 VNB N_A_182_321#_c_64_n 0.00415942f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_7 VNB N_A_182_321#_c_65_n 0.0566234f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.467
cc_8 VNB N_A_182_321#_c_66_n 0.00322995f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.467
cc_9 VNB N_A_182_321#_c_67_n 0.00763842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_182_321#_c_68_n 0.00267481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_TE_c_106_n 0.0151217f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.36
cc_12 VNB N_TE_c_107_n 0.00795244f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.595
cc_13 VNB N_TE_c_108_n 0.0157461f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.235
cc_14 VNB N_TE_M1003_g 0.0263287f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_15 VNB N_TE_c_110_n 0.0186459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB TE 0.00632145f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.43
cc_17 VNB N_TE_c_112_n 0.0185817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_TE_c_113_n 0.0436668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Z_c_148_n 0.0344595f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.595
cc_20 VNB N_VPWR_c_164_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_187_n 0.0182396f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.235
cc_22 VNB N_VGND_c_188_n 0.029547f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_23 VNB N_VGND_c_189_n 0.0337222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_190_n 0.17831f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.595
cc_25 VNB N_VGND_c_191_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.467
cc_26 VPB N_A_M1006_g 0.0499793f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_27 VPB N_A_182_321#_M1001_g 0.0280661f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.235
cc_28 VPB N_A_182_321#_c_64_n 0.0102393f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_29 VPB N_A_182_321#_c_71_n 0.0503247f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.43
cc_30 VPB N_A_182_321#_c_66_n 0.0029464f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.467
cc_31 VPB N_A_182_321#_c_67_n 0.023748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_182_321#_c_68_n 0.0054421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_TE_M1003_g 0.0541882f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_34 VPB N_Z_c_148_n 0.0557691f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.595
cc_35 VPB N_VPWR_c_165_n 0.00672007f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.235
cc_36 VPB N_VPWR_c_166_n 0.04412f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_37 VPB N_VPWR_c_167_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_168_n 0.018742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_164_n 0.0461163f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 N_A_M1006_g N_A_182_321#_c_66_n 0.00130581f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_41 N_A_M1006_g N_A_182_321#_c_67_n 0.0933949f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_42 A N_TE_c_106_n 7.41816e-19 $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_43 N_A_c_44_n N_TE_c_106_n 0.0205586f $X=0.505 $Y=0.43 $X2=-0.19 $Y2=-0.245
cc_44 N_A_M1005_g N_TE_c_107_n 0.0205586f $X=0.595 $Y=0.915 $X2=0 $Y2=0
cc_45 N_A_c_40_n N_Z_c_148_n 0.00621331f $X=0.545 $Y=1.36 $X2=0 $Y2=0
cc_46 N_A_M1006_g N_Z_c_148_n 0.0625761f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_47 N_A_M1005_g N_Z_c_148_n 0.00961968f $X=0.595 $Y=0.915 $X2=0 $Y2=0
cc_48 A N_Z_c_148_n 0.0272183f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_49 N_A_c_44_n N_Z_c_148_n 6.99102e-19 $X=0.505 $Y=0.43 $X2=0 $Y2=0
cc_50 N_A_M1006_g N_VPWR_c_166_n 0.00909457f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_51 N_A_M1006_g N_VPWR_c_164_n 0.0163322f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_52 N_A_M1005_g N_VGND_c_187_n 0.00176518f $X=0.595 $Y=0.915 $X2=0 $Y2=0
cc_53 A N_VGND_c_187_n 0.0251515f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_54 N_A_c_44_n N_VGND_c_187_n 0.00182601f $X=0.505 $Y=0.43 $X2=0 $Y2=0
cc_55 A N_VGND_c_188_n 0.0318703f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_56 N_A_c_44_n N_VGND_c_188_n 0.0021213f $X=0.505 $Y=0.43 $X2=0 $Y2=0
cc_57 A N_VGND_c_190_n 0.0251324f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_58 N_A_182_321#_c_66_n N_TE_c_107_n 0.00181553f $X=1.075 $Y=1.69 $X2=0 $Y2=0
cc_59 N_A_182_321#_c_67_n N_TE_c_107_n 0.0168769f $X=1.075 $Y=1.77 $X2=0 $Y2=0
cc_60 N_A_182_321#_M1001_g N_TE_M1003_g 0.0137874f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_61 N_A_182_321#_c_64_n N_TE_M1003_g 0.0235901f $X=1.95 $Y=1.69 $X2=0 $Y2=0
cc_62 N_A_182_321#_c_71_n N_TE_M1003_g 0.0427853f $X=2.115 $Y=2.24 $X2=0 $Y2=0
cc_63 N_A_182_321#_c_66_n N_TE_M1003_g 0.00103266f $X=1.075 $Y=1.69 $X2=0 $Y2=0
cc_64 N_A_182_321#_c_67_n N_TE_M1003_g 0.00795691f $X=1.075 $Y=1.77 $X2=0 $Y2=0
cc_65 N_A_182_321#_c_68_n N_TE_M1003_g 0.00506811f $X=2.115 $Y=1.69 $X2=0 $Y2=0
cc_66 N_A_182_321#_c_65_n N_TE_c_110_n 0.00349251f $X=2.07 $Y=0.715 $X2=0 $Y2=0
cc_67 N_A_182_321#_c_64_n TE 0.0245565f $X=1.95 $Y=1.69 $X2=0 $Y2=0
cc_68 N_A_182_321#_c_65_n TE 0.0507036f $X=2.07 $Y=0.715 $X2=0 $Y2=0
cc_69 N_A_182_321#_c_64_n N_TE_c_112_n 0.00570242f $X=1.95 $Y=1.69 $X2=0 $Y2=0
cc_70 N_A_182_321#_c_64_n N_TE_c_113_n 0.0033339f $X=1.95 $Y=1.69 $X2=0 $Y2=0
cc_71 N_A_182_321#_c_65_n N_TE_c_113_n 0.0205997f $X=2.07 $Y=0.715 $X2=0 $Y2=0
cc_72 N_A_182_321#_c_66_n N_Z_c_148_n 0.0114091f $X=1.075 $Y=1.69 $X2=0 $Y2=0
cc_73 N_A_182_321#_c_67_n N_Z_c_148_n 0.00594806f $X=1.075 $Y=1.77 $X2=0 $Y2=0
cc_74 N_A_182_321#_M1001_g N_VPWR_c_165_n 0.026706f $X=1.035 $Y=2.595 $X2=0
+ $Y2=0
cc_75 N_A_182_321#_c_64_n N_VPWR_c_165_n 0.0184442f $X=1.95 $Y=1.69 $X2=0 $Y2=0
cc_76 N_A_182_321#_c_71_n N_VPWR_c_165_n 0.0652318f $X=2.115 $Y=2.24 $X2=0 $Y2=0
cc_77 N_A_182_321#_M1001_g N_VPWR_c_166_n 0.00975641f $X=1.035 $Y=2.595 $X2=0
+ $Y2=0
cc_78 N_A_182_321#_c_71_n N_VPWR_c_168_n 0.019758f $X=2.115 $Y=2.24 $X2=0 $Y2=0
cc_79 N_A_182_321#_M1003_d N_VPWR_c_164_n 0.0023218f $X=1.975 $Y=2.095 $X2=0
+ $Y2=0
cc_80 N_A_182_321#_M1001_g N_VPWR_c_164_n 0.0177003f $X=1.035 $Y=2.595 $X2=0
+ $Y2=0
cc_81 N_A_182_321#_c_71_n N_VPWR_c_164_n 0.012508f $X=2.115 $Y=2.24 $X2=0 $Y2=0
cc_82 N_A_182_321#_c_64_n N_VGND_c_187_n 0.00185106f $X=1.95 $Y=1.69 $X2=0 $Y2=0
cc_83 N_A_182_321#_c_66_n N_VGND_c_187_n 0.00803444f $X=1.075 $Y=1.69 $X2=0
+ $Y2=0
cc_84 N_A_182_321#_c_67_n N_VGND_c_187_n 4.79785e-19 $X=1.075 $Y=1.77 $X2=0
+ $Y2=0
cc_85 N_A_182_321#_c_65_n N_VGND_c_189_n 0.00843139f $X=2.07 $Y=0.715 $X2=0
+ $Y2=0
cc_86 N_A_182_321#_c_65_n N_VGND_c_190_n 0.00990587f $X=2.07 $Y=0.715 $X2=0
+ $Y2=0
cc_87 N_TE_c_107_n N_Z_c_148_n 5.76476e-19 $X=1.06 $Y=1.275 $X2=0 $Y2=0
cc_88 N_TE_M1003_g N_VPWR_c_165_n 0.0246445f $X=1.85 $Y=2.595 $X2=0 $Y2=0
cc_89 N_TE_M1003_g N_VPWR_c_168_n 0.00840199f $X=1.85 $Y=2.595 $X2=0 $Y2=0
cc_90 N_TE_M1003_g N_VPWR_c_164_n 0.0145288f $X=1.85 $Y=2.595 $X2=0 $Y2=0
cc_91 N_TE_c_106_n N_VGND_c_187_n 0.0122889f $X=0.985 $Y=1.2 $X2=0 $Y2=0
cc_92 N_TE_c_108_n N_VGND_c_187_n 0.00940897f $X=1.495 $Y=1.035 $X2=0 $Y2=0
cc_93 TE N_VGND_c_187_n 0.0513509f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_94 N_TE_c_112_n N_VGND_c_187_n 0.00381987f $X=1.42 $Y=1.2 $X2=0 $Y2=0
cc_95 N_TE_c_106_n N_VGND_c_188_n 0.0031218f $X=0.985 $Y=1.2 $X2=0 $Y2=0
cc_96 N_TE_c_108_n N_VGND_c_189_n 0.00395107f $X=1.495 $Y=1.035 $X2=0 $Y2=0
cc_97 N_TE_c_110_n N_VGND_c_189_n 0.00472472f $X=1.855 $Y=1.035 $X2=0 $Y2=0
cc_98 TE N_VGND_c_189_n 0.0104128f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_99 N_TE_c_106_n N_VGND_c_190_n 0.00376215f $X=0.985 $Y=1.2 $X2=0 $Y2=0
cc_100 N_TE_c_108_n N_VGND_c_190_n 0.00503886f $X=1.495 $Y=1.035 $X2=0 $Y2=0
cc_101 N_TE_c_110_n N_VGND_c_190_n 0.00503886f $X=1.855 $Y=1.035 $X2=0 $Y2=0
cc_102 TE N_VGND_c_190_n 0.011321f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_103 N_Z_c_148_n N_VPWR_c_166_n 0.0210372f $X=0.3 $Y=1.015 $X2=0 $Y2=0
cc_104 N_Z_M1006_s N_VPWR_c_164_n 0.0023218f $X=0.135 $Y=2.095 $X2=0 $Y2=0
cc_105 N_Z_c_148_n N_VPWR_c_164_n 0.0131898f $X=0.3 $Y=1.015 $X2=0 $Y2=0
cc_106 N_Z_c_148_n N_VGND_c_187_n 0.00425379f $X=0.3 $Y=1.015 $X2=0 $Y2=0
cc_107 N_Z_c_148_n N_VGND_c_190_n 9.96765e-19 $X=0.3 $Y=1.015 $X2=0 $Y2=0
cc_108 A_134_419# N_VPWR_c_164_n 0.010279f $X=0.67 $Y=2.095 $X2=2.16 $Y2=3.33
