* File: sky130_fd_sc_lp__mux2_lp.pxi.spice
* Created: Wed Sep  2 10:00:40 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2_LP%A_84_29# N_A_84_29#_M1006_d N_A_84_29#_M1001_d
+ N_A_84_29#_M1009_g N_A_84_29#_c_92_n N_A_84_29#_c_103_n N_A_84_29#_M1000_g
+ N_A_84_29#_c_104_n N_A_84_29#_M1002_g N_A_84_29#_c_105_n N_A_84_29#_M1015_g
+ N_A_84_29#_c_94_n N_A_84_29#_c_95_n N_A_84_29#_c_106_n N_A_84_29#_c_129_p
+ N_A_84_29#_c_96_n N_A_84_29#_c_97_n N_A_84_29#_c_108_n N_A_84_29#_c_109_n
+ N_A_84_29#_c_98_n N_A_84_29#_c_99_n N_A_84_29#_c_110_n N_A_84_29#_c_100_n
+ N_A_84_29#_c_101_n PM_SKY130_FD_SC_LP__MUX2_LP%A_84_29#
x_PM_SKY130_FD_SC_LP__MUX2_LP%A_200_367# N_A_200_367#_M1014_d
+ N_A_200_367#_M1007_d N_A_200_367#_M1010_g N_A_200_367#_M1005_g
+ N_A_200_367#_c_188_n N_A_200_367#_c_193_n N_A_200_367#_c_194_n
+ N_A_200_367#_c_189_n N_A_200_367#_c_196_n N_A_200_367#_c_197_n
+ N_A_200_367#_c_198_n N_A_200_367#_c_190_n N_A_200_367#_c_191_n
+ PM_SKY130_FD_SC_LP__MUX2_LP%A_200_367#
x_PM_SKY130_FD_SC_LP__MUX2_LP%A1 N_A1_M1001_g N_A1_M1003_g N_A1_c_271_n
+ N_A1_c_272_n N_A1_c_273_n N_A1_c_274_n A1 N_A1_c_275_n N_A1_c_276_n
+ PM_SKY130_FD_SC_LP__MUX2_LP%A1
x_PM_SKY130_FD_SC_LP__MUX2_LP%A0 N_A0_c_332_n N_A0_M1006_g N_A0_M1011_g
+ N_A0_c_333_n A0 A0 A0 N_A0_c_335_n N_A0_c_336_n PM_SKY130_FD_SC_LP__MUX2_LP%A0
x_PM_SKY130_FD_SC_LP__MUX2_LP%S N_S_M1012_g N_S_c_391_n N_S_c_392_n N_S_M1008_g
+ N_S_c_394_n N_S_c_395_n N_S_M1004_g N_S_M1013_g N_S_M1007_g N_S_M1014_g
+ N_S_c_398_n N_S_c_387_n N_S_c_399_n S S N_S_c_389_n
+ PM_SKY130_FD_SC_LP__MUX2_LP%S
x_PM_SKY130_FD_SC_LP__MUX2_LP%X N_X_M1009_s N_X_M1000_s N_X_c_454_n X X X X X X
+ PM_SKY130_FD_SC_LP__MUX2_LP%X
x_PM_SKY130_FD_SC_LP__MUX2_LP%VPWR N_VPWR_M1015_d N_VPWR_M1012_d N_VPWR_c_473_n
+ N_VPWR_c_474_n N_VPWR_c_475_n VPWR N_VPWR_c_476_n N_VPWR_c_477_n
+ N_VPWR_c_472_n N_VPWR_c_479_n N_VPWR_c_480_n PM_SKY130_FD_SC_LP__MUX2_LP%VPWR
x_PM_SKY130_FD_SC_LP__MUX2_LP%VGND N_VGND_M1002_d N_VGND_M1008_d N_VGND_c_518_n
+ N_VGND_c_519_n N_VGND_c_520_n VGND N_VGND_c_521_n N_VGND_c_522_n
+ N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n PM_SKY130_FD_SC_LP__MUX2_LP%VGND
cc_1 VNB N_A_84_29#_M1009_g 0.022901f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.485
cc_2 VNB N_A_84_29#_c_92_n 0.00431346f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.375
cc_3 VNB N_A_84_29#_M1002_g 0.0210411f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_4 VNB N_A_84_29#_c_94_n 0.0183441f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.035
cc_5 VNB N_A_84_29#_c_95_n 0.0288136f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.555
cc_6 VNB N_A_84_29#_c_96_n 0.0270585f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.05
cc_7 VNB N_A_84_29#_c_97_n 0.00215769f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.375
cc_8 VNB N_A_84_29#_c_98_n 0.02242f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.94
cc_9 VNB N_A_84_29#_c_99_n 0.00320948f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.94
cc_10 VNB N_A_84_29#_c_100_n 0.0042089f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=0.485
cc_11 VNB N_A_84_29#_c_101_n 0.00281035f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.555
cc_12 VNB N_A_200_367#_M1005_g 0.021879f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.845
cc_13 VNB N_A_200_367#_c_188_n 0.028599f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_14 VNB N_A_200_367#_c_189_n 0.0453343f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.338
cc_15 VNB N_A_200_367#_c_190_n 0.0250713f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.375
cc_16 VNB N_A_200_367#_c_191_n 0.0388181f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.94
cc_17 VNB N_A1_M1001_g 0.00259188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1003_g 0.028228f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.885
cc_19 VNB N_A1_c_271_n 0.0125336f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.485
cc_20 VNB N_A1_c_272_n 0.0045472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_273_n 0.0107057f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.525
cc_22 VNB N_A1_c_274_n 0.0364004f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.845
cc_23 VNB N_A1_c_275_n 0.0344174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_276_n 0.00101293f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=2.525
cc_25 VNB N_A0_c_332_n 0.0175234f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.275
cc_26 VNB N_A0_c_333_n 0.0247521f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.375
cc_27 VNB A0 0.0180519f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.45
cc_28 VNB N_A0_c_335_n 0.0125103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A0_c_336_n 0.0388696f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=2.845
cc_30 VNB N_S_M1008_g 0.0657452f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.485
cc_31 VNB N_S_M1013_g 0.0338687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_S_M1014_g 0.0403933f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.555
cc_33 VNB N_S_c_387_n 0.0161183f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.05
cc_34 VNB S 0.0085604f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=2.46
cc_35 VNB N_S_c_389_n 0.0296656f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=2.845
cc_36 VNB X 0.0223563f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.375
cc_37 VNB X 0.0470948f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.525
cc_38 VNB N_VPWR_c_472_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.45
cc_39 VNB N_VGND_c_518_n 0.00397447f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.485
cc_40 VNB N_VGND_c_519_n 0.0541736f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.555
cc_41 VNB N_VGND_c_520_n 0.0126646f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.845
cc_42 VNB N_VGND_c_521_n 0.0269452f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_43 VNB N_VGND_c_522_n 0.0275816f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.885
cc_44 VNB N_VGND_c_523_n 0.27829f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.035
cc_45 VNB N_VGND_c_524_n 0.0054376f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.45
cc_46 VNB N_VGND_c_525_n 0.0048828f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.05
cc_47 VPB N_A_84_29#_c_92_n 0.042762f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.375
cc_48 VPB N_A_84_29#_c_103_n 0.0187966f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.525
cc_49 VPB N_A_84_29#_c_104_n 0.0238146f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=2.45
cc_50 VPB N_A_84_29#_c_105_n 0.0153956f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=2.525
cc_51 VPB N_A_84_29#_c_106_n 0.00606734f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.45
cc_52 VPB N_A_84_29#_c_97_n 0.0143799f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=2.375
cc_53 VPB N_A_84_29#_c_108_n 0.0135568f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=2.46
cc_54 VPB N_A_84_29#_c_109_n 0.00332868f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=2.46
cc_55 VPB N_A_84_29#_c_110_n 0.00203932f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=2.845
cc_56 VPB N_A_200_367#_M1010_g 0.0345898f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.555
cc_57 VPB N_A_200_367#_c_193_n 0.0494384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_200_367#_c_194_n 0.0374667f $X=-0.19 $Y=1.655 $X2=0.637 $Y2=1.035
cc_59 VPB N_A_200_367#_c_189_n 0.0180671f $X=-0.19 $Y=1.655 $X2=0.637 $Y2=1.338
cc_60 VPB N_A_200_367#_c_196_n 0.00936524f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.45
cc_61 VPB N_A_200_367#_c_197_n 0.0434588f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.025
cc_62 VPB N_A_200_367#_c_198_n 0.013449f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.05
cc_63 VPB N_A_200_367#_c_191_n 0.0114808f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.94
cc_64 VPB N_A1_M1001_g 0.0568091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A1_c_276_n 0.00404993f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=2.525
cc_66 VPB N_A0_M1011_g 0.0539231f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.485
cc_67 VPB A0 0.00771977f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=2.45
cc_68 VPB N_A0_c_335_n 0.0187733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_S_M1012_g 0.0425716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_S_c_391_n 0.0379206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_S_c_392_n 0.0087506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_S_M1008_g 0.00297809f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.485
cc_73 VPB N_S_c_394_n 0.0172047f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.375
cc_74 VPB N_S_c_395_n 0.00834675f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.525
cc_75 VPB N_S_M1004_g 0.0582988f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.45
cc_76 VPB N_S_M1007_g 0.0577266f $X=-0.19 $Y=1.655 $X2=0.637 $Y2=1.035
cc_77 VPB N_S_c_398_n 0.00655551f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.025
cc_78 VPB N_S_c_399_n 0.0128483f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.555
cc_79 VPB S 2.8175e-19 $X=-0.19 $Y=1.655 $X2=1.77 $Y2=2.46
cc_80 VPB N_S_c_389_n 0.00565502f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=2.845
cc_81 VPB N_X_c_454_n 0.025458f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.485
cc_82 VPB X 0.0493904f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.525
cc_83 VPB N_VPWR_c_473_n 0.00151893f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.485
cc_84 VPB N_VPWR_c_474_n 0.0367416f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.555
cc_85 VPB N_VPWR_c_475_n 0.00726902f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.845
cc_86 VPB N_VPWR_c_476_n 0.0279026f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.485
cc_87 VPB N_VPWR_c_477_n 0.0433865f $X=-0.19 $Y=1.655 $X2=0.637 $Y2=1.555
cc_88 VPB N_VPWR_c_472_n 0.0961433f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.45
cc_89 VPB N_VPWR_c_479_n 0.00485788f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.05
cc_90 VPB N_VPWR_c_480_n 0.00541171f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.555
cc_91 N_A_84_29#_c_92_n N_A_200_367#_M1010_g 0.00127901f $X=0.54 $Y=2.375 $X2=0
+ $Y2=0
cc_92 N_A_84_29#_c_104_n N_A_200_367#_M1010_g 0.0214164f $X=0.825 $Y=2.45 $X2=0
+ $Y2=0
cc_93 N_A_84_29#_c_97_n N_A_200_367#_M1010_g 0.00383149f $X=0.745 $Y=2.375 $X2=0
+ $Y2=0
cc_94 N_A_84_29#_c_108_n N_A_200_367#_M1010_g 0.011175f $X=1.77 $Y=2.46 $X2=0
+ $Y2=0
cc_95 N_A_84_29#_c_110_n N_A_200_367#_M1010_g 0.00185872f $X=1.935 $Y=2.845
+ $X2=0 $Y2=0
cc_96 N_A_84_29#_M1002_g N_A_200_367#_M1005_g 0.012931f $X=0.855 $Y=0.485 $X2=0
+ $Y2=0
cc_97 N_A_84_29#_c_98_n N_A_200_367#_M1005_g 0.00439052f $X=1.9 $Y=0.94 $X2=0
+ $Y2=0
cc_98 N_A_84_29#_c_100_n N_A_200_367#_M1005_g 0.00215374f $X=2.065 $Y=0.485
+ $X2=0 $Y2=0
cc_99 N_A_84_29#_M1002_g N_A_200_367#_c_188_n 0.00519362f $X=0.855 $Y=0.485
+ $X2=0 $Y2=0
cc_100 N_A_84_29#_c_98_n N_A_200_367#_c_188_n 0.0268822f $X=1.9 $Y=0.94 $X2=0
+ $Y2=0
cc_101 N_A_84_29#_c_108_n N_A_200_367#_c_193_n 0.0591181f $X=1.77 $Y=2.46 $X2=0
+ $Y2=0
cc_102 N_A_84_29#_c_97_n N_A_200_367#_c_196_n 0.0279729f $X=0.745 $Y=2.375 $X2=0
+ $Y2=0
cc_103 N_A_84_29#_c_108_n N_A_200_367#_c_196_n 0.0257749f $X=1.77 $Y=2.46 $X2=0
+ $Y2=0
cc_104 N_A_84_29#_c_92_n N_A_200_367#_c_197_n 0.00792907f $X=0.54 $Y=2.375 $X2=0
+ $Y2=0
cc_105 N_A_84_29#_c_97_n N_A_200_367#_c_197_n 0.00255116f $X=0.745 $Y=2.375
+ $X2=0 $Y2=0
cc_106 N_A_84_29#_c_108_n N_A_200_367#_c_197_n 0.00159168f $X=1.77 $Y=2.46 $X2=0
+ $Y2=0
cc_107 N_A_84_29#_c_92_n N_A_200_367#_c_191_n 0.00269529f $X=0.54 $Y=2.375 $X2=0
+ $Y2=0
cc_108 N_A_84_29#_c_94_n N_A_200_367#_c_191_n 0.00519362f $X=0.675 $Y=1.035
+ $X2=0 $Y2=0
cc_109 N_A_84_29#_c_129_p N_A_200_367#_c_191_n 0.00248894f $X=0.69 $Y=1.05 $X2=0
+ $Y2=0
cc_110 N_A_84_29#_c_96_n N_A_200_367#_c_191_n 0.0235225f $X=0.69 $Y=1.05 $X2=0
+ $Y2=0
cc_111 N_A_84_29#_c_97_n N_A_200_367#_c_191_n 0.0042122f $X=0.745 $Y=2.375 $X2=0
+ $Y2=0
cc_112 N_A_84_29#_c_108_n N_A1_M1001_g 0.0108481f $X=1.77 $Y=2.46 $X2=0 $Y2=0
cc_113 N_A_84_29#_c_110_n N_A1_M1001_g 0.0107772f $X=1.935 $Y=2.845 $X2=0 $Y2=0
cc_114 N_A_84_29#_c_98_n N_A1_M1003_g 0.00287586f $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_115 N_A_84_29#_c_100_n N_A1_M1003_g 0.0147316f $X=2.065 $Y=0.485 $X2=0 $Y2=0
cc_116 N_A_84_29#_c_98_n N_A1_c_271_n 0.0318229f $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_117 N_A_84_29#_c_129_p N_A1_c_272_n 0.00473167f $X=0.69 $Y=1.05 $X2=0 $Y2=0
cc_118 N_A_84_29#_c_98_n N_A1_c_272_n 0.0273939f $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_119 N_A_84_29#_c_98_n N_A1_c_273_n 0.00505999f $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_120 N_A_84_29#_c_98_n N_A1_c_274_n 3.67954e-19 $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_121 N_A_84_29#_c_98_n N_A1_c_275_n 0.00157992f $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_122 N_A_84_29#_c_129_p N_A1_c_276_n 0.00465591f $X=0.69 $Y=1.05 $X2=0 $Y2=0
cc_123 N_A_84_29#_c_97_n N_A1_c_276_n 0.00659313f $X=0.745 $Y=2.375 $X2=0 $Y2=0
cc_124 N_A_84_29#_c_100_n N_A0_c_332_n 0.0128985f $X=2.065 $Y=0.485 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_84_29#_c_108_n N_A0_M1011_g 0.00560383f $X=1.77 $Y=2.46 $X2=0 $Y2=0
cc_126 N_A_84_29#_c_110_n N_A0_M1011_g 0.010665f $X=1.935 $Y=2.845 $X2=0 $Y2=0
cc_127 N_A_84_29#_c_98_n N_A0_c_333_n 0.0118233f $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_128 N_A_84_29#_c_100_n N_A0_c_333_n 0.00832888f $X=2.065 $Y=0.485 $X2=0 $Y2=0
cc_129 N_A_84_29#_c_98_n N_A0_c_336_n 0.00454694f $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_130 N_A_84_29#_c_108_n N_S_M1012_g 8.3456e-19 $X=1.77 $Y=2.46 $X2=0 $Y2=0
cc_131 N_A_84_29#_c_110_n N_S_M1012_g 0.00164608f $X=1.935 $Y=2.845 $X2=0 $Y2=0
cc_132 N_A_84_29#_c_103_n N_X_c_454_n 0.0103221f $X=0.54 $Y=2.525 $X2=0 $Y2=0
cc_133 N_A_84_29#_c_105_n N_X_c_454_n 0.00147944f $X=0.9 $Y=2.525 $X2=0 $Y2=0
cc_134 N_A_84_29#_M1009_g X 0.0101577f $X=0.495 $Y=0.485 $X2=0 $Y2=0
cc_135 N_A_84_29#_M1002_g X 0.00132086f $X=0.855 $Y=0.485 $X2=0 $Y2=0
cc_136 N_A_84_29#_M1009_g X 0.0245267f $X=0.495 $Y=0.485 $X2=0 $Y2=0
cc_137 N_A_84_29#_c_92_n X 0.027183f $X=0.54 $Y=2.375 $X2=0 $Y2=0
cc_138 N_A_84_29#_c_129_p X 0.04075f $X=0.69 $Y=1.05 $X2=0 $Y2=0
cc_139 N_A_84_29#_c_97_n X 0.042135f $X=0.745 $Y=2.375 $X2=0 $Y2=0
cc_140 N_A_84_29#_c_109_n X 0.00906698f $X=0.83 $Y=2.46 $X2=0 $Y2=0
cc_141 N_A_84_29#_c_99_n X 0.0131023f $X=0.855 $Y=0.94 $X2=0 $Y2=0
cc_142 N_A_84_29#_c_103_n N_VPWR_c_473_n 0.00187407f $X=0.54 $Y=2.525 $X2=0
+ $Y2=0
cc_143 N_A_84_29#_c_105_n N_VPWR_c_473_n 0.0103548f $X=0.9 $Y=2.525 $X2=0 $Y2=0
cc_144 N_A_84_29#_c_108_n N_VPWR_c_473_n 0.0209144f $X=1.77 $Y=2.46 $X2=0 $Y2=0
cc_145 N_A_84_29#_c_110_n N_VPWR_c_473_n 0.011405f $X=1.935 $Y=2.845 $X2=0 $Y2=0
cc_146 N_A_84_29#_c_110_n N_VPWR_c_474_n 0.0233958f $X=1.935 $Y=2.845 $X2=0
+ $Y2=0
cc_147 N_A_84_29#_c_110_n N_VPWR_c_475_n 0.0145731f $X=1.935 $Y=2.845 $X2=0
+ $Y2=0
cc_148 N_A_84_29#_c_103_n N_VPWR_c_476_n 0.00511358f $X=0.54 $Y=2.525 $X2=0
+ $Y2=0
cc_149 N_A_84_29#_c_105_n N_VPWR_c_476_n 0.00452967f $X=0.9 $Y=2.525 $X2=0 $Y2=0
cc_150 N_A_84_29#_c_103_n N_VPWR_c_472_n 0.0102596f $X=0.54 $Y=2.525 $X2=0 $Y2=0
cc_151 N_A_84_29#_c_105_n N_VPWR_c_472_n 0.00414839f $X=0.9 $Y=2.525 $X2=0 $Y2=0
cc_152 N_A_84_29#_c_108_n N_VPWR_c_472_n 0.0205882f $X=1.77 $Y=2.46 $X2=0 $Y2=0
cc_153 N_A_84_29#_c_109_n N_VPWR_c_472_n 0.00697668f $X=0.83 $Y=2.46 $X2=0 $Y2=0
cc_154 N_A_84_29#_c_110_n N_VPWR_c_472_n 0.012542f $X=1.935 $Y=2.845 $X2=0 $Y2=0
cc_155 N_A_84_29#_M1009_g N_VGND_c_518_n 0.0020646f $X=0.495 $Y=0.485 $X2=0
+ $Y2=0
cc_156 N_A_84_29#_M1002_g N_VGND_c_518_n 0.0120518f $X=0.855 $Y=0.485 $X2=0
+ $Y2=0
cc_157 N_A_84_29#_c_98_n N_VGND_c_518_n 0.0238395f $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_158 N_A_84_29#_c_100_n N_VGND_c_518_n 0.0113006f $X=2.065 $Y=0.485 $X2=0
+ $Y2=0
cc_159 N_A_84_29#_c_100_n N_VGND_c_519_n 0.0234289f $X=2.065 $Y=0.485 $X2=0
+ $Y2=0
cc_160 N_A_84_29#_M1009_g N_VGND_c_521_n 0.00511358f $X=0.495 $Y=0.485 $X2=0
+ $Y2=0
cc_161 N_A_84_29#_M1002_g N_VGND_c_521_n 0.00452967f $X=0.855 $Y=0.485 $X2=0
+ $Y2=0
cc_162 N_A_84_29#_M1009_g N_VGND_c_523_n 0.0102307f $X=0.495 $Y=0.485 $X2=0
+ $Y2=0
cc_163 N_A_84_29#_M1002_g N_VGND_c_523_n 0.00429401f $X=0.855 $Y=0.485 $X2=0
+ $Y2=0
cc_164 N_A_84_29#_c_98_n N_VGND_c_523_n 0.0231253f $X=1.9 $Y=0.94 $X2=0 $Y2=0
cc_165 N_A_84_29#_c_99_n N_VGND_c_523_n 0.00604236f $X=0.855 $Y=0.94 $X2=0 $Y2=0
cc_166 N_A_84_29#_c_100_n N_VGND_c_523_n 0.0126421f $X=2.065 $Y=0.485 $X2=0
+ $Y2=0
cc_167 N_A_200_367#_c_193_n N_A1_M1001_g 0.0106402f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_168 N_A_200_367#_c_196_n N_A1_M1001_g 0.00118836f $X=1.165 $Y=2 $X2=0 $Y2=0
cc_169 N_A_200_367#_c_197_n N_A1_M1001_g 0.0729722f $X=1.165 $Y=2 $X2=0 $Y2=0
cc_170 N_A_200_367#_c_191_n N_A1_M1001_g 0.00767658f $X=1.202 $Y=1.835 $X2=0
+ $Y2=0
cc_171 N_A_200_367#_c_193_n N_A1_c_271_n 0.00605229f $X=3.845 $Y=2.12 $X2=0
+ $Y2=0
cc_172 N_A_200_367#_c_188_n N_A1_c_272_n 2.47634e-19 $X=1.46 $Y=0.95 $X2=0 $Y2=0
cc_173 N_A_200_367#_c_191_n N_A1_c_272_n 0.00216343f $X=1.202 $Y=1.835 $X2=0
+ $Y2=0
cc_174 N_A_200_367#_c_188_n N_A1_c_275_n 0.00195413f $X=1.46 $Y=0.95 $X2=0 $Y2=0
cc_175 N_A_200_367#_c_193_n N_A1_c_275_n 7.93964e-19 $X=3.845 $Y=2.12 $X2=0
+ $Y2=0
cc_176 N_A_200_367#_c_191_n N_A1_c_275_n 0.0201901f $X=1.202 $Y=1.835 $X2=0
+ $Y2=0
cc_177 N_A_200_367#_c_193_n N_A1_c_276_n 0.0193274f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_178 N_A_200_367#_c_191_n N_A1_c_276_n 0.00306172f $X=1.202 $Y=1.835 $X2=0
+ $Y2=0
cc_179 N_A_200_367#_M1005_g N_A0_c_332_n 0.0214178f $X=1.46 $Y=0.485 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A_200_367#_c_193_n N_A0_M1011_g 0.014926f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_181 N_A_200_367#_c_188_n N_A0_c_333_n 0.0214178f $X=1.46 $Y=0.95 $X2=0 $Y2=0
cc_182 N_A_200_367#_c_193_n A0 0.0910012f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_183 N_A_200_367#_c_193_n N_A0_c_335_n 0.0041736f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_184 N_A_200_367#_c_188_n N_A0_c_336_n 0.00132639f $X=1.46 $Y=0.95 $X2=0 $Y2=0
cc_185 N_A_200_367#_c_193_n N_S_c_391_n 0.0220819f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_186 N_A_200_367#_c_193_n N_S_c_392_n 0.0108594f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_187 N_A_200_367#_c_193_n N_S_c_394_n 0.00535869f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_188 N_A_200_367#_c_193_n N_S_c_395_n 0.00167556f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_189 N_A_200_367#_c_193_n N_S_M1004_g 0.0157124f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_190 N_A_200_367#_c_194_n N_S_M1004_g 0.00435841f $X=4.01 $Y=2.845 $X2=0 $Y2=0
cc_191 N_A_200_367#_c_190_n N_S_M1013_g 0.00125204f $X=4.02 $Y=0.485 $X2=0 $Y2=0
cc_192 N_A_200_367#_c_193_n N_S_M1007_g 0.0140344f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_193 N_A_200_367#_c_194_n N_S_M1007_g 0.025041f $X=4.01 $Y=2.845 $X2=0 $Y2=0
cc_194 N_A_200_367#_c_198_n N_S_M1007_g 0.00515835f $X=4.015 $Y=2.12 $X2=0 $Y2=0
cc_195 N_A_200_367#_c_189_n N_S_M1014_g 0.0191086f $X=4.1 $Y=2.035 $X2=0 $Y2=0
cc_196 N_A_200_367#_c_190_n N_S_M1014_g 0.0100964f $X=4.02 $Y=0.485 $X2=0 $Y2=0
cc_197 N_A_200_367#_c_198_n N_S_c_387_n 2.83435e-19 $X=4.015 $Y=2.12 $X2=0 $Y2=0
cc_198 N_A_200_367#_c_193_n N_S_c_399_n 2.08832e-19 $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_199 N_A_200_367#_c_193_n S 0.0257893f $X=3.845 $Y=2.12 $X2=0 $Y2=0
cc_200 N_A_200_367#_c_189_n S 0.0353805f $X=4.1 $Y=2.035 $X2=0 $Y2=0
cc_201 N_A_200_367#_c_189_n N_S_c_389_n 0.0182582f $X=4.1 $Y=2.035 $X2=0 $Y2=0
cc_202 N_A_200_367#_M1010_g N_VPWR_c_473_n 0.0105964f $X=1.33 $Y=2.845 $X2=0
+ $Y2=0
cc_203 N_A_200_367#_M1010_g N_VPWR_c_474_n 0.00452967f $X=1.33 $Y=2.845 $X2=0
+ $Y2=0
cc_204 N_A_200_367#_c_193_n N_VPWR_c_475_n 0.0136459f $X=3.845 $Y=2.12 $X2=0
+ $Y2=0
cc_205 N_A_200_367#_c_194_n N_VPWR_c_477_n 0.0241458f $X=4.01 $Y=2.845 $X2=0
+ $Y2=0
cc_206 N_A_200_367#_M1010_g N_VPWR_c_472_n 0.00424103f $X=1.33 $Y=2.845 $X2=0
+ $Y2=0
cc_207 N_A_200_367#_c_194_n N_VPWR_c_472_n 0.0130308f $X=4.01 $Y=2.845 $X2=0
+ $Y2=0
cc_208 N_A_200_367#_M1005_g N_VGND_c_518_n 0.00816797f $X=1.46 $Y=0.485 $X2=0
+ $Y2=0
cc_209 N_A_200_367#_c_188_n N_VGND_c_518_n 6.96729e-19 $X=1.46 $Y=0.95 $X2=0
+ $Y2=0
cc_210 N_A_200_367#_M1005_g N_VGND_c_519_n 0.00545548f $X=1.46 $Y=0.485 $X2=0
+ $Y2=0
cc_211 N_A_200_367#_c_190_n N_VGND_c_520_n 0.0153904f $X=4.02 $Y=0.485 $X2=0
+ $Y2=0
cc_212 N_A_200_367#_c_190_n N_VGND_c_522_n 0.0231046f $X=4.02 $Y=0.485 $X2=0
+ $Y2=0
cc_213 N_A_200_367#_M1005_g N_VGND_c_523_n 0.00637074f $X=1.46 $Y=0.485 $X2=0
+ $Y2=0
cc_214 N_A_200_367#_c_190_n N_VGND_c_523_n 0.0125807f $X=4.02 $Y=0.485 $X2=0
+ $Y2=0
cc_215 N_A1_M1003_g N_A0_c_332_n 0.00841288f $X=2.505 $Y=0.485 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A1_M1001_g N_A0_M1011_g 0.0444134f $X=1.72 $Y=2.845 $X2=0 $Y2=0
cc_217 N_A1_M1003_g N_A0_c_333_n 0.00798058f $X=2.505 $Y=0.485 $X2=0 $Y2=0
cc_218 N_A1_c_271_n N_A0_c_333_n 0.00124623f $X=2.4 $Y=1.28 $X2=0 $Y2=0
cc_219 N_A1_c_275_n N_A0_c_333_n 0.00220182f $X=1.665 $Y=1.43 $X2=0 $Y2=0
cc_220 N_A1_M1001_g A0 7.58552e-19 $X=1.72 $Y=2.845 $X2=0 $Y2=0
cc_221 N_A1_c_271_n A0 0.0266186f $X=2.4 $Y=1.28 $X2=0 $Y2=0
cc_222 N_A1_c_273_n A0 0.0278385f $X=2.565 $Y=1.13 $X2=0 $Y2=0
cc_223 N_A1_c_274_n A0 0.00200801f $X=2.565 $Y=1.13 $X2=0 $Y2=0
cc_224 N_A1_c_275_n A0 2.05067e-19 $X=1.665 $Y=1.43 $X2=0 $Y2=0
cc_225 N_A1_c_276_n A0 0.0172092f $X=1.665 $Y=1.43 $X2=0 $Y2=0
cc_226 N_A1_M1001_g N_A0_c_335_n 0.0140467f $X=1.72 $Y=2.845 $X2=0 $Y2=0
cc_227 N_A1_c_271_n N_A0_c_335_n 0.0041736f $X=2.4 $Y=1.28 $X2=0 $Y2=0
cc_228 N_A1_c_276_n N_A0_c_335_n 7.37089e-19 $X=1.665 $Y=1.43 $X2=0 $Y2=0
cc_229 N_A1_c_271_n N_A0_c_336_n 0.0111052f $X=2.4 $Y=1.28 $X2=0 $Y2=0
cc_230 N_A1_c_273_n N_A0_c_336_n 0.00157653f $X=2.565 $Y=1.13 $X2=0 $Y2=0
cc_231 N_A1_c_274_n N_A0_c_336_n 0.0211103f $X=2.565 $Y=1.13 $X2=0 $Y2=0
cc_232 N_A1_c_275_n N_A0_c_336_n 0.0211289f $X=1.665 $Y=1.43 $X2=0 $Y2=0
cc_233 N_A1_c_276_n N_A0_c_336_n 0.00113383f $X=1.665 $Y=1.43 $X2=0 $Y2=0
cc_234 N_A1_M1003_g N_S_M1008_g 0.0304651f $X=2.505 $Y=0.485 $X2=0 $Y2=0
cc_235 N_A1_c_273_n N_S_M1008_g 0.00358056f $X=2.565 $Y=1.13 $X2=0 $Y2=0
cc_236 N_A1_c_274_n N_S_M1008_g 0.0209433f $X=2.565 $Y=1.13 $X2=0 $Y2=0
cc_237 N_A1_c_273_n S 0.00461026f $X=2.565 $Y=1.13 $X2=0 $Y2=0
cc_238 N_A1_M1001_g N_VPWR_c_473_n 0.00188096f $X=1.72 $Y=2.845 $X2=0 $Y2=0
cc_239 N_A1_M1001_g N_VPWR_c_474_n 0.00511358f $X=1.72 $Y=2.845 $X2=0 $Y2=0
cc_240 N_A1_M1001_g N_VPWR_c_472_n 0.00574447f $X=1.72 $Y=2.845 $X2=0 $Y2=0
cc_241 N_A1_M1003_g N_VGND_c_519_n 0.00545548f $X=2.505 $Y=0.485 $X2=0 $Y2=0
cc_242 N_A1_M1003_g N_VGND_c_520_n 0.00290307f $X=2.505 $Y=0.485 $X2=0 $Y2=0
cc_243 N_A1_M1003_g N_VGND_c_523_n 0.0110623f $X=2.505 $Y=0.485 $X2=0 $Y2=0
cc_244 N_A0_M1011_g N_S_c_392_n 0.057384f $X=2.15 $Y=2.845 $X2=0 $Y2=0
cc_245 A0 N_S_c_392_n 0.00294036f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_246 A0 N_S_M1008_g 0.0142876f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_247 N_A0_c_335_n N_S_M1008_g 0.00502194f $X=2.205 $Y=1.7 $X2=0 $Y2=0
cc_248 A0 N_S_c_395_n 0.00612069f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_249 A0 N_S_c_398_n 0.00764755f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_250 A0 S 0.0269508f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_251 A0 N_S_c_389_n 0.00143053f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_252 N_A0_M1011_g N_VPWR_c_474_n 0.00511358f $X=2.15 $Y=2.845 $X2=0 $Y2=0
cc_253 N_A0_M1011_g N_VPWR_c_475_n 0.00216401f $X=2.15 $Y=2.845 $X2=0 $Y2=0
cc_254 N_A0_M1011_g N_VPWR_c_472_n 0.00961121f $X=2.15 $Y=2.845 $X2=0 $Y2=0
cc_255 N_A0_c_332_n N_VGND_c_519_n 0.00511358f $X=1.85 $Y=0.805 $X2=0 $Y2=0
cc_256 N_A0_c_332_n N_VGND_c_523_n 0.0062351f $X=1.85 $Y=0.805 $X2=0 $Y2=0
cc_257 N_S_M1012_g N_VPWR_c_474_n 0.00452967f $X=2.54 $Y=2.845 $X2=0 $Y2=0
cc_258 N_S_M1012_g N_VPWR_c_475_n 0.0146202f $X=2.54 $Y=2.845 $X2=0 $Y2=0
cc_259 N_S_c_391_n N_VPWR_c_475_n 0.00562326f $X=2.97 $Y=2.18 $X2=0 $Y2=0
cc_260 N_S_M1004_g N_VPWR_c_475_n 0.0148713f $X=3.435 $Y=2.845 $X2=0 $Y2=0
cc_261 N_S_M1004_g N_VPWR_c_477_n 0.00545548f $X=3.435 $Y=2.845 $X2=0 $Y2=0
cc_262 N_S_M1007_g N_VPWR_c_477_n 0.00511358f $X=3.795 $Y=2.845 $X2=0 $Y2=0
cc_263 N_S_M1012_g N_VPWR_c_472_n 0.00809218f $X=2.54 $Y=2.845 $X2=0 $Y2=0
cc_264 N_S_M1004_g N_VPWR_c_472_n 0.0113884f $X=3.435 $Y=2.845 $X2=0 $Y2=0
cc_265 N_S_M1007_g N_VPWR_c_472_n 0.0102504f $X=3.795 $Y=2.845 $X2=0 $Y2=0
cc_266 N_S_M1008_g N_VGND_c_519_n 0.00452967f $X=3.015 $Y=0.485 $X2=0 $Y2=0
cc_267 N_S_M1008_g N_VGND_c_520_n 0.0151547f $X=3.015 $Y=0.485 $X2=0 $Y2=0
cc_268 N_S_M1013_g N_VGND_c_520_n 0.0135085f $X=3.445 $Y=0.485 $X2=0 $Y2=0
cc_269 N_S_M1014_g N_VGND_c_520_n 0.00214625f $X=3.805 $Y=0.485 $X2=0 $Y2=0
cc_270 N_S_c_387_n N_VGND_c_520_n 3.49337e-19 $X=3.62 $Y=1.345 $X2=0 $Y2=0
cc_271 N_S_M1013_g N_VGND_c_522_n 0.00452967f $X=3.445 $Y=0.485 $X2=0 $Y2=0
cc_272 N_S_M1014_g N_VGND_c_522_n 0.00511358f $X=3.805 $Y=0.485 $X2=0 $Y2=0
cc_273 N_S_M1008_g N_VGND_c_523_n 0.00830881f $X=3.015 $Y=0.485 $X2=0 $Y2=0
cc_274 N_S_M1013_g N_VGND_c_523_n 0.00799963f $X=3.445 $Y=0.485 $X2=0 $Y2=0
cc_275 N_S_M1014_g N_VGND_c_523_n 0.010244f $X=3.805 $Y=0.485 $X2=0 $Y2=0
cc_276 N_X_c_454_n N_VPWR_c_473_n 0.0121636f $X=0.325 $Y=2.845 $X2=0 $Y2=0
cc_277 N_X_c_454_n N_VPWR_c_476_n 0.0263822f $X=0.325 $Y=2.845 $X2=0 $Y2=0
cc_278 N_X_c_454_n N_VPWR_c_472_n 0.0143399f $X=0.325 $Y=2.845 $X2=0 $Y2=0
cc_279 X N_VGND_c_518_n 0.0143867f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_280 X N_VGND_c_521_n 0.0232493f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_281 X N_VGND_c_523_n 0.0126078f $X=0.155 $Y=0.47 $X2=0 $Y2=0
