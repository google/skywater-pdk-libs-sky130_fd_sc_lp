* NGSPICE file created from sky130_fd_sc_lp__dlclkp_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlclkp_lp CLK GATE VGND VNB VPB VPWR GCLK
M1000 VGND a_80_21# a_110_47# VNB nshort w=420000u l=150000u
+  ad=5.061e+11p pd=5.77e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR a_584_21# a_526_419# VPB phighvt w=1e+06u l=250000u
+  ad=1.235e+12p pd=1.047e+07u as=3.2e+11p ps=2.64e+06u
M1002 a_1284_47# a_1147_419# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1003 VPWR a_80_21# a_27_47# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1004 VPWR a_584_21# a_1147_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1005 a_1147_419# a_584_21# a_1104_185# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1006 GCLK a_1147_419# a_1284_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1007 a_254_419# GATE VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1008 a_1147_419# CLK VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_284_47# GATE VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1010 a_352_419# a_80_21# a_284_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1011 VGND a_584_21# a_448_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.856e+11p ps=2.2e+06u
M1012 a_526_419# a_80_21# a_352_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=6.2e+11p ps=3.24e+06u
M1013 a_110_47# a_80_21# a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1014 VGND CLK a_923_185# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.365e+11p ps=1.49e+06u
M1015 a_584_21# a_352_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1016 a_923_185# CLK a_80_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1017 a_1104_185# CLK VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_352_419# a_27_47# a_254_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_700_47# a_352_419# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1020 VPWR CLK a_80_21# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1021 GCLK a_1147_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1022 a_448_47# a_27_47# a_352_419# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_584_21# a_352_419# a_700_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends

