* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__busdrivernovlpsleep_20 A SLEEP TE_B KAPWR VGND VNB VPB VPWR
+ Z
X0 VPWR SLEEP a_228_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VPWR A a_1492_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_407_491# a_280_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_2519_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND a_1486_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 KAPWR a_280_47# a_705_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_896_367# a_27_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_280_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VGND a_280_47# a_1053_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_2345_367# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 Z a_1486_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 VPWR SLEEP a_1172_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 a_1172_451# a_280_47# a_896_367# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 VGND A a_1486_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 VGND a_407_491# a_2063_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_110_47# SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1053_47# a_705_367# a_896_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_2519_47# a_2063_47# a_705_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_2033_373# a_1486_47# a_2063_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X24 a_27_47# SLEEP a_110_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 VGND A a_2519_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_705_367# a_2063_47# a_2519_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_705_367# A a_2345_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_228_491# TE_B a_280_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 a_2345_367# A a_705_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 VGND a_407_491# a_1486_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 Z a_1486_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X36 a_2063_47# a_1486_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VGND a_1486_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X38 a_896_367# a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X39 VGND a_1486_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X40 VGND SLEEP a_280_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X41 a_1486_47# a_407_491# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X42 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X43 a_1492_367# a_896_367# a_1486_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X44 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X45 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X46 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X47 Z a_1486_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X48 VGND a_1486_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X49 Z a_1486_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X50 Z a_1486_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X51 VGND a_1486_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X52 VPWR a_407_491# a_2033_373# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X53 a_280_47# SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X54 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X55 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X56 VGND a_1486_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X57 a_1492_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X58 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X59 Z a_1486_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X60 a_1486_47# a_896_367# a_1492_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X61 VGND TE_B a_280_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X62 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X63 KAPWR a_27_47# a_896_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X64 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X65 VGND a_1486_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X66 a_27_47# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X67 a_705_367# a_280_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X68 VPWR SLEEP a_2345_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X69 a_1486_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X70 Z a_1486_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X71 VPWR a_705_367# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X72 a_407_491# a_280_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X73 Z a_705_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
