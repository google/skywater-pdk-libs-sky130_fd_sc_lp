* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor2_lp A B VGND VNB VPB VPWR X
X0 a_159_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_84_93# B a_590_412# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_114_119# a_84_93# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 X a_84_93# a_159_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 VGND a_84_93# a_114_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_272_119# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 X B a_272_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_610_68# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_590_412# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VGND B a_446_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR B a_159_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_446_68# B a_84_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_84_93# A a_610_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
