* File: sky130_fd_sc_lp__nand3b_4.pxi.spice
* Created: Fri Aug 28 10:49:59 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3B_4%A_N N_A_N_c_109_n N_A_N_M1013_g N_A_N_c_112_n
+ N_A_N_M1016_g A_N A_N N_A_N_c_111_n PM_SKY130_FD_SC_LP__NAND3B_4%A_N
x_PM_SKY130_FD_SC_LP__NAND3B_4%A_35_74# N_A_35_74#_M1013_s N_A_35_74#_M1016_s
+ N_A_35_74#_M1001_g N_A_35_74#_c_145_n N_A_35_74#_M1000_g N_A_35_74#_M1009_g
+ N_A_35_74#_c_147_n N_A_35_74#_M1010_g N_A_35_74#_M1017_g N_A_35_74#_c_149_n
+ N_A_35_74#_M1014_g N_A_35_74#_M1023_g N_A_35_74#_c_151_n N_A_35_74#_M1025_g
+ N_A_35_74#_c_152_n N_A_35_74#_c_153_n N_A_35_74#_c_164_n N_A_35_74#_c_154_n
+ N_A_35_74#_c_155_n N_A_35_74#_c_156_n N_A_35_74#_c_157_n N_A_35_74#_c_158_n
+ N_A_35_74#_c_165_n PM_SKY130_FD_SC_LP__NAND3B_4%A_35_74#
x_PM_SKY130_FD_SC_LP__NAND3B_4%B N_B_c_274_n N_B_M1003_g N_B_M1007_g N_B_c_275_n
+ N_B_M1006_g N_B_M1008_g N_B_c_276_n N_B_M1012_g N_B_M1022_g N_B_c_277_n
+ N_B_M1021_g N_B_M1024_g B B B N_B_c_272_n N_B_c_273_n
+ PM_SKY130_FD_SC_LP__NAND3B_4%B
x_PM_SKY130_FD_SC_LP__NAND3B_4%C N_C_M1005_g N_C_M1002_g N_C_M1011_g N_C_M1004_g
+ N_C_M1018_g N_C_M1015_g N_C_M1020_g N_C_M1019_g C C C C C N_C_c_360_n
+ PM_SKY130_FD_SC_LP__NAND3B_4%C
x_PM_SKY130_FD_SC_LP__NAND3B_4%VPWR N_VPWR_M1016_d N_VPWR_M1009_s N_VPWR_M1023_s
+ N_VPWR_M1006_s N_VPWR_M1021_s N_VPWR_M1011_d N_VPWR_M1020_d N_VPWR_c_432_n
+ N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n
+ N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_442_n
+ N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n VPWR
+ N_VPWR_c_447_n N_VPWR_c_448_n N_VPWR_c_431_n N_VPWR_c_450_n N_VPWR_c_451_n
+ N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_454_n PM_SKY130_FD_SC_LP__NAND3B_4%VPWR
x_PM_SKY130_FD_SC_LP__NAND3B_4%Y N_Y_M1000_s N_Y_M1014_s N_Y_M1001_d N_Y_M1017_d
+ N_Y_M1003_d N_Y_M1012_d N_Y_M1005_s N_Y_M1018_s N_Y_c_549_n N_Y_c_550_n
+ N_Y_c_543_n N_Y_c_544_n N_Y_c_537_n N_Y_c_538_n N_Y_c_654_p N_Y_c_539_n
+ N_Y_c_580_n N_Y_c_545_n N_Y_c_588_n N_Y_c_589_n N_Y_c_592_n N_Y_c_605_n
+ N_Y_c_609_n N_Y_c_638_n N_Y_c_540_n N_Y_c_593_n N_Y_c_611_n Y Y N_Y_c_542_n Y
+ N_Y_c_640_n Y N_Y_c_642_n PM_SKY130_FD_SC_LP__NAND3B_4%Y
x_PM_SKY130_FD_SC_LP__NAND3B_4%VGND N_VGND_M1013_d N_VGND_M1002_s N_VGND_M1004_s
+ N_VGND_M1019_s N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n N_VGND_c_663_n
+ N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n VGND N_VGND_c_667_n
+ N_VGND_c_668_n N_VGND_c_669_n N_VGND_c_670_n N_VGND_c_671_n N_VGND_c_672_n
+ PM_SKY130_FD_SC_LP__NAND3B_4%VGND
x_PM_SKY130_FD_SC_LP__NAND3B_4%A_225_47# N_A_225_47#_M1000_d N_A_225_47#_M1010_d
+ N_A_225_47#_M1025_d N_A_225_47#_M1008_d N_A_225_47#_M1024_d
+ N_A_225_47#_c_758_n N_A_225_47#_c_767_n N_A_225_47#_c_759_n
+ N_A_225_47#_c_769_n N_A_225_47#_c_777_n N_A_225_47#_c_779_n
+ N_A_225_47#_c_771_n N_A_225_47#_c_775_n N_A_225_47#_c_783_n
+ N_A_225_47#_c_760_n PM_SKY130_FD_SC_LP__NAND3B_4%A_225_47#
x_PM_SKY130_FD_SC_LP__NAND3B_4%A_652_47# N_A_652_47#_M1007_s N_A_652_47#_M1022_s
+ N_A_652_47#_M1002_d N_A_652_47#_M1015_d N_A_652_47#_c_884_n
+ N_A_652_47#_c_840_n N_A_652_47#_c_841_n N_A_652_47#_c_889_n
+ N_A_652_47#_c_842_n N_A_652_47#_c_875_n N_A_652_47#_c_843_n
+ N_A_652_47#_c_880_n N_A_652_47#_c_844_n N_A_652_47#_c_845_n
+ PM_SKY130_FD_SC_LP__NAND3B_4%A_652_47#
cc_1 VNB N_A_N_c_109_n 0.023124f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.32
cc_2 VNB A_N 0.00135485f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_N_c_111_n 0.0365062f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.485
cc_4 VNB N_A_35_74#_M1001_g 0.00492033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_35_74#_c_145_n 0.0189677f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.52
cc_6 VNB N_A_35_74#_M1009_g 0.00452622f $X=-0.19 $Y=-0.245 $X2=0.702 $Y2=1.295
cc_7 VNB N_A_35_74#_c_147_n 0.0155844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_35_74#_M1017_g 0.00452622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_35_74#_c_149_n 0.0155672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_35_74#_M1023_g 0.00480072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_35_74#_c_151_n 0.01568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_35_74#_c_152_n 0.021539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_35_74#_c_153_n 0.0296277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_35_74#_c_154_n 0.013223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_35_74#_c_155_n 0.00543828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_35_74#_c_156_n 0.00125045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_35_74#_c_157_n 0.117368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_35_74#_c_158_n 0.00717518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_M1007_g 0.0240073f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=2.465
cc_20 VNB N_B_M1008_g 0.022958f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.485
cc_21 VNB N_B_M1022_g 0.0229704f $X=-0.19 $Y=-0.245 $X2=0.702 $Y2=1.665
cc_22 VNB N_B_M1024_g 0.0313016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_272_n 0.0794857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_273_n 0.00167635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C_M1002_g 0.0304352f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_26 VNB N_C_M1004_g 0.0227713f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.52
cc_27 VNB N_C_M1015_g 0.0227713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C_M1019_g 0.0343863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB C 0.0109037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_c_360_n 0.105041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_431_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_537_n 0.0030395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_538_n 0.00184201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_539_n 0.00158822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_540_n 0.00141162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB Y 0.00247066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_542_n 0.00304042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_660_n 0.00962729f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.52
cc_39 VNB N_VGND_c_661_n 0.00896055f $X=-0.19 $Y=-0.245 $X2=0.702 $Y2=1.485
cc_40 VNB N_VGND_c_662_n 3.15212e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_663_n 0.0112246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_664_n 0.0418664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_665_n 0.095439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_666_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_667_n 0.0179884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_668_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_669_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_670_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_671_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_672_n 0.369691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_225_47#_c_758_n 0.00271925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_225_47#_c_759_n 0.00181967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_225_47#_c_760_n 0.00644154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_652_47#_c_840_n 0.00307528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_652_47#_c_841_n 0.00308858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_652_47#_c_842_n 0.0213675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_652_47#_c_843_n 0.00693226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_652_47#_c_844_n 0.00142396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_652_47#_c_845_n 0.00144499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VPB N_A_N_c_112_n 0.0208574f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=1.72
cc_61 VPB A_N 0.0013541f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_62 VPB N_A_N_c_111_n 0.0134345f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.485
cc_63 VPB N_A_35_74#_M1001_g 0.0202883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_35_74#_M1009_g 0.0183705f $X=-0.19 $Y=1.655 $X2=0.702 $Y2=1.295
cc_65 VPB N_A_35_74#_M1017_g 0.0183705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_35_74#_M1023_g 0.0187971f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_35_74#_c_153_n 0.0146829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_35_74#_c_164_n 0.0463766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_35_74#_c_165_n 0.0171701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_B_c_274_n 0.0155917f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.32
cc_71 VPB N_B_c_275_n 0.0166498f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_72 VPB N_B_c_276_n 0.0166657f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=1.52
cc_73 VPB N_B_c_277_n 0.0175964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_B_c_272_n 0.0328556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_B_c_273_n 0.00929249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_C_M1005_g 0.0200551f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.79
cc_77 VPB N_C_M1011_g 0.0178551f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.52
cc_78 VPB N_C_M1018_g 0.0178551f $X=-0.19 $Y=1.655 $X2=0.702 $Y2=1.485
cc_79 VPB N_C_M1020_g 0.0233606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB C 0.0295264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_C_c_360_n 0.0307989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_432_n 0.00458851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_433_n 3.177e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_434_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_435_n 0.00212565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_436_n 0.0166272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_437_n 0.00445366f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_438_n 0.0176949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_439_n 0.00442504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_440_n 0.0162043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_441_n 3.26211e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_442_n 0.0478602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_443_n 0.0253043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_444_n 0.00525701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_445_n 0.0149762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_446_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_447_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_448_n 0.0183725f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_431_n 0.0658851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_450_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_451_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_452_n 0.00631492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_453_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_454_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_Y_c_543_n 0.00307336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_Y_c_544_n 0.00187063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_Y_c_545_n 0.00547399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB Y 3.76166e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 A_N N_A_35_74#_M1001_g 8.80292e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A_N_c_111_n N_A_35_74#_M1001_g 0.0193955f $X=0.685 $Y=1.485 $X2=0 $Y2=0
cc_111 N_A_N_c_109_n N_A_35_74#_c_152_n 0.00310755f $X=0.515 $Y=1.32 $X2=0 $Y2=0
cc_112 N_A_N_c_109_n N_A_35_74#_c_153_n 0.0138607f $X=0.515 $Y=1.32 $X2=0 $Y2=0
cc_113 N_A_N_c_112_n N_A_35_74#_c_153_n 0.00380806f $X=0.79 $Y=1.72 $X2=0 $Y2=0
cc_114 A_N N_A_35_74#_c_153_n 0.0371719f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A_N_c_112_n N_A_35_74#_c_164_n 0.0112657f $X=0.79 $Y=1.72 $X2=0 $Y2=0
cc_116 N_A_N_c_109_n N_A_35_74#_c_154_n 0.0186535f $X=0.515 $Y=1.32 $X2=0 $Y2=0
cc_117 A_N N_A_35_74#_c_154_n 0.0145315f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_118 N_A_N_c_111_n N_A_35_74#_c_154_n 0.0030827f $X=0.685 $Y=1.485 $X2=0 $Y2=0
cc_119 N_A_N_c_109_n N_A_35_74#_c_155_n 0.00307039f $X=0.515 $Y=1.32 $X2=0 $Y2=0
cc_120 A_N N_A_35_74#_c_155_n 0.0251878f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_121 N_A_N_c_111_n N_A_35_74#_c_155_n 0.00137692f $X=0.685 $Y=1.485 $X2=0
+ $Y2=0
cc_122 N_A_N_c_109_n N_A_35_74#_c_157_n 0.00256705f $X=0.515 $Y=1.32 $X2=0 $Y2=0
cc_123 A_N N_A_35_74#_c_157_n 8.44459e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_124 N_A_N_c_111_n N_A_35_74#_c_157_n 0.0159706f $X=0.685 $Y=1.485 $X2=0 $Y2=0
cc_125 N_A_N_c_112_n N_A_35_74#_c_165_n 0.00392704f $X=0.79 $Y=1.72 $X2=0 $Y2=0
cc_126 A_N N_A_35_74#_c_165_n 0.00968263f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A_N_c_111_n N_A_35_74#_c_165_n 0.00817539f $X=0.685 $Y=1.485 $X2=0
+ $Y2=0
cc_128 N_A_N_c_112_n N_VPWR_c_432_n 0.00372864f $X=0.79 $Y=1.72 $X2=0 $Y2=0
cc_129 N_A_N_c_112_n N_VPWR_c_443_n 0.0054895f $X=0.79 $Y=1.72 $X2=0 $Y2=0
cc_130 N_A_N_c_112_n N_VPWR_c_431_n 0.0110647f $X=0.79 $Y=1.72 $X2=0 $Y2=0
cc_131 A_N N_Y_c_544_n 0.00174642f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A_N_c_111_n N_Y_c_544_n 7.48019e-19 $X=0.685 $Y=1.485 $X2=0 $Y2=0
cc_133 A_N N_VGND_M1013_d 0.00223619f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_134 N_A_N_c_109_n N_VGND_c_660_n 0.0125811f $X=0.515 $Y=1.32 $X2=0 $Y2=0
cc_135 N_A_N_c_109_n N_VGND_c_667_n 0.00383152f $X=0.515 $Y=1.32 $X2=0 $Y2=0
cc_136 N_A_N_c_109_n N_VGND_c_672_n 0.00761264f $X=0.515 $Y=1.32 $X2=0 $Y2=0
cc_137 N_A_N_c_109_n N_A_225_47#_c_759_n 6.32428e-19 $X=0.515 $Y=1.32 $X2=0
+ $Y2=0
cc_138 N_A_35_74#_c_151_n N_B_M1007_g 0.0238063f $X=2.755 $Y=1.185 $X2=0 $Y2=0
cc_139 N_A_35_74#_c_157_n N_B_M1007_g 0.00749659f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_140 N_A_35_74#_M1023_g N_B_c_272_n 0.0492356f $X=2.575 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_35_74#_M1001_g N_VPWR_c_432_n 0.00240299f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_35_74#_c_155_n N_VPWR_c_432_n 0.00968272f $X=1.147 $Y=1.315 $X2=0
+ $Y2=0
cc_143 N_A_35_74#_c_157_n N_VPWR_c_432_n 0.00263451f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_144 N_A_35_74#_M1001_g N_VPWR_c_433_n 8.18924e-19 $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_35_74#_M1009_g N_VPWR_c_433_n 0.0142514f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_35_74#_M1017_g N_VPWR_c_433_n 0.0141286f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_35_74#_M1023_g N_VPWR_c_433_n 7.7769e-19 $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_35_74#_M1017_g N_VPWR_c_434_n 0.00486043f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_35_74#_M1023_g N_VPWR_c_434_n 0.00486043f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_35_74#_M1017_g N_VPWR_c_435_n 5.67328e-19 $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_35_74#_M1023_g N_VPWR_c_435_n 0.00976731f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_35_74#_c_164_n N_VPWR_c_443_n 0.0407605f $X=0.575 $Y=2.91 $X2=0 $Y2=0
cc_153 N_A_35_74#_M1001_g N_VPWR_c_445_n 0.00579312f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_154 N_A_35_74#_M1009_g N_VPWR_c_445_n 0.00486043f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_35_74#_M1016_s N_VPWR_c_431_n 0.00215158f $X=0.45 $Y=1.835 $X2=0
+ $Y2=0
cc_156 N_A_35_74#_M1001_g N_VPWR_c_431_n 0.0105992f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_35_74#_M1009_g N_VPWR_c_431_n 0.00824727f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A_35_74#_M1017_g N_VPWR_c_431_n 0.00824727f $X=2.145 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A_35_74#_M1023_g N_VPWR_c_431_n 0.00448966f $X=2.575 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_35_74#_c_164_n N_VPWR_c_431_n 0.0232603f $X=0.575 $Y=2.91 $X2=0 $Y2=0
cc_161 N_A_35_74#_M1001_g N_Y_c_549_n 0.011559f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_35_74#_c_145_n N_Y_c_550_n 0.00996943f $X=1.465 $Y=1.185 $X2=0 $Y2=0
cc_163 N_A_35_74#_c_154_n N_Y_c_550_n 0.0076384f $X=0.975 $Y=0.955 $X2=0 $Y2=0
cc_164 N_A_35_74#_M1009_g N_Y_c_543_n 0.0165106f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_35_74#_M1017_g N_Y_c_543_n 0.0165106f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A_35_74#_c_156_n N_Y_c_543_n 0.0489234f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_167 N_A_35_74#_c_157_n N_Y_c_543_n 0.00280127f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_168 N_A_35_74#_M1001_g N_Y_c_544_n 0.005961f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_35_74#_c_156_n N_Y_c_544_n 0.0195825f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_170 N_A_35_74#_c_157_n N_Y_c_544_n 0.00287397f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_171 N_A_35_74#_c_147_n N_Y_c_537_n 0.0120255f $X=1.895 $Y=1.185 $X2=0 $Y2=0
cc_172 N_A_35_74#_c_149_n N_Y_c_537_n 0.0119789f $X=2.325 $Y=1.185 $X2=0 $Y2=0
cc_173 N_A_35_74#_c_156_n N_Y_c_537_n 0.0473895f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_174 N_A_35_74#_c_157_n N_Y_c_537_n 0.00307213f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_175 N_A_35_74#_c_145_n N_Y_c_538_n 0.00431797f $X=1.465 $Y=1.185 $X2=0 $Y2=0
cc_176 N_A_35_74#_c_154_n N_Y_c_538_n 0.00510507f $X=0.975 $Y=0.955 $X2=0 $Y2=0
cc_177 N_A_35_74#_c_155_n N_Y_c_538_n 0.0078764f $X=1.147 $Y=1.315 $X2=0 $Y2=0
cc_178 N_A_35_74#_c_156_n N_Y_c_538_n 0.0207503f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_179 N_A_35_74#_c_157_n N_Y_c_538_n 0.00316311f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_180 N_A_35_74#_c_151_n N_Y_c_539_n 0.012084f $X=2.755 $Y=1.185 $X2=0 $Y2=0
cc_181 N_A_35_74#_c_156_n N_Y_c_539_n 0.00804017f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_182 N_A_35_74#_M1023_g N_Y_c_545_n 0.0302388f $X=2.575 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_35_74#_c_156_n N_Y_c_545_n 0.0389395f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_184 N_A_35_74#_c_157_n N_Y_c_545_n 0.00782277f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_185 N_A_35_74#_c_156_n N_Y_c_540_n 0.0152441f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_186 N_A_35_74#_c_157_n N_Y_c_540_n 0.00316311f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_187 N_A_35_74#_M1023_g Y 0.00256176f $X=2.575 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_35_74#_c_156_n Y 0.0138198f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_189 N_A_35_74#_c_157_n Y 0.00177702f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_190 N_A_35_74#_c_151_n N_Y_c_542_n 0.00454866f $X=2.755 $Y=1.185 $X2=0 $Y2=0
cc_191 N_A_35_74#_c_156_n N_Y_c_542_n 0.00300279f $X=2.585 $Y=1.4 $X2=0 $Y2=0
cc_192 N_A_35_74#_c_154_n N_VGND_M1013_d 0.00503415f $X=0.975 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_35_74#_c_145_n N_VGND_c_660_n 0.00296666f $X=1.465 $Y=1.185 $X2=0
+ $Y2=0
cc_194 N_A_35_74#_c_152_n N_VGND_c_660_n 0.0131188f $X=0.3 $Y=0.525 $X2=0 $Y2=0
cc_195 N_A_35_74#_c_154_n N_VGND_c_660_n 0.0220026f $X=0.975 $Y=0.955 $X2=0
+ $Y2=0
cc_196 N_A_35_74#_c_145_n N_VGND_c_665_n 0.00357877f $X=1.465 $Y=1.185 $X2=0
+ $Y2=0
cc_197 N_A_35_74#_c_147_n N_VGND_c_665_n 0.00357842f $X=1.895 $Y=1.185 $X2=0
+ $Y2=0
cc_198 N_A_35_74#_c_149_n N_VGND_c_665_n 0.00357842f $X=2.325 $Y=1.185 $X2=0
+ $Y2=0
cc_199 N_A_35_74#_c_151_n N_VGND_c_665_n 0.00357842f $X=2.755 $Y=1.185 $X2=0
+ $Y2=0
cc_200 N_A_35_74#_c_152_n N_VGND_c_667_n 0.0110678f $X=0.3 $Y=0.525 $X2=0 $Y2=0
cc_201 N_A_35_74#_c_145_n N_VGND_c_672_n 0.0068216f $X=1.465 $Y=1.185 $X2=0
+ $Y2=0
cc_202 N_A_35_74#_c_147_n N_VGND_c_672_n 0.00535118f $X=1.895 $Y=1.185 $X2=0
+ $Y2=0
cc_203 N_A_35_74#_c_149_n N_VGND_c_672_n 0.00535118f $X=2.325 $Y=1.185 $X2=0
+ $Y2=0
cc_204 N_A_35_74#_c_151_n N_VGND_c_672_n 0.00537652f $X=2.755 $Y=1.185 $X2=0
+ $Y2=0
cc_205 N_A_35_74#_c_152_n N_VGND_c_672_n 0.00947127f $X=0.3 $Y=0.525 $X2=0 $Y2=0
cc_206 N_A_35_74#_c_154_n N_A_225_47#_M1000_d 0.00512341f $X=0.975 $Y=0.955
+ $X2=-0.19 $Y2=-0.245
cc_207 N_A_35_74#_c_155_n N_A_225_47#_M1000_d 2.98003e-19 $X=1.147 $Y=1.315
+ $X2=-0.19 $Y2=-0.245
cc_208 N_A_35_74#_c_154_n N_A_225_47#_c_758_n 0.0205161f $X=0.975 $Y=0.955 $X2=0
+ $Y2=0
cc_209 N_A_35_74#_c_156_n N_A_225_47#_c_758_n 4.8513e-19 $X=2.585 $Y=1.4 $X2=0
+ $Y2=0
cc_210 N_A_35_74#_c_157_n N_A_225_47#_c_758_n 0.00139172f $X=2.585 $Y=1.4 $X2=0
+ $Y2=0
cc_211 N_A_35_74#_c_145_n N_A_225_47#_c_767_n 0.0132167f $X=1.465 $Y=1.185 $X2=0
+ $Y2=0
cc_212 N_A_35_74#_c_147_n N_A_225_47#_c_767_n 0.00826862f $X=1.895 $Y=1.185
+ $X2=0 $Y2=0
cc_213 N_A_35_74#_c_149_n N_A_225_47#_c_769_n 0.00826862f $X=2.325 $Y=1.185
+ $X2=0 $Y2=0
cc_214 N_A_35_74#_c_151_n N_A_225_47#_c_769_n 0.00826862f $X=2.755 $Y=1.185
+ $X2=0 $Y2=0
cc_215 N_A_35_74#_c_145_n N_A_225_47#_c_771_n 4.4915e-19 $X=1.465 $Y=1.185 $X2=0
+ $Y2=0
cc_216 N_A_35_74#_c_147_n N_A_225_47#_c_771_n 0.00616828f $X=1.895 $Y=1.185
+ $X2=0 $Y2=0
cc_217 N_A_35_74#_c_149_n N_A_225_47#_c_771_n 0.00598198f $X=2.325 $Y=1.185
+ $X2=0 $Y2=0
cc_218 N_A_35_74#_c_151_n N_A_225_47#_c_771_n 4.94237e-19 $X=2.755 $Y=1.185
+ $X2=0 $Y2=0
cc_219 N_A_35_74#_c_149_n N_A_225_47#_c_775_n 4.35384e-19 $X=2.325 $Y=1.185
+ $X2=0 $Y2=0
cc_220 N_A_35_74#_c_151_n N_A_225_47#_c_775_n 0.00598332f $X=2.755 $Y=1.185
+ $X2=0 $Y2=0
cc_221 N_B_c_277_n N_C_M1005_g 0.0306623f $X=4.405 $Y=1.725 $X2=0 $Y2=0
cc_222 N_B_c_273_n N_C_M1005_g 2.8199e-19 $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_223 N_B_c_272_n C 3.91936e-19 $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_224 N_B_c_273_n C 0.0248373f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_225 N_B_c_272_n N_C_c_360_n 0.0260773f $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_226 N_B_c_273_n N_C_c_360_n 0.00123583f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_227 N_B_c_274_n N_VPWR_c_435_n 0.00233948f $X=3.035 $Y=1.725 $X2=0 $Y2=0
cc_228 N_B_c_274_n N_VPWR_c_436_n 0.00585385f $X=3.035 $Y=1.725 $X2=0 $Y2=0
cc_229 N_B_c_275_n N_VPWR_c_436_n 0.00585385f $X=3.465 $Y=1.725 $X2=0 $Y2=0
cc_230 N_B_c_275_n N_VPWR_c_437_n 0.00293635f $X=3.465 $Y=1.725 $X2=0 $Y2=0
cc_231 N_B_c_276_n N_VPWR_c_437_n 0.00294627f $X=3.975 $Y=1.725 $X2=0 $Y2=0
cc_232 N_B_c_276_n N_VPWR_c_438_n 0.00585385f $X=3.975 $Y=1.725 $X2=0 $Y2=0
cc_233 N_B_c_277_n N_VPWR_c_438_n 0.00533769f $X=4.405 $Y=1.725 $X2=0 $Y2=0
cc_234 N_B_c_277_n N_VPWR_c_439_n 0.00712754f $X=4.405 $Y=1.725 $X2=0 $Y2=0
cc_235 N_B_c_274_n N_VPWR_c_431_n 0.00668526f $X=3.035 $Y=1.725 $X2=0 $Y2=0
cc_236 N_B_c_275_n N_VPWR_c_431_n 0.0107161f $X=3.465 $Y=1.725 $X2=0 $Y2=0
cc_237 N_B_c_276_n N_VPWR_c_431_n 0.0107435f $X=3.975 $Y=1.725 $X2=0 $Y2=0
cc_238 N_B_c_277_n N_VPWR_c_431_n 0.00996798f $X=4.405 $Y=1.725 $X2=0 $Y2=0
cc_239 N_B_c_275_n N_Y_c_580_n 0.0134371f $X=3.465 $Y=1.725 $X2=0 $Y2=0
cc_240 N_B_c_276_n N_Y_c_580_n 0.0134371f $X=3.975 $Y=1.725 $X2=0 $Y2=0
cc_241 N_B_c_272_n N_Y_c_580_n 0.00113876f $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_242 N_B_c_273_n N_Y_c_580_n 0.0457817f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_243 N_B_c_274_n N_Y_c_545_n 0.0257509f $X=3.035 $Y=1.725 $X2=0 $Y2=0
cc_244 N_B_c_275_n N_Y_c_545_n 0.00466478f $X=3.465 $Y=1.725 $X2=0 $Y2=0
cc_245 N_B_c_272_n N_Y_c_545_n 0.00633586f $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_246 N_B_c_273_n N_Y_c_545_n 0.00588587f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_247 N_B_c_277_n N_Y_c_588_n 0.0132259f $X=4.405 $Y=1.725 $X2=0 $Y2=0
cc_248 N_B_c_277_n N_Y_c_589_n 0.0112355f $X=4.405 $Y=1.725 $X2=0 $Y2=0
cc_249 N_B_c_272_n N_Y_c_589_n 0.00150636f $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_250 N_B_c_273_n N_Y_c_589_n 0.0261524f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_251 N_B_c_277_n N_Y_c_592_n 7.17653e-19 $X=4.405 $Y=1.725 $X2=0 $Y2=0
cc_252 N_B_c_277_n N_Y_c_593_n 0.00103713f $X=4.405 $Y=1.725 $X2=0 $Y2=0
cc_253 N_B_c_272_n N_Y_c_593_n 7.14461e-19 $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_254 N_B_c_273_n N_Y_c_593_n 0.0220533f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_255 N_B_c_272_n Y 0.0173936f $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_256 N_B_c_273_n Y 0.0213864f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_257 N_B_M1007_g N_Y_c_542_n 0.0101261f $X=3.185 $Y=0.655 $X2=0 $Y2=0
cc_258 N_B_M1008_g N_Y_c_542_n 6.35529e-19 $X=3.615 $Y=0.655 $X2=0 $Y2=0
cc_259 N_B_c_272_n N_Y_c_542_n 4.62069e-19 $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_260 N_B_M1024_g N_VGND_c_661_n 0.00333707f $X=4.475 $Y=0.655 $X2=0 $Y2=0
cc_261 N_B_M1007_g N_VGND_c_665_n 0.00357842f $X=3.185 $Y=0.655 $X2=0 $Y2=0
cc_262 N_B_M1008_g N_VGND_c_665_n 0.00357842f $X=3.615 $Y=0.655 $X2=0 $Y2=0
cc_263 N_B_M1022_g N_VGND_c_665_n 0.00357842f $X=4.045 $Y=0.655 $X2=0 $Y2=0
cc_264 N_B_M1024_g N_VGND_c_665_n 0.00357842f $X=4.475 $Y=0.655 $X2=0 $Y2=0
cc_265 N_B_M1007_g N_VGND_c_672_n 0.00537652f $X=3.185 $Y=0.655 $X2=0 $Y2=0
cc_266 N_B_M1008_g N_VGND_c_672_n 0.00535118f $X=3.615 $Y=0.655 $X2=0 $Y2=0
cc_267 N_B_M1022_g N_VGND_c_672_n 0.00535118f $X=4.045 $Y=0.655 $X2=0 $Y2=0
cc_268 N_B_M1024_g N_VGND_c_672_n 0.00665087f $X=4.475 $Y=0.655 $X2=0 $Y2=0
cc_269 N_B_M1007_g N_A_225_47#_c_777_n 0.0110641f $X=3.185 $Y=0.655 $X2=0 $Y2=0
cc_270 N_B_M1008_g N_A_225_47#_c_777_n 0.00862828f $X=3.615 $Y=0.655 $X2=0 $Y2=0
cc_271 N_B_M1022_g N_A_225_47#_c_779_n 0.00862828f $X=4.045 $Y=0.655 $X2=0 $Y2=0
cc_272 N_B_M1024_g N_A_225_47#_c_779_n 0.0089687f $X=4.475 $Y=0.655 $X2=0 $Y2=0
cc_273 N_B_M1007_g N_A_225_47#_c_775_n 0.00602808f $X=3.185 $Y=0.655 $X2=0 $Y2=0
cc_274 N_B_M1008_g N_A_225_47#_c_775_n 4.88603e-19 $X=3.615 $Y=0.655 $X2=0 $Y2=0
cc_275 N_B_M1007_g N_A_225_47#_c_783_n 4.82945e-19 $X=3.185 $Y=0.655 $X2=0 $Y2=0
cc_276 N_B_M1008_g N_A_225_47#_c_783_n 0.00562277f $X=3.615 $Y=0.655 $X2=0 $Y2=0
cc_277 N_B_M1022_g N_A_225_47#_c_783_n 0.00562277f $X=4.045 $Y=0.655 $X2=0 $Y2=0
cc_278 N_B_M1024_g N_A_225_47#_c_783_n 4.82945e-19 $X=4.475 $Y=0.655 $X2=0 $Y2=0
cc_279 N_B_M1022_g N_A_225_47#_c_760_n 5.14064e-19 $X=4.045 $Y=0.655 $X2=0 $Y2=0
cc_280 N_B_M1024_g N_A_225_47#_c_760_n 0.00724405f $X=4.475 $Y=0.655 $X2=0 $Y2=0
cc_281 N_B_M1008_g N_A_652_47#_c_840_n 0.0149929f $X=3.615 $Y=0.655 $X2=0 $Y2=0
cc_282 N_B_M1022_g N_A_652_47#_c_840_n 0.0156297f $X=4.045 $Y=0.655 $X2=0 $Y2=0
cc_283 N_B_c_272_n N_A_652_47#_c_840_n 0.00275226f $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_284 N_B_c_273_n N_A_652_47#_c_840_n 0.0513425f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_285 N_B_M1007_g N_A_652_47#_c_841_n 0.00150582f $X=3.185 $Y=0.655 $X2=0 $Y2=0
cc_286 N_B_c_272_n N_A_652_47#_c_841_n 0.00344977f $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_287 N_B_c_273_n N_A_652_47#_c_841_n 0.00925359f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_288 N_B_M1024_g N_A_652_47#_c_842_n 0.0142775f $X=4.475 $Y=0.655 $X2=0 $Y2=0
cc_289 N_B_c_272_n N_A_652_47#_c_842_n 0.00458275f $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_290 N_B_c_273_n N_A_652_47#_c_842_n 0.0281202f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_291 N_B_c_272_n N_A_652_47#_c_844_n 0.00280963f $X=4.475 $Y=1.535 $X2=0 $Y2=0
cc_292 N_B_c_273_n N_A_652_47#_c_844_n 0.015984f $X=4.57 $Y=1.51 $X2=0 $Y2=0
cc_293 N_C_M1005_g N_VPWR_c_439_n 0.00933988f $X=5.02 $Y=2.465 $X2=0 $Y2=0
cc_294 N_C_M1005_g N_VPWR_c_440_n 0.00495816f $X=5.02 $Y=2.465 $X2=0 $Y2=0
cc_295 N_C_M1011_g N_VPWR_c_440_n 0.00486043f $X=5.45 $Y=2.465 $X2=0 $Y2=0
cc_296 N_C_M1005_g N_VPWR_c_441_n 7.39816e-19 $X=5.02 $Y=2.465 $X2=0 $Y2=0
cc_297 N_C_M1011_g N_VPWR_c_441_n 0.0150308f $X=5.45 $Y=2.465 $X2=0 $Y2=0
cc_298 N_C_M1018_g N_VPWR_c_441_n 0.014798f $X=5.88 $Y=2.465 $X2=0 $Y2=0
cc_299 N_C_M1020_g N_VPWR_c_441_n 6.77662e-19 $X=6.31 $Y=2.465 $X2=0 $Y2=0
cc_300 N_C_M1018_g N_VPWR_c_442_n 7.26038e-19 $X=5.88 $Y=2.465 $X2=0 $Y2=0
cc_301 N_C_M1020_g N_VPWR_c_442_n 0.0200737f $X=6.31 $Y=2.465 $X2=0 $Y2=0
cc_302 C N_VPWR_c_442_n 0.0258892f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_303 N_C_c_360_n N_VPWR_c_442_n 0.0017771f $X=6.815 $Y=1.51 $X2=0 $Y2=0
cc_304 N_C_M1018_g N_VPWR_c_447_n 0.00486043f $X=5.88 $Y=2.465 $X2=0 $Y2=0
cc_305 N_C_M1020_g N_VPWR_c_447_n 0.00486043f $X=6.31 $Y=2.465 $X2=0 $Y2=0
cc_306 N_C_M1005_g N_VPWR_c_431_n 0.00910981f $X=5.02 $Y=2.465 $X2=0 $Y2=0
cc_307 N_C_M1011_g N_VPWR_c_431_n 0.00824727f $X=5.45 $Y=2.465 $X2=0 $Y2=0
cc_308 N_C_M1018_g N_VPWR_c_431_n 0.00824727f $X=5.88 $Y=2.465 $X2=0 $Y2=0
cc_309 N_C_M1020_g N_VPWR_c_431_n 0.00824727f $X=6.31 $Y=2.465 $X2=0 $Y2=0
cc_310 N_C_M1005_g N_Y_c_588_n 6.84592e-19 $X=5.02 $Y=2.465 $X2=0 $Y2=0
cc_311 N_C_M1005_g N_Y_c_589_n 0.00953547f $X=5.02 $Y=2.465 $X2=0 $Y2=0
cc_312 C N_Y_c_589_n 0.00607203f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_313 N_C_M1005_g N_Y_c_592_n 0.015037f $X=5.02 $Y=2.465 $X2=0 $Y2=0
cc_314 N_C_M1011_g N_Y_c_605_n 0.0122129f $X=5.45 $Y=2.465 $X2=0 $Y2=0
cc_315 N_C_M1018_g N_Y_c_605_n 0.0122595f $X=5.88 $Y=2.465 $X2=0 $Y2=0
cc_316 C N_Y_c_605_n 0.043087f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_317 N_C_c_360_n N_Y_c_605_n 5.62833e-19 $X=6.815 $Y=1.51 $X2=0 $Y2=0
cc_318 C N_Y_c_609_n 0.0154822f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_319 N_C_c_360_n N_Y_c_609_n 6.36061e-19 $X=6.815 $Y=1.51 $X2=0 $Y2=0
cc_320 N_C_M1005_g N_Y_c_611_n 0.00179973f $X=5.02 $Y=2.465 $X2=0 $Y2=0
cc_321 C N_Y_c_611_n 0.0221573f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_322 N_C_c_360_n N_Y_c_611_n 6.37898e-19 $X=6.815 $Y=1.51 $X2=0 $Y2=0
cc_323 N_C_M1002_g N_VGND_c_661_n 0.0123642f $X=5.425 $Y=0.655 $X2=0 $Y2=0
cc_324 N_C_M1004_g N_VGND_c_661_n 6.28154e-19 $X=5.855 $Y=0.655 $X2=0 $Y2=0
cc_325 N_C_M1002_g N_VGND_c_662_n 6.30983e-19 $X=5.425 $Y=0.655 $X2=0 $Y2=0
cc_326 N_C_M1004_g N_VGND_c_662_n 0.0115056f $X=5.855 $Y=0.655 $X2=0 $Y2=0
cc_327 N_C_M1015_g N_VGND_c_662_n 0.0115862f $X=6.285 $Y=0.655 $X2=0 $Y2=0
cc_328 N_C_M1019_g N_VGND_c_662_n 6.45202e-19 $X=6.715 $Y=0.655 $X2=0 $Y2=0
cc_329 N_C_M1019_g N_VGND_c_664_n 0.00707768f $X=6.715 $Y=0.655 $X2=0 $Y2=0
cc_330 C N_VGND_c_664_n 0.0135056f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_331 N_C_c_360_n N_VGND_c_664_n 0.00413353f $X=6.815 $Y=1.51 $X2=0 $Y2=0
cc_332 N_C_M1002_g N_VGND_c_668_n 0.00486043f $X=5.425 $Y=0.655 $X2=0 $Y2=0
cc_333 N_C_M1004_g N_VGND_c_668_n 0.00486043f $X=5.855 $Y=0.655 $X2=0 $Y2=0
cc_334 N_C_M1015_g N_VGND_c_669_n 0.00486043f $X=6.285 $Y=0.655 $X2=0 $Y2=0
cc_335 N_C_M1019_g N_VGND_c_669_n 0.00585385f $X=6.715 $Y=0.655 $X2=0 $Y2=0
cc_336 N_C_M1002_g N_VGND_c_672_n 0.00824727f $X=5.425 $Y=0.655 $X2=0 $Y2=0
cc_337 N_C_M1004_g N_VGND_c_672_n 0.00824727f $X=5.855 $Y=0.655 $X2=0 $Y2=0
cc_338 N_C_M1015_g N_VGND_c_672_n 0.00824727f $X=6.285 $Y=0.655 $X2=0 $Y2=0
cc_339 N_C_M1019_g N_VGND_c_672_n 0.0114643f $X=6.715 $Y=0.655 $X2=0 $Y2=0
cc_340 N_C_M1002_g N_A_225_47#_c_760_n 7.5311e-19 $X=5.425 $Y=0.655 $X2=0 $Y2=0
cc_341 N_C_M1002_g N_A_652_47#_c_842_n 0.0162256f $X=5.425 $Y=0.655 $X2=0 $Y2=0
cc_342 C N_A_652_47#_c_842_n 0.0443683f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_343 N_C_c_360_n N_A_652_47#_c_842_n 0.0111093f $X=6.815 $Y=1.51 $X2=0 $Y2=0
cc_344 N_C_M1004_g N_A_652_47#_c_843_n 0.0141287f $X=5.855 $Y=0.655 $X2=0 $Y2=0
cc_345 N_C_M1015_g N_A_652_47#_c_843_n 0.0138529f $X=6.285 $Y=0.655 $X2=0 $Y2=0
cc_346 N_C_M1019_g N_A_652_47#_c_843_n 0.00485766f $X=6.715 $Y=0.655 $X2=0 $Y2=0
cc_347 C N_A_652_47#_c_843_n 0.0685149f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_348 N_C_c_360_n N_A_652_47#_c_843_n 0.00501697f $X=6.815 $Y=1.51 $X2=0 $Y2=0
cc_349 C N_A_652_47#_c_845_n 0.0161049f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_350 N_C_c_360_n N_A_652_47#_c_845_n 0.00261053f $X=6.815 $Y=1.51 $X2=0 $Y2=0
cc_351 N_VPWR_c_431_n N_Y_M1001_d 0.00380103f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_352 N_VPWR_c_431_n N_Y_M1017_d 0.00536646f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_353 N_VPWR_c_431_n N_Y_M1003_d 0.00380103f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_354 N_VPWR_c_431_n N_Y_M1012_d 0.00223559f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_355 N_VPWR_c_431_n N_Y_M1005_s 0.00380103f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_356 N_VPWR_c_431_n N_Y_M1018_s 0.00536646f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_357 N_VPWR_c_445_n N_Y_c_549_n 0.0143246f $X=1.765 $Y=3.33 $X2=0 $Y2=0
cc_358 N_VPWR_c_431_n N_Y_c_549_n 0.00916141f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_359 N_VPWR_M1009_s N_Y_c_543_n 0.00178679f $X=1.79 $Y=1.835 $X2=0 $Y2=0
cc_360 N_VPWR_c_433_n N_Y_c_543_n 0.0175618f $X=1.93 $Y=2.2 $X2=0 $Y2=0
cc_361 N_VPWR_M1006_s N_Y_c_580_n 0.00484356f $X=3.54 $Y=1.835 $X2=0 $Y2=0
cc_362 N_VPWR_c_437_n N_Y_c_580_n 0.0200142f $X=3.715 $Y=2.38 $X2=0 $Y2=0
cc_363 N_VPWR_M1023_s N_Y_c_545_n 0.00213953f $X=2.65 $Y=1.835 $X2=0 $Y2=0
cc_364 N_VPWR_c_435_n N_Y_c_545_n 0.0191862f $X=2.79 $Y=2.78 $X2=0 $Y2=0
cc_365 N_VPWR_c_431_n N_Y_c_545_n 0.00956897f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_366 N_VPWR_c_438_n N_Y_c_588_n 0.0179664f $X=4.535 $Y=3.33 $X2=0 $Y2=0
cc_367 N_VPWR_c_431_n N_Y_c_588_n 0.01194f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_368 N_VPWR_M1021_s N_Y_c_589_n 0.0128837f $X=4.48 $Y=1.835 $X2=0 $Y2=0
cc_369 N_VPWR_c_439_n N_Y_c_589_n 0.0266042f $X=4.7 $Y=2.375 $X2=0 $Y2=0
cc_370 N_VPWR_c_439_n N_Y_c_592_n 0.0619736f $X=4.7 $Y=2.375 $X2=0 $Y2=0
cc_371 N_VPWR_c_440_n N_Y_c_592_n 0.0180741f $X=5.5 $Y=3.33 $X2=0 $Y2=0
cc_372 N_VPWR_c_431_n N_Y_c_592_n 0.011048f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_373 N_VPWR_M1011_d N_Y_c_605_n 0.00333177f $X=5.525 $Y=1.835 $X2=0 $Y2=0
cc_374 N_VPWR_c_441_n N_Y_c_605_n 0.0170777f $X=5.665 $Y=2.385 $X2=0 $Y2=0
cc_375 N_VPWR_c_447_n N_Y_c_638_n 0.0124525f $X=6.36 $Y=3.33 $X2=0 $Y2=0
cc_376 N_VPWR_c_431_n N_Y_c_638_n 0.00730901f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_377 N_VPWR_c_436_n N_Y_c_640_n 0.0140491f $X=3.55 $Y=3.33 $X2=0 $Y2=0
cc_378 N_VPWR_c_431_n N_Y_c_640_n 0.0090585f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_379 N_VPWR_c_434_n N_Y_c_642_n 0.0124525f $X=2.625 $Y=3.33 $X2=0 $Y2=0
cc_380 N_VPWR_c_431_n N_Y_c_642_n 0.00730901f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_381 N_Y_M1000_s N_VGND_c_672_n 0.00225186f $X=1.54 $Y=0.235 $X2=0 $Y2=0
cc_382 N_Y_M1014_s N_VGND_c_672_n 0.00225186f $X=2.4 $Y=0.235 $X2=0 $Y2=0
cc_383 N_Y_c_537_n N_A_225_47#_M1010_d 0.00176461f $X=2.445 $Y=1.06 $X2=0 $Y2=0
cc_384 N_Y_c_539_n N_A_225_47#_M1025_d 3.40166e-19 $X=2.92 $Y=1.06 $X2=0 $Y2=0
cc_385 N_Y_c_542_n N_A_225_47#_M1025_d 0.00157891f $X=3.062 $Y=1.352 $X2=0 $Y2=0
cc_386 N_Y_M1000_s N_A_225_47#_c_767_n 0.00332344f $X=1.54 $Y=0.235 $X2=0 $Y2=0
cc_387 N_Y_c_550_n N_A_225_47#_c_767_n 0.0140766f $X=1.68 $Y=0.76 $X2=0 $Y2=0
cc_388 N_Y_c_537_n N_A_225_47#_c_767_n 0.00321827f $X=2.445 $Y=1.06 $X2=0 $Y2=0
cc_389 N_Y_M1014_s N_A_225_47#_c_769_n 0.00332344f $X=2.4 $Y=0.235 $X2=0 $Y2=0
cc_390 N_Y_c_537_n N_A_225_47#_c_769_n 0.00321827f $X=2.445 $Y=1.06 $X2=0 $Y2=0
cc_391 N_Y_c_654_p N_A_225_47#_c_769_n 0.0124309f $X=2.54 $Y=0.76 $X2=0 $Y2=0
cc_392 N_Y_c_539_n N_A_225_47#_c_769_n 0.00321827f $X=2.92 $Y=1.06 $X2=0 $Y2=0
cc_393 N_Y_c_537_n N_A_225_47#_c_771_n 0.0167853f $X=2.445 $Y=1.06 $X2=0 $Y2=0
cc_394 N_Y_c_539_n N_A_225_47#_c_775_n 0.00435777f $X=2.92 $Y=1.06 $X2=0 $Y2=0
cc_395 N_Y_c_542_n N_A_225_47#_c_775_n 0.0132851f $X=3.062 $Y=1.352 $X2=0 $Y2=0
cc_396 N_Y_c_542_n N_A_652_47#_c_841_n 0.0108802f $X=3.062 $Y=1.352 $X2=0 $Y2=0
cc_397 N_VGND_c_672_n N_A_225_47#_M1000_d 0.00215965f $X=6.96 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_398 N_VGND_c_672_n N_A_225_47#_M1010_d 0.00223559f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_399 N_VGND_c_672_n N_A_225_47#_M1025_d 0.00223559f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_400 N_VGND_c_672_n N_A_225_47#_M1008_d 0.00223559f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_672_n N_A_225_47#_M1024_d 0.00215158f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_402 N_VGND_c_660_n N_A_225_47#_c_758_n 0.0207632f $X=0.73 $Y=0.585 $X2=0
+ $Y2=0
cc_403 N_VGND_c_665_n N_A_225_47#_c_767_n 0.0330185f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_404 N_VGND_c_672_n N_A_225_47#_c_767_n 0.0212998f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_405 N_VGND_c_660_n N_A_225_47#_c_759_n 0.0139f $X=0.73 $Y=0.585 $X2=0 $Y2=0
cc_406 N_VGND_c_665_n N_A_225_47#_c_759_n 0.0173895f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_407 N_VGND_c_672_n N_A_225_47#_c_759_n 0.0100003f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_c_665_n N_A_225_47#_c_769_n 0.0298674f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_672_n N_A_225_47#_c_769_n 0.0187823f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_665_n N_A_225_47#_c_777_n 0.0300582f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_672_n N_A_225_47#_c_777_n 0.0188286f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_c_665_n N_A_225_47#_c_779_n 0.0300582f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_672_n N_A_225_47#_c_779_n 0.0188286f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_665_n N_A_225_47#_c_771_n 0.0188331f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_672_n N_A_225_47#_c_771_n 0.0123854f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_665_n N_A_225_47#_c_775_n 0.0188331f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_c_672_n N_A_225_47#_c_775_n 0.0123854f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_665_n N_A_225_47#_c_783_n 0.0187942f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_c_672_n N_A_225_47#_c_783_n 0.0123736f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_661_n N_A_225_47#_c_760_n 0.0493778f $X=5.21 $Y=0.38 $X2=0 $Y2=0
cc_421 N_VGND_c_665_n N_A_225_47#_c_760_n 0.021102f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_672_n N_A_225_47#_c_760_n 0.0126219f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_672_n N_A_652_47#_M1007_s 0.00225186f $X=6.96 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_424 N_VGND_c_672_n N_A_652_47#_M1022_s 0.00225186f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_672_n N_A_652_47#_M1002_d 0.00536646f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_672_n N_A_652_47#_M1015_d 0.0041489f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_M1002_s N_A_652_47#_c_842_n 0.00230711f $X=5.085 $Y=0.235 $X2=0
+ $Y2=0
cc_428 N_VGND_c_661_n N_A_652_47#_c_842_n 0.021083f $X=5.21 $Y=0.38 $X2=0 $Y2=0
cc_429 N_VGND_c_668_n N_A_652_47#_c_875_n 0.0124525f $X=5.905 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_672_n N_A_652_47#_c_875_n 0.00730901f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_M1004_s N_A_652_47#_c_843_n 0.00176461f $X=5.93 $Y=0.235 $X2=0
+ $Y2=0
cc_432 N_VGND_c_662_n N_A_652_47#_c_843_n 0.0170777f $X=6.07 $Y=0.36 $X2=0 $Y2=0
cc_433 N_VGND_c_664_n N_A_652_47#_c_843_n 0.00166618f $X=6.93 $Y=0.38 $X2=0
+ $Y2=0
cc_434 N_VGND_c_669_n N_A_652_47#_c_880_n 0.0136943f $X=6.8 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_672_n N_A_652_47#_c_880_n 0.00866972f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_436 N_A_225_47#_c_777_n N_A_652_47#_M1007_s 0.00333487f $X=3.665 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_437 N_A_225_47#_c_779_n N_A_652_47#_M1022_s 0.00333487f $X=4.525 $Y=0.35
+ $X2=0 $Y2=0
cc_438 N_A_225_47#_c_777_n N_A_652_47#_c_884_n 0.0126051f $X=3.665 $Y=0.35 $X2=0
+ $Y2=0
cc_439 N_A_225_47#_M1008_d N_A_652_47#_c_840_n 0.00179194f $X=3.69 $Y=0.235
+ $X2=0 $Y2=0
cc_440 N_A_225_47#_c_777_n N_A_652_47#_c_840_n 0.00359357f $X=3.665 $Y=0.35
+ $X2=0 $Y2=0
cc_441 N_A_225_47#_c_779_n N_A_652_47#_c_840_n 0.00359357f $X=4.525 $Y=0.35
+ $X2=0 $Y2=0
cc_442 N_A_225_47#_c_783_n N_A_652_47#_c_840_n 0.0173351f $X=3.83 $Y=0.36 $X2=0
+ $Y2=0
cc_443 N_A_225_47#_c_779_n N_A_652_47#_c_889_n 0.0127003f $X=4.525 $Y=0.35 $X2=0
+ $Y2=0
cc_444 N_A_225_47#_M1024_d N_A_652_47#_c_842_n 0.00225342f $X=4.55 $Y=0.235
+ $X2=0 $Y2=0
cc_445 N_A_225_47#_c_779_n N_A_652_47#_c_842_n 0.00290962f $X=4.525 $Y=0.35
+ $X2=0 $Y2=0
cc_446 N_A_225_47#_c_760_n N_A_652_47#_c_842_n 0.0218936f $X=4.69 $Y=0.38 $X2=0
+ $Y2=0
