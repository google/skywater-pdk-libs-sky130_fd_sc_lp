* NGSPICE file created from sky130_fd_sc_lp__a211oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 VPWR A2 a_296_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0206e+12p pd=9.18e+06u as=1.0584e+12p ps=9.24e+06u
M1001 a_41_367# B1 a_296_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0206e+12p pd=9.18e+06u as=0p ps=0u
M1002 a_489_65# A1 Y VNB nshort w=840000u l=150000u
+  ad=6.804e+11p pd=6.66e+06u as=7.728e+11p ps=6.88e+06u
M1003 VPWR A1 a_296_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A2 a_489_65# VNB nshort w=840000u l=150000u
+  ad=1.05e+12p pd=9.22e+06u as=0p ps=0u
M1005 a_489_65# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_296_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y C1 a_41_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1009 a_296_367# B1 a_41_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_296_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_41_367# C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_489_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

