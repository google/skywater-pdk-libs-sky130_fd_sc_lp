# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o31a_m
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o31a_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.155000 1.285000 1.825000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.155000 1.765000 2.490000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.015000 2.275000 1.525000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 0.470000 2.735000 1.435000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 0.675000 0.580000 2.235000 ;
        RECT 0.370000 0.345000 0.580000 0.675000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.760000  2.095000 0.970000 3.245000 ;
      RECT 0.800000  0.085000 1.010000 0.545000 ;
      RECT 1.150000  2.670000 2.340000 2.840000 ;
      RECT 1.150000  2.840000 1.480000 3.025000 ;
      RECT 1.230000  0.345000 1.440000 0.665000 ;
      RECT 1.230000  0.665000 2.375000 0.835000 ;
      RECT 1.620000  0.085000 1.950000 0.485000 ;
      RECT 2.130000  1.805000 3.105000 1.975000 ;
      RECT 2.130000  1.975000 2.340000 2.670000 ;
      RECT 2.185000  0.345000 2.375000 0.665000 ;
      RECT 2.610000  2.155000 2.940000 3.245000 ;
      RECT 2.915000  0.345000 3.105000 1.805000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__o31a_m
