* File: sky130_fd_sc_lp__xor2_4.spice
* Created: Fri Aug 28 11:36:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xor2_4.pex.spice"
.subckt sky130_fd_sc_lp__xor2_4  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1012 N_A_110_47#_M1012_d N_A_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75009
+ A=0.126 P=1.98 MULT=1
MM1020 N_A_110_47#_M1012_d N_A_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75008.6 A=0.126 P=1.98 MULT=1
MM1030 N_A_110_47#_M1030_d N_A_M1030_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75008.1 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1007_d N_B_M1007_g N_A_110_47#_M1030_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75007.7 A=0.126 P=1.98 MULT=1
MM1016 N_X_M1007_d N_B_M1016_g N_A_110_47#_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75007.3 A=0.126 P=1.98 MULT=1
MM1019 N_X_M1019_d N_B_M1019_g N_A_110_47#_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75006.8 A=0.126 P=1.98 MULT=1
MM1033 N_X_M1019_d N_B_M1033_g N_A_110_47#_M1033_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75006.4 A=0.126 P=1.98 MULT=1
MM1039 N_A_110_47#_M1033_s N_A_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75003.2
+ SB=75006 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1039_s N_A_776_255#_M1013_g N_X_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.7 SB=75005.5
+ A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1024_d N_A_776_255#_M1024_g N_X_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.1
+ SB=75005.1 A=0.126 P=1.98 MULT=1
MM1026 N_VGND_M1024_d N_A_776_255#_M1026_g N_X_M1026_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.6
+ SB=75004.6 A=0.126 P=1.98 MULT=1
MM1031 N_VGND_M1031_d N_A_776_255#_M1031_g N_X_M1026_s VNB NSHORT L=0.15 W=0.84
+ AD=0.3528 AS=0.1176 PD=1.68 PS=1.12 NRD=26.664 NRS=0 M=1 R=5.6 SA=75005
+ SB=75004.2 A=0.126 P=1.98 MULT=1
MM1008 N_A_776_255#_M1008_d N_A_M1008_g N_VGND_M1031_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3528 PD=1.12 PS=1.68 NRD=0 NRS=53.328 M=1 R=5.6 SA=75006
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1017 N_A_776_255#_M1008_d N_A_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.4
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1018 N_A_776_255#_M1018_d N_A_M1018_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.8
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1034 N_A_776_255#_M1018_d N_A_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75007.3
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1034_s N_B_M1002_g N_A_776_255#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75007.7
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_B_M1015_g N_A_776_255#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75008.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1028 N_VGND_M1015_d N_B_M1028_g N_A_776_255#_M1028_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75008.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1029 N_VGND_M1029_d N_B_M1029_g N_A_776_255#_M1028_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75009 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_27_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2 SB=75005
+ A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1000_d N_A_M1004_g N_A_27_367#_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_A_27_367#_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1014_d N_B_M1003_g N_A_27_367#_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_B_M1009_g N_A_27_367#_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1009_d N_B_M1025_g N_A_27_367#_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1032 N_VPWR_M1032_d N_B_M1032_g N_A_27_367#_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1953 AS=0.1764 PD=1.57 PS=1.54 NRD=2.3443 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1032_d N_A_M1037_g N_A_27_367#_M1037_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1953 AS=0.1827 PD=1.57 PS=1.55 NRD=2.3443 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1005 N_A_27_367#_M1037_s N_A_776_255#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1827 AS=0.1764 PD=1.55 PS=1.54 NRD=1.5563 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_A_27_367#_M1010_d N_A_776_255#_M1010_g N_X_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1022 N_A_27_367#_M1010_d N_A_776_255#_M1022_g N_X_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1035 N_A_27_367#_M1035_d N_A_776_255#_M1035_g N_X_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_1199_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1006_d N_A_M1021_g N_A_1199_367#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1027 N_VPWR_M1027_d N_A_M1027_g N_A_1199_367#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1036 N_VPWR_M1027_d N_A_M1036_g N_A_1199_367#_M1036_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1001 N_A_776_255#_M1001_d N_B_M1001_g N_A_1199_367#_M1036_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_A_776_255#_M1001_d N_B_M1011_g N_A_1199_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1023 N_A_776_255#_M1023_d N_B_M1023_g N_A_1199_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1038 N_A_776_255#_M1023_d N_B_M1038_g N_A_1199_367#_M1038_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.5079 P=24.65
*
.include "sky130_fd_sc_lp__xor2_4.pxi.spice"
*
.ends
*
*
