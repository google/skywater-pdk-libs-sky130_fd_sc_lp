* File: sky130_fd_sc_lp__invlp_m.pxi.spice
* Created: Wed Sep  2 09:57:27 2020
* 
x_PM_SKY130_FD_SC_LP__INVLP_M%A N_A_M1000_g N_A_M1001_g N_A_c_28_n N_A_M1003_g
+ N_A_M1002_g N_A_c_31_n N_A_c_37_n N_A_c_32_n A A A N_A_c_34_n
+ PM_SKY130_FD_SC_LP__INVLP_M%A
x_PM_SKY130_FD_SC_LP__INVLP_M%VPWR N_VPWR_M1001_s N_VPWR_c_63_n N_VPWR_c_64_n
+ VPWR N_VPWR_c_65_n N_VPWR_c_62_n PM_SKY130_FD_SC_LP__INVLP_M%VPWR
x_PM_SKY130_FD_SC_LP__INVLP_M%Y N_Y_M1003_d N_Y_M1002_d Y Y Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__INVLP_M%Y
x_PM_SKY130_FD_SC_LP__INVLP_M%VGND N_VGND_M1000_s N_VGND_c_94_n N_VGND_c_95_n
+ VGND N_VGND_c_96_n N_VGND_c_97_n PM_SKY130_FD_SC_LP__INVLP_M%VGND
cc_1 VNB N_A_M1000_g 0.0350701f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.67
cc_2 VNB N_A_c_28_n 0.00722552f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.255
cc_3 VNB N_A_M1003_g 0.0299316f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.67
cc_4 VNB N_A_M1002_g 0.0171175f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.66
cc_5 VNB N_A_c_31_n 0.0146721f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.255
cc_6 VNB N_A_c_32_n 0.00615289f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.255
cc_7 VNB A 0.029322f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_A_c_34_n 0.024341f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.345
cc_9 VNB N_VPWR_c_62_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.67
cc_10 VNB Y 0.0235589f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.66
cc_11 VNB Y 0.038341f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_12 VNB N_VGND_c_94_n 0.0138117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_95_n 0.0370466f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.66
cc_14 VNB N_VGND_c_96_n 0.0300679f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.67
cc_15 VNB N_VGND_c_97_n 0.128946f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.67
cc_16 VPB N_A_M1001_g 0.0519149f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.66
cc_17 VPB N_A_M1002_g 0.0561364f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.66
cc_18 VPB N_A_c_37_n 0.0175337f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.85
cc_19 VPB A 0.0387193f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_20 VPB N_A_c_34_n 0.00217867f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.345
cc_21 VPB N_VPWR_c_63_n 0.0137858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_64_n 0.0372899f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.66
cc_23 VPB N_VPWR_c_65_n 0.0300679f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.67
cc_24 VPB N_VPWR_c_62_n 0.0647761f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.67
cc_25 VPB Y 0.0235489f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.67
cc_26 VPB Y 0.039355f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_27 N_A_M1001_g N_VPWR_c_64_n 0.0141994f $X=0.545 $Y=2.66 $X2=0 $Y2=0
cc_28 N_A_M1002_g N_VPWR_c_64_n 0.0018473f $X=0.935 $Y=2.66 $X2=0 $Y2=0
cc_29 N_A_c_37_n N_VPWR_c_64_n 7.66517e-19 $X=0.455 $Y=1.85 $X2=0 $Y2=0
cc_30 A N_VPWR_c_64_n 0.0214312f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_31 N_A_M1001_g N_VPWR_c_65_n 0.00426961f $X=0.545 $Y=2.66 $X2=0 $Y2=0
cc_32 N_A_M1002_g N_VPWR_c_65_n 0.00491683f $X=0.935 $Y=2.66 $X2=0 $Y2=0
cc_33 N_A_M1001_g N_VPWR_c_62_n 0.00434697f $X=0.545 $Y=2.66 $X2=0 $Y2=0
cc_34 N_A_M1002_g N_VPWR_c_62_n 0.00517496f $X=0.935 $Y=2.66 $X2=0 $Y2=0
cc_35 N_A_M1000_g Y 0.00130204f $X=0.545 $Y=0.67 $X2=0 $Y2=0
cc_36 N_A_M1003_g Y 0.0105259f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_37 N_A_M1001_g Y 0.00130204f $X=0.545 $Y=2.66 $X2=0 $Y2=0
cc_38 N_A_M1002_g Y 0.0105259f $X=0.935 $Y=2.66 $X2=0 $Y2=0
cc_39 N_A_M1003_g Y 0.0452709f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_40 A Y 0.0630741f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_41 N_A_M1000_g N_VGND_c_95_n 0.0141994f $X=0.545 $Y=0.67 $X2=0 $Y2=0
cc_42 N_A_M1003_g N_VGND_c_95_n 0.0018473f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_43 N_A_c_31_n N_VGND_c_95_n 0.00132932f $X=0.455 $Y=1.255 $X2=0 $Y2=0
cc_44 A N_VGND_c_95_n 0.0205783f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_45 N_A_M1000_g N_VGND_c_96_n 0.00426961f $X=0.545 $Y=0.67 $X2=0 $Y2=0
cc_46 N_A_M1003_g N_VGND_c_96_n 0.00491683f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_47 N_A_M1000_g N_VGND_c_97_n 0.00434697f $X=0.545 $Y=0.67 $X2=0 $Y2=0
cc_48 N_A_M1003_g N_VGND_c_97_n 0.00517496f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_49 N_VPWR_c_64_n Y 0.0145731f $X=0.33 $Y=2.66 $X2=0 $Y2=0
cc_50 N_VPWR_c_65_n Y 0.0105762f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_51 N_VPWR_c_62_n Y 0.011362f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_52 Y N_VGND_c_95_n 0.0145731f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_53 Y N_VGND_c_96_n 0.0105762f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_54 Y N_VGND_c_97_n 0.011362f $X=1.115 $Y=0.47 $X2=0 $Y2=0
