# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__fa_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__fa_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.636000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.220000 1.435000 5.475000 1.505000 ;
        RECT 3.220000 1.505000 4.495000 1.615000 ;
        RECT 4.325000 1.335000 5.475000 1.435000 ;
        RECT 5.305000 1.505000 5.475000 1.845000 ;
        RECT 5.305000 1.845000 6.445000 1.930000 ;
        RECT 5.305000 1.930000 6.935000 2.015000 ;
        RECT 6.115000 1.675000 6.445000 1.845000 ;
        RECT 6.275000 2.015000 6.935000 2.100000 ;
        RECT 6.765000 2.100000 6.935000 2.325000 ;
        RECT 6.765000 2.325000 8.005000 2.495000 ;
        RECT 7.815000 1.415000 8.265000 1.750000 ;
        RECT 7.815000 1.750000 8.005000 2.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.636000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.645000 1.335000 6.695000 1.505000 ;
        RECT 5.645000 1.505000 5.905000 1.665000 ;
        RECT 6.525000 0.525000 9.025000 0.695000 ;
        RECT 6.525000 0.695000 6.695000 1.335000 ;
        RECT 8.500000 0.255000 9.025000 0.525000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.830000 1.570000 2.570000 1.750000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.865000 0.865000 7.295000 1.750000 ;
        RECT 7.115000 1.750000 7.295000 1.815000 ;
        RECT 7.115000 1.815000 7.305000 2.145000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.725000 0.875000 0.905000 ;
        RECT 0.085000 0.905000 0.335000 2.320000 ;
        RECT 0.085000 2.320000 0.805000 2.490000 ;
        RECT 0.545000 0.255000 0.875000 0.725000 ;
        RECT 0.615000 2.490000 0.805000 3.075000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 9.120000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 9.310000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  0.085000 0.375000 0.555000 ;
      RECT 0.115000  2.660000 0.445000 3.245000 ;
      RECT 0.505000  1.075000 1.225000 1.245000 ;
      RECT 0.505000  1.245000 0.685000 1.920000 ;
      RECT 0.505000  1.920000 2.280000 2.150000 ;
      RECT 0.855000  1.425000 1.660000 1.595000 ;
      RECT 0.975000  2.320000 1.350000 3.245000 ;
      RECT 1.045000  0.085000 1.325000 0.710000 ;
      RECT 1.055000  0.880000 2.475000 1.050000 ;
      RECT 1.055000  1.050000 1.225000 1.075000 ;
      RECT 1.490000  1.230000 3.715000 1.255000 ;
      RECT 1.490000  1.255000 3.040000 1.400000 ;
      RECT 1.490000  1.400000 1.660000 1.425000 ;
      RECT 1.520000  2.320000 1.850000 2.820000 ;
      RECT 1.520000  2.820000 2.915000 2.990000 ;
      RECT 1.635000  0.370000 2.995000 0.540000 ;
      RECT 1.635000  0.540000 1.965000 0.710000 ;
      RECT 2.020000  2.150000 2.280000 2.640000 ;
      RECT 2.145000  0.710000 2.475000 0.880000 ;
      RECT 2.585000  2.145000 2.915000 2.820000 ;
      RECT 2.665000  0.540000 2.995000 0.915000 ;
      RECT 2.870000  1.085000 3.715000 1.230000 ;
      RECT 2.870000  1.400000 3.040000 1.785000 ;
      RECT 2.870000  1.785000 3.775000 1.955000 ;
      RECT 3.095000  2.145000 3.425000 3.245000 ;
      RECT 3.165000  0.085000 3.375000 0.915000 ;
      RECT 3.545000  0.640000 4.535000 0.970000 ;
      RECT 3.545000  0.970000 3.715000 1.085000 ;
      RECT 3.605000  1.955000 3.775000 2.075000 ;
      RECT 3.605000  2.075000 4.505000 2.245000 ;
      RECT 4.245000  2.245000 4.505000 2.745000 ;
      RECT 4.675000  1.675000 5.125000 2.120000 ;
      RECT 4.705000  0.640000 4.935000 0.995000 ;
      RECT 4.705000  0.995000 6.180000 1.165000 ;
      RECT 4.795000  2.290000 6.070000 2.470000 ;
      RECT 4.795000  2.470000 5.125000 2.890000 ;
      RECT 5.105000  0.085000 5.810000 0.825000 ;
      RECT 5.355000  2.640000 5.685000 3.245000 ;
      RECT 5.810000  2.200000 6.070000 2.290000 ;
      RECT 5.855000  2.470000 6.070000 2.870000 ;
      RECT 5.980000  0.705000 6.180000 0.995000 ;
      RECT 6.240000  2.270000 6.570000 2.665000 ;
      RECT 6.240000  2.665000 6.935000 3.245000 ;
      RECT 6.455000  0.085000 6.785000 0.355000 ;
      RECT 7.465000  1.075000 9.025000 1.245000 ;
      RECT 7.465000  1.245000 7.645000 1.545000 ;
      RECT 7.465000  2.665000 7.795000 3.245000 ;
      RECT 7.475000  0.085000 7.805000 0.355000 ;
      RECT 8.680000  0.865000 9.025000 1.075000 ;
      RECT 8.680000  1.245000 9.025000 2.495000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  1.950000 0.805000 2.120000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  1.950000 5.125000 2.120000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  1.950000 8.965000 2.120000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
    LAYER met1 ;
      RECT 0.575000 1.920000 0.865000 1.965000 ;
      RECT 0.575000 1.965000 9.025000 2.105000 ;
      RECT 0.575000 2.105000 0.865000 2.150000 ;
      RECT 4.895000 1.920000 5.185000 1.965000 ;
      RECT 4.895000 2.105000 5.185000 2.150000 ;
      RECT 8.735000 1.920000 9.025000 1.965000 ;
      RECT 8.735000 2.105000 9.025000 2.150000 ;
  END
END sky130_fd_sc_lp__fa_2
END LIBRARY
