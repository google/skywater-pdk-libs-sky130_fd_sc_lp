* File: sky130_fd_sc_lp__nor4bb_m.pxi.spice
* Created: Fri Aug 28 10:59:28 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4BB_M%D_N N_D_N_M1010_g N_D_N_M1002_g N_D_N_c_82_n
+ N_D_N_c_86_n D_N D_N N_D_N_c_88_n PM_SKY130_FD_SC_LP__NOR4BB_M%D_N
x_PM_SKY130_FD_SC_LP__NOR4BB_M%A_27_507# N_A_27_507#_M1002_s N_A_27_507#_M1010_s
+ N_A_27_507#_M1004_g N_A_27_507#_c_122_n N_A_27_507#_c_123_n
+ N_A_27_507#_M1003_g N_A_27_507#_c_116_n N_A_27_507#_c_117_n
+ N_A_27_507#_c_126_n N_A_27_507#_c_118_n N_A_27_507#_c_127_n
+ N_A_27_507#_c_128_n N_A_27_507#_c_119_n N_A_27_507#_c_129_n
+ N_A_27_507#_c_120_n N_A_27_507#_c_121_n N_A_27_507#_c_130_n
+ PM_SKY130_FD_SC_LP__NOR4BB_M%A_27_507#
x_PM_SKY130_FD_SC_LP__NOR4BB_M%B N_B_M1011_g N_B_M1009_g B B N_B_c_191_n
+ PM_SKY130_FD_SC_LP__NOR4BB_M%B
x_PM_SKY130_FD_SC_LP__NOR4BB_M%A N_A_M1001_g N_A_M1000_g N_A_c_223_n N_A_c_224_n
+ N_A_c_227_n A A N_A_c_225_n PM_SKY130_FD_SC_LP__NOR4BB_M%A
x_PM_SKY130_FD_SC_LP__NOR4BB_M%A_284_99# N_A_284_99#_M1005_d N_A_284_99#_M1007_d
+ N_A_284_99#_M1008_g N_A_284_99#_c_256_n N_A_284_99#_c_257_n
+ N_A_284_99#_M1006_g N_A_284_99#_c_262_n N_A_284_99#_c_263_n
+ N_A_284_99#_c_264_n N_A_284_99#_c_259_n N_A_284_99#_c_260_n
+ N_A_284_99#_c_266_n PM_SKY130_FD_SC_LP__NOR4BB_M%A_284_99#
x_PM_SKY130_FD_SC_LP__NOR4BB_M%C_N N_C_N_c_313_n N_C_N_M1005_g N_C_N_M1007_g
+ N_C_N_c_314_n C_N C_N C_N C_N N_C_N_c_316_n N_C_N_c_317_n
+ PM_SKY130_FD_SC_LP__NOR4BB_M%C_N
x_PM_SKY130_FD_SC_LP__NOR4BB_M%VPWR N_VPWR_M1010_d N_VPWR_M1001_d N_VPWR_c_350_n
+ N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n VPWR N_VPWR_c_354_n
+ N_VPWR_c_355_n N_VPWR_c_349_n N_VPWR_c_357_n PM_SKY130_FD_SC_LP__NOR4BB_M%VPWR
x_PM_SKY130_FD_SC_LP__NOR4BB_M%Y N_Y_M1004_d N_Y_M1011_d N_Y_M1003_s N_Y_c_383_n
+ N_Y_c_384_n N_Y_c_385_n N_Y_c_389_n N_Y_c_403_n N_Y_c_386_n Y N_Y_c_417_n
+ PM_SKY130_FD_SC_LP__NOR4BB_M%Y
x_PM_SKY130_FD_SC_LP__NOR4BB_M%VGND N_VGND_M1002_d N_VGND_M1008_d N_VGND_M1000_d
+ N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n
+ N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n VGND N_VGND_c_449_n
+ N_VGND_c_450_n N_VGND_c_451_n PM_SKY130_FD_SC_LP__NOR4BB_M%VGND
cc_1 VNB N_D_N_M1002_g 0.0449964f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.835
cc_2 VNB N_D_N_c_82_n 0.0214133f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.655
cc_3 VNB D_N 0.0103408f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_4 VNB N_A_27_507#_c_116_n 0.0178786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_27_507#_c_117_n 0.0229271f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.67
cc_6 VNB N_A_27_507#_c_118_n 0.0156262f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=2.035
cc_7 VNB N_A_27_507#_c_119_n 5.99582e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_507#_c_120_n 0.014624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_507#_c_121_n 0.0165244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_M1011_g 0.0364953f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.745
cc_11 VNB B 0.00944539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_c_191_n 0.0468021f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=2.01
cc_13 VNB N_A_c_223_n 0.0168416f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.655
cc_14 VNB N_A_c_224_n 0.0228339f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.505
cc_15 VNB N_A_c_225_n 0.0185374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_284_99#_M1008_g 0.0246985f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.655
cc_17 VNB N_A_284_99#_c_256_n 0.0244672f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.655
cc_18 VNB N_A_284_99#_c_257_n 0.0069866f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=2.01
cc_19 VNB N_A_284_99#_M1006_g 0.0130038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_284_99#_c_259_n 0.0324235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_284_99#_c_260_n 0.0104722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C_N_c_313_n 0.0234675f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.745
cc_23 VNB N_C_N_c_314_n 0.00135696f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.505
cc_24 VNB C_N 0.00267162f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.655
cc_25 VNB N_C_N_c_316_n 0.0210728f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.67
cc_26 VNB N_C_N_c_317_n 0.0227339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_349_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_383_n 6.62247e-19 $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.655
cc_29 VNB N_Y_c_384_n 0.00449412f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=2.175
cc_30 VNB N_Y_c_385_n 0.02186f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB N_Y_c_386_n 0.00123837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB Y 0.00279971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_441_n 0.0282592f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=2.01
cc_34 VNB N_VGND_c_442_n 0.0230073f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_VGND_c_443_n 0.0196472f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.67
cc_36 VNB N_VGND_c_444_n 0.0199916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_445_n 0.0252142f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.67
cc_38 VNB N_VGND_c_446_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=2.035
cc_39 VNB N_VGND_c_447_n 0.0275615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_448_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_449_n 0.0264871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_450_n 0.267456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_451_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_D_N_M1010_g 0.0452234f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.745
cc_45 VPB N_D_N_c_82_n 0.00612468f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.655
cc_46 VPB N_D_N_c_86_n 0.0194899f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.175
cc_47 VPB D_N 0.0216019f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_48 VPB N_D_N_c_88_n 0.030313f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.67
cc_49 VPB N_A_27_507#_c_122_n 0.0224976f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.505
cc_50 VPB N_A_27_507#_c_123_n 0.0167888f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.655
cc_51 VPB N_A_27_507#_M1003_g 0.0241925f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_52 VPB N_A_27_507#_c_117_n 0.00147314f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.67
cc_53 VPB N_A_27_507#_c_126_n 4.08405e-19 $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.665
cc_54 VPB N_A_27_507#_c_127_n 0.0103678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_27_507#_c_128_n 0.00869431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_27_507#_c_129_n 0.0113612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_27_507#_c_130_n 0.0121549f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_B_M1011_g 0.0251188f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.745
cc_59 VPB N_A_M1001_g 0.0203124f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.745
cc_60 VPB N_A_c_227_n 0.0173285f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.655
cc_61 VPB N_A_284_99#_M1006_g 0.0488767f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_284_99#_c_262_n 0.0868791f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_284_99#_c_263_n 0.0150294f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.67
cc_64 VPB N_A_284_99#_c_264_n 0.0126149f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.67
cc_65 VPB N_A_284_99#_c_259_n 0.0393042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_284_99#_c_266_n 0.0459483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_C_N_M1007_g 0.020557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_C_N_c_314_n 0.0204225f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.505
cc_69 VPB C_N 0.00430735f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.655
cc_70 VPB N_VPWR_c_350_n 0.0213814f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.655
cc_71 VPB N_VPWR_c_351_n 0.0275591f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.175
cc_72 VPB N_VPWR_c_352_n 0.0575342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_353_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_354_n 0.0175984f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.67
cc_75 VPB N_VPWR_c_355_n 0.0283247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_349_n 0.108032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_357_n 0.00617139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_Y_c_384_n 0.00262447f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.175
cc_79 VPB N_Y_c_389_n 0.00381568f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.67
cc_80 N_D_N_M1002_g N_A_27_507#_c_116_n 0.0105742f $X=0.595 $Y=0.835 $X2=0 $Y2=0
cc_81 N_D_N_c_82_n N_A_27_507#_c_117_n 0.0161578f $X=0.445 $Y=1.655 $X2=0 $Y2=0
cc_82 D_N N_A_27_507#_c_117_n 2.30985e-19 $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_83 N_D_N_c_88_n N_A_27_507#_c_117_n 0.00576198f $X=0.385 $Y=1.67 $X2=0 $Y2=0
cc_84 N_D_N_M1010_g N_A_27_507#_c_126_n 3.52891e-19 $X=0.475 $Y=2.745 $X2=0
+ $Y2=0
cc_85 N_D_N_M1002_g N_A_27_507#_c_118_n 0.00839396f $X=0.595 $Y=0.835 $X2=0
+ $Y2=0
cc_86 N_D_N_M1010_g N_A_27_507#_c_127_n 0.0165974f $X=0.475 $Y=2.745 $X2=0 $Y2=0
cc_87 N_D_N_c_86_n N_A_27_507#_c_127_n 3.7612e-19 $X=0.385 $Y=2.175 $X2=0 $Y2=0
cc_88 D_N N_A_27_507#_c_127_n 0.00918005f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_89 N_D_N_c_86_n N_A_27_507#_c_128_n 9.38953e-19 $X=0.385 $Y=2.175 $X2=0 $Y2=0
cc_90 D_N N_A_27_507#_c_128_n 0.0160032f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_91 N_D_N_M1002_g N_A_27_507#_c_119_n 0.00969611f $X=0.595 $Y=0.835 $X2=0
+ $Y2=0
cc_92 N_D_N_c_82_n N_A_27_507#_c_119_n 0.00202635f $X=0.445 $Y=1.655 $X2=0 $Y2=0
cc_93 D_N N_A_27_507#_c_119_n 0.0492293f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_94 N_D_N_c_86_n N_A_27_507#_c_129_n 0.00831589f $X=0.385 $Y=2.175 $X2=0 $Y2=0
cc_95 N_D_N_M1002_g N_A_27_507#_c_120_n 0.0182693f $X=0.595 $Y=0.835 $X2=0 $Y2=0
cc_96 N_D_N_c_82_n N_A_27_507#_c_120_n 0.00380652f $X=0.445 $Y=1.655 $X2=0 $Y2=0
cc_97 D_N N_A_27_507#_c_120_n 0.0194347f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_98 N_D_N_M1002_g N_A_27_507#_c_121_n 0.0161578f $X=0.595 $Y=0.835 $X2=0 $Y2=0
cc_99 N_D_N_c_82_n N_A_27_507#_c_130_n 0.00227311f $X=0.445 $Y=1.655 $X2=0 $Y2=0
cc_100 N_D_N_c_88_n N_A_27_507#_c_130_n 0.00831589f $X=0.385 $Y=1.67 $X2=0 $Y2=0
cc_101 N_D_N_M1010_g N_VPWR_c_350_n 0.0153836f $X=0.475 $Y=2.745 $X2=0 $Y2=0
cc_102 N_D_N_M1010_g N_VPWR_c_354_n 0.00379792f $X=0.475 $Y=2.745 $X2=0 $Y2=0
cc_103 N_D_N_M1010_g N_VPWR_c_349_n 0.00457201f $X=0.475 $Y=2.745 $X2=0 $Y2=0
cc_104 N_D_N_M1002_g N_VGND_c_441_n 0.0032771f $X=0.595 $Y=0.835 $X2=0 $Y2=0
cc_105 N_D_N_M1002_g N_VGND_c_445_n 0.00415323f $X=0.595 $Y=0.835 $X2=0 $Y2=0
cc_106 N_D_N_M1002_g N_VGND_c_450_n 0.00469432f $X=0.595 $Y=0.835 $X2=0 $Y2=0
cc_107 N_A_27_507#_c_116_n N_A_284_99#_M1008_g 0.0120484f $X=1.045 $Y=1.155
+ $X2=0 $Y2=0
cc_108 N_A_27_507#_c_121_n N_A_284_99#_M1008_g 0.00863618f $X=1.045 $Y=1.32
+ $X2=0 $Y2=0
cc_109 N_A_27_507#_c_122_n N_A_284_99#_c_257_n 0.00810936f $X=1.4 $Y=1.75 $X2=0
+ $Y2=0
cc_110 N_A_27_507#_c_117_n N_A_284_99#_c_257_n 0.00863618f $X=1.045 $Y=1.675
+ $X2=0 $Y2=0
cc_111 N_A_27_507#_c_122_n N_A_284_99#_M1006_g 0.0550193f $X=1.4 $Y=1.75 $X2=0
+ $Y2=0
cc_112 N_A_27_507#_c_117_n N_A_284_99#_M1006_g 0.00332356f $X=1.045 $Y=1.675
+ $X2=0 $Y2=0
cc_113 N_A_27_507#_c_127_n N_VPWR_c_350_n 0.0214292f $X=0.65 $Y=2.44 $X2=0 $Y2=0
cc_114 N_A_27_507#_c_126_n N_VPWR_c_354_n 0.00508656f $X=0.26 $Y=2.68 $X2=0
+ $Y2=0
cc_115 N_A_27_507#_M1003_g N_VPWR_c_349_n 0.00393927f $X=1.475 $Y=2.195 $X2=0
+ $Y2=0
cc_116 N_A_27_507#_c_126_n N_VPWR_c_349_n 0.00626512f $X=0.26 $Y=2.68 $X2=0
+ $Y2=0
cc_117 N_A_27_507#_c_127_n N_VPWR_c_349_n 0.00661368f $X=0.65 $Y=2.44 $X2=0
+ $Y2=0
cc_118 N_A_27_507#_c_116_n N_Y_c_383_n 0.00264399f $X=1.045 $Y=1.155 $X2=0 $Y2=0
cc_119 N_A_27_507#_c_122_n N_Y_c_384_n 0.0112403f $X=1.4 $Y=1.75 $X2=0 $Y2=0
cc_120 N_A_27_507#_M1003_g N_Y_c_384_n 0.00708909f $X=1.475 $Y=2.195 $X2=0 $Y2=0
cc_121 N_A_27_507#_c_119_n N_Y_c_384_n 0.0364061f $X=0.89 $Y=1.585 $X2=0 $Y2=0
cc_122 N_A_27_507#_c_129_n N_Y_c_384_n 0.00716176f $X=0.735 $Y=2.355 $X2=0 $Y2=0
cc_123 N_A_27_507#_c_120_n N_Y_c_384_n 0.00290726f $X=1.045 $Y=1.32 $X2=0 $Y2=0
cc_124 N_A_27_507#_c_121_n N_Y_c_384_n 0.00351801f $X=1.045 $Y=1.32 $X2=0 $Y2=0
cc_125 N_A_27_507#_c_122_n N_Y_c_385_n 3.89067e-19 $X=1.4 $Y=1.75 $X2=0 $Y2=0
cc_126 N_A_27_507#_c_122_n N_Y_c_389_n 3.96977e-19 $X=1.4 $Y=1.75 $X2=0 $Y2=0
cc_127 N_A_27_507#_c_123_n N_Y_c_389_n 0.00694507f $X=1.21 $Y=1.75 $X2=0 $Y2=0
cc_128 N_A_27_507#_M1003_g N_Y_c_389_n 0.00798574f $X=1.475 $Y=2.195 $X2=0 $Y2=0
cc_129 N_A_27_507#_c_129_n N_Y_c_389_n 0.0119873f $X=0.735 $Y=2.355 $X2=0 $Y2=0
cc_130 N_A_27_507#_c_130_n N_Y_c_389_n 0.00238204f $X=0.89 $Y=1.825 $X2=0 $Y2=0
cc_131 N_A_27_507#_c_116_n N_Y_c_403_n 0.00358665f $X=1.045 $Y=1.155 $X2=0 $Y2=0
cc_132 N_A_27_507#_c_118_n N_Y_c_403_n 0.00109094f $X=0.38 $Y=0.9 $X2=0 $Y2=0
cc_133 N_A_27_507#_c_120_n N_Y_c_403_n 9.87196e-19 $X=1.045 $Y=1.32 $X2=0 $Y2=0
cc_134 N_A_27_507#_c_121_n N_Y_c_403_n 0.00188037f $X=1.045 $Y=1.32 $X2=0 $Y2=0
cc_135 N_A_27_507#_c_116_n N_Y_c_386_n 0.00109821f $X=1.045 $Y=1.155 $X2=0 $Y2=0
cc_136 N_A_27_507#_c_120_n N_Y_c_386_n 0.0110105f $X=1.045 $Y=1.32 $X2=0 $Y2=0
cc_137 N_A_27_507#_c_121_n N_Y_c_386_n 9.63221e-19 $X=1.045 $Y=1.32 $X2=0 $Y2=0
cc_138 N_A_27_507#_c_116_n N_VGND_c_441_n 0.0032771f $X=1.045 $Y=1.155 $X2=0
+ $Y2=0
cc_139 N_A_27_507#_c_120_n N_VGND_c_441_n 0.0139845f $X=1.045 $Y=1.32 $X2=0
+ $Y2=0
cc_140 N_A_27_507#_c_121_n N_VGND_c_441_n 0.00140352f $X=1.045 $Y=1.32 $X2=0
+ $Y2=0
cc_141 N_A_27_507#_c_116_n N_VGND_c_442_n 0.00415323f $X=1.045 $Y=1.155 $X2=0
+ $Y2=0
cc_142 N_A_27_507#_c_116_n N_VGND_c_450_n 0.00469432f $X=1.045 $Y=1.155 $X2=0
+ $Y2=0
cc_143 N_A_27_507#_c_118_n N_VGND_c_450_n 0.0125263f $X=0.38 $Y=0.9 $X2=0 $Y2=0
cc_144 N_B_M1011_g N_A_c_223_n 0.0145431f $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_145 B N_A_c_223_n 0.0112934f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_146 N_B_c_191_n N_A_c_223_n 0.00129249f $X=2.175 $Y=0.35 $X2=0 $Y2=0
cc_147 N_B_M1011_g A 0.0033227f $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_148 B A 0.00401499f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_149 N_B_M1011_g N_A_c_225_n 0.0879648f $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_150 N_B_M1011_g N_A_284_99#_M1008_g 0.0092508f $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_151 N_B_c_191_n N_A_284_99#_M1008_g 4.18489e-19 $X=2.175 $Y=0.35 $X2=0 $Y2=0
cc_152 N_B_M1011_g N_A_284_99#_c_256_n 0.0801525f $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_153 N_B_M1011_g N_A_284_99#_c_262_n 0.00971367f $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_154 B N_Y_M1011_d 0.00189492f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_155 N_B_M1011_g N_Y_c_384_n 4.41091e-19 $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_156 N_B_M1011_g N_Y_c_385_n 6.53653e-19 $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_157 B N_Y_c_385_n 0.00221604f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_158 N_B_c_191_n N_Y_c_385_n 2.92753e-19 $X=2.175 $Y=0.35 $X2=0 $Y2=0
cc_159 N_B_M1011_g Y 0.0208781f $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_160 B Y 0.00833892f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_161 N_B_M1011_g N_Y_c_417_n 0.00243793f $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_162 B N_Y_c_417_n 0.0143434f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_163 N_B_c_191_n N_Y_c_417_n 2.51821e-19 $X=2.175 $Y=0.35 $X2=0 $Y2=0
cc_164 B N_VGND_M1008_d 0.00109537f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_165 N_B_M1011_g N_VGND_c_443_n 0.00464765f $X=2.195 $Y=0.835 $X2=0 $Y2=0
cc_166 B N_VGND_c_443_n 0.0291828f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_167 N_B_c_191_n N_VGND_c_443_n 0.00412556f $X=2.175 $Y=0.35 $X2=0 $Y2=0
cc_168 B N_VGND_c_444_n 0.0296805f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_169 N_B_c_191_n N_VGND_c_444_n 0.00210322f $X=2.175 $Y=0.35 $X2=0 $Y2=0
cc_170 B N_VGND_c_447_n 0.0447899f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_171 N_B_c_191_n N_VGND_c_447_n 0.00651318f $X=2.175 $Y=0.35 $X2=0 $Y2=0
cc_172 B N_VGND_c_450_n 0.0257035f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_173 N_B_c_191_n N_VGND_c_450_n 0.0100951f $X=2.175 $Y=0.35 $X2=0 $Y2=0
cc_174 N_A_M1001_g N_A_284_99#_c_262_n 0.00971367f $X=2.555 $Y=2.195 $X2=0 $Y2=0
cc_175 N_A_c_224_n N_C_N_c_313_n 0.0140329f $X=2.645 $Y=1.66 $X2=0 $Y2=0
cc_176 N_A_M1001_g N_C_N_M1007_g 0.00685291f $X=2.555 $Y=2.195 $X2=0 $Y2=0
cc_177 N_A_c_227_n N_C_N_c_314_n 0.0140329f $X=2.645 $Y=1.825 $X2=0 $Y2=0
cc_178 N_A_M1001_g C_N 0.00593542f $X=2.555 $Y=2.195 $X2=0 $Y2=0
cc_179 A C_N 0.0314511f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A_c_225_n C_N 0.00273341f $X=2.645 $Y=1.32 $X2=0 $Y2=0
cc_181 A N_C_N_c_316_n 0.00194131f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A_c_225_n N_C_N_c_316_n 0.0140329f $X=2.645 $Y=1.32 $X2=0 $Y2=0
cc_183 N_A_c_223_n N_C_N_c_317_n 0.0123825f $X=2.645 $Y=1.155 $X2=0 $Y2=0
cc_184 N_A_M1001_g N_VPWR_c_351_n 0.00374707f $X=2.555 $Y=2.195 $X2=0 $Y2=0
cc_185 N_A_c_227_n N_VPWR_c_351_n 0.00363594f $X=2.645 $Y=1.825 $X2=0 $Y2=0
cc_186 A N_VPWR_c_351_n 0.00626794f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_187 N_A_c_223_n Y 7.28744e-19 $X=2.645 $Y=1.155 $X2=0 $Y2=0
cc_188 A Y 0.00413485f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A_c_225_n Y 6.25133e-19 $X=2.645 $Y=1.32 $X2=0 $Y2=0
cc_190 N_A_c_223_n N_Y_c_417_n 0.00393005f $X=2.645 $Y=1.155 $X2=0 $Y2=0
cc_191 A N_Y_c_417_n 0.00476558f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A_c_225_n N_Y_c_417_n 0.00181669f $X=2.645 $Y=1.32 $X2=0 $Y2=0
cc_193 N_A_c_223_n N_VGND_c_444_n 0.00547814f $X=2.645 $Y=1.155 $X2=0 $Y2=0
cc_194 N_A_c_223_n N_VGND_c_447_n 5.42344e-19 $X=2.645 $Y=1.155 $X2=0 $Y2=0
cc_195 N_A_284_99#_c_264_n N_C_N_M1007_g 0.00177027f $X=3.45 $Y=2.94 $X2=0 $Y2=0
cc_196 N_A_284_99#_c_266_n N_C_N_M1007_g 0.00740777f $X=3.2 $Y=2.85 $X2=0 $Y2=0
cc_197 N_A_284_99#_c_264_n C_N 0.00902417f $X=3.45 $Y=2.94 $X2=0 $Y2=0
cc_198 N_A_284_99#_c_259_n C_N 0.0788738f $X=3.535 $Y=2.13 $X2=0 $Y2=0
cc_199 N_A_284_99#_c_260_n C_N 0.00103343f $X=3.545 $Y=0.87 $X2=0 $Y2=0
cc_200 N_A_284_99#_c_266_n C_N 0.00484813f $X=3.2 $Y=2.85 $X2=0 $Y2=0
cc_201 N_A_284_99#_c_259_n N_C_N_c_316_n 0.0259535f $X=3.535 $Y=2.13 $X2=0 $Y2=0
cc_202 N_A_284_99#_c_260_n N_C_N_c_316_n 0.00379389f $X=3.545 $Y=0.87 $X2=0
+ $Y2=0
cc_203 N_A_284_99#_c_259_n N_C_N_c_317_n 0.00504403f $X=3.535 $Y=2.13 $X2=0
+ $Y2=0
cc_204 N_A_284_99#_c_260_n N_C_N_c_317_n 0.00374612f $X=3.545 $Y=0.87 $X2=0
+ $Y2=0
cc_205 N_A_284_99#_c_262_n N_VPWR_c_351_n 0.0209757f $X=3.035 $Y=2.85 $X2=0
+ $Y2=0
cc_206 N_A_284_99#_c_264_n N_VPWR_c_351_n 0.0125751f $X=3.45 $Y=2.94 $X2=0 $Y2=0
cc_207 N_A_284_99#_c_259_n N_VPWR_c_351_n 0.0113502f $X=3.535 $Y=2.13 $X2=0
+ $Y2=0
cc_208 N_A_284_99#_c_266_n N_VPWR_c_351_n 0.00355239f $X=3.2 $Y=2.85 $X2=0 $Y2=0
cc_209 N_A_284_99#_c_263_n N_VPWR_c_352_n 0.023416f $X=1.91 $Y=2.85 $X2=0 $Y2=0
cc_210 N_A_284_99#_c_262_n N_VPWR_c_355_n 0.00445258f $X=3.035 $Y=2.85 $X2=0
+ $Y2=0
cc_211 N_A_284_99#_c_264_n N_VPWR_c_355_n 0.0297446f $X=3.45 $Y=2.94 $X2=0 $Y2=0
cc_212 N_A_284_99#_c_266_n N_VPWR_c_355_n 0.00593936f $X=3.2 $Y=2.85 $X2=0 $Y2=0
cc_213 N_A_284_99#_c_263_n N_VPWR_c_349_n 0.0295626f $X=1.91 $Y=2.85 $X2=0 $Y2=0
cc_214 N_A_284_99#_c_264_n N_VPWR_c_349_n 0.0207657f $X=3.45 $Y=2.94 $X2=0 $Y2=0
cc_215 N_A_284_99#_c_266_n N_VPWR_c_349_n 0.00809242f $X=3.2 $Y=2.85 $X2=0 $Y2=0
cc_216 N_A_284_99#_M1008_g N_Y_c_383_n 0.00386437f $X=1.495 $Y=0.835 $X2=0 $Y2=0
cc_217 N_A_284_99#_c_257_n N_Y_c_384_n 0.0050513f $X=1.57 $Y=1.36 $X2=0 $Y2=0
cc_218 N_A_284_99#_M1006_g N_Y_c_384_n 0.00685134f $X=1.835 $Y=2.195 $X2=0 $Y2=0
cc_219 N_A_284_99#_M1008_g N_Y_c_385_n 0.00996382f $X=1.495 $Y=0.835 $X2=0 $Y2=0
cc_220 N_A_284_99#_c_256_n N_Y_c_385_n 0.0152958f $X=1.76 $Y=1.36 $X2=0 $Y2=0
cc_221 N_A_284_99#_M1006_g N_Y_c_389_n 0.00117271f $X=1.835 $Y=2.195 $X2=0 $Y2=0
cc_222 N_A_284_99#_M1008_g N_Y_c_403_n 0.00448139f $X=1.495 $Y=0.835 $X2=0 $Y2=0
cc_223 N_A_284_99#_M1008_g N_Y_c_386_n 0.00180186f $X=1.495 $Y=0.835 $X2=0 $Y2=0
cc_224 N_A_284_99#_M1008_g Y 8.71479e-19 $X=1.495 $Y=0.835 $X2=0 $Y2=0
cc_225 N_A_284_99#_c_260_n N_Y_c_417_n 9.30852e-19 $X=3.545 $Y=0.87 $X2=0 $Y2=0
cc_226 N_A_284_99#_M1008_g N_VGND_c_442_n 0.00415323f $X=1.495 $Y=0.835 $X2=0
+ $Y2=0
cc_227 N_A_284_99#_M1008_g N_VGND_c_443_n 0.00645844f $X=1.495 $Y=0.835 $X2=0
+ $Y2=0
cc_228 N_A_284_99#_M1008_g N_VGND_c_450_n 0.00469432f $X=1.495 $Y=0.835 $X2=0
+ $Y2=0
cc_229 N_A_284_99#_c_260_n N_VGND_c_450_n 0.01437f $X=3.545 $Y=0.87 $X2=0 $Y2=0
cc_230 C_N N_VPWR_M1001_d 0.005299f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_231 N_C_N_M1007_g N_VPWR_c_351_n 0.00133958f $X=3.32 $Y=2.195 $X2=0 $Y2=0
cc_232 C_N N_VPWR_c_351_n 0.0272136f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_233 N_C_N_c_317_n N_Y_c_417_n 3.11132e-19 $X=3.207 $Y=1.155 $X2=0 $Y2=0
cc_234 C_N N_VGND_c_444_n 0.00268143f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_235 N_C_N_c_316_n N_VGND_c_444_n 0.00101269f $X=3.185 $Y=1.32 $X2=0 $Y2=0
cc_236 N_C_N_c_317_n N_VGND_c_444_n 0.00332466f $X=3.207 $Y=1.155 $X2=0 $Y2=0
cc_237 N_C_N_c_317_n N_VGND_c_449_n 0.00415323f $X=3.207 $Y=1.155 $X2=0 $Y2=0
cc_238 N_C_N_c_317_n N_VGND_c_450_n 0.00469432f $X=3.207 $Y=1.155 $X2=0 $Y2=0
cc_239 N_Y_c_385_n N_VGND_c_443_n 0.0133239f $X=2.075 $Y=1.2 $X2=0 $Y2=0
cc_240 N_Y_c_403_n N_VGND_c_443_n 0.0120901f $X=1.395 $Y=0.87 $X2=0 $Y2=0
cc_241 N_Y_c_417_n N_VGND_c_444_n 0.0044031f $X=2.41 $Y=0.92 $X2=0 $Y2=0
cc_242 N_Y_c_403_n N_VGND_c_450_n 0.0133746f $X=1.395 $Y=0.87 $X2=0 $Y2=0
