* File: sky130_fd_sc_lp__buflp_4.pxi.spice
* Created: Fri Aug 28 10:12:39 2020
* 
x_PM_SKY130_FD_SC_LP__BUFLP_4%A_84_21# N_A_84_21#_M1006_d N_A_84_21#_M1008_d
+ N_A_84_21#_M1003_g N_A_84_21#_M1000_g N_A_84_21#_M1004_g N_A_84_21#_M1011_g
+ N_A_84_21#_M1014_g N_A_84_21#_M1012_g N_A_84_21#_M1001_g N_A_84_21#_M1007_g
+ N_A_84_21#_M1002_g N_A_84_21#_M1010_g N_A_84_21#_M1009_g N_A_84_21#_M1013_g
+ N_A_84_21#_M1015_g N_A_84_21#_M1017_g N_A_84_21#_M1016_g N_A_84_21#_M1019_g
+ N_A_84_21#_c_171_p N_A_84_21#_c_91_n N_A_84_21#_c_107_p N_A_84_21#_c_217_p
+ N_A_84_21#_c_92_n N_A_84_21#_c_93_n N_A_84_21#_c_94_n N_A_84_21#_c_95_n
+ PM_SKY130_FD_SC_LP__BUFLP_4%A_84_21#
x_PM_SKY130_FD_SC_LP__BUFLP_4%A N_A_M1005_g N_A_M1018_g N_A_c_270_n N_A_c_271_n
+ N_A_M1006_g N_A_M1008_g N_A_c_273_n A N_A_c_274_n N_A_c_275_n N_A_c_276_n
+ PM_SKY130_FD_SC_LP__BUFLP_4%A
x_PM_SKY130_FD_SC_LP__BUFLP_4%VPWR N_VPWR_M1000_d N_VPWR_M1011_d N_VPWR_M1019_d
+ N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n VPWR
+ N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_314_n N_VPWR_c_323_n
+ N_VPWR_c_324_n PM_SKY130_FD_SC_LP__BUFLP_4%VPWR
x_PM_SKY130_FD_SC_LP__BUFLP_4%A_114_367# N_A_114_367#_M1000_s
+ N_A_114_367#_M1012_s N_A_114_367#_M1010_s N_A_114_367#_M1017_s
+ N_A_114_367#_c_383_n N_A_114_367#_c_385_n N_A_114_367#_c_387_n
+ N_A_114_367#_c_391_n N_A_114_367#_c_393_n N_A_114_367#_c_395_n
+ N_A_114_367#_c_397_n N_A_114_367#_c_399_n N_A_114_367#_c_382_n
+ N_A_114_367#_c_405_n N_A_114_367#_c_408_n
+ PM_SKY130_FD_SC_LP__BUFLP_4%A_114_367#
x_PM_SKY130_FD_SC_LP__BUFLP_4%X N_X_M1001_d N_X_M1009_d N_X_M1007_d N_X_M1013_d
+ N_X_c_440_n N_X_c_441_n N_X_c_445_n N_X_c_463_n N_X_c_442_n N_X_c_446_n
+ N_X_c_524_p N_X_c_443_n N_X_c_447_n N_X_c_448_n X X X
+ PM_SKY130_FD_SC_LP__BUFLP_4%X
x_PM_SKY130_FD_SC_LP__BUFLP_4%VGND N_VGND_M1003_d N_VGND_M1004_d N_VGND_M1016_d
+ N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n N_VGND_c_530_n N_VGND_c_531_n
+ N_VGND_c_532_n VGND N_VGND_c_533_n N_VGND_c_534_n N_VGND_c_535_n
+ N_VGND_c_536_n PM_SKY130_FD_SC_LP__BUFLP_4%VGND
x_PM_SKY130_FD_SC_LP__BUFLP_4%A_114_47# N_A_114_47#_M1003_s N_A_114_47#_M1014_s
+ N_A_114_47#_M1002_s N_A_114_47#_M1015_s N_A_114_47#_c_604_n
+ N_A_114_47#_c_605_n N_A_114_47#_c_607_n N_A_114_47#_c_608_n
+ N_A_114_47#_c_651_n N_A_114_47#_c_610_n N_A_114_47#_c_614_n
+ N_A_114_47#_c_616_n N_A_114_47#_c_603_n PM_SKY130_FD_SC_LP__BUFLP_4%A_114_47#
cc_1 VNB N_A_84_21#_M1003_g 0.0265231f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_2 VNB N_A_84_21#_M1000_g 4.92413e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_3 VNB N_A_84_21#_M1004_g 0.0219739f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_4 VNB N_A_84_21#_M1011_g 4.57346e-19 $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_5 VNB N_A_84_21#_M1014_g 0.0219982f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_6 VNB N_A_84_21#_M1012_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=2.465
cc_7 VNB N_A_84_21#_M1001_g 0.0221931f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.655
cc_8 VNB N_A_84_21#_M1007_g 4.82594e-19 $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=2.465
cc_9 VNB N_A_84_21#_M1002_g 0.0221973f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.655
cc_10 VNB N_A_84_21#_M1010_g 5.07481e-19 $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=2.465
cc_11 VNB N_A_84_21#_M1009_g 0.0221973f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_12 VNB N_A_84_21#_M1013_g 5.07481e-19 $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=2.465
cc_13 VNB N_A_84_21#_M1015_g 0.0226849f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=0.655
cc_14 VNB N_A_84_21#_M1017_g 5.07481e-19 $X=-0.19 $Y=-0.245 $X2=3.285 $Y2=2.465
cc_15 VNB N_A_84_21#_M1016_g 0.0265215f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=0.655
cc_16 VNB N_A_84_21#_M1019_g 5.41957e-19 $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=2.465
cc_17 VNB N_A_84_21#_c_91_n 0.00462096f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.315
cc_18 VNB N_A_84_21#_c_92_n 0.0223136f $X=-0.19 $Y=-0.245 $X2=4.96 $Y2=0.42
cc_19 VNB N_A_84_21#_c_93_n 0.026706f $X=-0.19 $Y=-0.245 $X2=4.96 $Y2=1.98
cc_20 VNB N_A_84_21#_c_94_n 0.00704942f $X=-0.19 $Y=-0.245 $X2=4.96 $Y2=0.925
cc_21 VNB N_A_84_21#_c_95_n 0.18684f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=1.48
cc_22 VNB N_A_M1018_g 0.00772229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_c_270_n 0.00795562f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_24 VNB N_A_c_271_n 0.0196285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_M1008_g 0.0192211f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.315
cc_26 VNB N_A_c_273_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_27 VNB N_A_c_274_n 0.0296313f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_28 VNB N_A_c_275_n 0.0186567f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_29 VNB N_A_c_276_n 0.00806568f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_30 VNB N_VPWR_c_314_n 0.223389f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.315
cc_31 VNB N_X_c_440_n 0.00852879f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_32 VNB N_X_c_441_n 0.00735212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_442_n 0.00524855f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.315
cc_34 VNB N_X_c_443_n 0.00177196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB X 0.0258508f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.315
cc_36 VNB N_VGND_c_527_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_528_n 0.0257496f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_38 VNB N_VGND_c_529_n 4.12476e-19 $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_39 VNB N_VGND_c_530_n 0.00558101f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_40 VNB N_VGND_c_531_n 0.0527389f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.315
cc_41 VNB N_VGND_c_532_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_42 VNB N_VGND_c_533_n 0.015032f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.645
cc_43 VNB N_VGND_c_534_n 0.0410942f $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=1.645
cc_44 VNB N_VGND_c_535_n 0.270983f $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=2.465
cc_45 VNB N_VGND_c_536_n 0.00436154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_114_47#_c_603_n 0.0025378f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.645
cc_47 VPB N_A_84_21#_M1000_g 0.0231375f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_48 VPB N_A_84_21#_M1011_g 0.0195909f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_49 VPB N_A_84_21#_M1012_g 0.0196149f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_50 VPB N_A_84_21#_M1007_g 0.0204614f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_51 VPB N_A_84_21#_M1010_g 0.0213036f $X=-0.19 $Y=1.655 $X2=2.285 $Y2=2.465
cc_52 VPB N_A_84_21#_M1013_g 0.0213079f $X=-0.19 $Y=1.655 $X2=2.785 $Y2=2.465
cc_53 VPB N_A_84_21#_M1017_g 0.0214038f $X=-0.19 $Y=1.655 $X2=3.285 $Y2=2.465
cc_54 VPB N_A_84_21#_M1019_g 0.0224232f $X=-0.19 $Y=1.655 $X2=3.785 $Y2=2.465
cc_55 VPB N_A_84_21#_c_93_n 0.0547566f $X=-0.19 $Y=1.655 $X2=4.96 $Y2=1.98
cc_56 VPB N_A_M1018_g 0.0211333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_M1008_g 0.0239109f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.315
cc_58 VPB N_VPWR_c_315_n 0.0106521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_316_n 0.0399534f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_60 VPB N_VPWR_c_317_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_61 VPB N_VPWR_c_318_n 0.0111167f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_62 VPB N_VPWR_c_319_n 0.0185788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_320_n 0.0624782f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=1.315
cc_64 VPB N_VPWR_c_321_n 0.0321841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_314_n 0.047538f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=1.315
cc_66 VPB N_VPWR_c_323_n 0.00324402f $X=-0.19 $Y=1.655 $X2=2.285 $Y2=2.465
cc_67 VPB N_VPWR_c_324_n 0.00631788f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=0.655
cc_68 VPB N_A_114_367#_c_382_n 0.00244912f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_69 VPB N_X_c_445_n 0.008933f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.315
cc_70 VPB N_X_c_446_n 0.00307912f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=0.655
cc_71 VPB N_X_c_447_n 0.00231148f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_72 VPB N_X_c_448_n 0.00231148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB X 4.43907e-19 $X=-0.19 $Y=1.655 $X2=2.215 $Y2=1.315
cc_74 VPB X 0.00889493f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=0.655
cc_75 N_A_84_21#_c_91_n N_A_M1018_g 6.48922e-19 $X=3.71 $Y=1.315 $X2=0 $Y2=0
cc_76 N_A_84_21#_c_95_n N_A_M1018_g 0.0389167f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_77 N_A_84_21#_c_107_p N_A_c_270_n 0.00204314f $X=4.795 $Y=0.925 $X2=0 $Y2=0
cc_78 N_A_84_21#_c_107_p N_A_c_271_n 0.0121759f $X=4.795 $Y=0.925 $X2=0 $Y2=0
cc_79 N_A_84_21#_c_92_n N_A_c_271_n 0.0129683f $X=4.96 $Y=0.42 $X2=0 $Y2=0
cc_80 N_A_84_21#_c_93_n N_A_c_271_n 0.00520624f $X=4.96 $Y=1.98 $X2=0 $Y2=0
cc_81 N_A_84_21#_c_94_n N_A_c_271_n 3.84191e-19 $X=4.96 $Y=0.925 $X2=0 $Y2=0
cc_82 N_A_84_21#_c_93_n N_A_M1008_g 0.0435091f $X=4.96 $Y=1.98 $X2=0 $Y2=0
cc_83 N_A_84_21#_c_93_n N_A_c_273_n 0.00657491f $X=4.96 $Y=1.98 $X2=0 $Y2=0
cc_84 N_A_84_21#_M1016_g N_A_c_274_n 0.00204876f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_85 N_A_84_21#_c_91_n N_A_c_274_n 5.22367e-19 $X=3.71 $Y=1.315 $X2=0 $Y2=0
cc_86 N_A_84_21#_c_107_p N_A_c_274_n 0.00112859f $X=4.795 $Y=0.925 $X2=0 $Y2=0
cc_87 N_A_84_21#_c_93_n N_A_c_274_n 0.00536769f $X=4.96 $Y=1.98 $X2=0 $Y2=0
cc_88 N_A_84_21#_c_95_n N_A_c_274_n 0.0110745f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_89 N_A_84_21#_M1016_g N_A_c_275_n 0.0126844f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_90 N_A_84_21#_c_91_n N_A_c_275_n 0.00283069f $X=3.71 $Y=1.315 $X2=0 $Y2=0
cc_91 N_A_84_21#_c_107_p N_A_c_275_n 0.0131732f $X=4.795 $Y=0.925 $X2=0 $Y2=0
cc_92 N_A_84_21#_c_92_n N_A_c_275_n 0.00289686f $X=4.96 $Y=0.42 $X2=0 $Y2=0
cc_93 N_A_84_21#_c_93_n N_A_c_275_n 8.44691e-19 $X=4.96 $Y=1.98 $X2=0 $Y2=0
cc_94 N_A_84_21#_c_91_n N_A_c_276_n 0.0281543f $X=3.71 $Y=1.315 $X2=0 $Y2=0
cc_95 N_A_84_21#_c_107_p N_A_c_276_n 0.0332393f $X=4.795 $Y=0.925 $X2=0 $Y2=0
cc_96 N_A_84_21#_c_93_n N_A_c_276_n 0.0138664f $X=4.96 $Y=1.98 $X2=0 $Y2=0
cc_97 N_A_84_21#_c_95_n N_A_c_276_n 0.00156678f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_98 N_A_84_21#_M1000_g N_VPWR_c_316_n 0.009097f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_84_21#_M1011_g N_VPWR_c_317_n 0.00359601f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_100 N_A_84_21#_M1012_g N_VPWR_c_317_n 0.00359601f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_101 N_A_84_21#_M1019_g N_VPWR_c_318_n 0.0109958f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_102 N_A_84_21#_c_93_n N_VPWR_c_318_n 0.0180682f $X=4.96 $Y=1.98 $X2=0 $Y2=0
cc_103 N_A_84_21#_M1000_g N_VPWR_c_319_n 0.0054895f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_A_84_21#_M1011_g N_VPWR_c_319_n 0.0054895f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_105 N_A_84_21#_M1012_g N_VPWR_c_320_n 0.00547432f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_106 N_A_84_21#_M1007_g N_VPWR_c_320_n 0.00357842f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_107 N_A_84_21#_M1010_g N_VPWR_c_320_n 0.00357877f $X=2.285 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_A_84_21#_M1013_g N_VPWR_c_320_n 0.00357842f $X=2.785 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_A_84_21#_M1017_g N_VPWR_c_320_n 0.00357877f $X=3.285 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_84_21#_M1019_g N_VPWR_c_320_n 0.00547432f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_111 N_A_84_21#_c_93_n N_VPWR_c_321_n 0.0210192f $X=4.96 $Y=1.98 $X2=0 $Y2=0
cc_112 N_A_84_21#_M1008_d N_VPWR_c_314_n 0.00231914f $X=4.82 $Y=1.835 $X2=0
+ $Y2=0
cc_113 N_A_84_21#_M1000_g N_VPWR_c_314_n 0.010744f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A_84_21#_M1011_g N_VPWR_c_314_n 0.00990036f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_115 N_A_84_21#_M1012_g N_VPWR_c_314_n 0.0098633f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_84_21#_M1007_g N_VPWR_c_314_n 0.00553547f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_84_21#_M1010_g N_VPWR_c_314_n 0.0057905f $X=2.285 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_84_21#_M1013_g N_VPWR_c_314_n 0.00570659f $X=2.785 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_A_84_21#_M1017_g N_VPWR_c_314_n 0.0057905f $X=3.285 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_84_21#_M1019_g N_VPWR_c_314_n 0.0103577f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_A_84_21#_c_93_n N_VPWR_c_314_n 0.0125689f $X=4.96 $Y=1.98 $X2=0 $Y2=0
cc_122 N_A_84_21#_M1011_g N_A_114_367#_c_383_n 0.01115f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_84_21#_M1012_g N_A_114_367#_c_383_n 0.01115f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_124 N_A_84_21#_M1012_g N_A_114_367#_c_385_n 7.32094e-19 $X=1.355 $Y=2.465
+ $X2=0 $Y2=0
cc_125 N_A_84_21#_M1007_g N_A_114_367#_c_385_n 0.00209265f $X=1.785 $Y=2.465
+ $X2=0 $Y2=0
cc_126 N_A_84_21#_M1011_g N_A_114_367#_c_387_n 6.2172e-19 $X=0.925 $Y=2.465
+ $X2=0 $Y2=0
cc_127 N_A_84_21#_M1012_g N_A_114_367#_c_387_n 0.00958318f $X=1.355 $Y=2.465
+ $X2=0 $Y2=0
cc_128 N_A_84_21#_M1007_g N_A_114_367#_c_387_n 0.00996263f $X=1.785 $Y=2.465
+ $X2=0 $Y2=0
cc_129 N_A_84_21#_M1010_g N_A_114_367#_c_387_n 5.82363e-19 $X=2.285 $Y=2.465
+ $X2=0 $Y2=0
cc_130 N_A_84_21#_M1007_g N_A_114_367#_c_391_n 0.0109138f $X=1.785 $Y=2.465
+ $X2=0 $Y2=0
cc_131 N_A_84_21#_M1010_g N_A_114_367#_c_391_n 0.0143648f $X=2.285 $Y=2.465
+ $X2=0 $Y2=0
cc_132 N_A_84_21#_M1012_g N_A_114_367#_c_393_n 0.00197018f $X=1.355 $Y=2.465
+ $X2=0 $Y2=0
cc_133 N_A_84_21#_M1007_g N_A_114_367#_c_393_n 5.89773e-19 $X=1.785 $Y=2.465
+ $X2=0 $Y2=0
cc_134 N_A_84_21#_M1013_g N_A_114_367#_c_395_n 0.0120553f $X=2.785 $Y=2.465
+ $X2=0 $Y2=0
cc_135 N_A_84_21#_M1017_g N_A_114_367#_c_395_n 6.92322e-19 $X=3.285 $Y=2.465
+ $X2=0 $Y2=0
cc_136 N_A_84_21#_M1013_g N_A_114_367#_c_397_n 0.0109138f $X=2.785 $Y=2.465
+ $X2=0 $Y2=0
cc_137 N_A_84_21#_M1017_g N_A_114_367#_c_397_n 0.0143648f $X=3.285 $Y=2.465
+ $X2=0 $Y2=0
cc_138 N_A_84_21#_M1019_g N_A_114_367#_c_399_n 0.00196648f $X=3.785 $Y=2.465
+ $X2=0 $Y2=0
cc_139 N_A_84_21#_M1017_g N_A_114_367#_c_382_n 0.00574467f $X=3.285 $Y=2.465
+ $X2=0 $Y2=0
cc_140 N_A_84_21#_M1019_g N_A_114_367#_c_382_n 0.0136231f $X=3.785 $Y=2.465
+ $X2=0 $Y2=0
cc_141 N_A_84_21#_c_171_p N_A_114_367#_c_382_n 0.0184323f $X=3.625 $Y=1.48 $X2=0
+ $Y2=0
cc_142 N_A_84_21#_c_91_n N_A_114_367#_c_382_n 0.00961143f $X=3.71 $Y=1.315 $X2=0
+ $Y2=0
cc_143 N_A_84_21#_c_95_n N_A_114_367#_c_382_n 0.004473f $X=3.785 $Y=1.48 $X2=0
+ $Y2=0
cc_144 N_A_84_21#_M1000_g N_A_114_367#_c_405_n 0.0129871f $X=0.495 $Y=2.465
+ $X2=0 $Y2=0
cc_145 N_A_84_21#_M1011_g N_A_114_367#_c_405_n 0.0122795f $X=0.925 $Y=2.465
+ $X2=0 $Y2=0
cc_146 N_A_84_21#_M1012_g N_A_114_367#_c_405_n 6.7275e-19 $X=1.355 $Y=2.465
+ $X2=0 $Y2=0
cc_147 N_A_84_21#_M1013_g N_A_114_367#_c_408_n 5.89773e-19 $X=2.785 $Y=2.465
+ $X2=0 $Y2=0
cc_148 N_A_84_21#_M1003_g N_X_c_440_n 0.017882f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_149 N_A_84_21#_M1004_g N_X_c_440_n 0.0104926f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_150 N_A_84_21#_M1014_g N_X_c_440_n 0.0104926f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_151 N_A_84_21#_M1001_g N_X_c_440_n 0.00889811f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_152 N_A_84_21#_c_171_p N_X_c_440_n 0.0803029f $X=3.625 $Y=1.48 $X2=0 $Y2=0
cc_153 N_A_84_21#_c_95_n N_X_c_440_n 0.00714474f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_154 N_A_84_21#_M1000_g N_X_c_445_n 0.0177123f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_84_21#_M1011_g N_X_c_445_n 0.010445f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A_84_21#_M1012_g N_X_c_445_n 0.0104915f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_84_21#_M1007_g N_X_c_445_n 0.0147025f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_84_21#_c_171_p N_X_c_445_n 0.0854672f $X=3.625 $Y=1.48 $X2=0 $Y2=0
cc_159 N_A_84_21#_c_95_n N_X_c_445_n 0.00714474f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_160 N_A_84_21#_M1014_g N_X_c_463_n 9.1803e-19 $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_161 N_A_84_21#_M1001_g N_X_c_463_n 0.00599327f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A_84_21#_M1002_g N_X_c_442_n 0.0111824f $X=2.215 $Y=0.655 $X2=0 $Y2=0
cc_163 N_A_84_21#_M1009_g N_X_c_442_n 0.0109305f $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_164 N_A_84_21#_M1015_g N_X_c_442_n 0.00189142f $X=3.075 $Y=0.655 $X2=0 $Y2=0
cc_165 N_A_84_21#_c_171_p N_X_c_442_n 0.0647563f $X=3.625 $Y=1.48 $X2=0 $Y2=0
cc_166 N_A_84_21#_c_95_n N_X_c_442_n 0.00522367f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_167 N_A_84_21#_M1010_g N_X_c_446_n 0.0115433f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A_84_21#_M1013_g N_X_c_446_n 0.0151263f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_84_21#_c_171_p N_X_c_446_n 0.0492574f $X=3.625 $Y=1.48 $X2=0 $Y2=0
cc_170 N_A_84_21#_c_95_n N_X_c_446_n 0.00436308f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_171 N_A_84_21#_M1001_g N_X_c_443_n 0.00199293f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_172 N_A_84_21#_c_171_p N_X_c_443_n 0.0206129f $X=3.625 $Y=1.48 $X2=0 $Y2=0
cc_173 N_A_84_21#_c_95_n N_X_c_443_n 0.00231141f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_174 N_A_84_21#_M1010_g N_X_c_447_n 0.0130701f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A_84_21#_M1013_g N_X_c_447_n 6.92322e-19 $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_84_21#_c_171_p N_X_c_447_n 0.02772f $X=3.625 $Y=1.48 $X2=0 $Y2=0
cc_177 N_A_84_21#_c_95_n N_X_c_447_n 0.00423635f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_178 N_A_84_21#_M1017_g N_X_c_448_n 0.0127819f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A_84_21#_M1019_g N_X_c_448_n 2.46243e-19 $X=3.785 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_84_21#_c_171_p N_X_c_448_n 0.02772f $X=3.625 $Y=1.48 $X2=0 $Y2=0
cc_181 N_A_84_21#_c_95_n N_X_c_448_n 0.00463077f $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_182 N_A_84_21#_M1003_g X 0.0184476f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_183 N_A_84_21#_c_171_p X 0.014323f $X=3.625 $Y=1.48 $X2=0 $Y2=0
cc_184 N_A_84_21#_M1000_g X 0.00593253f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_84_21#_c_91_n N_VGND_M1016_d 0.00152909f $X=3.71 $Y=1.315 $X2=0 $Y2=0
cc_186 N_A_84_21#_c_107_p N_VGND_M1016_d 0.0171548f $X=4.795 $Y=0.925 $X2=0
+ $Y2=0
cc_187 N_A_84_21#_c_217_p N_VGND_M1016_d 0.00321143f $X=3.795 $Y=0.925 $X2=0
+ $Y2=0
cc_188 N_A_84_21#_M1003_g N_VGND_c_528_n 0.00655014f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_189 N_A_84_21#_M1003_g N_VGND_c_529_n 6.17145e-19 $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_190 N_A_84_21#_M1004_g N_VGND_c_529_n 0.00666323f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_191 N_A_84_21#_M1014_g N_VGND_c_529_n 0.00765587f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_192 N_A_84_21#_M1001_g N_VGND_c_529_n 0.00121664f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_193 N_A_84_21#_M1016_g N_VGND_c_530_n 0.00741201f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_194 N_A_84_21#_c_107_p N_VGND_c_530_n 0.0126179f $X=4.795 $Y=0.925 $X2=0
+ $Y2=0
cc_195 N_A_84_21#_c_217_p N_VGND_c_530_n 0.0139023f $X=3.795 $Y=0.925 $X2=0
+ $Y2=0
cc_196 N_A_84_21#_c_95_n N_VGND_c_530_n 4.99323e-19 $X=3.785 $Y=1.48 $X2=0 $Y2=0
cc_197 N_A_84_21#_M1014_g N_VGND_c_531_n 0.00353537f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_198 N_A_84_21#_M1001_g N_VGND_c_531_n 0.00357877f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_199 N_A_84_21#_M1002_g N_VGND_c_531_n 0.00357842f $X=2.215 $Y=0.655 $X2=0
+ $Y2=0
cc_200 N_A_84_21#_M1009_g N_VGND_c_531_n 0.00357842f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_201 N_A_84_21#_M1015_g N_VGND_c_531_n 0.00357842f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_202 N_A_84_21#_M1016_g N_VGND_c_531_n 0.00547432f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_203 N_A_84_21#_M1003_g N_VGND_c_533_n 0.0054895f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_204 N_A_84_21#_M1004_g N_VGND_c_533_n 0.00353537f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_205 N_A_84_21#_c_92_n N_VGND_c_534_n 0.0210192f $X=4.96 $Y=0.42 $X2=0 $Y2=0
cc_206 N_A_84_21#_M1006_d N_VGND_c_535_n 0.00231914f $X=4.82 $Y=0.235 $X2=0
+ $Y2=0
cc_207 N_A_84_21#_M1003_g N_VGND_c_535_n 0.0109952f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_208 N_A_84_21#_M1004_g N_VGND_c_535_n 0.00419187f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_209 N_A_84_21#_M1014_g N_VGND_c_535_n 0.00419187f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_210 N_A_84_21#_M1001_g N_VGND_c_535_n 0.00542194f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_211 N_A_84_21#_M1002_g N_VGND_c_535_n 0.00542192f $X=2.215 $Y=0.655 $X2=0
+ $Y2=0
cc_212 N_A_84_21#_M1009_g N_VGND_c_535_n 0.00542192f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_213 N_A_84_21#_M1015_g N_VGND_c_535_n 0.00535118f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_214 N_A_84_21#_M1016_g N_VGND_c_535_n 0.0106313f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_215 N_A_84_21#_c_107_p N_VGND_c_535_n 0.0275875f $X=4.795 $Y=0.925 $X2=0
+ $Y2=0
cc_216 N_A_84_21#_c_217_p N_VGND_c_535_n 6.15084e-19 $X=3.795 $Y=0.925 $X2=0
+ $Y2=0
cc_217 N_A_84_21#_c_92_n N_VGND_c_535_n 0.0125689f $X=4.96 $Y=0.42 $X2=0 $Y2=0
cc_218 N_A_84_21#_M1003_g N_A_114_47#_c_604_n 0.00507277f $X=0.495 $Y=0.655
+ $X2=0 $Y2=0
cc_219 N_A_84_21#_M1004_g N_A_114_47#_c_605_n 0.0104796f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_220 N_A_84_21#_M1014_g N_A_114_47#_c_605_n 0.0102994f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_221 N_A_84_21#_M1003_g N_A_114_47#_c_607_n 0.00316993f $X=0.495 $Y=0.655
+ $X2=0 $Y2=0
cc_222 N_A_84_21#_M1001_g N_A_114_47#_c_608_n 0.00993982f $X=1.785 $Y=0.655
+ $X2=0 $Y2=0
cc_223 N_A_84_21#_M1002_g N_A_114_47#_c_608_n 0.00822205f $X=2.215 $Y=0.655
+ $X2=0 $Y2=0
cc_224 N_A_84_21#_M1001_g N_A_114_47#_c_610_n 6.036e-19 $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_225 N_A_84_21#_M1002_g N_A_114_47#_c_610_n 0.00663783f $X=2.215 $Y=0.655
+ $X2=0 $Y2=0
cc_226 N_A_84_21#_M1009_g N_A_114_47#_c_610_n 0.00642675f $X=2.645 $Y=0.655
+ $X2=0 $Y2=0
cc_227 N_A_84_21#_M1015_g N_A_114_47#_c_610_n 5.62335e-19 $X=3.075 $Y=0.655
+ $X2=0 $Y2=0
cc_228 N_A_84_21#_M1009_g N_A_114_47#_c_614_n 0.00826862f $X=2.645 $Y=0.655
+ $X2=0 $Y2=0
cc_229 N_A_84_21#_M1015_g N_A_114_47#_c_614_n 0.0105205f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_230 N_A_84_21#_M1002_g N_A_114_47#_c_616_n 0.00155283f $X=2.215 $Y=0.655
+ $X2=0 $Y2=0
cc_231 N_A_84_21#_M1009_g N_A_114_47#_c_616_n 0.00155283f $X=2.645 $Y=0.655
+ $X2=0 $Y2=0
cc_232 N_A_84_21#_M1009_g N_A_114_47#_c_603_n 6.73666e-19 $X=2.645 $Y=0.655
+ $X2=0 $Y2=0
cc_233 N_A_84_21#_M1015_g N_A_114_47#_c_603_n 0.0107672f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_234 N_A_84_21#_M1016_g N_A_114_47#_c_603_n 0.0167753f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_235 N_A_84_21#_c_171_p N_A_114_47#_c_603_n 0.0225884f $X=3.625 $Y=1.48 $X2=0
+ $Y2=0
cc_236 N_A_84_21#_c_91_n N_A_114_47#_c_603_n 0.00390425f $X=3.71 $Y=1.315 $X2=0
+ $Y2=0
cc_237 N_A_84_21#_c_95_n N_A_114_47#_c_603_n 0.00264294f $X=3.785 $Y=1.48 $X2=0
+ $Y2=0
cc_238 N_A_84_21#_c_107_p A_886_47# 0.00574972f $X=4.795 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_239 N_A_M1018_g N_VPWR_c_318_n 0.011107f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_c_274_n N_VPWR_c_318_n 0.00289631f $X=4.265 $Y=1.26 $X2=0 $Y2=0
cc_241 N_A_c_276_n N_VPWR_c_318_n 0.0154623f $X=4.265 $Y=1.35 $X2=0 $Y2=0
cc_242 N_A_M1018_g N_VPWR_c_321_n 0.00585385f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A_M1008_g N_VPWR_c_321_n 0.0054895f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A_M1018_g N_VPWR_c_314_n 0.0110668f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A_M1008_g N_VPWR_c_314_n 0.0108883f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A_c_275_n N_VGND_c_530_n 0.0117137f $X=4.265 $Y=1.185 $X2=0 $Y2=0
cc_247 N_A_c_271_n N_VGND_c_534_n 0.0054895f $X=4.745 $Y=1.185 $X2=0 $Y2=0
cc_248 N_A_c_275_n N_VGND_c_534_n 0.00585385f $X=4.265 $Y=1.185 $X2=0 $Y2=0
cc_249 N_A_c_271_n N_VGND_c_535_n 0.00713607f $X=4.745 $Y=1.185 $X2=0 $Y2=0
cc_250 N_A_c_275_n N_VGND_c_535_n 0.00721186f $X=4.265 $Y=1.185 $X2=0 $Y2=0
cc_251 N_VPWR_c_314_n N_A_114_367#_M1000_s 0.00223559f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_252 N_VPWR_c_314_n N_A_114_367#_M1012_s 0.00223559f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_314_n N_A_114_367#_M1010_s 0.00280658f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_314_n N_A_114_367#_M1017_s 0.00280658f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_255 N_VPWR_M1011_d N_A_114_367#_c_383_n 0.00341793f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_256 N_VPWR_c_317_n N_A_114_367#_c_383_n 0.0135055f $X=1.14 $Y=2.805 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_320_n N_A_114_367#_c_391_n 0.0374555f $X=3.905 $Y=3.33 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_314_n N_A_114_367#_c_391_n 0.0239316f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_320_n N_A_114_367#_c_393_n 0.01906f $X=3.905 $Y=3.33 $X2=0 $Y2=0
cc_260 N_VPWR_c_314_n N_A_114_367#_c_393_n 0.0124545f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_320_n N_A_114_367#_c_397_n 0.0374555f $X=3.905 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_314_n N_A_114_367#_c_397_n 0.0239316f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_320_n N_A_114_367#_c_399_n 0.0207136f $X=3.905 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_314_n N_A_114_367#_c_399_n 0.0126368f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_318_n N_A_114_367#_c_382_n 0.0416524f $X=4.07 $Y=1.98 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_319_n N_A_114_367#_c_405_n 0.0189236f $X=1.055 $Y=3.33 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_314_n N_A_114_367#_c_405_n 0.0123859f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_320_n N_A_114_367#_c_408_n 0.0207136f $X=3.905 $Y=3.33 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_314_n N_A_114_367#_c_408_n 0.0126421f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_314_n N_X_M1007_d 0.00281482f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_271 N_VPWR_c_314_n N_X_M1013_d 0.00281482f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_M1011_d N_X_c_445_n 0.00176891f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_273 N_VPWR_c_316_n N_X_c_445_n 6.14392e-19 $X=0.28 $Y=2.32 $X2=0 $Y2=0
cc_274 N_VPWR_M1000_d X 0.00910448f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_275 N_VPWR_c_316_n X 0.0184437f $X=0.28 $Y=2.32 $X2=0 $Y2=0
cc_276 N_VPWR_c_314_n A_886_367# 0.010279f $X=5.04 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_277 N_A_114_367#_c_391_n N_X_M1007_d 0.00472489f $X=2.405 $Y=2.99 $X2=0 $Y2=0
cc_278 N_A_114_367#_c_397_n N_X_M1013_d 0.00472489f $X=3.405 $Y=2.99 $X2=0 $Y2=0
cc_279 N_A_114_367#_M1000_s N_X_c_445_n 0.00176461f $X=0.57 $Y=1.835 $X2=0 $Y2=0
cc_280 N_A_114_367#_M1012_s N_X_c_445_n 0.00176461f $X=1.43 $Y=1.835 $X2=0 $Y2=0
cc_281 N_A_114_367#_c_383_n N_X_c_445_n 0.0289344f $X=1.405 $Y=2.24 $X2=0 $Y2=0
cc_282 N_A_114_367#_c_385_n N_X_c_445_n 0.01723f $X=1.57 $Y=2.325 $X2=0 $Y2=0
cc_283 N_A_114_367#_c_405_n N_X_c_445_n 0.01723f $X=0.71 $Y=2.32 $X2=0 $Y2=0
cc_284 N_A_114_367#_M1010_s N_X_c_446_n 0.00250873f $X=2.36 $Y=1.835 $X2=0 $Y2=0
cc_285 N_A_114_367#_c_395_n N_X_c_446_n 0.0209867f $X=2.57 $Y=2.32 $X2=0 $Y2=0
cc_286 N_A_114_367#_c_391_n N_X_c_447_n 0.0196355f $X=2.405 $Y=2.99 $X2=0 $Y2=0
cc_287 N_A_114_367#_c_397_n N_X_c_448_n 0.0196355f $X=3.405 $Y=2.99 $X2=0 $Y2=0
cc_288 N_A_114_367#_c_382_n N_X_c_448_n 0.00795492f $X=3.57 $Y=1.98 $X2=0 $Y2=0
cc_289 N_X_c_441_n N_VGND_M1003_d 0.00301575f $X=0.355 $Y=1.06 $X2=-0.19
+ $Y2=-0.245
cc_290 N_X_c_440_n N_VGND_M1004_d 0.00176891f $X=1.835 $Y=1.06 $X2=0 $Y2=0
cc_291 N_X_c_440_n N_VGND_c_528_n 6.14392e-19 $X=1.835 $Y=1.06 $X2=0 $Y2=0
cc_292 N_X_c_441_n N_VGND_c_528_n 0.0207726f $X=0.355 $Y=1.06 $X2=0 $Y2=0
cc_293 N_X_M1001_d N_VGND_c_535_n 0.00225186f $X=1.86 $Y=0.235 $X2=0 $Y2=0
cc_294 N_X_M1009_d N_VGND_c_535_n 0.00225186f $X=2.72 $Y=0.235 $X2=0 $Y2=0
cc_295 N_X_c_440_n N_A_114_47#_M1003_s 0.00176461f $X=1.835 $Y=1.06 $X2=-0.19
+ $Y2=-0.245
cc_296 N_X_c_440_n N_A_114_47#_M1014_s 0.00176461f $X=1.835 $Y=1.06 $X2=0 $Y2=0
cc_297 N_X_c_442_n N_A_114_47#_M1002_s 0.00176461f $X=2.775 $Y=1.06 $X2=0 $Y2=0
cc_298 N_X_c_440_n N_A_114_47#_c_605_n 0.045666f $X=1.835 $Y=1.06 $X2=0 $Y2=0
cc_299 N_X_c_440_n N_A_114_47#_c_607_n 0.015147f $X=1.835 $Y=1.06 $X2=0 $Y2=0
cc_300 N_X_M1001_d N_A_114_47#_c_608_n 0.00332344f $X=1.86 $Y=0.235 $X2=0 $Y2=0
cc_301 N_X_c_440_n N_A_114_47#_c_608_n 0.00320534f $X=1.835 $Y=1.06 $X2=0 $Y2=0
cc_302 N_X_c_463_n N_A_114_47#_c_608_n 0.0141126f $X=2 $Y=0.845 $X2=0 $Y2=0
cc_303 N_X_c_442_n N_A_114_47#_c_608_n 0.00320534f $X=2.775 $Y=1.06 $X2=0 $Y2=0
cc_304 N_X_c_442_n N_A_114_47#_c_610_n 0.0168669f $X=2.775 $Y=1.06 $X2=0 $Y2=0
cc_305 N_X_M1009_d N_A_114_47#_c_614_n 0.00332344f $X=2.72 $Y=0.235 $X2=0 $Y2=0
cc_306 N_X_c_442_n N_A_114_47#_c_614_n 0.00320534f $X=2.775 $Y=1.06 $X2=0 $Y2=0
cc_307 N_X_c_524_p N_A_114_47#_c_614_n 0.0124309f $X=2.86 $Y=0.845 $X2=0 $Y2=0
cc_308 N_X_c_442_n N_A_114_47#_c_603_n 0.00517071f $X=2.775 $Y=1.06 $X2=0 $Y2=0
cc_309 N_VGND_c_535_n N_A_114_47#_M1003_s 0.00244093f $X=5.04 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_310 N_VGND_c_535_n N_A_114_47#_M1014_s 0.002449f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_535_n N_A_114_47#_M1002_s 0.00225167f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_535_n N_A_114_47#_M1015_s 0.00223559f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_313 N_VGND_c_533_n N_A_114_47#_c_604_n 0.0151619f $X=0.975 $Y=0 $X2=0 $Y2=0
cc_314 N_VGND_c_535_n N_A_114_47#_c_604_n 0.00947388f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_M1004_d N_A_114_47#_c_605_n 0.00334936f $X=1 $Y=0.235 $X2=0 $Y2=0
cc_316 N_VGND_c_529_n N_A_114_47#_c_605_n 0.0159984f $X=1.14 $Y=0.38 $X2=0 $Y2=0
cc_317 N_VGND_c_531_n N_A_114_47#_c_605_n 0.00256318f $X=3.625 $Y=0 $X2=0 $Y2=0
cc_318 N_VGND_c_533_n N_A_114_47#_c_605_n 0.00256318f $X=0.975 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_c_535_n N_A_114_47#_c_605_n 0.0105226f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_320 N_VGND_c_531_n N_A_114_47#_c_608_n 0.0333712f $X=3.625 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_535_n N_A_114_47#_c_608_n 0.0216758f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_531_n N_A_114_47#_c_651_n 0.0116347f $X=3.625 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_535_n N_A_114_47#_c_651_n 0.00655263f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_324 N_VGND_c_531_n N_A_114_47#_c_614_n 0.0298674f $X=3.625 $Y=0 $X2=0 $Y2=0
cc_325 N_VGND_c_535_n N_A_114_47#_c_614_n 0.0187823f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_531_n N_A_114_47#_c_616_n 0.0188964f $X=3.625 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_535_n N_A_114_47#_c_616_n 0.0125309f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_c_531_n N_A_114_47#_c_603_n 0.01906f $X=3.625 $Y=0 $X2=0 $Y2=0
cc_329 N_VGND_c_535_n N_A_114_47#_c_603_n 0.0124545f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_330 N_VGND_c_535_n A_886_47# 0.00352191f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
