* File: sky130_fd_sc_lp__dlxtn_4.spice
* Created: Wed Sep  2 09:48:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxtn_4.pex.spice"
.subckt sky130_fd_sc_lp__dlxtn_4  VNB VPB D GATE_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_D_M1007_g N_A_27_481#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.1113 PD=0.72 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_200_481#_M1008_d N_GATE_N_M1008_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.063 PD=1.37 PS=0.72 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_200_481#_M1023_g N_A_310_485#_M1023_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1009 A_574_47# N_A_27_481#_M1009_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_609_485#_M1012_d N_A_200_481#_M1012_g A_574_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=12.852 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1015 A_754_47# N_A_310_485#_M1015_g N_A_609_485#_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_795_423#_M1022_g A_754_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.0819 PD=0.823333 PS=0.81 NRD=33.564 NRS=39.996 M=1 R=2.8
+ SA=75002.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1021 N_A_795_423#_M1021_d N_A_609_485#_M1021_g N_VGND_M1022_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1848 PD=2.21 PS=1.64667 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A_795_423#_M1000_g N_Q_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_A_795_423#_M1010_g N_Q_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1010_d N_A_795_423#_M1016_g N_Q_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1018 N_VGND_M1018_d N_A_795_423#_M1018_g N_Q_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1017 N_VPWR_M1017_d N_D_M1017_g N_A_27_481#_M1017_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=6.1464 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1003 N_A_200_481#_M1003_d N_GATE_N_M1003_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_VPWR_M1014_d N_A_200_481#_M1014_g N_A_310_485#_M1014_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.176 AS=0.1824 PD=1.19 PS=1.85 NRD=83.0946 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1004 A_537_485# N_A_27_481#_M1004_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.176 PD=0.85 PS=1.19 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.9
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1020 N_A_609_485#_M1020_d N_A_310_485#_M1020_g A_537_485# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.134098 AS=0.0672 PD=1.24377 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1005 A_717_485# N_A_200_481#_M1005_g N_A_609_485#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0880019 PD=0.81 PS=0.816226 NRD=65.6601 NRS=53.9386 M=1
+ R=2.8 SA=75001.8 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A_795_423#_M1013_g A_717_485# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.135975 AS=0.0819 PD=1.0125 PS=0.81 NRD=229.82 NRS=65.6601 M=1 R=2.8
+ SA=75002.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_795_423#_M1002_d N_A_609_485#_M1002_g N_VPWR_M1013_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.407925 PD=3.05 PS=3.0375 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A_795_423#_M1001_g N_Q_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_795_423#_M1006_g N_Q_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1006_d N_A_795_423#_M1011_g N_Q_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1019_d N_A_795_423#_M1019_g N_Q_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.1151 P=20.01
*
.include "sky130_fd_sc_lp__dlxtn_4.pxi.spice"
*
.ends
*
*
