* File: sky130_fd_sc_lp__a2111o_m.spice
* Created: Wed Sep  2 09:16:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111o_m.pex.spice"
.subckt sky130_fd_sc_lp__a2111o_m  VNB VPB D1 C1 B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_85_21#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.105 AS=0.1113 PD=0.92 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1001 N_A_85_21#_M1001_d N_D1_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.105 PD=0.7 PS=0.92 NRD=0 NRS=57.132 M=1 R=2.8 SA=75000.8
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_C1_M1006_g N_A_85_21#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.3 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_85_21#_M1009_d N_B1_M1009_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1000 A_503_47# N_A1_M1000_g N_A_85_21#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g A_503_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_85_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 A_267_369# N_D1_M1011_g N_A_85_21#_M1011_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1003 A_339_369# N_C1_M1003_g A_267_369# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1008 N_A_411_369#_M1008_d N_B1_M1008_g A_339_369# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.9
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_411_369#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_411_369#_M1004_d N_A2_M1004_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=18.7544 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a2111o_m.pxi.spice"
*
.ends
*
*
