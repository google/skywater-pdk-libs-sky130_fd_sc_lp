* File: sky130_fd_sc_lp__a221oi_m.pex.spice
* Created: Fri Aug 28 09:53:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221OI_M%C1 3 5 9 13 15 16 17 22
c40 22 0 1.46778e-19 $X=0.535 $Y=1.615
r41 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.535
+ $Y=1.615 $X2=0.535 $Y2=1.615
r42 16 17 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.627 $Y=1.665
+ $X2=0.627 $Y2=2.035
r43 16 23 1.62316 $w=3.53e-07 $l=5e-08 $layer=LI1_cond $X=0.627 $Y=1.665
+ $X2=0.627 $Y2=1.615
r44 15 23 10.3882 $w=3.53e-07 $l=3.2e-07 $layer=LI1_cond $X=0.627 $Y=1.295
+ $X2=0.627 $Y2=1.615
r45 13 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.535 $Y=1.955
+ $X2=0.535 $Y2=1.615
r46 13 14 59.7919 $w=3.3e-07 $l=3.77425e-07 $layer=POLY_cond $X=0.535 $Y=1.955
+ $X2=0.55 $Y2=2.325
r47 12 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.45
+ $X2=0.535 $Y2=1.615
r48 7 9 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.975 $Y=2.4
+ $X2=0.975 $Y2=2.885
r49 6 14 11.3495 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.7 $Y=2.325 $X2=0.55
+ $Y2=2.325
r50 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.9 $Y=2.325
+ $X2=0.975 $Y2=2.4
r51 5 6 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=0.9 $Y=2.325 $X2=0.7
+ $Y2=2.325
r52 3 12 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=0.625 $Y=0.485
+ $X2=0.625 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_M%B2 3 7 9 16
c42 9 0 3.35074e-19 $X=1.2 $Y=1.665
c43 7 0 7.46275e-20 $X=1.405 $Y=2.885
r44 14 16 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.15 $Y=1.845
+ $X2=1.405 $Y2=1.845
r45 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.845 $X2=1.15 $Y2=1.845
r46 11 14 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.055 $Y=1.845
+ $X2=1.15 $Y2=1.845
r47 9 15 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.845
r48 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=2.01
+ $X2=1.405 $Y2=1.845
r49 5 7 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.405 $Y=2.01
+ $X2=1.405 $Y2=2.885
r50 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.68
+ $X2=1.055 $Y2=1.845
r51 1 3 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=1.055 $Y=1.68
+ $X2=1.055 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_M%B1 3 7 10 12 14 16 17 20 21 25 32
c66 21 0 6.62111e-20 $X=3.12 $Y=1.665
c67 7 0 7.46275e-20 $X=2.885 $Y=2.885
r68 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.975
+ $Y=1.54 $X2=2.975 $Y2=1.54
r69 21 26 3.40061 $w=5.08e-07 $l=1.45e-07 $layer=LI1_cond $X=3.12 $Y=1.71
+ $X2=2.975 $Y2=1.71
r70 20 26 7.85659 $w=5.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.64 $Y=1.71
+ $X2=2.975 $Y2=1.71
r71 20 32 6.08875 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.71
+ $X2=2.555 $Y2=1.71
r72 17 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.275
+ $X2=1.505 $Y2=1.11
r73 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.505
+ $Y=1.275 $X2=1.505 $Y2=1.275
r74 14 32 47.4378 $w=2.13e-07 $l=8.85e-07 $layer=LI1_cond $X=1.67 $Y=1.857
+ $X2=2.555 $Y2=1.857
r75 12 14 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=1.585 $Y=1.75
+ $X2=1.67 $Y2=1.857
r76 11 16 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.585 $Y=1.36
+ $X2=1.505 $Y2=1.275
r77 11 12 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.585 $Y=1.36
+ $X2=1.585 $Y2=1.75
r78 9 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.975 $Y=1.88
+ $X2=2.975 $Y2=1.54
r79 9 10 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.88
+ $X2=2.975 $Y2=2.045
r80 7 10 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.885 $Y=2.885
+ $X2=2.885 $Y2=2.045
r81 3 29 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.415 $Y=0.485
+ $X2=1.415 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_M%A1 3 7 10 13 15 18
c46 18 0 6.62111e-20 $X=2.045 $Y=1.36
c47 15 0 3.13702e-20 $X=2.16 $Y=1.295
c48 13 0 1.43233e-19 $X=1.955 $Y=1.755
r49 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.045 $Y=1.36
+ $X2=2.045 $Y2=1.525
r50 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.045 $Y=1.36
+ $X2=2.045 $Y2=1.195
r51 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.045
+ $Y=1.36 $X2=2.045 $Y2=1.36
r52 15 19 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.36
+ $X2=2.045 $Y2=1.36
r53 11 13 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.835 $Y=1.755
+ $X2=1.955 $Y2=1.755
r54 10 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.955 $Y=1.68
+ $X2=1.955 $Y2=1.755
r55 10 21 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.955 $Y=1.68
+ $X2=1.955 $Y2=1.525
r56 7 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.955 $Y=0.485
+ $X2=1.955 $Y2=1.195
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.835 $Y=1.83
+ $X2=1.835 $Y2=1.755
r58 1 3 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=1.835 $Y=1.83
+ $X2=1.835 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_M%A2 1 3 6 10 11 12 13 17
c44 17 0 4.63965e-20 $X=2.495 $Y=0.97
r45 17 19 16.3083 $w=2.66e-07 $l=9e-08 $layer=POLY_cond $X=2.495 $Y=0.97
+ $X2=2.585 $Y2=0.97
r46 12 13 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=2.585 $Y=0.97
+ $X2=3.12 $Y2=0.97
r47 12 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=0.97 $X2=2.585 $Y2=0.97
r48 10 11 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=2.475 $Y=1.765
+ $X2=2.475 $Y2=1.915
r49 8 17 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.135
+ $X2=2.495 $Y2=0.97
r50 8 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.495 $Y=1.135
+ $X2=2.495 $Y2=1.765
r51 6 11 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.455 $Y=2.885
+ $X2=2.455 $Y2=1.915
r52 1 17 32.6165 $w=2.66e-07 $l=2.49199e-07 $layer=POLY_cond $X=2.315 $Y=0.805
+ $X2=2.495 $Y2=0.97
r53 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.315 $Y=0.805
+ $X2=2.315 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_M%Y 1 2 3 10 12 14 15 16 17 18 19 26 39 46
c56 46 0 1.50262e-20 $X=1.63 $Y=0.57
c57 26 0 1.46778e-19 $X=1.465 $Y=0.877
r58 46 48 10.7212 $w=3.28e-07 $l=3.07e-07 $layer=LI1_cond $X=1.63 $Y=0.57
+ $X2=1.63 $Y2=0.877
r59 39 41 9.0807 $w=4.13e-07 $l=3.27e-07 $layer=LI1_cond $X=0.307 $Y=0.55
+ $X2=0.307 $Y2=0.877
r60 32 48 2.04284 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0.877
+ $X2=1.63 $Y2=0.877
r61 27 41 3.3765 $w=2.65e-07 $l=2.08e-07 $layer=LI1_cond $X=0.515 $Y=0.877
+ $X2=0.307 $Y2=0.877
r62 26 48 2.04284 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0.877
+ $X2=1.63 $Y2=0.877
r63 19 32 15.8733 $w=2.63e-07 $l=3.65e-07 $layer=LI1_cond $X=2.16 $Y=0.877
+ $X2=1.795 $Y2=0.877
r64 18 48 1.67628 $w=3.28e-07 $l=4.8e-08 $layer=LI1_cond $X=1.63 $Y=0.925
+ $X2=1.63 $Y2=0.877
r65 17 26 11.5244 $w=2.63e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=0.877
+ $X2=1.465 $Y2=0.877
r66 16 17 20.8744 $w=2.63e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=0.877
+ $X2=1.2 $Y2=0.877
r67 16 27 8.91512 $w=2.63e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=0.877
+ $X2=0.515 $Y2=0.877
r68 15 41 1.33295 $w=4.13e-07 $l=4.8e-08 $layer=LI1_cond $X=0.307 $Y=0.925
+ $X2=0.307 $Y2=0.877
r69 14 15 67.7415 $w=2.83e-07 $l=1.645e-06 $layer=LI1_cond $X=0.185 $Y=2.655
+ $X2=0.185 $Y2=1.01
r70 10 14 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.27 $Y=2.82
+ $X2=0.185 $Y2=2.655
r71 10 12 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.27 $Y=2.82 $X2=0.76
+ $Y2=2.82
r72 3 12 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=2.675 $X2=0.76 $Y2=2.82
r73 2 46 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.275 $X2=1.63 $Y2=0.57
r74 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.285
+ $Y=0.275 $X2=0.41 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_M%A_210_535# 1 2 9 11 12 15
r36 13 15 26.671 $w=2.08e-07 $l=5.05e-07 $layer=LI1_cond $X=3.1 $Y=2.315 $X2=3.1
+ $Y2=2.82
r37 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.995 $Y=2.23
+ $X2=3.1 $Y2=2.315
r38 11 12 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=2.995 $Y=2.23
+ $X2=1.295 $Y2=2.23
r39 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.19 $Y=2.315
+ $X2=1.295 $Y2=2.23
r40 7 9 26.671 $w=2.08e-07 $l=5.05e-07 $layer=LI1_cond $X=1.19 $Y=2.315 $X2=1.19
+ $Y2=2.82
r41 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=2.675 $X2=3.1 $Y2=2.82
r42 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=2.675 $X2=1.19 $Y2=2.82
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_M%A_296_535# 1 2 9 11 12 15
c24 15 0 2.19644e-19 $X=2.67 $Y=2.82
c25 9 0 2.19644e-19 $X=1.62 $Y=2.82
r26 13 15 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=2.67 $Y=2.665
+ $X2=2.67 $Y2=2.82
r27 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.565 $Y=2.58
+ $X2=2.67 $Y2=2.665
r28 11 12 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.565 $Y=2.58
+ $X2=1.725 $Y2=2.58
r29 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.62 $Y=2.665
+ $X2=1.725 $Y2=2.58
r30 7 9 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.62 $Y=2.665
+ $X2=1.62 $Y2=2.82
r31 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=2.675 $X2=2.67 $Y2=2.82
r32 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=2.675 $X2=1.62 $Y2=2.82
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_M%VPWR 1 6 8 10 20 21 24
r39 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=3.33
+ $X2=2.145 $Y2=3.33
r43 18 20 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.31 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=3.33
+ $X2=2.145 $Y2=3.33
r47 10 16 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.98 $Y=3.33 $X2=1.68
+ $Y2=3.33
r48 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 8 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=3.245
+ $X2=2.145 $Y2=3.33
r52 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.145 $Y=3.245
+ $X2=2.145 $Y2=2.95
r53 1 6 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=2.675 $X2=2.145 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_M%VGND 1 2 9 13 16 17 19 20 21 34 35
r35 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r36 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r37 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 28 31 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r39 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r40 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r41 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r43 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r44 19 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.16
+ $Y2=0
r45 19 20 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.53
+ $Y2=0
r46 18 34 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.635 $Y=0 $X2=3.12
+ $Y2=0
r47 18 20 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.635 $Y=0 $X2=2.53
+ $Y2=0
r48 16 24 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=0 $X2=0.72
+ $Y2=0
r49 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.735 $Y=0 $X2=0.84
+ $Y2=0
r50 15 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r51 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.84
+ $Y2=0
r52 11 20 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0
r53 11 13 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0.42
r54 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=0.085
+ $X2=0.84 $Y2=0
r55 7 9 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=0.84 $Y=0.085
+ $X2=0.84 $Y2=0.4
r56 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.275 $X2=2.53 $Y2=0.42
r57 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.7
+ $Y=0.275 $X2=0.84 $Y2=0.4
.ends

