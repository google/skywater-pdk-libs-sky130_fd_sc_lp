* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_778_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0206e+12p pd=9.18e+06u as=7.056e+11p ps=6.16e+06u
M1001 VGND A1 a_39_65# VNB nshort w=840000u l=150000u
+  ad=1.176e+12p pd=7.84e+06u as=1.5288e+12p ps=1.372e+07u
M1002 VGND A2 a_39_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_778_365# A2 a_519_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.0458e+12p ps=9.22e+06u
M1004 a_39_65# B2 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=5.376e+11p ps=4.64e+06u
M1005 a_39_367# B2 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0206e+12p pd=9.18e+06u as=7.056e+11p ps=6.16e+06u
M1006 Y B1 a_39_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_39_65# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_39_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_778_365# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_39_65# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_519_365# A3 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_39_65# B1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_39_65# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_519_365# A2 a_778_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B2 a_39_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B1 a_39_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A3 a_519_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A3 a_39_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B2 a_39_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
