* File: sky130_fd_sc_lp__sdfxbp_1.pxi.spice
* Created: Wed Sep  2 10:36:09 2020
* 
x_PM_SKY130_FD_SC_LP__SDFXBP_1%SCD N_SCD_M1017_g N_SCD_M1012_g N_SCD_c_273_n
+ N_SCD_c_277_n SCD SCD SCD N_SCD_c_275_n PM_SKY130_FD_SC_LP__SDFXBP_1%SCD
x_PM_SKY130_FD_SC_LP__SDFXBP_1%D N_D_M1000_g N_D_M1014_g N_D_c_299_n N_D_c_304_n
+ D D N_D_c_300_n N_D_c_301_n PM_SKY130_FD_SC_LP__SDFXBP_1%D
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_324_431# N_A_324_431#_M1003_d
+ N_A_324_431#_M1008_s N_A_324_431#_c_336_n N_A_324_431#_M1020_g
+ N_A_324_431#_M1001_g N_A_324_431#_c_338_n N_A_324_431#_c_333_n
+ N_A_324_431#_c_334_n N_A_324_431#_c_335_n
+ PM_SKY130_FD_SC_LP__SDFXBP_1%A_324_431#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%SCE N_SCE_M1031_g N_SCE_M1032_g N_SCE_c_389_n
+ N_SCE_c_390_n N_SCE_M1003_g N_SCE_c_392_n N_SCE_M1008_g N_SCE_c_394_n
+ N_SCE_c_395_n SCE SCE SCE N_SCE_c_396_n N_SCE_c_397_n
+ PM_SKY130_FD_SC_LP__SDFXBP_1%SCE
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_767_121# N_A_767_121#_M1005_s
+ N_A_767_121#_M1029_s N_A_767_121#_M1004_s N_A_767_121#_M1035_d
+ N_A_767_121#_M1023_g N_A_767_121#_M1021_g N_A_767_121#_c_469_n
+ N_A_767_121#_c_464_n N_A_767_121#_c_471_n N_A_767_121#_c_472_n
+ N_A_767_121#_c_473_n N_A_767_121#_c_474_n N_A_767_121#_c_475_n
+ N_A_767_121#_c_465_n N_A_767_121#_c_477_n N_A_767_121#_c_478_n
+ N_A_767_121#_c_466_n N_A_767_121#_c_480_n N_A_767_121#_c_467_n
+ N_A_767_121#_c_489_p PM_SKY130_FD_SC_LP__SDFXBP_1%A_767_121#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_1075_95# N_A_1075_95#_M1013_s
+ N_A_1075_95#_M1028_s N_A_1075_95#_M1018_g N_A_1075_95#_c_599_n
+ N_A_1075_95#_c_600_n N_A_1075_95#_M1010_g N_A_1075_95#_c_601_n
+ N_A_1075_95#_c_602_n N_A_1075_95#_M1002_g N_A_1075_95#_c_619_n
+ N_A_1075_95#_c_620_n N_A_1075_95#_M1029_g N_A_1075_95#_c_604_n
+ N_A_1075_95#_c_605_n N_A_1075_95#_c_606_n N_A_1075_95#_c_607_n
+ N_A_1075_95#_c_608_n N_A_1075_95#_c_609_n N_A_1075_95#_c_610_n
+ N_A_1075_95#_c_611_n N_A_1075_95#_c_646_p N_A_1075_95#_c_612_n
+ N_A_1075_95#_c_624_n N_A_1075_95#_c_625_n N_A_1075_95#_c_613_n
+ N_A_1075_95#_c_614_n PM_SKY130_FD_SC_LP__SDFXBP_1%A_1075_95#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_722_23# N_A_722_23#_M1018_d N_A_722_23#_M1010_d
+ N_A_722_23#_c_762_n N_A_722_23#_c_763_n N_A_722_23#_c_764_n
+ N_A_722_23#_c_765_n N_A_722_23#_c_766_n N_A_722_23#_c_775_n
+ N_A_722_23#_c_776_n N_A_722_23#_c_767_n N_A_722_23#_M1005_g
+ N_A_722_23#_c_777_n N_A_722_23#_M1004_g N_A_722_23#_c_778_n
+ N_A_722_23#_c_779_n N_A_722_23#_c_768_n N_A_722_23#_c_780_n
+ N_A_722_23#_c_781_n N_A_722_23#_c_782_n N_A_722_23#_c_769_n
+ N_A_722_23#_c_770_n N_A_722_23#_c_771_n N_A_722_23#_c_783_n
+ N_A_722_23#_c_772_n N_A_722_23#_c_773_n PM_SKY130_FD_SC_LP__SDFXBP_1%A_722_23#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_1161_95# N_A_1161_95#_M1033_d
+ N_A_1161_95#_M1016_d N_A_1161_95#_c_893_n N_A_1161_95#_M1019_g
+ N_A_1161_95#_c_894_n N_A_1161_95#_c_895_n N_A_1161_95#_c_911_n
+ N_A_1161_95#_M1027_g N_A_1161_95#_c_912_n N_A_1161_95#_c_913_n
+ N_A_1161_95#_c_896_n N_A_1161_95#_M1028_g N_A_1161_95#_c_897_n
+ N_A_1161_95#_M1013_g N_A_1161_95#_c_898_n N_A_1161_95#_c_899_n
+ N_A_1161_95#_M1035_g N_A_1161_95#_M1015_g N_A_1161_95#_c_902_n
+ N_A_1161_95#_c_903_n N_A_1161_95#_c_904_n N_A_1161_95#_c_905_n
+ N_A_1161_95#_c_906_n N_A_1161_95#_c_907_n N_A_1161_95#_c_908_n
+ N_A_1161_95#_c_909_n N_A_1161_95#_c_910_n
+ PM_SKY130_FD_SC_LP__SDFXBP_1%A_1161_95#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%CLK N_CLK_M1033_g N_CLK_M1016_g CLK CLK
+ N_CLK_c_1051_n N_CLK_c_1052_n PM_SKY130_FD_SC_LP__SDFXBP_1%CLK
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_2082_99# N_A_2082_99#_M1007_d
+ N_A_2082_99#_M1022_d N_A_2082_99#_M1011_g N_A_2082_99#_c_1100_n
+ N_A_2082_99#_M1006_g N_A_2082_99#_M1030_g N_A_2082_99#_M1034_g
+ N_A_2082_99#_c_1088_n N_A_2082_99#_M1024_g N_A_2082_99#_c_1090_n
+ N_A_2082_99#_M1025_g N_A_2082_99#_c_1092_n N_A_2082_99#_c_1093_n
+ N_A_2082_99#_c_1094_n N_A_2082_99#_c_1095_n N_A_2082_99#_c_1103_n
+ N_A_2082_99#_c_1096_n N_A_2082_99#_c_1104_n N_A_2082_99#_c_1105_n
+ N_A_2082_99#_c_1097_n N_A_2082_99#_c_1098_n N_A_2082_99#_c_1106_n
+ N_A_2082_99#_c_1107_n N_A_2082_99#_c_1108_n
+ PM_SKY130_FD_SC_LP__SDFXBP_1%A_2082_99#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_1873_497# N_A_1873_497#_M1029_d
+ N_A_1873_497#_M1002_d N_A_1873_497#_c_1211_n N_A_1873_497#_M1007_g
+ N_A_1873_497#_M1022_g N_A_1873_497#_c_1212_n N_A_1873_497#_c_1213_n
+ N_A_1873_497#_c_1214_n N_A_1873_497#_c_1215_n N_A_1873_497#_c_1216_n
+ N_A_1873_497#_c_1217_n PM_SKY130_FD_SC_LP__SDFXBP_1%A_1873_497#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_2409_367# N_A_2409_367#_M1030_d
+ N_A_2409_367#_M1034_s N_A_2409_367#_M1009_g N_A_2409_367#_M1026_g
+ N_A_2409_367#_c_1272_n N_A_2409_367#_c_1279_n N_A_2409_367#_c_1273_n
+ N_A_2409_367#_c_1274_n N_A_2409_367#_c_1282_n N_A_2409_367#_c_1275_n
+ N_A_2409_367#_c_1276_n PM_SKY130_FD_SC_LP__SDFXBP_1%A_2409_367#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_27_483# N_A_27_483#_M1017_s N_A_27_483#_M1020_d
+ N_A_27_483#_c_1337_n N_A_27_483#_c_1338_n N_A_27_483#_c_1339_n
+ N_A_27_483#_c_1340_n PM_SKY130_FD_SC_LP__SDFXBP_1%A_27_483#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%VPWR N_VPWR_M1017_d N_VPWR_M1008_d N_VPWR_M1004_d
+ N_VPWR_M1028_d N_VPWR_M1006_d N_VPWR_M1034_d N_VPWR_M1026_s N_VPWR_c_1366_n
+ N_VPWR_c_1367_n N_VPWR_c_1368_n N_VPWR_c_1369_n N_VPWR_c_1370_n
+ N_VPWR_c_1371_n N_VPWR_c_1372_n N_VPWR_c_1373_n N_VPWR_c_1374_n VPWR
+ N_VPWR_c_1375_n N_VPWR_c_1376_n N_VPWR_c_1377_n N_VPWR_c_1378_n
+ N_VPWR_c_1379_n N_VPWR_c_1380_n N_VPWR_c_1381_n N_VPWR_c_1365_n
+ N_VPWR_c_1383_n N_VPWR_c_1384_n N_VPWR_c_1385_n N_VPWR_c_1386_n
+ N_VPWR_c_1387_n N_VPWR_c_1388_n PM_SKY130_FD_SC_LP__SDFXBP_1%VPWR
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_196_119# N_A_196_119#_M1031_d
+ N_A_196_119#_M1019_d N_A_196_119#_M1000_d N_A_196_119#_M1010_s
+ N_A_196_119#_c_1558_n N_A_196_119#_c_1515_n N_A_196_119#_c_1501_n
+ N_A_196_119#_c_1502_n N_A_196_119#_c_1503_n N_A_196_119#_c_1504_n
+ N_A_196_119#_c_1517_n N_A_196_119#_c_1518_n N_A_196_119#_c_1550_n
+ N_A_196_119#_c_1505_n N_A_196_119#_c_1506_n N_A_196_119#_c_1521_n
+ N_A_196_119#_c_1507_n N_A_196_119#_c_1508_n N_A_196_119#_c_1509_n
+ N_A_196_119#_c_1510_n N_A_196_119#_c_1511_n N_A_196_119#_c_1512_n
+ N_A_196_119#_c_1513_n N_A_196_119#_c_1514_n N_A_196_119#_c_1522_n
+ N_A_196_119#_c_1556_n N_A_196_119#_c_1523_n
+ PM_SKY130_FD_SC_LP__SDFXBP_1%A_196_119#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_974_425# N_A_974_425#_M1023_d
+ N_A_974_425#_M1027_d N_A_974_425#_c_1671_n N_A_974_425#_c_1672_n
+ N_A_974_425#_c_1673_n PM_SKY130_FD_SC_LP__SDFXBP_1%A_974_425#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%A_1786_497# N_A_1786_497#_M1002_s
+ N_A_1786_497#_M1006_s N_A_1786_497#_c_1705_n N_A_1786_497#_c_1706_n
+ N_A_1786_497#_c_1707_n PM_SKY130_FD_SC_LP__SDFXBP_1%A_1786_497#
x_PM_SKY130_FD_SC_LP__SDFXBP_1%Q N_Q_M1025_s N_Q_M1024_d Q Q Q Q Q N_Q_c_1738_n
+ Q PM_SKY130_FD_SC_LP__SDFXBP_1%Q
x_PM_SKY130_FD_SC_LP__SDFXBP_1%Q_N N_Q_N_M1009_d N_Q_N_M1026_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1761_n Q_N PM_SKY130_FD_SC_LP__SDFXBP_1%Q_N
x_PM_SKY130_FD_SC_LP__SDFXBP_1%VGND N_VGND_M1012_s N_VGND_M1001_d N_VGND_M1005_d
+ N_VGND_M1013_d N_VGND_M1011_d N_VGND_M1030_s N_VGND_M1025_d N_VGND_c_1774_n
+ N_VGND_c_1775_n N_VGND_c_1776_n N_VGND_c_1777_n N_VGND_c_1778_n
+ N_VGND_c_1779_n N_VGND_c_1780_n N_VGND_c_1781_n N_VGND_c_1782_n
+ N_VGND_c_1783_n N_VGND_c_1784_n N_VGND_c_1785_n VGND N_VGND_c_1786_n
+ N_VGND_c_1787_n N_VGND_c_1788_n N_VGND_c_1789_n N_VGND_c_1790_n
+ N_VGND_c_1791_n N_VGND_c_1792_n N_VGND_c_1793_n N_VGND_c_1794_n
+ N_VGND_c_1795_n PM_SKY130_FD_SC_LP__SDFXBP_1%VGND
cc_1 VNB N_SCD_M1012_g 0.0264852f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.805
cc_2 VNB N_SCD_c_273_n 0.0241817f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.36
cc_3 VNB SCD 0.0261231f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_SCD_c_275_n 0.0244506f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_5 VNB N_D_M1014_g 0.0221287f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.805
cc_6 VNB N_D_c_299_n 0.0132531f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.36
cc_7 VNB N_D_c_300_n 0.0151883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_D_c_301_n 0.00420856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_324_431#_M1001_g 0.0441697f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.715
cc_10 VNB N_A_324_431#_c_333_n 0.0157647f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_11 VNB N_A_324_431#_c_334_n 0.0177499f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_12 VNB N_A_324_431#_c_335_n 0.00754543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_M1031_g 0.0590503f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_14 VNB N_SCE_c_389_n 0.0855006f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.805
cc_15 VNB N_SCE_c_390_n 0.0125466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_M1003_g 0.0341864f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.36
cc_17 VNB N_SCE_c_392_n 0.0616406f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.88
cc_18 VNB N_SCE_M1008_g 0.0448384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_SCE_c_394_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_SCE_c_395_n 0.0203751f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_21 VNB N_SCE_c_396_n 0.0437222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCE_c_397_n 0.00509066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_767_121#_M1021_g 0.0417574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_767_121#_c_464_n 0.0114408f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_25 VNB N_A_767_121#_c_465_n 0.0107953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_767_121#_c_466_n 0.0160457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_767_121#_c_467_n 0.0100955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_1075_95#_M1018_g 0.0349832f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.36
cc_29 VNB N_A_1075_95#_c_599_n 0.0136134f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.36
cc_30 VNB N_A_1075_95#_c_600_n 0.0042931f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.715
cc_31 VNB N_A_1075_95#_c_601_n 0.17277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1075_95#_c_602_n 0.0185818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1075_95#_M1029_g 0.0471508f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_34 VNB N_A_1075_95#_c_604_n 0.15681f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=2.035
cc_35 VNB N_A_1075_95#_c_605_n 0.0465425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1075_95#_c_606_n 0.0268449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1075_95#_c_607_n 0.0161011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1075_95#_c_608_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1075_95#_c_609_n 0.0197538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1075_95#_c_610_n 0.0182734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1075_95#_c_611_n 0.0266027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1075_95#_c_612_n 0.0492003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1075_95#_c_613_n 0.00245478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1075_95#_c_614_n 0.00711857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_722_23#_c_762_n 0.059023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_722_23#_c_763_n 0.00691438f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.21
cc_47 VNB N_A_722_23#_c_764_n 0.214744f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.36
cc_48 VNB N_A_722_23#_c_765_n 0.0101054f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.715
cc_49 VNB N_A_722_23#_c_766_n 0.0321906f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.88
cc_50 VNB N_A_722_23#_c_767_n 0.0175039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_722_23#_c_768_n 0.00573254f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_52 VNB N_A_722_23#_c_769_n 0.00259441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_722_23#_c_770_n 0.0106107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_722_23#_c_771_n 0.00277256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_722_23#_c_772_n 0.00528136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_722_23#_c_773_n 0.0498484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1161_95#_c_893_n 0.0163001f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.805
cc_58 VNB N_A_1161_95#_c_894_n 0.0876272f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.21
cc_59 VNB N_A_1161_95#_c_895_n 0.00811462f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.36
cc_60 VNB N_A_1161_95#_c_896_n 0.0493701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1161_95#_c_897_n 0.0167877f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_62 VNB N_A_1161_95#_c_898_n 0.00537378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1161_95#_c_899_n 0.066608f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.375
cc_64 VNB N_A_1161_95#_M1035_g 0.00580346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1161_95#_M1015_g 0.0244287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1161_95#_c_902_n 0.01179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1161_95#_c_903_n 0.0254627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1161_95#_c_904_n 0.00296467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1161_95#_c_905_n 2.13406e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1161_95#_c_906_n 0.0146687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1161_95#_c_907_n 0.00145246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1161_95#_c_908_n 0.0505094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1161_95#_c_909_n 0.00385815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1161_95#_c_910_n 0.00761318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_CLK_M1016_g 0.0115142f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.805
cc_76 VNB CLK 0.0138758f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.36
cc_77 VNB N_CLK_c_1051_n 0.0295461f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.88
cc_78 VNB N_CLK_c_1052_n 0.0197192f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_79 VNB N_A_2082_99#_M1011_g 0.043537f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.36
cc_80 VNB N_A_2082_99#_M1034_g 5.21609e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_2082_99#_c_1088_n 0.016519f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_82 VNB N_A_2082_99#_M1024_g 5.82935e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2082_99#_c_1090_n 0.0240957f $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.665
cc_84 VNB N_A_2082_99#_M1025_g 0.0283683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2082_99#_c_1092_n 0.0208497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2082_99#_c_1093_n 0.0265738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2082_99#_c_1094_n 0.00958052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_2082_99#_c_1095_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2082_99#_c_1096_n 0.0194754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2082_99#_c_1097_n 0.00732918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2082_99#_c_1098_n 0.017713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1873_497#_c_1211_n 0.018422f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=0.805
cc_93 VNB N_A_1873_497#_c_1212_n 3.51036e-19 $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_94 VNB N_A_1873_497#_c_1213_n 0.00349342f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.375
cc_95 VNB N_A_1873_497#_c_1214_n 0.00282467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1873_497#_c_1215_n 2.51413e-19 $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.375
cc_97 VNB N_A_1873_497#_c_1216_n 0.0258324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1873_497#_c_1217_n 0.0337753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2409_367#_c_1272_n 0.0124991f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_100 VNB N_A_2409_367#_c_1273_n 0.00160827f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.375
cc_101 VNB N_A_2409_367#_c_1274_n 0.0312135f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.375
cc_102 VNB N_A_2409_367#_c_1275_n 0.00507539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2409_367#_c_1276_n 0.0205096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VPWR_c_1365_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_196_119#_c_1501_n 0.00664753f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.375
cc_106 VNB N_A_196_119#_c_1502_n 0.00547379f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.375
cc_107 VNB N_A_196_119#_c_1503_n 0.0242866f $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.295
cc_108 VNB N_A_196_119#_c_1504_n 0.00584413f $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.375
cc_109 VNB N_A_196_119#_c_1505_n 0.00547978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_196_119#_c_1506_n 0.00161772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_196_119#_c_1507_n 0.0204705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_196_119#_c_1508_n 0.0140231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_196_119#_c_1509_n 0.00251271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_196_119#_c_1510_n 0.00308258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_196_119#_c_1511_n 0.0444081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_196_119#_c_1512_n 0.00139048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_196_119#_c_1513_n 0.0073263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_196_119#_c_1514_n 0.00350047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB Q 0.00326131f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.36
cc_120 VNB Q 7.51475e-19 $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.21
cc_121 VNB N_Q_c_1738_n 0.00349105f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_122 VNB Q_N 0.0104405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB Q_N 0.0247429f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.36
cc_124 VNB N_Q_N_c_1761_n 0.0295912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1774_n 0.0138117f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_126 VNB N_VGND_c_1775_n 0.0384833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1776_n 0.00831555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1777_n 0.0100707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1778_n 0.0144623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1779_n 0.0178466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1780_n 0.0175986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1781_n 0.0102151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1782_n 0.0603864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1783_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1784_n 0.0332097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1785_n 0.00423165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1786_n 0.0407217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1787_n 0.0731728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1788_n 0.0754218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1789_n 0.0273229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1790_n 0.021682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1791_n 0.709254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1792_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1793_n 0.00366215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_1794_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_1795_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VPB N_SCD_M1017_g 0.0496546f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_148 VPB N_SCD_c_277_n 0.0188601f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.88
cc_149 VPB SCD 0.0215958f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_150 VPB N_SCD_c_275_n 0.00490676f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.375
cc_151 VPB N_D_M1000_g 0.0319787f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_152 VPB N_D_c_299_n 0.00767936f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.36
cc_153 VPB N_D_c_304_n 0.0153271f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.715
cc_154 VPB N_D_c_301_n 0.00917861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_324_431#_c_336_n 0.0540529f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.805
cc_156 VPB N_A_324_431#_M1001_g 0.0175832f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.715
cc_157 VPB N_A_324_431#_c_338_n 0.0626168f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_158 VPB N_A_324_431#_c_333_n 0.00156716f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.375
cc_159 VPB N_A_324_431#_c_334_n 0.0401913f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.375
cc_160 VPB N_SCE_M1031_g 0.0477083f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_161 VPB N_SCE_M1008_g 0.052458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_767_121#_M1023_g 0.0225294f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_163 VPB N_A_767_121#_c_469_n 0.00828865f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.375
cc_164 VPB N_A_767_121#_c_464_n 6.37513e-19 $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.295
cc_165 VPB N_A_767_121#_c_471_n 0.00882594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_767_121#_c_472_n 0.0162211f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_167 VPB N_A_767_121#_c_473_n 0.00744447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_767_121#_c_474_n 0.020785f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_767_121#_c_475_n 0.00200453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_767_121#_c_465_n 0.0144701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_767_121#_c_477_n 0.00993333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_767_121#_c_478_n 0.00210403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_767_121#_c_466_n 0.0351342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_767_121#_c_480_n 0.00578528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_1075_95#_c_599_n 0.00892486f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.36
cc_176 VPB N_A_1075_95#_c_600_n 0.00361206f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.715
cc_177 VPB N_A_1075_95#_M1010_g 0.030506f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_178 VPB N_A_1075_95#_M1002_g 0.0243023f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.375
cc_179 VPB N_A_1075_95#_c_619_n 0.185562f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.295
cc_180 VPB N_A_1075_95#_c_620_n 0.0107582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_1075_95#_c_606_n 0.089282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_1075_95#_c_607_n 0.0486195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_1075_95#_c_611_n 0.0726898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1075_95#_c_624_n 0.00248965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1075_95#_c_625_n 0.00391765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_722_23#_c_763_n 0.0816797f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.21
cc_187 VPB N_A_722_23#_c_775_n 0.0288653f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_188 VPB N_A_722_23#_c_776_n 0.0109077f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_189 VPB N_A_722_23#_c_777_n 0.0182711f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.375
cc_190 VPB N_A_722_23#_c_778_n 0.0808106f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.295
cc_191 VPB N_A_722_23#_c_779_n 0.0502275f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.375
cc_192 VPB N_A_722_23#_c_780_n 0.00732516f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_722_23#_c_781_n 0.00523552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_722_23#_c_782_n 0.0390763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_722_23#_c_783_n 0.00150584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1161_95#_c_911_n 0.015207f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.715
cc_197 VPB N_A_1161_95#_c_912_n 0.172556f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_198 VPB N_A_1161_95#_c_913_n 0.0125761f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_199 VPB N_A_1161_95#_c_896_n 0.0153285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_1161_95#_M1028_g 0.0244787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1161_95#_c_898_n 0.0836289f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1161_95#_M1035_g 0.0262288f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1161_95#_c_905_n 0.00294881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1161_95#_c_909_n 0.00699708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1161_95#_c_910_n 0.00613109f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_CLK_M1016_g 0.0274605f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.805
cc_207 VPB N_A_2082_99#_M1011_g 0.00402881f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.36
cc_208 VPB N_A_2082_99#_c_1100_n 0.018985f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.36
cc_209 VPB N_A_2082_99#_M1034_g 0.0229807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_2082_99#_M1024_g 0.0255873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_2082_99#_c_1103_n 0.00707426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_2082_99#_c_1104_n 0.00286812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_2082_99#_c_1105_n 0.00966172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_2082_99#_c_1106_n 0.0531024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_2082_99#_c_1107_n 0.00195376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_2082_99#_c_1108_n 0.00163348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_1873_497#_M1022_g 0.0222137f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.715
cc_218 VPB N_A_1873_497#_c_1212_n 0.00625249f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_219 VPB N_A_1873_497#_c_1217_n 0.0122286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_2409_367#_M1026_g 0.0255204f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.715
cc_221 VPB N_A_2409_367#_c_1272_n 0.00296432f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.58
cc_222 VPB N_A_2409_367#_c_1279_n 0.0149578f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_223 VPB N_A_2409_367#_c_1273_n 0.00133664f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.375
cc_224 VPB N_A_2409_367#_c_1274_n 0.00825223f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.375
cc_225 VPB N_A_2409_367#_c_1282_n 0.0212099f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.665
cc_226 VPB N_A_27_483#_c_1337_n 0.024775f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.36
cc_227 VPB N_A_27_483#_c_1338_n 0.0175257f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.36
cc_228 VPB N_A_27_483#_c_1339_n 0.00968134f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.715
cc_229 VPB N_A_27_483#_c_1340_n 0.003999f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.88
cc_230 VPB N_VPWR_c_1366_n 0.00151893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1367_n 0.0104717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1368_n 0.00446584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1369_n 0.0195479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1370_n 0.0130584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1371_n 0.010112f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1372_n 0.010125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1373_n 0.0605717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1374_n 0.00497553f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1375_n 0.0156862f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1376_n 0.022597f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1377_n 0.0812985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1378_n 0.0740088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1379_n 0.0355228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1380_n 0.0206876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1381_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1365_n 0.0944548f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1383_n 0.00485691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1384_n 0.00436918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1385_n 0.00485691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1386_n 0.00470161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1387_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1388_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_196_119#_c_1515_n 0.010186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_196_119#_c_1504_n 0.021778f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.375
cc_255 VPB N_A_196_119#_c_1517_n 0.00836731f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.665
cc_256 VPB N_A_196_119#_c_1518_n 0.00410578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_196_119#_c_1505_n 0.00530549f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_196_119#_c_1506_n 4.50165e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_196_119#_c_1521_n 0.0154976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_196_119#_c_1522_n 0.00333346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_196_119#_c_1523_n 0.00615882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_974_425#_c_1671_n 0.0095312f $X=-0.19 $Y=1.655 $X2=0.545
+ $Y2=0.805
cc_263 VPB N_A_974_425#_c_1672_n 0.00853039f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.21
cc_264 VPB N_A_974_425#_c_1673_n 0.0137786f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_265 VPB N_A_1786_497#_c_1705_n 0.020389f $X=-0.19 $Y=1.655 $X2=0.545
+ $Y2=0.805
cc_266 VPB N_A_1786_497#_c_1706_n 0.0061233f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.36
cc_267 VPB N_A_1786_497#_c_1707_n 0.00599342f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_268 VPB Q 0.00820185f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.21
cc_269 VPB Q_N 0.0570134f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.36
cc_270 SCD N_D_c_301_n 0.0302161f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_271 N_SCD_M1012_g N_SCE_M1031_g 0.0540046f $X=0.545 $Y=0.805 $X2=0 $Y2=0
cc_272 SCD N_SCE_M1031_g 0.00392268f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_273 N_SCD_c_275_n N_SCE_M1031_g 0.0630827f $X=0.385 $Y=1.375 $X2=0 $Y2=0
cc_274 N_SCD_M1017_g N_A_27_483#_c_1337_n 2.21843e-19 $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_275 N_SCD_M1017_g N_A_27_483#_c_1338_n 0.0146898f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_276 SCD N_A_27_483#_c_1338_n 0.015113f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_277 N_SCD_c_277_n N_A_27_483#_c_1339_n 6.17585e-19 $X=0.385 $Y=1.88 $X2=0
+ $Y2=0
cc_278 SCD N_A_27_483#_c_1339_n 0.0243611f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_279 N_SCD_M1017_g N_VPWR_c_1366_n 0.0111979f $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_280 N_SCD_M1017_g N_VPWR_c_1375_n 0.00452967f $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_281 N_SCD_M1017_g N_VPWR_c_1365_n 0.0088676f $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_282 SCD N_A_196_119#_c_1502_n 0.00143134f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_283 N_SCD_M1012_g N_VGND_c_1775_n 0.0124072f $X=0.545 $Y=0.805 $X2=0 $Y2=0
cc_284 N_SCD_c_273_n N_VGND_c_1775_n 0.0014799f $X=0.42 $Y=1.36 $X2=0 $Y2=0
cc_285 SCD N_VGND_c_1775_n 0.0274351f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_286 N_SCD_M1012_g N_VGND_c_1786_n 0.0035863f $X=0.545 $Y=0.805 $X2=0 $Y2=0
cc_287 N_SCD_M1012_g N_VGND_c_1791_n 0.00401353f $X=0.545 $Y=0.805 $X2=0 $Y2=0
cc_288 N_D_M1000_g N_A_324_431#_c_336_n 0.0407348f $X=1.265 $Y=2.735 $X2=0 $Y2=0
cc_289 N_D_c_301_n N_A_324_431#_c_336_n 0.0044882f $X=1.355 $Y=1.44 $X2=0 $Y2=0
cc_290 N_D_M1014_g N_A_324_431#_M1001_g 0.0918449f $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_291 N_D_c_301_n N_A_324_431#_M1001_g 0.00358213f $X=1.355 $Y=1.44 $X2=0 $Y2=0
cc_292 N_D_M1014_g N_SCE_M1031_g 0.0135652f $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_293 N_D_c_300_n N_SCE_M1031_g 0.116971f $X=1.355 $Y=1.44 $X2=0 $Y2=0
cc_294 N_D_c_301_n N_SCE_M1031_g 0.00947552f $X=1.355 $Y=1.44 $X2=0 $Y2=0
cc_295 N_D_M1014_g N_SCE_c_389_n 0.0104164f $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_296 N_D_M1000_g N_A_27_483#_c_1338_n 0.0139413f $X=1.265 $Y=2.735 $X2=0 $Y2=0
cc_297 N_D_c_304_n N_A_27_483#_c_1338_n 8.18438e-19 $X=1.355 $Y=1.945 $X2=0
+ $Y2=0
cc_298 N_D_c_301_n N_A_27_483#_c_1338_n 0.0408179f $X=1.355 $Y=1.44 $X2=0 $Y2=0
cc_299 N_D_M1000_g N_A_27_483#_c_1340_n 0.00108109f $X=1.265 $Y=2.735 $X2=0
+ $Y2=0
cc_300 N_D_M1000_g N_VPWR_c_1366_n 0.00260283f $X=1.265 $Y=2.735 $X2=0 $Y2=0
cc_301 N_D_M1000_g N_VPWR_c_1373_n 0.00510276f $X=1.265 $Y=2.735 $X2=0 $Y2=0
cc_302 N_D_M1000_g N_VPWR_c_1365_n 0.00951251f $X=1.265 $Y=2.735 $X2=0 $Y2=0
cc_303 N_D_M1000_g N_A_196_119#_c_1515_n 0.00445221f $X=1.265 $Y=2.735 $X2=0
+ $Y2=0
cc_304 N_D_M1014_g N_A_196_119#_c_1501_n 0.0140681f $X=1.445 $Y=0.805 $X2=0
+ $Y2=0
cc_305 N_D_c_300_n N_A_196_119#_c_1501_n 8.42502e-19 $X=1.355 $Y=1.44 $X2=0
+ $Y2=0
cc_306 N_D_c_301_n N_A_196_119#_c_1501_n 0.0137096f $X=1.355 $Y=1.44 $X2=0 $Y2=0
cc_307 N_D_c_300_n N_A_196_119#_c_1502_n 0.00440573f $X=1.355 $Y=1.44 $X2=0
+ $Y2=0
cc_308 N_D_c_301_n N_A_196_119#_c_1502_n 0.0286793f $X=1.355 $Y=1.44 $X2=0 $Y2=0
cc_309 N_D_M1014_g N_A_196_119#_c_1514_n 0.00389063f $X=1.445 $Y=0.805 $X2=0
+ $Y2=0
cc_310 N_D_c_301_n N_A_196_119#_c_1514_n 0.00520378f $X=1.355 $Y=1.44 $X2=0
+ $Y2=0
cc_311 N_D_M1014_g N_VGND_c_1776_n 0.00142485f $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_312 N_D_M1014_g N_VGND_c_1791_n 9.39239e-19 $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_313 N_A_324_431#_M1001_g N_SCE_c_389_n 0.0103107f $X=1.805 $Y=0.805 $X2=0
+ $Y2=0
cc_314 N_A_324_431#_M1001_g N_SCE_M1003_g 0.0159474f $X=1.805 $Y=0.805 $X2=0
+ $Y2=0
cc_315 N_A_324_431#_c_333_n N_SCE_M1003_g 0.00498355f $X=2.69 $Y=1.74 $X2=0
+ $Y2=0
cc_316 N_A_324_431#_c_335_n N_SCE_c_392_n 0.00742666f $X=2.7 $Y=0.805 $X2=0
+ $Y2=0
cc_317 N_A_324_431#_c_333_n N_SCE_M1008_g 0.00859961f $X=2.69 $Y=1.74 $X2=0
+ $Y2=0
cc_318 N_A_324_431#_c_334_n N_SCE_M1008_g 0.0364548f $X=2.69 $Y=1.74 $X2=0 $Y2=0
cc_319 N_A_324_431#_c_335_n N_SCE_c_396_n 0.0033891f $X=2.7 $Y=0.805 $X2=0 $Y2=0
cc_320 N_A_324_431#_c_333_n N_SCE_c_397_n 0.0329901f $X=2.69 $Y=1.74 $X2=0 $Y2=0
cc_321 N_A_324_431#_c_335_n N_SCE_c_397_n 0.0262483f $X=2.7 $Y=0.805 $X2=0 $Y2=0
cc_322 N_A_324_431#_c_336_n N_A_27_483#_c_1338_n 0.0119515f $X=1.695 $Y=2.305
+ $X2=0 $Y2=0
cc_323 N_A_324_431#_c_336_n N_A_27_483#_c_1340_n 0.0187758f $X=1.695 $Y=2.305
+ $X2=0 $Y2=0
cc_324 N_A_324_431#_c_338_n N_A_27_483#_c_1340_n 0.0106449f $X=2.525 $Y=2.23
+ $X2=0 $Y2=0
cc_325 N_A_324_431#_c_336_n N_VPWR_c_1373_n 0.00333919f $X=1.695 $Y=2.305 $X2=0
+ $Y2=0
cc_326 N_A_324_431#_c_336_n N_VPWR_c_1365_n 0.00600122f $X=1.695 $Y=2.305 $X2=0
+ $Y2=0
cc_327 N_A_324_431#_c_336_n N_A_196_119#_c_1515_n 0.0139015f $X=1.695 $Y=2.305
+ $X2=0 $Y2=0
cc_328 N_A_324_431#_c_338_n N_A_196_119#_c_1515_n 0.0043959f $X=2.525 $Y=2.23
+ $X2=0 $Y2=0
cc_329 N_A_324_431#_M1001_g N_A_196_119#_c_1501_n 3.55637e-19 $X=1.805 $Y=0.805
+ $X2=0 $Y2=0
cc_330 N_A_324_431#_c_336_n N_A_196_119#_c_1503_n 0.00106626f $X=1.695 $Y=2.305
+ $X2=0 $Y2=0
cc_331 N_A_324_431#_M1001_g N_A_196_119#_c_1503_n 0.0062431f $X=1.805 $Y=0.805
+ $X2=0 $Y2=0
cc_332 N_A_324_431#_c_333_n N_A_196_119#_c_1503_n 0.0177039f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_333 N_A_324_431#_c_335_n N_A_196_119#_c_1503_n 0.00443936f $X=2.7 $Y=0.805
+ $X2=0 $Y2=0
cc_334 N_A_324_431#_c_336_n N_A_196_119#_c_1504_n 0.00791176f $X=1.695 $Y=2.305
+ $X2=0 $Y2=0
cc_335 N_A_324_431#_M1001_g N_A_196_119#_c_1504_n 0.0112833f $X=1.805 $Y=0.805
+ $X2=0 $Y2=0
cc_336 N_A_324_431#_c_338_n N_A_196_119#_c_1504_n 0.0184308f $X=2.525 $Y=2.23
+ $X2=0 $Y2=0
cc_337 N_A_324_431#_c_333_n N_A_196_119#_c_1504_n 0.096333f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_338 N_A_324_431#_c_334_n N_A_196_119#_c_1504_n 0.00668186f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_339 N_A_324_431#_M1008_s N_A_196_119#_c_1517_n 0.0103924f $X=2.585 $Y=2.405
+ $X2=0 $Y2=0
cc_340 N_A_324_431#_c_338_n N_A_196_119#_c_1517_n 0.00649349f $X=2.525 $Y=2.23
+ $X2=0 $Y2=0
cc_341 N_A_324_431#_c_333_n N_A_196_119#_c_1517_n 0.0158656f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_342 N_A_324_431#_c_333_n N_A_196_119#_c_1518_n 0.047779f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_343 N_A_324_431#_c_334_n N_A_196_119#_c_1518_n 0.00379866f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_344 N_A_324_431#_M1008_s N_A_196_119#_c_1550_n 0.00479176f $X=2.585 $Y=2.405
+ $X2=0 $Y2=0
cc_345 N_A_324_431#_c_333_n N_A_196_119#_c_1550_n 0.01251f $X=2.69 $Y=1.74 $X2=0
+ $Y2=0
cc_346 N_A_324_431#_c_333_n N_A_196_119#_c_1506_n 0.0137774f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_347 N_A_324_431#_c_334_n N_A_196_119#_c_1506_n 0.00111674f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_348 N_A_324_431#_c_333_n N_A_196_119#_c_1507_n 0.0054798f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_349 N_A_324_431#_M1001_g N_A_196_119#_c_1514_n 0.0237668f $X=1.805 $Y=0.805
+ $X2=0 $Y2=0
cc_350 N_A_324_431#_M1008_s N_A_196_119#_c_1556_n 0.00166402f $X=2.585 $Y=2.405
+ $X2=0 $Y2=0
cc_351 N_A_324_431#_c_333_n N_A_196_119#_c_1556_n 0.0140936f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_352 N_A_324_431#_M1001_g N_VGND_c_1776_n 0.00843572f $X=1.805 $Y=0.805 $X2=0
+ $Y2=0
cc_353 N_A_324_431#_c_335_n N_VGND_c_1782_n 0.00821888f $X=2.7 $Y=0.805 $X2=0
+ $Y2=0
cc_354 N_A_324_431#_M1001_g N_VGND_c_1791_n 7.88961e-19 $X=1.805 $Y=0.805 $X2=0
+ $Y2=0
cc_355 N_A_324_431#_c_335_n N_VGND_c_1791_n 0.01139f $X=2.7 $Y=0.805 $X2=0 $Y2=0
cc_356 N_SCE_M1008_g N_A_767_121#_c_464_n 2.0567e-19 $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_357 N_SCE_c_396_n N_A_722_23#_c_762_n 0.0217552f $X=3.09 $Y=0.43 $X2=0 $Y2=0
cc_358 N_SCE_c_397_n N_A_722_23#_c_762_n 4.26349e-19 $X=3.09 $Y=0.43 $X2=0 $Y2=0
cc_359 N_SCE_M1008_g N_A_722_23#_c_763_n 0.0217552f $X=3.18 $Y=2.725 $X2=0 $Y2=0
cc_360 N_SCE_c_392_n N_A_722_23#_c_765_n 0.0217552f $X=2.925 $Y=0.18 $X2=0 $Y2=0
cc_361 N_SCE_c_395_n N_A_722_23#_c_768_n 0.0217552f $X=3.09 $Y=0.935 $X2=0 $Y2=0
cc_362 N_SCE_M1031_g N_A_27_483#_c_1338_n 0.0183727f $X=0.905 $Y=0.805 $X2=0
+ $Y2=0
cc_363 N_SCE_M1031_g N_VPWR_c_1366_n 0.0132475f $X=0.905 $Y=0.805 $X2=0 $Y2=0
cc_364 N_SCE_M1008_g N_VPWR_c_1367_n 0.00363022f $X=3.18 $Y=2.725 $X2=0 $Y2=0
cc_365 N_SCE_M1031_g N_VPWR_c_1373_n 0.00452967f $X=0.905 $Y=0.805 $X2=0 $Y2=0
cc_366 N_SCE_M1008_g N_VPWR_c_1373_n 0.00480426f $X=3.18 $Y=2.725 $X2=0 $Y2=0
cc_367 N_SCE_M1031_g N_VPWR_c_1365_n 0.00803025f $X=0.905 $Y=0.805 $X2=0 $Y2=0
cc_368 N_SCE_M1008_g N_VPWR_c_1365_n 0.00649402f $X=3.18 $Y=2.725 $X2=0 $Y2=0
cc_369 N_SCE_c_389_n N_A_196_119#_c_1558_n 0.00494997f $X=2.16 $Y=0.18 $X2=0
+ $Y2=0
cc_370 N_SCE_M1031_g N_A_196_119#_c_1515_n 6.17816e-19 $X=0.905 $Y=0.805 $X2=0
+ $Y2=0
cc_371 N_SCE_M1031_g N_A_196_119#_c_1502_n 0.00480083f $X=0.905 $Y=0.805 $X2=0
+ $Y2=0
cc_372 N_SCE_M1003_g N_A_196_119#_c_1503_n 0.00716278f $X=2.235 $Y=0.805 $X2=0
+ $Y2=0
cc_373 N_SCE_M1008_g N_A_196_119#_c_1504_n 8.4406e-19 $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_374 N_SCE_M1008_g N_A_196_119#_c_1517_n 0.00634426f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_375 N_SCE_M1008_g N_A_196_119#_c_1518_n 0.0182094f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_376 N_SCE_M1008_g N_A_196_119#_c_1550_n 0.0108942f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_377 N_SCE_M1008_g N_A_196_119#_c_1505_n 0.0095487f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_378 N_SCE_c_397_n N_A_196_119#_c_1505_n 0.00522204f $X=3.09 $Y=0.43 $X2=0
+ $Y2=0
cc_379 N_SCE_M1008_g N_A_196_119#_c_1506_n 0.00243228f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_380 N_SCE_c_395_n N_A_196_119#_c_1506_n 4.07083e-19 $X=3.09 $Y=0.935 $X2=0
+ $Y2=0
cc_381 N_SCE_c_397_n N_A_196_119#_c_1506_n 0.015473f $X=3.09 $Y=0.43 $X2=0 $Y2=0
cc_382 N_SCE_M1008_g N_A_196_119#_c_1521_n 0.0095342f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_383 N_SCE_c_396_n N_A_196_119#_c_1507_n 0.00886248f $X=3.09 $Y=0.43 $X2=0
+ $Y2=0
cc_384 N_SCE_c_397_n N_A_196_119#_c_1507_n 0.0699547f $X=3.09 $Y=0.43 $X2=0
+ $Y2=0
cc_385 N_SCE_c_396_n N_A_196_119#_c_1509_n 0.00146874f $X=3.09 $Y=0.43 $X2=0
+ $Y2=0
cc_386 N_SCE_c_397_n N_A_196_119#_c_1509_n 0.0140305f $X=3.09 $Y=0.43 $X2=0
+ $Y2=0
cc_387 N_SCE_M1003_g N_A_196_119#_c_1514_n 8.66828e-19 $X=2.235 $Y=0.805 $X2=0
+ $Y2=0
cc_388 N_SCE_M1008_g N_A_196_119#_c_1522_n 3.2832e-19 $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_389 N_SCE_M1008_g N_A_196_119#_c_1556_n 0.00351786f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_390 N_SCE_M1031_g N_VGND_c_1775_n 0.00180362f $X=0.905 $Y=0.805 $X2=0 $Y2=0
cc_391 N_SCE_c_390_n N_VGND_c_1775_n 0.0101515f $X=0.98 $Y=0.18 $X2=0 $Y2=0
cc_392 N_SCE_c_389_n N_VGND_c_1776_n 0.0182317f $X=2.16 $Y=0.18 $X2=0 $Y2=0
cc_393 N_SCE_M1003_g N_VGND_c_1776_n 0.0249022f $X=2.235 $Y=0.805 $X2=0 $Y2=0
cc_394 N_SCE_c_394_n N_VGND_c_1776_n 0.00460513f $X=2.235 $Y=0.18 $X2=0 $Y2=0
cc_395 N_SCE_c_394_n N_VGND_c_1782_n 0.0317094f $X=2.235 $Y=0.18 $X2=0 $Y2=0
cc_396 N_SCE_c_397_n N_VGND_c_1782_n 0.0152228f $X=3.09 $Y=0.43 $X2=0 $Y2=0
cc_397 N_SCE_c_390_n N_VGND_c_1786_n 0.0335445f $X=0.98 $Y=0.18 $X2=0 $Y2=0
cc_398 N_SCE_c_389_n N_VGND_c_1791_n 0.0326485f $X=2.16 $Y=0.18 $X2=0 $Y2=0
cc_399 N_SCE_c_390_n N_VGND_c_1791_n 0.0116041f $X=0.98 $Y=0.18 $X2=0 $Y2=0
cc_400 N_SCE_c_392_n N_VGND_c_1791_n 0.0347351f $X=2.925 $Y=0.18 $X2=0 $Y2=0
cc_401 N_SCE_c_394_n N_VGND_c_1791_n 0.00749832f $X=2.235 $Y=0.18 $X2=0 $Y2=0
cc_402 N_SCE_c_397_n N_VGND_c_1791_n 0.00811271f $X=3.09 $Y=0.43 $X2=0 $Y2=0
cc_403 N_A_767_121#_c_474_n N_A_1075_95#_M1028_s 0.00514762f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_404 N_A_767_121#_M1021_g N_A_1075_95#_M1018_g 0.0380545f $X=5.09 $Y=0.815
+ $X2=0 $Y2=0
cc_405 N_A_767_121#_c_472_n N_A_1075_95#_c_600_n 0.007886f $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_406 N_A_767_121#_c_466_n N_A_1075_95#_c_600_n 0.0380545f $X=4.885 $Y=1.77
+ $X2=0 $Y2=0
cc_407 N_A_767_121#_c_473_n N_A_1075_95#_M1010_g 6.6777e-19 $X=6.65 $Y=2.345
+ $X2=0 $Y2=0
cc_408 N_A_767_121#_c_467_n N_A_1075_95#_c_601_n 0.00796081f $X=9.48 $Y=0.835
+ $X2=0 $Y2=0
cc_409 N_A_767_121#_c_477_n N_A_1075_95#_M1002_g 0.0075087f $X=10.02 $Y=2.43
+ $X2=0 $Y2=0
cc_410 N_A_767_121#_c_489_p N_A_1075_95#_M1002_g 0.0044856f $X=9.17 $Y=2.43
+ $X2=0 $Y2=0
cc_411 N_A_767_121#_c_465_n N_A_1075_95#_M1029_g 0.00136687f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_412 N_A_767_121#_c_472_n N_A_1075_95#_c_607_n 0.0247508f $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_413 N_A_767_121#_c_472_n N_A_1075_95#_c_610_n 0.0133403f $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_414 N_A_767_121#_c_473_n N_A_1075_95#_c_610_n 0.00833792f $X=6.65 $Y=2.345
+ $X2=0 $Y2=0
cc_415 N_A_767_121#_c_472_n N_A_1075_95#_c_611_n 0.016548f $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_416 N_A_767_121#_c_473_n N_A_1075_95#_c_611_n 0.0217807f $X=6.65 $Y=2.345
+ $X2=0 $Y2=0
cc_417 N_A_767_121#_c_474_n N_A_1075_95#_c_611_n 0.00868563f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_418 N_A_767_121#_c_473_n N_A_1075_95#_c_624_n 0.0144733f $X=6.65 $Y=2.345
+ $X2=0 $Y2=0
cc_419 N_A_767_121#_c_474_n N_A_1075_95#_c_624_n 0.0198939f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_420 N_A_767_121#_c_474_n N_A_1075_95#_c_625_n 0.0292389f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_421 N_A_767_121#_c_464_n N_A_722_23#_c_762_n 0.00640311f $X=3.98 $Y=0.78
+ $X2=0 $Y2=0
cc_422 N_A_767_121#_c_469_n N_A_722_23#_c_763_n 0.0137939f $X=3.93 $Y=1.685
+ $X2=0 $Y2=0
cc_423 N_A_767_121#_c_464_n N_A_722_23#_c_763_n 0.00215263f $X=3.98 $Y=0.78
+ $X2=0 $Y2=0
cc_424 N_A_767_121#_M1021_g N_A_722_23#_c_764_n 0.0104353f $X=5.09 $Y=0.815
+ $X2=0 $Y2=0
cc_425 N_A_767_121#_c_464_n N_A_722_23#_c_766_n 0.0182748f $X=3.98 $Y=0.78 $X2=0
+ $Y2=0
cc_426 N_A_767_121#_c_471_n N_A_722_23#_c_766_n 0.00730549f $X=4.785 $Y=1.95
+ $X2=0 $Y2=0
cc_427 N_A_767_121#_c_464_n N_A_722_23#_c_767_n 0.00214601f $X=3.98 $Y=0.78
+ $X2=0 $Y2=0
cc_428 N_A_767_121#_M1023_g N_A_722_23#_c_777_n 0.0222249f $X=4.795 $Y=2.335
+ $X2=0 $Y2=0
cc_429 N_A_767_121#_c_471_n N_A_722_23#_c_777_n 0.0143299f $X=4.785 $Y=1.95
+ $X2=0 $Y2=0
cc_430 N_A_767_121#_M1023_g N_A_722_23#_c_778_n 0.00456925f $X=4.795 $Y=2.335
+ $X2=0 $Y2=0
cc_431 N_A_767_121#_c_472_n N_A_722_23#_c_781_n 0.0734513f $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_432 N_A_767_121#_c_473_n N_A_722_23#_c_781_n 0.0142392f $X=6.65 $Y=2.345
+ $X2=0 $Y2=0
cc_433 N_A_767_121#_c_480_n N_A_722_23#_c_781_n 0.00979869f $X=5.05 $Y=1.95
+ $X2=0 $Y2=0
cc_434 N_A_767_121#_M1023_g N_A_722_23#_c_782_n 0.0179462f $X=4.795 $Y=2.335
+ $X2=0 $Y2=0
cc_435 N_A_767_121#_c_472_n N_A_722_23#_c_782_n 0.00377378f $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_436 N_A_767_121#_c_480_n N_A_722_23#_c_782_n 0.00370573f $X=5.05 $Y=1.95
+ $X2=0 $Y2=0
cc_437 N_A_767_121#_M1021_g N_A_722_23#_c_769_n 0.00147723f $X=5.09 $Y=0.815
+ $X2=0 $Y2=0
cc_438 N_A_767_121#_c_473_n N_A_722_23#_c_783_n 0.00982387f $X=6.65 $Y=2.345
+ $X2=0 $Y2=0
cc_439 N_A_767_121#_c_475_n N_A_722_23#_c_783_n 0.0133632f $X=6.735 $Y=2.43
+ $X2=0 $Y2=0
cc_440 N_A_767_121#_c_474_n N_A_1161_95#_M1016_d 0.00444638f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_441 N_A_767_121#_c_472_n N_A_1161_95#_c_894_n 0.00253857f $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_442 N_A_767_121#_c_472_n N_A_1161_95#_c_911_n 5.33412e-19 $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_443 N_A_767_121#_c_475_n N_A_1161_95#_c_911_n 0.00320944f $X=6.735 $Y=2.43
+ $X2=0 $Y2=0
cc_444 N_A_767_121#_c_474_n N_A_1161_95#_c_912_n 0.0259161f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_445 N_A_767_121#_c_475_n N_A_1161_95#_c_912_n 5.18472e-19 $X=6.735 $Y=2.43
+ $X2=0 $Y2=0
cc_446 N_A_767_121#_c_474_n N_A_1161_95#_M1028_g 0.0140973f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_447 N_A_767_121#_c_474_n N_A_1161_95#_c_898_n 0.012717f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_448 N_A_767_121#_c_465_n N_A_1161_95#_c_898_n 0.00915956f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_449 N_A_767_121#_c_465_n N_A_1161_95#_c_899_n 0.0149561f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_450 N_A_767_121#_c_467_n N_A_1161_95#_c_899_n 0.00907382f $X=9.48 $Y=0.835
+ $X2=0 $Y2=0
cc_451 N_A_767_121#_c_465_n N_A_1161_95#_M1035_g 0.00468757f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_452 N_A_767_121#_c_477_n N_A_1161_95#_M1035_g 0.0132994f $X=10.02 $Y=2.43
+ $X2=0 $Y2=0
cc_453 N_A_767_121#_c_478_n N_A_1161_95#_c_903_n 0.00110116f $X=10.125 $Y=2.04
+ $X2=0 $Y2=0
cc_454 N_A_767_121#_c_474_n N_A_1161_95#_c_905_n 5.78535e-19 $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_455 N_A_767_121#_c_467_n N_A_1161_95#_c_906_n 0.0247864f $X=9.48 $Y=0.835
+ $X2=0 $Y2=0
cc_456 N_A_767_121#_c_465_n N_A_1161_95#_c_907_n 0.0452704f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_457 N_A_767_121#_c_467_n N_A_1161_95#_c_907_n 0.00428086f $X=9.48 $Y=0.835
+ $X2=0 $Y2=0
cc_458 N_A_767_121#_c_465_n N_A_1161_95#_c_908_n 0.00785067f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_459 N_A_767_121#_c_467_n N_A_1161_95#_c_908_n 0.00127742f $X=9.48 $Y=0.835
+ $X2=0 $Y2=0
cc_460 N_A_767_121#_c_474_n N_A_1161_95#_c_909_n 0.0180439f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_461 N_A_767_121#_c_474_n N_A_1161_95#_c_910_n 0.042292f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_462 N_A_767_121#_c_465_n N_A_1161_95#_c_910_n 0.0459271f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_463 N_A_767_121#_c_474_n N_CLK_M1016_g 0.0124284f $X=9.085 $Y=2.43 $X2=0
+ $Y2=0
cc_464 N_A_767_121#_c_478_n N_A_2082_99#_c_1100_n 0.00320565f $X=10.125 $Y=2.04
+ $X2=0 $Y2=0
cc_465 N_A_767_121#_c_478_n N_A_2082_99#_c_1106_n 0.00333917f $X=10.125 $Y=2.04
+ $X2=0 $Y2=0
cc_466 N_A_767_121#_c_478_n N_A_2082_99#_c_1107_n 0.00792506f $X=10.125 $Y=2.04
+ $X2=0 $Y2=0
cc_467 N_A_767_121#_c_477_n N_A_1873_497#_M1002_d 0.00675231f $X=10.02 $Y=2.43
+ $X2=0 $Y2=0
cc_468 N_A_767_121#_c_465_n N_A_1873_497#_c_1212_n 0.0317569f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_469 N_A_767_121#_c_477_n N_A_1873_497#_c_1212_n 0.0220026f $X=10.02 $Y=2.43
+ $X2=0 $Y2=0
cc_470 N_A_767_121#_c_478_n N_A_1873_497#_c_1212_n 0.0119949f $X=10.125 $Y=2.04
+ $X2=0 $Y2=0
cc_471 N_A_767_121#_c_465_n N_A_1873_497#_c_1213_n 0.015973f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_472 N_A_767_121#_c_465_n N_A_1873_497#_c_1214_n 0.00923121f $X=9.17 $Y=2.345
+ $X2=0 $Y2=0
cc_473 N_A_767_121#_c_478_n N_A_1873_497#_c_1214_n 0.00305742f $X=10.125 $Y=2.04
+ $X2=0 $Y2=0
cc_474 N_A_767_121#_c_467_n N_A_1873_497#_c_1214_n 0.00151885f $X=9.48 $Y=0.835
+ $X2=0 $Y2=0
cc_475 N_A_767_121#_c_478_n N_A_1873_497#_c_1216_n 0.0102608f $X=10.125 $Y=2.04
+ $X2=0 $Y2=0
cc_476 N_A_767_121#_c_471_n N_VPWR_M1004_d 0.00295406f $X=4.785 $Y=1.95 $X2=0
+ $Y2=0
cc_477 N_A_767_121#_c_474_n N_VPWR_M1028_d 0.00978495f $X=9.085 $Y=2.43 $X2=0
+ $Y2=0
cc_478 N_A_767_121#_c_474_n N_VPWR_c_1369_n 0.0254559f $X=9.085 $Y=2.43 $X2=0
+ $Y2=0
cc_479 N_A_767_121#_M1023_g N_VPWR_c_1365_n 9.73184e-19 $X=4.795 $Y=2.335 $X2=0
+ $Y2=0
cc_480 N_A_767_121#_c_474_n N_VPWR_c_1365_n 0.0534381f $X=9.085 $Y=2.43 $X2=0
+ $Y2=0
cc_481 N_A_767_121#_c_475_n N_VPWR_c_1365_n 3.36104e-19 $X=6.735 $Y=2.43 $X2=0
+ $Y2=0
cc_482 N_A_767_121#_c_469_n N_A_196_119#_c_1518_n 0.0140399f $X=3.93 $Y=1.685
+ $X2=0 $Y2=0
cc_483 N_A_767_121#_c_469_n N_A_196_119#_c_1505_n 0.00326221f $X=3.93 $Y=1.685
+ $X2=0 $Y2=0
cc_484 N_A_767_121#_c_464_n N_A_196_119#_c_1505_n 0.0084081f $X=3.98 $Y=0.78
+ $X2=0 $Y2=0
cc_485 N_A_767_121#_M1004_s N_A_196_119#_c_1521_n 0.00681899f $X=3.835 $Y=1.975
+ $X2=0 $Y2=0
cc_486 N_A_767_121#_M1023_g N_A_196_119#_c_1521_n 0.0110012f $X=4.795 $Y=2.335
+ $X2=0 $Y2=0
cc_487 N_A_767_121#_c_469_n N_A_196_119#_c_1521_n 0.0220442f $X=3.93 $Y=1.685
+ $X2=0 $Y2=0
cc_488 N_A_767_121#_c_471_n N_A_196_119#_c_1521_n 0.0584519f $X=4.785 $Y=1.95
+ $X2=0 $Y2=0
cc_489 N_A_767_121#_c_472_n N_A_196_119#_c_1521_n 0.0111591f $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_490 N_A_767_121#_c_466_n N_A_196_119#_c_1521_n 0.00110549f $X=4.885 $Y=1.77
+ $X2=0 $Y2=0
cc_491 N_A_767_121#_c_464_n N_A_196_119#_c_1507_n 0.0572543f $X=3.98 $Y=0.78
+ $X2=0 $Y2=0
cc_492 N_A_767_121#_c_464_n N_A_196_119#_c_1508_n 0.0198509f $X=3.98 $Y=0.78
+ $X2=0 $Y2=0
cc_493 N_A_767_121#_M1021_g N_A_196_119#_c_1510_n 0.00436128f $X=5.09 $Y=0.815
+ $X2=0 $Y2=0
cc_494 N_A_767_121#_c_464_n N_A_196_119#_c_1510_n 0.0279592f $X=3.98 $Y=0.78
+ $X2=0 $Y2=0
cc_495 N_A_767_121#_M1021_g N_A_196_119#_c_1511_n 0.0166739f $X=5.09 $Y=0.815
+ $X2=0 $Y2=0
cc_496 N_A_767_121#_c_471_n N_A_196_119#_c_1511_n 0.113866f $X=4.785 $Y=1.95
+ $X2=0 $Y2=0
cc_497 N_A_767_121#_c_472_n N_A_196_119#_c_1511_n 0.0176162f $X=6.565 $Y=1.77
+ $X2=0 $Y2=0
cc_498 N_A_767_121#_c_466_n N_A_196_119#_c_1511_n 0.00833538f $X=4.885 $Y=1.77
+ $X2=0 $Y2=0
cc_499 N_A_767_121#_c_464_n N_A_196_119#_c_1512_n 0.0134135f $X=3.98 $Y=0.78
+ $X2=0 $Y2=0
cc_500 N_A_767_121#_c_471_n N_A_196_119#_c_1512_n 0.0147867f $X=4.785 $Y=1.95
+ $X2=0 $Y2=0
cc_501 N_A_767_121#_c_480_n N_A_974_425#_M1023_d 0.00244319f $X=5.05 $Y=1.95
+ $X2=-0.19 $Y2=-0.245
cc_502 N_A_767_121#_c_474_n N_A_974_425#_M1027_d 0.00117312f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_503 N_A_767_121#_c_475_n N_A_974_425#_M1027_d 0.00176768f $X=6.735 $Y=2.43
+ $X2=0 $Y2=0
cc_504 N_A_767_121#_c_474_n N_A_974_425#_c_1673_n 0.0121102f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_505 N_A_767_121#_c_475_n N_A_974_425#_c_1673_n 0.0141193f $X=6.735 $Y=2.43
+ $X2=0 $Y2=0
cc_506 N_A_767_121#_c_474_n N_A_1786_497#_M1002_s 0.00161549f $X=9.085 $Y=2.43
+ $X2=-0.19 $Y2=-0.245
cc_507 N_A_767_121#_c_489_p N_A_1786_497#_M1002_s 7.97188e-19 $X=9.17 $Y=2.43
+ $X2=-0.19 $Y2=-0.245
cc_508 N_A_767_121#_M1035_d N_A_1786_497#_c_1705_n 0.00254685f $X=9.985 $Y=1.895
+ $X2=0 $Y2=0
cc_509 N_A_767_121#_c_477_n N_A_1786_497#_c_1705_n 0.0517263f $X=10.02 $Y=2.43
+ $X2=0 $Y2=0
cc_510 N_A_767_121#_c_489_p N_A_1786_497#_c_1705_n 9.01554e-19 $X=9.17 $Y=2.43
+ $X2=0 $Y2=0
cc_511 N_A_767_121#_c_477_n N_A_1786_497#_c_1706_n 0.0139779f $X=10.02 $Y=2.43
+ $X2=0 $Y2=0
cc_512 N_A_767_121#_c_478_n N_A_1786_497#_c_1706_n 0.00615079f $X=10.125 $Y=2.04
+ $X2=0 $Y2=0
cc_513 N_A_767_121#_c_474_n N_A_1786_497#_c_1707_n 0.012801f $X=9.085 $Y=2.43
+ $X2=0 $Y2=0
cc_514 N_A_767_121#_c_489_p N_A_1786_497#_c_1707_n 0.00780602f $X=9.17 $Y=2.43
+ $X2=0 $Y2=0
cc_515 N_A_767_121#_M1021_g N_VGND_c_1777_n 0.0207078f $X=5.09 $Y=0.815 $X2=0
+ $Y2=0
cc_516 N_A_767_121#_c_467_n N_VGND_c_1788_n 0.00842906f $X=9.48 $Y=0.835 $X2=0
+ $Y2=0
cc_517 N_A_767_121#_M1021_g N_VGND_c_1791_n 9.27138e-19 $X=5.09 $Y=0.815 $X2=0
+ $Y2=0
cc_518 N_A_767_121#_c_467_n N_VGND_c_1791_n 0.0120887f $X=9.48 $Y=0.835 $X2=0
+ $Y2=0
cc_519 N_A_1075_95#_M1018_g N_A_722_23#_c_764_n 0.0103221f $X=5.45 $Y=0.815
+ $X2=0 $Y2=0
cc_520 N_A_1075_95#_c_602_n N_A_722_23#_c_764_n 0.020224f $X=7.28 $Y=0.18 $X2=0
+ $Y2=0
cc_521 N_A_1075_95#_c_646_p N_A_722_23#_c_764_n 2.28803e-19 $X=7.115 $Y=0.35
+ $X2=0 $Y2=0
cc_522 N_A_1075_95#_M1010_g N_A_722_23#_c_779_n 0.0181902f $X=6.005 $Y=2.715
+ $X2=0 $Y2=0
cc_523 N_A_1075_95#_M1010_g N_A_722_23#_c_781_n 0.00765135f $X=6.005 $Y=2.715
+ $X2=0 $Y2=0
cc_524 N_A_1075_95#_c_607_n N_A_722_23#_c_781_n 0.0224753f $X=6.415 $Y=1.83
+ $X2=0 $Y2=0
cc_525 N_A_1075_95#_c_600_n N_A_722_23#_c_782_n 0.0138299f $X=5.525 $Y=1.6 $X2=0
+ $Y2=0
cc_526 N_A_1075_95#_c_607_n N_A_722_23#_c_782_n 0.0225216f $X=6.415 $Y=1.83
+ $X2=0 $Y2=0
cc_527 N_A_1075_95#_M1018_g N_A_722_23#_c_769_n 0.0112892f $X=5.45 $Y=0.815
+ $X2=0 $Y2=0
cc_528 N_A_1075_95#_M1010_g N_A_722_23#_c_783_n 0.0119183f $X=6.005 $Y=2.715
+ $X2=0 $Y2=0
cc_529 N_A_1075_95#_c_646_p N_A_722_23#_c_772_n 0.0210298f $X=7.115 $Y=0.35
+ $X2=0 $Y2=0
cc_530 N_A_1075_95#_c_612_n N_A_722_23#_c_772_n 0.00160003f $X=7.115 $Y=0.35
+ $X2=0 $Y2=0
cc_531 N_A_1075_95#_c_614_n N_A_722_23#_c_772_n 0.0182583f $X=7.092 $Y=0.78
+ $X2=0 $Y2=0
cc_532 N_A_1075_95#_c_646_p N_A_722_23#_c_773_n 6.62023e-19 $X=7.115 $Y=0.35
+ $X2=0 $Y2=0
cc_533 N_A_1075_95#_c_612_n N_A_722_23#_c_773_n 0.020224f $X=7.115 $Y=0.35 $X2=0
+ $Y2=0
cc_534 N_A_1075_95#_c_614_n N_A_722_23#_c_773_n 0.00158695f $X=7.092 $Y=0.78
+ $X2=0 $Y2=0
cc_535 N_A_1075_95#_M1018_g N_A_1161_95#_c_893_n 0.0194169f $X=5.45 $Y=0.815
+ $X2=0 $Y2=0
cc_536 N_A_1075_95#_c_607_n N_A_1161_95#_c_894_n 0.0811446f $X=6.415 $Y=1.83
+ $X2=0 $Y2=0
cc_537 N_A_1075_95#_c_610_n N_A_1161_95#_c_894_n 0.0188557f $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_538 N_A_1075_95#_c_612_n N_A_1161_95#_c_894_n 0.0151757f $X=7.115 $Y=0.35
+ $X2=0 $Y2=0
cc_539 N_A_1075_95#_c_625_n N_A_1161_95#_c_894_n 0.00485686f $X=7.47 $Y=2.08
+ $X2=0 $Y2=0
cc_540 N_A_1075_95#_c_613_n N_A_1161_95#_c_894_n 0.0045017f $X=7.515 $Y=0.78
+ $X2=0 $Y2=0
cc_541 N_A_1075_95#_c_614_n N_A_1161_95#_c_894_n 0.00305495f $X=7.092 $Y=0.78
+ $X2=0 $Y2=0
cc_542 N_A_1075_95#_c_599_n N_A_1161_95#_c_895_n 0.00712379f $X=5.93 $Y=1.6
+ $X2=0 $Y2=0
cc_543 N_A_1075_95#_M1010_g N_A_1161_95#_c_911_n 0.0162864f $X=6.005 $Y=2.715
+ $X2=0 $Y2=0
cc_544 N_A_1075_95#_c_607_n N_A_1161_95#_c_911_n 0.0115285f $X=6.415 $Y=1.83
+ $X2=0 $Y2=0
cc_545 N_A_1075_95#_c_620_n N_A_1161_95#_c_912_n 0.0118762f $X=9.365 $Y=3.15
+ $X2=0 $Y2=0
cc_546 N_A_1075_95#_c_610_n N_A_1161_95#_c_896_n 0.00563203f $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_547 N_A_1075_95#_c_611_n N_A_1161_95#_c_896_n 0.0168162f $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_548 N_A_1075_95#_c_625_n N_A_1161_95#_c_896_n 0.00129042f $X=7.47 $Y=2.08
+ $X2=0 $Y2=0
cc_549 N_A_1075_95#_c_613_n N_A_1161_95#_c_896_n 0.00156316f $X=7.515 $Y=0.78
+ $X2=0 $Y2=0
cc_550 N_A_1075_95#_c_610_n N_A_1161_95#_M1028_g 9.37869e-19 $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_551 N_A_1075_95#_c_611_n N_A_1161_95#_M1028_g 0.00778849f $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_552 N_A_1075_95#_c_625_n N_A_1161_95#_M1028_g 0.00486957f $X=7.47 $Y=2.08
+ $X2=0 $Y2=0
cc_553 N_A_1075_95#_c_601_n N_A_1161_95#_c_897_n 0.0104164f $X=9.62 $Y=0.18
+ $X2=0 $Y2=0
cc_554 N_A_1075_95#_c_610_n N_A_1161_95#_c_897_n 0.00417183f $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_555 N_A_1075_95#_c_646_p N_A_1161_95#_c_897_n 5.10414e-19 $X=7.115 $Y=0.35
+ $X2=0 $Y2=0
cc_556 N_A_1075_95#_c_612_n N_A_1161_95#_c_897_n 0.00801451f $X=7.115 $Y=0.35
+ $X2=0 $Y2=0
cc_557 N_A_1075_95#_M1002_g N_A_1161_95#_c_898_n 0.0118762f $X=9.29 $Y=2.695
+ $X2=0 $Y2=0
cc_558 N_A_1075_95#_M1029_g N_A_1161_95#_c_899_n 0.00874073f $X=9.695 $Y=0.835
+ $X2=0 $Y2=0
cc_559 N_A_1075_95#_M1002_g N_A_1161_95#_M1035_g 0.0127273f $X=9.29 $Y=2.695
+ $X2=0 $Y2=0
cc_560 N_A_1075_95#_c_619_n N_A_1161_95#_M1035_g 0.00886347f $X=11.82 $Y=3.15
+ $X2=0 $Y2=0
cc_561 N_A_1075_95#_M1029_g N_A_1161_95#_M1015_g 0.0163664f $X=9.695 $Y=0.835
+ $X2=0 $Y2=0
cc_562 N_A_1075_95#_c_604_n N_A_1161_95#_M1015_g 0.00899284f $X=11.7 $Y=0.18
+ $X2=0 $Y2=0
cc_563 N_A_1075_95#_c_610_n N_A_1161_95#_c_904_n 0.0282538f $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_564 N_A_1075_95#_c_611_n N_A_1161_95#_c_904_n 5.5547e-19 $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_565 N_A_1075_95#_c_613_n N_A_1161_95#_c_904_n 0.0166011f $X=7.515 $Y=0.78
+ $X2=0 $Y2=0
cc_566 N_A_1075_95#_c_610_n N_A_1161_95#_c_905_n 0.0101131f $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_567 N_A_1075_95#_c_611_n N_A_1161_95#_c_905_n 7.2548e-19 $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_568 N_A_1075_95#_c_625_n N_A_1161_95#_c_905_n 0.0152844f $X=7.47 $Y=2.08
+ $X2=0 $Y2=0
cc_569 N_A_1075_95#_c_601_n N_A_1161_95#_c_906_n 0.0101058f $X=9.62 $Y=0.18
+ $X2=0 $Y2=0
cc_570 N_A_1075_95#_c_601_n N_A_1161_95#_c_908_n 0.00492978f $X=9.62 $Y=0.18
+ $X2=0 $Y2=0
cc_571 N_A_1075_95#_M1029_g N_A_1161_95#_c_908_n 0.0023854f $X=9.695 $Y=0.835
+ $X2=0 $Y2=0
cc_572 N_A_1075_95#_c_625_n N_CLK_M1016_g 8.44954e-19 $X=7.47 $Y=2.08 $X2=0
+ $Y2=0
cc_573 N_A_1075_95#_c_601_n N_CLK_c_1052_n 0.0104164f $X=9.62 $Y=0.18 $X2=0
+ $Y2=0
cc_574 N_A_1075_95#_c_604_n N_A_2082_99#_M1011_g 0.00907339f $X=11.7 $Y=0.18
+ $X2=0 $Y2=0
cc_575 N_A_1075_95#_c_619_n N_A_2082_99#_c_1100_n 0.00646075f $X=11.82 $Y=3.15
+ $X2=0 $Y2=0
cc_576 N_A_1075_95#_c_606_n N_A_2082_99#_M1034_g 0.0195948f $X=11.895 $Y=3.075
+ $X2=0 $Y2=0
cc_577 N_A_1075_95#_c_605_n N_A_2082_99#_c_1092_n 0.00924313f $X=11.775 $Y=0.94
+ $X2=0 $Y2=0
cc_578 N_A_1075_95#_c_609_n N_A_2082_99#_c_1092_n 0.00138657f $X=11.895 $Y=1.015
+ $X2=0 $Y2=0
cc_579 N_A_1075_95#_c_606_n N_A_2082_99#_c_1093_n 0.0183461f $X=11.895 $Y=3.075
+ $X2=0 $Y2=0
cc_580 N_A_1075_95#_c_604_n N_A_2082_99#_c_1096_n 0.00857044f $X=11.7 $Y=0.18
+ $X2=0 $Y2=0
cc_581 N_A_1075_95#_c_605_n N_A_2082_99#_c_1096_n 0.00888262f $X=11.775 $Y=0.94
+ $X2=0 $Y2=0
cc_582 N_A_1075_95#_c_609_n N_A_2082_99#_c_1096_n 0.00951405f $X=11.895 $Y=1.015
+ $X2=0 $Y2=0
cc_583 N_A_1075_95#_c_606_n N_A_2082_99#_c_1104_n 0.00443353f $X=11.895 $Y=3.075
+ $X2=0 $Y2=0
cc_584 N_A_1075_95#_c_619_n N_A_2082_99#_c_1105_n 0.00455019f $X=11.82 $Y=3.15
+ $X2=0 $Y2=0
cc_585 N_A_1075_95#_c_606_n N_A_2082_99#_c_1105_n 0.012253f $X=11.895 $Y=3.075
+ $X2=0 $Y2=0
cc_586 N_A_1075_95#_c_606_n N_A_2082_99#_c_1097_n 0.0298663f $X=11.895 $Y=3.075
+ $X2=0 $Y2=0
cc_587 N_A_1075_95#_c_609_n N_A_2082_99#_c_1097_n 0.0124531f $X=11.895 $Y=1.015
+ $X2=0 $Y2=0
cc_588 N_A_1075_95#_c_609_n N_A_2082_99#_c_1098_n 0.0183461f $X=11.895 $Y=1.015
+ $X2=0 $Y2=0
cc_589 N_A_1075_95#_c_606_n N_A_2082_99#_c_1108_n 0.00204323f $X=11.895 $Y=3.075
+ $X2=0 $Y2=0
cc_590 N_A_1075_95#_c_604_n N_A_1873_497#_c_1211_n 0.00905501f $X=11.7 $Y=0.18
+ $X2=0 $Y2=0
cc_591 N_A_1075_95#_c_605_n N_A_1873_497#_c_1211_n 0.00581219f $X=11.775 $Y=0.94
+ $X2=0 $Y2=0
cc_592 N_A_1075_95#_c_606_n N_A_1873_497#_c_1211_n 0.00212002f $X=11.895
+ $Y=3.075 $X2=0 $Y2=0
cc_593 N_A_1075_95#_c_619_n N_A_1873_497#_M1022_g 0.0103107f $X=11.82 $Y=3.15
+ $X2=0 $Y2=0
cc_594 N_A_1075_95#_M1029_g N_A_1873_497#_c_1213_n 0.00781692f $X=9.695 $Y=0.835
+ $X2=0 $Y2=0
cc_595 N_A_1075_95#_c_604_n N_A_1873_497#_c_1213_n 0.0044536f $X=11.7 $Y=0.18
+ $X2=0 $Y2=0
cc_596 N_A_1075_95#_M1029_g N_A_1873_497#_c_1214_n 8.77705e-19 $X=9.695 $Y=0.835
+ $X2=0 $Y2=0
cc_597 N_A_1075_95#_c_606_n N_A_1873_497#_c_1217_n 0.0310914f $X=11.895 $Y=3.075
+ $X2=0 $Y2=0
cc_598 N_A_1075_95#_c_606_n N_A_2409_367#_c_1282_n 0.00697666f $X=11.895
+ $Y=3.075 $X2=0 $Y2=0
cc_599 N_A_1075_95#_c_619_n N_VPWR_c_1370_n 0.0271239f $X=11.82 $Y=3.15 $X2=0
+ $Y2=0
cc_600 N_A_1075_95#_c_606_n N_VPWR_c_1370_n 0.00629238f $X=11.895 $Y=3.075 $X2=0
+ $Y2=0
cc_601 N_A_1075_95#_c_606_n N_VPWR_c_1371_n 0.0126056f $X=11.895 $Y=3.075 $X2=0
+ $Y2=0
cc_602 N_A_1075_95#_M1010_g N_VPWR_c_1377_n 9.29198e-19 $X=6.005 $Y=2.715 $X2=0
+ $Y2=0
cc_603 N_A_1075_95#_c_620_n N_VPWR_c_1378_n 0.0416934f $X=9.365 $Y=3.15 $X2=0
+ $Y2=0
cc_604 N_A_1075_95#_c_619_n N_VPWR_c_1379_n 0.0201276f $X=11.82 $Y=3.15 $X2=0
+ $Y2=0
cc_605 N_A_1075_95#_c_619_n N_VPWR_c_1365_n 0.068374f $X=11.82 $Y=3.15 $X2=0
+ $Y2=0
cc_606 N_A_1075_95#_c_620_n N_VPWR_c_1365_n 0.00525952f $X=9.365 $Y=3.15 $X2=0
+ $Y2=0
cc_607 N_A_1075_95#_M1018_g N_A_196_119#_c_1511_n 0.0152693f $X=5.45 $Y=0.815
+ $X2=0 $Y2=0
cc_608 N_A_1075_95#_c_599_n N_A_196_119#_c_1511_n 0.00762725f $X=5.93 $Y=1.6
+ $X2=0 $Y2=0
cc_609 N_A_1075_95#_c_607_n N_A_196_119#_c_1511_n 0.00487031f $X=6.415 $Y=1.83
+ $X2=0 $Y2=0
cc_610 N_A_1075_95#_M1018_g N_A_196_119#_c_1513_n 0.00201325f $X=5.45 $Y=0.815
+ $X2=0 $Y2=0
cc_611 N_A_1075_95#_M1010_g N_A_196_119#_c_1523_n 0.00250845f $X=6.005 $Y=2.715
+ $X2=0 $Y2=0
cc_612 N_A_1075_95#_M1010_g N_A_974_425#_c_1671_n 0.0146842f $X=6.005 $Y=2.715
+ $X2=0 $Y2=0
cc_613 N_A_1075_95#_c_611_n N_A_974_425#_c_1673_n 8.31485e-19 $X=7 $Y=1.66 $X2=0
+ $Y2=0
cc_614 N_A_1075_95#_M1002_g N_A_1786_497#_c_1705_n 0.0104796f $X=9.29 $Y=2.695
+ $X2=0 $Y2=0
cc_615 N_A_1075_95#_c_619_n N_A_1786_497#_c_1705_n 0.0274679f $X=11.82 $Y=3.15
+ $X2=0 $Y2=0
cc_616 N_A_1075_95#_M1002_g N_A_1786_497#_c_1707_n 0.00247782f $X=9.29 $Y=2.695
+ $X2=0 $Y2=0
cc_617 N_A_1075_95#_c_601_n N_VGND_c_1778_n 0.0229587f $X=9.62 $Y=0.18 $X2=0
+ $Y2=0
cc_618 N_A_1075_95#_c_646_p N_VGND_c_1778_n 0.0119608f $X=7.115 $Y=0.35 $X2=0
+ $Y2=0
cc_619 N_A_1075_95#_c_612_n N_VGND_c_1778_n 0.00407101f $X=7.115 $Y=0.35 $X2=0
+ $Y2=0
cc_620 N_A_1075_95#_c_604_n N_VGND_c_1779_n 0.0260628f $X=11.7 $Y=0.18 $X2=0
+ $Y2=0
cc_621 N_A_1075_95#_c_605_n N_VGND_c_1779_n 0.00567278f $X=11.775 $Y=0.94 $X2=0
+ $Y2=0
cc_622 N_A_1075_95#_c_604_n N_VGND_c_1780_n 0.0166171f $X=11.7 $Y=0.18 $X2=0
+ $Y2=0
cc_623 N_A_1075_95#_c_602_n N_VGND_c_1787_n 0.0228632f $X=7.28 $Y=0.18 $X2=0
+ $Y2=0
cc_624 N_A_1075_95#_c_646_p N_VGND_c_1787_n 0.0223688f $X=7.115 $Y=0.35 $X2=0
+ $Y2=0
cc_625 N_A_1075_95#_c_613_n N_VGND_c_1787_n 0.00653584f $X=7.515 $Y=0.78 $X2=0
+ $Y2=0
cc_626 N_A_1075_95#_c_614_n N_VGND_c_1787_n 9.50445e-19 $X=7.092 $Y=0.78 $X2=0
+ $Y2=0
cc_627 N_A_1075_95#_c_601_n N_VGND_c_1788_n 0.0806179f $X=9.62 $Y=0.18 $X2=0
+ $Y2=0
cc_628 N_A_1075_95#_c_604_n N_VGND_c_1789_n 0.0249021f $X=11.7 $Y=0.18 $X2=0
+ $Y2=0
cc_629 N_A_1075_95#_M1018_g N_VGND_c_1791_n 7.7504e-19 $X=5.45 $Y=0.815 $X2=0
+ $Y2=0
cc_630 N_A_1075_95#_c_601_n N_VGND_c_1791_n 0.064007f $X=9.62 $Y=0.18 $X2=0
+ $Y2=0
cc_631 N_A_1075_95#_c_602_n N_VGND_c_1791_n 0.00903939f $X=7.28 $Y=0.18 $X2=0
+ $Y2=0
cc_632 N_A_1075_95#_c_604_n N_VGND_c_1791_n 0.0675119f $X=11.7 $Y=0.18 $X2=0
+ $Y2=0
cc_633 N_A_1075_95#_c_608_n N_VGND_c_1791_n 0.0085374f $X=9.695 $Y=0.18 $X2=0
+ $Y2=0
cc_634 N_A_1075_95#_c_646_p N_VGND_c_1791_n 0.0112528f $X=7.115 $Y=0.35 $X2=0
+ $Y2=0
cc_635 N_A_1075_95#_c_613_n N_VGND_c_1791_n 0.009153f $X=7.515 $Y=0.78 $X2=0
+ $Y2=0
cc_636 N_A_1075_95#_c_614_n N_VGND_c_1791_n 0.00138582f $X=7.092 $Y=0.78 $X2=0
+ $Y2=0
cc_637 N_A_722_23#_c_764_n N_A_1161_95#_c_893_n 0.00976298f $X=6.38 $Y=0.19
+ $X2=0 $Y2=0
cc_638 N_A_722_23#_c_769_n N_A_1161_95#_c_893_n 0.00194566f $X=5.665 $Y=0.815
+ $X2=0 $Y2=0
cc_639 N_A_722_23#_c_770_n N_A_1161_95#_c_893_n 0.0037576f $X=6.38 $Y=0.345
+ $X2=0 $Y2=0
cc_640 N_A_722_23#_c_772_n N_A_1161_95#_c_893_n 6.38665e-19 $X=6.545 $Y=0.35
+ $X2=0 $Y2=0
cc_641 N_A_722_23#_c_773_n N_A_1161_95#_c_893_n 0.00640003f $X=6.545 $Y=0.35
+ $X2=0 $Y2=0
cc_642 N_A_722_23#_c_772_n N_A_1161_95#_c_894_n 0.00204259f $X=6.545 $Y=0.35
+ $X2=0 $Y2=0
cc_643 N_A_722_23#_c_773_n N_A_1161_95#_c_894_n 0.0138504f $X=6.545 $Y=0.35
+ $X2=0 $Y2=0
cc_644 N_A_722_23#_c_783_n N_A_1161_95#_c_911_n 0.0113948f $X=6.22 $Y=2.63 $X2=0
+ $Y2=0
cc_645 N_A_722_23#_c_763_n N_VPWR_c_1367_n 0.0142425f $X=3.685 $Y=3.075 $X2=0
+ $Y2=0
cc_646 N_A_722_23#_c_763_n N_VPWR_c_1368_n 0.00117707f $X=3.685 $Y=3.075 $X2=0
+ $Y2=0
cc_647 N_A_722_23#_c_777_n N_VPWR_c_1368_n 0.0117333f $X=4.27 $Y=3.075 $X2=0
+ $Y2=0
cc_648 N_A_722_23#_c_778_n N_VPWR_c_1368_n 0.0180829f $X=5.34 $Y=3.15 $X2=0
+ $Y2=0
cc_649 N_A_722_23#_c_779_n N_VPWR_c_1368_n 2.18997e-19 $X=5.415 $Y=3.075 $X2=0
+ $Y2=0
cc_650 N_A_722_23#_c_780_n N_VPWR_c_1368_n 0.00460513f $X=4.27 $Y=3.15 $X2=0
+ $Y2=0
cc_651 N_A_722_23#_c_776_n N_VPWR_c_1376_n 0.0266976f $X=3.76 $Y=3.15 $X2=0
+ $Y2=0
cc_652 N_A_722_23#_c_778_n N_VPWR_c_1377_n 0.0222665f $X=5.34 $Y=3.15 $X2=0
+ $Y2=0
cc_653 N_A_722_23#_c_775_n N_VPWR_c_1365_n 0.0128304f $X=4.195 $Y=3.15 $X2=0
+ $Y2=0
cc_654 N_A_722_23#_c_776_n N_VPWR_c_1365_n 0.0060156f $X=3.76 $Y=3.15 $X2=0
+ $Y2=0
cc_655 N_A_722_23#_c_778_n N_VPWR_c_1365_n 0.0235189f $X=5.34 $Y=3.15 $X2=0
+ $Y2=0
cc_656 N_A_722_23#_c_780_n N_VPWR_c_1365_n 0.00362613f $X=4.27 $Y=3.15 $X2=0
+ $Y2=0
cc_657 N_A_722_23#_c_763_n N_A_196_119#_c_1518_n 0.00238952f $X=3.685 $Y=3.075
+ $X2=0 $Y2=0
cc_658 N_A_722_23#_c_763_n N_A_196_119#_c_1550_n 8.68806e-19 $X=3.685 $Y=3.075
+ $X2=0 $Y2=0
cc_659 N_A_722_23#_c_763_n N_A_196_119#_c_1505_n 0.00181197f $X=3.685 $Y=3.075
+ $X2=0 $Y2=0
cc_660 N_A_722_23#_c_763_n N_A_196_119#_c_1521_n 0.0174657f $X=3.685 $Y=3.075
+ $X2=0 $Y2=0
cc_661 N_A_722_23#_c_775_n N_A_196_119#_c_1521_n 0.00605291f $X=4.195 $Y=3.15
+ $X2=0 $Y2=0
cc_662 N_A_722_23#_c_777_n N_A_196_119#_c_1521_n 0.0127764f $X=4.27 $Y=3.075
+ $X2=0 $Y2=0
cc_663 N_A_722_23#_c_778_n N_A_196_119#_c_1521_n 0.00515367f $X=5.34 $Y=3.15
+ $X2=0 $Y2=0
cc_664 N_A_722_23#_c_779_n N_A_196_119#_c_1521_n 0.0120133f $X=5.415 $Y=3.075
+ $X2=0 $Y2=0
cc_665 N_A_722_23#_c_781_n N_A_196_119#_c_1521_n 0.0108022f $X=6.055 $Y=2.12
+ $X2=0 $Y2=0
cc_666 N_A_722_23#_c_782_n N_A_196_119#_c_1521_n 0.00133948f $X=5.555 $Y=2.12
+ $X2=0 $Y2=0
cc_667 N_A_722_23#_c_762_n N_A_196_119#_c_1507_n 0.0135221f $X=3.685 $Y=1.355
+ $X2=0 $Y2=0
cc_668 N_A_722_23#_c_762_n N_A_196_119#_c_1508_n 0.0139907f $X=3.685 $Y=1.355
+ $X2=0 $Y2=0
cc_669 N_A_722_23#_c_764_n N_A_196_119#_c_1508_n 0.0108395f $X=6.38 $Y=0.19
+ $X2=0 $Y2=0
cc_670 N_A_722_23#_c_767_n N_A_196_119#_c_1508_n 0.00283033f $X=4.195 $Y=1.355
+ $X2=0 $Y2=0
cc_671 N_A_722_23#_c_762_n N_A_196_119#_c_1510_n 0.00181273f $X=3.685 $Y=1.355
+ $X2=0 $Y2=0
cc_672 N_A_722_23#_c_767_n N_A_196_119#_c_1510_n 0.0255334f $X=4.195 $Y=1.355
+ $X2=0 $Y2=0
cc_673 N_A_722_23#_c_769_n N_A_196_119#_c_1511_n 0.0114123f $X=5.665 $Y=0.815
+ $X2=0 $Y2=0
cc_674 N_A_722_23#_c_766_n N_A_196_119#_c_1512_n 0.00643356f $X=4.12 $Y=1.43
+ $X2=0 $Y2=0
cc_675 N_A_722_23#_c_767_n N_A_196_119#_c_1512_n 6.75682e-19 $X=4.195 $Y=1.355
+ $X2=0 $Y2=0
cc_676 N_A_722_23#_c_777_n N_A_196_119#_c_1512_n 3.32747e-19 $X=4.27 $Y=3.075
+ $X2=0 $Y2=0
cc_677 N_A_722_23#_c_764_n N_A_196_119#_c_1513_n 0.0011448f $X=6.38 $Y=0.19
+ $X2=0 $Y2=0
cc_678 N_A_722_23#_c_770_n N_A_196_119#_c_1513_n 0.0134624f $X=6.38 $Y=0.345
+ $X2=0 $Y2=0
cc_679 N_A_722_23#_c_772_n N_A_196_119#_c_1513_n 0.0148369f $X=6.545 $Y=0.35
+ $X2=0 $Y2=0
cc_680 N_A_722_23#_c_773_n N_A_196_119#_c_1513_n 0.00165671f $X=6.545 $Y=0.35
+ $X2=0 $Y2=0
cc_681 N_A_722_23#_c_779_n N_A_196_119#_c_1523_n 0.00546122f $X=5.415 $Y=3.075
+ $X2=0 $Y2=0
cc_682 N_A_722_23#_c_781_n N_A_196_119#_c_1523_n 0.0257321f $X=6.055 $Y=2.12
+ $X2=0 $Y2=0
cc_683 N_A_722_23#_c_782_n N_A_196_119#_c_1523_n 0.00431683f $X=5.555 $Y=2.12
+ $X2=0 $Y2=0
cc_684 N_A_722_23#_c_783_n N_A_196_119#_c_1523_n 0.0169412f $X=6.22 $Y=2.63
+ $X2=0 $Y2=0
cc_685 N_A_722_23#_M1010_d N_A_974_425#_c_1671_n 0.00176461f $X=6.08 $Y=2.505
+ $X2=0 $Y2=0
cc_686 N_A_722_23#_c_779_n N_A_974_425#_c_1671_n 0.0121427f $X=5.415 $Y=3.075
+ $X2=0 $Y2=0
cc_687 N_A_722_23#_c_782_n N_A_974_425#_c_1671_n 2.99023e-19 $X=5.555 $Y=2.12
+ $X2=0 $Y2=0
cc_688 N_A_722_23#_c_783_n N_A_974_425#_c_1671_n 0.0160508f $X=6.22 $Y=2.63
+ $X2=0 $Y2=0
cc_689 N_A_722_23#_c_777_n N_A_974_425#_c_1672_n 8.5977e-19 $X=4.27 $Y=3.075
+ $X2=0 $Y2=0
cc_690 N_A_722_23#_c_778_n N_A_974_425#_c_1672_n 0.00739395f $X=5.34 $Y=3.15
+ $X2=0 $Y2=0
cc_691 N_A_722_23#_c_779_n N_A_974_425#_c_1672_n 0.00841291f $X=5.415 $Y=3.075
+ $X2=0 $Y2=0
cc_692 N_A_722_23#_c_764_n N_VGND_c_1777_n 0.0265021f $X=6.38 $Y=0.19 $X2=0
+ $Y2=0
cc_693 N_A_722_23#_c_767_n N_VGND_c_1777_n 0.00371944f $X=4.195 $Y=1.355 $X2=0
+ $Y2=0
cc_694 N_A_722_23#_c_769_n N_VGND_c_1777_n 0.0160574f $X=5.665 $Y=0.815 $X2=0
+ $Y2=0
cc_695 N_A_722_23#_c_771_n N_VGND_c_1777_n 0.00656011f $X=5.795 $Y=0.345 $X2=0
+ $Y2=0
cc_696 N_A_722_23#_c_765_n N_VGND_c_1782_n 0.0225456f $X=3.76 $Y=0.19 $X2=0
+ $Y2=0
cc_697 N_A_722_23#_c_764_n N_VGND_c_1787_n 0.0460284f $X=6.38 $Y=0.19 $X2=0
+ $Y2=0
cc_698 N_A_722_23#_c_770_n N_VGND_c_1787_n 0.0360645f $X=6.38 $Y=0.345 $X2=0
+ $Y2=0
cc_699 N_A_722_23#_c_771_n N_VGND_c_1787_n 0.0201108f $X=5.795 $Y=0.345 $X2=0
+ $Y2=0
cc_700 N_A_722_23#_c_772_n N_VGND_c_1787_n 0.0222946f $X=6.545 $Y=0.35 $X2=0
+ $Y2=0
cc_701 N_A_722_23#_c_764_n N_VGND_c_1791_n 0.0801906f $X=6.38 $Y=0.19 $X2=0
+ $Y2=0
cc_702 N_A_722_23#_c_765_n N_VGND_c_1791_n 0.0047315f $X=3.76 $Y=0.19 $X2=0
+ $Y2=0
cc_703 N_A_722_23#_c_770_n N_VGND_c_1791_n 0.0193217f $X=6.38 $Y=0.345 $X2=0
+ $Y2=0
cc_704 N_A_722_23#_c_771_n N_VGND_c_1791_n 0.0101191f $X=5.795 $Y=0.345 $X2=0
+ $Y2=0
cc_705 N_A_722_23#_c_772_n N_VGND_c_1791_n 0.0112784f $X=6.545 $Y=0.35 $X2=0
+ $Y2=0
cc_706 N_A_1161_95#_c_912_n N_CLK_M1016_g 0.00635107f $X=8.705 $Y=3.11 $X2=0
+ $Y2=0
cc_707 N_A_1161_95#_c_896_n N_CLK_M1016_g 0.0358542f $X=7.685 $Y=1.795 $X2=0
+ $Y2=0
cc_708 N_A_1161_95#_c_898_n N_CLK_M1016_g 0.0344673f $X=8.78 $Y=3.035 $X2=0
+ $Y2=0
cc_709 N_A_1161_95#_c_902_n N_CLK_M1016_g 0.00486215f $X=8.82 $Y=1.49 $X2=0
+ $Y2=0
cc_710 N_A_1161_95#_c_904_n N_CLK_M1016_g 7.69803e-19 $X=7.57 $Y=1.29 $X2=0
+ $Y2=0
cc_711 N_A_1161_95#_c_907_n N_CLK_M1016_g 0.0017016f $X=8.82 $Y=1.06 $X2=0 $Y2=0
cc_712 N_A_1161_95#_c_909_n N_CLK_M1016_g 0.00960692f $X=8.32 $Y=1.9 $X2=0 $Y2=0
cc_713 N_A_1161_95#_c_910_n N_CLK_M1016_g 0.0141112f $X=8.802 $Y=1.9 $X2=0 $Y2=0
cc_714 N_A_1161_95#_c_897_n CLK 0.00341247f $X=7.73 $Y=1.125 $X2=0 $Y2=0
cc_715 N_A_1161_95#_c_904_n CLK 0.0272748f $X=7.57 $Y=1.29 $X2=0 $Y2=0
cc_716 N_A_1161_95#_c_906_n CLK 0.0200185f $X=8.69 $Y=0.78 $X2=0 $Y2=0
cc_717 N_A_1161_95#_c_907_n CLK 0.0273811f $X=8.82 $Y=1.06 $X2=0 $Y2=0
cc_718 N_A_1161_95#_c_908_n CLK 0.00237033f $X=8.82 $Y=1.06 $X2=0 $Y2=0
cc_719 N_A_1161_95#_c_909_n CLK 0.0546571f $X=8.32 $Y=1.9 $X2=0 $Y2=0
cc_720 N_A_1161_95#_c_896_n N_CLK_c_1051_n 0.0133365f $X=7.685 $Y=1.795 $X2=0
+ $Y2=0
cc_721 N_A_1161_95#_c_906_n N_CLK_c_1051_n 0.00106896f $X=8.69 $Y=0.78 $X2=0
+ $Y2=0
cc_722 N_A_1161_95#_c_907_n N_CLK_c_1051_n 3.57422e-19 $X=8.82 $Y=1.06 $X2=0
+ $Y2=0
cc_723 N_A_1161_95#_c_908_n N_CLK_c_1051_n 0.0174512f $X=8.82 $Y=1.06 $X2=0
+ $Y2=0
cc_724 N_A_1161_95#_c_909_n N_CLK_c_1051_n 0.00291648f $X=8.32 $Y=1.9 $X2=0
+ $Y2=0
cc_725 N_A_1161_95#_c_910_n N_CLK_c_1051_n 0.00162667f $X=8.802 $Y=1.9 $X2=0
+ $Y2=0
cc_726 N_A_1161_95#_c_897_n N_CLK_c_1052_n 0.0131156f $X=7.73 $Y=1.125 $X2=0
+ $Y2=0
cc_727 N_A_1161_95#_c_904_n N_CLK_c_1052_n 2.23938e-19 $X=7.57 $Y=1.29 $X2=0
+ $Y2=0
cc_728 N_A_1161_95#_c_907_n N_CLK_c_1052_n 8.52579e-19 $X=8.82 $Y=1.06 $X2=0
+ $Y2=0
cc_729 N_A_1161_95#_c_908_n N_CLK_c_1052_n 0.00604227f $X=8.82 $Y=1.06 $X2=0
+ $Y2=0
cc_730 N_A_1161_95#_M1035_g N_A_2082_99#_M1011_g 0.0114537f $X=9.91 $Y=2.315
+ $X2=0 $Y2=0
cc_731 N_A_1161_95#_M1015_g N_A_2082_99#_M1011_g 0.0595632f $X=10.125 $Y=0.835
+ $X2=0 $Y2=0
cc_732 N_A_1161_95#_c_903_n N_A_2082_99#_M1011_g 0.00470649f $X=9.91 $Y=1.445
+ $X2=0 $Y2=0
cc_733 N_A_1161_95#_M1035_g N_A_2082_99#_c_1107_n 3.63407e-19 $X=9.91 $Y=2.315
+ $X2=0 $Y2=0
cc_734 N_A_1161_95#_M1035_g N_A_1873_497#_c_1212_n 0.0142092f $X=9.91 $Y=2.315
+ $X2=0 $Y2=0
cc_735 N_A_1161_95#_c_899_n N_A_1873_497#_c_1213_n 0.00271982f $X=9.835 $Y=1.49
+ $X2=0 $Y2=0
cc_736 N_A_1161_95#_M1015_g N_A_1873_497#_c_1213_n 0.0143184f $X=10.125 $Y=0.835
+ $X2=0 $Y2=0
cc_737 N_A_1161_95#_c_903_n N_A_1873_497#_c_1213_n 0.00975805f $X=9.91 $Y=1.445
+ $X2=0 $Y2=0
cc_738 N_A_1161_95#_c_899_n N_A_1873_497#_c_1214_n 0.0150945f $X=9.835 $Y=1.49
+ $X2=0 $Y2=0
cc_739 N_A_1161_95#_M1035_g N_A_1873_497#_c_1214_n 0.0089518f $X=9.91 $Y=2.315
+ $X2=0 $Y2=0
cc_740 N_A_1161_95#_c_903_n N_A_1873_497#_c_1214_n 0.00406439f $X=9.91 $Y=1.445
+ $X2=0 $Y2=0
cc_741 N_A_1161_95#_c_903_n N_A_1873_497#_c_1216_n 0.00972088f $X=9.91 $Y=1.445
+ $X2=0 $Y2=0
cc_742 N_A_1161_95#_c_912_n N_VPWR_c_1369_n 0.027252f $X=8.705 $Y=3.11 $X2=0
+ $Y2=0
cc_743 N_A_1161_95#_M1028_g N_VPWR_c_1369_n 0.00113877f $X=7.685 $Y=2.275 $X2=0
+ $Y2=0
cc_744 N_A_1161_95#_c_898_n N_VPWR_c_1369_n 0.00784876f $X=8.78 $Y=3.035 $X2=0
+ $Y2=0
cc_745 N_A_1161_95#_c_913_n N_VPWR_c_1377_n 0.0416312f $X=6.51 $Y=3.11 $X2=0
+ $Y2=0
cc_746 N_A_1161_95#_c_912_n N_VPWR_c_1378_n 0.0236603f $X=8.705 $Y=3.11 $X2=0
+ $Y2=0
cc_747 N_A_1161_95#_c_912_n N_VPWR_c_1365_n 0.0582731f $X=8.705 $Y=3.11 $X2=0
+ $Y2=0
cc_748 N_A_1161_95#_c_913_n N_VPWR_c_1365_n 0.00542714f $X=6.51 $Y=3.11 $X2=0
+ $Y2=0
cc_749 N_A_1161_95#_M1028_g N_VPWR_c_1365_n 9.21552e-19 $X=7.685 $Y=2.275 $X2=0
+ $Y2=0
cc_750 N_A_1161_95#_c_895_n N_A_196_119#_c_1511_n 0.00397153f $X=5.955 $Y=1.21
+ $X2=0 $Y2=0
cc_751 N_A_1161_95#_c_893_n N_A_196_119#_c_1513_n 0.00492241f $X=5.88 $Y=1.135
+ $X2=0 $Y2=0
cc_752 N_A_1161_95#_c_894_n N_A_196_119#_c_1513_n 0.019793f $X=7.405 $Y=1.21
+ $X2=0 $Y2=0
cc_753 N_A_1161_95#_c_911_n N_A_974_425#_c_1671_n 0.0112597f $X=6.435 $Y=3.035
+ $X2=0 $Y2=0
cc_754 N_A_1161_95#_c_912_n N_A_974_425#_c_1671_n 6.78191e-19 $X=8.705 $Y=3.11
+ $X2=0 $Y2=0
cc_755 N_A_1161_95#_c_913_n N_A_974_425#_c_1671_n 0.00209531f $X=6.51 $Y=3.11
+ $X2=0 $Y2=0
cc_756 N_A_1161_95#_c_911_n N_A_974_425#_c_1673_n 0.00123565f $X=6.435 $Y=3.035
+ $X2=0 $Y2=0
cc_757 N_A_1161_95#_c_912_n N_A_974_425#_c_1673_n 0.0112325f $X=8.705 $Y=3.11
+ $X2=0 $Y2=0
cc_758 N_A_1161_95#_M1035_g N_A_1786_497#_c_1705_n 0.0105479f $X=9.91 $Y=2.315
+ $X2=0 $Y2=0
cc_759 N_A_1161_95#_M1035_g N_A_1786_497#_c_1706_n 0.00418845f $X=9.91 $Y=2.315
+ $X2=0 $Y2=0
cc_760 N_A_1161_95#_c_898_n N_A_1786_497#_c_1707_n 0.00825403f $X=8.78 $Y=3.035
+ $X2=0 $Y2=0
cc_761 N_A_1161_95#_c_897_n N_VGND_c_1778_n 0.00178847f $X=7.73 $Y=1.125 $X2=0
+ $Y2=0
cc_762 N_A_1161_95#_c_906_n N_VGND_c_1788_n 0.0129231f $X=8.69 $Y=0.78 $X2=0
+ $Y2=0
cc_763 N_A_1161_95#_c_897_n N_VGND_c_1791_n 9.39239e-19 $X=7.73 $Y=1.125 $X2=0
+ $Y2=0
cc_764 N_A_1161_95#_M1015_g N_VGND_c_1791_n 9.49986e-19 $X=10.125 $Y=0.835 $X2=0
+ $Y2=0
cc_765 N_A_1161_95#_c_906_n N_VGND_c_1791_n 0.0174119f $X=8.69 $Y=0.78 $X2=0
+ $Y2=0
cc_766 N_CLK_M1016_g N_VPWR_c_1369_n 0.00119146f $X=8.27 $Y=2.275 $X2=0 $Y2=0
cc_767 N_CLK_M1016_g N_VPWR_c_1365_n 9.21552e-19 $X=8.27 $Y=2.275 $X2=0 $Y2=0
cc_768 CLK N_VGND_c_1778_n 0.018094f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_769 N_CLK_c_1052_n N_VGND_c_1778_n 0.00360122f $X=8.25 $Y=1.13 $X2=0 $Y2=0
cc_770 N_CLK_c_1052_n N_VGND_c_1791_n 9.39239e-19 $X=8.25 $Y=1.13 $X2=0 $Y2=0
cc_771 N_A_2082_99#_M1011_g N_A_1873_497#_c_1211_n 0.021727f $X=10.485 $Y=0.835
+ $X2=0 $Y2=0
cc_772 N_A_2082_99#_c_1096_n N_A_1873_497#_c_1211_n 0.00308846f $X=11.645
+ $Y=1.645 $X2=0 $Y2=0
cc_773 N_A_2082_99#_c_1103_n N_A_1873_497#_M1022_g 0.0155487f $X=11.505 $Y=1.89
+ $X2=0 $Y2=0
cc_774 N_A_2082_99#_c_1105_n N_A_1873_497#_M1022_g 0.00102156f $X=11.62 $Y=2.04
+ $X2=0 $Y2=0
cc_775 N_A_2082_99#_c_1106_n N_A_1873_497#_M1022_g 0.0166017f $X=10.575 $Y=1.88
+ $X2=0 $Y2=0
cc_776 N_A_2082_99#_M1011_g N_A_1873_497#_c_1212_n 8.08117e-19 $X=10.485
+ $Y=0.835 $X2=0 $Y2=0
cc_777 N_A_2082_99#_c_1107_n N_A_1873_497#_c_1212_n 0.00266857f $X=10.74 $Y=1.88
+ $X2=0 $Y2=0
cc_778 N_A_2082_99#_M1011_g N_A_1873_497#_c_1213_n 0.0023806f $X=10.485 $Y=0.835
+ $X2=0 $Y2=0
cc_779 N_A_2082_99#_c_1103_n N_A_1873_497#_c_1215_n 0.0237005f $X=11.505 $Y=1.89
+ $X2=0 $Y2=0
cc_780 N_A_2082_99#_c_1096_n N_A_1873_497#_c_1215_n 0.0270793f $X=11.645
+ $Y=1.645 $X2=0 $Y2=0
cc_781 N_A_2082_99#_M1011_g N_A_1873_497#_c_1216_n 0.015806f $X=10.485 $Y=0.835
+ $X2=0 $Y2=0
cc_782 N_A_2082_99#_c_1103_n N_A_1873_497#_c_1216_n 0.0183826f $X=11.505 $Y=1.89
+ $X2=0 $Y2=0
cc_783 N_A_2082_99#_c_1106_n N_A_1873_497#_c_1216_n 0.0054842f $X=10.575 $Y=1.88
+ $X2=0 $Y2=0
cc_784 N_A_2082_99#_c_1107_n N_A_1873_497#_c_1216_n 0.0232333f $X=10.74 $Y=1.88
+ $X2=0 $Y2=0
cc_785 N_A_2082_99#_c_1103_n N_A_1873_497#_c_1217_n 0.00806573f $X=11.505
+ $Y=1.89 $X2=0 $Y2=0
cc_786 N_A_2082_99#_c_1096_n N_A_1873_497#_c_1217_n 0.013149f $X=11.645 $Y=1.645
+ $X2=0 $Y2=0
cc_787 N_A_2082_99#_c_1104_n N_A_1873_497#_c_1217_n 0.0044637f $X=11.645
+ $Y=1.805 $X2=0 $Y2=0
cc_788 N_A_2082_99#_M1034_g N_A_2409_367#_c_1272_n 0.0036316f $X=12.385 $Y=2.155
+ $X2=0 $Y2=0
cc_789 N_A_2082_99#_c_1088_n N_A_2409_367#_c_1272_n 0.012368f $X=12.835 $Y=1.57
+ $X2=0 $Y2=0
cc_790 N_A_2082_99#_M1024_g N_A_2409_367#_c_1272_n 0.00150362f $X=12.91 $Y=2.465
+ $X2=0 $Y2=0
cc_791 N_A_2082_99#_M1025_g N_A_2409_367#_c_1272_n 0.00147751f $X=13.31 $Y=0.815
+ $X2=0 $Y2=0
cc_792 N_A_2082_99#_c_1092_n N_A_2409_367#_c_1272_n 0.00510044f $X=12.375
+ $Y=0.975 $X2=0 $Y2=0
cc_793 N_A_2082_99#_c_1097_n N_A_2409_367#_c_1272_n 0.0504652f $X=12.375 $Y=1.14
+ $X2=0 $Y2=0
cc_794 N_A_2082_99#_c_1098_n N_A_2409_367#_c_1272_n 0.00641283f $X=12.375
+ $Y=1.14 $X2=0 $Y2=0
cc_795 N_A_2082_99#_M1024_g N_A_2409_367#_c_1279_n 0.0189233f $X=12.91 $Y=2.465
+ $X2=0 $Y2=0
cc_796 N_A_2082_99#_c_1090_n N_A_2409_367#_c_1279_n 9.84987e-19 $X=13.235
+ $Y=1.57 $X2=0 $Y2=0
cc_797 N_A_2082_99#_M1024_g N_A_2409_367#_c_1273_n 0.00426383f $X=12.91 $Y=2.465
+ $X2=0 $Y2=0
cc_798 N_A_2082_99#_M1025_g N_A_2409_367#_c_1273_n 3.7339e-19 $X=13.31 $Y=0.815
+ $X2=0 $Y2=0
cc_799 N_A_2082_99#_M1024_g N_A_2409_367#_c_1274_n 3.13166e-19 $X=12.91 $Y=2.465
+ $X2=0 $Y2=0
cc_800 N_A_2082_99#_M1025_g N_A_2409_367#_c_1274_n 0.0160765f $X=13.31 $Y=0.815
+ $X2=0 $Y2=0
cc_801 N_A_2082_99#_M1034_g N_A_2409_367#_c_1282_n 0.0249937f $X=12.385 $Y=2.155
+ $X2=0 $Y2=0
cc_802 N_A_2082_99#_c_1088_n N_A_2409_367#_c_1282_n 0.00480667f $X=12.835
+ $Y=1.57 $X2=0 $Y2=0
cc_803 N_A_2082_99#_M1024_g N_A_2409_367#_c_1282_n 0.00301479f $X=12.91 $Y=2.465
+ $X2=0 $Y2=0
cc_804 N_A_2082_99#_c_1094_n N_A_2409_367#_c_1282_n 0.00268875f $X=12.375
+ $Y=1.57 $X2=0 $Y2=0
cc_805 N_A_2082_99#_c_1105_n N_A_2409_367#_c_1282_n 0.0377683f $X=11.62 $Y=2.04
+ $X2=0 $Y2=0
cc_806 N_A_2082_99#_c_1097_n N_A_2409_367#_c_1282_n 0.040399f $X=12.375 $Y=1.14
+ $X2=0 $Y2=0
cc_807 N_A_2082_99#_c_1108_n N_A_2409_367#_c_1282_n 0.0123981f $X=11.645 $Y=1.89
+ $X2=0 $Y2=0
cc_808 N_A_2082_99#_c_1088_n N_A_2409_367#_c_1275_n 5.23078e-19 $X=12.835
+ $Y=1.57 $X2=0 $Y2=0
cc_809 N_A_2082_99#_M1025_g N_A_2409_367#_c_1275_n 7.45467e-19 $X=13.31 $Y=0.815
+ $X2=0 $Y2=0
cc_810 N_A_2082_99#_c_1098_n N_A_2409_367#_c_1275_n 0.0033862f $X=12.375 $Y=1.14
+ $X2=0 $Y2=0
cc_811 N_A_2082_99#_M1025_g N_A_2409_367#_c_1276_n 0.0123497f $X=13.31 $Y=0.815
+ $X2=0 $Y2=0
cc_812 N_A_2082_99#_c_1103_n N_VPWR_M1006_d 0.00227667f $X=11.505 $Y=1.89 $X2=0
+ $Y2=0
cc_813 N_A_2082_99#_c_1100_n N_VPWR_c_1370_n 0.00519336f $X=10.86 $Y=2.095 $X2=0
+ $Y2=0
cc_814 N_A_2082_99#_c_1103_n N_VPWR_c_1370_n 0.0241141f $X=11.505 $Y=1.89 $X2=0
+ $Y2=0
cc_815 N_A_2082_99#_c_1105_n N_VPWR_c_1370_n 0.023917f $X=11.62 $Y=2.04 $X2=0
+ $Y2=0
cc_816 N_A_2082_99#_M1024_g N_VPWR_c_1371_n 0.0272495f $X=12.91 $Y=2.465 $X2=0
+ $Y2=0
cc_817 N_A_2082_99#_M1024_g N_VPWR_c_1372_n 0.0123669f $X=12.91 $Y=2.465 $X2=0
+ $Y2=0
cc_818 N_A_2082_99#_M1034_g N_VPWR_c_1379_n 0.00312414f $X=12.385 $Y=2.155 $X2=0
+ $Y2=0
cc_819 N_A_2082_99#_c_1105_n N_VPWR_c_1379_n 0.00640219f $X=11.62 $Y=2.04 $X2=0
+ $Y2=0
cc_820 N_A_2082_99#_M1024_g N_VPWR_c_1380_n 0.00486043f $X=12.91 $Y=2.465 $X2=0
+ $Y2=0
cc_821 N_A_2082_99#_c_1100_n N_VPWR_c_1365_n 8.0667e-19 $X=10.86 $Y=2.095 $X2=0
+ $Y2=0
cc_822 N_A_2082_99#_M1034_g N_VPWR_c_1365_n 0.00410284f $X=12.385 $Y=2.155 $X2=0
+ $Y2=0
cc_823 N_A_2082_99#_M1024_g N_VPWR_c_1365_n 0.00600853f $X=12.91 $Y=2.465 $X2=0
+ $Y2=0
cc_824 N_A_2082_99#_c_1105_n N_VPWR_c_1365_n 0.00771299f $X=11.62 $Y=2.04 $X2=0
+ $Y2=0
cc_825 N_A_2082_99#_c_1100_n N_A_1786_497#_c_1705_n 0.00126569f $X=10.86
+ $Y=2.095 $X2=0 $Y2=0
cc_826 N_A_2082_99#_c_1106_n N_A_1786_497#_c_1705_n 0.00183976f $X=10.575
+ $Y=1.88 $X2=0 $Y2=0
cc_827 N_A_2082_99#_c_1100_n N_A_1786_497#_c_1706_n 0.00775432f $X=10.86
+ $Y=2.095 $X2=0 $Y2=0
cc_828 N_A_2082_99#_c_1106_n N_A_1786_497#_c_1706_n 0.0077637f $X=10.575 $Y=1.88
+ $X2=0 $Y2=0
cc_829 N_A_2082_99#_c_1107_n N_A_1786_497#_c_1706_n 0.0164339f $X=10.74 $Y=1.88
+ $X2=0 $Y2=0
cc_830 N_A_2082_99#_c_1090_n Q 0.00679927f $X=13.235 $Y=1.57 $X2=0 $Y2=0
cc_831 N_A_2082_99#_M1025_g Q 0.0100467f $X=13.31 $Y=0.815 $X2=0 $Y2=0
cc_832 N_A_2082_99#_M1024_g Q 0.00428114f $X=12.91 $Y=2.465 $X2=0 $Y2=0
cc_833 N_A_2082_99#_c_1090_n Q 0.0138226f $X=13.235 $Y=1.57 $X2=0 $Y2=0
cc_834 N_A_2082_99#_M1025_g N_Q_c_1738_n 0.0185425f $X=13.31 $Y=0.815 $X2=0
+ $Y2=0
cc_835 N_A_2082_99#_c_1092_n N_Q_c_1738_n 0.00278156f $X=12.375 $Y=0.975 $X2=0
+ $Y2=0
cc_836 N_A_2082_99#_M1011_g N_VGND_c_1779_n 0.013886f $X=10.485 $Y=0.835 $X2=0
+ $Y2=0
cc_837 N_A_2082_99#_c_1096_n N_VGND_c_1779_n 0.0246671f $X=11.645 $Y=1.645 $X2=0
+ $Y2=0
cc_838 N_A_2082_99#_c_1092_n N_VGND_c_1780_n 0.00386049f $X=12.375 $Y=0.975
+ $X2=0 $Y2=0
cc_839 N_A_2082_99#_c_1096_n N_VGND_c_1780_n 0.0122143f $X=11.645 $Y=1.645 $X2=0
+ $Y2=0
cc_840 N_A_2082_99#_c_1097_n N_VGND_c_1780_n 0.0242884f $X=12.375 $Y=1.14 $X2=0
+ $Y2=0
cc_841 N_A_2082_99#_c_1098_n N_VGND_c_1780_n 0.00145897f $X=12.375 $Y=1.14 $X2=0
+ $Y2=0
cc_842 N_A_2082_99#_M1025_g N_VGND_c_1781_n 0.00543974f $X=13.31 $Y=0.815 $X2=0
+ $Y2=0
cc_843 N_A_2082_99#_M1025_g N_VGND_c_1784_n 0.00507333f $X=13.31 $Y=0.815 $X2=0
+ $Y2=0
cc_844 N_A_2082_99#_c_1092_n N_VGND_c_1784_n 0.00523993f $X=12.375 $Y=0.975
+ $X2=0 $Y2=0
cc_845 N_A_2082_99#_c_1096_n N_VGND_c_1789_n 0.0111137f $X=11.645 $Y=1.645 $X2=0
+ $Y2=0
cc_846 N_A_2082_99#_M1011_g N_VGND_c_1791_n 9.49986e-19 $X=10.485 $Y=0.835 $X2=0
+ $Y2=0
cc_847 N_A_2082_99#_M1025_g N_VGND_c_1791_n 0.00537853f $X=13.31 $Y=0.815 $X2=0
+ $Y2=0
cc_848 N_A_2082_99#_c_1092_n N_VGND_c_1791_n 0.0052212f $X=12.375 $Y=0.975 $X2=0
+ $Y2=0
cc_849 N_A_2082_99#_c_1096_n N_VGND_c_1791_n 0.0137775f $X=11.645 $Y=1.645 $X2=0
+ $Y2=0
cc_850 N_A_1873_497#_M1022_g N_VPWR_c_1370_n 0.0114703f $X=11.385 $Y=2.315 $X2=0
+ $Y2=0
cc_851 N_A_1873_497#_M1022_g N_VPWR_c_1365_n 7.88961e-19 $X=11.385 $Y=2.315
+ $X2=0 $Y2=0
cc_852 N_A_1873_497#_M1002_d N_A_1786_497#_c_1705_n 0.00527944f $X=9.365
+ $Y=2.485 $X2=0 $Y2=0
cc_853 N_A_1873_497#_M1022_g N_A_1786_497#_c_1705_n 4.54107e-19 $X=11.385
+ $Y=2.315 $X2=0 $Y2=0
cc_854 N_A_1873_497#_c_1211_n N_VGND_c_1779_n 0.00953128f $X=11.08 $Y=1.375
+ $X2=0 $Y2=0
cc_855 N_A_1873_497#_c_1213_n N_VGND_c_1779_n 0.0122365f $X=9.91 $Y=0.9 $X2=0
+ $Y2=0
cc_856 N_A_1873_497#_c_1216_n N_VGND_c_1779_n 0.0197316f $X=11.005 $Y=1.54 $X2=0
+ $Y2=0
cc_857 N_A_1873_497#_c_1211_n N_VGND_c_1791_n 9.24653e-19 $X=11.08 $Y=1.375
+ $X2=0 $Y2=0
cc_858 N_A_1873_497#_c_1213_n N_VGND_c_1791_n 0.01192f $X=9.91 $Y=0.9 $X2=0
+ $Y2=0
cc_859 N_A_2409_367#_c_1282_n N_VPWR_M1034_d 0.00493955f $X=12.81 $Y=2.155 $X2=0
+ $Y2=0
cc_860 N_A_2409_367#_c_1279_n N_VPWR_M1026_s 0.00450523f $X=13.625 $Y=2.41 $X2=0
+ $Y2=0
cc_861 N_A_2409_367#_c_1273_n N_VPWR_M1026_s 0.0078218f $X=13.79 $Y=1.51 $X2=0
+ $Y2=0
cc_862 N_A_2409_367#_c_1282_n N_VPWR_c_1371_n 0.0234949f $X=12.81 $Y=2.155 $X2=0
+ $Y2=0
cc_863 N_A_2409_367#_M1026_g N_VPWR_c_1372_n 0.0138465f $X=13.925 $Y=2.465 $X2=0
+ $Y2=0
cc_864 N_A_2409_367#_c_1279_n N_VPWR_c_1372_n 0.0230391f $X=13.625 $Y=2.41 $X2=0
+ $Y2=0
cc_865 N_A_2409_367#_M1026_g N_VPWR_c_1381_n 0.00486043f $X=13.925 $Y=2.465
+ $X2=0 $Y2=0
cc_866 N_A_2409_367#_M1026_g N_VPWR_c_1365_n 0.00917987f $X=13.925 $Y=2.465
+ $X2=0 $Y2=0
cc_867 N_A_2409_367#_c_1279_n N_VPWR_c_1365_n 0.0240967f $X=13.625 $Y=2.41 $X2=0
+ $Y2=0
cc_868 N_A_2409_367#_c_1282_n N_VPWR_c_1365_n 0.0213928f $X=12.81 $Y=2.155 $X2=0
+ $Y2=0
cc_869 N_A_2409_367#_c_1279_n N_Q_M1024_d 0.00706161f $X=13.625 $Y=2.41 $X2=0
+ $Y2=0
cc_870 N_A_2409_367#_c_1273_n Q 0.0535947f $X=13.79 $Y=1.51 $X2=0 $Y2=0
cc_871 N_A_2409_367#_c_1274_n Q 0.00221851f $X=13.79 $Y=1.51 $X2=0 $Y2=0
cc_872 N_A_2409_367#_M1026_g Q 0.0021663f $X=13.925 $Y=2.465 $X2=0 $Y2=0
cc_873 N_A_2409_367#_c_1279_n Q 0.0287045f $X=13.625 $Y=2.41 $X2=0 $Y2=0
cc_874 N_A_2409_367#_c_1282_n Q 0.00155324f $X=12.81 $Y=2.155 $X2=0 $Y2=0
cc_875 N_A_2409_367#_c_1272_n N_Q_c_1738_n 0.0752625f $X=12.725 $Y=1.815 $X2=0
+ $Y2=0
cc_876 N_A_2409_367#_c_1275_n N_Q_c_1738_n 0.025858f $X=12.725 $Y=0.64 $X2=0
+ $Y2=0
cc_877 N_A_2409_367#_c_1276_n N_Q_c_1738_n 0.00102315f $X=13.812 $Y=1.345 $X2=0
+ $Y2=0
cc_878 N_A_2409_367#_c_1274_n Q_N 0.00578206f $X=13.79 $Y=1.51 $X2=0 $Y2=0
cc_879 N_A_2409_367#_c_1273_n Q_N 0.0549046f $X=13.79 $Y=1.51 $X2=0 $Y2=0
cc_880 N_A_2409_367#_c_1274_n Q_N 0.0154054f $X=13.79 $Y=1.51 $X2=0 $Y2=0
cc_881 N_A_2409_367#_c_1276_n Q_N 0.00582627f $X=13.812 $Y=1.345 $X2=0 $Y2=0
cc_882 N_A_2409_367#_c_1276_n N_Q_N_c_1761_n 0.00147405f $X=13.812 $Y=1.345
+ $X2=0 $Y2=0
cc_883 N_A_2409_367#_c_1276_n N_VGND_c_1781_n 0.0035146f $X=13.812 $Y=1.345
+ $X2=0 $Y2=0
cc_884 N_A_2409_367#_c_1275_n N_VGND_c_1784_n 0.00950487f $X=12.725 $Y=0.64
+ $X2=0 $Y2=0
cc_885 N_A_2409_367#_c_1276_n N_VGND_c_1790_n 0.00559701f $X=13.812 $Y=1.345
+ $X2=0 $Y2=0
cc_886 N_A_2409_367#_c_1275_n N_VGND_c_1791_n 0.0122344f $X=12.725 $Y=0.64 $X2=0
+ $Y2=0
cc_887 N_A_2409_367#_c_1276_n N_VGND_c_1791_n 0.00537853f $X=13.812 $Y=1.345
+ $X2=0 $Y2=0
cc_888 N_A_27_483#_c_1338_n N_VPWR_M1017_d 0.00176461f $X=1.745 $Y=2.375
+ $X2=-0.19 $Y2=1.655
cc_889 N_A_27_483#_c_1337_n N_VPWR_c_1366_n 0.0166834f $X=0.26 $Y=2.56 $X2=0
+ $Y2=0
cc_890 N_A_27_483#_c_1338_n N_VPWR_c_1366_n 0.0170436f $X=1.745 $Y=2.375 $X2=0
+ $Y2=0
cc_891 N_A_27_483#_c_1337_n N_VPWR_c_1375_n 0.0173955f $X=0.26 $Y=2.56 $X2=0
+ $Y2=0
cc_892 N_A_27_483#_c_1337_n N_VPWR_c_1365_n 0.00998284f $X=0.26 $Y=2.56 $X2=0
+ $Y2=0
cc_893 N_A_27_483#_c_1338_n A_196_483# 0.00366293f $X=1.745 $Y=2.375 $X2=-0.19
+ $Y2=1.655
cc_894 N_A_27_483#_c_1338_n N_A_196_119#_M1000_d 0.00257467f $X=1.745 $Y=2.375
+ $X2=0 $Y2=0
cc_895 N_A_27_483#_M1020_d N_A_196_119#_c_1515_n 0.00303242f $X=1.77 $Y=2.415
+ $X2=0 $Y2=0
cc_896 N_A_27_483#_c_1338_n N_A_196_119#_c_1515_n 0.0123684f $X=1.745 $Y=2.375
+ $X2=0 $Y2=0
cc_897 N_A_27_483#_c_1340_n N_A_196_119#_c_1515_n 0.0204042f $X=1.91 $Y=2.375
+ $X2=0 $Y2=0
cc_898 N_A_27_483#_c_1340_n N_A_196_119#_c_1504_n 0.0284387f $X=1.91 $Y=2.375
+ $X2=0 $Y2=0
cc_899 N_VPWR_c_1366_n N_A_196_119#_c_1515_n 0.0080909f $X=0.69 $Y=2.755 $X2=0
+ $Y2=0
cc_900 N_VPWR_c_1373_n N_A_196_119#_c_1515_n 0.0576265f $X=3.315 $Y=3.33 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_1365_n N_A_196_119#_c_1515_n 0.0345592f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_902 N_VPWR_c_1367_n N_A_196_119#_c_1517_n 0.0137976f $X=3.41 $Y=2.89 $X2=0
+ $Y2=0
cc_903 N_VPWR_c_1373_n N_A_196_119#_c_1517_n 0.044618f $X=3.315 $Y=3.33 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_1365_n N_A_196_119#_c_1517_n 0.0269405f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_905 N_VPWR_c_1367_n N_A_196_119#_c_1550_n 0.0123063f $X=3.41 $Y=2.89 $X2=0
+ $Y2=0
cc_906 N_VPWR_M1008_d N_A_196_119#_c_1521_n 0.00228329f $X=3.255 $Y=2.405 $X2=0
+ $Y2=0
cc_907 N_VPWR_M1004_d N_A_196_119#_c_1521_n 0.00489664f $X=4.345 $Y=2.125 $X2=0
+ $Y2=0
cc_908 N_VPWR_c_1367_n N_A_196_119#_c_1521_n 0.0205461f $X=3.41 $Y=2.89 $X2=0
+ $Y2=0
cc_909 N_VPWR_c_1368_n N_A_196_119#_c_1521_n 0.0214123f $X=4.485 $Y=2.82 $X2=0
+ $Y2=0
cc_910 N_VPWR_c_1365_n N_A_196_119#_c_1521_n 0.0414544f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_911 N_VPWR_c_1373_n N_A_196_119#_c_1522_n 0.0113943f $X=3.315 $Y=3.33 $X2=0
+ $Y2=0
cc_912 N_VPWR_c_1365_n N_A_196_119#_c_1522_n 0.00656694f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_913 N_VPWR_c_1377_n N_A_974_425#_c_1671_n 0.0774805f $X=7.83 $Y=3.33 $X2=0
+ $Y2=0
cc_914 N_VPWR_c_1365_n N_A_974_425#_c_1671_n 0.0464317f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_915 N_VPWR_c_1368_n N_A_974_425#_c_1672_n 0.0195442f $X=4.485 $Y=2.82 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1377_n N_A_974_425#_c_1672_n 0.0210061f $X=7.83 $Y=3.33 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1365_n N_A_974_425#_c_1672_n 0.0111577f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_918 N_VPWR_c_1377_n N_A_974_425#_c_1673_n 0.0201327f $X=7.83 $Y=3.33 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1365_n N_A_974_425#_c_1673_n 0.0109922f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1370_n N_A_1786_497#_c_1705_n 0.0194269f $X=11.17 $Y=2.23 $X2=0
+ $Y2=0
cc_921 N_VPWR_c_1378_n N_A_1786_497#_c_1705_n 0.0129199f $X=10.98 $Y=3.33 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1365_n N_A_1786_497#_c_1705_n 0.0106163f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1370_n N_A_1786_497#_c_1706_n 0.0221379f $X=11.17 $Y=2.23 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1378_n N_A_1786_497#_c_1707_n 0.0562509f $X=10.98 $Y=3.33 $X2=0
+ $Y2=0
cc_925 N_VPWR_c_1365_n N_A_1786_497#_c_1707_n 0.0494203f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1365_n N_Q_M1024_d 0.00389753f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_927 N_VPWR_c_1365_n N_Q_N_M1026_d 0.00371702f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_928 N_VPWR_c_1381_n Q_N 0.018528f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_929 N_VPWR_c_1365_n Q_N 0.0104192f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_930 N_A_196_119#_c_1521_n N_A_974_425#_M1023_d 0.00761826f $X=5.545 $Y=2.47
+ $X2=-0.19 $Y2=-0.245
cc_931 N_A_196_119#_M1010_s N_A_974_425#_c_1671_n 0.0032654f $X=5.565 $Y=2.505
+ $X2=0 $Y2=0
cc_932 N_A_196_119#_c_1521_n N_A_974_425#_c_1671_n 0.010204f $X=5.545 $Y=2.47
+ $X2=0 $Y2=0
cc_933 N_A_196_119#_c_1523_n N_A_974_425#_c_1671_n 0.0237223f $X=5.71 $Y=2.47
+ $X2=0 $Y2=0
cc_934 N_A_196_119#_c_1521_n N_A_974_425#_c_1672_n 0.0247179f $X=5.545 $Y=2.47
+ $X2=0 $Y2=0
cc_935 N_A_196_119#_c_1510_n N_VGND_M1005_d 0.0068223f $X=4.32 $Y=1.335 $X2=0
+ $Y2=0
cc_936 N_A_196_119#_c_1503_n N_VGND_c_1776_n 0.0120188f $X=2.255 $Y=1.31 $X2=0
+ $Y2=0
cc_937 N_A_196_119#_c_1514_n N_VGND_c_1776_n 0.00105969f $X=1.785 $Y=1.09 $X2=0
+ $Y2=0
cc_938 N_A_196_119#_c_1508_n N_VGND_c_1777_n 0.0150385f $X=4.235 $Y=0.35 $X2=0
+ $Y2=0
cc_939 N_A_196_119#_c_1510_n N_VGND_c_1777_n 0.0562361f $X=4.32 $Y=1.335 $X2=0
+ $Y2=0
cc_940 N_A_196_119#_c_1511_n N_VGND_c_1777_n 0.0271222f $X=5.965 $Y=1.42 $X2=0
+ $Y2=0
cc_941 N_A_196_119#_c_1508_n N_VGND_c_1782_n 0.0516118f $X=4.235 $Y=0.35 $X2=0
+ $Y2=0
cc_942 N_A_196_119#_c_1509_n N_VGND_c_1782_n 0.0114622f $X=3.555 $Y=0.35 $X2=0
+ $Y2=0
cc_943 N_A_196_119#_c_1558_n N_VGND_c_1786_n 0.00567329f $X=1.175 $Y=0.805 $X2=0
+ $Y2=0
cc_944 N_A_196_119#_c_1558_n N_VGND_c_1791_n 0.00851804f $X=1.175 $Y=0.805 $X2=0
+ $Y2=0
cc_945 N_A_196_119#_c_1508_n N_VGND_c_1791_n 0.0285895f $X=4.235 $Y=0.35 $X2=0
+ $Y2=0
cc_946 N_A_196_119#_c_1509_n N_VGND_c_1791_n 0.00657784f $X=3.555 $Y=0.35 $X2=0
+ $Y2=0
cc_947 N_A_196_119#_c_1501_n A_304_119# 0.00366293f $X=1.7 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_948 N_Q_c_1738_n N_VGND_c_1781_n 0.0597301f $X=13.095 $Y=0.54 $X2=0 $Y2=0
cc_949 N_Q_c_1738_n N_VGND_c_1784_n 0.0117388f $X=13.095 $Y=0.54 $X2=0 $Y2=0
cc_950 N_Q_c_1738_n N_VGND_c_1791_n 0.0106146f $X=13.095 $Y=0.54 $X2=0 $Y2=0
cc_951 N_Q_N_c_1761_n N_VGND_c_1781_n 0.00157726f $X=13.97 $Y=0.54 $X2=0 $Y2=0
cc_952 N_Q_N_c_1761_n N_VGND_c_1790_n 0.0189751f $X=13.97 $Y=0.54 $X2=0 $Y2=0
cc_953 N_Q_N_c_1761_n N_VGND_c_1791_n 0.017022f $X=13.97 $Y=0.54 $X2=0 $Y2=0
