* File: sky130_fd_sc_lp__and2_1.spice
* Created: Wed Sep  2 09:30:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and2_1.pex.spice"
.subckt sky130_fd_sc_lp__and2_1  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 A_175_131# N_A_M1005_g N_A_92_131#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g A_175_131# VNB NSHORT L=0.15 W=0.42 AD=0.0973
+ AS=0.0441 PD=0.82 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_92_131#_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2478 AS=0.1946 PD=2.27 PS=1.64 NRD=0 NRS=7.848 M=1 R=5.6 SA=75000.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_92_131#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=32.8202 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_B_M1002_g N_A_92_131#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.101325 AS=0.0819 PD=0.8475 PS=0.81 NRD=87.3498 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_92_131#_M1001_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.303975 PD=3.05 PS=2.5425 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__and2_1.pxi.spice"
*
.ends
*
*
