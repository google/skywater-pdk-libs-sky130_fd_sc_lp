* File: sky130_fd_sc_lp__srsdfrtp_1.pex.spice
* Created: Wed Sep  2 10:39:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%SCE 3 7 9 11 15 19 22 24 25 26 30
c59 11 0 6.29175e-20 $X=1.415 $Y=2.095
c60 9 0 1.01062e-19 $X=1.51 $Y=1.525
c61 3 0 2.11477e-20 $X=0.485 $Y=0.76
r62 25 26 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.77 $Y=1.665
+ $X2=0.77 $Y2=2.035
r63 25 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.77
+ $Y=1.665 $X2=0.77 $Y2=1.665
r64 23 30 42.9206 $w=4.6e-07 $l=3.55e-07 $layer=POLY_cond $X=0.72 $Y=2.02
+ $X2=0.72 $Y2=1.665
r65 23 24 10.9339 $w=3.05e-07 $l=7.5e-08 $layer=POLY_cond $X=0.72 $Y=2.02
+ $X2=0.72 $Y2=2.095
r66 21 30 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=0.72 $Y=1.6 $X2=0.72
+ $Y2=1.665
r67 21 22 10.9339 $w=3.05e-07 $l=9.28709e-08 $layer=POLY_cond $X=0.72 $Y=1.6
+ $X2=0.68 $Y2=1.525
r68 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.585 $Y=1.45
+ $X2=1.585 $Y2=0.89
r69 13 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.49 $Y=2.17
+ $X2=1.49 $Y2=2.65
r70 12 24 15.748 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=0.95 $Y=2.095
+ $X2=0.72 $Y2=2.095
r71 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.415 $Y=2.095
+ $X2=1.49 $Y2=2.17
r72 11 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.415 $Y=2.095
+ $X2=0.95 $Y2=2.095
r73 10 22 15.748 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.95 $Y=1.525
+ $X2=0.68 $Y2=1.525
r74 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.51 $Y=1.525
+ $X2=1.585 $Y2=1.45
r75 9 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.51 $Y=1.525
+ $X2=0.95 $Y2=1.525
r76 5 24 10.9339 $w=3.05e-07 $l=1.88812e-07 $layer=POLY_cond $X=0.565 $Y=2.17
+ $X2=0.72 $Y2=2.095
r77 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.565 $Y=2.17
+ $X2=0.565 $Y2=2.65
r78 1 22 10.9339 $w=3.05e-07 $l=2.29456e-07 $layer=POLY_cond $X=0.485 $Y=1.45
+ $X2=0.68 $Y2=1.525
r79 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.485 $Y=1.45
+ $X2=0.485 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%D 3 7 9 13 14
c38 14 0 5.74567e-20 $X=1.97 $Y=2.005
c39 7 0 1.29647e-19 $X=2.235 $Y=0.89
r40 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=2.005 $X2=1.97 $Y2=2.005
r41 11 13 16.2472 $w=2.67e-07 $l=9e-08 $layer=POLY_cond $X=1.88 $Y=2.005
+ $X2=1.97 $Y2=2.005
r42 9 14 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=2.005
+ $X2=1.97 $Y2=2.005
r43 5 13 47.839 $w=2.67e-07 $l=3.37565e-07 $layer=POLY_cond $X=2.235 $Y=1.84
+ $X2=1.97 $Y2=2.005
r44 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.235 $Y=1.84
+ $X2=2.235 $Y2=0.89
r45 1 11 16.2448 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=2.17
+ $X2=1.88 $Y2=2.005
r46 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.88 $Y=2.17 $X2=1.88
+ $Y2=2.65
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_27_110# 1 2 9 13 17 21 23 26 27 28 30
+ 31 35 36
c86 36 0 5.74567e-20 $X=2.715 $Y=1.765
c87 30 0 1.01062e-19 $X=2.39 $Y=1.6
c88 23 0 6.29175e-20 $X=1.49 $Y=1.245
c89 9 0 1.84393e-19 $X=2.595 $Y=0.89
r90 36 40 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.765
+ $X2=2.7 $Y2=1.93
r91 36 39 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.765
+ $X2=2.7 $Y2=1.6
r92 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.715
+ $Y=1.765 $X2=2.715 $Y2=1.765
r93 32 35 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.39 $Y=1.765
+ $X2=2.715 $Y2=1.765
r94 30 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=1.6 $X2=2.39
+ $Y2=1.765
r95 29 30 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.39 $Y=0.765
+ $X2=2.39 $Y2=1.6
r96 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.305 $Y=0.68
+ $X2=2.39 $Y2=0.765
r97 27 28 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.305 $Y=0.68
+ $X2=1.66 $Y2=0.68
r98 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.575 $Y=0.765
+ $X2=1.66 $Y2=0.68
r99 25 26 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.575 $Y=0.765
+ $X2=1.575 $Y2=1.16
r100 24 31 3.3199 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=1.245
+ $X2=0.27 $Y2=1.245
r101 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.49 $Y=1.245
+ $X2=1.575 $Y2=1.16
r102 23 24 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=1.49 $Y=1.245
+ $X2=0.435 $Y2=1.245
r103 19 31 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=1.33
+ $X2=0.27 $Y2=1.245
r104 19 21 39.9863 $w=3.28e-07 $l=1.145e-06 $layer=LI1_cond $X=0.27 $Y=1.33
+ $X2=0.27 $Y2=2.475
r105 15 31 3.24686 $w=2.9e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.23 $Y=1.16
+ $X2=0.27 $Y2=1.245
r106 15 17 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.23 $Y=1.16 $X2=0.23
+ $Y2=0.76
r107 13 40 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.685 $Y=2.65
+ $X2=2.685 $Y2=1.93
r108 9 39 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.595 $Y=0.89
+ $X2=2.595 $Y2=1.6
r109 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.205
+ $Y=2.33 $X2=0.35 $Y2=2.475
r110 1 17 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.55 $X2=0.27 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%SCD 1 3 5 8 12 14 19
c37 14 0 1.84393e-19 $X=3.6 $Y=1.665
r38 16 19 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=3.195 $Y=1.715
+ $X2=3.515 $Y2=1.715
r39 14 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.515
+ $Y=1.715 $X2=3.515 $Y2=1.715
r40 10 12 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.025 $Y=1.285
+ $X2=3.195 $Y2=1.285
r41 6 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.88
+ $X2=3.195 $Y2=1.715
r42 6 8 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.195 $Y=1.88 $X2=3.195
+ $Y2=2.65
r43 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.55
+ $X2=3.195 $Y2=1.715
r44 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.195 $Y=1.36
+ $X2=3.195 $Y2=1.285
r45 4 5 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.195 $Y=1.36
+ $X2=3.195 $Y2=1.55
r46 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.025 $Y=1.21
+ $X2=3.025 $Y2=1.285
r47 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.025 $Y=1.21
+ $X2=3.025 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_969_318# 1 2 9 13 15 17 18 19 20 22 23
+ 25 27 29 30 31 32 34 37 39 40 42 45 49 53 61 63 65 72 73 80
c190 65 0 9.57414e-20 $X=9.375 $Y=1.58
c191 61 0 1.33414e-19 $X=8.99 $Y=1.5
c192 45 0 1.01483e-19 $X=5.05 $Y=1.755
c193 30 0 8.61052e-20 $X=5.78 $Y=2.685
r194 73 86 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=13.29 $Y=2.91
+ $X2=13.29 $Y2=3.135
r195 72 75 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=13.29 $Y=2.91
+ $X2=13.29 $Y2=2.99
r196 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.29
+ $Y=2.91 $X2=13.29 $Y2=2.91
r197 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.375
+ $Y=1.66 $X2=9.375 $Y2=1.66
r198 65 68 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.375 $Y=1.58
+ $X2=9.375 $Y2=1.66
r199 60 61 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.825 $Y=1.5
+ $X2=8.99 $Y2=1.5
r200 57 60 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=8.56 $Y=1.5
+ $X2=8.825 $Y2=1.5
r201 53 55 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=2.35
+ $X2=7.595 $Y2=2.515
r202 49 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.865 $Y=2.515
+ $X2=5.865 $Y2=2.685
r203 46 80 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.05 $Y=1.755
+ $X2=5.175 $Y2=1.755
r204 46 77 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.05 $Y=1.755
+ $X2=4.92 $Y2=1.755
r205 45 48 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.05 $Y=1.755
+ $X2=5.05 $Y2=1.92
r206 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=1.755 $X2=5.05 $Y2=1.755
r207 42 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.21 $Y=1.58
+ $X2=9.375 $Y2=1.58
r208 42 61 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.21 $Y=1.58
+ $X2=8.99 $Y2=1.58
r209 41 64 2.58477 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=2.99
+ $X2=8.56 $Y2=2.99
r210 40 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.125 $Y=2.99
+ $X2=13.29 $Y2=2.99
r211 40 41 287.059 $w=1.68e-07 $l=4.4e-06 $layer=LI1_cond $X=13.125 $Y=2.99
+ $X2=8.725 $Y2=2.99
r212 39 64 13.2697 $w=3.3e-07 $l=3.3e-07 $layer=LI1_cond $X=8.56 $Y=2.66
+ $X2=8.56 $Y2=2.99
r213 38 63 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.56 $Y=2.435
+ $X2=8.56 $Y2=2.35
r214 38 39 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=8.56 $Y=2.435
+ $X2=8.56 $Y2=2.66
r215 37 63 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.56 $Y=2.265
+ $X2=8.56 $Y2=2.35
r216 36 57 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.56 $Y=1.665
+ $X2=8.56 $Y2=1.5
r217 36 37 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=8.56 $Y=1.665
+ $X2=8.56 $Y2=2.265
r218 35 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.68 $Y=2.35
+ $X2=7.595 $Y2=2.35
r219 34 63 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.395 $Y=2.35
+ $X2=8.56 $Y2=2.35
r220 34 35 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=8.395 $Y=2.35
+ $X2=7.68 $Y2=2.35
r221 33 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=2.515
+ $X2=5.865 $Y2=2.515
r222 32 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.51 $Y=2.515
+ $X2=7.595 $Y2=2.515
r223 32 33 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=7.51 $Y=2.515
+ $X2=5.95 $Y2=2.515
r224 30 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.78 $Y=2.685
+ $X2=5.865 $Y2=2.685
r225 30 31 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.78 $Y=2.685
+ $X2=5.095 $Y2=2.685
r226 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.01 $Y=2.6
+ $X2=5.095 $Y2=2.685
r227 29 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.01 $Y=2.6
+ $X2=5.01 $Y2=1.92
r228 25 27 117.608 $w=2.5e-07 $l=6.1e-07 $layer=POLY_cond $X=14.055 $Y=3.06
+ $X2=14.055 $Y2=2.45
r229 24 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.455 $Y=3.135
+ $X2=13.29 $Y2=3.135
r230 23 25 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=13.93 $Y=3.135
+ $X2=14.055 $Y2=3.06
r231 23 24 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=13.93 $Y=3.135
+ $X2=13.455 $Y2=3.135
r232 20 22 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=9.94 $Y=1.365
+ $X2=9.94 $Y2=0.945
r233 19 69 29.374 $w=3.61e-07 $l=3.14307e-07 $layer=POLY_cond $X=9.655 $Y=1.44
+ $X2=9.432 $Y2=1.66
r234 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.865 $Y=1.44
+ $X2=9.94 $Y2=1.365
r235 18 19 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.865 $Y=1.44
+ $X2=9.655 $Y2=1.44
r236 15 19 26.9074 $w=3.61e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.58 $Y=1.365
+ $X2=9.655 $Y2=1.44
r237 15 17 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=9.58 $Y=1.365
+ $X2=9.58 $Y2=0.945
r238 11 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.175 $Y=1.59
+ $X2=5.175 $Y2=1.755
r239 11 13 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.175 $Y=1.59
+ $X2=5.175 $Y2=1.035
r240 7 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.92 $Y=1.92
+ $X2=4.92 $Y2=1.755
r241 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.92 $Y=1.92 $X2=4.92
+ $Y2=2.33
r242 2 63 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.42
+ $Y=2.165 $X2=8.56 $Y2=2.31
r243 1 60 182 $w=1.7e-07 $l=7.98154e-07 $layer=licon1_NDIFF $count=1 $X=8.58
+ $Y=0.815 $X2=8.825 $Y2=1.5
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_1176_349# 1 2 3 4 15 21 23 24 28 29 31
+ 32 36 40 41 46 47 48 51 55 57
c156 32 0 1.40585e-19 $X=7.965 $Y=1.97
c157 15 0 8.61052e-20 $X=5.955 $Y=2.33
r158 56 57 5.28416 $w=1.78e-07 $l=8.5e-08 $layer=LI1_cond $X=8.05 $Y=1.085
+ $X2=8.135 $Y2=1.085
r159 49 51 80.4405 $w=2.48e-07 $l=1.745e-06 $layer=LI1_cond $X=10.805 $Y=0.435
+ $X2=10.805 $Y2=2.18
r160 47 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.68 $Y=0.35
+ $X2=10.805 $Y2=0.435
r161 47 48 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=10.68 $Y=0.35
+ $X2=9.53 $Y2=0.35
r162 44 46 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=9.365 $Y=0.995
+ $X2=9.365 $Y2=0.77
r163 43 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.365 $Y=0.435
+ $X2=9.53 $Y2=0.35
r164 43 46 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.365 $Y=0.435
+ $X2=9.365 $Y2=0.77
r165 41 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.2 $Y=1.08
+ $X2=9.365 $Y2=0.995
r166 41 57 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=9.2 $Y=1.08
+ $X2=8.135 $Y2=1.08
r167 39 56 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.05 $Y=1.175 $X2=8.05
+ $Y2=1.085
r168 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.05 $Y=1.175
+ $X2=8.05 $Y2=1.845
r169 36 56 20.6414 $w=1.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.715 $Y=1.085
+ $X2=8.05 $Y2=1.085
r170 36 55 7.7488 $w=1.78e-07 $l=1.25e-07 $layer=LI1_cond $X=7.715 $Y=1.085
+ $X2=7.59 $Y2=1.085
r171 36 38 5.856 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=7.715 $Y=0.995
+ $X2=7.715 $Y2=0.875
r172 32 40 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.965 $Y=1.97
+ $X2=8.05 $Y2=1.845
r173 32 34 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=7.965 $Y=1.97
+ $X2=7.505 $Y2=1.97
r174 31 55 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.61 $Y=1.09
+ $X2=7.59 $Y2=1.09
r175 29 60 37.1502 $w=2.53e-07 $l=1.95e-07 $layer=POLY_cond $X=6.445 $Y=1.32
+ $X2=6.64 $Y2=1.32
r176 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.445
+ $Y=1.32 $X2=6.445 $Y2=1.32
r177 25 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.445 $Y=1.175
+ $X2=6.61 $Y2=1.09
r178 25 28 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.445 $Y=1.175
+ $X2=6.445 $Y2=1.32
r179 23 24 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=6.085 $Y=1.745
+ $X2=6.085 $Y2=1.895
r180 19 60 14.9957 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.64 $Y=1.155
+ $X2=6.64 $Y2=1.32
r181 19 21 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.64 $Y=1.155
+ $X2=6.64 $Y2=0.805
r182 17 29 60.9644 $w=2.53e-07 $l=3.93954e-07 $layer=POLY_cond $X=6.125 $Y=1.485
+ $X2=6.445 $Y2=1.32
r183 17 23 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=6.125 $Y=1.485
+ $X2=6.125 $Y2=1.745
r184 15 24 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.955 $Y=2.33
+ $X2=5.955 $Y2=1.895
r185 4 51 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=10.705
+ $Y=1.985 $X2=10.845 $Y2=2.18
r186 3 34 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.36
+ $Y=1.865 $X2=7.505 $Y2=2.01
r187 2 46 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=9.23
+ $Y=0.625 $X2=9.365 $Y2=0.77
r188 1 38 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=7.62
+ $Y=0.595 $X2=7.755 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_999_424# 1 2 3 12 14 16 18 19 22 23 25
+ 32 34 40
c95 12 0 1.43917e-19 $X=7.72 $Y=2.285
r96 34 36 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=1.1
+ $X2=5.465 $Y2=1.265
r97 31 32 5.76029 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=5.47 $Y=2.26
+ $X2=5.555 $Y2=2.26
r98 29 31 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=5.35 $Y=2.26
+ $X2=5.47 $Y2=2.26
r99 26 40 17.2143 $w=2.52e-07 $l=9e-08 $layer=POLY_cond $X=7.63 $Y=1.51 $X2=7.72
+ $Y2=1.51
r100 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.63
+ $Y=1.51 $X2=7.63 $Y2=1.51
r101 23 25 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=7.11 $Y=1.51
+ $X2=7.63 $Y2=1.51
r102 22 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.945 $Y=2.09
+ $X2=6.945 $Y2=2.175
r103 21 23 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=6.945 $Y=1.675
+ $X2=7.11 $Y2=1.51
r104 21 22 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=6.945 $Y=1.675
+ $X2=6.945 $Y2=2.09
r105 19 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=2.175
+ $X2=6.945 $Y2=2.175
r106 19 32 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=6.78 $Y=2.175
+ $X2=5.555 $Y2=2.175
r107 18 31 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.47 $Y=2.09
+ $X2=5.47 $Y2=2.26
r108 18 36 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.47 $Y=2.09
+ $X2=5.47 $Y2=1.265
r109 14 40 47.8175 $w=2.52e-07 $l=3.22102e-07 $layer=POLY_cond $X=7.97 $Y=1.345
+ $X2=7.72 $Y2=1.51
r110 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.97 $Y=1.345
+ $X2=7.97 $Y2=0.915
r111 10 40 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.72 $Y=1.675
+ $X2=7.72 $Y2=1.51
r112 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.72 $Y=1.675
+ $X2=7.72 $Y2=2.285
r113 3 38 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=6.69
+ $Y=2.12 $X2=6.945 $Y2=2.095
r114 2 29 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=4.995
+ $Y=2.12 $X2=5.35 $Y2=2.265
r115 1 34 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=5.25
+ $Y=0.825 $X2=5.46 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_2176_99# 1 2 7 9 10 12 15 21 23 24 25
+ 27 28 31 33 34 35 38 41 44 48
r123 45 48 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=15.73 $Y=2.055
+ $X2=15.915 $Y2=2.055
r124 44 52 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=14.79 $Y=1.445
+ $X2=14.545 $Y2=1.445
r125 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.79
+ $Y=1.445 $X2=14.79 $Y2=1.445
r126 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.265
+ $Y=1.32 $X2=11.265 $Y2=1.32
r127 38 45 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.73 $Y=1.93
+ $X2=15.73 $Y2=2.055
r128 37 38 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=15.73 $Y=1.61
+ $X2=15.73 $Y2=1.93
r129 36 43 4.03884 $w=1.7e-07 $l=1.65227e-07 $layer=LI1_cond $X=14.955 $Y=1.525
+ $X2=14.825 $Y2=1.445
r130 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.645 $Y=1.525
+ $X2=15.73 $Y2=1.61
r131 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=15.645 $Y=1.525
+ $X2=14.955 $Y2=1.525
r132 33 43 3.17338 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=14.825 $Y=1.61
+ $X2=14.825 $Y2=1.445
r133 33 34 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=14.825 $Y=1.61
+ $X2=14.825 $Y2=2.01
r134 29 31 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=12.07 $Y=1.155
+ $X2=12.07 $Y2=0.805
r135 27 34 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=14.695 $Y=2.095
+ $X2=14.825 $Y2=2.01
r136 27 28 213.011 $w=1.68e-07 $l=3.265e-06 $layer=LI1_cond $X=14.695 $Y=2.095
+ $X2=11.43 $Y2=2.095
r137 26 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.43 $Y=1.24
+ $X2=11.265 $Y2=1.24
r138 25 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.905 $Y=1.24
+ $X2=12.07 $Y2=1.155
r139 25 26 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=11.905 $Y=1.24
+ $X2=11.43 $Y2=1.24
r140 24 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.265 $Y=2.01
+ $X2=11.43 $Y2=2.095
r141 23 40 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.265 $Y=1.325
+ $X2=11.265 $Y2=1.24
r142 23 24 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=11.265 $Y=1.325
+ $X2=11.265 $Y2=2.01
r143 20 41 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=11.265 $Y=1.305
+ $X2=11.265 $Y2=1.32
r144 20 21 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=11.265 $Y=1.23
+ $X2=11.315 $Y2=1.23
r145 17 20 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=10.955 $Y=1.23
+ $X2=11.265 $Y2=1.23
r146 13 52 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.545 $Y=1.61
+ $X2=14.545 $Y2=1.445
r147 13 15 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=14.545 $Y=1.61
+ $X2=14.545 $Y2=2.45
r148 10 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.315 $Y=1.155
+ $X2=11.315 $Y2=1.23
r149 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.315 $Y=1.155
+ $X2=11.315 $Y2=0.835
r150 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.955 $Y=1.155
+ $X2=10.955 $Y2=1.23
r151 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.955 $Y=1.155
+ $X2=10.955 $Y2=0.835
r152 2 48 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.775
+ $Y=1.95 $X2=15.915 $Y2=2.095
r153 1 31 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=11.935
+ $Y=0.595 $X2=12.07 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_1098_271# 1 2 10 11 13 14 15 19 20 24
+ 29 30 31 32 36 41 42 45 48 52 54 55 56 57 58 61 62 63 66 68 69 70 75 77 78
c227 62 0 4.89312e-20 $X=16.105 $Y=1.025
c228 52 0 1.33414e-19 $X=8.505 $Y=1.98
c229 48 0 6.30553e-20 $X=5.675 $Y=1.43
c230 31 0 9.57414e-20 $X=10.345 $Y=1.8
c231 29 0 1.3677e-19 $X=10.27 $Y=2.405
r232 78 85 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.805 $Y=1.675
+ $X2=11.805 $Y2=1.84
r233 77 80 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=11.805 $Y=1.675
+ $X2=11.805 $Y2=1.755
r234 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.805
+ $Y=1.675 $X2=11.805 $Y2=1.675
r235 74 75 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=17.41 $Y=1.29
+ $X2=17.41 $Y2=2.01
r236 70 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.325 $Y=2.095
+ $X2=17.41 $Y2=2.01
r237 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=17.325 $Y=2.095
+ $X2=17.02 $Y2=2.095
r238 68 74 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.325 $Y=1.205
+ $X2=17.41 $Y2=1.29
r239 68 69 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=17.325 $Y=1.205
+ $X2=16.76 $Y2=1.205
r240 64 69 27.9399 $w=2.19e-07 $l=5.33104e-07 $layer=LI1_cond $X=16.27 $Y=1.115
+ $X2=16.76 $Y2=1.205
r241 64 66 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=16.27 $Y=0.94
+ $X2=16.27 $Y2=0.76
r242 62 64 9.83486 $w=2.19e-07 $l=2.05122e-07 $layer=LI1_cond $X=16.105 $Y=1.025
+ $X2=16.27 $Y2=1.115
r243 62 63 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=16.105 $Y=1.025
+ $X2=14.525 $Y2=1.025
r244 60 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.44 $Y=1.11
+ $X2=14.525 $Y2=1.025
r245 60 61 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=14.44 $Y=1.11
+ $X2=14.44 $Y2=1.67
r246 59 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.97 $Y=1.755
+ $X2=11.805 $Y2=1.755
r247 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.355 $Y=1.755
+ $X2=14.44 $Y2=1.67
r248 58 59 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=14.355 $Y=1.755
+ $X2=11.97 $Y2=1.755
r249 50 52 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=8.345 $Y=1.98
+ $X2=8.505 $Y2=1.98
r250 46 48 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=5.565 $Y=1.43
+ $X2=5.675 $Y2=1.43
r251 45 85 633.266 $w=1.5e-07 $l=1.235e-06 $layer=POLY_cond $X=11.715 $Y=3.075
+ $X2=11.715 $Y2=1.84
r252 43 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.705 $Y=3.15
+ $X2=10.63 $Y2=3.15
r253 42 45 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.64 $Y=3.15
+ $X2=11.715 $Y2=3.075
r254 42 43 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=11.64 $Y=3.15
+ $X2=10.705 $Y2=3.15
r255 39 57 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.63 $Y=3.075
+ $X2=10.63 $Y2=3.15
r256 39 41 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=10.63 $Y=3.075
+ $X2=10.63 $Y2=2.405
r257 38 56 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=10.63 $Y=1.875
+ $X2=10.612 $Y2=1.8
r258 38 41 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.63 $Y=1.875
+ $X2=10.63 $Y2=2.405
r259 34 56 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=10.595 $Y=1.725
+ $X2=10.612 $Y2=1.8
r260 34 36 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=10.595 $Y=1.725
+ $X2=10.595 $Y2=0.835
r261 33 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.345 $Y=3.15
+ $X2=10.27 $Y2=3.15
r262 32 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.555 $Y=3.15
+ $X2=10.63 $Y2=3.15
r263 32 33 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.555 $Y=3.15
+ $X2=10.345 $Y2=3.15
r264 30 56 5.30422 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=10.52 $Y=1.8
+ $X2=10.612 $Y2=1.8
r265 30 31 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=10.52 $Y=1.8
+ $X2=10.345 $Y2=1.8
r266 27 55 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.27 $Y=3.075
+ $X2=10.27 $Y2=3.15
r267 27 29 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=10.27 $Y=3.075
+ $X2=10.27 $Y2=2.405
r268 26 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.27 $Y=1.875
+ $X2=10.345 $Y2=1.8
r269 26 29 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.27 $Y=1.875
+ $X2=10.27 $Y2=2.405
r270 22 52 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.505 $Y=1.905
+ $X2=8.505 $Y2=1.98
r271 22 24 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=8.505 $Y=1.905
+ $X2=8.505 $Y2=1.025
r272 21 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.42 $Y=3.15
+ $X2=8.345 $Y2=3.15
r273 20 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.195 $Y=3.15
+ $X2=10.27 $Y2=3.15
r274 20 21 910.16 $w=1.5e-07 $l=1.775e-06 $layer=POLY_cond $X=10.195 $Y=3.15
+ $X2=8.42 $Y2=3.15
r275 17 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.345 $Y=3.075
+ $X2=8.345 $Y2=3.15
r276 17 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.345 $Y=3.075
+ $X2=8.345 $Y2=2.485
r277 16 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.345 $Y=2.055
+ $X2=8.345 $Y2=1.98
r278 16 19 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.345 $Y=2.055
+ $X2=8.345 $Y2=2.485
r279 14 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.27 $Y=3.15
+ $X2=8.345 $Y2=3.15
r280 14 15 1348.57 $w=1.5e-07 $l=2.63e-06 $layer=POLY_cond $X=8.27 $Y=3.15
+ $X2=5.64 $Y2=3.15
r281 11 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.675 $Y=1.355
+ $X2=5.675 $Y2=1.43
r282 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.675 $Y=1.355
+ $X2=5.675 $Y2=1.035
r283 8 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.565 $Y=3.075
+ $X2=5.64 $Y2=3.15
r284 8 10 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=5.565 $Y=3.075
+ $X2=5.565 $Y2=2.33
r285 7 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.565 $Y=1.505
+ $X2=5.565 $Y2=1.43
r286 7 10 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=5.565 $Y=1.505
+ $X2=5.565 $Y2=2.33
r287 2 72 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=16.85
+ $Y=1.95 $X2=17.02 $Y2=2.095
r288 1 66 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=16.125
+ $Y=0.485 $X2=16.27 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_1982_397# 1 2 3 12 16 20 24 28 32 34 36
+ 40 42 45 46 49 51 55 59 62 65 67 69 71 72
c198 59 0 8.2015e-20 $X=12.375 $Y=2.515
c199 49 0 1.20173e-19 $X=19.24 $Y=2.35
c200 34 0 1.3677e-19 $X=12.21 $Y=2.65
c201 28 0 5.48677e-20 $X=19.185 $Y=0.575
c202 20 0 4.39729e-20 $X=16.18 $Y=2.45
r203 72 83 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=19.207 $Y=1.48
+ $X2=19.207 $Y2=1.645
r204 72 82 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=19.207 $Y=1.48
+ $X2=19.207 $Y2=1.315
r205 71 74 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=19.21 $Y=1.48
+ $X2=19.21 $Y2=1.645
r206 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=19.21
+ $Y=1.48 $X2=19.21 $Y2=1.48
r207 65 80 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=16.15 $Y=1.575
+ $X2=16.15 $Y2=1.74
r208 64 67 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=16.15 $Y=1.575
+ $X2=16.335 $Y2=1.575
r209 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.15
+ $Y=1.575 $X2=16.15 $Y2=1.575
r210 59 75 16.3083 $w=2.66e-07 $l=9e-08 $layer=POLY_cond $X=12.375 $Y=2.515
+ $X2=12.285 $Y2=2.515
r211 58 60 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=12.375 $Y=2.515
+ $X2=12.375 $Y2=2.65
r212 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.375
+ $Y=2.515 $X2=12.375 $Y2=2.515
r213 55 58 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=12.375 $Y=2.435
+ $X2=12.375 $Y2=2.515
r214 51 53 10.1961 $w=6.08e-07 $l=5.2e-07 $layer=LI1_cond $X=10.195 $Y=2.13
+ $X2=10.195 $Y2=2.65
r215 51 52 4.65126 $w=6.08e-07 $l=9e-08 $layer=LI1_cond $X=10.195 $Y=2.13
+ $X2=10.195 $Y2=2.04
r216 49 74 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=19.24 $Y=2.35
+ $X2=19.24 $Y2=1.645
r217 47 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.42 $Y=2.435
+ $X2=16.335 $Y2=2.435
r218 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=19.155 $Y=2.435
+ $X2=19.24 $Y2=2.35
r219 46 47 178.433 $w=1.68e-07 $l=2.735e-06 $layer=LI1_cond $X=19.155 $Y=2.435
+ $X2=16.42 $Y2=2.435
r220 45 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.335 $Y=2.35
+ $X2=16.335 $Y2=2.435
r221 44 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.335 $Y=1.74
+ $X2=16.335 $Y2=1.575
r222 44 45 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=16.335 $Y=1.74
+ $X2=16.335 $Y2=2.35
r223 43 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.955 $Y=2.435
+ $X2=13.79 $Y2=2.435
r224 42 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.25 $Y=2.435
+ $X2=16.335 $Y2=2.435
r225 42 43 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=16.25 $Y=2.435
+ $X2=13.955 $Y2=2.435
r226 38 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.79 $Y=2.52
+ $X2=13.79 $Y2=2.435
r227 38 40 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=13.79 $Y=2.52
+ $X2=13.79 $Y2=2.66
r228 37 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.54 $Y=2.435
+ $X2=12.375 $Y2=2.435
r229 36 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.625 $Y=2.435
+ $X2=13.79 $Y2=2.435
r230 36 37 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=13.625 $Y=2.435
+ $X2=12.54 $Y2=2.435
r231 35 53 8.42348 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=10.5 $Y=2.65
+ $X2=10.195 $Y2=2.65
r232 34 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.21 $Y=2.65
+ $X2=12.375 $Y2=2.65
r233 34 35 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=12.21 $Y=2.65
+ $X2=10.5 $Y2=2.65
r234 32 52 47.213 $w=3.08e-07 $l=1.27e-06 $layer=LI1_cond $X=10.345 $Y=0.77
+ $X2=10.345 $Y2=2.04
r235 28 82 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=19.185 $Y=0.575
+ $X2=19.185 $Y2=1.315
r236 24 83 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=19.115 $Y=2.155
+ $X2=19.115 $Y2=1.645
r237 20 80 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=16.18 $Y=2.45
+ $X2=16.18 $Y2=1.74
r238 14 59 48.9248 $w=2.66e-07 $l=3.4271e-07 $layer=POLY_cond $X=12.645 $Y=2.35
+ $X2=12.375 $Y2=2.515
r239 14 16 792.223 $w=1.5e-07 $l=1.545e-06 $layer=POLY_cond $X=12.645 $Y=2.35
+ $X2=12.645 $Y2=0.805
r240 10 75 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.285 $Y=2.35
+ $X2=12.285 $Y2=2.515
r241 10 12 792.223 $w=1.5e-07 $l=1.545e-06 $layer=POLY_cond $X=12.285 $Y=2.35
+ $X2=12.285 $Y2=0.805
r242 3 40 600 $w=1.7e-07 $l=7.79134e-07 $layer=licon1_PDIFF $count=1 $X=13.645
+ $Y=1.95 $X2=13.79 $Y2=2.66
r243 2 51 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.91
+ $Y=1.985 $X2=10.055 $Y2=2.13
r244 1 32 91 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=2 $X=10.015
+ $Y=0.625 $X2=10.275 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_2586_249# 1 2 9 11 13 16 17 20 23 24 25
+ 27 28 29 31 32 33 35 38 42 43 47
r152 44 47 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=17.98 $Y=2.015
+ $X2=18.325 $Y2=2.015
r153 42 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.15 $Y=0.63
+ $X2=15.15 $Y2=0.795
r154 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.15
+ $Y=0.63 $X2=15.15 $Y2=0.63
r155 36 43 3.70735 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=18.18 $Y=0.78
+ $X2=18.12 $Y2=0.865
r156 36 38 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=18.18 $Y=0.78
+ $X2=18.18 $Y2=0.575
r157 35 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.98 $Y=1.85
+ $X2=17.98 $Y2=2.015
r158 34 43 3.70735 $w=2.5e-07 $l=1.77482e-07 $layer=LI1_cond $X=17.98 $Y=0.95
+ $X2=18.12 $Y2=0.865
r159 34 35 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=17.98 $Y=0.95
+ $X2=17.98 $Y2=1.85
r160 32 43 2.76166 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=17.895 $Y=0.865
+ $X2=18.12 $Y2=0.865
r161 32 33 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=17.895 $Y=0.865
+ $X2=17.1 $Y2=0.865
r162 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.015 $Y=0.78
+ $X2=17.1 $Y2=0.865
r163 30 31 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=17.015 $Y=0.425
+ $X2=17.015 $Y2=0.78
r164 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=16.93 $Y=0.34
+ $X2=17.015 $Y2=0.425
r165 28 29 105.364 $w=1.68e-07 $l=1.615e-06 $layer=LI1_cond $X=16.93 $Y=0.34
+ $X2=15.315 $Y2=0.34
r166 27 41 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.15 $Y=0.6
+ $X2=15.15 $Y2=0.685
r167 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=15.15 $Y=0.425
+ $X2=15.315 $Y2=0.34
r168 26 27 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=15.15 $Y=0.425
+ $X2=15.15 $Y2=0.6
r169 24 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.985 $Y=0.685
+ $X2=15.15 $Y2=0.685
r170 24 25 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=14.985 $Y=0.685
+ $X2=14.185 $Y2=0.685
r171 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.1 $Y=0.77
+ $X2=14.185 $Y2=0.685
r172 22 23 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=14.1 $Y=0.77
+ $X2=14.1 $Y2=1.32
r173 20 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.095 $Y=1.41
+ $X2=13.095 $Y2=1.245
r174 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.095
+ $Y=1.41 $X2=13.095 $Y2=1.41
r175 17 23 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=14.015 $Y=1.41
+ $X2=14.1 $Y2=1.32
r176 17 19 56.6869 $w=1.78e-07 $l=9.2e-07 $layer=LI1_cond $X=14.015 $Y=1.41
+ $X2=13.095 $Y2=1.41
r177 16 54 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=15.24 $Y=1.82
+ $X2=15.24 $Y2=0.795
r178 11 16 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=15.19 $Y=1.945
+ $X2=15.19 $Y2=1.82
r179 11 13 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=15.19 $Y=1.945
+ $X2=15.19 $Y2=2.45
r180 9 50 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=13.075 $Y=0.805
+ $X2=13.075 $Y2=1.245
r181 2 47 600 $w=1.7e-07 $l=2.85657e-07 $layer=licon1_PDIFF $count=1 $X=18.07
+ $Y=1.95 $X2=18.325 $Y2=2.015
r182 1 38 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=18.045
+ $Y=0.365 $X2=18.18 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%RESET_B 3 7 10 11 12 15 17 18 22 24 25 29
+ 31 33 35 39 41 42 43 44 50
c167 50 0 1.01483e-19 $X=4.375 $Y=1.715
c168 31 0 4.89312e-20 $X=15.625 $Y=0.18
c169 17 0 1.40585e-19 $X=6.955 $Y=1.8
r170 48 50 47.223 $w=2.96e-07 $l=2.9e-07 $layer=POLY_cond $X=4.085 $Y=1.715
+ $X2=4.375 $Y2=1.715
r171 46 48 14.6554 $w=2.96e-07 $l=9e-08 $layer=POLY_cond $X=3.995 $Y=1.715
+ $X2=4.085 $Y2=1.715
r172 44 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.085
+ $Y=1.715 $X2=4.085 $Y2=1.715
r173 40 41 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=7.015 $Y=1.125
+ $X2=7.015 $Y2=1.275
r174 37 43 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=15.7 $Y=0.255
+ $X2=15.7 $Y2=1.035
r175 33 43 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=15.65 $Y=1.16
+ $X2=15.65 $Y2=1.035
r176 33 35 320.505 $w=2.5e-07 $l=1.29e-06 $layer=POLY_cond $X=15.65 $Y=1.16
+ $X2=15.65 $Y2=2.45
r177 32 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.62 $Y=0.18
+ $X2=13.545 $Y2=0.18
r178 31 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.625 $Y=0.18
+ $X2=15.7 $Y2=0.255
r179 31 32 1028.1 $w=1.5e-07 $l=2.005e-06 $layer=POLY_cond $X=15.625 $Y=0.18
+ $X2=13.62 $Y2=0.18
r180 27 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.545 $Y=0.255
+ $X2=13.545 $Y2=0.18
r181 27 29 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=13.545 $Y=0.255
+ $X2=13.545 $Y2=0.805
r182 26 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.075 $Y=0.18 $X2=7
+ $Y2=0.18
r183 25 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.47 $Y=0.18
+ $X2=13.545 $Y2=0.18
r184 25 26 3279.14 $w=1.5e-07 $l=6.395e-06 $layer=POLY_cond $X=13.47 $Y=0.18
+ $X2=7.075 $Y2=0.18
r185 24 41 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.03 $Y=1.725
+ $X2=7.03 $Y2=1.275
r186 22 40 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7 $Y=0.805 $X2=7
+ $Y2=1.125
r187 19 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7 $Y=0.255 $X2=7
+ $Y2=0.18
r188 19 22 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7 $Y=0.255 $X2=7
+ $Y2=0.805
r189 17 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.955 $Y=1.8
+ $X2=7.03 $Y2=1.725
r190 17 18 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=6.955 $Y=1.8
+ $X2=6.69 $Y2=1.8
r191 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.615 $Y=1.875
+ $X2=6.69 $Y2=1.8
r192 13 15 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.615 $Y=1.875
+ $X2=6.615 $Y2=2.33
r193 11 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.925 $Y=0.18 $X2=7
+ $Y2=0.18
r194 11 12 1207.56 $w=1.5e-07 $l=2.355e-06 $layer=POLY_cond $X=6.925 $Y=0.18
+ $X2=4.57 $Y2=0.18
r195 10 50 19.5405 $w=2.96e-07 $l=2.16852e-07 $layer=POLY_cond $X=4.495 $Y=1.55
+ $X2=4.375 $Y2=1.715
r196 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.495 $Y=0.255
+ $X2=4.57 $Y2=0.18
r197 9 10 664.032 $w=1.5e-07 $l=1.295e-06 $layer=POLY_cond $X=4.495 $Y=0.255
+ $X2=4.495 $Y2=1.55
r198 5 50 18.6531 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.88
+ $X2=4.375 $Y2=1.715
r199 5 7 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=4.375 $Y=1.88
+ $X2=4.375 $Y2=2.65
r200 1 46 18.6531 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.55
+ $X2=3.995 $Y2=1.715
r201 1 3 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.995 $Y=1.55
+ $X2=3.995 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%CLK 3 7 9 12
c44 9 0 4.39729e-20 $X=17.04 $Y=1.665
r45 12 15 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=16.722 $Y=1.625
+ $X2=16.722 $Y2=1.79
r46 12 14 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=16.722 $Y=1.625
+ $X2=16.722 $Y2=1.46
r47 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.755
+ $Y=1.625 $X2=16.755 $Y2=1.625
r48 9 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=17.04 $Y=1.625
+ $X2=16.755 $Y2=1.625
r49 7 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=16.775 $Y=2.27
+ $X2=16.775 $Y2=1.79
r50 3 14 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=16.6 $Y=0.695
+ $X2=16.6 $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%SLEEP_B 1 3 6 8 10 11 12 15 17 19 23 27
+ 32 33 34 38
c90 34 0 5.48677e-20 $X=18.48 $Y=1.295
r91 36 38 0.730303 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=18.395 $Y=1.187
+ $X2=18.4 $Y2=1.187
r92 34 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.4
+ $Y=1.285 $X2=18.4 $Y2=1.285
r93 30 31 14.5801 $w=2.81e-07 $l=8.5e-08 $layer=POLY_cond $X=17.235 $Y=1.307
+ $X2=17.32 $Y2=1.307
r94 25 38 51.8515 $w=3.3e-07 $l=4.68012e-07 $layer=POLY_cond $X=18.755 $Y=0.925
+ $X2=18.4 $Y2=1.187
r95 25 27 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=18.755 $Y=0.925
+ $X2=18.755 $Y2=0.575
r96 21 36 21.2229 $w=1.5e-07 $l=2.62e-07 $layer=POLY_cond $X=18.395 $Y=0.925
+ $X2=18.395 $Y2=1.187
r97 21 23 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=18.395 $Y=0.925
+ $X2=18.395 $Y2=0.575
r98 20 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.97 $Y=1.375
+ $X2=17.895 $Y2=1.375
r99 19 36 37.8699 $w=3.3e-07 $l=2.55781e-07 $layer=POLY_cond $X=18.235 $Y=1.375
+ $X2=18.395 $Y2=1.187
r100 19 20 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=18.235 $Y=1.375
+ $X2=17.97 $Y2=1.375
r101 15 33 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=17.945 $Y=1.815
+ $X2=17.945 $Y2=1.69
r102 15 17 157.768 $w=2.5e-07 $l=6.35e-07 $layer=POLY_cond $X=17.945 $Y=1.815
+ $X2=17.945 $Y2=2.45
r103 13 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.895 $Y=1.45
+ $X2=17.895 $Y2=1.375
r104 13 33 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=17.895 $Y=1.45
+ $X2=17.895 $Y2=1.69
r105 12 31 23.2782 $w=2.81e-07 $l=1.03562e-07 $layer=POLY_cond $X=17.395
+ $Y=1.375 $X2=17.32 $Y2=1.307
r106 11 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.82 $Y=1.375
+ $X2=17.895 $Y2=1.375
r107 11 12 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=17.82 $Y=1.375
+ $X2=17.395 $Y2=1.375
r108 8 31 17.4353 $w=1.5e-07 $l=2.92e-07 $layer=POLY_cond $X=17.32 $Y=1.015
+ $X2=17.32 $Y2=1.307
r109 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=17.32 $Y=1.015
+ $X2=17.32 $Y2=0.695
r110 4 30 17.4353 $w=1.5e-07 $l=1.43e-07 $layer=POLY_cond $X=17.235 $Y=1.45
+ $X2=17.235 $Y2=1.307
r111 4 6 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=17.235 $Y=1.45
+ $X2=17.235 $Y2=2.27
r112 1 30 47.1708 $w=2.81e-07 $l=4.06896e-07 $layer=POLY_cond $X=16.96 $Y=1.015
+ $X2=17.235 $Y2=1.307
r113 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=16.96 $Y=1.015
+ $X2=16.96 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_3751_367# 1 2 9 13 17 18 21 24 26 27 29
+ 33 37
r72 34 37 16.6846 $w=2.6e-07 $l=9e-08 $layer=POLY_cond $X=19.855 $Y=1.48
+ $X2=19.945 $Y2=1.48
r73 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=19.855
+ $Y=1.48 $X2=19.855 $Y2=1.48
r74 30 33 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=19.6 $Y=1.48
+ $X2=19.855 $Y2=1.48
r75 26 27 9.48474 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=18.86 $Y=1.995
+ $X2=18.86 $Y2=1.815
r76 24 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.6 $Y=1.315
+ $X2=19.6 $Y2=1.48
r77 23 29 3.05675 $w=3.1e-07 $l=1.77482e-07 $layer=LI1_cond $X=19.6 $Y=1.145
+ $X2=19.46 $Y2=1.06
r78 23 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=19.6 $Y=1.145
+ $X2=19.6 $Y2=1.315
r79 19 29 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=19.46 $Y=0.975
+ $X2=19.46 $Y2=1.06
r80 19 21 10.6318 $w=4.48e-07 $l=4e-07 $layer=LI1_cond $X=19.46 $Y=0.975
+ $X2=19.46 $Y2=0.575
r81 17 29 3.57226 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=19.235 $Y=1.06
+ $X2=19.46 $Y2=1.06
r82 17 18 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=19.235 $Y=1.06
+ $X2=18.905 $Y2=1.06
r83 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=18.82 $Y=1.145
+ $X2=18.905 $Y2=1.06
r84 15 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=18.82 $Y=1.145
+ $X2=18.82 $Y2=1.815
r85 11 37 38.9308 $w=2.6e-07 $l=2.80624e-07 $layer=POLY_cond $X=20.155 $Y=1.315
+ $X2=19.945 $Y2=1.48
r86 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=20.155 $Y=1.315
+ $X2=20.155 $Y2=0.705
r87 7 37 15.628 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=19.945 $Y=1.645
+ $X2=19.945 $Y2=1.48
r88 7 9 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=19.945 $Y=1.645
+ $X2=19.945 $Y2=2.465
r89 2 26 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=18.755
+ $Y=1.835 $X2=18.9 $Y2=1.995
r90 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=19.26
+ $Y=0.365 $X2=19.4 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%VPWR 1 2 3 4 5 18 22 26 30 34 39 40 42 43
+ 45 46 47 49 67 79 80 83 86 100
c144 80 0 1.43917e-19 $X=20.4 $Y=3.33
c145 1 0 1.4905e-19 $X=0.64 $Y=2.33
r146 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r147 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r148 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.4 $Y=3.33
+ $X2=20.4 $Y2=3.33
r149 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=19.44 $Y=3.33
+ $X2=20.4 $Y2=3.33
r150 77 100 2.47516 $w=4.9e-07 $l=8.88e-06 $layer=MET1_cond $X=19.44 $Y=3.33
+ $X2=10.56 $Y2=3.33
r151 76 77 0.775 $w=1.7e-07 $l=2.04e-06 $layer=mcon $count=12 $X=19.44 $Y=3.33
+ $X2=19.44 $Y2=3.33
r152 74 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r153 73 76 720.257 $w=1.68e-07 $l=1.104e-05 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=19.44 $Y2=3.33
r154 73 74 0.775 $w=1.7e-07 $l=2.04e-06 $layer=mcon $count=12 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 71 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.18 $Y=3.33
+ $X2=8.015 $Y2=3.33
r156 71 73 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.18 $Y=3.33
+ $X2=8.4 $Y2=3.33
r157 70 87 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r158 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r159 67 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.85 $Y=3.33
+ $X2=8.015 $Y2=3.33
r160 67 69 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=7.85 $Y=3.33
+ $X2=6.48 $Y2=3.33
r161 66 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r162 65 66 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r163 63 66 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r164 62 65 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r165 62 63 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r166 60 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r167 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r168 57 60 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r169 57 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r170 56 59 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r171 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r172 54 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.785 $Y2=3.33
r173 54 56 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=1.2 $Y2=3.33
r174 52 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r175 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r176 49 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.785 $Y2=3.33
r177 49 51 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.24 $Y2=3.33
r178 47 100 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.56 $Y2=3.33
r179 47 74 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=8.4 $Y2=3.33
r180 45 76 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=19.495 $Y=3.33
+ $X2=19.44 $Y2=3.33
r181 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.495 $Y=3.33
+ $X2=19.66 $Y2=3.33
r182 44 79 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=19.825 $Y=3.33
+ $X2=20.4 $Y2=3.33
r183 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.825 $Y=3.33
+ $X2=19.66 $Y2=3.33
r184 42 65 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.12 $Y=3.33 $X2=6
+ $Y2=3.33
r185 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.12 $Y=3.33
+ $X2=6.285 $Y2=3.33
r186 41 69 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=6.45 $Y=3.33 $X2=6.48
+ $Y2=3.33
r187 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.45 $Y=3.33
+ $X2=6.285 $Y2=3.33
r188 39 59 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.12 $Y2=3.33
r189 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.41 $Y2=3.33
r190 38 62 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=3.6 $Y2=3.33
r191 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=3.41 $Y2=3.33
r192 34 37 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=19.66 $Y=1.98
+ $X2=19.66 $Y2=2.465
r193 32 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.66 $Y=3.245
+ $X2=19.66 $Y2=3.33
r194 32 37 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=19.66 $Y=3.245
+ $X2=19.66 $Y2=2.465
r195 28 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=3.245
+ $X2=8.015 $Y2=3.33
r196 28 30 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=8.015 $Y=3.245
+ $X2=8.015 $Y2=2.77
r197 24 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.285 $Y=3.245
+ $X2=6.285 $Y2=3.33
r198 24 26 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.285 $Y=3.245
+ $X2=6.285 $Y2=2.855
r199 20 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=3.245
+ $X2=3.41 $Y2=3.33
r200 20 22 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.41 $Y=3.245
+ $X2=3.41 $Y2=2.715
r201 16 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r202 16 18 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.665
r203 5 37 300 $w=1.7e-07 $l=8.32466e-07 $layer=licon1_PDIFF $count=2 $X=19.19
+ $Y=1.835 $X2=19.66 $Y2=2.465
r204 5 34 600 $w=1.7e-07 $l=5.37634e-07 $layer=licon1_PDIFF $count=1 $X=19.19
+ $Y=1.835 $X2=19.66 $Y2=1.98
r205 4 30 600 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.865 $X2=8.015 $Y2=2.77
r206 3 26 600 $w=1.7e-07 $l=8.53024e-07 $layer=licon1_PDIFF $count=1 $X=6.03
+ $Y=2.12 $X2=6.285 $Y2=2.855
r207 2 22 600 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=2.33 $X2=3.41 $Y2=2.715
r208 1 18 600 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=2.33 $X2=0.785 $Y2=2.665
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_332_136# 1 2 3 4 14 15 16 17 18 21 25
+ 29 32 33 34 36 37 38 41 43 47 48
c133 33 0 6.30553e-20 $X=5.035 $Y=1.335
c134 16 0 1.73039e-19 $X=1.395 $Y=1.585
c135 14 0 1.4905e-19 $X=1.31 $Y=2.34
r136 45 47 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.47 $Y=2.425
+ $X2=2.47 $Y2=2.475
r137 43 45 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.47 $Y=2.185
+ $X2=2.47 $Y2=2.425
r138 39 41 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=5.89 $Y=0.765
+ $X2=5.89 $Y2=1.035
r139 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.725 $Y=0.68
+ $X2=5.89 $Y2=0.765
r140 37 38 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.725 $Y=0.68
+ $X2=5.205 $Y2=0.68
r141 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.12 $Y=0.765
+ $X2=5.205 $Y2=0.68
r142 35 36 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.12 $Y=0.765
+ $X2=5.12 $Y2=1.25
r143 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.035 $Y=1.335
+ $X2=5.12 $Y2=1.25
r144 33 34 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.035 $Y=1.335
+ $X2=4.715 $Y2=1.335
r145 32 48 3.70735 $w=2.5e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.63 $Y=2.1
+ $X2=4.59 $Y2=2.185
r146 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.63 $Y=1.42
+ $X2=4.715 $Y2=1.335
r147 31 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.63 $Y=1.42
+ $X2=4.63 $Y2=2.1
r148 27 48 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=2.27
+ $X2=4.59 $Y2=2.185
r149 27 29 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.59 $Y=2.27
+ $X2=4.59 $Y2=2.475
r150 26 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=2.185
+ $X2=2.47 $Y2=2.185
r151 25 48 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=2.185
+ $X2=4.59 $Y2=2.185
r152 25 26 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=4.425 $Y=2.185
+ $X2=2.635 $Y2=2.185
r153 19 21 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=1.955 $Y=1.5
+ $X2=1.955 $Y2=1.1
r154 17 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=2.425
+ $X2=2.47 $Y2=2.425
r155 17 18 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.305 $Y=2.425
+ $X2=1.395 $Y2=2.425
r156 15 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.83 $Y=1.585
+ $X2=1.955 $Y2=1.5
r157 15 16 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.83 $Y=1.585
+ $X2=1.395 $Y2=1.585
r158 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.31 $Y=2.34
+ $X2=1.395 $Y2=2.425
r159 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.31 $Y=1.67
+ $X2=1.395 $Y2=1.585
r160 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.31 $Y=1.67
+ $X2=1.31 $Y2=2.34
r161 4 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.45
+ $Y=2.33 $X2=4.59 $Y2=2.475
r162 3 47 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.955
+ $Y=2.33 $X2=2.47 $Y2=2.475
r163 2 41 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.75
+ $Y=0.825 $X2=5.89 $Y2=1.035
r164 1 21 182 $w=1.7e-07 $l=5.32447e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.68 $X2=1.915 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%KAPWR 1 2 3 10 13 19 26 29 34
c122 26 0 8.2015e-20 $X=17.04 $Y=2.82
r123 25 29 18.0607 $w=3.33e-07 $l=5.25e-07 $layer=LI1_cond $X=17.04 $Y=2.857
+ $X2=17.565 $Y2=2.857
r124 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=2.82
+ $X2=17.04 $Y2=2.82
r125 22 26 0.262345 $w=2.7e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=2.81
+ $X2=17.04 $Y2=2.81
r126 19 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=2.82
+ $X2=16.56 $Y2=2.82
r127 14 22 1.04938 $w=2.7e-07 $l=1.92e-06 $layer=MET1_cond $X=14.64 $Y=2.81
+ $X2=16.56 $Y2=2.81
r128 14 34 2.22993 $w=2.7e-07 $l=4.08e-06 $layer=MET1_cond $X=14.64 $Y=2.81
+ $X2=10.56 $Y2=2.81
r129 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=2.82
+ $X2=14.64 $Y2=2.82
r130 10 34 0.131172 $w=2.7e-07 $l=2.4e-07 $layer=MET1_cond $X=10.32 $Y=2.81
+ $X2=10.56 $Y2=2.81
r131 3 29 600 $w=1.7e-07 $l=1.0246e-06 $layer=licon1_PDIFF $count=1 $X=17.31
+ $Y=1.95 $X2=17.565 $Y2=2.855
r132 2 19 600 $w=1.7e-07 $l=9.07304e-07 $layer=licon1_PDIFF $count=1 $X=16.305
+ $Y=1.95 $X2=16.445 $Y2=2.79
r133 1 13 600 $w=1.7e-07 $l=9.07304e-07 $layer=licon1_PDIFF $count=1 $X=14.67
+ $Y=1.95 $X2=14.81 $Y2=2.79
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%Q 1 2 9 11 12 13 14 15 23
c22 15 0 1.3383e-19 $X=20.4 $Y=2.035
r23 21 34 7.22427 $w=3.33e-07 $l=2.1e-07 $layer=LI1_cond $X=20.37 $Y=1.982
+ $X2=20.16 $Y2=1.982
r24 15 21 1.03204 $w=3.33e-07 $l=3e-08 $layer=LI1_cond $X=20.4 $Y=1.982
+ $X2=20.37 $Y2=1.982
r25 14 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=20.37 $Y=1.665
+ $X2=20.37 $Y2=1.815
r26 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=20.37 $Y=1.295
+ $X2=20.37 $Y2=1.665
r27 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=20.37 $Y=0.925
+ $X2=20.37 $Y2=1.295
r28 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=20.37 $Y=0.555
+ $X2=20.37 $Y2=0.925
r29 11 23 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=20.37 $Y=0.555
+ $X2=20.37 $Y2=0.43
r30 7 34 0.808037 $w=3.3e-07 $l=1.68e-07 $layer=LI1_cond $X=20.16 $Y=2.15
+ $X2=20.16 $Y2=1.982
r31 7 9 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=20.16 $Y=2.15
+ $X2=20.16 $Y2=2.91
r32 2 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=20.02
+ $Y=1.835 $X2=20.16 $Y2=1.98
r33 2 9 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=20.02
+ $Y=1.835 $X2=20.16 $Y2=2.91
r34 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=20.23
+ $Y=0.285 $X2=20.37 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50
+ 54 58 60 64 67 68 70 71 73 74 76 77 78 80 107 111 116 123 124 127 130 133 136
+ 139 151
c172 64 0 1.3383e-19 $X=19.94 $Y=0.43
r173 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.92 $Y=0
+ $X2=19.92 $Y2=0
r174 137 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=18.96 $Y=0
+ $X2=19.92 $Y2=0
r175 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.96 $Y=0
+ $X2=18.96 $Y2=0
r176 133 134 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r177 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r178 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r179 124 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=20.4 $Y=0
+ $X2=19.92 $Y2=0
r180 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.4 $Y=0
+ $X2=20.4 $Y2=0
r181 121 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.025 $Y=0
+ $X2=19.94 $Y2=0
r182 121 123 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=20.025 $Y=0
+ $X2=20.4 $Y2=0
r183 120 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=18.48 $Y=0
+ $X2=18.96 $Y2=0
r184 120 134 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=18.48 $Y=0
+ $X2=17.52 $Y2=0
r185 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.48 $Y=0
+ $X2=18.48 $Y2=0
r186 117 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.805 $Y=0
+ $X2=17.64 $Y2=0
r187 117 119 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=17.805 $Y=0
+ $X2=18.48 $Y2=0
r188 116 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=18.805 $Y=0
+ $X2=18.93 $Y2=0
r189 116 119 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=18.805 $Y=0
+ $X2=18.48 $Y2=0
r190 115 134 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=17.52 $Y2=0
r191 115 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r192 114 115 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r193 112 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.29 $Y2=0
r194 112 114 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.68 $Y2=0
r195 111 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.475 $Y=0
+ $X2=17.64 $Y2=0
r196 111 114 247.588 $w=1.68e-07 $l=3.795e-06 $layer=LI1_cond $X=17.475 $Y=0
+ $X2=13.68 $Y2=0
r197 110 131 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r198 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r199 107 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.125 $Y=0
+ $X2=13.29 $Y2=0
r200 107 109 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=13.125 $Y=0
+ $X2=11.76 $Y2=0
r201 106 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r202 105 106 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r203 103 151 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=10.08 $Y2=0
r204 102 105 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=8.4 $Y=0
+ $X2=11.28 $Y2=0
r205 102 103 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r206 100 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r207 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r208 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.92 $Y2=0
r209 96 97 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r210 94 97 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=6.96 $Y2=0
r211 93 96 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6.96
+ $Y2=0
r212 93 94 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r213 91 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r214 90 91 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r215 88 91 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r216 88 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r217 87 90 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r218 87 88 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r219 85 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.7
+ $Y2=0
r220 85 87 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r221 83 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r222 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r223 80 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.7
+ $Y2=0
r224 80 82 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r225 78 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r226 78 151 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.08 $Y2=0
r227 76 105 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=11.365 $Y=0
+ $X2=11.28 $Y2=0
r228 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.365 $Y=0
+ $X2=11.53 $Y2=0
r229 75 109 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=11.695 $Y=0
+ $X2=11.76 $Y2=0
r230 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.695 $Y=0
+ $X2=11.53 $Y2=0
r231 73 99 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=8.02 $Y=0 $X2=7.92
+ $Y2=0
r232 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.02 $Y=0 $X2=8.185
+ $Y2=0
r233 72 102 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=8.35 $Y=0 $X2=8.4
+ $Y2=0
r234 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.35 $Y=0 $X2=8.185
+ $Y2=0
r235 70 96 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.05 $Y=0 $X2=6.96
+ $Y2=0
r236 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.05 $Y=0 $X2=7.215
+ $Y2=0
r237 69 99 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=7.38 $Y=0 $X2=7.92
+ $Y2=0
r238 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.38 $Y=0 $X2=7.215
+ $Y2=0
r239 67 90 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.6
+ $Y2=0
r240 67 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.74
+ $Y2=0
r241 66 93 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.865 $Y=0
+ $X2=4.08 $Y2=0
r242 66 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.865 $Y=0 $X2=3.74
+ $Y2=0
r243 62 139 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.94 $Y=0.085
+ $X2=19.94 $Y2=0
r244 62 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=19.94 $Y=0.085
+ $X2=19.94 $Y2=0.43
r245 61 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=19.055 $Y=0
+ $X2=18.93 $Y2=0
r246 60 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.855 $Y=0
+ $X2=19.94 $Y2=0
r247 60 61 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=19.855 $Y=0
+ $X2=19.055 $Y2=0
r248 56 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=18.93 $Y=0.085
+ $X2=18.93 $Y2=0
r249 56 58 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=18.93 $Y=0.085
+ $X2=18.93 $Y2=0.575
r250 52 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.64 $Y=0.085
+ $X2=17.64 $Y2=0
r251 52 54 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=17.64 $Y=0.085
+ $X2=17.64 $Y2=0.43
r252 48 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.29 $Y=0.085
+ $X2=13.29 $Y2=0
r253 48 50 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=13.29 $Y=0.085
+ $X2=13.29 $Y2=0.725
r254 44 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.53 $Y=0.085
+ $X2=11.53 $Y2=0
r255 44 46 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=11.53 $Y=0.085
+ $X2=11.53 $Y2=0.795
r256 40 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.185 $Y=0.085
+ $X2=8.185 $Y2=0
r257 40 42 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=8.185 $Y=0.085
+ $X2=8.185 $Y2=0.74
r258 36 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=0.085
+ $X2=7.215 $Y2=0
r259 36 38 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=7.215 $Y=0.085
+ $X2=7.215 $Y2=0.745
r260 32 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=0.085
+ $X2=3.74 $Y2=0
r261 32 34 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=3.74 $Y=0.085
+ $X2=3.74 $Y2=0.81
r262 28 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0
r263 28 30 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.76
r264 9 64 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=19.805
+ $Y=0.285 $X2=19.94 $Y2=0.43
r265 8 58 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=18.83
+ $Y=0.365 $X2=18.97 $Y2=0.575
r266 7 54 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=17.395
+ $Y=0.485 $X2=17.64 $Y2=0.43
r267 6 50 182 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_NDIFF $count=1 $X=13.15
+ $Y=0.595 $X2=13.29 $Y2=0.725
r268 5 46 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=11.39
+ $Y=0.625 $X2=11.53 $Y2=0.795
r269 4 42 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.045
+ $Y=0.595 $X2=8.185 $Y2=0.74
r270 3 38 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=7.075
+ $Y=0.595 $X2=7.215 $Y2=0.745
r271 2 34 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.645
+ $Y=0.6 $X2=3.78 $Y2=0.81
r272 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.55 $X2=0.7 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%noxref_29 1 2 9 11 12 15
c26 12 0 2.11477e-20 $X=1.32 $Y=0.34
r27 13 15 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=3.28 $Y=0.425
+ $X2=3.28 $Y2=0.85
r28 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.155 $Y=0.34
+ $X2=3.28 $Y2=0.425
r29 11 12 119.717 $w=1.68e-07 $l=1.835e-06 $layer=LI1_cond $X=3.155 $Y=0.34
+ $X2=1.32 $Y2=0.34
r30 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.195 $Y=0.425
+ $X2=1.32 $Y2=0.34
r31 7 9 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=1.195 $Y=0.425 $X2=1.195
+ $Y2=0.825
r32 2 15 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=3.1
+ $Y=0.68 $X2=3.24 $Y2=0.85
r33 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.68 $X2=1.235 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%noxref_31 1 2 9 11 12 15
c32 12 0 1.29647e-19 $X=2.975 $Y=1.295
r33 13 15 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.21 $Y=1.21 $X2=4.21
+ $Y2=0.81
r34 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.045 $Y=1.295
+ $X2=4.21 $Y2=1.21
r35 11 12 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.045 $Y=1.295
+ $X2=2.975 $Y2=1.295
r36 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.81 $Y=1.21
+ $X2=2.975 $Y2=1.295
r37 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.81 $Y=1.21 $X2=2.81
+ $Y2=0.89
r38 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.07
+ $Y=0.6 $X2=4.21 $Y2=0.81
r39 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.67
+ $Y=0.68 $X2=2.81 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_929_152# 1 2 9 11 12 15
r35 13 15 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6.425 $Y=0.425
+ $X2=6.425 $Y2=0.745
r36 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.26 $Y=0.34
+ $X2=6.425 $Y2=0.425
r37 11 12 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=6.26 $Y=0.34
+ $X2=4.865 $Y2=0.34
r38 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.74 $Y=0.425
+ $X2=4.865 $Y2=0.34
r39 7 9 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=4.74 $Y=0.425
+ $X2=4.74 $Y2=0.91
r40 2 15 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=6.29
+ $Y=0.595 $X2=6.425 $Y2=0.745
r41 1 9 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=4.645
+ $Y=0.76 $X2=4.78 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTP_1%A_2544_119# 1 2 9 11 12 15
r32 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=13.76 $Y=0.98
+ $X2=13.76 $Y2=0.805
r33 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.675 $Y=1.065
+ $X2=13.76 $Y2=0.98
r34 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=13.675 $Y=1.065
+ $X2=12.945 $Y2=1.065
r35 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.82 $Y=0.98
+ $X2=12.945 $Y2=1.065
r36 7 9 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=12.82 $Y=0.98
+ $X2=12.82 $Y2=0.805
r37 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.62
+ $Y=0.595 $X2=13.76 $Y2=0.805
r38 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.72
+ $Y=0.595 $X2=12.86 $Y2=0.805
.ends

