* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_85_367# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 Y C1 a_85_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_1334_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_546_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_85_367# B1 a_533_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_85_367# B1 a_533_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR A2 a_533_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 Y B1 a_546_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND A2 a_1334_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VGND B2 a_546_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 Y C1 a_85_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 Y A1 a_1334_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_1334_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_533_367# B1 a_85_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VPWR A2 a_533_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VGND A2 a_1334_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_533_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 a_533_367# B1 a_85_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND B2 a_546_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_546_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 Y B1 a_546_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_85_367# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_1334_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_533_367# B2 a_85_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 a_533_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VPWR A1 a_533_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_1334_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 a_546_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 a_85_367# B2 a_533_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 a_533_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 a_533_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 a_546_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 a_533_367# B2 a_85_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 VPWR A1 a_533_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 a_85_367# B2 a_533_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 Y A1 a_1334_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
