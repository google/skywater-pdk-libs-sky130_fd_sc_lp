* File: sky130_fd_sc_lp__bufbuf_16.pex.spice
* Created: Wed Sep  2 09:35:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFBUF_16%A 3 7 9 12 13
r31 12 15 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.352 $Y=1.46
+ $X2=0.352 $Y2=1.625
r32 12 14 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.352 $Y=1.46
+ $X2=0.352 $Y2=1.295
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.46 $X2=0.32 $Y2=1.46
r34 9 13 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.32 $Y=1.665
+ $X2=0.32 $Y2=1.46
r35 7 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.625
r36 3 14 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.475 $Y=0.665
+ $X2=0.475 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_16%A_27_49# 1 2 9 13 17 21 25 29 33 35 37 39
+ 40 41 44 46 52 53 57 58
c103 53 0 9.40868e-20 $X=2.015 $Y=1.49
c104 52 0 1.2152e-19 $X=2.015 $Y=1.49
r105 64 65 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.335 $Y=1.49
+ $X2=1.765 $Y2=1.49
r106 58 65 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.49
+ $X2=1.765 $Y2=1.49
r107 53 58 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.015 $Y=1.49
+ $X2=1.84 $Y2=1.49
r108 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.015
+ $Y=1.49 $X2=2.015 $Y2=1.49
r109 50 64 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.995 $Y=1.49
+ $X2=1.335 $Y2=1.49
r110 50 61 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.995 $Y=1.49
+ $X2=0.905 $Y2=1.49
r111 49 52 61.1499 $w=1.83e-07 $l=1.02e-06 $layer=LI1_cond $X=0.995 $Y=1.497
+ $X2=2.015 $Y2=1.497
r112 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.995
+ $Y=1.49 $X2=0.995 $Y2=1.49
r113 47 57 1.03991 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=1.497
+ $X2=0.75 $Y2=1.497
r114 47 49 9.59214 $w=1.83e-07 $l=1.6e-07 $layer=LI1_cond $X=0.835 $Y=1.497
+ $X2=0.995 $Y2=1.497
r115 45 57 5.53942 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=0.75 $Y=1.59
+ $X2=0.75 $Y2=1.497
r116 45 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.75 $Y=1.59
+ $X2=0.75 $Y2=1.92
r117 44 57 5.53942 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=0.75 $Y=1.405
+ $X2=0.75 $Y2=1.497
r118 43 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.75 $Y=1.185
+ $X2=0.75 $Y2=1.405
r119 42 56 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.39 $Y=2.005
+ $X2=0.242 $Y2=2.005
r120 41 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=2.005
+ $X2=0.75 $Y2=1.92
r121 41 42 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.665 $Y=2.005
+ $X2=0.39 $Y2=2.005
r122 39 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=1.1
+ $X2=0.75 $Y2=1.185
r123 39 40 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.665 $Y=1.1
+ $X2=0.355 $Y2=1.1
r124 35 56 2.72785 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.242 $Y=2.09
+ $X2=0.242 $Y2=2.005
r125 35 37 30.276 $w=2.93e-07 $l=7.75e-07 $layer=LI1_cond $X=0.242 $Y=2.09
+ $X2=0.242 $Y2=2.865
r126 31 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=1.015
+ $X2=0.355 $Y2=1.1
r127 31 33 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=0.225 $Y=1.015
+ $X2=0.225 $Y2=0.42
r128 27 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.655
+ $X2=1.765 $Y2=1.49
r129 27 29 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.765 $Y=1.655
+ $X2=1.765 $Y2=2.465
r130 23 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.325
+ $X2=1.765 $Y2=1.49
r131 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.765 $Y=1.325
+ $X2=1.765 $Y2=0.665
r132 19 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.655
+ $X2=1.335 $Y2=1.49
r133 19 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.335 $Y=1.655
+ $X2=1.335 $Y2=2.465
r134 15 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.325
+ $X2=1.335 $Y2=1.49
r135 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.325
+ $X2=1.335 $Y2=0.665
r136 11 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.655
+ $X2=0.905 $Y2=1.49
r137 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.905 $Y=1.655
+ $X2=0.905 $Y2=2.465
r138 7 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.49
r139 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=0.665
r140 2 56 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.085
r141 2 37 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.865
r142 1 33 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.245 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_16%A_196_49# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 69 71 72 73 74 77 81 85 87 90 96 99 100 113
c169 113 0 1.2152e-19 $X=5.125 $Y=1.48
c170 96 0 1.58852e-19 $X=4.97 $Y=1.48
c171 19 0 9.40868e-20 $X=2.975 $Y=2.465
r172 110 111 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.265 $Y=1.48
+ $X2=4.695 $Y2=1.48
r173 109 110 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.835 $Y=1.48
+ $X2=4.265 $Y2=1.48
r174 108 109 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.405 $Y=1.48
+ $X2=3.835 $Y2=1.48
r175 107 108 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.975 $Y=1.48
+ $X2=3.405 $Y2=1.48
r176 103 104 7.88995 $w=5.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.602 $Y=1.48
+ $X2=2.602 $Y2=1.575
r177 97 113 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=4.97 $Y=1.48
+ $X2=5.125 $Y2=1.48
r178 97 111 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=4.97 $Y=1.48
+ $X2=4.695 $Y2=1.48
r179 96 97 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=4.97
+ $Y=1.48 $X2=4.97 $Y2=1.48
r180 94 107 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=2.93 $Y=1.48
+ $X2=2.975 $Y2=1.48
r181 93 96 119.081 $w=1.88e-07 $l=2.04e-06 $layer=LI1_cond $X=2.93 $Y=1.48
+ $X2=4.97 $Y2=1.48
r182 93 94 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=2.93
+ $Y=1.48 $X2=2.93 $Y2=1.48
r183 91 103 6.52558 $w=1.9e-07 $l=2.53e-07 $layer=LI1_cond $X=2.855 $Y=1.48
+ $X2=2.602 $Y2=1.48
r184 91 93 4.37799 $w=1.88e-07 $l=7.5e-08 $layer=LI1_cond $X=2.855 $Y=1.48
+ $X2=2.93 $Y2=1.48
r185 90 104 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.435 $Y=1.76
+ $X2=2.435 $Y2=1.575
r186 88 100 7.00709 $w=1.77e-07 $l=1.33454e-07 $layer=LI1_cond $X=2.145 $Y=1.845
+ $X2=2.015 $Y2=1.852
r187 87 90 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.35 $Y=1.845
+ $X2=2.435 $Y2=1.76
r188 87 88 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.35 $Y=1.845
+ $X2=2.145 $Y2=1.845
r189 86 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.145 $Y=1.15
+ $X2=2.015 $Y2=1.15
r190 85 103 7.81596 $w=5.03e-07 $l=3.3e-07 $layer=LI1_cond $X=2.602 $Y=1.15
+ $X2=2.602 $Y2=1.48
r191 85 86 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.35 $Y=1.15
+ $X2=2.145 $Y2=1.15
r192 81 83 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=2.015 $Y=2.025
+ $X2=2.015 $Y2=2.865
r193 79 100 0.0115521 $w=2.6e-07 $l=9.3e-08 $layer=LI1_cond $X=2.015 $Y=1.945
+ $X2=2.015 $Y2=1.852
r194 79 81 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=2.015 $Y=1.945
+ $X2=2.015 $Y2=2.025
r195 75 99 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=1.065
+ $X2=2.015 $Y2=1.15
r196 75 77 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=2.015 $Y=1.065
+ $X2=2.015 $Y2=0.42
r197 73 100 7.00709 $w=1.77e-07 $l=1.3e-07 $layer=LI1_cond $X=1.885 $Y=1.852
+ $X2=2.015 $Y2=1.852
r198 73 74 40.1671 $w=1.83e-07 $l=6.7e-07 $layer=LI1_cond $X=1.885 $Y=1.852
+ $X2=1.215 $Y2=1.852
r199 71 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.885 $Y=1.15
+ $X2=2.015 $Y2=1.15
r200 71 72 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.885 $Y=1.15
+ $X2=1.215 $Y2=1.15
r201 67 72 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.12 $Y=1.065
+ $X2=1.215 $Y2=1.15
r202 67 69 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=1.12 $Y=1.065
+ $X2=1.12 $Y2=0.42
r203 63 65 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=1.11 $Y=2.025
+ $X2=1.11 $Y2=2.865
r204 61 74 6.85207 $w=1.85e-07 $l=1.44187e-07 $layer=LI1_cond $X=1.11 $Y=1.945
+ $X2=1.215 $Y2=1.852
r205 61 63 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.11 $Y=1.945
+ $X2=1.11 $Y2=2.025
r206 57 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.125 $Y=1.645
+ $X2=5.125 $Y2=1.48
r207 57 59 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.125 $Y=1.645
+ $X2=5.125 $Y2=2.465
r208 53 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.125 $Y=1.315
+ $X2=5.125 $Y2=1.48
r209 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.125 $Y=1.315
+ $X2=5.125 $Y2=0.655
r210 49 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.695 $Y=1.645
+ $X2=4.695 $Y2=1.48
r211 49 51 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=4.695 $Y=1.645
+ $X2=4.695 $Y2=2.465
r212 45 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.695 $Y=1.315
+ $X2=4.695 $Y2=1.48
r213 45 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.695 $Y=1.315
+ $X2=4.695 $Y2=0.655
r214 41 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.645
+ $X2=4.265 $Y2=1.48
r215 41 43 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=4.265 $Y=1.645
+ $X2=4.265 $Y2=2.465
r216 37 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.315
+ $X2=4.265 $Y2=1.48
r217 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.265 $Y=1.315
+ $X2=4.265 $Y2=0.655
r218 33 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.835 $Y=1.645
+ $X2=3.835 $Y2=1.48
r219 33 35 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.835 $Y=1.645
+ $X2=3.835 $Y2=2.465
r220 29 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.835 $Y=1.315
+ $X2=3.835 $Y2=1.48
r221 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.835 $Y=1.315
+ $X2=3.835 $Y2=0.655
r222 25 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.405 $Y=1.645
+ $X2=3.405 $Y2=1.48
r223 25 27 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.405 $Y=1.645
+ $X2=3.405 $Y2=2.465
r224 21 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.405 $Y=1.315
+ $X2=3.405 $Y2=1.48
r225 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.405 $Y=1.315
+ $X2=3.405 $Y2=0.655
r226 17 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.645
+ $X2=2.975 $Y2=1.48
r227 17 19 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.975 $Y=1.645
+ $X2=2.975 $Y2=2.465
r228 13 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.315
+ $X2=2.975 $Y2=1.48
r229 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.975 $Y=1.315
+ $X2=2.975 $Y2=0.655
r230 4 83 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.865
r231 4 81 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.025
r232 3 65 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.865
r233 3 63 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.025
r234 2 77 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.245 $X2=1.98 $Y2=0.42
r235 1 69 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.245 $X2=1.12 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_16%A_610_47# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 53 57 61 65 69 73 77 81 85 89 93 97 101 105 109 113 117 121 125 129 133 137
+ 141 145 149 153 157 158 159 160 163 167 171 173 177 181 185 187 189 190 191
+ 192 197 218 226 231 236 241 246 251 256 258
c382 258 0 1.58852e-19 $X=12.005 $Y=1.48
c383 187 0 1.55749e-19 $X=5.305 $Y=1.835
r384 257 258 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=11.575 $Y=1.48
+ $X2=12.005 $Y2=1.48
r385 255 257 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=11.36 $Y=1.48
+ $X2=11.575 $Y2=1.48
r386 255 256 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.36
+ $Y=1.48 $X2=11.36 $Y2=1.48
r387 253 255 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=11.145 $Y=1.48
+ $X2=11.36 $Y2=1.48
r388 252 253 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=10.715 $Y=1.48
+ $X2=11.145 $Y2=1.48
r389 250 252 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=10.5 $Y=1.48
+ $X2=10.715 $Y2=1.48
r390 250 251 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.5
+ $Y=1.48 $X2=10.5 $Y2=1.48
r391 248 250 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=10.285 $Y=1.48
+ $X2=10.5 $Y2=1.48
r392 247 248 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=9.855 $Y=1.48
+ $X2=10.285 $Y2=1.48
r393 245 247 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=9.64 $Y=1.48
+ $X2=9.855 $Y2=1.48
r394 245 246 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.64
+ $Y=1.48 $X2=9.64 $Y2=1.48
r395 243 245 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=9.425 $Y=1.48
+ $X2=9.64 $Y2=1.48
r396 242 243 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=8.995 $Y=1.48
+ $X2=9.425 $Y2=1.48
r397 240 242 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=8.78 $Y=1.48
+ $X2=8.995 $Y2=1.48
r398 240 241 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.78
+ $Y=1.48 $X2=8.78 $Y2=1.48
r399 238 240 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=8.565 $Y=1.48
+ $X2=8.78 $Y2=1.48
r400 237 238 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=8.135 $Y=1.48
+ $X2=8.565 $Y2=1.48
r401 235 237 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.92 $Y=1.48
+ $X2=8.135 $Y2=1.48
r402 235 236 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.92
+ $Y=1.48 $X2=7.92 $Y2=1.48
r403 233 235 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.705 $Y=1.48
+ $X2=7.92 $Y2=1.48
r404 232 233 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.275 $Y=1.48
+ $X2=7.705 $Y2=1.48
r405 230 232 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.06 $Y=1.48
+ $X2=7.275 $Y2=1.48
r406 230 231 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.06
+ $Y=1.48 $X2=7.06 $Y2=1.48
r407 228 230 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.845 $Y=1.48
+ $X2=7.06 $Y2=1.48
r408 227 228 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.415 $Y=1.48
+ $X2=6.845 $Y2=1.48
r409 225 227 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.2 $Y=1.48
+ $X2=6.415 $Y2=1.48
r410 225 226 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.2
+ $Y=1.48 $X2=6.2 $Y2=1.48
r411 223 225 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.985 $Y=1.48
+ $X2=6.2 $Y2=1.48
r412 221 223 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.555 $Y=1.48
+ $X2=5.985 $Y2=1.48
r413 219 256 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=11.36 $Y=1.665
+ $X2=11.36 $Y2=1.48
r414 218 219 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.36 $Y=1.665
+ $X2=11.36 $Y2=1.665
r415 216 251 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=10.5 $Y=1.665
+ $X2=10.5 $Y2=1.48
r416 215 218 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=10.5 $Y=1.665
+ $X2=11.36 $Y2=1.665
r417 215 216 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.5 $Y=1.665
+ $X2=10.5 $Y2=1.665
r418 213 246 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=9.64 $Y=1.665
+ $X2=9.64 $Y2=1.48
r419 212 215 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=9.64 $Y=1.665
+ $X2=10.5 $Y2=1.665
r420 212 213 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.64 $Y=1.665
+ $X2=9.64 $Y2=1.665
r421 210 241 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=8.78 $Y=1.665
+ $X2=8.78 $Y2=1.48
r422 209 212 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=8.78 $Y=1.665
+ $X2=9.64 $Y2=1.665
r423 209 210 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.78 $Y=1.665
+ $X2=8.78 $Y2=1.665
r424 207 236 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.48
r425 206 209 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.92 $Y=1.665
+ $X2=8.78 $Y2=1.665
r426 206 207 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.665
r427 204 231 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=7.06 $Y=1.665
+ $X2=7.06 $Y2=1.48
r428 203 206 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.06 $Y=1.665
+ $X2=7.92 $Y2=1.665
r429 203 204 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.06 $Y=1.665
+ $X2=7.06 $Y2=1.665
r430 201 226 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=6.2 $Y=1.665
+ $X2=6.2 $Y2=1.48
r431 200 203 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.2 $Y=1.665
+ $X2=7.06 $Y2=1.665
r432 200 201 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.2 $Y=1.665
+ $X2=6.2 $Y2=1.665
r433 196 200 0.513283 $w=2.3e-07 $l=8e-07 $layer=MET1_cond $X=5.4 $Y=1.665
+ $X2=6.2 $Y2=1.665
r434 196 197 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.4 $Y=1.665
+ $X2=5.4 $Y2=1.665
r435 194 197 4.66986 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=5.4 $Y=1.745
+ $X2=5.4 $Y2=1.665
r436 193 197 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=5.4 $Y=1.215
+ $X2=5.4 $Y2=1.665
r437 188 192 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=5.04 $Y=1.835
+ $X2=4.91 $Y2=1.835
r438 187 194 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=5.305 $Y=1.835
+ $X2=5.4 $Y2=1.745
r439 187 188 16.3283 $w=1.78e-07 $l=2.65e-07 $layer=LI1_cond $X=5.305 $Y=1.835
+ $X2=5.04 $Y2=1.835
r440 186 191 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.04 $Y=1.13
+ $X2=4.91 $Y2=1.13
r441 185 193 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.305 $Y=1.13
+ $X2=5.4 $Y2=1.215
r442 185 186 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.305 $Y=1.13
+ $X2=5.04 $Y2=1.13
r443 181 183 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=4.91 $Y=2.045
+ $X2=4.91 $Y2=2.885
r444 179 192 0.0585112 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=4.91 $Y=1.925
+ $X2=4.91 $Y2=1.835
r445 179 181 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=4.91 $Y=1.925
+ $X2=4.91 $Y2=2.045
r446 175 191 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=1.045
+ $X2=4.91 $Y2=1.13
r447 175 177 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=4.91 $Y=1.045
+ $X2=4.91 $Y2=0.45
r448 174 190 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=4.18 $Y=1.835
+ $X2=4.05 $Y2=1.835
r449 173 192 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=4.78 $Y=1.835
+ $X2=4.91 $Y2=1.835
r450 173 174 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=4.78 $Y=1.835
+ $X2=4.18 $Y2=1.835
r451 172 189 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.18 $Y=1.13
+ $X2=4.05 $Y2=1.13
r452 171 191 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.78 $Y=1.13
+ $X2=4.91 $Y2=1.13
r453 171 172 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.78 $Y=1.13
+ $X2=4.18 $Y2=1.13
r454 167 169 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=4.05 $Y=2.045
+ $X2=4.05 $Y2=2.885
r455 165 190 0.0585112 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=4.05 $Y=1.925
+ $X2=4.05 $Y2=1.835
r456 165 167 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=4.05 $Y=1.925
+ $X2=4.05 $Y2=2.045
r457 161 189 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=1.045
+ $X2=4.05 $Y2=1.13
r458 161 163 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=4.05 $Y=1.045
+ $X2=4.05 $Y2=0.45
r459 159 190 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=3.92 $Y=1.835
+ $X2=4.05 $Y2=1.835
r460 159 160 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=3.92 $Y=1.835
+ $X2=3.32 $Y2=1.835
r461 157 189 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.92 $Y=1.13
+ $X2=4.05 $Y2=1.13
r462 157 158 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.92 $Y=1.13
+ $X2=3.285 $Y2=1.13
r463 153 155 43.0245 $w=2.23e-07 $l=8.4e-07 $layer=LI1_cond $X=3.207 $Y=2.045
+ $X2=3.207 $Y2=2.885
r464 151 160 6.92652 $w=1.8e-07 $l=1.51456e-07 $layer=LI1_cond $X=3.207 $Y=1.925
+ $X2=3.32 $Y2=1.835
r465 151 153 6.14636 $w=2.23e-07 $l=1.2e-07 $layer=LI1_cond $X=3.207 $Y=1.925
+ $X2=3.207 $Y2=2.045
r466 147 158 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.17 $Y=1.045
+ $X2=3.285 $Y2=1.13
r467 147 149 29.8132 $w=2.28e-07 $l=5.95e-07 $layer=LI1_cond $X=3.17 $Y=1.045
+ $X2=3.17 $Y2=0.45
r468 143 258 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.005 $Y=1.645
+ $X2=12.005 $Y2=1.48
r469 143 145 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=12.005 $Y=1.645
+ $X2=12.005 $Y2=2.465
r470 139 258 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.005 $Y=1.315
+ $X2=12.005 $Y2=1.48
r471 139 141 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.005 $Y=1.315
+ $X2=12.005 $Y2=0.655
r472 135 257 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.575 $Y=1.645
+ $X2=11.575 $Y2=1.48
r473 135 137 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=11.575 $Y=1.645
+ $X2=11.575 $Y2=2.465
r474 131 257 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.575 $Y=1.315
+ $X2=11.575 $Y2=1.48
r475 131 133 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.575 $Y=1.315
+ $X2=11.575 $Y2=0.655
r476 127 253 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.145 $Y=1.645
+ $X2=11.145 $Y2=1.48
r477 127 129 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=11.145 $Y=1.645
+ $X2=11.145 $Y2=2.465
r478 123 253 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.145 $Y=1.315
+ $X2=11.145 $Y2=1.48
r479 123 125 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.145 $Y=1.315
+ $X2=11.145 $Y2=0.655
r480 119 252 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.715 $Y=1.645
+ $X2=10.715 $Y2=1.48
r481 119 121 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=10.715 $Y=1.645
+ $X2=10.715 $Y2=2.465
r482 115 252 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.715 $Y=1.315
+ $X2=10.715 $Y2=1.48
r483 115 117 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.715 $Y=1.315
+ $X2=10.715 $Y2=0.655
r484 111 248 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.285 $Y=1.645
+ $X2=10.285 $Y2=1.48
r485 111 113 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=10.285 $Y=1.645
+ $X2=10.285 $Y2=2.465
r486 107 248 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.285 $Y=1.315
+ $X2=10.285 $Y2=1.48
r487 107 109 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.285 $Y=1.315
+ $X2=10.285 $Y2=0.655
r488 103 247 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.855 $Y=1.645
+ $X2=9.855 $Y2=1.48
r489 103 105 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=9.855 $Y=1.645
+ $X2=9.855 $Y2=2.465
r490 99 247 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.855 $Y=1.315
+ $X2=9.855 $Y2=1.48
r491 99 101 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.855 $Y=1.315
+ $X2=9.855 $Y2=0.655
r492 95 243 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.425 $Y=1.645
+ $X2=9.425 $Y2=1.48
r493 95 97 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=9.425 $Y=1.645
+ $X2=9.425 $Y2=2.465
r494 91 243 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.425 $Y=1.315
+ $X2=9.425 $Y2=1.48
r495 91 93 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.425 $Y=1.315
+ $X2=9.425 $Y2=0.655
r496 87 242 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.995 $Y=1.645
+ $X2=8.995 $Y2=1.48
r497 87 89 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=8.995 $Y=1.645
+ $X2=8.995 $Y2=2.465
r498 83 242 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.995 $Y=1.315
+ $X2=8.995 $Y2=1.48
r499 83 85 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.995 $Y=1.315
+ $X2=8.995 $Y2=0.655
r500 79 238 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.645
+ $X2=8.565 $Y2=1.48
r501 79 81 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=8.565 $Y=1.645
+ $X2=8.565 $Y2=2.465
r502 75 238 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.315
+ $X2=8.565 $Y2=1.48
r503 75 77 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.565 $Y=1.315
+ $X2=8.565 $Y2=0.655
r504 71 237 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.135 $Y=1.645
+ $X2=8.135 $Y2=1.48
r505 71 73 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=8.135 $Y=1.645
+ $X2=8.135 $Y2=2.465
r506 67 237 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.135 $Y=1.315
+ $X2=8.135 $Y2=1.48
r507 67 69 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.135 $Y=1.315
+ $X2=8.135 $Y2=0.655
r508 63 233 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.705 $Y=1.645
+ $X2=7.705 $Y2=1.48
r509 63 65 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.705 $Y=1.645
+ $X2=7.705 $Y2=2.465
r510 59 233 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.705 $Y=1.315
+ $X2=7.705 $Y2=1.48
r511 59 61 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.705 $Y=1.315
+ $X2=7.705 $Y2=0.655
r512 55 232 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.275 $Y=1.645
+ $X2=7.275 $Y2=1.48
r513 55 57 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.275 $Y=1.645
+ $X2=7.275 $Y2=2.465
r514 51 232 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.275 $Y=1.315
+ $X2=7.275 $Y2=1.48
r515 51 53 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.275 $Y=1.315
+ $X2=7.275 $Y2=0.655
r516 47 228 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.845 $Y=1.645
+ $X2=6.845 $Y2=1.48
r517 47 49 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.845 $Y=1.645
+ $X2=6.845 $Y2=2.465
r518 43 228 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.845 $Y=1.315
+ $X2=6.845 $Y2=1.48
r519 43 45 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.845 $Y=1.315
+ $X2=6.845 $Y2=0.655
r520 39 227 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.415 $Y=1.645
+ $X2=6.415 $Y2=1.48
r521 39 41 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.415 $Y=1.645
+ $X2=6.415 $Y2=2.465
r522 35 227 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.415 $Y=1.315
+ $X2=6.415 $Y2=1.48
r523 35 37 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.415 $Y=1.315
+ $X2=6.415 $Y2=0.655
r524 31 223 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.985 $Y=1.645
+ $X2=5.985 $Y2=1.48
r525 31 33 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.985 $Y=1.645
+ $X2=5.985 $Y2=2.465
r526 27 223 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.985 $Y=1.315
+ $X2=5.985 $Y2=1.48
r527 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.985 $Y=1.315
+ $X2=5.985 $Y2=0.655
r528 23 221 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.555 $Y=1.645
+ $X2=5.555 $Y2=1.48
r529 23 25 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.555 $Y=1.645
+ $X2=5.555 $Y2=2.465
r530 19 221 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.555 $Y=1.315
+ $X2=5.555 $Y2=1.48
r531 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.555 $Y=1.315
+ $X2=5.555 $Y2=0.655
r532 6 183 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=4.77
+ $Y=1.835 $X2=4.91 $Y2=2.885
r533 6 181 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.77
+ $Y=1.835 $X2=4.91 $Y2=2.045
r534 5 169 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.835 $X2=4.05 $Y2=2.885
r535 5 167 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.835 $X2=4.05 $Y2=2.045
r536 4 155 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=3.05
+ $Y=1.835 $X2=3.19 $Y2=2.885
r537 4 153 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.05
+ $Y=1.835 $X2=3.19 $Y2=2.045
r538 3 177 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=4.77
+ $Y=0.235 $X2=4.91 $Y2=0.45
r539 2 163 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=3.91
+ $Y=0.235 $X2=4.05 $Y2=0.45
r540 1 149 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=3.05
+ $Y=0.235 $X2=3.19 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14 45
+ 49 53 57 63 69 75 81 85 89 95 101 107 113 117 121 125 127 132 133 135 136 137
+ 138 140 141 143 144 145 146 147 149 154 159 174 189 195 198 201 204 207 210
+ 213 217
r233 216 217 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r234 213 214 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r235 210 211 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r236 207 208 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r237 204 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r238 201 202 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r239 199 202 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r240 198 199 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r241 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r242 193 217 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r243 193 214 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r244 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r245 190 213 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.49 $Y=3.33
+ $X2=11.36 $Y2=3.33
r246 190 192 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.49 $Y=3.33
+ $X2=11.76 $Y2=3.33
r247 189 216 4.44548 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.09 $Y=3.33
+ $X2=12.285 $Y2=3.33
r248 189 192 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=12.09 $Y=3.33
+ $X2=11.76 $Y2=3.33
r249 188 214 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r250 187 188 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r251 185 188 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r252 184 185 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r253 182 185 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r254 182 211 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r255 181 182 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r256 179 210 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.05 $Y=3.33
+ $X2=7.92 $Y2=3.33
r257 179 181 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.05 $Y=3.33
+ $X2=8.4 $Y2=3.33
r258 178 211 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r259 178 208 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r260 177 178 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r261 175 207 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.19 $Y=3.33
+ $X2=7.06 $Y2=3.33
r262 175 177 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.19 $Y=3.33
+ $X2=7.44 $Y2=3.33
r263 174 210 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.79 $Y=3.33
+ $X2=7.92 $Y2=3.33
r264 174 177 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.79 $Y=3.33
+ $X2=7.44 $Y2=3.33
r265 172 173 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r266 170 173 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r267 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r268 167 170 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r269 167 205 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r270 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r271 164 204 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.75 $Y=3.33
+ $X2=3.62 $Y2=3.33
r272 164 166 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.75 $Y=3.33
+ $X2=4.08 $Y2=3.33
r273 163 205 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r274 163 202 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r275 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r276 160 201 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=2.76 $Y2=3.33
r277 160 162 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=3.12 $Y2=3.33
r278 159 204 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.49 $Y=3.33
+ $X2=3.62 $Y2=3.33
r279 159 162 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.49 $Y=3.33
+ $X2=3.12 $Y2=3.33
r280 158 199 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r281 158 196 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r282 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r283 155 195 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.69 $Y2=3.33
r284 155 157 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=1.2 $Y2=3.33
r285 154 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.55 $Y2=3.33
r286 154 157 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.2 $Y2=3.33
r287 152 196 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r288 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r289 149 195 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.69 $Y2=3.33
r290 149 151 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r291 147 208 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=6.96 $Y2=3.33
r292 147 173 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=6 $Y2=3.33
r293 145 187 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=10.37 $Y=3.33
+ $X2=10.32 $Y2=3.33
r294 145 146 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.37 $Y=3.33
+ $X2=10.5 $Y2=3.33
r295 143 184 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=9.51 $Y=3.33
+ $X2=9.36 $Y2=3.33
r296 143 144 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.51 $Y=3.33
+ $X2=9.64 $Y2=3.33
r297 142 187 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=9.77 $Y=3.33
+ $X2=10.32 $Y2=3.33
r298 142 144 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.77 $Y=3.33
+ $X2=9.64 $Y2=3.33
r299 140 181 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.65 $Y=3.33
+ $X2=8.4 $Y2=3.33
r300 140 141 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.65 $Y=3.33
+ $X2=8.78 $Y2=3.33
r301 139 184 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.91 $Y=3.33
+ $X2=9.36 $Y2=3.33
r302 139 141 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.91 $Y=3.33
+ $X2=8.78 $Y2=3.33
r303 137 172 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.07 $Y=3.33 $X2=6
+ $Y2=3.33
r304 137 138 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.07 $Y=3.33
+ $X2=6.2 $Y2=3.33
r305 135 169 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.04 $Y2=3.33
r306 135 136 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.34 $Y2=3.33
r307 134 172 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.47 $Y=3.33
+ $X2=6 $Y2=3.33
r308 134 136 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.47 $Y=3.33
+ $X2=5.34 $Y2=3.33
r309 132 166 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.35 $Y=3.33
+ $X2=4.08 $Y2=3.33
r310 132 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.35 $Y=3.33
+ $X2=4.48 $Y2=3.33
r311 131 169 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.61 $Y=3.33
+ $X2=5.04 $Y2=3.33
r312 131 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.61 $Y=3.33
+ $X2=4.48 $Y2=3.33
r313 127 130 31.8387 $w=2.93e-07 $l=8.15e-07 $layer=LI1_cond $X=12.237 $Y=2.09
+ $X2=12.237 $Y2=2.905
r314 125 216 3.03205 $w=2.95e-07 $l=1.06325e-07 $layer=LI1_cond $X=12.237
+ $Y=3.245 $X2=12.285 $Y2=3.33
r315 125 130 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=12.237 $Y=3.245
+ $X2=12.237 $Y2=2.905
r316 121 124 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=11.36 $Y=2.09
+ $X2=11.36 $Y2=2.905
r317 119 213 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=11.36 $Y=3.245
+ $X2=11.36 $Y2=3.33
r318 119 124 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=11.36 $Y=3.245
+ $X2=11.36 $Y2=2.905
r319 118 146 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.63 $Y=3.33
+ $X2=10.5 $Y2=3.33
r320 117 213 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.23 $Y=3.33
+ $X2=11.36 $Y2=3.33
r321 117 118 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=11.23 $Y=3.33
+ $X2=10.63 $Y2=3.33
r322 113 116 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=10.5 $Y=2.09
+ $X2=10.5 $Y2=2.905
r323 111 146 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.5 $Y=3.245
+ $X2=10.5 $Y2=3.33
r324 111 116 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=10.5 $Y=3.245
+ $X2=10.5 $Y2=2.905
r325 107 110 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=9.64 $Y=2.09
+ $X2=9.64 $Y2=2.905
r326 105 144 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.64 $Y=3.245
+ $X2=9.64 $Y2=3.33
r327 105 110 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=9.64 $Y=3.245
+ $X2=9.64 $Y2=2.905
r328 101 104 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=8.78 $Y=2.09
+ $X2=8.78 $Y2=2.905
r329 99 141 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.78 $Y=3.245
+ $X2=8.78 $Y2=3.33
r330 99 104 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=8.78 $Y=3.245
+ $X2=8.78 $Y2=2.905
r331 95 98 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=7.92 $Y=2.09
+ $X2=7.92 $Y2=2.905
r332 93 210 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=3.33
r333 93 98 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=2.905
r334 89 92 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=7.06 $Y=2.09
+ $X2=7.06 $Y2=2.905
r335 87 207 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.06 $Y=3.245
+ $X2=7.06 $Y2=3.33
r336 87 92 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=7.06 $Y=3.245
+ $X2=7.06 $Y2=2.905
r337 86 138 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.33 $Y=3.33
+ $X2=6.2 $Y2=3.33
r338 85 207 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.93 $Y=3.33
+ $X2=7.06 $Y2=3.33
r339 85 86 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.93 $Y=3.33 $X2=6.33
+ $Y2=3.33
r340 81 84 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=6.2 $Y=2.09
+ $X2=6.2 $Y2=2.905
r341 79 138 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.2 $Y=3.245
+ $X2=6.2 $Y2=3.33
r342 79 84 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=6.2 $Y=3.245
+ $X2=6.2 $Y2=2.905
r343 75 78 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=5.34 $Y=2.26
+ $X2=5.34 $Y2=2.94
r344 73 136 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=3.245
+ $X2=5.34 $Y2=3.33
r345 73 78 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=5.34 $Y=3.245
+ $X2=5.34 $Y2=2.94
r346 69 72 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=4.48 $Y=2.26
+ $X2=4.48 $Y2=2.94
r347 67 133 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=3.33
r348 67 72 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=2.94
r349 63 66 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=3.62 $Y=2.26
+ $X2=3.62 $Y2=2.94
r350 61 204 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=3.245
+ $X2=3.62 $Y2=3.33
r351 61 66 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=3.62 $Y=3.245
+ $X2=3.62 $Y2=2.94
r352 57 60 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.76 $Y=2.225
+ $X2=2.76 $Y2=2.905
r353 55 201 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=3.245
+ $X2=2.76 $Y2=3.33
r354 55 60 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.76 $Y=3.245
+ $X2=2.76 $Y2=2.905
r355 54 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.55 $Y2=3.33
r356 53 201 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=2.76 $Y2=3.33
r357 53 54 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=1.715 $Y2=3.33
r358 49 52 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.25
+ $X2=1.55 $Y2=2.93
r359 47 198 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.55 $Y2=3.33
r360 47 52 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.55 $Y2=2.93
r361 43 195 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r362 43 45 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.425
r363 14 130 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=12.08
+ $Y=1.835 $X2=12.22 $Y2=2.905
r364 14 127 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=12.08
+ $Y=1.835 $X2=12.22 $Y2=2.09
r365 13 124 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=11.22
+ $Y=1.835 $X2=11.36 $Y2=2.905
r366 13 121 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=11.22
+ $Y=1.835 $X2=11.36 $Y2=2.09
r367 12 116 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=10.36
+ $Y=1.835 $X2=10.5 $Y2=2.905
r368 12 113 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=10.36
+ $Y=1.835 $X2=10.5 $Y2=2.09
r369 11 110 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=9.5
+ $Y=1.835 $X2=9.64 $Y2=2.905
r370 11 107 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=9.5
+ $Y=1.835 $X2=9.64 $Y2=2.09
r371 10 104 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=8.64
+ $Y=1.835 $X2=8.78 $Y2=2.905
r372 10 101 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=8.64
+ $Y=1.835 $X2=8.78 $Y2=2.09
r373 9 98 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=7.78
+ $Y=1.835 $X2=7.92 $Y2=2.905
r374 9 95 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=7.78
+ $Y=1.835 $X2=7.92 $Y2=2.09
r375 8 92 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=6.92
+ $Y=1.835 $X2=7.06 $Y2=2.905
r376 8 89 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=6.92
+ $Y=1.835 $X2=7.06 $Y2=2.09
r377 7 84 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=6.06
+ $Y=1.835 $X2=6.2 $Y2=2.905
r378 7 81 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=6.06
+ $Y=1.835 $X2=6.2 $Y2=2.09
r379 6 78 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.835 $X2=5.34 $Y2=2.94
r380 6 75 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.835 $X2=5.34 $Y2=2.26
r381 5 72 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=4.34
+ $Y=1.835 $X2=4.48 $Y2=2.94
r382 5 69 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=4.34
+ $Y=1.835 $X2=4.48 $Y2=2.26
r383 4 66 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=1.835 $X2=3.62 $Y2=2.94
r384 4 63 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=1.835 $X2=3.62 $Y2=2.26
r385 3 60 400 $w=1.7e-07 $l=1.13077e-06 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.835 $X2=2.76 $Y2=2.905
r386 3 57 400 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.835 $X2=2.76 $Y2=2.225
r387 2 52 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.93
r388 2 49 400 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.25
r389 1 45 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 49 52 62 72 82 92 102 112 122 126
c185 126 0 1.55749e-19 $X=11.79 $Y=2.035
r186 125 129 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=11.79 $Y=2.035
+ $X2=11.79 $Y2=2.885
r187 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.79 $Y=2.035
+ $X2=11.79 $Y2=2.035
r188 122 125 70.2547 $w=2.58e-07 $l=1.585e-06 $layer=LI1_cond $X=11.79 $Y=0.45
+ $X2=11.79 $Y2=2.035
r189 116 126 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=10.93 $Y=2.035
+ $X2=11.79 $Y2=2.035
r190 115 119 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=10.93 $Y=2.035
+ $X2=10.93 $Y2=2.885
r191 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.93 $Y=2.035
+ $X2=10.93 $Y2=2.035
r192 112 115 70.2547 $w=2.58e-07 $l=1.585e-06 $layer=LI1_cond $X=10.93 $Y=0.45
+ $X2=10.93 $Y2=2.035
r193 106 116 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=10.07 $Y=2.035
+ $X2=10.93 $Y2=2.035
r194 105 109 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=10.07 $Y=2.035
+ $X2=10.07 $Y2=2.885
r195 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.07 $Y=2.035
+ $X2=10.07 $Y2=2.035
r196 102 105 70.2547 $w=2.58e-07 $l=1.585e-06 $layer=LI1_cond $X=10.07 $Y=0.45
+ $X2=10.07 $Y2=2.035
r197 96 106 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=9.21 $Y=2.035
+ $X2=10.07 $Y2=2.035
r198 95 99 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=9.21 $Y=2.035
+ $X2=9.21 $Y2=2.885
r199 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.21 $Y=2.035
+ $X2=9.21 $Y2=2.035
r200 92 95 70.2547 $w=2.58e-07 $l=1.585e-06 $layer=LI1_cond $X=9.21 $Y=0.45
+ $X2=9.21 $Y2=2.035
r201 85 89 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=8.35 $Y=2.035
+ $X2=8.35 $Y2=2.885
r202 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.35 $Y=2.035
+ $X2=8.35 $Y2=2.035
r203 82 85 70.2547 $w=2.58e-07 $l=1.585e-06 $layer=LI1_cond $X=8.35 $Y=0.45
+ $X2=8.35 $Y2=2.035
r204 76 86 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.49 $Y=2.035
+ $X2=8.35 $Y2=2.035
r205 75 79 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=7.49 $Y=2.035
+ $X2=7.49 $Y2=2.885
r206 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.49 $Y=2.035
+ $X2=7.49 $Y2=2.035
r207 72 75 70.2547 $w=2.58e-07 $l=1.585e-06 $layer=LI1_cond $X=7.49 $Y=0.45
+ $X2=7.49 $Y2=2.035
r208 66 76 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.63 $Y=2.035
+ $X2=7.49 $Y2=2.035
r209 65 69 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=6.63 $Y=2.035
+ $X2=6.63 $Y2=2.885
r210 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.63 $Y=2.035
+ $X2=6.63 $Y2=2.035
r211 62 65 70.2547 $w=2.58e-07 $l=1.585e-06 $layer=LI1_cond $X=6.63 $Y=0.45
+ $X2=6.63 $Y2=2.035
r212 56 66 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=5.77 $Y=2.035
+ $X2=6.63 $Y2=2.035
r213 55 59 41.6841 $w=2.33e-07 $l=8.5e-07 $layer=LI1_cond $X=5.782 $Y=2.035
+ $X2=5.782 $Y2=2.885
r214 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.77 $Y=2.035
+ $X2=5.77 $Y2=2.035
r215 52 55 77.7286 $w=2.33e-07 $l=1.585e-06 $layer=LI1_cond $X=5.782 $Y=0.45
+ $X2=5.782 $Y2=2.035
r216 49 96 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=8.78 $Y=2.035
+ $X2=9.21 $Y2=2.035
r217 49 86 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=8.78 $Y=2.035
+ $X2=8.35 $Y2=2.035
r218 16 129 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=11.65
+ $Y=1.835 $X2=11.79 $Y2=2.885
r219 16 125 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.65
+ $Y=1.835 $X2=11.79 $Y2=2.045
r220 15 119 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=10.79
+ $Y=1.835 $X2=10.93 $Y2=2.885
r221 15 115 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=10.79
+ $Y=1.835 $X2=10.93 $Y2=2.045
r222 14 109 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=1.835 $X2=10.07 $Y2=2.885
r223 14 105 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=1.835 $X2=10.07 $Y2=2.045
r224 13 99 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=9.07
+ $Y=1.835 $X2=9.21 $Y2=2.885
r225 13 95 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=9.07
+ $Y=1.835 $X2=9.21 $Y2=2.045
r226 12 89 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.835 $X2=8.35 $Y2=2.885
r227 12 85 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.835 $X2=8.35 $Y2=2.045
r228 11 79 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=7.35
+ $Y=1.835 $X2=7.49 $Y2=2.885
r229 11 75 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.35
+ $Y=1.835 $X2=7.49 $Y2=2.045
r230 10 69 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=6.49
+ $Y=1.835 $X2=6.63 $Y2=2.885
r231 10 65 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.49
+ $Y=1.835 $X2=6.63 $Y2=2.045
r232 9 59 400 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=5.63
+ $Y=1.835 $X2=5.77 $Y2=2.885
r233 9 55 400 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.63
+ $Y=1.835 $X2=5.77 $Y2=2.045
r234 8 122 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=11.65
+ $Y=0.235 $X2=11.79 $Y2=0.45
r235 7 112 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=10.79
+ $Y=0.235 $X2=10.93 $Y2=0.45
r236 6 102 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=9.93
+ $Y=0.235 $X2=10.07 $Y2=0.45
r237 5 92 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=9.07
+ $Y=0.235 $X2=9.21 $Y2=0.45
r238 4 82 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=8.21
+ $Y=0.235 $X2=8.35 $Y2=0.45
r239 3 72 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=7.35
+ $Y=0.235 $X2=7.49 $Y2=0.45
r240 2 62 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=6.49
+ $Y=0.235 $X2=6.63 $Y2=0.45
r241 1 52 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=5.63
+ $Y=0.235 $X2=5.77 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14 45
+ 49 51 55 59 63 67 71 73 77 81 85 89 93 95 99 101 103 106 107 109 110 111 112
+ 114 115 117 118 119 120 121 123 128 133 148 163 169 172 175 178 181 184 187
+ 191
r202 190 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r203 187 188 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r204 184 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r205 181 182 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r206 178 179 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r207 175 176 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r208 173 176 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.64 $Y2=0
r209 172 173 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r210 169 170 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r211 167 191 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r212 167 188 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r213 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r214 164 187 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.49 $Y=0
+ $X2=11.36 $Y2=0
r215 164 166 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.49 $Y=0
+ $X2=11.76 $Y2=0
r216 163 190 4.44548 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.09 $Y=0
+ $X2=12.285 $Y2=0
r217 163 166 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=12.09 $Y=0
+ $X2=11.76 $Y2=0
r218 162 188 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r219 161 162 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r220 159 162 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.32 $Y2=0
r221 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r222 156 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=9.36 $Y2=0
r223 156 185 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=7.92 $Y2=0
r224 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r225 153 184 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.05 $Y=0 $X2=7.92
+ $Y2=0
r226 153 155 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.05 $Y=0 $X2=8.4
+ $Y2=0
r227 152 185 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r228 152 182 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r229 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r230 149 181 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.19 $Y=0 $X2=7.06
+ $Y2=0
r231 149 151 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.19 $Y=0
+ $X2=7.44 $Y2=0
r232 148 184 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.79 $Y=0 $X2=7.92
+ $Y2=0
r233 148 151 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.79 $Y=0
+ $X2=7.44 $Y2=0
r234 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r235 144 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r236 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r237 141 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r238 141 179 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=3.6 $Y2=0
r239 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r240 138 178 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.75 $Y=0
+ $X2=3.602 $Y2=0
r241 138 140 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.75 $Y=0
+ $X2=4.08 $Y2=0
r242 137 179 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=3.6 $Y2=0
r243 137 176 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=2.64 $Y2=0
r244 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r245 134 175 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.885 $Y=0
+ $X2=2.74 $Y2=0
r246 134 136 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.885 $Y=0
+ $X2=3.12 $Y2=0
r247 133 178 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=3.455 $Y=0
+ $X2=3.602 $Y2=0
r248 133 136 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.455 $Y=0
+ $X2=3.12 $Y2=0
r249 132 173 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=1.68 $Y2=0
r250 132 170 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=0.72 $Y2=0
r251 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r252 129 169 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0
+ $X2=0.69 $Y2=0
r253 129 131 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0
+ $X2=1.2 $Y2=0
r254 128 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=1.55 $Y2=0
r255 128 131 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=1.2 $Y2=0
r256 126 170 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r257 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r258 123 169 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.69 $Y2=0
r259 123 125 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.24 $Y2=0
r260 121 182 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.24 $Y=0
+ $X2=6.96 $Y2=0
r261 121 147 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=0 $X2=6
+ $Y2=0
r262 119 161 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=10.37 $Y=0
+ $X2=10.32 $Y2=0
r263 119 120 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.37 $Y=0
+ $X2=10.5 $Y2=0
r264 117 158 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=9.51 $Y=0 $X2=9.36
+ $Y2=0
r265 117 118 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.51 $Y=0 $X2=9.64
+ $Y2=0
r266 116 161 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=9.77 $Y=0
+ $X2=10.32 $Y2=0
r267 116 118 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.77 $Y=0 $X2=9.64
+ $Y2=0
r268 114 155 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.65 $Y=0 $X2=8.4
+ $Y2=0
r269 114 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.65 $Y=0 $X2=8.78
+ $Y2=0
r270 113 158 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.91 $Y=0
+ $X2=9.36 $Y2=0
r271 113 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.91 $Y=0 $X2=8.78
+ $Y2=0
r272 111 146 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.07 $Y=0 $X2=6
+ $Y2=0
r273 111 112 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.07 $Y=0 $X2=6.2
+ $Y2=0
r274 109 143 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.21 $Y=0
+ $X2=5.04 $Y2=0
r275 109 110 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.34
+ $Y2=0
r276 108 146 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.47 $Y=0 $X2=6
+ $Y2=0
r277 108 110 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.47 $Y=0 $X2=5.34
+ $Y2=0
r278 106 140 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.35 $Y=0 $X2=4.08
+ $Y2=0
r279 106 107 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.35 $Y=0 $X2=4.48
+ $Y2=0
r280 105 143 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.61 $Y=0
+ $X2=5.04 $Y2=0
r281 105 107 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.61 $Y=0 $X2=4.48
+ $Y2=0
r282 101 190 3.03205 $w=2.95e-07 $l=1.06325e-07 $layer=LI1_cond $X=12.237
+ $Y=0.085 $X2=12.285 $Y2=0
r283 101 103 14.259 $w=2.93e-07 $l=3.65e-07 $layer=LI1_cond $X=12.237 $Y=0.085
+ $X2=12.237 $Y2=0.45
r284 97 187 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=11.36 $Y=0.085
+ $X2=11.36 $Y2=0
r285 97 99 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=11.36 $Y=0.085
+ $X2=11.36 $Y2=0.45
r286 96 120 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.63 $Y=0 $X2=10.5
+ $Y2=0
r287 95 187 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.23 $Y=0
+ $X2=11.36 $Y2=0
r288 95 96 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=11.23 $Y=0 $X2=10.63
+ $Y2=0
r289 91 120 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0
r290 91 93 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0.45
r291 87 118 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.64 $Y=0.085
+ $X2=9.64 $Y2=0
r292 87 89 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=9.64 $Y=0.085
+ $X2=9.64 $Y2=0.45
r293 83 115 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.78 $Y=0.085
+ $X2=8.78 $Y2=0
r294 83 85 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=8.78 $Y=0.085
+ $X2=8.78 $Y2=0.45
r295 79 184 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=0.085
+ $X2=7.92 $Y2=0
r296 79 81 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=7.92 $Y=0.085
+ $X2=7.92 $Y2=0.45
r297 75 181 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.06 $Y=0.085
+ $X2=7.06 $Y2=0
r298 75 77 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=7.06 $Y=0.085
+ $X2=7.06 $Y2=0.45
r299 74 112 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.33 $Y=0 $X2=6.2
+ $Y2=0
r300 73 181 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.93 $Y=0 $X2=7.06
+ $Y2=0
r301 73 74 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.93 $Y=0 $X2=6.33
+ $Y2=0
r302 69 112 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.2 $Y=0.085
+ $X2=6.2 $Y2=0
r303 69 71 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=6.2 $Y=0.085
+ $X2=6.2 $Y2=0.45
r304 65 110 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.34 $Y2=0
r305 65 67 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.34 $Y2=0.37
r306 61 107 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.48 $Y2=0
r307 61 63 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.48 $Y2=0.37
r308 57 178 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.602 $Y=0.085
+ $X2=3.602 $Y2=0
r309 57 59 11.1338 $w=2.93e-07 $l=2.85e-07 $layer=LI1_cond $X=3.602 $Y=0.085
+ $X2=3.602 $Y2=0.37
r310 53 175 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0
r311 53 55 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0.39
r312 52 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=0
+ $X2=1.55 $Y2=0
r313 51 175 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.595 $Y=0
+ $X2=2.74 $Y2=0
r314 51 52 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.595 $Y=0
+ $X2=1.715 $Y2=0
r315 47 172 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0
r316 47 49 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0.425
r317 43 169 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r318 43 45 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.39
r319 14 103 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=12.08
+ $Y=0.235 $X2=12.22 $Y2=0.45
r320 13 99 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=11.22
+ $Y=0.235 $X2=11.36 $Y2=0.45
r321 12 93 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=10.36
+ $Y=0.235 $X2=10.5 $Y2=0.45
r322 11 89 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=9.5
+ $Y=0.235 $X2=9.64 $Y2=0.45
r323 10 85 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=8.64
+ $Y=0.235 $X2=8.78 $Y2=0.45
r324 9 81 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=7.78
+ $Y=0.235 $X2=7.92 $Y2=0.45
r325 8 77 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=6.92
+ $Y=0.235 $X2=7.06 $Y2=0.45
r326 7 71 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=6.06
+ $Y=0.235 $X2=6.2 $Y2=0.45
r327 6 67 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=5.2
+ $Y=0.235 $X2=5.34 $Y2=0.37
r328 5 63 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=4.34
+ $Y=0.235 $X2=4.48 $Y2=0.37
r329 4 59 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.48
+ $Y=0.235 $X2=3.62 $Y2=0.37
r330 3 55 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=2.635
+ $Y=0.235 $X2=2.76 $Y2=0.39
r331 2 49 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=1.41 $Y=0.245
+ $X2=1.55 $Y2=0.425
r332 1 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.245 $X2=0.69 $Y2=0.39
.ends

