* File: sky130_fd_sc_lp__and2_0.pxi.spice
* Created: Wed Sep  2 09:30:08 2020
* 
x_PM_SKY130_FD_SC_LP__AND2_0%A N_A_c_47_n N_A_M1003_g N_A_M1000_g N_A_c_53_n A A
+ A N_A_c_50_n PM_SKY130_FD_SC_LP__AND2_0%A
x_PM_SKY130_FD_SC_LP__AND2_0%B N_B_M1001_g N_B_c_84_n N_B_M1005_g N_B_c_86_n B B
+ N_B_c_83_n PM_SKY130_FD_SC_LP__AND2_0%B
x_PM_SKY130_FD_SC_LP__AND2_0%A_63_47# N_A_63_47#_M1003_s N_A_63_47#_M1000_d
+ N_A_63_47#_c_120_n N_A_63_47#_M1004_g N_A_63_47#_c_121_n N_A_63_47#_M1002_g
+ N_A_63_47#_c_123_n N_A_63_47#_c_124_n N_A_63_47#_c_125_n N_A_63_47#_c_166_p
+ N_A_63_47#_c_126_n N_A_63_47#_c_134_n N_A_63_47#_c_127_n
+ PM_SKY130_FD_SC_LP__AND2_0%A_63_47#
x_PM_SKY130_FD_SC_LP__AND2_0%VPWR N_VPWR_M1000_s N_VPWR_M1005_d N_VPWR_c_184_n
+ N_VPWR_c_185_n N_VPWR_c_186_n N_VPWR_c_187_n N_VPWR_c_188_n VPWR
+ N_VPWR_c_189_n N_VPWR_c_183_n N_VPWR_c_191_n PM_SKY130_FD_SC_LP__AND2_0%VPWR
x_PM_SKY130_FD_SC_LP__AND2_0%X N_X_M1004_d N_X_M1002_d X X X X X X X X
+ N_X_c_213_n N_X_c_214_n X PM_SKY130_FD_SC_LP__AND2_0%X
x_PM_SKY130_FD_SC_LP__AND2_0%VGND N_VGND_M1001_d N_VGND_c_238_n VGND
+ N_VGND_c_239_n N_VGND_c_240_n N_VGND_c_241_n N_VGND_c_242_n
+ PM_SKY130_FD_SC_LP__AND2_0%VGND
cc_1 VNB N_A_c_47_n 0.0192731f $X=-0.19 $Y=-0.245 $X2=0.512 $Y2=1.663
cc_2 VNB N_A_M1003_g 0.0473927f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.445
cc_3 VNB A 0.0298913f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_50_n 0.0264522f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.375
cc_5 VNB N_B_M1001_g 0.0557488f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.21
cc_6 VNB B 0.00587928f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_B_c_83_n 0.0158916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_63_47#_c_120_n 0.0202947f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.88
cc_9 VNB N_A_63_47#_c_121_n 0.103315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_63_47#_M1002_g 0.0143622f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A_63_47#_c_123_n 0.0224476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_63_47#_c_124_n 0.00841248f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.375
cc_13 VNB N_A_63_47#_c_125_n 0.0133891f $X=-0.19 $Y=-0.245 $X2=0.512 $Y2=1.21
cc_14 VNB N_A_63_47#_c_126_n 0.00856635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_63_47#_c_127_n 0.00569337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_183_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=2.035
cc_17 VNB X 0.0515609f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.605
cc_18 VNB N_X_c_213_n 0.0117488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_X_c_214_n 0.0216375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_238_n 0.0025812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_239_n 0.0322723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_240_n 0.0284434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_241_n 0.160554f $X=-0.19 $Y=-0.245 $X2=0.512 $Y2=1.375
cc_24 VNB N_VGND_c_242_n 0.00424349f $X=-0.19 $Y=-0.245 $X2=0.512 $Y2=1.21
cc_25 VPB N_A_c_47_n 5.94326e-19 $X=-0.19 $Y=1.655 $X2=0.512 $Y2=1.663
cc_26 VPB N_A_M1000_g 0.0407716f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.605
cc_27 VPB N_A_c_53_n 0.0275066f $X=-0.19 $Y=1.655 $X2=0.512 $Y2=1.88
cc_28 VPB A 0.0380837f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_29 VPB N_B_c_84_n 0.021736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_B_M1005_g 0.0238112f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.605
cc_31 VPB N_B_c_86_n 0.0221807f $X=-0.19 $Y=1.655 $X2=0.512 $Y2=1.88
cc_32 VPB B 0.0085289f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_33 VPB N_B_c_83_n 0.00551053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_A_63_47#_M1002_g 0.062731f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_35 VPB N_A_63_47#_c_127_n 0.00498759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_184_n 0.0350471f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.605
cc_37 VPB N_VPWR_c_185_n 0.01783f $X=-0.19 $Y=1.655 $X2=0.512 $Y2=1.88
cc_38 VPB N_VPWR_c_186_n 0.0269571f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_187_n 0.0108943f $X=-0.19 $Y=1.655 $X2=0.512 $Y2=1.375
cc_40 VPB N_VPWR_c_188_n 0.00516749f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.375
cc_41 VPB N_VPWR_c_189_n 0.0189304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_183_n 0.0644913f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=2.035
cc_43 VPB N_VPWR_c_191_n 0.0118035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB X 0.0401172f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.605
cc_45 VPB X 0.0234139f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_46 VPB X 0.0134315f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 N_A_M1003_g N_B_M1001_g 0.031938f $X=0.655 $Y=0.445 $X2=0 $Y2=0
cc_48 N_A_c_47_n N_B_c_84_n 0.031938f $X=0.512 $Y=1.663 $X2=0 $Y2=0
cc_49 N_A_M1000_g N_B_M1005_g 0.0141941f $X=0.655 $Y=2.605 $X2=0 $Y2=0
cc_50 N_A_c_53_n N_B_c_86_n 0.031938f $X=0.512 $Y=1.88 $X2=0 $Y2=0
cc_51 N_A_c_47_n B 5.07445e-19 $X=0.512 $Y=1.663 $X2=0 $Y2=0
cc_52 N_A_c_50_n N_B_c_83_n 0.031938f $X=0.46 $Y=1.375 $X2=0 $Y2=0
cc_53 N_A_M1003_g N_A_63_47#_c_123_n 0.0136593f $X=0.655 $Y=0.445 $X2=0 $Y2=0
cc_54 N_A_M1003_g N_A_63_47#_c_125_n 0.0163848f $X=0.655 $Y=0.445 $X2=0 $Y2=0
cc_55 A N_A_63_47#_c_125_n 0.020605f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A_c_50_n N_A_63_47#_c_125_n 0.00302286f $X=0.46 $Y=1.375 $X2=0 $Y2=0
cc_57 N_A_M1000_g N_A_63_47#_c_134_n 0.00350009f $X=0.655 $Y=2.605 $X2=0 $Y2=0
cc_58 N_A_c_47_n N_A_63_47#_c_127_n 0.00492123f $X=0.512 $Y=1.663 $X2=0 $Y2=0
cc_59 N_A_M1003_g N_A_63_47#_c_127_n 0.00821367f $X=0.655 $Y=0.445 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_A_63_47#_c_127_n 0.0153569f $X=0.655 $Y=2.605 $X2=0 $Y2=0
cc_61 N_A_c_53_n N_A_63_47#_c_127_n 0.00456371f $X=0.512 $Y=1.88 $X2=0 $Y2=0
cc_62 A N_A_63_47#_c_127_n 0.0783676f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A_c_50_n N_A_63_47#_c_127_n 0.00456371f $X=0.46 $Y=1.375 $X2=0 $Y2=0
cc_64 N_A_M1000_g N_VPWR_c_184_n 0.00405922f $X=0.655 $Y=2.605 $X2=0 $Y2=0
cc_65 N_A_c_53_n N_VPWR_c_184_n 9.18505e-19 $X=0.512 $Y=1.88 $X2=0 $Y2=0
cc_66 A N_VPWR_c_184_n 0.0203872f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A_M1000_g N_VPWR_c_185_n 0.00467362f $X=0.655 $Y=2.605 $X2=0 $Y2=0
cc_68 N_A_M1000_g N_VPWR_c_186_n 5.70571e-19 $X=0.655 $Y=2.605 $X2=0 $Y2=0
cc_69 N_A_M1000_g N_VPWR_c_183_n 0.00500913f $X=0.655 $Y=2.605 $X2=0 $Y2=0
cc_70 N_A_M1003_g N_VGND_c_238_n 0.00224374f $X=0.655 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_M1003_g N_VGND_c_239_n 0.0054978f $X=0.655 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A_M1003_g N_VGND_c_241_n 0.00734508f $X=0.655 $Y=0.445 $X2=0 $Y2=0
cc_73 N_B_M1001_g N_A_63_47#_c_120_n 0.0332827f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_74 N_B_M1001_g N_A_63_47#_c_121_n 0.00637197f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_75 B N_A_63_47#_c_121_n 6.18306e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_76 N_B_M1001_g N_A_63_47#_M1002_g 0.00217846f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_77 N_B_M1005_g N_A_63_47#_M1002_g 0.00675648f $X=1.085 $Y=2.605 $X2=0 $Y2=0
cc_78 B N_A_63_47#_M1002_g 0.00609346f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_79 N_B_c_83_n N_A_63_47#_M1002_g 0.0143527f $X=1.16 $Y=1.7 $X2=0 $Y2=0
cc_80 N_B_M1001_g N_A_63_47#_c_123_n 0.00207889f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_81 N_B_M1001_g N_A_63_47#_c_124_n 0.0156386f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_82 B N_A_63_47#_c_124_n 0.0110391f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_83 N_B_c_83_n N_A_63_47#_c_124_n 0.00125128f $X=1.16 $Y=1.7 $X2=0 $Y2=0
cc_84 N_B_M1001_g N_A_63_47#_c_126_n 0.00138367f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_85 N_B_c_86_n N_A_63_47#_c_134_n 0.00112532f $X=1.132 $Y=2.205 $X2=0 $Y2=0
cc_86 N_B_M1001_g N_A_63_47#_c_127_n 0.0123446f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_87 N_B_M1005_g N_A_63_47#_c_127_n 0.00431054f $X=1.085 $Y=2.605 $X2=0 $Y2=0
cc_88 B N_A_63_47#_c_127_n 0.048251f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_89 N_B_M1005_g N_VPWR_c_185_n 0.00445291f $X=1.085 $Y=2.605 $X2=0 $Y2=0
cc_90 N_B_M1005_g N_VPWR_c_186_n 0.0110698f $X=1.085 $Y=2.605 $X2=0 $Y2=0
cc_91 N_B_c_86_n N_VPWR_c_186_n 0.00128253f $X=1.132 $Y=2.205 $X2=0 $Y2=0
cc_92 B N_VPWR_c_186_n 0.0209962f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_93 N_B_M1005_g N_VPWR_c_183_n 0.00470859f $X=1.085 $Y=2.605 $X2=0 $Y2=0
cc_94 B X 0.0206606f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_95 N_B_M1001_g N_VGND_c_238_n 0.0111072f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_96 N_B_M1001_g N_VGND_c_239_n 0.00486043f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_97 N_B_M1001_g N_VGND_c_241_n 0.00446184f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_63_47#_c_134_n N_VPWR_c_185_n 0.00501806f $X=0.87 $Y=2.605 $X2=0 $Y2=0
cc_99 N_A_63_47#_M1002_g N_VPWR_c_186_n 0.00867858f $X=1.855 $Y=2.715 $X2=0
+ $Y2=0
cc_100 N_A_63_47#_c_127_n N_VPWR_c_186_n 0.0031228f $X=0.847 $Y=2.44 $X2=0 $Y2=0
cc_101 N_A_63_47#_M1002_g N_VPWR_c_189_n 0.00526658f $X=1.855 $Y=2.715 $X2=0
+ $Y2=0
cc_102 N_A_63_47#_M1002_g N_VPWR_c_183_n 0.0114972f $X=1.855 $Y=2.715 $X2=0
+ $Y2=0
cc_103 N_A_63_47#_c_134_n N_VPWR_c_183_n 0.00831973f $X=0.87 $Y=2.605 $X2=0
+ $Y2=0
cc_104 N_A_63_47#_c_120_n X 0.00215699f $X=1.445 $Y=0.765 $X2=0 $Y2=0
cc_105 N_A_63_47#_c_121_n X 0.0207791f $X=1.855 $Y=1.435 $X2=0 $Y2=0
cc_106 N_A_63_47#_M1002_g X 0.0277048f $X=1.855 $Y=2.715 $X2=0 $Y2=0
cc_107 N_A_63_47#_c_166_p X 0.0139714f $X=1.73 $Y=1.015 $X2=0 $Y2=0
cc_108 N_A_63_47#_c_126_n X 0.0324771f $X=1.73 $Y=1.27 $X2=0 $Y2=0
cc_109 N_A_63_47#_c_120_n N_X_c_213_n 0.00168379f $X=1.445 $Y=0.765 $X2=0 $Y2=0
cc_110 N_A_63_47#_c_121_n N_X_c_213_n 0.0162988f $X=1.855 $Y=1.435 $X2=0 $Y2=0
cc_111 N_A_63_47#_c_124_n N_X_c_213_n 0.00334238f $X=1.565 $Y=0.93 $X2=0 $Y2=0
cc_112 N_A_63_47#_c_166_p N_X_c_213_n 0.0271191f $X=1.73 $Y=1.015 $X2=0 $Y2=0
cc_113 N_A_63_47#_M1002_g X 7.11522e-19 $X=1.855 $Y=2.715 $X2=0 $Y2=0
cc_114 N_A_63_47#_c_120_n N_VGND_c_238_n 0.0031293f $X=1.445 $Y=0.765 $X2=0
+ $Y2=0
cc_115 N_A_63_47#_c_123_n N_VGND_c_238_n 0.0108521f $X=0.44 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_63_47#_c_124_n N_VGND_c_238_n 0.0141266f $X=1.565 $Y=0.93 $X2=0 $Y2=0
cc_117 N_A_63_47#_c_123_n N_VGND_c_239_n 0.0164055f $X=0.44 $Y=0.445 $X2=0 $Y2=0
cc_118 N_A_63_47#_c_120_n N_VGND_c_240_n 0.00585385f $X=1.445 $Y=0.765 $X2=0
+ $Y2=0
cc_119 N_A_63_47#_M1003_s N_VGND_c_241_n 0.00216892f $X=0.315 $Y=0.235 $X2=0
+ $Y2=0
cc_120 N_A_63_47#_c_120_n N_VGND_c_241_n 0.00775698f $X=1.445 $Y=0.765 $X2=0
+ $Y2=0
cc_121 N_A_63_47#_c_123_n N_VGND_c_241_n 0.0114541f $X=0.44 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_63_47#_c_124_n N_VGND_c_241_n 0.00585106f $X=1.565 $Y=0.93 $X2=0
+ $Y2=0
cc_123 N_A_63_47#_c_125_n N_VGND_c_241_n 0.0141135f $X=0.895 $Y=0.93 $X2=0 $Y2=0
cc_124 N_VPWR_c_189_n X 0.0240432f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_125 N_VPWR_c_183_n X 0.014552f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_126 N_VPWR_c_186_n X 0.00246979f $X=1.3 $Y=2.55 $X2=0 $Y2=0
cc_127 N_X_c_213_n N_VGND_c_240_n 0.0303259f $X=2.065 $Y=0.477 $X2=0 $Y2=0
cc_128 N_X_c_214_n N_VGND_c_240_n 0.0154715f $X=2.19 $Y=0.675 $X2=0 $Y2=0
cc_129 N_X_M1004_d N_VGND_c_241_n 0.0021695f $X=1.52 $Y=0.235 $X2=0 $Y2=0
cc_130 N_X_c_213_n N_VGND_c_241_n 0.0205961f $X=2.065 $Y=0.477 $X2=0 $Y2=0
cc_131 N_X_c_214_n N_VGND_c_241_n 0.00960138f $X=2.19 $Y=0.675 $X2=0 $Y2=0
cc_132 A_146_47# N_VGND_c_241_n 0.00309736f $X=0.73 $Y=0.235 $X2=2.16 $Y2=0
