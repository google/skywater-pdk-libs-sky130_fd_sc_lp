* File: sky130_fd_sc_lp__bushold0_1.pxi.spice
* Created: Wed Sep  2 09:37:40 2020
* 
x_PM_SKY130_FD_SC_LP__BUSHOLD0_1%X N_X_M1000_d N_X_M1001_d N_X_M1005_g
+ N_X_M1003_g N_X_c_60_n N_X_c_61_n N_X_c_52_n N_X_c_53_n N_X_c_64_n N_X_c_65_n
+ N_X_c_54_n N_X_c_55_n N_X_c_56_n X X X X X X N_X_c_58_n
+ PM_SKY130_FD_SC_LP__BUSHOLD0_1%X
x_PM_SKY130_FD_SC_LP__BUSHOLD0_1%RESET N_RESET_M1000_g N_RESET_M1002_g
+ N_RESET_c_135_n N_RESET_c_136_n RESET RESET N_RESET_c_133_n
+ PM_SKY130_FD_SC_LP__BUSHOLD0_1%RESET
x_PM_SKY130_FD_SC_LP__BUSHOLD0_1%A_27_535# N_A_27_535#_M1005_s
+ N_A_27_535#_M1003_s N_A_27_535#_c_171_n N_A_27_535#_M1004_g
+ N_A_27_535#_c_178_n N_A_27_535#_M1001_g N_A_27_535#_c_172_n
+ N_A_27_535#_c_173_n N_A_27_535#_c_174_n N_A_27_535#_c_194_n
+ N_A_27_535#_c_196_n N_A_27_535#_c_175_n N_A_27_535#_c_179_n
+ N_A_27_535#_c_176_n N_A_27_535#_c_177_n
+ PM_SKY130_FD_SC_LP__BUSHOLD0_1%A_27_535#
x_PM_SKY130_FD_SC_LP__BUSHOLD0_1%VPWR N_VPWR_M1003_d N_VPWR_c_236_n
+ N_VPWR_c_237_n N_VPWR_c_238_n VPWR N_VPWR_c_239_n N_VPWR_c_235_n VPWR
+ PM_SKY130_FD_SC_LP__BUSHOLD0_1%VPWR
x_PM_SKY130_FD_SC_LP__BUSHOLD0_1%VGND N_VGND_M1005_d N_VGND_M1004_d
+ N_VGND_c_261_n N_VGND_c_262_n N_VGND_c_263_n N_VGND_c_264_n N_VGND_c_265_n
+ VGND N_VGND_c_266_n N_VGND_c_267_n VGND PM_SKY130_FD_SC_LP__BUSHOLD0_1%VGND
cc_1 VNB N_X_M1005_g 0.0630483f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.445
cc_2 VNB N_X_c_52_n 0.00167151f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.69
cc_3 VNB N_X_c_53_n 0.0149328f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.69
cc_4 VNB N_X_c_54_n 0.00231913f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=0.42
cc_5 VNB N_X_c_55_n 0.00141805f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=0.927
cc_6 VNB N_X_c_56_n 0.00477548f $X=-0.19 $Y=-0.245 $X2=1.525 $Y2=0.927
cc_7 VNB X 0.0334475f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_8 VNB N_X_c_58_n 0.0109864f $X=-0.19 $Y=-0.245 $X2=2.17 $Y2=1.015
cc_9 VNB N_RESET_M1000_g 0.0570323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB RESET 0.00167108f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.885
cc_11 VNB N_RESET_c_133_n 0.0139525f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.23
cc_12 VNB N_A_27_535#_c_171_n 0.0374571f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.525
cc_13 VNB N_A_27_535#_c_172_n 0.0284125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_535#_c_173_n 0.0385907f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.69
cc_15 VNB N_A_27_535#_c_174_n 0.0241611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_535#_c_175_n 0.0353116f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_17 VNB N_A_27_535#_c_176_n 0.0164984f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=2.32
cc_18 VNB N_A_27_535#_c_177_n 0.0605905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_235_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.69
cc_20 VNB N_VGND_c_261_n 0.00522139f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.445
cc_21 VNB N_VGND_c_262_n 0.0103405f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.23
cc_22 VNB N_VGND_c_263_n 0.0175269f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.885
cc_23 VNB N_VGND_c_264_n 0.0246812f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.525
cc_24 VNB N_VGND_c_265_n 0.00497572f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.065
cc_25 VNB N_VGND_c_266_n 0.0252348f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.45
cc_26 VNB N_VGND_c_267_n 0.157588f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=0.927
cc_27 VPB N_X_M1003_g 0.0411489f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.885
cc_28 VPB N_X_c_60_n 0.0282697f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.065
cc_29 VPB N_X_c_61_n 0.0177793f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.23
cc_30 VPB N_X_c_52_n 0.00124518f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.69
cc_31 VPB N_X_c_53_n 0.00265265f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.69
cc_32 VPB N_X_c_64_n 0.0232556f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=2.45
cc_33 VPB N_X_c_65_n 0.00512466f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=2.45
cc_34 VPB X 0.0371619f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_35 VPB X 0.00777251f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=2.32
cc_36 VPB X 0.0219272f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=2.69
cc_37 VPB N_RESET_M1002_g 0.0343164f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=1.525
cc_38 VPB N_RESET_c_135_n 0.0230674f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.23
cc_39 VPB N_RESET_c_136_n 0.0163411f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.885
cc_40 VPB RESET 0.00167108f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.885
cc_41 VPB N_RESET_c_133_n 0.00238864f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.23
cc_42 VPB N_A_27_535#_c_178_n 0.0565522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_27_535#_c_179_n 0.0133144f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.95
cc_44 VPB N_A_27_535#_c_176_n 0.0535154f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=2.32
cc_45 VPB N_A_27_535#_c_177_n 0.0653024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_236_n 0.00283171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_237_n 0.0256865f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.445
cc_48 VPB N_VPWR_c_238_n 0.00510915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_239_n 0.0378164f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.69
cc_50 VPB N_VPWR_c_235_n 0.0442239f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.69
cc_51 N_X_M1005_g N_RESET_M1000_g 0.0466991f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_52 N_X_c_54_n N_RESET_M1000_g 0.00292047f $X=1.36 $Y=0.42 $X2=0 $Y2=0
cc_53 N_X_c_56_n N_RESET_M1000_g 0.00304368f $X=1.525 $Y=0.927 $X2=0 $Y2=0
cc_54 N_X_c_61_n N_RESET_M1002_g 0.0254671f $X=0.65 $Y=2.23 $X2=0 $Y2=0
cc_55 N_X_c_52_n N_RESET_M1002_g 0.00102052f $X=0.65 $Y=1.69 $X2=0 $Y2=0
cc_56 N_X_c_64_n N_RESET_M1002_g 0.0114924f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_57 N_X_c_60_n N_RESET_c_135_n 0.0135694f $X=0.65 $Y=2.065 $X2=0 $Y2=0
cc_58 N_X_c_61_n N_RESET_c_136_n 0.0135694f $X=0.65 $Y=2.23 $X2=0 $Y2=0
cc_59 N_X_c_64_n N_RESET_c_136_n 0.00123898f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_60 N_X_c_52_n RESET 0.0423335f $X=0.65 $Y=1.69 $X2=0 $Y2=0
cc_61 N_X_c_53_n RESET 0.00232658f $X=0.65 $Y=1.69 $X2=0 $Y2=0
cc_62 N_X_c_64_n RESET 0.0256202f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_63 N_X_c_52_n N_RESET_c_133_n 0.00232658f $X=0.65 $Y=1.69 $X2=0 $Y2=0
cc_64 N_X_c_53_n N_RESET_c_133_n 0.0135694f $X=0.65 $Y=1.69 $X2=0 $Y2=0
cc_65 N_X_c_54_n N_A_27_535#_c_171_n 0.0158755f $X=1.36 $Y=0.42 $X2=0 $Y2=0
cc_66 N_X_c_64_n N_A_27_535#_c_178_n 0.0224084f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_67 X N_A_27_535#_c_178_n 0.00718359f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_68 N_X_c_54_n N_A_27_535#_c_172_n 0.00644612f $X=1.36 $Y=0.42 $X2=0 $Y2=0
cc_69 N_X_c_55_n N_A_27_535#_c_172_n 0.0205305f $X=2.025 $Y=0.927 $X2=0 $Y2=0
cc_70 N_X_c_56_n N_A_27_535#_c_172_n 0.00203562f $X=1.525 $Y=0.927 $X2=0 $Y2=0
cc_71 N_X_M1005_g N_A_27_535#_c_173_n 0.0133024f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_72 N_X_c_54_n N_A_27_535#_c_173_n 0.00614532f $X=1.36 $Y=0.42 $X2=0 $Y2=0
cc_73 N_X_c_56_n N_A_27_535#_c_173_n 0.0062567f $X=1.525 $Y=0.927 $X2=0 $Y2=0
cc_74 N_X_M1005_g N_A_27_535#_c_174_n 0.0168724f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_75 N_X_c_55_n N_A_27_535#_c_174_n 0.00566377f $X=2.025 $Y=0.927 $X2=0 $Y2=0
cc_76 N_X_c_56_n N_A_27_535#_c_174_n 0.0253377f $X=1.525 $Y=0.927 $X2=0 $Y2=0
cc_77 N_X_c_55_n N_A_27_535#_c_194_n 0.0190819f $X=2.025 $Y=0.927 $X2=0 $Y2=0
cc_78 X N_A_27_535#_c_194_n 0.0141259f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_79 N_X_c_64_n N_A_27_535#_c_196_n 0.0188915f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_80 X N_A_27_535#_c_196_n 0.0644409f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_81 N_X_M1005_g N_A_27_535#_c_175_n 0.00604826f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_82 N_X_c_52_n N_A_27_535#_c_175_n 0.0260863f $X=0.65 $Y=1.69 $X2=0 $Y2=0
cc_83 N_X_c_53_n N_A_27_535#_c_175_n 0.00111169f $X=0.65 $Y=1.69 $X2=0 $Y2=0
cc_84 N_X_M1003_g N_A_27_535#_c_179_n 0.00680076f $X=0.74 $Y=2.885 $X2=0 $Y2=0
cc_85 N_X_M1005_g N_A_27_535#_c_176_n 0.00509974f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_86 N_X_M1003_g N_A_27_535#_c_176_n 0.00686558f $X=0.74 $Y=2.885 $X2=0 $Y2=0
cc_87 N_X_c_52_n N_A_27_535#_c_176_n 0.0650573f $X=0.65 $Y=1.69 $X2=0 $Y2=0
cc_88 N_X_c_53_n N_A_27_535#_c_176_n 0.0158776f $X=0.65 $Y=1.69 $X2=0 $Y2=0
cc_89 N_X_c_65_n N_A_27_535#_c_176_n 0.0146597f $X=0.815 $Y=2.45 $X2=0 $Y2=0
cc_90 N_X_c_64_n N_A_27_535#_c_177_n 0.0144293f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_91 N_X_c_55_n N_A_27_535#_c_177_n 0.0132019f $X=2.025 $Y=0.927 $X2=0 $Y2=0
cc_92 X N_A_27_535#_c_177_n 0.0452244f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_93 N_X_M1003_g N_VPWR_c_236_n 0.00325608f $X=0.74 $Y=2.885 $X2=0 $Y2=0
cc_94 N_X_c_64_n N_VPWR_c_236_n 0.0205709f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_95 N_X_M1003_g N_VPWR_c_237_n 0.00585385f $X=0.74 $Y=2.885 $X2=0 $Y2=0
cc_96 X N_VPWR_c_239_n 0.0165867f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_97 N_X_M1001_d N_VPWR_c_235_n 0.00230893f $X=2 $Y=2.675 $X2=0 $Y2=0
cc_98 N_X_M1003_g N_VPWR_c_235_n 0.00753316f $X=0.74 $Y=2.885 $X2=0 $Y2=0
cc_99 N_X_c_64_n N_VPWR_c_235_n 0.0282627f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_100 N_X_c_65_n N_VPWR_c_235_n 0.0123558f $X=0.815 $Y=2.45 $X2=0 $Y2=0
cc_101 X N_VPWR_c_235_n 0.0110608f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_102 N_X_M1005_g N_VGND_c_261_n 0.00319241f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_103 N_X_c_54_n N_VGND_c_263_n 0.012019f $X=1.36 $Y=0.42 $X2=0 $Y2=0
cc_104 N_X_c_55_n N_VGND_c_263_n 0.00199564f $X=2.025 $Y=0.927 $X2=0 $Y2=0
cc_105 N_X_c_58_n N_VGND_c_263_n 0.0184241f $X=2.17 $Y=1.015 $X2=0 $Y2=0
cc_106 N_X_M1005_g N_VGND_c_264_n 0.00585385f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_107 N_X_c_54_n N_VGND_c_266_n 0.0171073f $X=1.36 $Y=0.42 $X2=0 $Y2=0
cc_108 N_X_M1000_d N_VGND_c_267_n 0.00240953f $X=1.22 $Y=0.235 $X2=0 $Y2=0
cc_109 N_X_M1005_g N_VGND_c_267_n 0.0117375f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_110 N_X_c_54_n N_VGND_c_267_n 0.0114026f $X=1.36 $Y=0.42 $X2=0 $Y2=0
cc_111 N_X_c_55_n N_VGND_c_267_n 0.0125445f $X=2.025 $Y=0.927 $X2=0 $Y2=0
cc_112 N_X_c_58_n N_VGND_c_267_n 0.00161861f $X=2.17 $Y=1.015 $X2=0 $Y2=0
cc_113 N_RESET_M1000_g N_A_27_535#_c_171_n 0.0211178f $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_114 N_RESET_M1002_g N_A_27_535#_c_178_n 0.0561123f $X=1.215 $Y=2.885 $X2=0
+ $Y2=0
cc_115 N_RESET_M1000_g N_A_27_535#_c_174_n 0.0153288f $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_116 RESET N_A_27_535#_c_174_n 0.0256202f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_117 N_RESET_c_133_n N_A_27_535#_c_174_n 0.00123898f $X=1.19 $Y=1.69 $X2=0
+ $Y2=0
cc_118 N_RESET_M1000_g N_A_27_535#_c_196_n 9.37527e-19 $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_119 RESET N_A_27_535#_c_196_n 0.0361219f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_120 N_RESET_c_133_n N_A_27_535#_c_196_n 0.00219599f $X=1.19 $Y=1.69 $X2=0
+ $Y2=0
cc_121 N_RESET_M1000_g N_A_27_535#_c_177_n 0.0215869f $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_122 N_RESET_M1002_g N_A_27_535#_c_177_n 0.011358f $X=1.215 $Y=2.885 $X2=0
+ $Y2=0
cc_123 RESET N_A_27_535#_c_177_n 0.00252912f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_124 N_RESET_c_133_n N_A_27_535#_c_177_n 0.0419327f $X=1.19 $Y=1.69 $X2=0
+ $Y2=0
cc_125 N_RESET_M1002_g N_VPWR_c_236_n 0.0117776f $X=1.215 $Y=2.885 $X2=0 $Y2=0
cc_126 N_RESET_M1002_g N_VPWR_c_239_n 0.00486043f $X=1.215 $Y=2.885 $X2=0 $Y2=0
cc_127 N_RESET_M1002_g N_VPWR_c_235_n 0.00435698f $X=1.215 $Y=2.885 $X2=0 $Y2=0
cc_128 N_RESET_M1000_g N_VGND_c_261_n 0.00313081f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_129 N_RESET_M1000_g N_VGND_c_266_n 0.00585385f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_130 N_RESET_M1000_g N_VGND_c_267_n 0.010696f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_27_535#_c_178_n N_VPWR_c_236_n 0.00325895f $X=1.75 $Y=2.655 $X2=0
+ $Y2=0
cc_132 N_A_27_535#_c_179_n N_VPWR_c_237_n 0.0202039f $X=0.26 $Y=2.885 $X2=0
+ $Y2=0
cc_133 N_A_27_535#_c_178_n N_VPWR_c_239_n 0.0195128f $X=1.75 $Y=2.655 $X2=0
+ $Y2=0
cc_134 N_A_27_535#_M1003_s N_VPWR_c_235_n 0.00758182f $X=0.135 $Y=2.675 $X2=0
+ $Y2=0
cc_135 N_A_27_535#_c_178_n N_VPWR_c_235_n 0.0182509f $X=1.75 $Y=2.655 $X2=0
+ $Y2=0
cc_136 N_A_27_535#_c_179_n N_VPWR_c_235_n 0.0128998f $X=0.26 $Y=2.885 $X2=0
+ $Y2=0
cc_137 N_A_27_535#_c_174_n N_VGND_c_261_n 0.00717784f $X=1.605 $Y=1.27 $X2=0
+ $Y2=0
cc_138 N_A_27_535#_c_171_n N_VGND_c_263_n 0.0170555f $X=1.75 $Y=0.725 $X2=0
+ $Y2=0
cc_139 N_A_27_535#_c_173_n N_VGND_c_264_n 0.0188755f $X=0.5 $Y=0.42 $X2=0 $Y2=0
cc_140 N_A_27_535#_c_171_n N_VGND_c_266_n 0.0181551f $X=1.75 $Y=0.725 $X2=0
+ $Y2=0
cc_141 N_A_27_535#_M1005_s N_VGND_c_267_n 0.0026734f $X=0.375 $Y=0.235 $X2=0
+ $Y2=0
cc_142 N_A_27_535#_c_171_n N_VGND_c_267_n 0.0156372f $X=1.75 $Y=0.725 $X2=0
+ $Y2=0
cc_143 N_A_27_535#_c_173_n N_VGND_c_267_n 0.0111968f $X=0.5 $Y=0.42 $X2=0 $Y2=0
cc_144 N_VPWR_c_235_n A_258_535# 0.0029401f $X=2.16 $Y=3.33 $X2=-0.19 $Y2=-0.245
