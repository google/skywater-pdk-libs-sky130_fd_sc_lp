* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor2_lp A B VGND VNB VPB VPWR Y
X0 a_280_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 Y B a_280_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_510_125# B a_82_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_112_92# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_82_66# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VGND B a_112_92# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_82_66# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 VGND A a_510_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Y a_82_66# a_112_92# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR A a_82_66# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
