* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or2_0 A B VGND VNB VPB VPWR X
M1000 a_159_473# B a_76_473# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.113e+11p ps=1.37e+06u
M1001 X a_76_473# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=3.627e+11p ps=2.52e+06u
M1002 a_76_473# B VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.289e+11p ps=2.77e+06u
M1003 VPWR A a_159_473# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A a_76_473# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_76_473# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends
