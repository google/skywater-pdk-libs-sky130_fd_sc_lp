* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
X0 a_27_463# a_306_277# a_336_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR CLK_N a_306_277# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_294_35# a_306_277# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_336_463# a_294_35# a_447_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND RESET_B a_142_121# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_540_123# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND RESET_B a_1465_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1099_447# a_306_277# a_1229_531# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1275_125# a_1287_276# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_1832_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_294_35# a_306_277# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VPWR a_336_463# a_501_229# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 a_438_123# a_501_229# a_540_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1832_367# a_1099_447# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_27_463# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VPWR D a_27_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VPWR RESET_B a_1287_276# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_1099_447# a_294_35# a_1275_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1287_276# a_1099_447# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_142_121# D a_27_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_336_463# a_501_229# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_501_229# a_306_277# a_1099_447# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_27_463# a_294_35# a_336_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_306_277# CLK_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_1229_531# a_1287_276# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VPWR RESET_B a_336_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_336_463# a_306_277# a_438_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_1465_125# a_1099_447# a_1287_276# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_447_463# a_501_229# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_501_229# a_294_35# a_1099_447# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X30 a_1832_367# a_1099_447# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VGND a_1832_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
