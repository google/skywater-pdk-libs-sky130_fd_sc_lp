* File: sky130_fd_sc_lp__dfbbn_1.pxi.spice
* Created: Wed Sep  2 09:42:54 2020
* 
x_PM_SKY130_FD_SC_LP__DFBBN_1%CLK_N N_CLK_N_M1029_g N_CLK_N_M1027_g CLK_N CLK_N
+ CLK_N N_CLK_N_c_281_n N_CLK_N_c_282_n PM_SKY130_FD_SC_LP__DFBBN_1%CLK_N
x_PM_SKY130_FD_SC_LP__DFBBN_1%D N_D_c_303_n N_D_c_304_n N_D_c_305_n N_D_c_309_n
+ N_D_M1008_g N_D_c_306_n N_D_M1022_g N_D_c_310_n D N_D_c_307_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%D
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_113_67# N_A_113_67#_M1029_d N_A_113_67#_M1027_d
+ N_A_113_67#_M1009_g N_A_113_67#_M1032_g N_A_113_67#_c_357_n
+ N_A_113_67#_c_358_n N_A_113_67#_c_378_n N_A_113_67#_c_379_n
+ N_A_113_67#_M1036_g N_A_113_67#_M1038_g N_A_113_67#_M1025_g
+ N_A_113_67#_c_381_n N_A_113_67#_M1039_g N_A_113_67#_c_382_n
+ N_A_113_67#_c_360_n N_A_113_67#_c_383_n N_A_113_67#_c_384_n
+ N_A_113_67#_c_361_n N_A_113_67#_c_362_n N_A_113_67#_c_363_n
+ N_A_113_67#_c_364_n N_A_113_67#_c_365_n N_A_113_67#_c_366_n
+ N_A_113_67#_c_367_n N_A_113_67#_c_368_n N_A_113_67#_c_369_n
+ N_A_113_67#_c_370_n N_A_113_67#_c_387_n N_A_113_67#_c_388_n
+ N_A_113_67#_c_389_n N_A_113_67#_c_390_n N_A_113_67#_c_391_n
+ N_A_113_67#_c_371_n N_A_113_67#_c_372_n N_A_113_67#_c_373_n
+ N_A_113_67#_c_392_n N_A_113_67#_c_374_n N_A_113_67#_c_375_n
+ N_A_113_67#_c_376_n PM_SKY130_FD_SC_LP__DFBBN_1%A_113_67#
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_755_398# N_A_755_398#_M1017_d
+ N_A_755_398#_M1037_d N_A_755_398#_c_615_n N_A_755_398#_M1010_g
+ N_A_755_398#_M1031_g N_A_755_398#_c_608_n N_A_755_398#_M1004_g
+ N_A_755_398#_M1005_g N_A_755_398#_c_619_n N_A_755_398#_c_649_p
+ N_A_755_398#_c_716_p N_A_755_398#_c_650_p N_A_755_398#_c_651_p
+ N_A_755_398#_c_610_n N_A_755_398#_c_659_p N_A_755_398#_c_611_n
+ N_A_755_398#_c_620_n N_A_755_398#_c_612_n N_A_755_398#_c_613_n
+ N_A_755_398#_c_614_n N_A_755_398#_c_623_n N_A_755_398#_c_624_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%A_755_398#
x_PM_SKY130_FD_SC_LP__DFBBN_1%SET_B N_SET_B_M1024_g N_SET_B_M1037_g
+ N_SET_B_M1026_g N_SET_B_c_769_n N_SET_B_c_770_n N_SET_B_M1015_g
+ N_SET_B_c_771_n SET_B N_SET_B_c_762_n N_SET_B_c_763_n N_SET_B_c_764_n
+ N_SET_B_c_765_n N_SET_B_c_766_n N_SET_B_c_767_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%SET_B
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_546_449# N_A_546_449#_M1023_d
+ N_A_546_449#_M1036_d N_A_546_449#_M1017_g N_A_546_449#_M1003_g
+ N_A_546_449#_c_901_n N_A_546_449#_c_911_n N_A_546_449#_c_902_n
+ N_A_546_449#_c_903_n N_A_546_449#_c_904_n N_A_546_449#_c_905_n
+ N_A_546_449#_c_958_n N_A_546_449#_c_914_n N_A_546_449#_c_915_n
+ N_A_546_449#_c_906_n N_A_546_449#_c_917_n N_A_546_449#_c_907_n
+ N_A_546_449#_c_908_n N_A_546_449#_c_919_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%A_546_449#
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_223_119# N_A_223_119#_M1009_s
+ N_A_223_119#_M1032_s N_A_223_119#_M1023_g N_A_223_119#_c_1056_n
+ N_A_223_119#_c_1057_n N_A_223_119#_c_1058_n N_A_223_119#_M1033_g
+ N_A_223_119#_c_1060_n N_A_223_119#_c_1061_n N_A_223_119#_M1021_g
+ N_A_223_119#_c_1063_n N_A_223_119#_c_1064_n N_A_223_119#_c_1047_n
+ N_A_223_119#_c_1048_n N_A_223_119#_c_1049_n N_A_223_119#_c_1050_n
+ N_A_223_119#_M1018_g N_A_223_119#_c_1051_n N_A_223_119#_c_1052_n
+ N_A_223_119#_c_1068_n N_A_223_119#_c_1069_n N_A_223_119#_c_1053_n
+ N_A_223_119#_c_1070_n N_A_223_119#_c_1054_n N_A_223_119#_c_1055_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%A_223_119#
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_1741_137# N_A_1741_137#_M1001_d
+ N_A_1741_137#_M1015_d N_A_1741_137#_c_1212_n N_A_1741_137#_M1006_g
+ N_A_1741_137#_M1000_g N_A_1741_137#_M1030_g N_A_1741_137#_M1011_g
+ N_A_1741_137#_c_1214_n N_A_1741_137#_c_1215_n N_A_1741_137#_M1034_g
+ N_A_1741_137#_M1019_g N_A_1741_137#_c_1217_n N_A_1741_137#_c_1218_n
+ N_A_1741_137#_c_1228_n N_A_1741_137#_c_1229_n N_A_1741_137#_c_1260_n
+ N_A_1741_137#_c_1230_n N_A_1741_137#_c_1219_n N_A_1741_137#_c_1232_n
+ N_A_1741_137#_c_1220_n N_A_1741_137#_c_1234_n N_A_1741_137#_c_1269_p
+ N_A_1741_137#_c_1292_p N_A_1741_137#_c_1221_n N_A_1741_137#_c_1222_n
+ N_A_1741_137#_c_1223_n N_A_1741_137#_c_1224_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%A_1741_137#
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_1531_428# N_A_1531_428#_M1025_d
+ N_A_1531_428#_M1021_d N_A_1531_428#_M1001_g N_A_1531_428#_M1028_g
+ N_A_1531_428#_c_1389_n N_A_1531_428#_c_1381_n N_A_1531_428#_c_1382_n
+ N_A_1531_428#_c_1383_n N_A_1531_428#_c_1384_n N_A_1531_428#_c_1385_n
+ N_A_1531_428#_c_1386_n N_A_1531_428#_c_1387_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%A_1531_428#
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_1186_21# N_A_1186_21#_M1002_s
+ N_A_1186_21#_M1007_s N_A_1186_21#_M1012_g N_A_1186_21#_c_1477_n
+ N_A_1186_21#_c_1478_n N_A_1186_21#_c_1479_n N_A_1186_21#_c_1480_n
+ N_A_1186_21#_M1020_g N_A_1186_21#_M1014_g N_A_1186_21#_c_1490_n
+ N_A_1186_21#_M1013_g N_A_1186_21#_c_1483_n N_A_1186_21#_c_1484_n
+ N_A_1186_21#_c_1485_n N_A_1186_21#_c_1492_n N_A_1186_21#_c_1486_n
+ N_A_1186_21#_c_1487_n N_A_1186_21#_c_1494_n N_A_1186_21#_c_1495_n
+ N_A_1186_21#_c_1488_n PM_SKY130_FD_SC_LP__DFBBN_1%A_1186_21#
x_PM_SKY130_FD_SC_LP__DFBBN_1%RESET_B N_RESET_B_M1002_g N_RESET_B_M1007_g
+ RESET_B N_RESET_B_c_1598_n N_RESET_B_c_1599_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%RESET_B
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_2511_137# N_A_2511_137#_M1034_s
+ N_A_2511_137#_M1019_s N_A_2511_137#_M1035_g N_A_2511_137#_M1016_g
+ N_A_2511_137#_c_1630_n N_A_2511_137#_c_1635_n N_A_2511_137#_c_1631_n
+ N_A_2511_137#_c_1632_n N_A_2511_137#_c_1633_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%A_2511_137#
x_PM_SKY130_FD_SC_LP__DFBBN_1%VPWR N_VPWR_M1027_s N_VPWR_M1032_d N_VPWR_M1010_d
+ N_VPWR_M1020_d N_VPWR_M1000_d N_VPWR_M1013_d N_VPWR_M1007_d N_VPWR_M1019_d
+ N_VPWR_c_1678_n N_VPWR_c_1679_n N_VPWR_c_1680_n N_VPWR_c_1681_n
+ N_VPWR_c_1682_n N_VPWR_c_1683_n N_VPWR_c_1684_n N_VPWR_c_1685_n
+ N_VPWR_c_1686_n N_VPWR_c_1687_n N_VPWR_c_1688_n N_VPWR_c_1689_n
+ N_VPWR_c_1690_n N_VPWR_c_1691_n N_VPWR_c_1692_n VPWR N_VPWR_c_1693_n
+ N_VPWR_c_1694_n N_VPWR_c_1695_n N_VPWR_c_1696_n N_VPWR_c_1697_n
+ N_VPWR_c_1677_n N_VPWR_c_1699_n N_VPWR_c_1700_n N_VPWR_c_1701_n
+ N_VPWR_c_1702_n PM_SKY130_FD_SC_LP__DFBBN_1%VPWR
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_460_449# N_A_460_449#_M1022_d
+ N_A_460_449#_M1008_d N_A_460_449#_c_1820_n N_A_460_449#_c_1821_n
+ N_A_460_449#_c_1824_n N_A_460_449#_c_1822_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%A_460_449#
x_PM_SKY130_FD_SC_LP__DFBBN_1%Q_N N_Q_N_M1030_d N_Q_N_M1011_d N_Q_N_c_1872_n
+ N_Q_N_c_1873_n N_Q_N_c_1875_n N_Q_N_c_1874_n Q_N Q_N Q_N
+ PM_SKY130_FD_SC_LP__DFBBN_1%Q_N
x_PM_SKY130_FD_SC_LP__DFBBN_1%Q N_Q_M1035_d N_Q_M1016_d N_Q_c_1910_n
+ N_Q_c_1911_n N_Q_c_1907_n Q Q N_Q_c_1909_n Q PM_SKY130_FD_SC_LP__DFBBN_1%Q
x_PM_SKY130_FD_SC_LP__DFBBN_1%VGND N_VGND_M1029_s N_VGND_M1009_d N_VGND_M1031_d
+ N_VGND_M1005_s N_VGND_M1006_d N_VGND_M1002_d N_VGND_M1034_d N_VGND_c_1930_n
+ N_VGND_c_1931_n N_VGND_c_1932_n N_VGND_c_1933_n N_VGND_c_1934_n
+ N_VGND_c_1935_n N_VGND_c_1936_n N_VGND_c_1937_n N_VGND_c_1938_n
+ N_VGND_c_1939_n N_VGND_c_1940_n N_VGND_c_1941_n VGND N_VGND_c_1942_n
+ N_VGND_c_1943_n N_VGND_c_1944_n N_VGND_c_1945_n N_VGND_c_1946_n
+ N_VGND_c_1947_n N_VGND_c_1948_n N_VGND_c_1949_n N_VGND_c_1950_n
+ N_VGND_c_1951_n PM_SKY130_FD_SC_LP__DFBBN_1%VGND
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_1013_66# N_A_1013_66#_M1024_d
+ N_A_1013_66#_M1012_d N_A_1013_66#_c_2066_n N_A_1013_66#_c_2059_n
+ N_A_1013_66#_c_2064_n PM_SKY130_FD_SC_LP__DFBBN_1%A_1013_66#
x_PM_SKY130_FD_SC_LP__DFBBN_1%A_1896_119# N_A_1896_119#_M1026_d
+ N_A_1896_119#_M1014_d N_A_1896_119#_c_2086_n N_A_1896_119#_c_2087_n
+ N_A_1896_119#_c_2088_n N_A_1896_119#_c_2089_n
+ PM_SKY130_FD_SC_LP__DFBBN_1%A_1896_119#
cc_1 VNB N_CLK_N_M1029_g 0.0320033f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.545
cc_2 VNB N_CLK_N_M1027_g 0.00176087f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.725
cc_3 VNB N_CLK_N_c_281_n 0.0979208f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_4 VNB N_CLK_N_c_282_n 0.00572117f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_5 VNB N_D_c_303_n 0.0419615f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.955
cc_6 VNB N_D_c_304_n 0.00797105f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.545
cc_7 VNB N_D_c_305_n 0.0260713f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.545
cc_8 VNB N_D_c_306_n 0.0159307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_D_c_307_n 0.00839529f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_10 VNB N_A_113_67#_M1009_g 0.0371364f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB N_A_113_67#_c_357_n 0.149962f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.12
cc_12 VNB N_A_113_67#_c_358_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_13 VNB N_A_113_67#_M1038_g 0.0320059f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.035
cc_14 VNB N_A_113_67#_c_360_n 0.00136476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_113_67#_c_361_n 0.0494568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_113_67#_c_362_n 0.044249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_113_67#_c_363_n 0.0044511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_113_67#_c_364_n 0.00240362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_113_67#_c_365_n 0.0139653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_113_67#_c_366_n 0.00199013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_113_67#_c_367_n 0.0142191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_113_67#_c_368_n 0.00925362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_113_67#_c_369_n 0.00105008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_113_67#_c_370_n 0.00825304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_113_67#_c_371_n 0.0104635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_113_67#_c_372_n 0.00921001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_113_67#_c_373_n 0.00809138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_113_67#_c_374_n 0.0224609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_113_67#_c_375_n 0.0680099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_113_67#_c_376_n 0.0198839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_755_398#_M1031_g 0.0564711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_755_398#_c_608_n 0.0233465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_755_398#_M1005_g 0.0210529f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_34 VNB N_A_755_398#_c_610_n 0.00330454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_755_398#_c_611_n 0.00323308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_755_398#_c_612_n 0.00126966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_755_398#_c_613_n 0.00337175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_755_398#_c_614_n 0.00703299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_SET_B_M1024_g 0.0419489f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.545
cc_40 VNB N_SET_B_M1026_g 0.0237568f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_41 VNB SET_B 0.00589365f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_42 VNB N_SET_B_c_762_n 0.014964f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_43 VNB N_SET_B_c_763_n 6.81341e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_SET_B_c_764_n 0.00123986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_SET_B_c_765_n 0.0234283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_SET_B_c_766_n 0.00424424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_SET_B_c_767_n 0.0133434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_546_449#_M1017_g 0.0375209f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_49 VNB N_A_546_449#_c_901_n 0.0114516f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_50 VNB N_A_546_449#_c_902_n 4.7162e-19 $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_51 VNB N_A_546_449#_c_903_n 0.0159305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_546_449#_c_904_n 0.00228237f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_53 VNB N_A_546_449#_c_905_n 0.00163477f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_54 VNB N_A_546_449#_c_906_n 0.00113099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_546_449#_c_907_n 0.0464728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_546_449#_c_908_n 0.00347569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_223_119#_M1023_g 0.0373527f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_58 VNB N_A_223_119#_c_1047_n 0.0119617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_223_119#_c_1048_n 0.0238153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_223_119#_c_1049_n 0.00823124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_223_119#_c_1050_n 0.0153732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_223_119#_c_1051_n 0.0199525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_223_119#_c_1052_n 0.00629432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_223_119#_c_1053_n 0.001848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_223_119#_c_1054_n 0.00264715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_223_119#_c_1055_n 0.00944102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1741_137#_c_1212_n 0.0148407f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=2.725
cc_68 VNB N_A_1741_137#_M1011_g 0.00105396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1741_137#_c_1214_n 0.057322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1741_137#_c_1215_n 0.0183925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1741_137#_M1019_g 0.0176658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1741_137#_c_1217_n 0.0201028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1741_137#_c_1218_n 0.00545278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1741_137#_c_1219_n 0.00780338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1741_137#_c_1220_n 2.80413e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1741_137#_c_1221_n 0.00420852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1741_137#_c_1222_n 0.0119783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1741_137#_c_1223_n 0.0308271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1741_137#_c_1224_n 0.022685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1531_428#_M1001_g 0.0231662f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_81 VNB N_A_1531_428#_c_1381_n 0.00865036f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=1.12
cc_82 VNB N_A_1531_428#_c_1382_n 0.0119644f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.035
cc_83 VNB N_A_1531_428#_c_1383_n 0.00151555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1531_428#_c_1384_n 0.00194526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1531_428#_c_1385_n 7.20997e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1531_428#_c_1386_n 0.00147634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1531_428#_c_1387_n 0.0227393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1186_21#_M1012_g 0.00558136f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_89 VNB N_A_1186_21#_c_1477_n 0.338708f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_90 VNB N_A_1186_21#_c_1478_n 0.0118327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1186_21#_c_1479_n 0.0294239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1186_21#_c_1480_n 0.00716914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1186_21#_M1020_g 0.0240485f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_94 VNB N_A_1186_21#_M1014_g 0.0145337f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_95 VNB N_A_1186_21#_c_1483_n 0.0179221f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.035
cc_96 VNB N_A_1186_21#_c_1484_n 0.0100796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1186_21#_c_1485_n 0.00866839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1186_21#_c_1486_n 0.0152594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1186_21#_c_1487_n 0.00193209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1186_21#_c_1488_n 0.041276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_RESET_B_M1007_g 0.00123868f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.725
cc_102 VNB RESET_B 0.0072784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_RESET_B_c_1598_n 0.0282557f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_104 VNB N_RESET_B_c_1599_n 0.0197197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2511_137#_M1035_g 0.0292121f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_106 VNB N_A_2511_137#_M1016_g 0.00114141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2511_137#_c_1630_n 0.00388384f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=1.12
cc_108 VNB N_A_2511_137#_c_1631_n 0.00708653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2511_137#_c_1632_n 0.0344463f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.035
cc_110 VNB N_A_2511_137#_c_1633_n 0.00248805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VPWR_c_1677_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_460_449#_c_1820_n 0.0022778f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_113 VNB N_A_460_449#_c_1821_n 0.0025387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_460_449#_c_1822_n 0.00589038f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=1.12
cc_115 VNB N_Q_N_c_1872_n 0.0106682f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_116 VNB N_Q_N_c_1873_n 0.00289167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_Q_N_c_1874_n 0.00515846f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_118 VNB N_Q_c_1907_n 0.0250313f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.12
cc_119 VNB Q 0.0126596f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_120 VNB N_Q_c_1909_n 0.0287706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1930_n 0.0105185f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_122 VNB N_VGND_c_1931_n 0.0286338f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_123 VNB N_VGND_c_1932_n 0.0150651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1933_n 0.0120256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1934_n 0.0117815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1935_n 0.0229387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1936_n 0.0168508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1937_n 0.0152123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1938_n 0.0672053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1939_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1940_n 0.0553869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1941_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1942_n 0.0338008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1943_n 0.054773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1944_n 0.0572163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1945_n 0.0344484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1946_n 0.0187754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1947_n 0.717459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1948_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1949_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1950_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1951_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_1013_66#_c_2059_n 0.00448151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_1896_119#_c_2086_n 0.00267609f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_145 VNB N_A_1896_119#_c_2087_n 0.00823192f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_146 VNB N_A_1896_119#_c_2088_n 0.00408722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_1896_119#_c_2089_n 0.0151349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VPB N_CLK_N_M1027_g 0.0675323f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.725
cc_149 VPB N_CLK_N_c_282_n 0.0232389f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_150 VPB N_D_c_304_n 0.020057f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.545
cc_151 VPB N_D_c_309_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.625
cc_152 VPB N_D_c_310_n 0.0280654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_113_67#_M1032_g 0.0289613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_113_67#_c_378_n 0.076227f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_155 VPB N_A_113_67#_c_379_n 0.0130423f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=0.955
cc_156 VPB N_A_113_67#_M1036_g 0.0348794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_113_67#_c_381_n 0.0194056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_113_67#_c_382_n 0.0347325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_113_67#_c_383_n 0.0222167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_113_67#_c_384_n 0.00220155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_113_67#_c_361_n 0.0141661f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_113_67#_c_370_n 0.00275943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_113_67#_c_387_n 0.0041844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_113_67#_c_388_n 0.00763822f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_113_67#_c_389_n 0.00192422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_113_67#_c_390_n 0.00388454f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_113_67#_c_391_n 0.049662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_113_67#_c_392_n 0.00125702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_113_67#_c_374_n 0.00640373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_113_67#_c_375_n 0.0611419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_755_398#_c_615_n 0.0177181f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.725
cc_172 VPB N_A_755_398#_M1031_g 0.00536732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_755_398#_c_608_n 0.0118431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_755_398#_M1004_g 0.0199714f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_175 VPB N_A_755_398#_c_619_n 0.00405338f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.665
cc_176 VPB N_A_755_398#_c_620_n 0.00429896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_755_398#_c_612_n 9.54123e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_755_398#_c_613_n 0.00289718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_755_398#_c_623_n 0.00285448f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_755_398#_c_624_n 0.0750783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_SET_B_M1037_g 0.0238422f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.725
cc_182 VPB N_SET_B_c_769_n 0.0128672f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_SET_B_c_770_n 0.0166356f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.12
cc_184 VPB N_SET_B_c_771_n 0.0236785f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_185 VPB SET_B 0.00721479f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.295
cc_186 VPB N_SET_B_c_762_n 0.0325696f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.665
cc_187 VPB N_SET_B_c_763_n 0.00134298f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_SET_B_c_764_n 0.00254874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_SET_B_c_765_n 0.0111757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_SET_B_c_766_n 0.00138662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_SET_B_c_767_n 0.0150079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_546_449#_M1003_g 0.0223817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_546_449#_c_901_n 0.00475902f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_194 VPB N_A_546_449#_c_911_n 0.00486065f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_195 VPB N_A_546_449#_c_902_n 0.00392785f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_196 VPB N_A_546_449#_c_905_n 0.00561856f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.665
cc_197 VPB N_A_546_449#_c_914_n 0.002616f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=2.035
cc_198 VPB N_A_546_449#_c_915_n 0.00389173f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_546_449#_c_906_n 2.8428e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_546_449#_c_917_n 0.00102307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_546_449#_c_907_n 0.0192506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_546_449#_c_919_n 0.00615795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_223_119#_c_1056_n 0.0135504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_223_119#_c_1057_n 0.0281061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_223_119#_c_1058_n 0.0132768f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_223_119#_M1033_g 0.0385361f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=0.955
cc_207 VPB N_A_223_119#_c_1060_n 0.320682f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.625
cc_208 VPB N_A_223_119#_c_1061_n 0.0119033f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_209 VPB N_A_223_119#_M1021_g 0.0103807f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.665
cc_210 VPB N_A_223_119#_c_1063_n 0.0303276f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_223_119#_c_1064_n 0.00720376f $X=-0.19 $Y=1.655 $X2=0.28
+ $Y2=2.035
cc_212 VPB N_A_223_119#_c_1047_n 0.0166665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_223_119#_c_1051_n 0.0207303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_223_119#_c_1052_n 0.0291904f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_223_119#_c_1068_n 0.00387725f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_223_119#_c_1069_n 0.00974231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_223_119#_c_1070_n 0.0134351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_223_119#_c_1054_n 0.00113365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1741_137#_M1000_g 0.0252516f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_1741_137#_M1011_g 0.0262959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_1741_137#_M1019_g 0.0257009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_1741_137#_c_1228_n 0.00644791f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_1741_137#_c_1229_n 0.0339934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_1741_137#_c_1230_n 0.00408807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1741_137#_c_1219_n 0.00802394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_1741_137#_c_1232_n 0.0263393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_1741_137#_c_1220_n 0.00173733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_1741_137#_c_1234_n 0.00302308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_1741_137#_c_1222_n 0.0214239f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_1531_428#_M1028_g 0.0359044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_1531_428#_c_1389_n 0.00244956f $X=-0.19 $Y=1.655 $X2=0.342
+ $Y2=1.12
cc_232 VPB N_A_1531_428#_c_1384_n 0.00364636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_1531_428#_c_1386_n 0.00102512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_1531_428#_c_1387_n 0.0169443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_1186_21#_M1020_g 0.021241f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_236 VPB N_A_1186_21#_c_1490_n 0.0165555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_1186_21#_c_1485_n 0.0196904f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_1186_21#_c_1492_n 0.0298429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_1186_21#_c_1487_n 0.0019898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_1186_21#_c_1494_n 0.00351305f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_1186_21#_c_1495_n 0.010603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_RESET_B_M1007_g 0.0284531f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.725
cc_243 VPB N_A_2511_137#_M1016_g 0.0281049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_2511_137#_c_1635_n 0.00641237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1678_n 0.0113568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1679_n 0.0336858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1680_n 0.0109364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1681_n 0.0224016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1682_n 0.0143437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1683_n 0.00686995f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1684_n 0.0234361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1685_n 0.0254247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1686_n 0.0188927f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1687_n 0.0338092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1688_n 0.00522307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1689_n 0.076882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1690_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1691_n 0.0267309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1692_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1693_n 0.0531593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1694_n 0.0560467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1695_n 0.0228482f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1696_n 0.0333948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1697_n 0.0187754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1677_n 0.148098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1699_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1700_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1701_n 0.00601829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1702_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_460_449#_c_1821_n 0.00736134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_460_449#_c_1824_n 0.0028426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_Q_N_c_1875_n 0.00492543f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_273 VPB N_Q_N_c_1874_n 0.00299801f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.12
cc_274 VPB Q_N 0.0209594f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=0.955
cc_275 VPB N_Q_c_1910_n 0.0423813f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_276 VPB N_Q_c_1911_n 0.0126596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_Q_c_1907_n 0.00769959f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.12
cc_278 N_CLK_N_M1027_g N_A_113_67#_c_360_n 0.0203015f $X=0.495 $Y=2.725 $X2=0
+ $Y2=0
cc_279 N_CLK_N_M1029_g N_A_113_67#_c_371_n 0.00784668f $X=0.49 $Y=0.545 $X2=0
+ $Y2=0
cc_280 N_CLK_N_c_281_n N_A_113_67#_c_371_n 2.27703e-19 $X=0.28 $Y=1.12 $X2=0
+ $Y2=0
cc_281 N_CLK_N_M1029_g N_A_113_67#_c_373_n 0.00721658f $X=0.49 $Y=0.545 $X2=0
+ $Y2=0
cc_282 N_CLK_N_c_281_n N_A_113_67#_c_373_n 0.0203015f $X=0.28 $Y=1.12 $X2=0
+ $Y2=0
cc_283 N_CLK_N_c_282_n N_A_113_67#_c_373_n 0.0911511f $X=0.28 $Y=1.12 $X2=0
+ $Y2=0
cc_284 N_CLK_N_c_281_n N_A_113_67#_c_375_n 0.0434121f $X=0.28 $Y=1.12 $X2=0
+ $Y2=0
cc_285 N_CLK_N_c_282_n N_A_113_67#_c_375_n 5.50353e-19 $X=0.28 $Y=1.12 $X2=0
+ $Y2=0
cc_286 N_CLK_N_M1029_g N_A_223_119#_c_1055_n 4.13043e-19 $X=0.49 $Y=0.545 $X2=0
+ $Y2=0
cc_287 N_CLK_N_M1027_g N_VPWR_c_1679_n 0.0140908f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_288 N_CLK_N_c_282_n N_VPWR_c_1679_n 0.0242307f $X=0.28 $Y=1.12 $X2=0 $Y2=0
cc_289 N_CLK_N_M1027_g N_VPWR_c_1687_n 0.00445056f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_290 N_CLK_N_M1027_g N_VPWR_c_1677_n 0.00899805f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_291 N_CLK_N_M1029_g N_VGND_c_1931_n 0.00566738f $X=0.49 $Y=0.545 $X2=0 $Y2=0
cc_292 N_CLK_N_c_281_n N_VGND_c_1931_n 0.00188881f $X=0.28 $Y=1.12 $X2=0 $Y2=0
cc_293 N_CLK_N_c_282_n N_VGND_c_1931_n 0.0207432f $X=0.28 $Y=1.12 $X2=0 $Y2=0
cc_294 N_CLK_N_M1029_g N_VGND_c_1942_n 0.00461273f $X=0.49 $Y=0.545 $X2=0 $Y2=0
cc_295 N_CLK_N_M1029_g N_VGND_c_1947_n 0.00945239f $X=0.49 $Y=0.545 $X2=0 $Y2=0
cc_296 N_D_c_303_n N_A_113_67#_M1009_g 0.0246666f $X=1.975 $Y=1.51 $X2=0 $Y2=0
cc_297 N_D_c_307_n N_A_113_67#_M1009_g 0.00272531f $X=1.915 $Y=1.345 $X2=0 $Y2=0
cc_298 N_D_c_309_n N_A_113_67#_M1032_g 0.00992098f $X=2.225 $Y=2.17 $X2=0 $Y2=0
cc_299 N_D_c_310_n N_A_113_67#_M1032_g 0.0118992f $X=2.225 $Y=2.095 $X2=0 $Y2=0
cc_300 N_D_c_306_n N_A_113_67#_c_357_n 0.0103003f $X=2.36 $Y=1.09 $X2=0 $Y2=0
cc_301 N_D_c_309_n N_A_113_67#_c_378_n 0.0104235f $X=2.225 $Y=2.17 $X2=0 $Y2=0
cc_302 N_D_c_310_n N_A_113_67#_M1036_g 0.0134153f $X=2.225 $Y=2.095 $X2=0 $Y2=0
cc_303 N_D_c_304_n N_A_113_67#_c_375_n 0.0216468f $X=1.975 $Y=2.02 $X2=0 $Y2=0
cc_304 N_D_c_307_n N_A_113_67#_c_375_n 0.00174536f $X=1.915 $Y=1.345 $X2=0 $Y2=0
cc_305 N_D_c_303_n N_A_223_119#_M1023_g 0.00308966f $X=1.975 $Y=1.51 $X2=0 $Y2=0
cc_306 N_D_c_306_n N_A_223_119#_M1023_g 0.0177992f $X=2.36 $Y=1.09 $X2=0 $Y2=0
cc_307 N_D_c_307_n N_A_223_119#_M1023_g 7.87828e-19 $X=1.915 $Y=1.345 $X2=0
+ $Y2=0
cc_308 N_D_c_310_n N_A_223_119#_c_1058_n 0.00109874f $X=2.225 $Y=2.095 $X2=0
+ $Y2=0
cc_309 N_D_c_303_n N_A_223_119#_c_1051_n 0.00197912f $X=1.975 $Y=1.51 $X2=0
+ $Y2=0
cc_310 N_D_c_304_n N_A_223_119#_c_1051_n 0.0177905f $X=1.975 $Y=2.02 $X2=0 $Y2=0
cc_311 N_D_c_305_n N_A_223_119#_c_1051_n 0.008189f $X=2.285 $Y=1.165 $X2=0 $Y2=0
cc_312 N_D_c_310_n N_A_223_119#_c_1051_n 6.56187e-19 $X=2.225 $Y=2.095 $X2=0
+ $Y2=0
cc_313 N_D_c_310_n N_A_223_119#_c_1068_n 6.84014e-19 $X=2.225 $Y=2.095 $X2=0
+ $Y2=0
cc_314 N_D_c_303_n N_A_223_119#_c_1053_n 7.46008e-19 $X=1.975 $Y=1.51 $X2=0
+ $Y2=0
cc_315 N_D_c_304_n N_A_223_119#_c_1053_n 0.0016349f $X=1.975 $Y=2.02 $X2=0 $Y2=0
cc_316 N_D_c_307_n N_A_223_119#_c_1053_n 0.0245882f $X=1.915 $Y=1.345 $X2=0
+ $Y2=0
cc_317 N_D_c_303_n N_A_223_119#_c_1070_n 0.00316172f $X=1.975 $Y=1.51 $X2=0
+ $Y2=0
cc_318 N_D_c_304_n N_A_223_119#_c_1070_n 0.00981452f $X=1.975 $Y=2.02 $X2=0
+ $Y2=0
cc_319 N_D_c_305_n N_A_223_119#_c_1070_n 0.00443558f $X=2.285 $Y=1.165 $X2=0
+ $Y2=0
cc_320 N_D_c_310_n N_A_223_119#_c_1070_n 0.0168112f $X=2.225 $Y=2.095 $X2=0
+ $Y2=0
cc_321 N_D_c_307_n N_A_223_119#_c_1070_n 0.0204418f $X=1.915 $Y=1.345 $X2=0
+ $Y2=0
cc_322 N_D_c_304_n N_A_223_119#_c_1054_n 0.00410242f $X=1.975 $Y=2.02 $X2=0
+ $Y2=0
cc_323 N_D_c_305_n N_A_223_119#_c_1054_n 9.30981e-19 $X=2.285 $Y=1.165 $X2=0
+ $Y2=0
cc_324 N_D_c_307_n N_A_223_119#_c_1054_n 0.00186833f $X=1.915 $Y=1.345 $X2=0
+ $Y2=0
cc_325 N_D_c_309_n N_VPWR_c_1680_n 0.00905793f $X=2.225 $Y=2.17 $X2=0 $Y2=0
cc_326 N_D_c_310_n N_VPWR_c_1680_n 0.00453517f $X=2.225 $Y=2.095 $X2=0 $Y2=0
cc_327 N_D_c_309_n N_VPWR_c_1677_n 8.60012e-19 $X=2.225 $Y=2.17 $X2=0 $Y2=0
cc_328 N_D_c_305_n N_A_460_449#_c_1820_n 0.00230027f $X=2.285 $Y=1.165 $X2=0
+ $Y2=0
cc_329 N_D_c_306_n N_A_460_449#_c_1820_n 0.0134879f $X=2.36 $Y=1.09 $X2=0 $Y2=0
cc_330 N_D_c_304_n N_A_460_449#_c_1821_n 4.53732e-19 $X=1.975 $Y=2.02 $X2=0
+ $Y2=0
cc_331 N_D_c_310_n N_A_460_449#_c_1821_n 0.00168156f $X=2.225 $Y=2.095 $X2=0
+ $Y2=0
cc_332 N_D_c_307_n N_A_460_449#_c_1821_n 0.00312695f $X=1.915 $Y=1.345 $X2=0
+ $Y2=0
cc_333 N_D_c_309_n N_A_460_449#_c_1824_n 0.00569074f $X=2.225 $Y=2.17 $X2=0
+ $Y2=0
cc_334 N_D_c_303_n N_A_460_449#_c_1822_n 2.92269e-19 $X=1.975 $Y=1.51 $X2=0
+ $Y2=0
cc_335 N_D_c_305_n N_A_460_449#_c_1822_n 0.00521064f $X=2.285 $Y=1.165 $X2=0
+ $Y2=0
cc_336 N_D_c_307_n N_A_460_449#_c_1822_n 0.00585641f $X=1.915 $Y=1.345 $X2=0
+ $Y2=0
cc_337 N_D_c_303_n N_VGND_c_1932_n 0.00412711f $X=1.975 $Y=1.51 $X2=0 $Y2=0
cc_338 N_D_c_306_n N_VGND_c_1932_n 0.0111394f $X=2.36 $Y=1.09 $X2=0 $Y2=0
cc_339 N_D_c_307_n N_VGND_c_1932_n 0.0265089f $X=1.915 $Y=1.345 $X2=0 $Y2=0
cc_340 N_D_c_306_n N_VGND_c_1947_n 9.39239e-19 $X=2.36 $Y=1.09 $X2=0 $Y2=0
cc_341 N_A_113_67#_c_365_n N_A_755_398#_M1017_d 0.00385177f $X=6.485 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_342 N_A_113_67#_M1038_g N_A_755_398#_M1031_g 0.0188647f $X=3.435 $Y=0.76
+ $X2=0 $Y2=0
cc_343 N_A_113_67#_c_384_n N_A_755_398#_M1031_g 0.00131637f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_344 N_A_113_67#_c_361_n N_A_755_398#_M1031_g 0.0360344f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_345 N_A_113_67#_c_362_n N_A_755_398#_M1031_g 0.0167805f $X=4.69 $Y=1.14 $X2=0
+ $Y2=0
cc_346 N_A_113_67#_c_364_n N_A_755_398#_M1031_g 0.00435336f $X=4.775 $Y=1.055
+ $X2=0 $Y2=0
cc_347 N_A_113_67#_c_368_n N_A_755_398#_c_608_n 0.00499615f $X=7.36 $Y=1.17
+ $X2=0 $Y2=0
cc_348 N_A_113_67#_c_370_n N_A_755_398#_c_608_n 3.79349e-19 $X=7.445 $Y=1.675
+ $X2=0 $Y2=0
cc_349 N_A_113_67#_c_387_n N_A_755_398#_c_608_n 0.0138212f $X=7.445 $Y=2.895
+ $X2=0 $Y2=0
cc_350 N_A_113_67#_c_374_n N_A_755_398#_c_608_n 0.00687547f $X=7.585 $Y=1.51
+ $X2=0 $Y2=0
cc_351 N_A_113_67#_c_367_n N_A_755_398#_M1005_g 0.00503526f $X=6.57 $Y=1.085
+ $X2=0 $Y2=0
cc_352 N_A_113_67#_c_368_n N_A_755_398#_M1005_g 0.0153878f $X=7.36 $Y=1.17 $X2=0
+ $Y2=0
cc_353 N_A_113_67#_c_370_n N_A_755_398#_M1005_g 0.00491325f $X=7.445 $Y=1.675
+ $X2=0 $Y2=0
cc_354 N_A_113_67#_c_374_n N_A_755_398#_M1005_g 0.0126247f $X=7.585 $Y=1.51
+ $X2=0 $Y2=0
cc_355 N_A_113_67#_c_376_n N_A_755_398#_M1005_g 0.0297824f $X=7.585 $Y=1.345
+ $X2=0 $Y2=0
cc_356 N_A_113_67#_c_369_n N_A_755_398#_c_610_n 0.0103611f $X=6.655 $Y=1.17
+ $X2=0 $Y2=0
cc_357 N_A_113_67#_c_369_n N_A_755_398#_c_612_n 0.0127695f $X=6.655 $Y=1.17
+ $X2=0 $Y2=0
cc_358 N_A_113_67#_c_368_n N_A_755_398#_c_613_n 0.0348891f $X=7.36 $Y=1.17 $X2=0
+ $Y2=0
cc_359 N_A_113_67#_c_370_n N_A_755_398#_c_613_n 0.0182607f $X=7.445 $Y=1.675
+ $X2=0 $Y2=0
cc_360 N_A_113_67#_c_387_n N_A_755_398#_c_613_n 0.00119187f $X=7.445 $Y=2.895
+ $X2=0 $Y2=0
cc_361 N_A_113_67#_c_374_n N_A_755_398#_c_613_n 3.12197e-19 $X=7.585 $Y=1.51
+ $X2=0 $Y2=0
cc_362 N_A_113_67#_c_367_n N_A_755_398#_c_614_n 0.00363818f $X=6.57 $Y=1.085
+ $X2=0 $Y2=0
cc_363 N_A_113_67#_c_369_n N_A_755_398#_c_614_n 0.00128241f $X=6.655 $Y=1.17
+ $X2=0 $Y2=0
cc_364 N_A_113_67#_c_362_n N_SET_B_M1024_g 0.00792239f $X=4.69 $Y=1.14 $X2=0
+ $Y2=0
cc_365 N_A_113_67#_c_364_n N_SET_B_M1024_g 0.0132062f $X=4.775 $Y=1.055 $X2=0
+ $Y2=0
cc_366 N_A_113_67#_c_365_n N_SET_B_M1024_g 0.0144163f $X=6.485 $Y=0.35 $X2=0
+ $Y2=0
cc_367 N_A_113_67#_c_390_n SET_B 0.0070688f $X=8.485 $Y=1.895 $X2=0 $Y2=0
cc_368 N_A_113_67#_c_391_n SET_B 5.98535e-19 $X=8.485 $Y=1.895 $X2=0 $Y2=0
cc_369 N_A_113_67#_c_382_n N_SET_B_c_762_n 0.00427915f $X=8.485 $Y=2.305 $X2=0
+ $Y2=0
cc_370 N_A_113_67#_c_368_n N_SET_B_c_762_n 0.00952633f $X=7.36 $Y=1.17 $X2=0
+ $Y2=0
cc_371 N_A_113_67#_c_369_n N_SET_B_c_762_n 9.98332e-19 $X=6.655 $Y=1.17 $X2=0
+ $Y2=0
cc_372 N_A_113_67#_c_370_n N_SET_B_c_762_n 0.0266024f $X=7.445 $Y=1.675 $X2=0
+ $Y2=0
cc_373 N_A_113_67#_c_387_n N_SET_B_c_762_n 0.0121524f $X=7.445 $Y=2.895 $X2=0
+ $Y2=0
cc_374 N_A_113_67#_c_390_n N_SET_B_c_762_n 0.0193206f $X=8.485 $Y=1.895 $X2=0
+ $Y2=0
cc_375 N_A_113_67#_c_391_n N_SET_B_c_762_n 0.00365763f $X=8.485 $Y=1.895 $X2=0
+ $Y2=0
cc_376 N_A_113_67#_c_374_n N_SET_B_c_762_n 4.36452e-19 $X=7.585 $Y=1.51 $X2=0
+ $Y2=0
cc_377 N_A_113_67#_c_390_n N_SET_B_c_764_n 0.00136161f $X=8.485 $Y=1.895 $X2=0
+ $Y2=0
cc_378 N_A_113_67#_c_391_n N_SET_B_c_764_n 7.27604e-19 $X=8.485 $Y=1.895 $X2=0
+ $Y2=0
cc_379 N_A_113_67#_c_362_n N_SET_B_c_765_n 0.0021982f $X=4.69 $Y=1.14 $X2=0
+ $Y2=0
cc_380 N_A_113_67#_c_365_n N_A_546_449#_M1017_g 0.0101774f $X=6.485 $Y=0.35
+ $X2=0 $Y2=0
cc_381 N_A_113_67#_c_384_n N_A_546_449#_c_901_n 0.0361961f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_382 N_A_113_67#_c_361_n N_A_546_449#_c_901_n 0.0103658f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_383 N_A_113_67#_c_363_n N_A_546_449#_c_901_n 0.0129661f $X=3.62 $Y=1.14 $X2=0
+ $Y2=0
cc_384 N_A_113_67#_c_384_n N_A_546_449#_c_911_n 0.00652275f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_385 N_A_113_67#_c_361_n N_A_546_449#_c_911_n 0.0026796f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_386 N_A_113_67#_c_384_n N_A_546_449#_c_902_n 0.0120512f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_387 N_A_113_67#_c_361_n N_A_546_449#_c_902_n 0.00114065f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_388 N_A_113_67#_c_362_n N_A_546_449#_c_903_n 0.0530348f $X=4.69 $Y=1.14 $X2=0
+ $Y2=0
cc_389 N_A_113_67#_c_384_n N_A_546_449#_c_904_n 0.0132341f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_390 N_A_113_67#_c_361_n N_A_546_449#_c_904_n 0.0012848f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_391 N_A_113_67#_c_362_n N_A_546_449#_c_904_n 0.0134534f $X=4.69 $Y=1.14 $X2=0
+ $Y2=0
cc_392 N_A_113_67#_c_357_n N_A_546_449#_c_908_n 0.0067834f $X=3.36 $Y=0.18 $X2=0
+ $Y2=0
cc_393 N_A_113_67#_M1038_g N_A_546_449#_c_908_n 0.0103658f $X=3.435 $Y=0.76
+ $X2=0 $Y2=0
cc_394 N_A_113_67#_M1036_g N_A_546_449#_c_919_n 0.00295918f $X=2.655 $Y=2.455
+ $X2=0 $Y2=0
cc_395 N_A_113_67#_c_361_n N_A_546_449#_c_919_n 2.29269e-19 $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_396 N_A_113_67#_c_357_n N_A_223_119#_M1023_g 0.0103003f $X=3.36 $Y=0.18 $X2=0
+ $Y2=0
cc_397 N_A_113_67#_M1038_g N_A_223_119#_M1023_g 0.010274f $X=3.435 $Y=0.76 $X2=0
+ $Y2=0
cc_398 N_A_113_67#_c_384_n N_A_223_119#_c_1057_n 5.05812e-19 $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_399 N_A_113_67#_c_361_n N_A_223_119#_c_1057_n 0.00923753f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_400 N_A_113_67#_M1036_g N_A_223_119#_c_1058_n 0.00265089f $X=2.655 $Y=2.455
+ $X2=0 $Y2=0
cc_401 N_A_113_67#_M1036_g N_A_223_119#_M1033_g 0.00708051f $X=2.655 $Y=2.455
+ $X2=0 $Y2=0
cc_402 N_A_113_67#_c_381_n N_A_223_119#_c_1060_n 0.00922235f $X=8.17 $Y=2.455
+ $X2=0 $Y2=0
cc_403 N_A_113_67#_c_389_n N_A_223_119#_c_1060_n 0.00135484f $X=7.53 $Y=2.98
+ $X2=0 $Y2=0
cc_404 N_A_113_67#_c_378_n N_A_223_119#_c_1061_n 0.00708051f $X=2.58 $Y=3.08
+ $X2=0 $Y2=0
cc_405 N_A_113_67#_c_382_n N_A_223_119#_M1021_g 0.00922235f $X=8.485 $Y=2.305
+ $X2=0 $Y2=0
cc_406 N_A_113_67#_c_387_n N_A_223_119#_M1021_g 0.0178895f $X=7.445 $Y=2.895
+ $X2=0 $Y2=0
cc_407 N_A_113_67#_c_388_n N_A_223_119#_M1021_g 0.0113053f $X=8.32 $Y=2.98 $X2=0
+ $Y2=0
cc_408 N_A_113_67#_c_389_n N_A_223_119#_M1021_g 0.0035501f $X=7.53 $Y=2.98 $X2=0
+ $Y2=0
cc_409 N_A_113_67#_c_391_n N_A_223_119#_M1021_g 0.00238264f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_410 N_A_113_67#_c_382_n N_A_223_119#_c_1063_n 0.00102066f $X=8.485 $Y=2.305
+ $X2=0 $Y2=0
cc_411 N_A_113_67#_c_370_n N_A_223_119#_c_1064_n 0.00233248f $X=7.445 $Y=1.675
+ $X2=0 $Y2=0
cc_412 N_A_113_67#_c_387_n N_A_223_119#_c_1064_n 0.00511403f $X=7.445 $Y=2.895
+ $X2=0 $Y2=0
cc_413 N_A_113_67#_c_374_n N_A_223_119#_c_1064_n 0.013269f $X=7.585 $Y=1.51
+ $X2=0 $Y2=0
cc_414 N_A_113_67#_c_387_n N_A_223_119#_c_1047_n 0.00127287f $X=7.445 $Y=2.895
+ $X2=0 $Y2=0
cc_415 N_A_113_67#_c_390_n N_A_223_119#_c_1047_n 0.0011518f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_416 N_A_113_67#_c_391_n N_A_223_119#_c_1047_n 0.0202912f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_417 N_A_113_67#_c_390_n N_A_223_119#_c_1048_n 8.68712e-19 $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_418 N_A_113_67#_c_391_n N_A_223_119#_c_1048_n 0.00713933f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_419 N_A_113_67#_c_370_n N_A_223_119#_c_1049_n 4.41579e-19 $X=7.445 $Y=1.675
+ $X2=0 $Y2=0
cc_420 N_A_113_67#_c_374_n N_A_223_119#_c_1049_n 0.0213403f $X=7.585 $Y=1.51
+ $X2=0 $Y2=0
cc_421 N_A_113_67#_c_376_n N_A_223_119#_c_1049_n 0.0017406f $X=7.585 $Y=1.345
+ $X2=0 $Y2=0
cc_422 N_A_113_67#_c_376_n N_A_223_119#_c_1050_n 0.00720201f $X=7.585 $Y=1.345
+ $X2=0 $Y2=0
cc_423 N_A_113_67#_M1036_g N_A_223_119#_c_1051_n 0.00767437f $X=2.655 $Y=2.455
+ $X2=0 $Y2=0
cc_424 N_A_113_67#_c_361_n N_A_223_119#_c_1052_n 0.0149941f $X=3.525 $Y=1.245
+ $X2=0 $Y2=0
cc_425 N_A_113_67#_M1032_g N_A_223_119#_c_1068_n 0.00958839f $X=1.585 $Y=2.565
+ $X2=0 $Y2=0
cc_426 N_A_113_67#_c_383_n N_A_223_119#_c_1068_n 0.0206743f $X=0.79 $Y=2.55
+ $X2=0 $Y2=0
cc_427 N_A_113_67#_c_375_n N_A_223_119#_c_1068_n 0.0160241f $X=1.465 $Y=1.547
+ $X2=0 $Y2=0
cc_428 N_A_113_67#_M1032_g N_A_223_119#_c_1069_n 0.00896663f $X=1.585 $Y=2.565
+ $X2=0 $Y2=0
cc_429 N_A_113_67#_c_383_n N_A_223_119#_c_1069_n 0.0442049f $X=0.79 $Y=2.55
+ $X2=0 $Y2=0
cc_430 N_A_113_67#_M1009_g N_A_223_119#_c_1053_n 0.00787087f $X=1.465 $Y=0.805
+ $X2=0 $Y2=0
cc_431 N_A_113_67#_c_383_n N_A_223_119#_c_1053_n 4.19374e-19 $X=0.79 $Y=2.55
+ $X2=0 $Y2=0
cc_432 N_A_113_67#_c_372_n N_A_223_119#_c_1053_n 0.0467084f $X=0.945 $Y=1.36
+ $X2=0 $Y2=0
cc_433 N_A_113_67#_c_373_n N_A_223_119#_c_1053_n 0.00802392f $X=0.845 $Y=1.195
+ $X2=0 $Y2=0
cc_434 N_A_113_67#_c_375_n N_A_223_119#_c_1053_n 0.0318862f $X=1.465 $Y=1.547
+ $X2=0 $Y2=0
cc_435 N_A_113_67#_M1032_g N_A_223_119#_c_1070_n 0.00860984f $X=1.585 $Y=2.565
+ $X2=0 $Y2=0
cc_436 N_A_113_67#_c_375_n N_A_223_119#_c_1070_n 0.00350336f $X=1.465 $Y=1.547
+ $X2=0 $Y2=0
cc_437 N_A_113_67#_M1009_g N_A_223_119#_c_1055_n 0.00680518f $X=1.465 $Y=0.805
+ $X2=0 $Y2=0
cc_438 N_A_113_67#_c_371_n N_A_223_119#_c_1055_n 0.0306756f $X=0.705 $Y=0.545
+ $X2=0 $Y2=0
cc_439 N_A_113_67#_c_375_n N_A_223_119#_c_1055_n 0.00718807f $X=1.465 $Y=1.547
+ $X2=0 $Y2=0
cc_440 N_A_113_67#_c_381_n N_A_1741_137#_M1000_g 0.00717512f $X=8.17 $Y=2.455
+ $X2=0 $Y2=0
cc_441 N_A_113_67#_c_382_n N_A_1741_137#_M1000_g 0.00321678f $X=8.485 $Y=2.305
+ $X2=0 $Y2=0
cc_442 N_A_113_67#_c_388_n N_A_1741_137#_M1000_g 0.00223055f $X=8.32 $Y=2.98
+ $X2=0 $Y2=0
cc_443 N_A_113_67#_c_390_n N_A_1741_137#_M1000_g 0.00690445f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_444 N_A_113_67#_c_390_n N_A_1741_137#_c_1228_n 0.0193387f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_445 N_A_113_67#_c_391_n N_A_1741_137#_c_1228_n 0.00120179f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_446 N_A_113_67#_c_382_n N_A_1741_137#_c_1229_n 0.0213378f $X=8.485 $Y=2.305
+ $X2=0 $Y2=0
cc_447 N_A_113_67#_c_390_n N_A_1741_137#_c_1229_n 3.92283e-19 $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_448 N_A_113_67#_c_390_n N_A_1741_137#_c_1222_n 0.00158688f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_449 N_A_113_67#_c_391_n N_A_1741_137#_c_1222_n 0.0213378f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_450 N_A_113_67#_c_388_n N_A_1531_428#_M1021_d 0.00392154f $X=8.32 $Y=2.98
+ $X2=0 $Y2=0
cc_451 N_A_113_67#_c_381_n N_A_1531_428#_c_1389_n 0.00659397f $X=8.17 $Y=2.455
+ $X2=0 $Y2=0
cc_452 N_A_113_67#_c_382_n N_A_1531_428#_c_1389_n 0.00468001f $X=8.485 $Y=2.305
+ $X2=0 $Y2=0
cc_453 N_A_113_67#_c_370_n N_A_1531_428#_c_1389_n 9.03112e-19 $X=7.445 $Y=1.675
+ $X2=0 $Y2=0
cc_454 N_A_113_67#_c_387_n N_A_1531_428#_c_1389_n 0.0200399f $X=7.445 $Y=2.895
+ $X2=0 $Y2=0
cc_455 N_A_113_67#_c_388_n N_A_1531_428#_c_1389_n 0.0237862f $X=8.32 $Y=2.98
+ $X2=0 $Y2=0
cc_456 N_A_113_67#_c_376_n N_A_1531_428#_c_1381_n 0.0147003f $X=7.585 $Y=1.345
+ $X2=0 $Y2=0
cc_457 N_A_113_67#_c_390_n N_A_1531_428#_c_1382_n 0.00624077f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_458 N_A_113_67#_c_391_n N_A_1531_428#_c_1382_n 0.0018745f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_459 N_A_113_67#_c_370_n N_A_1531_428#_c_1384_n 0.0244806f $X=7.445 $Y=1.675
+ $X2=0 $Y2=0
cc_460 N_A_113_67#_c_387_n N_A_1531_428#_c_1384_n 0.0164042f $X=7.445 $Y=2.895
+ $X2=0 $Y2=0
cc_461 N_A_113_67#_c_390_n N_A_1531_428#_c_1384_n 0.0606006f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_462 N_A_113_67#_c_391_n N_A_1531_428#_c_1384_n 0.00365056f $X=8.485 $Y=1.895
+ $X2=0 $Y2=0
cc_463 N_A_113_67#_c_374_n N_A_1531_428#_c_1384_n 9.39256e-19 $X=7.585 $Y=1.51
+ $X2=0 $Y2=0
cc_464 N_A_113_67#_c_370_n N_A_1531_428#_c_1385_n 0.00605747f $X=7.445 $Y=1.675
+ $X2=0 $Y2=0
cc_465 N_A_113_67#_c_376_n N_A_1531_428#_c_1385_n 0.00199747f $X=7.585 $Y=1.345
+ $X2=0 $Y2=0
cc_466 N_A_113_67#_c_365_n N_A_1186_21#_M1012_g 0.0106317f $X=6.485 $Y=0.35
+ $X2=0 $Y2=0
cc_467 N_A_113_67#_c_367_n N_A_1186_21#_M1012_g 0.00439847f $X=6.57 $Y=1.085
+ $X2=0 $Y2=0
cc_468 N_A_113_67#_c_365_n N_A_1186_21#_c_1477_n 0.0115412f $X=6.485 $Y=0.35
+ $X2=0 $Y2=0
cc_469 N_A_113_67#_c_376_n N_A_1186_21#_c_1477_n 0.0104164f $X=7.585 $Y=1.345
+ $X2=0 $Y2=0
cc_470 N_A_113_67#_c_365_n N_A_1186_21#_c_1479_n 0.00457315f $X=6.485 $Y=0.35
+ $X2=0 $Y2=0
cc_471 N_A_113_67#_c_367_n N_A_1186_21#_c_1479_n 0.00269204f $X=6.57 $Y=1.085
+ $X2=0 $Y2=0
cc_472 N_A_113_67#_c_369_n N_A_1186_21#_c_1479_n 0.00454105f $X=6.655 $Y=1.17
+ $X2=0 $Y2=0
cc_473 N_A_113_67#_c_369_n N_A_1186_21#_M1020_g 0.00246138f $X=6.655 $Y=1.17
+ $X2=0 $Y2=0
cc_474 N_A_113_67#_c_383_n N_VPWR_c_1679_n 0.0258905f $X=0.79 $Y=2.55 $X2=0
+ $Y2=0
cc_475 N_A_113_67#_M1032_g N_VPWR_c_1680_n 0.0102682f $X=1.585 $Y=2.565 $X2=0
+ $Y2=0
cc_476 N_A_113_67#_c_378_n N_VPWR_c_1680_n 0.0284081f $X=2.58 $Y=3.08 $X2=0
+ $Y2=0
cc_477 N_A_113_67#_M1036_g N_VPWR_c_1680_n 0.00549858f $X=2.655 $Y=2.455 $X2=0
+ $Y2=0
cc_478 N_A_113_67#_c_387_n N_VPWR_c_1682_n 0.0482063f $X=7.445 $Y=2.895 $X2=0
+ $Y2=0
cc_479 N_A_113_67#_c_389_n N_VPWR_c_1682_n 0.0098469f $X=7.53 $Y=2.98 $X2=0
+ $Y2=0
cc_480 N_A_113_67#_c_388_n N_VPWR_c_1683_n 0.00588632f $X=8.32 $Y=2.98 $X2=0
+ $Y2=0
cc_481 N_A_113_67#_c_390_n N_VPWR_c_1683_n 0.00969659f $X=8.485 $Y=1.895 $X2=0
+ $Y2=0
cc_482 N_A_113_67#_c_379_n N_VPWR_c_1687_n 0.00675559f $X=1.66 $Y=3.08 $X2=0
+ $Y2=0
cc_483 N_A_113_67#_c_383_n N_VPWR_c_1687_n 0.0221152f $X=0.79 $Y=2.55 $X2=0
+ $Y2=0
cc_484 N_A_113_67#_c_378_n N_VPWR_c_1689_n 0.0189178f $X=2.58 $Y=3.08 $X2=0
+ $Y2=0
cc_485 N_A_113_67#_c_381_n N_VPWR_c_1694_n 0.00290313f $X=8.17 $Y=2.455 $X2=0
+ $Y2=0
cc_486 N_A_113_67#_c_388_n N_VPWR_c_1694_n 0.0669521f $X=8.32 $Y=2.98 $X2=0
+ $Y2=0
cc_487 N_A_113_67#_c_389_n N_VPWR_c_1694_n 0.0113436f $X=7.53 $Y=2.98 $X2=0
+ $Y2=0
cc_488 N_A_113_67#_c_378_n N_VPWR_c_1677_n 0.0272517f $X=2.58 $Y=3.08 $X2=0
+ $Y2=0
cc_489 N_A_113_67#_c_379_n N_VPWR_c_1677_n 0.00953141f $X=1.66 $Y=3.08 $X2=0
+ $Y2=0
cc_490 N_A_113_67#_c_381_n N_VPWR_c_1677_n 0.0040605f $X=8.17 $Y=2.455 $X2=0
+ $Y2=0
cc_491 N_A_113_67#_c_382_n N_VPWR_c_1677_n 9.0413e-19 $X=8.485 $Y=2.305 $X2=0
+ $Y2=0
cc_492 N_A_113_67#_c_383_n N_VPWR_c_1677_n 0.0126914f $X=0.79 $Y=2.55 $X2=0
+ $Y2=0
cc_493 N_A_113_67#_c_388_n N_VPWR_c_1677_n 0.0396725f $X=8.32 $Y=2.98 $X2=0
+ $Y2=0
cc_494 N_A_113_67#_c_389_n N_VPWR_c_1677_n 0.00585025f $X=7.53 $Y=2.98 $X2=0
+ $Y2=0
cc_495 N_A_113_67#_c_357_n N_A_460_449#_c_1820_n 0.00582439f $X=3.36 $Y=0.18
+ $X2=0 $Y2=0
cc_496 N_A_113_67#_M1036_g N_A_460_449#_c_1821_n 0.00371878f $X=2.655 $Y=2.455
+ $X2=0 $Y2=0
cc_497 N_A_113_67#_c_378_n N_A_460_449#_c_1824_n 0.00389513f $X=2.58 $Y=3.08
+ $X2=0 $Y2=0
cc_498 N_A_113_67#_M1036_g N_A_460_449#_c_1824_n 0.0151046f $X=2.655 $Y=2.455
+ $X2=0 $Y2=0
cc_499 N_A_113_67#_c_387_n A_1436_379# 0.0107406f $X=7.445 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_500 N_A_113_67#_c_389_n A_1436_379# 0.00123794f $X=7.53 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_501 N_A_113_67#_c_388_n A_1649_512# 0.00246644f $X=8.32 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_502 N_A_113_67#_c_390_n A_1649_512# 0.0117371f $X=8.485 $Y=1.895 $X2=-0.19
+ $Y2=-0.245
cc_503 N_A_113_67#_c_364_n N_VGND_M1031_d 0.00971632f $X=4.775 $Y=1.055 $X2=0
+ $Y2=0
cc_504 N_A_113_67#_c_366_n N_VGND_M1031_d 0.00144038f $X=4.86 $Y=0.35 $X2=0
+ $Y2=0
cc_505 N_A_113_67#_c_368_n N_VGND_M1005_s 0.00501179f $X=7.36 $Y=1.17 $X2=0
+ $Y2=0
cc_506 N_A_113_67#_c_371_n N_VGND_c_1931_n 0.0179429f $X=0.705 $Y=0.545 $X2=0
+ $Y2=0
cc_507 N_A_113_67#_M1009_g N_VGND_c_1932_n 0.0216434f $X=1.465 $Y=0.805 $X2=0
+ $Y2=0
cc_508 N_A_113_67#_c_357_n N_VGND_c_1932_n 0.0248025f $X=3.36 $Y=0.18 $X2=0
+ $Y2=0
cc_509 N_A_113_67#_c_357_n N_VGND_c_1933_n 0.00663125f $X=3.36 $Y=0.18 $X2=0
+ $Y2=0
cc_510 N_A_113_67#_c_362_n N_VGND_c_1933_n 0.0260135f $X=4.69 $Y=1.14 $X2=0
+ $Y2=0
cc_511 N_A_113_67#_c_364_n N_VGND_c_1933_n 0.0321918f $X=4.775 $Y=1.055 $X2=0
+ $Y2=0
cc_512 N_A_113_67#_c_366_n N_VGND_c_1933_n 0.0140894f $X=4.86 $Y=0.35 $X2=0
+ $Y2=0
cc_513 N_A_113_67#_c_365_n N_VGND_c_1934_n 0.0141601f $X=6.485 $Y=0.35 $X2=0
+ $Y2=0
cc_514 N_A_113_67#_c_367_n N_VGND_c_1934_n 0.0345265f $X=6.57 $Y=1.085 $X2=0
+ $Y2=0
cc_515 N_A_113_67#_c_368_n N_VGND_c_1934_n 0.0147238f $X=7.36 $Y=1.17 $X2=0
+ $Y2=0
cc_516 N_A_113_67#_c_376_n N_VGND_c_1934_n 0.00207662f $X=7.585 $Y=1.345 $X2=0
+ $Y2=0
cc_517 N_A_113_67#_c_357_n N_VGND_c_1938_n 0.0492316f $X=3.36 $Y=0.18 $X2=0
+ $Y2=0
cc_518 N_A_113_67#_c_358_n N_VGND_c_1942_n 0.00768994f $X=1.54 $Y=0.18 $X2=0
+ $Y2=0
cc_519 N_A_113_67#_c_371_n N_VGND_c_1942_n 0.0168228f $X=0.705 $Y=0.545 $X2=0
+ $Y2=0
cc_520 N_A_113_67#_c_365_n N_VGND_c_1943_n 0.108638f $X=6.485 $Y=0.35 $X2=0
+ $Y2=0
cc_521 N_A_113_67#_c_366_n N_VGND_c_1943_n 0.0114622f $X=4.86 $Y=0.35 $X2=0
+ $Y2=0
cc_522 N_A_113_67#_c_357_n N_VGND_c_1947_n 0.0689974f $X=3.36 $Y=0.18 $X2=0
+ $Y2=0
cc_523 N_A_113_67#_c_358_n N_VGND_c_1947_n 0.0106678f $X=1.54 $Y=0.18 $X2=0
+ $Y2=0
cc_524 N_A_113_67#_c_365_n N_VGND_c_1947_n 0.0629179f $X=6.485 $Y=0.35 $X2=0
+ $Y2=0
cc_525 N_A_113_67#_c_366_n N_VGND_c_1947_n 0.00657784f $X=4.86 $Y=0.35 $X2=0
+ $Y2=0
cc_526 N_A_113_67#_c_371_n N_VGND_c_1947_n 0.0122116f $X=0.705 $Y=0.545 $X2=0
+ $Y2=0
cc_527 N_A_113_67#_c_376_n N_VGND_c_1947_n 9.39239e-19 $X=7.585 $Y=1.345 $X2=0
+ $Y2=0
cc_528 N_A_113_67#_c_365_n N_A_1013_66#_M1024_d 0.00186629f $X=6.485 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_529 N_A_113_67#_c_365_n N_A_1013_66#_M1012_d 0.00330037f $X=6.485 $Y=0.35
+ $X2=0 $Y2=0
cc_530 N_A_113_67#_c_364_n N_A_1013_66#_c_2059_n 0.0148023f $X=4.775 $Y=1.055
+ $X2=0 $Y2=0
cc_531 N_A_113_67#_c_365_n N_A_1013_66#_c_2059_n 0.0522087f $X=6.485 $Y=0.35
+ $X2=0 $Y2=0
cc_532 N_A_113_67#_c_365_n N_A_1013_66#_c_2064_n 0.0114888f $X=6.485 $Y=0.35
+ $X2=0 $Y2=0
cc_533 N_A_113_67#_c_367_n N_A_1013_66#_c_2064_n 0.0234193f $X=6.57 $Y=1.085
+ $X2=0 $Y2=0
cc_534 N_A_113_67#_c_368_n A_1442_119# 0.00351031f $X=7.36 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_535 N_A_113_67#_c_370_n A_1442_119# 0.00744656f $X=7.445 $Y=1.675 $X2=-0.19
+ $Y2=-0.245
cc_536 N_A_755_398#_c_619_n N_SET_B_M1037_g 0.00380294f $X=4.245 $Y=1.92 $X2=0
+ $Y2=0
cc_537 N_A_755_398#_c_649_p N_SET_B_M1037_g 0.0139161f $X=5.685 $Y=2.395 $X2=0
+ $Y2=0
cc_538 N_A_755_398#_c_650_p N_SET_B_M1037_g 5.52917e-19 $X=5.85 $Y=2.085 $X2=0
+ $Y2=0
cc_539 N_A_755_398#_c_651_p N_SET_B_M1037_g 0.0046913f $X=5.85 $Y=2.31 $X2=0
+ $Y2=0
cc_540 N_A_755_398#_c_623_n N_SET_B_M1037_g 0.00728481f $X=5.85 $Y=2.395 $X2=0
+ $Y2=0
cc_541 N_A_755_398#_c_624_n N_SET_B_M1037_g 0.00541027f $X=4.005 $Y=1.947 $X2=0
+ $Y2=0
cc_542 N_A_755_398#_c_608_n N_SET_B_c_762_n 0.00390004f $X=7.105 $Y=1.73 $X2=0
+ $Y2=0
cc_543 N_A_755_398#_M1004_g N_SET_B_c_762_n 0.00538523f $X=7.105 $Y=2.315 $X2=0
+ $Y2=0
cc_544 N_A_755_398#_c_649_p N_SET_B_c_762_n 0.00392284f $X=5.685 $Y=2.395 $X2=0
+ $Y2=0
cc_545 N_A_755_398#_c_650_p N_SET_B_c_762_n 0.00777916f $X=5.85 $Y=2.085 $X2=0
+ $Y2=0
cc_546 N_A_755_398#_c_610_n N_SET_B_c_762_n 0.00459857f $X=6.135 $Y=1.21 $X2=0
+ $Y2=0
cc_547 N_A_755_398#_c_659_p N_SET_B_c_762_n 0.00922921f $X=6.375 $Y=2 $X2=0
+ $Y2=0
cc_548 N_A_755_398#_c_611_n N_SET_B_c_762_n 8.66912e-19 $X=6.22 $Y=1.435 $X2=0
+ $Y2=0
cc_549 N_A_755_398#_c_620_n N_SET_B_c_762_n 0.0108555f $X=6.46 $Y=1.915 $X2=0
+ $Y2=0
cc_550 N_A_755_398#_c_612_n N_SET_B_c_762_n 0.01559f $X=6.545 $Y=1.565 $X2=0
+ $Y2=0
cc_551 N_A_755_398#_c_613_n N_SET_B_c_762_n 0.0230842f $X=7.015 $Y=1.565 $X2=0
+ $Y2=0
cc_552 N_A_755_398#_c_614_n N_SET_B_c_762_n 0.00200222f $X=5.715 $Y=1.13 $X2=0
+ $Y2=0
cc_553 N_A_755_398#_c_611_n N_A_546_449#_M1017_g 0.00230702f $X=6.22 $Y=1.435
+ $X2=0 $Y2=0
cc_554 N_A_755_398#_c_614_n N_A_546_449#_M1017_g 0.0104431f $X=5.715 $Y=1.13
+ $X2=0 $Y2=0
cc_555 N_A_755_398#_c_649_p N_A_546_449#_M1003_g 2.90452e-19 $X=5.685 $Y=2.395
+ $X2=0 $Y2=0
cc_556 N_A_755_398#_c_650_p N_A_546_449#_M1003_g 9.18867e-19 $X=5.85 $Y=2.085
+ $X2=0 $Y2=0
cc_557 N_A_755_398#_c_651_p N_A_546_449#_M1003_g 0.00463691f $X=5.85 $Y=2.31
+ $X2=0 $Y2=0
cc_558 N_A_755_398#_c_659_p N_A_546_449#_M1003_g 0.0118106f $X=6.375 $Y=2 $X2=0
+ $Y2=0
cc_559 N_A_755_398#_c_623_n N_A_546_449#_M1003_g 0.0102814f $X=5.85 $Y=2.395
+ $X2=0 $Y2=0
cc_560 N_A_755_398#_M1031_g N_A_546_449#_c_901_n 0.00102235f $X=4.005 $Y=0.76
+ $X2=0 $Y2=0
cc_561 N_A_755_398#_c_624_n N_A_546_449#_c_901_n 6.43471e-19 $X=4.005 $Y=1.947
+ $X2=0 $Y2=0
cc_562 N_A_755_398#_c_615_n N_A_546_449#_c_911_n 0.0109704f $X=3.85 $Y=2.14
+ $X2=0 $Y2=0
cc_563 N_A_755_398#_c_619_n N_A_546_449#_c_911_n 0.00387559f $X=4.245 $Y=1.92
+ $X2=0 $Y2=0
cc_564 N_A_755_398#_c_615_n N_A_546_449#_c_902_n 0.00324677f $X=3.85 $Y=2.14
+ $X2=0 $Y2=0
cc_565 N_A_755_398#_M1031_g N_A_546_449#_c_902_n 0.00479542f $X=4.005 $Y=0.76
+ $X2=0 $Y2=0
cc_566 N_A_755_398#_c_619_n N_A_546_449#_c_902_n 0.0313677f $X=4.245 $Y=1.92
+ $X2=0 $Y2=0
cc_567 N_A_755_398#_c_624_n N_A_546_449#_c_902_n 0.0184119f $X=4.005 $Y=1.947
+ $X2=0 $Y2=0
cc_568 N_A_755_398#_M1031_g N_A_546_449#_c_903_n 0.0117891f $X=4.005 $Y=0.76
+ $X2=0 $Y2=0
cc_569 N_A_755_398#_c_619_n N_A_546_449#_c_903_n 0.0147674f $X=4.245 $Y=1.92
+ $X2=0 $Y2=0
cc_570 N_A_755_398#_c_624_n N_A_546_449#_c_903_n 0.00652965f $X=4.005 $Y=1.947
+ $X2=0 $Y2=0
cc_571 N_A_755_398#_M1031_g N_A_546_449#_c_904_n 0.00224778f $X=4.005 $Y=0.76
+ $X2=0 $Y2=0
cc_572 N_A_755_398#_M1031_g N_A_546_449#_c_905_n 0.00294159f $X=4.005 $Y=0.76
+ $X2=0 $Y2=0
cc_573 N_A_755_398#_c_619_n N_A_546_449#_c_905_n 0.0140935f $X=4.245 $Y=1.92
+ $X2=0 $Y2=0
cc_574 N_A_755_398#_c_624_n N_A_546_449#_c_905_n 0.00236092f $X=4.005 $Y=1.947
+ $X2=0 $Y2=0
cc_575 N_A_755_398#_M1037_d N_A_546_449#_c_958_n 0.00871375f $X=5.14 $Y=1.895
+ $X2=0 $Y2=0
cc_576 N_A_755_398#_c_649_p N_A_546_449#_c_958_n 0.047819f $X=5.685 $Y=2.395
+ $X2=0 $Y2=0
cc_577 N_A_755_398#_c_650_p N_A_546_449#_c_958_n 0.0107957f $X=5.85 $Y=2.085
+ $X2=0 $Y2=0
cc_578 N_A_755_398#_c_651_p N_A_546_449#_c_958_n 0.00363338f $X=5.85 $Y=2.31
+ $X2=0 $Y2=0
cc_579 N_A_755_398#_c_619_n N_A_546_449#_c_914_n 0.0132567f $X=4.245 $Y=1.92
+ $X2=0 $Y2=0
cc_580 N_A_755_398#_c_649_p N_A_546_449#_c_914_n 0.0133439f $X=5.685 $Y=2.395
+ $X2=0 $Y2=0
cc_581 N_A_755_398#_c_624_n N_A_546_449#_c_914_n 0.00221666f $X=4.005 $Y=1.947
+ $X2=0 $Y2=0
cc_582 N_A_755_398#_M1037_d N_A_546_449#_c_915_n 0.00214809f $X=5.14 $Y=1.895
+ $X2=0 $Y2=0
cc_583 N_A_755_398#_c_650_p N_A_546_449#_c_915_n 0.00347295f $X=5.85 $Y=2.085
+ $X2=0 $Y2=0
cc_584 N_A_755_398#_c_649_p N_A_546_449#_c_917_n 0.00299167f $X=5.685 $Y=2.395
+ $X2=0 $Y2=0
cc_585 N_A_755_398#_c_650_p N_A_546_449#_c_917_n 0.0168101f $X=5.85 $Y=2.085
+ $X2=0 $Y2=0
cc_586 N_A_755_398#_c_610_n N_A_546_449#_c_917_n 0.00488729f $X=6.135 $Y=1.21
+ $X2=0 $Y2=0
cc_587 N_A_755_398#_c_620_n N_A_546_449#_c_917_n 9.58716e-19 $X=6.46 $Y=1.915
+ $X2=0 $Y2=0
cc_588 N_A_755_398#_c_612_n N_A_546_449#_c_917_n 0.0157219f $X=6.545 $Y=1.565
+ $X2=0 $Y2=0
cc_589 N_A_755_398#_c_614_n N_A_546_449#_c_917_n 0.0225561f $X=5.715 $Y=1.13
+ $X2=0 $Y2=0
cc_590 N_A_755_398#_c_649_p N_A_546_449#_c_907_n 6.25207e-19 $X=5.685 $Y=2.395
+ $X2=0 $Y2=0
cc_591 N_A_755_398#_c_650_p N_A_546_449#_c_907_n 0.00523169f $X=5.85 $Y=2.085
+ $X2=0 $Y2=0
cc_592 N_A_755_398#_c_610_n N_A_546_449#_c_907_n 0.00342752f $X=6.135 $Y=1.21
+ $X2=0 $Y2=0
cc_593 N_A_755_398#_c_611_n N_A_546_449#_c_907_n 0.00153031f $X=6.22 $Y=1.435
+ $X2=0 $Y2=0
cc_594 N_A_755_398#_c_620_n N_A_546_449#_c_907_n 0.00325965f $X=6.46 $Y=1.915
+ $X2=0 $Y2=0
cc_595 N_A_755_398#_c_612_n N_A_546_449#_c_907_n 0.00743425f $X=6.545 $Y=1.565
+ $X2=0 $Y2=0
cc_596 N_A_755_398#_c_614_n N_A_546_449#_c_907_n 0.00782124f $X=5.715 $Y=1.13
+ $X2=0 $Y2=0
cc_597 N_A_755_398#_c_615_n N_A_546_449#_c_919_n 0.00143523f $X=3.85 $Y=2.14
+ $X2=0 $Y2=0
cc_598 N_A_755_398#_c_624_n N_A_223_119#_c_1056_n 3.96836e-19 $X=4.005 $Y=1.947
+ $X2=0 $Y2=0
cc_599 N_A_755_398#_c_624_n N_A_223_119#_c_1057_n 0.0212381f $X=4.005 $Y=1.947
+ $X2=0 $Y2=0
cc_600 N_A_755_398#_c_615_n N_A_223_119#_M1033_g 0.0212381f $X=3.85 $Y=2.14
+ $X2=0 $Y2=0
cc_601 N_A_755_398#_c_615_n N_A_223_119#_c_1060_n 0.00729606f $X=3.85 $Y=2.14
+ $X2=0 $Y2=0
cc_602 N_A_755_398#_M1004_g N_A_223_119#_c_1060_n 0.0103107f $X=7.105 $Y=2.315
+ $X2=0 $Y2=0
cc_603 N_A_755_398#_c_649_p N_A_223_119#_c_1060_n 0.0185756f $X=5.685 $Y=2.395
+ $X2=0 $Y2=0
cc_604 N_A_755_398#_c_716_p N_A_223_119#_c_1060_n 0.0051239f $X=4.345 $Y=2.395
+ $X2=0 $Y2=0
cc_605 N_A_755_398#_c_623_n N_A_223_119#_c_1060_n 0.00624358f $X=5.85 $Y=2.395
+ $X2=0 $Y2=0
cc_606 N_A_755_398#_M1004_g N_A_223_119#_c_1064_n 0.0315699f $X=7.105 $Y=2.315
+ $X2=0 $Y2=0
cc_607 N_A_755_398#_c_614_n N_A_1186_21#_M1012_g 0.0028641f $X=5.715 $Y=1.13
+ $X2=0 $Y2=0
cc_608 N_A_755_398#_M1005_g N_A_1186_21#_c_1477_n 0.0103107f $X=7.135 $Y=0.915
+ $X2=0 $Y2=0
cc_609 N_A_755_398#_M1005_g N_A_1186_21#_c_1479_n 0.00773473f $X=7.135 $Y=0.915
+ $X2=0 $Y2=0
cc_610 N_A_755_398#_c_610_n N_A_1186_21#_c_1479_n 0.00775278f $X=6.135 $Y=1.21
+ $X2=0 $Y2=0
cc_611 N_A_755_398#_c_612_n N_A_1186_21#_c_1479_n 0.00317609f $X=6.545 $Y=1.565
+ $X2=0 $Y2=0
cc_612 N_A_755_398#_c_610_n N_A_1186_21#_c_1480_n 0.00514288f $X=6.135 $Y=1.21
+ $X2=0 $Y2=0
cc_613 N_A_755_398#_c_608_n N_A_1186_21#_M1020_g 0.0128587f $X=7.105 $Y=1.73
+ $X2=0 $Y2=0
cc_614 N_A_755_398#_M1004_g N_A_1186_21#_M1020_g 0.0136878f $X=7.105 $Y=2.315
+ $X2=0 $Y2=0
cc_615 N_A_755_398#_c_651_p N_A_1186_21#_M1020_g 0.00331525f $X=5.85 $Y=2.31
+ $X2=0 $Y2=0
cc_616 N_A_755_398#_c_610_n N_A_1186_21#_M1020_g 0.00301824f $X=6.135 $Y=1.21
+ $X2=0 $Y2=0
cc_617 N_A_755_398#_c_659_p N_A_1186_21#_M1020_g 0.0127206f $X=6.375 $Y=2 $X2=0
+ $Y2=0
cc_618 N_A_755_398#_c_611_n N_A_1186_21#_M1020_g 0.00483974f $X=6.22 $Y=1.435
+ $X2=0 $Y2=0
cc_619 N_A_755_398#_c_620_n N_A_1186_21#_M1020_g 0.00505703f $X=6.46 $Y=1.915
+ $X2=0 $Y2=0
cc_620 N_A_755_398#_c_612_n N_A_1186_21#_M1020_g 0.0147602f $X=6.545 $Y=1.565
+ $X2=0 $Y2=0
cc_621 N_A_755_398#_c_619_n N_VPWR_M1010_d 0.00169035f $X=4.245 $Y=1.92 $X2=0
+ $Y2=0
cc_622 N_A_755_398#_c_649_p N_VPWR_M1010_d 0.0191732f $X=5.685 $Y=2.395 $X2=0
+ $Y2=0
cc_623 N_A_755_398#_c_716_p N_VPWR_M1010_d 0.00572186f $X=4.345 $Y=2.395 $X2=0
+ $Y2=0
cc_624 N_A_755_398#_c_615_n N_VPWR_c_1681_n 0.00296255f $X=3.85 $Y=2.14 $X2=0
+ $Y2=0
cc_625 N_A_755_398#_c_649_p N_VPWR_c_1681_n 0.0248544f $X=5.685 $Y=2.395 $X2=0
+ $Y2=0
cc_626 N_A_755_398#_c_608_n N_VPWR_c_1682_n 0.00340166f $X=7.105 $Y=1.73 $X2=0
+ $Y2=0
cc_627 N_A_755_398#_M1004_g N_VPWR_c_1682_n 0.0182665f $X=7.105 $Y=2.315 $X2=0
+ $Y2=0
cc_628 N_A_755_398#_c_620_n N_VPWR_c_1682_n 0.00225528f $X=6.46 $Y=1.915 $X2=0
+ $Y2=0
cc_629 N_A_755_398#_c_613_n N_VPWR_c_1682_n 0.0218994f $X=7.015 $Y=1.565 $X2=0
+ $Y2=0
cc_630 N_A_755_398#_c_623_n N_VPWR_c_1693_n 0.00749462f $X=5.85 $Y=2.395 $X2=0
+ $Y2=0
cc_631 N_A_755_398#_c_615_n N_VPWR_c_1677_n 9.6081e-19 $X=3.85 $Y=2.14 $X2=0
+ $Y2=0
cc_632 N_A_755_398#_M1004_g N_VPWR_c_1677_n 7.88961e-19 $X=7.105 $Y=2.315 $X2=0
+ $Y2=0
cc_633 N_A_755_398#_c_649_p N_VPWR_c_1677_n 0.0313826f $X=5.685 $Y=2.395 $X2=0
+ $Y2=0
cc_634 N_A_755_398#_c_716_p N_VPWR_c_1677_n 0.00684441f $X=4.345 $Y=2.395 $X2=0
+ $Y2=0
cc_635 N_A_755_398#_c_623_n N_VPWR_c_1677_n 0.00907254f $X=5.85 $Y=2.395 $X2=0
+ $Y2=0
cc_636 N_A_755_398#_c_659_p A_1228_379# 0.0059188f $X=6.375 $Y=2 $X2=-0.19
+ $Y2=-0.245
cc_637 N_A_755_398#_M1031_g N_VGND_c_1933_n 0.0182126f $X=4.005 $Y=0.76 $X2=0
+ $Y2=0
cc_638 N_A_755_398#_M1005_g N_VGND_c_1934_n 0.0113215f $X=7.135 $Y=0.915 $X2=0
+ $Y2=0
cc_639 N_A_755_398#_M1031_g N_VGND_c_1938_n 0.00457115f $X=4.005 $Y=0.76 $X2=0
+ $Y2=0
cc_640 N_A_755_398#_M1031_g N_VGND_c_1947_n 0.00490658f $X=4.005 $Y=0.76 $X2=0
+ $Y2=0
cc_641 N_A_755_398#_M1005_g N_VGND_c_1947_n 7.88961e-19 $X=7.135 $Y=0.915 $X2=0
+ $Y2=0
cc_642 N_A_755_398#_M1017_d N_A_1013_66#_c_2066_n 0.00710661f $X=5.5 $Y=0.33
+ $X2=0 $Y2=0
cc_643 N_A_755_398#_c_610_n N_A_1013_66#_c_2066_n 0.00800995f $X=6.135 $Y=1.21
+ $X2=0 $Y2=0
cc_644 N_A_755_398#_c_614_n N_A_1013_66#_c_2066_n 0.0232515f $X=5.715 $Y=1.13
+ $X2=0 $Y2=0
cc_645 N_A_755_398#_c_614_n N_A_1013_66#_c_2059_n 0.00158693f $X=5.715 $Y=1.13
+ $X2=0 $Y2=0
cc_646 N_A_755_398#_c_610_n N_A_1013_66#_c_2064_n 0.0125012f $X=6.135 $Y=1.21
+ $X2=0 $Y2=0
cc_647 N_SET_B_M1024_g N_A_546_449#_M1017_g 0.0364448f $X=4.99 $Y=0.65 $X2=0
+ $Y2=0
cc_648 N_SET_B_c_763_n N_A_546_449#_c_903_n 2.00503e-19 $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_649 N_SET_B_c_765_n N_A_546_449#_c_903_n 0.0042644f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_650 N_SET_B_c_766_n N_A_546_449#_c_903_n 0.0133619f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_651 N_SET_B_M1037_g N_A_546_449#_c_905_n 0.00205036f $X=5.065 $Y=2.315 $X2=0
+ $Y2=0
cc_652 N_SET_B_c_763_n N_A_546_449#_c_905_n 0.00142005f $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_653 N_SET_B_c_765_n N_A_546_449#_c_905_n 0.0038462f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_654 N_SET_B_c_766_n N_A_546_449#_c_905_n 0.0132798f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_655 N_SET_B_M1037_g N_A_546_449#_c_958_n 0.013025f $X=5.065 $Y=2.315 $X2=0
+ $Y2=0
cc_656 N_SET_B_c_762_n N_A_546_449#_c_958_n 0.0064047f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_657 N_SET_B_c_763_n N_A_546_449#_c_958_n 0.00335371f $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_658 N_SET_B_c_765_n N_A_546_449#_c_958_n 0.00291689f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_659 N_SET_B_c_766_n N_A_546_449#_c_958_n 0.0147665f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_660 N_SET_B_M1037_g N_A_546_449#_c_915_n 0.00443444f $X=5.065 $Y=2.315 $X2=0
+ $Y2=0
cc_661 N_SET_B_c_763_n N_A_546_449#_c_915_n 0.00132093f $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_662 N_SET_B_c_766_n N_A_546_449#_c_915_n 0.00277181f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_663 N_SET_B_c_762_n N_A_546_449#_c_906_n 0.0108805f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_664 N_SET_B_c_763_n N_A_546_449#_c_906_n 0.00136642f $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_665 N_SET_B_c_765_n N_A_546_449#_c_906_n 9.39653e-19 $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_666 N_SET_B_c_766_n N_A_546_449#_c_906_n 0.0189935f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_667 N_SET_B_c_762_n N_A_546_449#_c_917_n 0.0168568f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_762_n N_A_546_449#_c_907_n 0.0039909f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_669 N_SET_B_c_765_n N_A_546_449#_c_907_n 0.0135659f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_670 N_SET_B_c_766_n N_A_546_449#_c_907_n 0.00208451f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_671 N_SET_B_M1037_g N_A_223_119#_c_1060_n 0.0100607f $X=5.065 $Y=2.315 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_762_n N_A_223_119#_c_1064_n 0.00665641f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_673 SET_B N_A_223_119#_c_1047_n 0.00355556f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_674 N_SET_B_c_762_n N_A_223_119#_c_1047_n 0.00248701f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_764_n N_A_223_119#_c_1047_n 8.21853e-19 $X=8.88 $Y=1.665 $X2=0
+ $Y2=0
cc_676 N_SET_B_c_762_n N_A_223_119#_c_1048_n 0.00661355f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_677 N_SET_B_M1026_g N_A_1741_137#_c_1212_n 0.0134836f $X=9.405 $Y=0.915 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_770_n N_A_1741_137#_M1000_g 0.010713f $X=9.675 $Y=2.18 $X2=0
+ $Y2=0
cc_679 N_SET_B_M1026_g N_A_1741_137#_c_1217_n 0.00880682f $X=9.405 $Y=0.915
+ $X2=0 $Y2=0
cc_680 SET_B N_A_1741_137#_c_1217_n 0.00199736f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_681 N_SET_B_c_762_n N_A_1741_137#_c_1217_n 8.4248e-19 $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_764_n N_A_1741_137#_c_1217_n 0.00186167f $X=8.88 $Y=1.665 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_770_n N_A_1741_137#_c_1228_n 0.011858f $X=9.675 $Y=2.18 $X2=0
+ $Y2=0
cc_684 N_SET_B_c_771_n N_A_1741_137#_c_1228_n 0.0156276f $X=9.675 $Y=2.105 $X2=0
+ $Y2=0
cc_685 SET_B N_A_1741_137#_c_1228_n 0.0418816f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_686 N_SET_B_c_764_n N_A_1741_137#_c_1228_n 0.00104962f $X=8.88 $Y=1.665 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_767_n N_A_1741_137#_c_1228_n 0.00429286f $X=9.415 $Y=1.665
+ $X2=0 $Y2=0
cc_688 N_SET_B_c_770_n N_A_1741_137#_c_1229_n 0.00588305f $X=9.675 $Y=2.18 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_771_n N_A_1741_137#_c_1229_n 0.00606012f $X=9.675 $Y=2.105
+ $X2=0 $Y2=0
cc_690 SET_B N_A_1741_137#_c_1229_n 0.00403704f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_691 N_SET_B_c_770_n N_A_1741_137#_c_1260_n 0.0107117f $X=9.675 $Y=2.18 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_770_n N_A_1741_137#_c_1234_n 0.00135358f $X=9.675 $Y=2.18 $X2=0
+ $Y2=0
cc_693 N_SET_B_c_771_n N_A_1741_137#_c_1234_n 0.00264702f $X=9.675 $Y=2.105
+ $X2=0 $Y2=0
cc_694 N_SET_B_c_769_n N_A_1741_137#_c_1222_n 0.00847531f $X=9.505 $Y=2.03 $X2=0
+ $Y2=0
cc_695 SET_B N_A_1741_137#_c_1222_n 0.0165421f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_696 N_SET_B_c_767_n N_A_1741_137#_c_1222_n 0.0180926f $X=9.415 $Y=1.665 $X2=0
+ $Y2=0
cc_697 N_SET_B_M1026_g N_A_1531_428#_M1001_g 0.0269478f $X=9.405 $Y=0.915 $X2=0
+ $Y2=0
cc_698 N_SET_B_c_771_n N_A_1531_428#_M1028_g 0.0218f $X=9.675 $Y=2.105 $X2=0
+ $Y2=0
cc_699 SET_B N_A_1531_428#_M1028_g 2.11699e-19 $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_700 N_SET_B_c_767_n N_A_1531_428#_M1028_g 0.00746385f $X=9.415 $Y=1.665 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_762_n N_A_1531_428#_c_1389_n 0.00851774f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_702 N_SET_B_M1026_g N_A_1531_428#_c_1382_n 0.015516f $X=9.405 $Y=0.915 $X2=0
+ $Y2=0
cc_703 SET_B N_A_1531_428#_c_1382_n 0.0550286f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_704 N_SET_B_c_762_n N_A_1531_428#_c_1382_n 0.0143652f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_764_n N_A_1531_428#_c_1382_n 0.00389788f $X=8.88 $Y=1.665 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_767_n N_A_1531_428#_c_1382_n 0.00436857f $X=9.415 $Y=1.665
+ $X2=0 $Y2=0
cc_707 N_SET_B_M1026_g N_A_1531_428#_c_1383_n 0.0025476f $X=9.405 $Y=0.915 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_762_n N_A_1531_428#_c_1384_n 0.0252389f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_762_n N_A_1531_428#_c_1385_n 0.00688499f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_710 N_SET_B_M1026_g N_A_1531_428#_c_1386_n 8.07861e-19 $X=9.405 $Y=0.915
+ $X2=0 $Y2=0
cc_711 SET_B N_A_1531_428#_c_1386_n 0.0219534f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_712 N_SET_B_c_767_n N_A_1531_428#_c_1386_n 9.91162e-19 $X=9.415 $Y=1.665
+ $X2=0 $Y2=0
cc_713 N_SET_B_M1026_g N_A_1531_428#_c_1387_n 0.00145966f $X=9.405 $Y=0.915
+ $X2=0 $Y2=0
cc_714 SET_B N_A_1531_428#_c_1387_n 3.48211e-19 $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_715 N_SET_B_c_767_n N_A_1531_428#_c_1387_n 0.0188435f $X=9.415 $Y=1.665 $X2=0
+ $Y2=0
cc_716 N_SET_B_M1026_g N_A_1186_21#_c_1477_n 0.0101494f $X=9.405 $Y=0.915 $X2=0
+ $Y2=0
cc_717 N_SET_B_M1037_g N_VPWR_c_1681_n 0.0068806f $X=5.065 $Y=2.315 $X2=0 $Y2=0
cc_718 N_SET_B_c_762_n N_VPWR_c_1682_n 0.00884806f $X=8.735 $Y=1.665 $X2=0 $Y2=0
cc_719 N_SET_B_c_770_n N_VPWR_c_1683_n 0.00827993f $X=9.675 $Y=2.18 $X2=0 $Y2=0
cc_720 N_SET_B_c_771_n N_VPWR_c_1683_n 5.42704e-19 $X=9.675 $Y=2.105 $X2=0 $Y2=0
cc_721 N_SET_B_c_770_n N_VPWR_c_1691_n 0.00549284f $X=9.675 $Y=2.18 $X2=0 $Y2=0
cc_722 N_SET_B_M1037_g N_VPWR_c_1677_n 9.39239e-19 $X=5.065 $Y=2.315 $X2=0 $Y2=0
cc_723 N_SET_B_c_770_n N_VPWR_c_1677_n 0.011183f $X=9.675 $Y=2.18 $X2=0 $Y2=0
cc_724 N_SET_B_M1024_g N_VGND_c_1933_n 0.00296535f $X=4.99 $Y=0.65 $X2=0 $Y2=0
cc_725 N_SET_B_M1026_g N_VGND_c_1935_n 0.00652941f $X=9.405 $Y=0.915 $X2=0 $Y2=0
cc_726 N_SET_B_M1024_g N_VGND_c_1943_n 0.0030132f $X=4.99 $Y=0.65 $X2=0 $Y2=0
cc_727 N_SET_B_M1024_g N_VGND_c_1947_n 0.00472126f $X=4.99 $Y=0.65 $X2=0 $Y2=0
cc_728 N_SET_B_M1026_g N_VGND_c_1947_n 7.85159e-19 $X=9.405 $Y=0.915 $X2=0 $Y2=0
cc_729 N_SET_B_M1024_g N_A_1013_66#_c_2059_n 0.00540799f $X=4.99 $Y=0.65 $X2=0
+ $Y2=0
cc_730 N_SET_B_c_762_n N_A_1013_66#_c_2059_n 0.00509508f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_731 N_SET_B_c_763_n N_A_1013_66#_c_2059_n 0.00176133f $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_732 N_SET_B_c_765_n N_A_1013_66#_c_2059_n 4.7521e-19 $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_733 N_SET_B_c_766_n N_A_1013_66#_c_2059_n 0.00393097f $X=4.975 $Y=1.57 $X2=0
+ $Y2=0
cc_734 N_SET_B_M1026_g N_A_1896_119#_c_2086_n 0.00754224f $X=9.405 $Y=0.915
+ $X2=0 $Y2=0
cc_735 N_A_546_449#_c_901_n N_A_223_119#_M1023_g 0.00340072f $X=3.165 $Y=2.225
+ $X2=0 $Y2=0
cc_736 N_A_546_449#_c_908_n N_A_223_119#_M1023_g 0.00395169f $X=3.085 $Y=0.74
+ $X2=0 $Y2=0
cc_737 N_A_546_449#_c_901_n N_A_223_119#_c_1056_n 0.00590579f $X=3.165 $Y=2.225
+ $X2=0 $Y2=0
cc_738 N_A_546_449#_c_901_n N_A_223_119#_c_1057_n 0.00969738f $X=3.165 $Y=2.225
+ $X2=0 $Y2=0
cc_739 N_A_546_449#_c_902_n N_A_223_119#_c_1057_n 8.72087e-19 $X=3.885 $Y=2.225
+ $X2=0 $Y2=0
cc_740 N_A_546_449#_c_919_n N_A_223_119#_c_1057_n 0.00594646f $X=3.41 $Y=2.455
+ $X2=0 $Y2=0
cc_741 N_A_546_449#_c_901_n N_A_223_119#_c_1058_n 0.00235928f $X=3.165 $Y=2.225
+ $X2=0 $Y2=0
cc_742 N_A_546_449#_c_919_n N_A_223_119#_c_1058_n 0.0014858f $X=3.41 $Y=2.455
+ $X2=0 $Y2=0
cc_743 N_A_546_449#_c_901_n N_A_223_119#_M1033_g 7.50406e-19 $X=3.165 $Y=2.225
+ $X2=0 $Y2=0
cc_744 N_A_546_449#_c_911_n N_A_223_119#_M1033_g 0.0111711f $X=3.8 $Y=2.31 $X2=0
+ $Y2=0
cc_745 N_A_546_449#_c_919_n N_A_223_119#_M1033_g 0.00768742f $X=3.41 $Y=2.455
+ $X2=0 $Y2=0
cc_746 N_A_546_449#_M1003_g N_A_223_119#_c_1060_n 0.0103003f $X=6.065 $Y=2.315
+ $X2=0 $Y2=0
cc_747 N_A_546_449#_c_911_n N_A_223_119#_c_1060_n 0.00290732f $X=3.8 $Y=2.31
+ $X2=0 $Y2=0
cc_748 N_A_546_449#_c_901_n N_A_223_119#_c_1052_n 0.00518338f $X=3.165 $Y=2.225
+ $X2=0 $Y2=0
cc_749 N_A_546_449#_c_902_n N_A_223_119#_c_1052_n 0.00103004f $X=3.885 $Y=2.225
+ $X2=0 $Y2=0
cc_750 N_A_546_449#_M1017_g N_A_1186_21#_c_1478_n 0.0262411f $X=5.425 $Y=0.65
+ $X2=0 $Y2=0
cc_751 N_A_546_449#_c_907_n N_A_1186_21#_c_1480_n 0.0135778f $X=5.79 $Y=1.57
+ $X2=0 $Y2=0
cc_752 N_A_546_449#_c_917_n N_A_1186_21#_M1020_g 2.5542e-19 $X=5.79 $Y=1.57
+ $X2=0 $Y2=0
cc_753 N_A_546_449#_c_907_n N_A_1186_21#_M1020_g 0.0762995f $X=5.79 $Y=1.57
+ $X2=0 $Y2=0
cc_754 N_A_546_449#_c_905_n N_VPWR_M1010_d 0.00117613f $X=4.61 $Y=1.96 $X2=0
+ $Y2=0
cc_755 N_A_546_449#_c_958_n N_VPWR_M1010_d 0.00925932f $X=5.335 $Y=2.045 $X2=0
+ $Y2=0
cc_756 N_A_546_449#_c_914_n N_VPWR_M1010_d 0.00144282f $X=4.695 $Y=2.045 $X2=0
+ $Y2=0
cc_757 N_A_546_449#_c_919_n N_VPWR_c_1689_n 0.00627379f $X=3.41 $Y=2.455 $X2=0
+ $Y2=0
cc_758 N_A_546_449#_M1003_g N_VPWR_c_1677_n 9.39239e-19 $X=6.065 $Y=2.315 $X2=0
+ $Y2=0
cc_759 N_A_546_449#_c_919_n N_VPWR_c_1677_n 0.00961952f $X=3.41 $Y=2.455 $X2=0
+ $Y2=0
cc_760 N_A_546_449#_c_901_n N_A_460_449#_c_1820_n 0.00792442f $X=3.165 $Y=2.225
+ $X2=0 $Y2=0
cc_761 N_A_546_449#_c_908_n N_A_460_449#_c_1820_n 0.0141997f $X=3.085 $Y=0.74
+ $X2=0 $Y2=0
cc_762 N_A_546_449#_M1036_d N_A_460_449#_c_1821_n 5.87996e-19 $X=2.73 $Y=2.245
+ $X2=0 $Y2=0
cc_763 N_A_546_449#_c_919_n N_A_460_449#_c_1821_n 0.00657775f $X=3.41 $Y=2.455
+ $X2=0 $Y2=0
cc_764 N_A_546_449#_M1036_d N_A_460_449#_c_1824_n 0.00439139f $X=2.73 $Y=2.245
+ $X2=0 $Y2=0
cc_765 N_A_546_449#_c_919_n N_A_460_449#_c_1824_n 0.0216238f $X=3.41 $Y=2.455
+ $X2=0 $Y2=0
cc_766 N_A_546_449#_c_901_n N_A_460_449#_c_1822_n 0.078061f $X=3.165 $Y=2.225
+ $X2=0 $Y2=0
cc_767 N_A_546_449#_c_911_n A_707_449# 0.00291917f $X=3.8 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_768 N_A_546_449#_c_908_n N_VGND_c_1938_n 0.00825626f $X=3.085 $Y=0.74 $X2=0
+ $Y2=0
cc_769 N_A_546_449#_M1017_g N_VGND_c_1943_n 0.0030132f $X=5.425 $Y=0.65 $X2=0
+ $Y2=0
cc_770 N_A_546_449#_M1017_g N_VGND_c_1947_n 0.00439052f $X=5.425 $Y=0.65 $X2=0
+ $Y2=0
cc_771 N_A_546_449#_c_908_n N_VGND_c_1947_n 0.00933227f $X=3.085 $Y=0.74 $X2=0
+ $Y2=0
cc_772 N_A_546_449#_M1017_g N_A_1013_66#_c_2066_n 0.0122347f $X=5.425 $Y=0.65
+ $X2=0 $Y2=0
cc_773 N_A_546_449#_c_907_n N_A_1013_66#_c_2066_n 8.77006e-19 $X=5.79 $Y=1.57
+ $X2=0 $Y2=0
cc_774 N_A_546_449#_M1017_g N_A_1013_66#_c_2059_n 0.00536738f $X=5.425 $Y=0.65
+ $X2=0 $Y2=0
cc_775 N_A_546_449#_c_906_n N_A_1013_66#_c_2059_n 0.00111074f $X=5.505 $Y=1.605
+ $X2=0 $Y2=0
cc_776 N_A_223_119#_c_1050_n N_A_1741_137#_c_1212_n 0.0211871f $X=8.39 $Y=1.31
+ $X2=0 $Y2=0
cc_777 N_A_223_119#_c_1048_n N_A_1741_137#_c_1217_n 0.0211871f $X=8.315 $Y=1.385
+ $X2=0 $Y2=0
cc_778 N_A_223_119#_M1021_g N_A_1531_428#_c_1389_n 0.00418066f $X=7.58 $Y=2.56
+ $X2=0 $Y2=0
cc_779 N_A_223_119#_c_1063_n N_A_1531_428#_c_1389_n 0.00926013f $X=7.96 $Y=1.99
+ $X2=0 $Y2=0
cc_780 N_A_223_119#_c_1050_n N_A_1531_428#_c_1381_n 0.00660346f $X=8.39 $Y=1.31
+ $X2=0 $Y2=0
cc_781 N_A_223_119#_c_1048_n N_A_1531_428#_c_1382_n 0.00392507f $X=8.315
+ $Y=1.385 $X2=0 $Y2=0
cc_782 N_A_223_119#_c_1050_n N_A_1531_428#_c_1382_n 0.0127472f $X=8.39 $Y=1.31
+ $X2=0 $Y2=0
cc_783 N_A_223_119#_M1021_g N_A_1531_428#_c_1384_n 5.16583e-19 $X=7.58 $Y=2.56
+ $X2=0 $Y2=0
cc_784 N_A_223_119#_c_1063_n N_A_1531_428#_c_1384_n 0.0110069f $X=7.96 $Y=1.99
+ $X2=0 $Y2=0
cc_785 N_A_223_119#_c_1047_n N_A_1531_428#_c_1384_n 0.018037f $X=8.035 $Y=1.915
+ $X2=0 $Y2=0
cc_786 N_A_223_119#_c_1049_n N_A_1531_428#_c_1384_n 0.00475344f $X=8.11 $Y=1.385
+ $X2=0 $Y2=0
cc_787 N_A_223_119#_c_1048_n N_A_1531_428#_c_1385_n 0.0063708f $X=8.315 $Y=1.385
+ $X2=0 $Y2=0
cc_788 N_A_223_119#_c_1049_n N_A_1531_428#_c_1385_n 0.00414556f $X=8.11 $Y=1.385
+ $X2=0 $Y2=0
cc_789 N_A_223_119#_c_1050_n N_A_1186_21#_c_1477_n 0.00495681f $X=8.39 $Y=1.31
+ $X2=0 $Y2=0
cc_790 N_A_223_119#_c_1060_n N_A_1186_21#_M1020_g 0.0104164f $X=7.505 $Y=3.15
+ $X2=0 $Y2=0
cc_791 N_A_223_119#_c_1069_n N_VPWR_c_1680_n 0.0258905f $X=1.37 $Y=2.39 $X2=0
+ $Y2=0
cc_792 N_A_223_119#_c_1070_n N_VPWR_c_1680_n 0.0260518f $X=2.29 $Y=1.96 $X2=0
+ $Y2=0
cc_793 N_A_223_119#_c_1060_n N_VPWR_c_1681_n 0.0253641f $X=7.505 $Y=3.15 $X2=0
+ $Y2=0
cc_794 N_A_223_119#_c_1060_n N_VPWR_c_1682_n 0.0256899f $X=7.505 $Y=3.15 $X2=0
+ $Y2=0
cc_795 N_A_223_119#_M1021_g N_VPWR_c_1682_n 0.00130027f $X=7.58 $Y=2.56 $X2=0
+ $Y2=0
cc_796 N_A_223_119#_c_1064_n N_VPWR_c_1682_n 8.45453e-19 $X=7.655 $Y=1.99 $X2=0
+ $Y2=0
cc_797 N_A_223_119#_c_1069_n N_VPWR_c_1687_n 0.0111657f $X=1.37 $Y=2.39 $X2=0
+ $Y2=0
cc_798 N_A_223_119#_c_1061_n N_VPWR_c_1689_n 0.0436552f $X=3.535 $Y=3.15 $X2=0
+ $Y2=0
cc_799 N_A_223_119#_c_1060_n N_VPWR_c_1693_n 0.0594415f $X=7.505 $Y=3.15 $X2=0
+ $Y2=0
cc_800 N_A_223_119#_c_1060_n N_VPWR_c_1694_n 0.0175991f $X=7.505 $Y=3.15 $X2=0
+ $Y2=0
cc_801 N_A_223_119#_c_1060_n N_VPWR_c_1677_n 0.130228f $X=7.505 $Y=3.15 $X2=0
+ $Y2=0
cc_802 N_A_223_119#_c_1061_n N_VPWR_c_1677_n 0.0104273f $X=3.535 $Y=3.15 $X2=0
+ $Y2=0
cc_803 N_A_223_119#_c_1069_n N_VPWR_c_1677_n 0.0114323f $X=1.37 $Y=2.39 $X2=0
+ $Y2=0
cc_804 N_A_223_119#_M1023_g N_A_460_449#_c_1820_n 0.00882143f $X=2.79 $Y=0.805
+ $X2=0 $Y2=0
cc_805 N_A_223_119#_M1023_g N_A_460_449#_c_1821_n 0.00570686f $X=2.79 $Y=0.805
+ $X2=0 $Y2=0
cc_806 N_A_223_119#_c_1056_n N_A_460_449#_c_1821_n 0.00627643f $X=3.045 $Y=2.02
+ $X2=0 $Y2=0
cc_807 N_A_223_119#_M1033_g N_A_460_449#_c_1821_n 2.38835e-19 $X=3.46 $Y=2.455
+ $X2=0 $Y2=0
cc_808 N_A_223_119#_c_1052_n N_A_460_449#_c_1821_n 0.0174195f $X=2.79 $Y=1.66
+ $X2=0 $Y2=0
cc_809 N_A_223_119#_c_1070_n N_A_460_449#_c_1821_n 0.0137875f $X=2.29 $Y=1.96
+ $X2=0 $Y2=0
cc_810 N_A_223_119#_c_1054_n N_A_460_449#_c_1821_n 0.0269053f $X=2.455 $Y=1.645
+ $X2=0 $Y2=0
cc_811 N_A_223_119#_c_1051_n N_A_460_449#_c_1824_n 0.00164568f $X=2.715 $Y=1.645
+ $X2=0 $Y2=0
cc_812 N_A_223_119#_c_1070_n N_A_460_449#_c_1824_n 0.0147448f $X=2.29 $Y=1.96
+ $X2=0 $Y2=0
cc_813 N_A_223_119#_M1023_g N_A_460_449#_c_1822_n 0.0130223f $X=2.79 $Y=0.805
+ $X2=0 $Y2=0
cc_814 N_A_223_119#_c_1051_n N_A_460_449#_c_1822_n 0.00826811f $X=2.715 $Y=1.645
+ $X2=0 $Y2=0
cc_815 N_A_223_119#_c_1054_n N_A_460_449#_c_1822_n 0.0116251f $X=2.455 $Y=1.645
+ $X2=0 $Y2=0
cc_816 N_A_223_119#_c_1055_n N_VGND_c_1932_n 0.0159918f $X=1.25 $Y=0.795 $X2=0
+ $Y2=0
cc_817 N_A_223_119#_c_1055_n N_VGND_c_1942_n 0.00738991f $X=1.25 $Y=0.795 $X2=0
+ $Y2=0
cc_818 N_A_223_119#_M1023_g N_VGND_c_1947_n 9.39239e-19 $X=2.79 $Y=0.805 $X2=0
+ $Y2=0
cc_819 N_A_223_119#_c_1050_n N_VGND_c_1947_n 9.72468e-19 $X=8.39 $Y=1.31 $X2=0
+ $Y2=0
cc_820 N_A_223_119#_c_1055_n N_VGND_c_1947_n 0.0101824f $X=1.25 $Y=0.795 $X2=0
+ $Y2=0
cc_821 N_A_1741_137#_c_1219_n N_A_1531_428#_M1001_g 0.00382463f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_822 N_A_1741_137#_c_1269_p N_A_1531_428#_M1001_g 0.00391488f $X=10.13 $Y=0.79
+ $X2=0 $Y2=0
cc_823 N_A_1741_137#_c_1260_n N_A_1531_428#_M1028_g 0.0122826f $X=9.89 $Y=2.4
+ $X2=0 $Y2=0
cc_824 N_A_1741_137#_c_1230_n N_A_1531_428#_M1028_g 0.0130346f $X=10.3 $Y=2.29
+ $X2=0 $Y2=0
cc_825 N_A_1741_137#_c_1234_n N_A_1531_428#_M1028_g 0.0050702f $X=9.89 $Y=2.235
+ $X2=0 $Y2=0
cc_826 N_A_1741_137#_c_1212_n N_A_1531_428#_c_1382_n 0.0127607f $X=8.78 $Y=1.31
+ $X2=0 $Y2=0
cc_827 N_A_1741_137#_c_1217_n N_A_1531_428#_c_1382_n 0.0071292f $X=8.935
+ $Y=1.385 $X2=0 $Y2=0
cc_828 N_A_1741_137#_c_1219_n N_A_1531_428#_c_1382_n 0.00742332f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_829 N_A_1741_137#_c_1219_n N_A_1531_428#_c_1383_n 0.00575516f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_830 N_A_1741_137#_c_1217_n N_A_1531_428#_c_1384_n 4.90084e-19 $X=8.935
+ $Y=1.385 $X2=0 $Y2=0
cc_831 N_A_1741_137#_c_1230_n N_A_1531_428#_c_1386_n 0.00224246f $X=10.3 $Y=2.29
+ $X2=0 $Y2=0
cc_832 N_A_1741_137#_c_1219_n N_A_1531_428#_c_1386_n 0.0238005f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_833 N_A_1741_137#_c_1234_n N_A_1531_428#_c_1386_n 0.016233f $X=9.89 $Y=2.235
+ $X2=0 $Y2=0
cc_834 N_A_1741_137#_c_1269_p N_A_1531_428#_c_1386_n 0.00425108f $X=10.13
+ $Y=0.79 $X2=0 $Y2=0
cc_835 N_A_1741_137#_c_1219_n N_A_1531_428#_c_1387_n 0.011765f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_836 N_A_1741_137#_c_1234_n N_A_1531_428#_c_1387_n 0.00578013f $X=9.89
+ $Y=2.235 $X2=0 $Y2=0
cc_837 N_A_1741_137#_c_1269_p N_A_1531_428#_c_1387_n 0.00476386f $X=10.13
+ $Y=0.79 $X2=0 $Y2=0
cc_838 N_A_1741_137#_c_1232_n N_A_1186_21#_M1007_s 0.00307548f $X=11.725 $Y=2.29
+ $X2=0 $Y2=0
cc_839 N_A_1741_137#_c_1212_n N_A_1186_21#_c_1477_n 0.00495681f $X=8.78 $Y=1.31
+ $X2=0 $Y2=0
cc_840 N_A_1741_137#_c_1219_n N_A_1186_21#_M1014_g 0.0040442f $X=10.385 $Y=2.205
+ $X2=0 $Y2=0
cc_841 N_A_1741_137#_c_1269_p N_A_1186_21#_M1014_g 0.0084807f $X=10.13 $Y=0.79
+ $X2=0 $Y2=0
cc_842 N_A_1741_137#_c_1260_n N_A_1186_21#_c_1490_n 0.00216242f $X=9.89 $Y=2.4
+ $X2=0 $Y2=0
cc_843 N_A_1741_137#_c_1219_n N_A_1186_21#_c_1490_n 0.00112394f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_844 N_A_1741_137#_c_1232_n N_A_1186_21#_c_1490_n 0.0101369f $X=11.725 $Y=2.29
+ $X2=0 $Y2=0
cc_845 N_A_1741_137#_c_1292_p N_A_1186_21#_c_1490_n 0.0069047f $X=10.385 $Y=2.29
+ $X2=0 $Y2=0
cc_846 N_A_1741_137#_c_1219_n N_A_1186_21#_c_1483_n 0.00344532f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_847 N_A_1741_137#_c_1219_n N_A_1186_21#_c_1484_n 0.00718731f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_848 N_A_1741_137#_c_1219_n N_A_1186_21#_c_1485_n 9.13136e-19 $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_849 N_A_1741_137#_c_1219_n N_A_1186_21#_c_1492_n 0.00975664f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_850 N_A_1741_137#_c_1232_n N_A_1186_21#_c_1492_n 0.00912637f $X=11.725
+ $Y=2.29 $X2=0 $Y2=0
cc_851 N_A_1741_137#_c_1219_n N_A_1186_21#_c_1487_n 0.0487934f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_852 N_A_1741_137#_c_1219_n N_A_1186_21#_c_1494_n 0.0252514f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_853 N_A_1741_137#_c_1232_n N_A_1186_21#_c_1494_n 0.0259892f $X=11.725 $Y=2.29
+ $X2=0 $Y2=0
cc_854 N_A_1741_137#_M1011_g N_A_1186_21#_c_1495_n 2.92461e-19 $X=11.945
+ $Y=2.345 $X2=0 $Y2=0
cc_855 N_A_1741_137#_c_1232_n N_A_1186_21#_c_1495_n 0.0259734f $X=11.725 $Y=2.29
+ $X2=0 $Y2=0
cc_856 N_A_1741_137#_c_1220_n N_A_1186_21#_c_1495_n 0.0152803f $X=11.81 $Y=2.205
+ $X2=0 $Y2=0
cc_857 N_A_1741_137#_c_1219_n N_A_1186_21#_c_1488_n 0.00304667f $X=10.385
+ $Y=2.205 $X2=0 $Y2=0
cc_858 N_A_1741_137#_c_1232_n N_A_1186_21#_c_1488_n 4.62084e-19 $X=11.725
+ $Y=2.29 $X2=0 $Y2=0
cc_859 N_A_1741_137#_M1011_g N_RESET_B_M1007_g 0.0299287f $X=11.945 $Y=2.345
+ $X2=0 $Y2=0
cc_860 N_A_1741_137#_c_1232_n N_RESET_B_M1007_g 0.0203522f $X=11.725 $Y=2.29
+ $X2=0 $Y2=0
cc_861 N_A_1741_137#_c_1220_n N_RESET_B_M1007_g 0.00984648f $X=11.81 $Y=2.205
+ $X2=0 $Y2=0
cc_862 N_A_1741_137#_c_1221_n RESET_B 0.0230292f $X=11.92 $Y=1.35 $X2=0 $Y2=0
cc_863 N_A_1741_137#_c_1223_n RESET_B 3.9254e-19 $X=11.92 $Y=1.26 $X2=0 $Y2=0
cc_864 N_A_1741_137#_c_1221_n N_RESET_B_c_1598_n 0.00117707f $X=11.92 $Y=1.35
+ $X2=0 $Y2=0
cc_865 N_A_1741_137#_c_1223_n N_RESET_B_c_1598_n 0.0186835f $X=11.92 $Y=1.26
+ $X2=0 $Y2=0
cc_866 N_A_1741_137#_c_1224_n N_RESET_B_c_1599_n 0.0133137f $X=11.92 $Y=1.185
+ $X2=0 $Y2=0
cc_867 N_A_1741_137#_c_1215_n N_A_2511_137#_M1035_g 0.0153889f $X=12.915
+ $Y=1.185 $X2=0 $Y2=0
cc_868 N_A_1741_137#_M1019_g N_A_2511_137#_M1016_g 0.0167472f $X=12.915 $Y=2.155
+ $X2=0 $Y2=0
cc_869 N_A_1741_137#_c_1214_n N_A_2511_137#_c_1630_n 0.0072312f $X=12.84 $Y=1.26
+ $X2=0 $Y2=0
cc_870 N_A_1741_137#_c_1215_n N_A_2511_137#_c_1630_n 0.00878607f $X=12.915
+ $Y=1.185 $X2=0 $Y2=0
cc_871 N_A_1741_137#_c_1218_n N_A_2511_137#_c_1630_n 0.00226016f $X=12.915
+ $Y=1.26 $X2=0 $Y2=0
cc_872 N_A_1741_137#_c_1224_n N_A_2511_137#_c_1630_n 4.17281e-19 $X=11.92
+ $Y=1.185 $X2=0 $Y2=0
cc_873 N_A_1741_137#_M1011_g N_A_2511_137#_c_1635_n 0.00155041f $X=11.945
+ $Y=2.345 $X2=0 $Y2=0
cc_874 N_A_1741_137#_M1019_g N_A_2511_137#_c_1635_n 0.0151894f $X=12.915
+ $Y=2.155 $X2=0 $Y2=0
cc_875 N_A_1741_137#_M1019_g N_A_2511_137#_c_1631_n 0.0120704f $X=12.915
+ $Y=2.155 $X2=0 $Y2=0
cc_876 N_A_1741_137#_c_1218_n N_A_2511_137#_c_1631_n 0.00652629f $X=12.915
+ $Y=1.26 $X2=0 $Y2=0
cc_877 N_A_1741_137#_c_1218_n N_A_2511_137#_c_1632_n 0.0213246f $X=12.915
+ $Y=1.26 $X2=0 $Y2=0
cc_878 N_A_1741_137#_c_1214_n N_A_2511_137#_c_1633_n 0.00657016f $X=12.84
+ $Y=1.26 $X2=0 $Y2=0
cc_879 N_A_1741_137#_M1019_g N_A_2511_137#_c_1633_n 0.00634186f $X=12.915
+ $Y=2.155 $X2=0 $Y2=0
cc_880 N_A_1741_137#_c_1228_n N_VPWR_M1000_d 0.00225286f $X=9.725 $Y=2.235 $X2=0
+ $Y2=0
cc_881 N_A_1741_137#_c_1232_n N_VPWR_M1013_d 0.00308676f $X=11.725 $Y=2.29 $X2=0
+ $Y2=0
cc_882 N_A_1741_137#_c_1232_n N_VPWR_M1007_d 0.00824504f $X=11.725 $Y=2.29 $X2=0
+ $Y2=0
cc_883 N_A_1741_137#_c_1220_n N_VPWR_M1007_d 0.00561339f $X=11.81 $Y=2.205 $X2=0
+ $Y2=0
cc_884 N_A_1741_137#_M1000_g N_VPWR_c_1683_n 0.00755813f $X=8.965 $Y=2.77 $X2=0
+ $Y2=0
cc_885 N_A_1741_137#_c_1228_n N_VPWR_c_1683_n 0.026891f $X=9.725 $Y=2.235 $X2=0
+ $Y2=0
cc_886 N_A_1741_137#_c_1260_n N_VPWR_c_1684_n 0.0170632f $X=9.89 $Y=2.4 $X2=0
+ $Y2=0
cc_887 N_A_1741_137#_c_1232_n N_VPWR_c_1684_n 0.0210759f $X=11.725 $Y=2.29 $X2=0
+ $Y2=0
cc_888 N_A_1741_137#_M1011_g N_VPWR_c_1685_n 0.0132198f $X=11.945 $Y=2.345 $X2=0
+ $Y2=0
cc_889 N_A_1741_137#_c_1232_n N_VPWR_c_1685_n 0.0219318f $X=11.725 $Y=2.29 $X2=0
+ $Y2=0
cc_890 N_A_1741_137#_M1019_g N_VPWR_c_1686_n 0.00524354f $X=12.915 $Y=2.155
+ $X2=0 $Y2=0
cc_891 N_A_1741_137#_c_1260_n N_VPWR_c_1691_n 0.0177952f $X=9.89 $Y=2.4 $X2=0
+ $Y2=0
cc_892 N_A_1741_137#_M1000_g N_VPWR_c_1694_n 0.00478016f $X=8.965 $Y=2.77 $X2=0
+ $Y2=0
cc_893 N_A_1741_137#_M1011_g N_VPWR_c_1696_n 0.00393414f $X=11.945 $Y=2.345
+ $X2=0 $Y2=0
cc_894 N_A_1741_137#_M1019_g N_VPWR_c_1696_n 0.00312414f $X=12.915 $Y=2.155
+ $X2=0 $Y2=0
cc_895 N_A_1741_137#_M1015_d N_VPWR_c_1677_n 0.00223819f $X=9.75 $Y=2.255 $X2=0
+ $Y2=0
cc_896 N_A_1741_137#_M1000_g N_VPWR_c_1677_n 0.00969176f $X=8.965 $Y=2.77 $X2=0
+ $Y2=0
cc_897 N_A_1741_137#_M1011_g N_VPWR_c_1677_n 0.00787963f $X=11.945 $Y=2.345
+ $X2=0 $Y2=0
cc_898 N_A_1741_137#_M1019_g N_VPWR_c_1677_n 0.00410284f $X=12.915 $Y=2.155
+ $X2=0 $Y2=0
cc_899 N_A_1741_137#_c_1260_n N_VPWR_c_1677_n 0.0123247f $X=9.89 $Y=2.4 $X2=0
+ $Y2=0
cc_900 N_A_1741_137#_c_1230_n A_2036_451# 0.00236564f $X=10.3 $Y=2.29 $X2=-0.19
+ $Y2=-0.245
cc_901 N_A_1741_137#_c_1292_p A_2036_451# 0.00148865f $X=10.385 $Y=2.29
+ $X2=-0.19 $Y2=-0.245
cc_902 N_A_1741_137#_c_1215_n N_Q_N_c_1872_n 0.00334021f $X=12.915 $Y=1.185
+ $X2=0 $Y2=0
cc_903 N_A_1741_137#_c_1224_n N_Q_N_c_1872_n 0.00609048f $X=11.92 $Y=1.185 $X2=0
+ $Y2=0
cc_904 N_A_1741_137#_c_1214_n N_Q_N_c_1873_n 0.00711665f $X=12.84 $Y=1.26 $X2=0
+ $Y2=0
cc_905 N_A_1741_137#_c_1221_n N_Q_N_c_1873_n 0.00605347f $X=11.92 $Y=1.35 $X2=0
+ $Y2=0
cc_906 N_A_1741_137#_c_1224_n N_Q_N_c_1873_n 0.00279956f $X=11.92 $Y=1.185 $X2=0
+ $Y2=0
cc_907 N_A_1741_137#_M1011_g N_Q_N_c_1875_n 0.00453786f $X=11.945 $Y=2.345 $X2=0
+ $Y2=0
cc_908 N_A_1741_137#_c_1214_n N_Q_N_c_1875_n 0.00605641f $X=12.84 $Y=1.26 $X2=0
+ $Y2=0
cc_909 N_A_1741_137#_c_1220_n N_Q_N_c_1875_n 0.0172466f $X=11.81 $Y=2.205 $X2=0
+ $Y2=0
cc_910 N_A_1741_137#_c_1221_n N_Q_N_c_1875_n 7.27024e-19 $X=11.92 $Y=1.35 $X2=0
+ $Y2=0
cc_911 N_A_1741_137#_c_1223_n N_Q_N_c_1875_n 2.43744e-19 $X=11.92 $Y=1.26 $X2=0
+ $Y2=0
cc_912 N_A_1741_137#_M1011_g N_Q_N_c_1874_n 0.00250731f $X=11.945 $Y=2.345 $X2=0
+ $Y2=0
cc_913 N_A_1741_137#_c_1214_n N_Q_N_c_1874_n 0.0146609f $X=12.84 $Y=1.26 $X2=0
+ $Y2=0
cc_914 N_A_1741_137#_M1019_g N_Q_N_c_1874_n 0.00341839f $X=12.915 $Y=2.155 $X2=0
+ $Y2=0
cc_915 N_A_1741_137#_c_1220_n N_Q_N_c_1874_n 0.00519375f $X=11.81 $Y=2.205 $X2=0
+ $Y2=0
cc_916 N_A_1741_137#_c_1221_n N_Q_N_c_1874_n 0.0233178f $X=11.92 $Y=1.35 $X2=0
+ $Y2=0
cc_917 N_A_1741_137#_c_1223_n N_Q_N_c_1874_n 0.00124625f $X=11.92 $Y=1.26 $X2=0
+ $Y2=0
cc_918 N_A_1741_137#_c_1224_n N_Q_N_c_1874_n 0.00400465f $X=11.92 $Y=1.185 $X2=0
+ $Y2=0
cc_919 N_A_1741_137#_M1019_g Q_N 0.00202202f $X=12.915 $Y=2.155 $X2=0 $Y2=0
cc_920 N_A_1741_137#_c_1212_n N_VGND_c_1935_n 0.00803036f $X=8.78 $Y=1.31 $X2=0
+ $Y2=0
cc_921 N_A_1741_137#_c_1217_n N_VGND_c_1935_n 3.43708e-19 $X=8.935 $Y=1.385
+ $X2=0 $Y2=0
cc_922 N_A_1741_137#_c_1221_n N_VGND_c_1936_n 0.00541978f $X=11.92 $Y=1.35 $X2=0
+ $Y2=0
cc_923 N_A_1741_137#_c_1223_n N_VGND_c_1936_n 8.98567e-19 $X=11.92 $Y=1.26 $X2=0
+ $Y2=0
cc_924 N_A_1741_137#_c_1224_n N_VGND_c_1936_n 0.00483983f $X=11.92 $Y=1.185
+ $X2=0 $Y2=0
cc_925 N_A_1741_137#_c_1215_n N_VGND_c_1937_n 0.00409263f $X=12.915 $Y=1.185
+ $X2=0 $Y2=0
cc_926 N_A_1741_137#_c_1215_n N_VGND_c_1945_n 0.00371502f $X=12.915 $Y=1.185
+ $X2=0 $Y2=0
cc_927 N_A_1741_137#_c_1224_n N_VGND_c_1945_n 0.00549284f $X=11.92 $Y=1.185
+ $X2=0 $Y2=0
cc_928 N_A_1741_137#_c_1212_n N_VGND_c_1947_n 9.72468e-19 $X=8.78 $Y=1.31 $X2=0
+ $Y2=0
cc_929 N_A_1741_137#_c_1215_n N_VGND_c_1947_n 0.00453162f $X=12.915 $Y=1.185
+ $X2=0 $Y2=0
cc_930 N_A_1741_137#_c_1224_n N_VGND_c_1947_n 0.0123926f $X=11.92 $Y=1.185 $X2=0
+ $Y2=0
cc_931 N_A_1741_137#_M1001_d N_A_1896_119#_c_2087_n 0.00229129f $X=9.97 $Y=0.595
+ $X2=0 $Y2=0
cc_932 N_A_1741_137#_c_1269_p N_A_1896_119#_c_2087_n 0.0218947f $X=10.13 $Y=0.79
+ $X2=0 $Y2=0
cc_933 N_A_1531_428#_M1001_g N_A_1186_21#_c_1477_n 0.00881852f $X=9.895 $Y=0.915
+ $X2=0 $Y2=0
cc_934 N_A_1531_428#_c_1381_n N_A_1186_21#_c_1477_n 0.00666278f $X=8.095 $Y=0.74
+ $X2=0 $Y2=0
cc_935 N_A_1531_428#_M1001_g N_A_1186_21#_M1014_g 0.014615f $X=9.895 $Y=0.915
+ $X2=0 $Y2=0
cc_936 N_A_1531_428#_c_1382_n N_A_1186_21#_c_1484_n 4.49431e-19 $X=9.775
+ $Y=1.235 $X2=0 $Y2=0
cc_937 N_A_1531_428#_M1028_g N_A_1186_21#_c_1485_n 0.00446321f $X=10.105
+ $Y=2.675 $X2=0 $Y2=0
cc_938 N_A_1531_428#_M1028_g N_A_1186_21#_c_1492_n 0.0720151f $X=10.105 $Y=2.675
+ $X2=0 $Y2=0
cc_939 N_A_1531_428#_M1001_g N_A_1186_21#_c_1488_n 0.00120779f $X=9.895 $Y=0.915
+ $X2=0 $Y2=0
cc_940 N_A_1531_428#_c_1387_n N_A_1186_21#_c_1488_n 0.00446321f $X=10.105
+ $Y=1.625 $X2=0 $Y2=0
cc_941 N_A_1531_428#_M1028_g N_VPWR_c_1684_n 0.00267012f $X=10.105 $Y=2.675
+ $X2=0 $Y2=0
cc_942 N_A_1531_428#_M1028_g N_VPWR_c_1691_n 0.00549284f $X=10.105 $Y=2.675
+ $X2=0 $Y2=0
cc_943 N_A_1531_428#_M1028_g N_VPWR_c_1677_n 0.00987829f $X=10.105 $Y=2.675
+ $X2=0 $Y2=0
cc_944 N_A_1531_428#_c_1382_n N_VGND_M1006_d 0.00485776f $X=9.775 $Y=1.235 $X2=0
+ $Y2=0
cc_945 N_A_1531_428#_c_1382_n N_VGND_c_1935_n 0.025283f $X=9.775 $Y=1.235 $X2=0
+ $Y2=0
cc_946 N_A_1531_428#_c_1381_n N_VGND_c_1940_n 0.00755126f $X=8.095 $Y=0.74 $X2=0
+ $Y2=0
cc_947 N_A_1531_428#_c_1381_n N_VGND_c_1947_n 0.00910022f $X=8.095 $Y=0.74 $X2=0
+ $Y2=0
cc_948 N_A_1531_428#_c_1382_n A_1693_163# 0.0048076f $X=9.775 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_949 N_A_1531_428#_c_1382_n N_A_1896_119#_M1026_d 0.00246076f $X=9.775
+ $Y=1.235 $X2=-0.19 $Y2=-0.245
cc_950 N_A_1531_428#_M1001_g N_A_1896_119#_c_2086_n 0.00564135f $X=9.895
+ $Y=0.915 $X2=0 $Y2=0
cc_951 N_A_1531_428#_c_1382_n N_A_1896_119#_c_2086_n 0.0194208f $X=9.775
+ $Y=1.235 $X2=0 $Y2=0
cc_952 N_A_1531_428#_M1001_g N_A_1896_119#_c_2087_n 0.00368088f $X=9.895
+ $Y=0.915 $X2=0 $Y2=0
cc_953 N_A_1186_21#_c_1485_n N_RESET_B_M1007_g 0.00941845f $X=10.725 $Y=2.03
+ $X2=0 $Y2=0
cc_954 N_A_1186_21#_c_1487_n N_RESET_B_M1007_g 0.00361871f $X=10.815 $Y=1.35
+ $X2=0 $Y2=0
cc_955 N_A_1186_21#_c_1495_n N_RESET_B_M1007_g 0.00566222f $X=11.225 $Y=1.86
+ $X2=0 $Y2=0
cc_956 N_A_1186_21#_c_1486_n RESET_B 0.0134492f $X=10.815 $Y=1 $X2=0 $Y2=0
cc_957 N_A_1186_21#_c_1487_n RESET_B 0.0249904f $X=10.815 $Y=1.35 $X2=0 $Y2=0
cc_958 N_A_1186_21#_c_1495_n RESET_B 0.0170778f $X=11.225 $Y=1.86 $X2=0 $Y2=0
cc_959 N_A_1186_21#_c_1488_n RESET_B 0.00200279f $X=10.815 $Y=1.175 $X2=0 $Y2=0
cc_960 N_A_1186_21#_c_1486_n N_RESET_B_c_1598_n 9.4527e-19 $X=10.815 $Y=1 $X2=0
+ $Y2=0
cc_961 N_A_1186_21#_c_1487_n N_RESET_B_c_1598_n 3.92584e-19 $X=10.815 $Y=1.35
+ $X2=0 $Y2=0
cc_962 N_A_1186_21#_c_1495_n N_RESET_B_c_1598_n 0.00406126f $X=11.225 $Y=1.86
+ $X2=0 $Y2=0
cc_963 N_A_1186_21#_c_1488_n N_RESET_B_c_1598_n 0.0212551f $X=10.815 $Y=1.175
+ $X2=0 $Y2=0
cc_964 N_A_1186_21#_c_1486_n N_RESET_B_c_1599_n 0.00490526f $X=10.815 $Y=1 $X2=0
+ $Y2=0
cc_965 N_A_1186_21#_c_1487_n N_RESET_B_c_1599_n 0.00335526f $X=10.815 $Y=1.35
+ $X2=0 $Y2=0
cc_966 N_A_1186_21#_c_1488_n N_RESET_B_c_1599_n 0.00330647f $X=10.815 $Y=1.175
+ $X2=0 $Y2=0
cc_967 N_A_1186_21#_M1020_g N_VPWR_c_1682_n 0.0202718f $X=6.455 $Y=2.315 $X2=0
+ $Y2=0
cc_968 N_A_1186_21#_c_1490_n N_VPWR_c_1684_n 0.0179417f $X=10.465 $Y=2.18 $X2=0
+ $Y2=0
cc_969 N_A_1186_21#_c_1490_n N_VPWR_c_1691_n 0.00486043f $X=10.465 $Y=2.18 $X2=0
+ $Y2=0
cc_970 N_A_1186_21#_M1020_g N_VPWR_c_1677_n 9.39239e-19 $X=6.455 $Y=2.315 $X2=0
+ $Y2=0
cc_971 N_A_1186_21#_c_1490_n N_VPWR_c_1677_n 0.00818711f $X=10.465 $Y=2.18 $X2=0
+ $Y2=0
cc_972 N_A_1186_21#_c_1477_n N_VGND_c_1934_n 0.0211465f $X=10.295 $Y=0.18 $X2=0
+ $Y2=0
cc_973 N_A_1186_21#_c_1477_n N_VGND_c_1935_n 0.026083f $X=10.295 $Y=0.18 $X2=0
+ $Y2=0
cc_974 N_A_1186_21#_c_1486_n N_VGND_c_1936_n 0.0146485f $X=10.815 $Y=1 $X2=0
+ $Y2=0
cc_975 N_A_1186_21#_c_1477_n N_VGND_c_1940_n 0.0619124f $X=10.295 $Y=0.18 $X2=0
+ $Y2=0
cc_976 N_A_1186_21#_c_1478_n N_VGND_c_1943_n 0.0219031f $X=6.08 $Y=0.18 $X2=0
+ $Y2=0
cc_977 N_A_1186_21#_c_1477_n N_VGND_c_1944_n 0.0272727f $X=10.295 $Y=0.18 $X2=0
+ $Y2=0
cc_978 N_A_1186_21#_c_1486_n N_VGND_c_1944_n 0.00632222f $X=10.815 $Y=1 $X2=0
+ $Y2=0
cc_979 N_A_1186_21#_c_1477_n N_VGND_c_1947_n 0.135053f $X=10.295 $Y=0.18 $X2=0
+ $Y2=0
cc_980 N_A_1186_21#_c_1478_n N_VGND_c_1947_n 0.00569756f $X=6.08 $Y=0.18 $X2=0
+ $Y2=0
cc_981 N_A_1186_21#_c_1486_n N_VGND_c_1947_n 0.0189337f $X=10.815 $Y=1 $X2=0
+ $Y2=0
cc_982 N_A_1186_21#_M1012_g N_A_1013_66#_c_2066_n 0.00996469f $X=6.005 $Y=0.65
+ $X2=0 $Y2=0
cc_983 N_A_1186_21#_M1012_g N_A_1013_66#_c_2059_n 8.27039e-19 $X=6.005 $Y=0.65
+ $X2=0 $Y2=0
cc_984 N_A_1186_21#_c_1479_n N_A_1013_66#_c_2064_n 0.00358134f $X=6.38 $Y=1.12
+ $X2=0 $Y2=0
cc_985 N_A_1186_21#_c_1486_n N_A_1896_119#_M1014_d 0.00371196f $X=10.815 $Y=1
+ $X2=0 $Y2=0
cc_986 N_A_1186_21#_c_1487_n N_A_1896_119#_M1014_d 2.12115e-19 $X=10.815 $Y=1.35
+ $X2=0 $Y2=0
cc_987 N_A_1186_21#_M1014_g N_A_1896_119#_c_2086_n 0.00103384f $X=10.37 $Y=0.705
+ $X2=0 $Y2=0
cc_988 N_A_1186_21#_c_1477_n N_A_1896_119#_c_2087_n 0.00732302f $X=10.295
+ $Y=0.18 $X2=0 $Y2=0
cc_989 N_A_1186_21#_M1014_g N_A_1896_119#_c_2087_n 0.0127219f $X=10.37 $Y=0.705
+ $X2=0 $Y2=0
cc_990 N_A_1186_21#_c_1477_n N_A_1896_119#_c_2088_n 0.00770783f $X=10.295
+ $Y=0.18 $X2=0 $Y2=0
cc_991 N_A_1186_21#_M1014_g N_A_1896_119#_c_2089_n 0.00140971f $X=10.37 $Y=0.705
+ $X2=0 $Y2=0
cc_992 N_A_1186_21#_c_1483_n N_A_1896_119#_c_2089_n 0.00450911f $X=10.65
+ $Y=1.175 $X2=0 $Y2=0
cc_993 N_A_1186_21#_c_1486_n N_A_1896_119#_c_2089_n 0.0134462f $X=10.815 $Y=1
+ $X2=0 $Y2=0
cc_994 N_A_1186_21#_c_1488_n N_A_1896_119#_c_2089_n 6.26375e-19 $X=10.815
+ $Y=1.175 $X2=0 $Y2=0
cc_995 N_RESET_B_M1007_g N_VPWR_c_1677_n 0.0038268f $X=11.44 $Y=2.035 $X2=0
+ $Y2=0
cc_996 N_RESET_B_c_1599_n N_VGND_c_1936_n 0.00490854f $X=11.355 $Y=1.185 $X2=0
+ $Y2=0
cc_997 N_RESET_B_c_1599_n N_VGND_c_1944_n 0.00384813f $X=11.355 $Y=1.185 $X2=0
+ $Y2=0
cc_998 N_RESET_B_c_1599_n N_VGND_c_1947_n 0.0046122f $X=11.355 $Y=1.185 $X2=0
+ $Y2=0
cc_999 N_RESET_B_c_1599_n N_A_1896_119#_c_2089_n 0.0028454f $X=11.355 $Y=1.185
+ $X2=0 $Y2=0
cc_1000 N_A_2511_137#_M1016_g N_VPWR_c_1686_n 0.00698192f $X=13.425 $Y=2.465
+ $X2=0 $Y2=0
cc_1001 N_A_2511_137#_c_1635_n N_VPWR_c_1686_n 0.0248129f $X=12.7 $Y=1.98 $X2=0
+ $Y2=0
cc_1002 N_A_2511_137#_c_1631_n N_VPWR_c_1686_n 0.0206753f $X=13.365 $Y=1.47
+ $X2=0 $Y2=0
cc_1003 N_A_2511_137#_c_1632_n N_VPWR_c_1686_n 0.002179f $X=13.365 $Y=1.47 $X2=0
+ $Y2=0
cc_1004 N_A_2511_137#_M1016_g N_VPWR_c_1697_n 0.00549284f $X=13.425 $Y=2.465
+ $X2=0 $Y2=0
cc_1005 N_A_2511_137#_M1016_g N_VPWR_c_1677_n 0.0120439f $X=13.425 $Y=2.465
+ $X2=0 $Y2=0
cc_1006 N_A_2511_137#_c_1635_n N_VPWR_c_1677_n 0.00972751f $X=12.7 $Y=1.98 $X2=0
+ $Y2=0
cc_1007 N_A_2511_137#_c_1630_n N_Q_N_c_1872_n 0.0484357f $X=12.7 $Y=0.895 $X2=0
+ $Y2=0
cc_1008 N_A_2511_137#_c_1635_n N_Q_N_c_1874_n 0.06692f $X=12.7 $Y=1.98 $X2=0
+ $Y2=0
cc_1009 N_A_2511_137#_c_1633_n N_Q_N_c_1874_n 0.0265131f $X=12.74 $Y=1.47 $X2=0
+ $Y2=0
cc_1010 N_A_2511_137#_M1016_g N_Q_c_1910_n 0.0145249f $X=13.425 $Y=2.465 $X2=0
+ $Y2=0
cc_1011 N_A_2511_137#_M1016_g N_Q_c_1911_n 0.00349143f $X=13.425 $Y=2.465 $X2=0
+ $Y2=0
cc_1012 N_A_2511_137#_c_1632_n N_Q_c_1911_n 0.00131892f $X=13.365 $Y=1.47 $X2=0
+ $Y2=0
cc_1013 N_A_2511_137#_M1035_g N_Q_c_1907_n 0.00448208f $X=13.425 $Y=0.685 $X2=0
+ $Y2=0
cc_1014 N_A_2511_137#_M1016_g N_Q_c_1907_n 0.00448208f $X=13.425 $Y=2.465 $X2=0
+ $Y2=0
cc_1015 N_A_2511_137#_c_1631_n N_Q_c_1907_n 0.0250952f $X=13.365 $Y=1.47 $X2=0
+ $Y2=0
cc_1016 N_A_2511_137#_c_1632_n N_Q_c_1907_n 0.00782465f $X=13.365 $Y=1.47 $X2=0
+ $Y2=0
cc_1017 N_A_2511_137#_M1035_g Q 0.00349143f $X=13.425 $Y=0.685 $X2=0 $Y2=0
cc_1018 N_A_2511_137#_c_1632_n Q 0.00131892f $X=13.365 $Y=1.47 $X2=0 $Y2=0
cc_1019 N_A_2511_137#_M1035_g N_Q_c_1909_n 0.010351f $X=13.425 $Y=0.685 $X2=0
+ $Y2=0
cc_1020 N_A_2511_137#_M1035_g N_VGND_c_1937_n 0.0055345f $X=13.425 $Y=0.685
+ $X2=0 $Y2=0
cc_1021 N_A_2511_137#_c_1630_n N_VGND_c_1937_n 0.0172562f $X=12.7 $Y=0.895 $X2=0
+ $Y2=0
cc_1022 N_A_2511_137#_c_1631_n N_VGND_c_1937_n 0.0206753f $X=13.365 $Y=1.47
+ $X2=0 $Y2=0
cc_1023 N_A_2511_137#_c_1632_n N_VGND_c_1937_n 0.002179f $X=13.365 $Y=1.47 $X2=0
+ $Y2=0
cc_1024 N_A_2511_137#_c_1630_n N_VGND_c_1945_n 0.00467036f $X=12.7 $Y=0.895
+ $X2=0 $Y2=0
cc_1025 N_A_2511_137#_M1035_g N_VGND_c_1946_n 0.00520813f $X=13.425 $Y=0.685
+ $X2=0 $Y2=0
cc_1026 N_A_2511_137#_M1035_g N_VGND_c_1947_n 0.0115451f $X=13.425 $Y=0.685
+ $X2=0 $Y2=0
cc_1027 N_A_2511_137#_c_1630_n N_VGND_c_1947_n 0.00733137f $X=12.7 $Y=0.895
+ $X2=0 $Y2=0
cc_1028 N_VPWR_c_1680_n N_A_460_449#_c_1824_n 0.0240212f $X=1.88 $Y=2.39 $X2=0
+ $Y2=0
cc_1029 N_VPWR_c_1689_n N_A_460_449#_c_1824_n 0.006147f $X=4.605 $Y=3.33 $X2=0
+ $Y2=0
cc_1030 N_VPWR_c_1677_n N_A_460_449#_c_1824_n 0.0182625f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1031 N_VPWR_c_1677_n A_2036_451# 0.00899413f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1032 N_VPWR_c_1685_n Q_N 0.0165395f $X=11.73 $Y=2.775 $X2=0 $Y2=0
cc_1033 N_VPWR_c_1686_n Q_N 0.0168408f $X=13.21 $Y=1.98 $X2=0 $Y2=0
cc_1034 N_VPWR_c_1696_n Q_N 0.0169956f $X=13.045 $Y=3.33 $X2=0 $Y2=0
cc_1035 N_VPWR_c_1677_n Q_N 0.0133402f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1036 N_VPWR_c_1677_n N_Q_M1016_d 0.0023218f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1037 N_VPWR_c_1697_n N_Q_c_1910_n 0.0214436f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1038 N_VPWR_c_1677_n N_Q_c_1910_n 0.0134754f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1039 N_VPWR_c_1686_n N_Q_c_1911_n 0.045997f $X=13.21 $Y=1.98 $X2=0 $Y2=0
cc_1040 N_A_460_449#_c_1820_n N_VGND_c_1932_n 0.01467f $X=2.575 $Y=0.805 $X2=0
+ $Y2=0
cc_1041 N_A_460_449#_c_1820_n N_VGND_c_1938_n 0.00743798f $X=2.575 $Y=0.805
+ $X2=0 $Y2=0
cc_1042 N_A_460_449#_c_1820_n N_VGND_c_1947_n 0.00904485f $X=2.575 $Y=0.805
+ $X2=0 $Y2=0
cc_1043 N_Q_N_c_1872_n N_VGND_c_1937_n 0.0137265f $X=12.14 $Y=0.43 $X2=0 $Y2=0
cc_1044 N_Q_N_c_1872_n N_VGND_c_1945_n 0.0285232f $X=12.14 $Y=0.43 $X2=0 $Y2=0
cc_1045 N_Q_N_M1030_d N_VGND_c_1947_n 0.0023218f $X=12 $Y=0.235 $X2=0 $Y2=0
cc_1046 N_Q_N_c_1872_n N_VGND_c_1947_n 0.0175381f $X=12.14 $Y=0.43 $X2=0 $Y2=0
cc_1047 N_Q_c_1909_n N_VGND_c_1937_n 0.0318617f $X=13.64 $Y=0.43 $X2=0 $Y2=0
cc_1048 N_Q_c_1909_n N_VGND_c_1946_n 0.0214436f $X=13.64 $Y=0.43 $X2=0 $Y2=0
cc_1049 N_Q_c_1909_n N_VGND_c_1947_n 0.0135379f $X=13.64 $Y=0.43 $X2=0 $Y2=0
cc_1050 N_VGND_c_1935_n N_A_1896_119#_c_2086_n 0.0256141f $X=9.11 $Y=0.77 $X2=0
+ $Y2=0
cc_1051 N_VGND_c_1944_n N_A_1896_119#_c_2087_n 0.0413713f $X=11.545 $Y=0 $X2=0
+ $Y2=0
cc_1052 N_VGND_c_1947_n N_A_1896_119#_c_2087_n 0.023033f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1053 N_VGND_c_1935_n N_A_1896_119#_c_2088_n 0.0144411f $X=9.11 $Y=0.77 $X2=0
+ $Y2=0
cc_1054 N_VGND_c_1944_n N_A_1896_119#_c_2088_n 0.0223013f $X=11.545 $Y=0 $X2=0
+ $Y2=0
cc_1055 N_VGND_c_1947_n N_A_1896_119#_c_2088_n 0.0114651f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1056 N_VGND_c_1944_n N_A_1896_119#_c_2089_n 0.0212031f $X=11.545 $Y=0 $X2=0
+ $Y2=0
cc_1057 N_VGND_c_1947_n N_A_1896_119#_c_2089_n 0.0125042f $X=13.68 $Y=0 $X2=0
+ $Y2=0
