* File: sky130_fd_sc_lp__sdfrbp_2.spice
* Created: Wed Sep  2 10:34:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfrbp_2.pex.spice"
.subckt sky130_fd_sc_lp__sdfrbp_2  VNB VPB SCE D SCD CLK RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_SCE_M1014_g N_A_27_81#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1033 noxref_26 N_A_27_81#_M1033_g N_noxref_25_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1035 N_A_359_489#_M1035_d N_D_M1035_g noxref_26 VNB NSHORT L=0.15 W=0.42
+ AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=7.14 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1024 noxref_27 N_SCE_M1024_g N_A_359_489#_M1035_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.06405 PD=0.715 PS=0.725 NRD=26.424 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1047 N_noxref_25_M1047_d N_SCD_M1047_g noxref_27 VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.06195 PD=0.7 PS=0.715 NRD=0 NRS=26.424 M=1 R=2.8 SA=75001.4
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_RESET_B_M1015_g N_noxref_25_M1047_d VNB NSHORT L=0.15
+ W=0.42 AD=0.08945 AS=0.0588 PD=0.95 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1019 N_A_759_119#_M1019_d N_CLK_M1019_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.08945 PD=0.7 PS=0.95 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1022 N_A_759_119#_M1019_d N_CLK_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.103375 PD=0.7 PS=0.975 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_934_367#_M1013_d N_A_759_119#_M1013_g N_VGND_M1022_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.103375 PD=0.7 PS=0.975 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75002.4 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1027 N_A_934_367#_M1013_d N_A_759_119#_M1027_g N_VGND_M1027_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1043 N_A_1162_463#_M1043_d N_A_759_119#_M1043_g N_A_359_489#_M1043_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1028 A_1349_119# N_A_934_367#_M1028_g N_A_1162_463#_M1043_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1036 A_1421_119# N_A_1290_365#_M1036_g A_1349_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_RESET_B_M1025_g A_1421_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.136104 AS=0.0441 PD=0.978679 PS=0.63 NRD=76.872 NRS=14.28 M=1 R=2.8
+ SA=75001.3 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_1290_365#_M1005_d N_A_1162_463#_M1005_g N_VGND_M1025_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.23415 AS=0.207396 PD=1.51 PS=1.49132 NRD=58.284 NRS=23.436
+ M=1 R=4.26667 SA=75001.4 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1046 N_A_1770_412#_M1046_d N_A_934_367#_M1046_g N_A_1290_365#_M1005_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.125283 AS=0.23415 PD=1.19547 PS=1.51 NRD=13.116
+ NRS=58.284 M=1 R=4.26667 SA=75002.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1040 A_1879_68# N_A_759_119#_M1040_g N_A_1770_412#_M1046_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.082217 PD=0.78 PS=0.784528 NRD=35.712 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1044 N_VGND_M1044_d N_A_1923_174#_M1044_g A_1879_68# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=35.712 M=1 R=2.8 SA=75002.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1016 A_2067_68# N_RESET_B_M1016_g N_VGND_M1044_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_A_1923_174#_M1020_d N_A_1770_412#_M1020_g A_2067_68# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_1770_412#_M1003_g N_Q_N_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1037 N_VGND_M1037_d N_A_1770_412#_M1037_g N_Q_N_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1792 AS=0.1176 PD=1.62 PS=1.12 NRD=6.78 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.5 A=0.126 P=1.98 MULT=1
MM1011 N_A_2516_367#_M1011_d N_A_1770_412#_M1011_g N_VGND_M1037_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0896 PD=1.37 PS=0.81 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_2516_367#_M1006_g N_Q_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1030 N_VGND_M1030_d N_A_2516_367#_M1030_g N_Q_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_VPWR_M1021_d N_SCE_M1021_g N_A_27_81#_M1021_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1004 A_287_489# N_SCE_M1004_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1009 N_A_359_489#_M1009_d N_D_M1009_g A_287_489# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1041 A_445_489# N_A_27_81#_M1041_g N_A_359_489#_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=32.308 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1034 N_VPWR_M1034_d N_SCD_M1034_g A_445_489# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.1024 PD=1.03 PS=0.96 NRD=0 NRS=32.308 M=1 R=4.26667 SA=75001.9
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_359_489#_M1002_d N_RESET_B_M1002_g N_VPWR_M1034_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1248 PD=1.81 PS=1.03 NRD=0 NRS=33.8446 M=1 R=4.26667
+ SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1042 N_VPWR_M1042_d N_CLK_M1042_g N_A_759_119#_M1042_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_A_934_367#_M1017_d N_A_759_119#_M1017_g N_VPWR_M1042_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1038 N_A_1162_463#_M1038_d N_A_934_367#_M1038_g N_A_359_489#_M1038_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1218 PD=0.7 PS=1.42 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1023 A_1248_463# N_A_759_119#_M1023_g N_A_1162_463#_M1038_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_1290_365#_M1000_g A_1248_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1395 AS=0.0441 PD=1.11 PS=0.63 NRD=56.2829 NRS=23.443 M=1 R=2.8
+ SA=75001 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1018 N_A_1162_463#_M1018_d N_RESET_B_M1018_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1395 PD=1.37 PS=1.11 NRD=0 NRS=129.981 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_A_1290_365#_M1031_d N_A_1162_463#_M1031_g N_VPWR_M1031_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.192937 AS=0.2604 PD=1.43 PS=2.3 NRD=8.1952 NRS=10.5395 M=1
+ R=5.6 SA=75000.2 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1010 N_A_1770_412#_M1010_d N_A_759_119#_M1010_g N_A_1290_365#_M1031_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1932 AS=0.192937 PD=1.68667 PS=1.43 NRD=0
+ NRS=25.7873 M=1 R=5.6 SA=75000.7 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1032 A_1885_496# N_A_934_367#_M1032_g N_A_1770_412#_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0966 PD=0.81 PS=0.843333 NRD=65.6601 NRS=68.0044 M=1
+ R=2.8 SA=75001.2 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_1923_174#_M1001_g A_1885_496# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09975 AS=0.0819 PD=0.895 PS=0.81 NRD=39.8531 NRS=65.6601 M=1 R=2.8
+ SA=75001.7 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1012 N_A_1923_174#_M1012_d N_RESET_B_M1012_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.09975 PD=0.7 PS=0.895 NRD=0 NRS=51.5943 M=1 R=2.8
+ SA=75002.3 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1045 N_VPWR_M1045_d N_A_1770_412#_M1045_g N_A_1923_174#_M1012_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.111825 AS=0.0588 PD=0.8575 PS=0.7 NRD=99.0713 NRS=0 M=1
+ R=2.8 SA=75002.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1007 N_Q_N_M1007_d N_A_1770_412#_M1007_g N_VPWR_M1045_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.335475 PD=1.54 PS=2.5725 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75001.3 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1039 N_Q_N_M1007_d N_A_1770_412#_M1039_g N_VPWR_M1039_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.268115 PD=1.54 PS=2.16853 NRD=0 NRS=2.3443 M=1 R=8.4
+ SA=75001.7 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1029 N_A_2516_367#_M1029_d N_A_1770_412#_M1029_g N_VPWR_M1039_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.136185 PD=1.81 PS=1.10147 NRD=0 NRS=23.0687 M=1
+ R=4.26667 SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A_2516_367#_M1008_g N_Q_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1026_d N_A_2516_367#_M1026_g N_Q_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX48_noxref VNB VPB NWDIODE A=27.5647 P=33.29
c_150 VNB 0 8.72856e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__sdfrbp_2.pxi.spice"
*
.ends
*
*
