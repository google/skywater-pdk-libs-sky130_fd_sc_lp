* File: sky130_fd_sc_lp__maj3_lp.pex.spice
* Created: Wed Sep  2 09:59:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MAJ3_LP%A 3 7 11 15 17 18 26
r52 26 27 7.32523 $w=3.29e-07 $l=5e-08 $layer=POLY_cond $X=1.625 $Y=1.77
+ $X2=1.675 $Y2=1.77
r53 24 26 5.86018 $w=3.29e-07 $l=4e-08 $layer=POLY_cond $X=1.585 $Y=1.77
+ $X2=1.625 $Y2=1.77
r54 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=1.77 $X2=1.585 $Y2=1.77
r55 22 24 71.7872 $w=3.29e-07 $l=4.9e-07 $layer=POLY_cond $X=1.095 $Y=1.77
+ $X2=1.585 $Y2=1.77
r56 21 22 1.46505 $w=3.29e-07 $l=1e-08 $layer=POLY_cond $X=1.085 $Y=1.77
+ $X2=1.095 $Y2=1.77
r57 18 25 2.08491 $w=5.43e-07 $l=9.5e-08 $layer=LI1_cond $X=1.68 $Y=1.877
+ $X2=1.585 $Y2=1.877
r58 17 25 8.44936 $w=5.43e-07 $l=3.85e-07 $layer=LI1_cond $X=1.2 $Y=1.877
+ $X2=1.585 $Y2=1.877
r59 13 27 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.605
+ $X2=1.675 $Y2=1.77
r60 13 15 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.675 $Y=1.605
+ $X2=1.675 $Y2=0.835
r61 9 26 9.27491 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=1.935
+ $X2=1.625 $Y2=1.77
r62 9 11 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.625 $Y=1.935
+ $X2=1.625 $Y2=2.595
r63 5 21 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.605
+ $X2=1.085 $Y2=1.77
r64 5 7 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.085 $Y=1.605
+ $X2=1.085 $Y2=0.835
r65 1 22 9.27491 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.935
+ $X2=1.095 $Y2=1.77
r66 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.095 $Y=1.935
+ $X2=1.095 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_LP%B 3 8 9 10 13 15 17 20 22 27 31 32 35 36 37
+ 44 46
c98 13 0 2.67377e-20 $X=2.615 $Y=2.595
r99 37 46 6.54083 $w=2.33e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.297
+ $X2=1.315 $Y2=1.297
r100 37 44 6.0959 $w=2.33e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.297
+ $X2=1.085 $Y2=1.297
r101 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.595
+ $Y=1.39 $X2=0.595 $Y2=1.39
r102 32 42 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=1.75
+ $X2=2.585 $Y2=1.915
r103 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=1.75 $X2=2.585 $Y2=1.75
r104 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.585 $Y=1.415
+ $X2=2.585 $Y2=1.75
r105 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.42 $Y=1.33
+ $X2=2.585 $Y2=1.415
r106 27 46 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.42 $Y=1.33
+ $X2=1.315 $Y2=1.33
r107 26 35 4.64874 $w=1.9e-07 $l=1.6e-07 $layer=LI1_cond $X=0.76 $Y=1.32 $X2=0.6
+ $Y2=1.32
r108 26 44 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=0.76 $Y=1.32
+ $X2=1.085 $Y2=1.32
r109 21 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.595 $Y=1.73
+ $X2=0.595 $Y2=1.39
r110 21 22 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.73
+ $X2=0.595 $Y2=1.895
r111 20 36 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.595 $Y=1.375
+ $X2=0.595 $Y2=1.39
r112 19 20 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.6 $Y=1.225
+ $X2=0.6 $Y2=1.375
r113 15 17 94.7933 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.575 $Y=0.255
+ $X2=2.575 $Y2=0.55
r114 13 42 168.948 $w=2.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.615 $Y=2.595
+ $X2=2.615 $Y2=1.915
r115 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.5 $Y=0.18
+ $X2=2.575 $Y2=0.255
r116 9 10 887.085 $w=1.5e-07 $l=1.73e-06 $layer=POLY_cond $X=2.5 $Y=0.18
+ $X2=0.77 $Y2=0.18
r117 8 19 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=0.695 $Y=0.835
+ $X2=0.695 $Y2=1.225
r118 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.695 $Y=0.255
+ $X2=0.77 $Y2=0.18
r119 5 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.695 $Y=0.255
+ $X2=0.695 $Y2=0.835
r120 3 22 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.635 $Y=2.595
+ $X2=0.635 $Y2=1.895
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_LP%C 3 7 9 13 17 19 21 23 24 27 28
r71 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.125
+ $Y=1.41 $X2=3.125 $Y2=1.41
r72 24 28 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.125 $Y=1.665
+ $X2=3.125 $Y2=1.41
r73 22 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.125 $Y=1.75
+ $X2=3.125 $Y2=1.41
r74 22 23 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.75
+ $X2=3.125 $Y2=1.915
r75 20 27 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.125 $Y=1.375
+ $X2=3.125 $Y2=1.41
r76 20 21 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=3.125 $Y=1.375
+ $X2=3.125 $Y2=1.3
r77 17 23 168.948 $w=2.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.115 $Y=2.595
+ $X2=3.115 $Y2=1.915
r78 11 21 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.035 $Y=1.225
+ $X2=3.125 $Y2=1.3
r79 11 13 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.035 $Y=1.225
+ $X2=3.035 $Y2=0.55
r80 10 19 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.21 $Y=1.3
+ $X2=2.085 $Y2=1.3
r81 9 21 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.96 $Y=1.3
+ $X2=3.125 $Y2=1.3
r82 9 10 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.96 $Y=1.3 $X2=2.21
+ $Y2=1.3
r83 5 19 15.9654 $w=2e-07 $l=8.44097e-08 $layer=POLY_cond $X=2.065 $Y=1.225
+ $X2=2.085 $Y2=1.3
r84 5 7 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.065 $Y=1.225
+ $X2=2.065 $Y2=0.835
r85 1 19 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=2.085 $Y=1.375
+ $X2=2.085 $Y2=1.3
r86 1 3 303.113 $w=2.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.085 $Y=1.375
+ $X2=2.085 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_LP%A_29_419# 1 2 3 4 13 15 18 20 22 27 30 35 37
+ 40 41 47 49 53 54 60 61 63 64 66 68 69
c135 37 0 2.67377e-20 $X=2.185 $Y=2.415
r136 66 68 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.35 $Y=2.26
+ $X2=2.35 $Y2=2.415
r137 63 64 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=1.495 $Y=0.947
+ $X2=1.665 $Y2=0.947
r138 60 62 5.52541 $w=3.63e-07 $l=1.75e-07 $layer=LI1_cond $X=0.272 $Y=2.24
+ $X2=0.272 $Y2=2.415
r139 60 61 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=2.24
+ $X2=0.272 $Y2=2.075
r140 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.695
+ $Y=1.15 $X2=3.695 $Y2=1.15
r141 51 53 2.92411 $w=3.33e-07 $l=8.5e-08 $layer=LI1_cond $X=3.692 $Y=1.065
+ $X2=3.692 $Y2=1.15
r142 50 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=0.98
+ $X2=2.36 $Y2=0.98
r143 49 51 20.8151 $w=9.4e-08 $l=2.05144e-07 $layer=LI1_cond $X=3.525 $Y=0.98
+ $X2=3.692 $Y2=1.065
r144 49 50 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.525 $Y=0.98
+ $X2=2.525 $Y2=0.98
r145 45 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.895
+ $X2=2.36 $Y2=0.98
r146 45 47 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.36 $Y=0.895
+ $X2=2.36 $Y2=0.55
r147 41 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0.98
+ $X2=2.36 $Y2=0.98
r148 41 64 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.195 $Y=0.98
+ $X2=1.665 $Y2=0.98
r149 40 58 8.95823 $w=3.3e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.645 $Y=0.915
+ $X2=0.48 $Y2=0.825
r150 40 63 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.645 $Y=0.915
+ $X2=1.495 $Y2=0.915
r151 38 62 5.2253 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.455 $Y=2.415
+ $X2=0.272 $Y2=2.415
r152 37 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=2.415
+ $X2=2.35 $Y2=2.415
r153 37 38 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=2.185 $Y=2.415
+ $X2=0.455 $Y2=2.415
r154 33 62 2.68377 $w=3.63e-07 $l=8.5e-08 $layer=LI1_cond $X=0.272 $Y=2.5
+ $X2=0.272 $Y2=2.415
r155 33 35 12.6295 $w=3.63e-07 $l=4e-07 $layer=LI1_cond $X=0.272 $Y=2.5
+ $X2=0.272 $Y2=2.9
r156 31 58 11.2758 $w=3.3e-07 $l=4.00156e-07 $layer=LI1_cond $X=0.175 $Y=1.045
+ $X2=0.48 $Y2=0.825
r157 31 61 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.175 $Y=1.045
+ $X2=0.175 $Y2=2.075
r158 29 54 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.695 $Y=1.49
+ $X2=3.695 $Y2=1.15
r159 29 30 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.49
+ $X2=3.695 $Y2=1.655
r160 26 54 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=0.985
+ $X2=3.695 $Y2=1.15
r161 26 27 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=3.695 $Y=0.91
+ $X2=3.825 $Y2=0.91
r162 23 26 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.465 $Y=0.91
+ $X2=3.695 $Y2=0.91
r163 20 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.825 $Y=0.835
+ $X2=3.825 $Y2=0.91
r164 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.825 $Y=0.835
+ $X2=3.825 $Y2=0.55
r165 18 30 233.546 $w=2.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.655 $Y=2.595
+ $X2=3.655 $Y2=1.655
r166 13 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.465 $Y=0.835
+ $X2=3.465 $Y2=0.91
r167 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.465 $Y=0.835
+ $X2=3.465 $Y2=0.55
r168 4 66 300 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=2 $X=2.21
+ $Y=2.095 $X2=2.35 $Y2=2.26
r169 3 60 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=2.095 $X2=0.29 $Y2=2.24
r170 3 35 600 $w=1.7e-07 $l=8.745e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=2.095 $X2=0.29 $Y2=2.9
r171 2 47 182 $w=1.7e-07 $l=2.54755e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.625 $X2=2.36 $Y2=0.55
r172 1 58 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.335
+ $Y=0.625 $X2=0.48 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_LP%VPWR 1 2 9 13 18 19 20 22 35 36 39
r50 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 29 32 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.36 $Y2=3.33
r58 27 29 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 25 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.36 $Y2=3.33
r62 22 24 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 20 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r64 20 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 18 32 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.215 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=3.33
+ $X2=3.38 $Y2=3.33
r67 17 35 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=4.08 $Y2=3.33
r68 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=3.38 $Y2=3.33
r69 13 16 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.38 $Y=2.26
+ $X2=3.38 $Y2=2.95
r70 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.38 $Y=3.245
+ $X2=3.38 $Y2=3.33
r71 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.38 $Y=3.245
+ $X2=3.38 $Y2=2.95
r72 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=3.245 $X2=1.36
+ $Y2=3.33
r73 7 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.36 $Y=3.245 $X2=1.36
+ $Y2=2.895
r74 2 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=2.095 $X2=3.38 $Y2=2.95
r75 2 13 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=2.095 $X2=3.38 $Y2=2.26
r76 1 9 600 $w=1.7e-07 $l=8.67179e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=2.095 $X2=1.36 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_LP%X 1 2 10 13 14 15 21 28
r24 19 21 2.44473 $w=4.53e-07 $l=9.3e-08 $layer=LI1_cond $X=3.982 $Y=2.147
+ $X2=3.982 $Y2=2.24
r25 14 15 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.982 $Y=2.405
+ $X2=3.982 $Y2=2.775
r26 14 21 4.33743 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.982 $Y=2.405
+ $X2=3.982 $Y2=2.24
r27 13 19 2.94419 $w=4.53e-07 $l=1.12e-07 $layer=LI1_cond $X=3.982 $Y=2.035
+ $X2=3.982 $Y2=2.147
r28 13 28 7.93754 $w=4.53e-07 $l=1.15e-07 $layer=LI1_cond $X=3.982 $Y=2.035
+ $X2=3.982 $Y2=1.92
r29 12 28 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=4.125 $Y=0.78
+ $X2=4.125 $Y2=1.92
r30 10 12 10.7022 $w=3.33e-07 $l=2.3e-07 $layer=LI1_cond $X=4.042 $Y=0.55
+ $X2=4.042 $Y2=0.78
r31 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.78
+ $Y=2.095 $X2=3.92 $Y2=2.24
r32 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.34 $X2=4.04 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_LP%VGND 1 2 9 13 16 17 18 27 33 34 37
r46 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 34 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r48 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r49 31 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.25
+ $Y2=0
r50 31 33 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=4.08
+ $Y2=0
r51 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 27 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.25
+ $Y2=0
r53 27 29 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=3.085 $Y=0
+ $X2=1.68 $Y2=0
r54 26 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r55 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r56 22 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r57 21 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r58 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 18 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r60 18 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r61 16 25 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.215 $Y=0 $X2=1.2
+ $Y2=0
r62 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=0 $X2=1.38
+ $Y2=0
r63 15 29 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.68
+ $Y2=0
r64 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.38
+ $Y2=0
r65 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0
r66 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0.515
r67 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=0.085 $X2=1.38
+ $Y2=0
r68 7 9 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=1.38 $Y=0.085 $X2=1.38
+ $Y2=0.485
r69 2 13 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3.11
+ $Y=0.34 $X2=3.25 $Y2=0.515
r70 1 9 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.625 $X2=1.38 $Y2=0.485
.ends

