# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o31a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o31a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.375000 1.210000 6.095000 1.535000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.850000 1.345000 5.205000 1.705000 ;
        RECT 4.850000 1.705000 6.595000 1.750000 ;
        RECT 4.920000 1.750000 6.595000 1.875000 ;
        RECT 6.265000 1.295000 6.595000 1.705000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.425000 4.680000 1.750000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.425000 3.335000 2.120000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 1.750000 1.225000 ;
        RECT 0.085000 1.225000 0.335000 1.755000 ;
        RECT 0.085000 1.755000 1.975000 1.925000 ;
        RECT 0.700000 0.255000 0.890000 1.055000 ;
        RECT 0.925000 1.925000 1.115000 3.075000 ;
        RECT 1.560000 0.255000 1.750000 1.055000 ;
        RECT 1.795000 1.925000 1.975000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.200000  0.085000 0.530000 0.885000 ;
      RECT 0.425000  2.095000 0.755000 3.245000 ;
      RECT 0.505000  1.405000 2.835000 1.575000 ;
      RECT 1.060000  0.085000 1.390000 0.885000 ;
      RECT 1.285000  2.095000 1.615000 3.245000 ;
      RECT 1.920000  0.085000 2.250000 1.105000 ;
      RECT 2.145000  1.815000 2.475000 3.245000 ;
      RECT 2.620000  0.255000 3.820000 0.435000 ;
      RECT 2.620000  0.435000 2.950000 0.905000 ;
      RECT 2.635000  1.075000 3.460000 1.245000 ;
      RECT 2.635000  1.245000 2.835000 1.405000 ;
      RECT 2.645000  1.575000 2.835000 2.290000 ;
      RECT 2.645000  2.290000 4.260000 2.460000 ;
      RECT 2.645000  2.460000 2.825000 3.075000 ;
      RECT 3.005000  2.630000 3.335000 3.245000 ;
      RECT 3.130000  0.605000 3.460000 1.075000 ;
      RECT 3.560000  1.920000 4.750000 2.045000 ;
      RECT 3.560000  2.045000 6.625000 2.120000 ;
      RECT 3.630000  0.435000 3.820000 1.075000 ;
      RECT 3.630000  1.075000 4.710000 1.245000 ;
      RECT 3.990000  0.085000 4.320000 0.895000 ;
      RECT 3.990000  2.460000 4.260000 3.075000 ;
      RECT 4.430000  2.120000 6.625000 2.265000 ;
      RECT 4.430000  2.265000 4.750000 3.075000 ;
      RECT 4.490000  0.305000 4.750000 0.870000 ;
      RECT 4.490000  0.870000 6.625000 1.040000 ;
      RECT 4.490000  1.040000 4.710000 1.075000 ;
      RECT 4.925000  0.085000 5.255000 0.700000 ;
      RECT 4.925000  2.435000 5.255000 2.835000 ;
      RECT 4.925000  2.835000 6.195000 3.075000 ;
      RECT 5.425000  2.435000 6.625000 2.665000 ;
      RECT 5.435000  0.305000 5.695000 0.870000 ;
      RECT 5.865000  0.085000 6.195000 0.700000 ;
      RECT 6.365000  0.305000 6.625000 0.870000 ;
      RECT 6.365000  2.665000 6.625000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__o31a_4
END LIBRARY
