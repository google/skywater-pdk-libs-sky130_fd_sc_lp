* File: sky130_fd_sc_lp__mux2i_lp2.pxi.spice
* Created: Wed Sep  2 10:01:24 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2I_LP2%S N_S_M1006_g N_S_c_72_n N_S_c_73_n N_S_M1005_g
+ N_S_c_75_n N_S_M1000_g N_S_c_76_n N_S_M1003_g N_S_c_78_n N_S_M1009_g
+ N_S_c_79_n N_S_c_80_n N_S_c_81_n N_S_c_82_n N_S_c_83_n N_S_c_84_n S N_S_c_85_n
+ N_S_c_86_n PM_SKY130_FD_SC_LP__MUX2I_LP2%S
x_PM_SKY130_FD_SC_LP__MUX2I_LP2%A0 N_A0_M1007_g N_A0_M1010_g N_A0_c_185_n
+ N_A0_c_186_n N_A0_c_187_n N_A0_c_188_n A0 N_A0_c_189_n
+ PM_SKY130_FD_SC_LP__MUX2I_LP2%A0
x_PM_SKY130_FD_SC_LP__MUX2I_LP2%A1 N_A1_M1004_g N_A1_M1008_g A1 N_A1_c_249_n
+ N_A1_c_250_n PM_SKY130_FD_SC_LP__MUX2I_LP2%A1
x_PM_SKY130_FD_SC_LP__MUX2I_LP2%A_490_21# N_A_490_21#_M1009_d
+ N_A_490_21#_M1003_d N_A_490_21#_M1002_g N_A_490_21#_M1001_g
+ N_A_490_21#_c_292_n N_A_490_21#_c_293_n N_A_490_21#_c_294_n
+ N_A_490_21#_c_295_n N_A_490_21#_c_302_n N_A_490_21#_c_296_n
+ N_A_490_21#_c_297_n N_A_490_21#_c_298_n
+ PM_SKY130_FD_SC_LP__MUX2I_LP2%A_490_21#
x_PM_SKY130_FD_SC_LP__MUX2I_LP2%VPWR N_VPWR_M1006_s N_VPWR_M1001_d
+ N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n N_VPWR_c_361_n
+ VPWR N_VPWR_c_362_n N_VPWR_c_356_n PM_SKY130_FD_SC_LP__MUX2I_LP2%VPWR
x_PM_SKY130_FD_SC_LP__MUX2I_LP2%Y N_Y_M1004_d N_Y_M1007_d N_Y_c_401_n
+ N_Y_c_402_n N_Y_c_403_n N_Y_c_406_n N_Y_c_407_n N_Y_c_404_n N_Y_c_468_p
+ N_Y_c_425_n N_Y_c_445_n N_Y_c_430_n N_Y_c_437_n Y Y N_Y_c_408_n Y
+ PM_SKY130_FD_SC_LP__MUX2I_LP2%Y
x_PM_SKY130_FD_SC_LP__MUX2I_LP2%VGND N_VGND_M1005_s N_VGND_M1002_d
+ N_VGND_c_487_n N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n VGND
+ N_VGND_c_491_n N_VGND_c_492_n N_VGND_c_493_n N_VGND_c_494_n
+ PM_SKY130_FD_SC_LP__MUX2I_LP2%VGND
cc_1 VNB N_S_c_72_n 0.02783f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.15
cc_2 VNB N_S_c_73_n 0.0189524f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.15
cc_3 VNB N_S_M1005_g 0.0386251f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.445
cc_4 VNB N_S_c_75_n 0.015126f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=0.765
cc_5 VNB N_S_c_76_n 0.053738f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=1.28
cc_6 VNB N_S_M1003_g 0.0253179f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.595
cc_7 VNB N_S_c_78_n 0.0192926f $X=-0.19 $Y=-0.245 $X2=3.33 $Y2=0.765
cc_8 VNB N_S_c_79_n 0.00569476f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.745
cc_9 VNB N_S_c_80_n 0.0111557f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.16
cc_10 VNB N_S_c_81_n 0.00173406f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.075
cc_11 VNB N_S_c_82_n 8.77584e-19 $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.8
cc_12 VNB N_S_c_83_n 0.00475825f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.24
cc_13 VNB N_S_c_84_n 0.0346434f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.24
cc_14 VNB N_S_c_85_n 0.00871636f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=0.93
cc_15 VNB N_S_c_86_n 0.0222552f $X=-0.19 $Y=-0.245 $X2=2.525 $Y2=0.905
cc_16 VNB N_A0_M1010_g 0.0324788f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.075
cc_17 VNB N_A0_c_185_n 0.00845209f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.445
cc_18 VNB N_A0_c_186_n 0.00767059f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=0.765
cc_19 VNB N_A0_c_187_n 0.0290467f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=0.445
cc_20 VNB N_A0_c_188_n 0.00419156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A0_c_189_n 0.0166974f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.58
cc_22 VNB N_A1_M1004_g 0.0636929f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.595
cc_23 VNB N_A1_c_249_n 0.0144903f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=0.445
cc_24 VNB N_A1_c_250_n 0.003868f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.595
cc_25 VNB N_A_490_21#_c_292_n 0.014996f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.595
cc_26 VNB N_A_490_21#_c_293_n 0.00870458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_490_21#_c_294_n 0.0112412f $X=-0.19 $Y=-0.245 $X2=3.33 $Y2=0.765
cc_28 VNB N_A_490_21#_c_295_n 0.0269215f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.225
cc_29 VNB N_A_490_21#_c_296_n 0.0480436f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.075
cc_30 VNB N_A_490_21#_c_297_n 0.0168844f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.8
cc_31 VNB N_A_490_21#_c_298_n 0.0241736f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.24
cc_32 VNB N_VPWR_c_356_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.8
cc_33 VNB N_Y_c_401_n 0.0404991f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.445
cc_34 VNB N_Y_c_402_n 0.0222511f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.445
cc_35 VNB N_Y_c_403_n 0.0104961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_404_n 0.00322783f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=1.28
cc_37 VNB N_VGND_c_487_n 0.0173524f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.445
cc_38 VNB N_VGND_c_488_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=0.445
cc_39 VNB N_VGND_c_489_n 0.012318f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.595
cc_40 VNB N_VGND_c_490_n 0.006319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_491_n 0.0461021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_492_n 0.0265702f $X=-0.19 $Y=-0.245 $X2=2.525 $Y2=0.8
cc_43 VNB N_VGND_c_493_n 0.212473f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.8
cc_44 VNB N_VGND_c_494_n 0.00436557f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.24
cc_45 VPB N_S_M1006_g 0.0415053f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.595
cc_46 VPB N_S_M1003_g 0.0516649f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=2.595
cc_47 VPB N_S_c_79_n 0.00906011f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.745
cc_48 VPB N_S_c_83_n 7.46168e-19 $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.24
cc_49 VPB N_A0_M1007_g 0.0382448f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.595
cc_50 VPB N_A0_c_185_n 0.00290646f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=0.445
cc_51 VPB N_A0_c_188_n 0.0090307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A0_c_189_n 0.0102922f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.58
cc_53 VPB N_A1_M1008_g 0.0290761f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=1.075
cc_54 VPB N_A1_c_249_n 0.0389121f $X=-0.19 $Y=1.655 $X2=2.97 $Y2=0.445
cc_55 VPB N_A1_c_250_n 0.00467449f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=2.595
cc_56 VPB N_A_490_21#_M1001_g 0.0450227f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=1.28
cc_57 VPB N_A_490_21#_c_294_n 0.00364207f $X=-0.19 $Y=1.655 $X2=3.33 $Y2=0.765
cc_58 VPB N_A_490_21#_c_295_n 0.00285041f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.225
cc_59 VPB N_A_490_21#_c_302_n 0.0629326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_490_21#_c_297_n 4.92344e-19 $X=-0.19 $Y=1.655 $X2=1.38 $Y2=0.8
cc_61 VPB N_VPWR_c_357_n 0.012566f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=1.075
cc_62 VPB N_VPWR_c_358_n 0.0352579f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=0.445
cc_63 VPB N_VPWR_c_359_n 0.00684629f $X=-0.19 $Y=1.655 $X2=2.97 $Y2=0.445
cc_64 VPB N_VPWR_c_360_n 0.0601917f $X=-0.19 $Y=1.655 $X2=3.33 $Y2=0.765
cc_65 VPB N_VPWR_c_361_n 0.00510842f $X=-0.19 $Y=1.655 $X2=3.33 $Y2=0.445
cc_66 VPB N_VPWR_c_362_n 0.0237525f $X=-0.19 $Y=1.655 $X2=2.525 $Y2=0.8
cc_67 VPB N_VPWR_c_356_n 0.0500474f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=0.8
cc_68 VPB N_Y_c_401_n 0.0132621f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=0.445
cc_69 VPB N_Y_c_406_n 0.0105794f $X=-0.19 $Y=1.655 $X2=2.97 $Y2=0.765
cc_70 VPB N_Y_c_407_n 0.0116422f $X=-0.19 $Y=1.655 $X2=2.97 $Y2=0.445
cc_71 VPB N_Y_c_408_n 0.00761768f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 N_S_c_85_n N_A0_M1010_g 9.61099e-19 $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_73 N_S_c_86_n N_A0_M1010_g 0.0122794f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_74 N_S_c_80_n N_A0_c_185_n 0.0131393f $X=1.21 $Y=1.16 $X2=0 $Y2=0
cc_75 N_S_c_81_n N_A0_c_185_n 6.49003e-19 $X=1.295 $Y=1.075 $X2=0 $Y2=0
cc_76 N_S_c_86_n N_A0_c_185_n 0.0127141f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_77 N_S_c_85_n N_A0_c_186_n 0.00152791f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_78 N_S_c_86_n N_A0_c_186_n 0.0368978f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_79 N_S_c_86_n N_A0_c_187_n 0.00400978f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_80 N_S_M1006_g N_A0_c_188_n 3.28058e-19 $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_81 N_S_c_72_n N_A0_c_188_n 3.71966e-19 $X=1.13 $Y=1.15 $X2=0 $Y2=0
cc_82 N_S_c_80_n N_A0_c_188_n 0.0260927f $X=1.21 $Y=1.16 $X2=0 $Y2=0
cc_83 N_S_c_83_n N_A0_c_188_n 0.018521f $X=0.605 $Y=1.24 $X2=0 $Y2=0
cc_84 N_S_c_84_n N_A0_c_188_n 9.67814e-19 $X=0.605 $Y=1.24 $X2=0 $Y2=0
cc_85 N_S_c_86_n N_A0_c_188_n 0.00575618f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_86 N_S_M1006_g N_A0_c_189_n 0.0824779f $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_87 N_S_c_72_n N_A0_c_189_n 0.016729f $X=1.13 $Y=1.15 $X2=0 $Y2=0
cc_88 N_S_c_80_n N_A0_c_189_n 0.00258061f $X=1.21 $Y=1.16 $X2=0 $Y2=0
cc_89 N_S_c_83_n N_A0_c_189_n 3.51769e-19 $X=0.605 $Y=1.24 $X2=0 $Y2=0
cc_90 N_S_c_84_n N_A0_c_189_n 0.0175938f $X=0.605 $Y=1.24 $X2=0 $Y2=0
cc_91 N_S_M1005_g N_A1_M1004_g 0.0602007f $X=1.205 $Y=0.445 $X2=0 $Y2=0
cc_92 N_S_c_80_n N_A1_M1004_g 0.00139318f $X=1.21 $Y=1.16 $X2=0 $Y2=0
cc_93 N_S_c_81_n N_A1_M1004_g 0.00381449f $X=1.295 $Y=1.075 $X2=0 $Y2=0
cc_94 N_S_c_86_n N_A1_M1004_g 0.0108054f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_95 N_S_M1003_g N_A_490_21#_M1001_g 0.024008f $X=3.175 $Y=2.595 $X2=0 $Y2=0
cc_96 N_S_c_75_n N_A_490_21#_c_292_n 0.011181f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_97 N_S_c_85_n N_A_490_21#_c_292_n 0.00190353f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_98 N_S_c_86_n N_A_490_21#_c_292_n 0.00212273f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_99 N_S_c_75_n N_A_490_21#_c_293_n 0.00166604f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_100 N_S_c_76_n N_A_490_21#_c_293_n 0.0180844f $X=3.175 $Y=1.28 $X2=0 $Y2=0
cc_101 N_S_c_85_n N_A_490_21#_c_293_n 0.0034705f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_102 N_S_c_86_n N_A_490_21#_c_293_n 0.00350991f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_103 N_S_c_76_n N_A_490_21#_c_294_n 0.00488496f $X=3.175 $Y=1.28 $X2=0 $Y2=0
cc_104 N_S_M1003_g N_A_490_21#_c_294_n 0.0247486f $X=3.175 $Y=2.595 $X2=0 $Y2=0
cc_105 N_S_c_85_n N_A_490_21#_c_294_n 0.040927f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_106 N_S_c_86_n N_A_490_21#_c_294_n 0.00144497f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_107 N_S_M1003_g N_A_490_21#_c_295_n 0.0181444f $X=3.175 $Y=2.595 $X2=0 $Y2=0
cc_108 N_S_c_85_n N_A_490_21#_c_295_n 0.00431096f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_109 N_S_M1003_g N_A_490_21#_c_302_n 0.0381513f $X=3.175 $Y=2.595 $X2=0 $Y2=0
cc_110 N_S_c_75_n N_A_490_21#_c_296_n 0.00168463f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_111 N_S_c_76_n N_A_490_21#_c_296_n 0.0174313f $X=3.175 $Y=1.28 $X2=0 $Y2=0
cc_112 N_S_c_78_n N_A_490_21#_c_296_n 0.0105728f $X=3.33 $Y=0.765 $X2=0 $Y2=0
cc_113 N_S_c_85_n N_A_490_21#_c_296_n 0.0297299f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_114 N_S_c_76_n N_A_490_21#_c_297_n 0.00310225f $X=3.175 $Y=1.28 $X2=0 $Y2=0
cc_115 N_S_M1003_g N_A_490_21#_c_297_n 0.00835871f $X=3.175 $Y=2.595 $X2=0 $Y2=0
cc_116 N_S_c_76_n N_A_490_21#_c_298_n 0.00866032f $X=3.175 $Y=1.28 $X2=0 $Y2=0
cc_117 N_S_c_85_n N_A_490_21#_c_298_n 0.00938609f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_118 N_S_c_86_n N_A_490_21#_c_298_n 0.00102836f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_119 N_S_M1006_g N_VPWR_c_358_n 0.0101011f $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_120 N_S_M1003_g N_VPWR_c_359_n 0.00345323f $X=3.175 $Y=2.595 $X2=0 $Y2=0
cc_121 N_S_M1006_g N_VPWR_c_360_n 0.00772576f $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_122 N_S_M1003_g N_VPWR_c_362_n 0.00939541f $X=3.175 $Y=2.595 $X2=0 $Y2=0
cc_123 N_S_M1006_g N_VPWR_c_356_n 0.0128874f $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_124 N_S_M1003_g N_VPWR_c_356_n 0.0170272f $X=3.175 $Y=2.595 $X2=0 $Y2=0
cc_125 N_S_M1006_g N_Y_c_401_n 0.00609602f $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_126 N_S_c_73_n N_Y_c_401_n 0.00116522f $X=0.77 $Y=1.15 $X2=0 $Y2=0
cc_127 N_S_c_83_n N_Y_c_401_n 0.0488899f $X=0.605 $Y=1.24 $X2=0 $Y2=0
cc_128 N_S_c_84_n N_Y_c_401_n 0.0111183f $X=0.605 $Y=1.24 $X2=0 $Y2=0
cc_129 N_S_c_72_n N_Y_c_402_n 0.00505358f $X=1.13 $Y=1.15 $X2=0 $Y2=0
cc_130 N_S_c_73_n N_Y_c_402_n 0.00226817f $X=0.77 $Y=1.15 $X2=0 $Y2=0
cc_131 N_S_M1005_g N_Y_c_402_n 0.00372938f $X=1.205 $Y=0.445 $X2=0 $Y2=0
cc_132 N_S_c_80_n N_Y_c_402_n 0.0191515f $X=1.21 $Y=1.16 $X2=0 $Y2=0
cc_133 N_S_c_81_n N_Y_c_402_n 7.40334e-19 $X=1.295 $Y=1.075 $X2=0 $Y2=0
cc_134 N_S_c_82_n N_Y_c_402_n 0.0136564f $X=1.38 $Y=0.8 $X2=0 $Y2=0
cc_135 N_S_c_83_n N_Y_c_402_n 0.0252203f $X=0.605 $Y=1.24 $X2=0 $Y2=0
cc_136 N_S_M1006_g N_Y_c_406_n 0.0120586f $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_137 N_S_c_79_n N_Y_c_406_n 3.37098e-19 $X=0.605 $Y=1.745 $X2=0 $Y2=0
cc_138 N_S_c_83_n N_Y_c_406_n 0.0120673f $X=0.605 $Y=1.24 $X2=0 $Y2=0
cc_139 N_S_M1005_g N_Y_c_404_n 0.00683717f $X=1.205 $Y=0.445 $X2=0 $Y2=0
cc_140 N_S_c_82_n N_Y_c_404_n 7.28787e-19 $X=1.38 $Y=0.8 $X2=0 $Y2=0
cc_141 N_S_c_72_n N_Y_c_425_n 0.00128461f $X=1.13 $Y=1.15 $X2=0 $Y2=0
cc_142 N_S_M1005_g N_Y_c_425_n 0.0162518f $X=1.205 $Y=0.445 $X2=0 $Y2=0
cc_143 N_S_c_80_n N_Y_c_425_n 0.00415947f $X=1.21 $Y=1.16 $X2=0 $Y2=0
cc_144 N_S_c_82_n N_Y_c_425_n 0.0104502f $X=1.38 $Y=0.8 $X2=0 $Y2=0
cc_145 N_S_c_86_n N_Y_c_425_n 0.0346132f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_146 N_S_M1006_g N_Y_c_430_n 0.00655714f $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_147 N_S_M1006_g Y 0.013895f $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_148 N_S_M1006_g N_Y_c_408_n 0.022409f $X=0.615 $Y=2.595 $X2=0 $Y2=0
cc_149 N_S_c_79_n N_Y_c_408_n 2.25414e-19 $X=0.605 $Y=1.745 $X2=0 $Y2=0
cc_150 N_S_c_83_n N_Y_c_408_n 0.0133705f $X=0.605 $Y=1.24 $X2=0 $Y2=0
cc_151 N_S_M1005_g N_VGND_c_487_n 0.00412089f $X=1.205 $Y=0.445 $X2=0 $Y2=0
cc_152 N_S_c_75_n N_VGND_c_488_n 0.00941898f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_153 N_S_c_78_n N_VGND_c_488_n 0.00198038f $X=3.33 $Y=0.765 $X2=0 $Y2=0
cc_154 N_S_c_85_n N_VGND_c_488_n 0.0210298f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_155 N_S_M1005_g N_VGND_c_491_n 0.00359964f $X=1.205 $Y=0.445 $X2=0 $Y2=0
cc_156 N_S_c_86_n N_VGND_c_491_n 0.0088477f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_157 N_S_c_75_n N_VGND_c_492_n 0.00392053f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_158 N_S_c_78_n N_VGND_c_492_n 0.00549284f $X=3.33 $Y=0.765 $X2=0 $Y2=0
cc_159 N_S_c_85_n N_VGND_c_492_n 0.00449058f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_160 N_S_M1005_g N_VGND_c_493_n 0.00674206f $X=1.205 $Y=0.445 $X2=0 $Y2=0
cc_161 N_S_c_75_n N_VGND_c_493_n 0.00444666f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_162 N_S_c_78_n N_VGND_c_493_n 0.0109191f $X=3.33 $Y=0.765 $X2=0 $Y2=0
cc_163 N_S_c_85_n N_VGND_c_493_n 0.00880474f $X=3.035 $Y=0.93 $X2=0 $Y2=0
cc_164 N_S_c_86_n N_VGND_c_493_n 0.0159135f $X=2.525 $Y=0.905 $X2=0 $Y2=0
cc_165 N_A0_M1010_g N_A1_M1004_g 0.0262049f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A0_c_185_n N_A1_M1004_g 0.0212466f $X=1.73 $Y=1.23 $X2=0 $Y2=0
cc_167 N_A0_c_186_n N_A1_M1004_g 5.48191e-19 $X=2.075 $Y=1.23 $X2=0 $Y2=0
cc_168 N_A0_c_187_n N_A1_M1004_g 0.0180888f $X=2.075 $Y=1.23 $X2=0 $Y2=0
cc_169 N_A0_c_188_n N_A1_M1004_g 0.0032969f $X=1.56 $Y=1.63 $X2=0 $Y2=0
cc_170 N_A0_c_189_n N_A1_M1004_g 0.0187929f $X=1.145 $Y=1.63 $X2=0 $Y2=0
cc_171 N_A0_M1007_g N_A1_c_249_n 0.0195235f $X=1.105 $Y=2.595 $X2=0 $Y2=0
cc_172 N_A0_c_185_n N_A1_c_249_n 0.00920573f $X=1.73 $Y=1.23 $X2=0 $Y2=0
cc_173 N_A0_c_186_n N_A1_c_249_n 0.00757552f $X=2.075 $Y=1.23 $X2=0 $Y2=0
cc_174 N_A0_c_187_n N_A1_c_249_n 0.0213824f $X=2.075 $Y=1.23 $X2=0 $Y2=0
cc_175 N_A0_c_188_n N_A1_c_249_n 0.00300457f $X=1.56 $Y=1.63 $X2=0 $Y2=0
cc_176 N_A0_c_189_n N_A1_c_249_n 7.58987e-19 $X=1.145 $Y=1.63 $X2=0 $Y2=0
cc_177 N_A0_M1007_g N_A1_c_250_n 0.00142537f $X=1.105 $Y=2.595 $X2=0 $Y2=0
cc_178 N_A0_c_185_n N_A1_c_250_n 0.013217f $X=1.73 $Y=1.23 $X2=0 $Y2=0
cc_179 N_A0_c_186_n N_A1_c_250_n 0.0217701f $X=2.075 $Y=1.23 $X2=0 $Y2=0
cc_180 N_A0_c_187_n N_A1_c_250_n 0.00122829f $X=2.075 $Y=1.23 $X2=0 $Y2=0
cc_181 N_A0_M1010_g N_A_490_21#_c_292_n 0.028558f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_182 N_A0_c_186_n N_A_490_21#_c_294_n 0.00363714f $X=2.075 $Y=1.23 $X2=0 $Y2=0
cc_183 N_A0_M1010_g N_A_490_21#_c_298_n 0.00618656f $X=2.035 $Y=0.445 $X2=0
+ $Y2=0
cc_184 N_A0_c_186_n N_A_490_21#_c_298_n 0.00165119f $X=2.075 $Y=1.23 $X2=0 $Y2=0
cc_185 N_A0_c_187_n N_A_490_21#_c_298_n 0.0169187f $X=2.075 $Y=1.23 $X2=0 $Y2=0
cc_186 N_A0_M1007_g N_VPWR_c_360_n 0.00599594f $X=1.105 $Y=2.595 $X2=0 $Y2=0
cc_187 N_A0_M1007_g N_VPWR_c_356_n 0.00844577f $X=1.105 $Y=2.595 $X2=0 $Y2=0
cc_188 N_A0_M1010_g N_Y_c_425_n 0.00542874f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A0_M1007_g N_Y_c_430_n 0.0112312f $X=1.105 $Y=2.595 $X2=0 $Y2=0
cc_190 N_A0_M1007_g N_Y_c_437_n 0.00197775f $X=1.105 $Y=2.595 $X2=0 $Y2=0
cc_191 N_A0_c_185_n N_Y_c_437_n 0.00674879f $X=1.73 $Y=1.23 $X2=0 $Y2=0
cc_192 N_A0_c_188_n N_Y_c_437_n 0.00242777f $X=1.56 $Y=1.63 $X2=0 $Y2=0
cc_193 N_A0_M1007_g Y 0.0197514f $X=1.105 $Y=2.595 $X2=0 $Y2=0
cc_194 N_A0_M1007_g N_Y_c_408_n 0.0251909f $X=1.105 $Y=2.595 $X2=0 $Y2=0
cc_195 N_A0_c_188_n N_Y_c_408_n 0.0155231f $X=1.56 $Y=1.63 $X2=0 $Y2=0
cc_196 N_A0_c_189_n N_Y_c_408_n 0.0015016f $X=1.145 $Y=1.63 $X2=0 $Y2=0
cc_197 N_A0_M1010_g N_VGND_c_488_n 0.00190478f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_198 N_A0_M1010_g N_VGND_c_491_n 0.00426284f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_199 N_A0_M1010_g N_VGND_c_493_n 0.00633491f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_200 N_A1_M1008_g N_A_490_21#_M1001_g 0.0361781f $X=1.925 $Y=2.595 $X2=0 $Y2=0
cc_201 N_A1_c_250_n N_A_490_21#_c_294_n 0.00433137f $X=2.075 $Y=1.77 $X2=0 $Y2=0
cc_202 N_A1_c_249_n N_A_490_21#_c_295_n 0.0173541f $X=1.925 $Y=1.77 $X2=0 $Y2=0
cc_203 N_A1_c_250_n N_A_490_21#_c_295_n 0.0107328f $X=2.075 $Y=1.77 $X2=0 $Y2=0
cc_204 N_A1_M1008_g N_VPWR_c_359_n 0.00465423f $X=1.925 $Y=2.595 $X2=0 $Y2=0
cc_205 N_A1_c_250_n N_VPWR_c_359_n 0.00290078f $X=2.075 $Y=1.77 $X2=0 $Y2=0
cc_206 N_A1_M1008_g N_VPWR_c_360_n 0.00938036f $X=1.925 $Y=2.595 $X2=0 $Y2=0
cc_207 N_A1_M1008_g N_VPWR_c_356_n 0.0171214f $X=1.925 $Y=2.595 $X2=0 $Y2=0
cc_208 N_A1_M1004_g N_Y_c_425_n 0.00998242f $X=1.595 $Y=0.445 $X2=0 $Y2=0
cc_209 N_A1_M1008_g N_Y_c_445_n 0.00437649f $X=1.925 $Y=2.595 $X2=0 $Y2=0
cc_210 N_A1_M1008_g N_Y_c_437_n 0.0141775f $X=1.925 $Y=2.595 $X2=0 $Y2=0
cc_211 N_A1_c_249_n N_Y_c_437_n 0.00228483f $X=1.925 $Y=1.77 $X2=0 $Y2=0
cc_212 N_A1_M1008_g Y 8.04506e-19 $X=1.925 $Y=2.595 $X2=0 $Y2=0
cc_213 N_A1_M1008_g N_Y_c_408_n 0.00421796f $X=1.925 $Y=2.595 $X2=0 $Y2=0
cc_214 N_A1_c_250_n N_Y_c_408_n 0.00171599f $X=2.075 $Y=1.77 $X2=0 $Y2=0
cc_215 N_A1_c_250_n A_410_419# 0.00812675f $X=2.075 $Y=1.77 $X2=-0.19 $Y2=-0.245
cc_216 N_A1_M1004_g N_VGND_c_491_n 0.00359964f $X=1.595 $Y=0.445 $X2=0 $Y2=0
cc_217 N_A1_M1004_g N_VGND_c_493_n 0.00538649f $X=1.595 $Y=0.445 $X2=0 $Y2=0
cc_218 N_A_490_21#_M1001_g N_VPWR_c_359_n 0.0284387f $X=2.605 $Y=2.595 $X2=0
+ $Y2=0
cc_219 N_A_490_21#_c_294_n N_VPWR_c_359_n 0.0152032f $X=3.275 $Y=1.5 $X2=0 $Y2=0
cc_220 N_A_490_21#_c_295_n N_VPWR_c_359_n 0.00160278f $X=2.645 $Y=1.5 $X2=0
+ $Y2=0
cc_221 N_A_490_21#_c_302_n N_VPWR_c_359_n 0.0300392f $X=3.44 $Y=2.24 $X2=0 $Y2=0
cc_222 N_A_490_21#_M1001_g N_VPWR_c_360_n 0.008763f $X=2.605 $Y=2.595 $X2=0
+ $Y2=0
cc_223 N_A_490_21#_c_302_n N_VPWR_c_362_n 0.0268376f $X=3.44 $Y=2.24 $X2=0 $Y2=0
cc_224 N_A_490_21#_M1003_d N_VPWR_c_356_n 0.0023218f $X=3.3 $Y=2.095 $X2=0 $Y2=0
cc_225 N_A_490_21#_M1001_g N_VPWR_c_356_n 0.0149113f $X=2.605 $Y=2.595 $X2=0
+ $Y2=0
cc_226 N_A_490_21#_c_302_n N_VPWR_c_356_n 0.0165708f $X=3.44 $Y=2.24 $X2=0 $Y2=0
cc_227 N_A_490_21#_c_292_n N_Y_c_425_n 8.1197e-19 $X=2.54 $Y=0.73 $X2=0 $Y2=0
cc_228 N_A_490_21#_M1001_g N_Y_c_445_n 6.96967e-19 $X=2.605 $Y=2.595 $X2=0 $Y2=0
cc_229 N_A_490_21#_M1001_g N_Y_c_437_n 0.00233049f $X=2.605 $Y=2.595 $X2=0 $Y2=0
cc_230 N_A_490_21#_c_292_n N_VGND_c_488_n 0.010508f $X=2.54 $Y=0.73 $X2=0 $Y2=0
cc_231 N_A_490_21#_c_296_n N_VGND_c_488_n 0.00886789f $X=3.545 $Y=0.47 $X2=0
+ $Y2=0
cc_232 N_A_490_21#_c_292_n N_VGND_c_491_n 0.00377504f $X=2.54 $Y=0.73 $X2=0
+ $Y2=0
cc_233 N_A_490_21#_c_296_n N_VGND_c_492_n 0.0197885f $X=3.545 $Y=0.47 $X2=0
+ $Y2=0
cc_234 N_A_490_21#_M1009_d N_VGND_c_493_n 0.00232985f $X=3.405 $Y=0.235 $X2=0
+ $Y2=0
cc_235 N_A_490_21#_c_292_n N_VGND_c_493_n 0.00468318f $X=2.54 $Y=0.73 $X2=0
+ $Y2=0
cc_236 N_A_490_21#_c_296_n N_VGND_c_493_n 0.0125808f $X=3.545 $Y=0.47 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_356_n A_148_419# 0.00193225f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_238 N_VPWR_c_356_n N_Y_M1007_d 0.00465189f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_c_358_n N_Y_c_406_n 0.0129704f $X=0.34 $Y=2.44 $X2=0 $Y2=0
cc_240 N_VPWR_M1006_s N_Y_c_407_n 7.36937e-19 $X=0.195 $Y=2.095 $X2=0 $Y2=0
cc_241 N_VPWR_c_358_n N_Y_c_407_n 0.00732286f $X=0.34 $Y=2.44 $X2=0 $Y2=0
cc_242 N_VPWR_c_360_n N_Y_c_445_n 0.0305392f $X=2.705 $Y=3.33 $X2=0 $Y2=0
cc_243 N_VPWR_c_356_n N_Y_c_445_n 0.0192996f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_358_n N_Y_c_430_n 0.0131326f $X=0.34 $Y=2.44 $X2=0 $Y2=0
cc_245 N_VPWR_c_360_n N_Y_c_430_n 0.0405279f $X=2.705 $Y=3.33 $X2=0 $Y2=0
cc_246 N_VPWR_c_356_n N_Y_c_430_n 0.0256988f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_247 N_VPWR_c_358_n Y 0.034258f $X=0.34 $Y=2.44 $X2=0 $Y2=0
cc_248 N_VPWR_c_358_n N_Y_c_408_n 0.0135653f $X=0.34 $Y=2.44 $X2=0 $Y2=0
cc_249 N_VPWR_c_356_n A_410_419# 0.0184401f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_250 A_148_419# N_Y_c_430_n 0.00125965f $X=0.74 $Y=2.095 $X2=0 $Y2=3.085
cc_251 A_148_419# N_Y_c_408_n 0.00568393f $X=0.74 $Y=2.095 $X2=0.24 $Y2=3.33
cc_252 N_Y_c_404_n N_VGND_M1005_s 0.0062092f $X=0.945 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_253 N_Y_c_468_p N_VGND_M1005_s 0.00610898f $X=1.03 $Y=0.4 $X2=-0.19
+ $Y2=-0.245
cc_254 N_Y_c_425_n N_VGND_M1005_s 0.00109276f $X=1.815 $Y=0.44 $X2=-0.19
+ $Y2=-0.245
cc_255 N_Y_c_402_n N_VGND_c_487_n 0.0248587f $X=0.86 $Y=0.81 $X2=0 $Y2=0
cc_256 N_Y_c_404_n N_VGND_c_487_n 6.97618e-19 $X=0.945 $Y=0.725 $X2=0 $Y2=0
cc_257 N_Y_c_468_p N_VGND_c_487_n 0.0220318f $X=1.03 $Y=0.4 $X2=0 $Y2=0
cc_258 N_Y_c_425_n N_VGND_c_488_n 0.00751108f $X=1.815 $Y=0.44 $X2=0 $Y2=0
cc_259 N_Y_c_402_n N_VGND_c_489_n 0.00135325f $X=0.86 $Y=0.81 $X2=0 $Y2=0
cc_260 N_Y_c_403_n N_VGND_c_489_n 0.0028865f $X=0.26 $Y=0.81 $X2=0 $Y2=0
cc_261 N_Y_c_402_n N_VGND_c_491_n 0.00272171f $X=0.86 $Y=0.81 $X2=0 $Y2=0
cc_262 N_Y_c_468_p N_VGND_c_491_n 0.0111686f $X=1.03 $Y=0.4 $X2=0 $Y2=0
cc_263 N_Y_c_425_n N_VGND_c_491_n 0.0496931f $X=1.815 $Y=0.44 $X2=0 $Y2=0
cc_264 N_Y_M1004_d N_VGND_c_493_n 0.00231907f $X=1.67 $Y=0.235 $X2=0 $Y2=0
cc_265 N_Y_c_402_n N_VGND_c_493_n 0.00854741f $X=0.86 $Y=0.81 $X2=0 $Y2=0
cc_266 N_Y_c_403_n N_VGND_c_493_n 0.0048263f $X=0.26 $Y=0.81 $X2=0 $Y2=0
cc_267 N_Y_c_468_p N_VGND_c_493_n 0.00656418f $X=1.03 $Y=0.4 $X2=0 $Y2=0
cc_268 N_Y_c_425_n N_VGND_c_493_n 0.0342648f $X=1.815 $Y=0.44 $X2=0 $Y2=0
cc_269 N_Y_c_425_n A_256_47# 0.00262077f $X=1.815 $Y=0.44 $X2=-0.19 $Y2=-0.245
cc_270 N_VGND_c_493_n A_256_47# 0.00193256f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_271 N_VGND_c_493_n A_422_47# 0.00435305f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_272 N_VGND_c_493_n A_609_47# 0.00434009f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
