* NGSPICE file created from sky130_fd_sc_lp__o2111a_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o2111a_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VPWR C1 a_80_21# VPB phighvt w=640000u l=150000u
+  ad=7.904e+11p pd=6.31e+06u as=3.584e+11p ps=3.68e+06u
M1001 a_315_47# D1 a_80_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1002 VPWR a_80_21# X VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1003 VGND a_80_21# X VNB nshort w=420000u l=150000u
+  ad=2.583e+11p pd=2.91e+06u as=1.113e+11p ps=1.37e+06u
M1004 a_387_47# C1 a_315_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 a_459_47# B1 a_387_47# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1006 a_585_481# A2 a_80_21# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1007 VPWR A1 a_585_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_80_21# D1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_459_47# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_459_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_80_21# B1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

