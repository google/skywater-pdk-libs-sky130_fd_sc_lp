* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_478_47# A2 a_550_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_346_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 X a_113_237# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 X a_113_237# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR A4 a_346_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND B1 a_113_237# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR A2 a_346_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_550_47# A3 a_658_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_658_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_346_367# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_113_237# A1 a_478_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_113_237# B1 a_346_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
