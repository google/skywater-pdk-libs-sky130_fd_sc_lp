# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfrtp_lp2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfrtp_lp2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.32000 BY  3.330000 ;
  SYMMETRY R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 1.510000 0.905000 1.840000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.645000 1.920000 16.205000 2.960000 ;
        RECT 15.875000 0.430000 16.205000 1.920000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.939000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  2.975000 1.550000  3.265000 1.595000 ;
        RECT  2.975000 1.595000 12.865000 1.735000 ;
        RECT  2.975000 1.735000  3.265000 1.780000 ;
        RECT  8.735000 1.550000  9.025000 1.595000 ;
        RECT  8.735000 1.735000  9.025000 1.780000 ;
        RECT 12.575000 1.550000 12.865000 1.595000 ;
        RECT 12.575000 1.735000 12.865000 1.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 1.450000 2.255000 1.780000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.550000 1.685000 1.960000 ;
        RECT 1.085000 1.960000 3.655000 2.130000 ;
        RECT 3.485000 1.555000 3.875000 1.885000 ;
        RECT 3.485000 1.885000 3.655000 1.960000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.825000 1.170000 5.155000 1.500000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 16.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.320000 0.085000 ;
      RECT  0.000000  3.245000 16.320000 3.415000 ;
      RECT  0.090000  0.620000  1.480000 0.790000 ;
      RECT  0.090000  0.790000  0.260000 2.075000 ;
      RECT  0.090000  2.075000  0.890000 2.310000 ;
      RECT  0.090000  2.310000  3.020000 2.480000 ;
      RECT  0.090000  2.480000  0.890000 3.065000 ;
      RECT  0.170000  0.265000  2.380000 0.435000 ;
      RECT  0.170000  0.435000  0.500000 0.440000 ;
      RECT  0.440000  0.970000  0.735000 1.100000 ;
      RECT  0.440000  1.100000  4.225000 1.270000 ;
      RECT  0.440000  1.270000  0.735000 1.300000 ;
      RECT  1.150000  0.615000  1.480000 0.620000 ;
      RECT  1.150000  0.790000  1.480000 0.865000 ;
      RECT  1.580000  2.660000  1.910000 3.245000 ;
      RECT  2.050000  0.435000  2.380000 0.880000 ;
      RECT  2.435000  1.270000  2.765000 1.780000 ;
      RECT  2.560000  0.085000  2.890000 0.880000 ;
      RECT  2.690000  2.480000  3.020000 2.505000 ;
      RECT  2.690000  2.505000  3.900000 2.675000 ;
      RECT  2.690000  2.675000  3.020000 3.065000 ;
      RECT  2.975000  1.450000  3.305000 1.780000 ;
      RECT  3.220000  2.855000  3.550000 3.245000 ;
      RECT  3.730000  2.675000  3.900000 2.895000 ;
      RECT  3.730000  2.895000  5.010000 3.065000 ;
      RECT  3.820000  0.595000  4.225000 1.100000 ;
      RECT  3.835000  2.075000  4.225000 2.325000 ;
      RECT  4.055000  1.270000  4.225000 2.075000 ;
      RECT  4.420000  0.635000  4.590000 1.680000 ;
      RECT  4.420000  1.680000  5.805000 1.850000 ;
      RECT  4.420000  1.850000  4.670000 2.715000 ;
      RECT  4.840000  2.460000  7.035000 2.630000 ;
      RECT  4.840000  2.630000  5.010000 2.895000 ;
      RECT  5.180000  2.810000  5.510000 3.245000 ;
      RECT  5.210000  0.085000  5.540000 0.725000 ;
      RECT  5.475000  1.180000  5.805000 1.680000 ;
      RECT  5.710000  2.030000  6.290000 2.280000 ;
      RECT  5.975000  1.450000  6.685000 1.780000 ;
      RECT  5.975000  1.780000  6.290000 2.030000 ;
      RECT  6.070000  0.595000  6.455000 1.450000 ;
      RECT  6.705000  0.595000  7.035000 1.145000 ;
      RECT  6.865000  1.145000  7.035000 2.460000 ;
      RECT  6.865000  2.630000  7.035000 2.755000 ;
      RECT  7.215000  0.625000  7.385000 1.790000 ;
      RECT  7.215000  1.790000  7.790000 1.960000 ;
      RECT  7.215000  1.960000  9.700000 2.130000 ;
      RECT  7.215000  2.130000  7.790000 2.755000 ;
      RECT  7.555000  0.625000 10.425000 0.795000 ;
      RECT  7.555000  0.795000  7.725000 1.525000 ;
      RECT  8.225000  0.975000 10.040000 1.145000 ;
      RECT  8.225000  1.145000  8.555000 1.525000 ;
      RECT  8.585000  2.310000  8.915000 3.245000 ;
      RECT  8.765000  1.325000  9.200000 1.645000 ;
      RECT  8.765000  1.645000  9.185000 1.780000 ;
      RECT  8.850000  0.085000  9.180000 0.445000 ;
      RECT  9.275000  2.130000  9.700000 2.755000 ;
      RECT  9.355000  1.715000  9.700000 1.960000 ;
      RECT  9.370000  1.325000  9.700000 1.715000 ;
      RECT  9.870000  1.145000 10.040000 1.275000 ;
      RECT  9.870000  1.275000 10.775000 1.445000 ;
      RECT 10.005000  0.275000 10.775000 0.445000 ;
      RECT 10.080000  1.685000 10.410000 3.245000 ;
      RECT 10.210000  0.795000 10.425000 1.095000 ;
      RECT 10.605000  0.445000 10.775000 1.275000 ;
      RECT 10.605000  1.445000 10.775000 1.685000 ;
      RECT 10.605000  1.685000 11.020000 2.725000 ;
      RECT 10.955000  1.120000 12.105000 1.450000 ;
      RECT 11.300000  1.685000 12.455000 1.855000 ;
      RECT 11.300000  1.855000 11.630000 3.065000 ;
      RECT 11.510000  0.265000 11.840000 0.505000 ;
      RECT 11.510000  0.505000 12.455000 0.675000 ;
      RECT 11.815000  0.910000 12.105000 1.120000 ;
      RECT 12.285000  0.675000 12.455000 0.690000 ;
      RECT 12.285000  0.690000 13.845000 0.860000 ;
      RECT 12.285000  0.860000 12.455000 1.685000 ;
      RECT 12.400000  2.075000 12.650000 3.245000 ;
      RECT 12.635000  0.085000 12.965000 0.510000 ;
      RECT 12.635000  1.040000 13.185000 1.265000 ;
      RECT 12.635000  1.265000 14.195000 1.370000 ;
      RECT 12.635000  1.550000 12.835000 1.615000 ;
      RECT 12.635000  1.615000 13.485000 1.785000 ;
      RECT 13.015000  1.370000 14.195000 1.435000 ;
      RECT 13.085000  1.785000 13.485000 1.935000 ;
      RECT 13.085000  1.935000 13.315000 2.890000 ;
      RECT 13.495000  2.115000 13.835000 3.065000 ;
      RECT 13.515000  0.860000 13.845000 1.085000 ;
      RECT 13.665000  1.435000 13.835000 2.115000 ;
      RECT 13.670000  0.295000 14.195000 0.510000 ;
      RECT 14.025000  0.510000 14.195000 1.265000 ;
      RECT 14.025000  2.075000 14.355000 3.245000 ;
      RECT 14.375000  0.430000 14.705000 0.890000 ;
      RECT 14.535000  0.890000 14.705000 1.570000 ;
      RECT 14.535000  1.570000 15.680000 1.740000 ;
      RECT 14.535000  1.740000 14.915000 2.960000 ;
      RECT 15.085000  0.085000 15.415000 0.890000 ;
      RECT 15.115000  1.920000 15.445000 3.245000 ;
      RECT 15.350000  1.070000 15.680000 1.570000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.580000  3.205000 1.750000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.580000  8.965000 1.750000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  1.580000 12.805000 1.750000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfrtp_lp2
