* File: sky130_fd_sc_lp__a21boi_2.pxi.spice
* Created: Wed Sep  2 09:19:24 2020
* 
x_PM_SKY130_FD_SC_LP__A21BOI_2%B1_N N_B1_N_M1011_g N_B1_N_c_83_n N_B1_N_c_84_n
+ N_B1_N_c_85_n N_B1_N_M1012_g N_B1_N_c_86_n B1_N B1_N B1_N B1_N B1_N B1_N
+ N_B1_N_c_88_n PM_SKY130_FD_SC_LP__A21BOI_2%B1_N
x_PM_SKY130_FD_SC_LP__A21BOI_2%A_119_500# N_A_119_500#_M1012_s
+ N_A_119_500#_M1011_d N_A_119_500#_c_117_n N_A_119_500#_c_118_n
+ N_A_119_500#_M1002_g N_A_119_500#_M1004_g N_A_119_500#_c_120_n
+ N_A_119_500#_c_121_n N_A_119_500#_M1007_g N_A_119_500#_M1010_g
+ N_A_119_500#_c_123_n N_A_119_500#_c_124_n N_A_119_500#_c_125_n
+ N_A_119_500#_c_126_n N_A_119_500#_c_127_n N_A_119_500#_c_128_n
+ PM_SKY130_FD_SC_LP__A21BOI_2%A_119_500#
x_PM_SKY130_FD_SC_LP__A21BOI_2%A2 N_A2_M1001_g N_A2_M1009_g N_A2_M1013_g
+ N_A2_M1008_g N_A2_c_196_n N_A2_c_197_n N_A2_c_198_n N_A2_c_199_n N_A2_c_200_n
+ N_A2_c_201_n A2 A2 A2 A2 PM_SKY130_FD_SC_LP__A21BOI_2%A2
x_PM_SKY130_FD_SC_LP__A21BOI_2%A1 N_A1_M1003_g N_A1_M1000_g N_A1_M1005_g
+ N_A1_M1006_g A1 N_A1_c_290_n PM_SKY130_FD_SC_LP__A21BOI_2%A1
x_PM_SKY130_FD_SC_LP__A21BOI_2%VPWR N_VPWR_M1011_s N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_348_n VPWR
+ N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_344_n N_VPWR_c_353_n
+ N_VPWR_c_354_n PM_SKY130_FD_SC_LP__A21BOI_2%VPWR
x_PM_SKY130_FD_SC_LP__A21BOI_2%A_231_367# N_A_231_367#_M1004_d
+ N_A_231_367#_M1010_d N_A_231_367#_M1000_s N_A_231_367#_M1008_s
+ N_A_231_367#_c_402_n N_A_231_367#_c_403_n N_A_231_367#_c_413_n
+ N_A_231_367#_c_404_n N_A_231_367#_c_420_n N_A_231_367#_c_421_n
+ N_A_231_367#_c_425_n N_A_231_367#_c_426_n N_A_231_367#_c_405_n
+ N_A_231_367#_c_434_n N_A_231_367#_c_435_n N_A_231_367#_c_406_n
+ PM_SKY130_FD_SC_LP__A21BOI_2%A_231_367#
x_PM_SKY130_FD_SC_LP__A21BOI_2%Y N_Y_M1002_d N_Y_M1003_d N_Y_M1004_s N_Y_c_466_n
+ N_Y_c_502_n Y Y Y Y Y Y N_Y_c_467_n Y Y PM_SKY130_FD_SC_LP__A21BOI_2%Y
x_PM_SKY130_FD_SC_LP__A21BOI_2%VGND N_VGND_M1012_d N_VGND_M1007_s N_VGND_M1013_s
+ N_VGND_c_522_n N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n VGND
+ N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n N_VGND_c_530_n
+ N_VGND_c_531_n PM_SKY130_FD_SC_LP__A21BOI_2%VGND
x_PM_SKY130_FD_SC_LP__A21BOI_2%A_502_65# N_A_502_65#_M1009_d N_A_502_65#_M1005_s
+ N_A_502_65#_c_582_n N_A_502_65#_c_579_n N_A_502_65#_c_580_n
+ N_A_502_65#_c_581_n PM_SKY130_FD_SC_LP__A21BOI_2%A_502_65#
cc_1 VNB N_B1_N_M1011_g 0.00816182f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.71
cc_2 VNB N_B1_N_c_83_n 0.030621f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.93
cc_3 VNB N_B1_N_c_84_n 0.022726f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.93
cc_4 VNB N_B1_N_c_85_n 0.0223715f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.855
cc_5 VNB N_B1_N_c_86_n 0.0224829f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.525
cc_6 VNB B1_N 0.0628231f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_7 VNB N_B1_N_c_88_n 0.0300086f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.02
cc_8 VNB N_A_119_500#_c_117_n 0.0182331f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.855
cc_9 VNB N_A_119_500#_c_118_n 0.0178732f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.535
cc_10 VNB N_A_119_500#_M1004_g 0.0110173f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_11 VNB N_A_119_500#_c_120_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_A_119_500#_c_121_n 0.0162997f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_13 VNB N_A_119_500#_M1010_g 0.0116313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_119_500#_c_123_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.02
cc_15 VNB N_A_119_500#_c_124_n 0.0055116f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.02
cc_16 VNB N_A_119_500#_c_125_n 0.00605282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_119_500#_c_126_n 0.0013732f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.02
cc_18 VNB N_A_119_500#_c_127_n 0.00408685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_119_500#_c_128_n 0.0399477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_M1009_g 0.0208387f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.855
cc_21 VNB N_A2_M1013_g 0.0269357f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.338
cc_22 VNB N_A2_c_196_n 4.19707e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_23 VNB N_A2_c_197_n 6.84753e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_198_n 0.0235074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A2_c_199_n 0.0027694f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.02
cc_26 VNB N_A2_c_200_n 0.0167799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A2_c_201_n 0.0290222f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=0.925
cc_28 VNB N_A1_M1003_g 0.0203468f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.71
cc_29 VNB N_A1_M1005_g 0.0208263f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.338
cc_30 VNB A1 0.00148046f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_31 VNB N_A1_c_290_n 0.0358454f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.02
cc_32 VNB N_VPWR_c_344_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=2.405
cc_33 VNB N_Y_c_466_n 0.0161811f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.005
cc_34 VNB N_Y_c_467_n 0.00209028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB Y 0.0022815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_522_n 0.012771f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.525
cc_37 VNB N_VGND_c_523_n 0.00464497f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_38 VNB N_VGND_c_524_n 0.0121815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_525_n 0.0463167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_526_n 0.0323636f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.02
cc_41 VNB N_VGND_c_527_n 0.0162863f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=0.925
cc_42 VNB N_VGND_c_528_n 0.0389928f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.665
cc_43 VNB N_VGND_c_529_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_530_n 0.00581671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_531_n 0.254937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_502_65#_c_579_n 0.00513958f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.338
cc_47 VNB N_A_502_65#_c_580_n 0.00207236f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.525
cc_48 VNB N_A_502_65#_c_581_n 0.00300049f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_49 VPB N_B1_N_M1011_g 0.069264f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.71
cc_50 VPB B1_N 0.0407406f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.47
cc_51 VPB N_A_119_500#_M1004_g 0.023601f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_52 VPB N_A_119_500#_M1010_g 0.0199541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_119_500#_c_126_n 0.0228807f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.02
cc_54 VPB N_A2_M1001_g 0.0200092f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.71
cc_55 VPB N_A2_M1008_g 0.0247293f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_56 VPB N_A2_c_196_n 0.0015121f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_57 VPB N_A2_c_197_n 0.00150234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A2_c_198_n 0.00654571f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A2_c_201_n 0.00656679f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=0.925
cc_60 VPB N_A1_M1000_g 0.0198787f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=0.855
cc_61 VPB N_A1_M1006_g 0.0184692f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_62 VPB A1 0.00402995f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_63 VPB N_A1_c_290_n 0.00713887f $X=-0.19 $Y=1.655 $X2=0.407 $Y2=1.02
cc_64 VPB N_VPWR_c_345_n 0.0129883f $X=-0.19 $Y=1.655 $X2=0.407 $Y2=1.005
cc_65 VPB N_VPWR_c_346_n 0.0230554f $X=-0.19 $Y=1.655 $X2=0.407 $Y2=1.525
cc_66 VPB N_VPWR_c_347_n 0.00495471f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_67 VPB N_VPWR_c_348_n 4.12476e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_349_n 0.050759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_350_n 0.016248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_351_n 0.0166487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_344_n 0.0620912f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=2.405
cc_72 VPB N_VPWR_c_353_n 0.00631788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_354_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_231_367#_c_402_n 0.00276803f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.47
cc_75 VPB N_A_231_367#_c_403_n 0.0129436f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_76 VPB N_A_231_367#_c_404_n 0.00323528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_231_367#_c_405_n 0.021061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_231_367#_c_406_n 0.0305687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB Y 7.57264e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB Y 0.00153678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 N_B1_N_c_85_n N_A_119_500#_c_118_n 0.0095716f $X=0.97 $Y=0.855 $X2=0 $Y2=0
cc_82 N_B1_N_c_83_n N_A_119_500#_c_125_n 0.017881f $X=0.895 $Y=0.93 $X2=0 $Y2=0
cc_83 N_B1_N_c_85_n N_A_119_500#_c_125_n 0.00793581f $X=0.97 $Y=0.855 $X2=0
+ $Y2=0
cc_84 B1_N N_A_119_500#_c_125_n 0.0774505f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_85 N_B1_N_c_88_n N_A_119_500#_c_125_n 0.00778306f $X=0.385 $Y=1.02 $X2=0
+ $Y2=0
cc_86 N_B1_N_M1011_g N_A_119_500#_c_126_n 0.0205915f $X=0.52 $Y=2.71 $X2=0 $Y2=0
cc_87 B1_N N_A_119_500#_c_126_n 0.0695153f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_88 N_B1_N_c_83_n N_A_119_500#_c_127_n 0.00149094f $X=0.895 $Y=0.93 $X2=0
+ $Y2=0
cc_89 N_B1_N_c_86_n N_A_119_500#_c_127_n 0.00210931f $X=0.407 $Y=1.525 $X2=0
+ $Y2=0
cc_90 B1_N N_A_119_500#_c_127_n 0.0219066f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_91 N_B1_N_c_83_n N_A_119_500#_c_128_n 0.010963f $X=0.895 $Y=0.93 $X2=0 $Y2=0
cc_92 B1_N N_A_119_500#_c_128_n 2.42458e-19 $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_93 N_B1_N_c_88_n N_A_119_500#_c_128_n 0.0170499f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_94 N_B1_N_M1011_g N_VPWR_c_346_n 0.00956706f $X=0.52 $Y=2.71 $X2=0 $Y2=0
cc_95 B1_N N_VPWR_c_346_n 0.0266999f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_96 N_B1_N_M1011_g N_VPWR_c_349_n 0.00455951f $X=0.52 $Y=2.71 $X2=0 $Y2=0
cc_97 N_B1_N_M1011_g N_VPWR_c_344_n 0.00447788f $X=0.52 $Y=2.71 $X2=0 $Y2=0
cc_98 B1_N N_VPWR_c_344_n 0.00335395f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_99 N_B1_N_M1011_g N_A_231_367#_c_402_n 0.00246733f $X=0.52 $Y=2.71 $X2=0
+ $Y2=0
cc_100 N_B1_N_c_85_n N_VGND_c_522_n 0.00781693f $X=0.97 $Y=0.855 $X2=0 $Y2=0
cc_101 B1_N N_VGND_c_522_n 0.00154784f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_102 N_B1_N_c_85_n N_VGND_c_526_n 0.0047088f $X=0.97 $Y=0.855 $X2=0 $Y2=0
cc_103 B1_N N_VGND_c_526_n 0.0194208f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_104 N_B1_N_c_84_n N_VGND_c_531_n 0.00411719f $X=0.595 $Y=0.93 $X2=0 $Y2=0
cc_105 N_B1_N_c_85_n N_VGND_c_531_n 0.00955492f $X=0.97 $Y=0.855 $X2=0 $Y2=0
cc_106 B1_N N_VGND_c_531_n 0.0143955f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_107 N_A_119_500#_M1010_g N_A2_M1001_g 0.0181634f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_A_119_500#_c_121_n N_A2_M1009_g 0.0242958f $X=1.925 $Y=1.275 $X2=0
+ $Y2=0
cc_109 N_A_119_500#_M1010_g N_A2_c_196_n 7.03961e-19 $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_119_500#_c_124_n N_A2_c_198_n 0.0171939f $X=1.925 $Y=1.35 $X2=0 $Y2=0
cc_111 N_A_119_500#_M1010_g N_A2_c_199_n 6.17958e-19 $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_112 N_A_119_500#_M1004_g N_VPWR_c_349_n 0.00357877f $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_119_500#_M1010_g N_VPWR_c_349_n 0.00357877f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_119_500#_c_126_n N_VPWR_c_349_n 0.00768407f $X=0.735 $Y=2.71 $X2=0
+ $Y2=0
cc_115 N_A_119_500#_M1004_g N_VPWR_c_344_n 0.00665089f $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_119_500#_M1010_g N_VPWR_c_344_n 0.00537654f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_119_500#_c_126_n N_VPWR_c_344_n 0.0089047f $X=0.735 $Y=2.71 $X2=0
+ $Y2=0
cc_118 N_A_119_500#_c_117_n N_A_231_367#_c_403_n 0.00410225f $X=1.42 $Y=1.35
+ $X2=0 $Y2=0
cc_119 N_A_119_500#_M1004_g N_A_231_367#_c_403_n 0.00272392f $X=1.495 $Y=2.465
+ $X2=0 $Y2=0
cc_120 N_A_119_500#_c_126_n N_A_231_367#_c_403_n 0.0712055f $X=0.735 $Y=2.71
+ $X2=0 $Y2=0
cc_121 N_A_119_500#_c_127_n N_A_231_367#_c_403_n 0.00330209f $X=1 $Y=1.44 $X2=0
+ $Y2=0
cc_122 N_A_119_500#_c_128_n N_A_231_367#_c_403_n 0.00110876f $X=1 $Y=1.35 $X2=0
+ $Y2=0
cc_123 N_A_119_500#_M1004_g N_A_231_367#_c_413_n 0.011508f $X=1.495 $Y=2.465
+ $X2=0 $Y2=0
cc_124 N_A_119_500#_M1010_g N_A_231_367#_c_413_n 0.011508f $X=1.925 $Y=2.465
+ $X2=0 $Y2=0
cc_125 N_A_119_500#_M1010_g N_A_231_367#_c_404_n 3.12571e-19 $X=1.925 $Y=2.465
+ $X2=0 $Y2=0
cc_126 N_A_119_500#_c_121_n N_Y_c_466_n 0.01769f $X=1.925 $Y=1.275 $X2=0 $Y2=0
cc_127 N_A_119_500#_c_118_n Y 0.00358065f $X=1.495 $Y=1.275 $X2=0 $Y2=0
cc_128 N_A_119_500#_c_125_n Y 0.00229748f $X=0.755 $Y=0.535 $X2=0 $Y2=0
cc_129 N_A_119_500#_M1004_g Y 0.00199061f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A_119_500#_M1010_g Y 0.00248941f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A_119_500#_c_118_n N_Y_c_467_n 0.00993108f $X=1.495 $Y=1.275 $X2=0
+ $Y2=0
cc_132 N_A_119_500#_c_121_n N_Y_c_467_n 8.74036e-19 $X=1.925 $Y=1.275 $X2=0
+ $Y2=0
cc_133 N_A_119_500#_c_118_n Y 8.57102e-19 $X=1.495 $Y=1.275 $X2=0 $Y2=0
cc_134 N_A_119_500#_M1004_g Y 0.0108745f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_119_500#_c_120_n Y 0.0105871f $X=1.85 $Y=1.35 $X2=0 $Y2=0
cc_136 N_A_119_500#_c_121_n Y 7.45058e-19 $X=1.925 $Y=1.275 $X2=0 $Y2=0
cc_137 N_A_119_500#_M1010_g Y 0.00496417f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A_119_500#_c_123_n Y 0.00399874f $X=1.495 $Y=1.35 $X2=0 $Y2=0
cc_139 N_A_119_500#_c_125_n Y 0.00243272f $X=0.755 $Y=0.535 $X2=0 $Y2=0
cc_140 N_A_119_500#_c_126_n Y 0.00621679f $X=0.735 $Y=2.71 $X2=0 $Y2=0
cc_141 N_A_119_500#_c_127_n Y 0.0105074f $X=1 $Y=1.44 $X2=0 $Y2=0
cc_142 N_A_119_500#_M1004_g Y 0.00825888f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_119_500#_M1010_g Y 0.00784738f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_119_500#_c_118_n N_VGND_c_522_n 0.00245325f $X=1.495 $Y=1.275 $X2=0
+ $Y2=0
cc_145 N_A_119_500#_c_125_n N_VGND_c_522_n 0.0554673f $X=0.755 $Y=0.535 $X2=0
+ $Y2=0
cc_146 N_A_119_500#_c_127_n N_VGND_c_522_n 0.00407089f $X=1 $Y=1.44 $X2=0 $Y2=0
cc_147 N_A_119_500#_c_128_n N_VGND_c_522_n 0.00732175f $X=1 $Y=1.35 $X2=0 $Y2=0
cc_148 N_A_119_500#_c_118_n N_VGND_c_523_n 5.48845e-19 $X=1.495 $Y=1.275 $X2=0
+ $Y2=0
cc_149 N_A_119_500#_c_121_n N_VGND_c_523_n 0.0101045f $X=1.925 $Y=1.275 $X2=0
+ $Y2=0
cc_150 N_A_119_500#_c_125_n N_VGND_c_526_n 0.0100258f $X=0.755 $Y=0.535 $X2=0
+ $Y2=0
cc_151 N_A_119_500#_c_118_n N_VGND_c_527_n 0.0046877f $X=1.495 $Y=1.275 $X2=0
+ $Y2=0
cc_152 N_A_119_500#_c_121_n N_VGND_c_527_n 0.00414769f $X=1.925 $Y=1.275 $X2=0
+ $Y2=0
cc_153 N_A_119_500#_c_118_n N_VGND_c_531_n 0.00898771f $X=1.495 $Y=1.275 $X2=0
+ $Y2=0
cc_154 N_A_119_500#_c_121_n N_VGND_c_531_n 0.00787505f $X=1.925 $Y=1.275 $X2=0
+ $Y2=0
cc_155 N_A_119_500#_c_125_n N_VGND_c_531_n 0.0100136f $X=0.755 $Y=0.535 $X2=0
+ $Y2=0
cc_156 N_A2_M1009_g N_A1_M1003_g 0.0216198f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_157 N_A2_M1001_g N_A1_M1000_g 0.0355065f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A2_c_196_n N_A1_M1000_g 0.00364947f $X=2.51 $Y=1.925 $X2=0 $Y2=0
cc_159 A2 N_A1_M1000_g 0.0123339f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_160 N_A2_M1013_g N_A1_M1005_g 0.0285162f $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_161 N_A2_M1008_g N_A1_M1006_g 0.0285162f $X=3.805 $Y=2.465 $X2=0 $Y2=0
cc_162 A2 N_A1_M1006_g 0.0156248f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_163 N_A2_M1001_g A1 2.22272e-19 $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A2_c_196_n A1 0.0111965f $X=2.51 $Y=1.925 $X2=0 $Y2=0
cc_165 N_A2_c_197_n A1 0.00732665f $X=3.63 $Y=1.925 $X2=0 $Y2=0
cc_166 N_A2_c_198_n A1 3.01865e-19 $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_167 N_A2_c_199_n A1 0.0125605f $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_168 N_A2_c_200_n A1 0.0165705f $X=3.895 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A2_c_201_n A1 2.41291e-19 $X=3.895 $Y=1.51 $X2=0 $Y2=0
cc_170 A2 A1 0.0331228f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_171 N_A2_c_196_n N_A1_c_290_n 2.41156e-19 $X=2.51 $Y=1.925 $X2=0 $Y2=0
cc_172 N_A2_c_197_n N_A1_c_290_n 0.00519784f $X=3.63 $Y=1.925 $X2=0 $Y2=0
cc_173 N_A2_c_198_n N_A1_c_290_n 0.0225706f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_174 N_A2_c_199_n N_A1_c_290_n 5.76239e-19 $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_175 N_A2_c_200_n N_A1_c_290_n 0.00434328f $X=3.895 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A2_c_201_n N_A1_c_290_n 0.0285162f $X=3.895 $Y=1.51 $X2=0 $Y2=0
cc_177 A2 N_A1_c_290_n 9.29551e-19 $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_178 N_A2_c_196_n N_VPWR_M1001_d 0.00229751f $X=2.51 $Y=1.925 $X2=0 $Y2=0
cc_179 A2 N_VPWR_M1001_d 0.0109043f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_180 N_A2_c_197_n N_VPWR_M1006_d 0.0027396f $X=3.63 $Y=1.925 $X2=0 $Y2=0
cc_181 A2 N_VPWR_M1006_d 3.46473e-19 $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_182 N_A2_M1001_g N_VPWR_c_347_n 0.00593682f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A2_M1008_g N_VPWR_c_348_n 0.0120491f $X=3.805 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A2_M1001_g N_VPWR_c_349_n 0.00532251f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A2_M1008_g N_VPWR_c_351_n 0.00486043f $X=3.805 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A2_M1001_g N_VPWR_c_344_n 0.00990847f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A2_M1008_g N_VPWR_c_344_n 0.00921558f $X=3.805 $Y=2.465 $X2=0 $Y2=0
cc_188 A2 N_A_231_367#_M1000_s 0.00336231f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_189 N_A2_M1001_g N_A_231_367#_c_413_n 0.00217191f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A2_M1001_g N_A_231_367#_c_404_n 3.19814e-19 $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A2_c_196_n N_A_231_367#_c_404_n 0.00319111f $X=2.51 $Y=1.925 $X2=0
+ $Y2=0
cc_192 N_A2_M1001_g N_A_231_367#_c_420_n 0.00734737f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_A2_M1001_g N_A_231_367#_c_421_n 0.0142247f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_A2_c_196_n N_A_231_367#_c_421_n 0.00889332f $X=2.51 $Y=1.925 $X2=0
+ $Y2=0
cc_195 N_A2_c_198_n N_A_231_367#_c_421_n 3.70402e-19 $X=2.415 $Y=1.51 $X2=0
+ $Y2=0
cc_196 A2 N_A_231_367#_c_421_n 0.0238056f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_197 N_A2_M1001_g N_A_231_367#_c_425_n 6.36091e-19 $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A2_M1008_g N_A_231_367#_c_426_n 0.0141605f $X=3.805 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A2_c_197_n N_A_231_367#_c_426_n 0.0135138f $X=3.63 $Y=1.925 $X2=0 $Y2=0
cc_200 N_A2_c_200_n N_A_231_367#_c_426_n 0.00358451f $X=3.895 $Y=1.51 $X2=0
+ $Y2=0
cc_201 A2 N_A_231_367#_c_426_n 0.0107917f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_202 N_A2_M1008_g N_A_231_367#_c_405_n 0.00201949f $X=3.805 $Y=2.465 $X2=0
+ $Y2=0
cc_203 N_A2_c_197_n N_A_231_367#_c_405_n 0.00463659f $X=3.63 $Y=1.925 $X2=0
+ $Y2=0
cc_204 N_A2_c_200_n N_A_231_367#_c_405_n 0.0120338f $X=3.895 $Y=1.51 $X2=0 $Y2=0
cc_205 N_A2_c_201_n N_A_231_367#_c_405_n 0.00347745f $X=3.895 $Y=1.51 $X2=0
+ $Y2=0
cc_206 N_A2_M1001_g N_A_231_367#_c_434_n 0.00230939f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_207 A2 N_A_231_367#_c_435_n 0.0162808f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_208 N_A2_M1009_g N_Y_c_466_n 0.0147359f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_209 N_A2_M1013_g N_Y_c_466_n 3.20368e-19 $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_210 N_A2_c_198_n N_Y_c_466_n 0.00474835f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_211 N_A2_c_199_n N_Y_c_466_n 0.0231284f $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_212 N_A2_c_196_n Y 2.72222e-19 $X=2.51 $Y=1.925 $X2=0 $Y2=0
cc_213 N_A2_M1009_g Y 2.86632e-19 $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_214 N_A2_c_196_n Y 0.00607868f $X=2.51 $Y=1.925 $X2=0 $Y2=0
cc_215 N_A2_c_198_n Y 3.69884e-19 $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_216 N_A2_c_199_n Y 0.00623774f $X=2.51 $Y=1.51 $X2=0 $Y2=0
cc_217 N_A2_M1009_g N_VGND_c_523_n 0.00524298f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_218 N_A2_M1013_g N_VGND_c_525_n 0.00783332f $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_219 N_A2_c_200_n N_VGND_c_525_n 0.0141273f $X=3.895 $Y=1.51 $X2=0 $Y2=0
cc_220 N_A2_c_201_n N_VGND_c_525_n 0.00398458f $X=3.895 $Y=1.51 $X2=0 $Y2=0
cc_221 N_A2_M1009_g N_VGND_c_528_n 0.00466948f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_222 N_A2_M1013_g N_VGND_c_528_n 0.00499542f $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_223 N_A2_M1009_g N_VGND_c_531_n 0.00896985f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_224 N_A2_M1013_g N_VGND_c_531_n 0.0100884f $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_225 N_A2_M1009_g N_A_502_65#_c_582_n 0.00524231f $X=2.435 $Y=0.745 $X2=0
+ $Y2=0
cc_226 N_A2_M1013_g N_A_502_65#_c_579_n 5.28944e-19 $X=3.805 $Y=0.745 $X2=0
+ $Y2=0
cc_227 N_A2_M1009_g N_A_502_65#_c_580_n 0.00264416f $X=2.435 $Y=0.745 $X2=0
+ $Y2=0
cc_228 N_A2_M1013_g N_A_502_65#_c_581_n 8.9451e-19 $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_229 N_A2_c_200_n N_A_502_65#_c_581_n 0.017881f $X=3.895 $Y=1.51 $X2=0 $Y2=0
cc_230 N_A1_M1000_g N_VPWR_c_347_n 0.00451811f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A1_M1000_g N_VPWR_c_348_n 7.72556e-19 $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A1_M1006_g N_VPWR_c_348_n 0.0114585f $X=3.375 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A1_M1000_g N_VPWR_c_350_n 0.00538529f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A1_M1006_g N_VPWR_c_350_n 0.00486043f $X=3.375 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A1_M1000_g N_VPWR_c_344_n 0.0100061f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A1_M1006_g N_VPWR_c_344_n 0.00835506f $X=3.375 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A1_M1000_g N_A_231_367#_c_420_n 6.23203e-19 $X=2.945 $Y=2.465 $X2=0
+ $Y2=0
cc_238 N_A1_M1000_g N_A_231_367#_c_421_n 0.0111411f $X=2.945 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A1_M1000_g N_A_231_367#_c_425_n 0.00822731f $X=2.945 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_A1_M1006_g N_A_231_367#_c_426_n 0.0122129f $X=3.375 $Y=2.465 $X2=0
+ $Y2=0
cc_241 N_A1_M1000_g N_A_231_367#_c_435_n 0.00102264f $X=2.945 $Y=2.465 $X2=0
+ $Y2=0
cc_242 N_A1_M1003_g N_Y_c_466_n 0.0127523f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_243 N_A1_M1005_g N_Y_c_466_n 0.00414996f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_244 A1 N_Y_c_466_n 0.0397651f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_245 N_A1_c_290_n N_Y_c_466_n 0.00492218f $X=3.375 $Y=1.51 $X2=0 $Y2=0
cc_246 N_A1_M1005_g N_Y_c_502_n 0.00506691f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_247 N_A1_M1003_g N_VGND_c_528_n 0.00304113f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_248 N_A1_M1005_g N_VGND_c_528_n 0.0030414f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_249 N_A1_M1003_g N_VGND_c_531_n 0.00443262f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_250 N_A1_M1005_g N_VGND_c_531_n 0.00443266f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_251 N_A1_M1003_g N_A_502_65#_c_582_n 0.00676031f $X=2.865 $Y=0.745 $X2=0
+ $Y2=0
cc_252 N_A1_M1005_g N_A_502_65#_c_582_n 5.37284e-19 $X=3.375 $Y=0.745 $X2=0
+ $Y2=0
cc_253 N_A1_M1003_g N_A_502_65#_c_579_n 0.00875863f $X=2.865 $Y=0.745 $X2=0
+ $Y2=0
cc_254 N_A1_M1005_g N_A_502_65#_c_579_n 0.0122692f $X=3.375 $Y=0.745 $X2=0 $Y2=0
cc_255 N_A1_M1003_g N_A_502_65#_c_580_n 0.00124108f $X=2.865 $Y=0.745 $X2=0
+ $Y2=0
cc_256 N_A1_M1005_g N_A_502_65#_c_581_n 8.30663e-19 $X=3.375 $Y=0.745 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_344_n N_A_231_367#_M1004_d 0.00215161f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_258 N_VPWR_c_344_n N_A_231_367#_M1010_d 0.00223562f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_344_n N_A_231_367#_M1000_s 0.0039448f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_344_n N_A_231_367#_M1008_s 0.00371702f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_346_n N_A_231_367#_c_402_n 0.00532082f $X=0.305 $Y=2.765 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_349_n N_A_231_367#_c_402_n 0.0179183f $X=2.485 $Y=3.33 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_344_n N_A_231_367#_c_402_n 0.0101029f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_346_n N_A_231_367#_c_403_n 8.29431e-19 $X=0.305 $Y=2.765 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_349_n N_A_231_367#_c_413_n 0.0525906f $X=2.485 $Y=3.33 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_344_n N_A_231_367#_c_413_n 0.0339238f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_267 N_VPWR_M1001_d N_A_231_367#_c_421_n 0.00765266f $X=2.43 $Y=1.835 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_347_n N_A_231_367#_c_421_n 0.0254128f $X=2.65 $Y=2.78 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_350_n N_A_231_367#_c_425_n 0.00976751f $X=3.425 $Y=3.33 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_344_n N_A_231_367#_c_425_n 0.00966132f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_271 N_VPWR_M1006_d N_A_231_367#_c_426_n 0.0035188f $X=3.45 $Y=1.835 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_348_n N_A_231_367#_c_426_n 0.0170777f $X=3.59 $Y=2.765 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_351_n N_A_231_367#_c_406_n 0.0178111f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_344_n N_A_231_367#_c_406_n 0.0100304f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_344_n N_Y_M1004_s 0.00225186f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_276 N_A_231_367#_c_413_n N_Y_M1004_s 0.00334491f $X=2.045 $Y=2.99 $X2=0 $Y2=0
cc_277 N_A_231_367#_c_404_n N_Y_c_466_n 0.0070672f $X=2.14 $Y=1.995 $X2=0 $Y2=0
cc_278 N_A_231_367#_c_403_n Y 0.0338931f $X=1.28 $Y=1.995 $X2=0 $Y2=0
cc_279 N_A_231_367#_c_404_n Y 0.017377f $X=2.14 $Y=1.995 $X2=0 $Y2=0
cc_280 N_A_231_367#_c_413_n Y 0.0155817f $X=2.045 $Y=2.99 $X2=0 $Y2=0
cc_281 N_A_231_367#_c_403_n N_VGND_c_522_n 0.0074605f $X=1.28 $Y=1.995 $X2=0
+ $Y2=0
cc_282 N_A_231_367#_c_405_n N_VGND_c_525_n 0.00463729f $X=4.02 $Y=1.98 $X2=0
+ $Y2=0
cc_283 N_Y_c_466_n N_VGND_M1007_s 0.00261503f $X=2.995 $Y=1.16 $X2=0 $Y2=0
cc_284 Y N_VGND_c_522_n 0.00416299f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_285 N_Y_c_467_n N_VGND_c_522_n 0.0301083f $X=1.71 $Y=0.45 $X2=0 $Y2=0
cc_286 N_Y_c_466_n N_VGND_c_523_n 0.0218003f $X=2.995 $Y=1.16 $X2=0 $Y2=0
cc_287 N_Y_c_467_n N_VGND_c_523_n 0.0248289f $X=1.71 $Y=0.45 $X2=0 $Y2=0
cc_288 N_Y_c_467_n N_VGND_c_527_n 0.0154596f $X=1.71 $Y=0.45 $X2=0 $Y2=0
cc_289 N_Y_c_467_n N_VGND_c_531_n 0.00977127f $X=1.71 $Y=0.45 $X2=0 $Y2=0
cc_290 N_Y_c_466_n N_A_502_65#_M1009_d 0.00176461f $X=2.995 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_291 N_Y_c_466_n N_A_502_65#_c_582_n 0.0169932f $X=2.995 $Y=1.16 $X2=0 $Y2=0
cc_292 N_Y_M1003_d N_A_502_65#_c_579_n 0.00261503f $X=2.94 $Y=0.325 $X2=0 $Y2=0
cc_293 N_Y_c_466_n N_A_502_65#_c_579_n 0.00280043f $X=2.995 $Y=1.16 $X2=0 $Y2=0
cc_294 N_Y_c_502_n N_A_502_65#_c_579_n 0.020345f $X=3.16 $Y=0.69 $X2=0 $Y2=0
cc_295 N_Y_c_466_n N_A_502_65#_c_581_n 0.00538273f $X=2.995 $Y=1.16 $X2=0 $Y2=0
cc_296 N_VGND_c_525_n N_A_502_65#_c_579_n 0.00517394f $X=4.02 $Y=0.47 $X2=0
+ $Y2=0
cc_297 N_VGND_c_528_n N_A_502_65#_c_579_n 0.0555626f $X=3.89 $Y=0 $X2=0 $Y2=0
cc_298 N_VGND_c_531_n N_A_502_65#_c_579_n 0.032853f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_299 N_VGND_c_523_n N_A_502_65#_c_580_n 0.00920528f $X=2.14 $Y=0.45 $X2=0
+ $Y2=0
cc_300 N_VGND_c_528_n N_A_502_65#_c_580_n 0.0219773f $X=3.89 $Y=0 $X2=0 $Y2=0
cc_301 N_VGND_c_531_n N_A_502_65#_c_580_n 0.0125175f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_302 N_VGND_c_525_n N_A_502_65#_c_581_n 0.0015231f $X=4.02 $Y=0.47 $X2=0 $Y2=0
