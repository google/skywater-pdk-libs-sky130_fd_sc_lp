* File: sky130_fd_sc_lp__or4_m.spice
* Created: Wed Sep  2 10:32:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4_m.pex.spice"
.subckt sky130_fd_sc_lp__or4_m  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1006 N_A_116_397#_M1006_d N_D_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_C_M1009_g N_A_116_397#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1344 AS=0.0588 PD=1.06 PS=0.7 NRD=102.852 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1001 N_A_116_397#_M1001_d N_B_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1344 PD=0.7 PS=1.06 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_116_397#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0966 AS=0.0588 PD=0.88 PS=0.7 NRD=28.56 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_116_397#_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0966 PD=1.37 PS=0.88 NRD=0 NRS=22.848 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_199_397# N_D_M1003_g N_A_116_397#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1002 A_271_397# N_C_M1002_g A_199_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1005 A_343_397# N_B_M1005_g A_271_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.9
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_343_397# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.12495 AS=0.0441 PD=1.015 PS=0.63 NRD=110.222 NRS=23.443 M=1 R=2.8
+ SA=75001.3 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1008 N_X_M1008_d N_A_116_397#_M1008_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.12495 PD=1.37 PS=1.015 NRD=0 NRS=37.5088 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__or4_m.pxi.spice"
*
.ends
*
*
