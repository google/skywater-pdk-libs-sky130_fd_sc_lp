* File: sky130_fd_sc_lp__nor4b_lp.pex.spice
* Created: Wed Sep  2 10:11:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4B_LP%D_N 2 5 7 9 12 14 16 17 18 19 20 24 26
c52 2 0 7.95967e-20 $X=0.627 $Y=1.658
r53 24 26 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.627 $Y=1.34
+ $X2=0.627 $Y2=1.175
r54 19 20 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.66 $Y=1.295
+ $X2=0.66 $Y2=1.665
r55 19 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.65
+ $Y=1.34 $X2=0.65 $Y2=1.34
r56 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.005 $Y=0.78
+ $X2=1.005 $Y2=0.495
r57 13 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.72 $Y=0.855
+ $X2=0.645 $Y2=0.855
r58 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.93 $Y=0.855
+ $X2=1.005 $Y2=0.78
r59 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.93 $Y=0.855
+ $X2=0.72 $Y2=0.855
r60 10 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.645 $Y=0.93
+ $X2=0.645 $Y2=0.855
r61 10 26 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=0.645 $Y=0.93
+ $X2=0.645 $Y2=1.175
r62 7 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.645 $Y=0.78
+ $X2=0.645 $Y2=0.855
r63 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.645 $Y=0.78 $X2=0.645
+ $Y2=0.495
r64 5 17 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.565 $Y=2.545
+ $X2=0.565 $Y2=1.845
r65 2 17 33.9275 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.627 $Y=1.658
+ $X2=0.627 $Y2=1.845
r66 1 24 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.627 $Y=1.362
+ $X2=0.627 $Y2=1.34
r67 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.627 $Y=1.362
+ $X2=0.627 $Y2=1.658
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_LP%A_31_409# 1 2 8 11 13 14 17 19 21 23 24 27
+ 33 35 37 41 42 44 45
r83 42 47 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.282 $Y=1.34
+ $X2=1.282 $Y2=1.175
r84 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.22
+ $Y=1.34 $X2=1.22 $Y2=1.34
r85 39 41 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.22 $Y=0.995
+ $X2=1.22 $Y2=1.34
r86 38 44 3.63293 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.595 $Y=0.91
+ $X2=0.365 $Y2=0.91
r87 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.055 $Y=0.91
+ $X2=1.22 $Y2=0.995
r88 37 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.055 $Y=0.91
+ $X2=0.595 $Y2=0.91
r89 33 45 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.3 $Y=2.19 $X2=0.3
+ $Y2=2.025
r90 33 35 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.3 $Y=2.19 $X2=0.3
+ $Y2=2.9
r91 29 44 3.01263 $w=3.15e-07 $l=1.8262e-07 $layer=LI1_cond $X=0.22 $Y=0.995
+ $X2=0.365 $Y2=0.91
r92 29 45 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.22 $Y=0.995
+ $X2=0.22 $Y2=2.025
r93 25 44 3.01263 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.365 $Y=0.825
+ $X2=0.365 $Y2=0.91
r94 25 27 8.58056 $w=4.58e-07 $l=3.3e-07 $layer=LI1_cond $X=0.365 $Y=0.825
+ $X2=0.365 $Y2=0.495
r95 21 23 117.608 $w=2.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.56 $Y=1.935
+ $X2=2.56 $Y2=2.545
r96 20 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.9 $Y=1.86
+ $X2=1.825 $Y2=1.86
r97 19 21 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=2.435 $Y=1.86
+ $X2=2.56 $Y2=1.935
r98 19 20 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.435 $Y=1.86
+ $X2=1.9 $Y2=1.86
r99 15 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.825 $Y=1.785
+ $X2=1.825 $Y2=1.86
r100 15 17 661.468 $w=1.5e-07 $l=1.29e-06 $layer=POLY_cond $X=1.825 $Y=1.785
+ $X2=1.825 $Y2=0.495
r101 13 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=1.86
+ $X2=1.825 $Y2=1.86
r102 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.75 $Y=1.86
+ $X2=1.51 $Y2=1.86
r103 11 47 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.435 $Y=0.495
+ $X2=1.435 $Y2=1.175
r104 8 14 36.9868 $w=1.5e-07 $l=2.62838e-07 $layer=POLY_cond $X=1.282 $Y=1.785
+ $X2=1.51 $Y2=1.86
r105 7 42 7.57836 $w=4.55e-07 $l=6.2e-08 $layer=POLY_cond $X=1.282 $Y=1.402
+ $X2=1.282 $Y2=1.34
r106 7 8 46.8147 $w=4.55e-07 $l=3.83e-07 $layer=POLY_cond $X=1.282 $Y=1.402
+ $X2=1.282 $Y2=1.785
r107 2 35 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=2.045 $X2=0.3 $Y2=2.9
r108 2 33 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=2.045 $X2=0.3 $Y2=2.19
r109 1 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.285
+ $Y=0.285 $X2=0.43 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_LP%C 3 5 6 9 13 15 16 17 18 33 34
c50 13 0 6.63748e-20 $X=3.05 $Y=2.545
r51 33 35 50.8532 $w=3.27e-07 $l=3.45e-07 $layer=POLY_cond $X=2.705 $Y=1.442
+ $X2=3.05 $Y2=1.442
r52 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=1.38 $X2=2.705 $Y2=1.38
r53 31 33 13.2661 $w=3.27e-07 $l=9e-08 $layer=POLY_cond $X=2.615 $Y=1.442
+ $X2=2.705 $Y2=1.442
r54 17 18 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=2.405
+ $X2=2.88 $Y2=2.775
r55 16 17 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=2.035
+ $X2=2.88 $Y2=2.405
r56 15 16 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=2.035
r57 15 34 4.80116 $w=7.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=1.38
r58 11 35 9.13417 $w=2.5e-07 $l=2.28e-07 $layer=POLY_cond $X=3.05 $Y=1.67
+ $X2=3.05 $Y2=1.442
r59 11 13 217.397 $w=2.5e-07 $l=8.75e-07 $layer=POLY_cond $X=3.05 $Y=1.67
+ $X2=3.05 $Y2=2.545
r60 7 31 21.0057 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=2.615 $Y=1.215
+ $X2=2.615 $Y2=1.442
r61 7 9 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.615 $Y=1.215
+ $X2=2.615 $Y2=0.495
r62 5 31 25.3157 $w=3.27e-07 $l=1.85753e-07 $layer=POLY_cond $X=2.54 $Y=1.29
+ $X2=2.615 $Y2=1.442
r63 5 6 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.54 $Y=1.29 $X2=2.33
+ $Y2=1.29
r64 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.255 $Y=1.215
+ $X2=2.33 $Y2=1.29
r65 1 3 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.255 $Y=1.215
+ $X2=2.255 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_LP%B 1 3 4 5 6 8 13 15 17 18 19 20 21 22 23 29
+ 30
c61 15 0 5.91563e-20 $X=3.49 $Y=0.855
r62 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.58
+ $Y=1.38 $X2=3.58 $Y2=1.38
r63 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.58 $Y=2.405
+ $X2=3.58 $Y2=2.775
r64 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.58 $Y=2.035
+ $X2=3.58 $Y2=2.405
r65 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.58 $Y=1.665
+ $X2=3.58 $Y2=2.035
r66 20 30 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.58 $Y=1.665
+ $X2=3.58 $Y2=1.38
r67 18 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.58 $Y=1.72
+ $X2=3.58 $Y2=1.38
r68 18 19 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.72
+ $X2=3.58 $Y2=1.885
r69 17 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.215
+ $X2=3.58 $Y2=1.38
r70 13 19 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.54 $Y=2.545
+ $X2=3.54 $Y2=1.885
r71 9 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=0.93 $X2=3.49
+ $Y2=0.855
r72 9 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.49 $Y=0.93
+ $X2=3.49 $Y2=1.215
r73 6 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=0.78 $X2=3.49
+ $Y2=0.855
r74 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.49 $Y=0.78 $X2=3.49
+ $Y2=0.495
r75 4 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.415 $Y=0.855
+ $X2=3.49 $Y2=0.855
r76 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.415 $Y=0.855
+ $X2=3.205 $Y2=0.855
r77 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.13 $Y=0.78
+ $X2=3.205 $Y2=0.855
r78 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.13 $Y=0.78 $X2=3.13
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_LP%A 1 3 6 8 11 14 16 17 18 20 27
c37 20 0 5.91563e-20 $X=4.56 $Y=1.665
r38 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.19
+ $Y=1.07 $X2=4.19 $Y2=1.07
r39 20 28 5.15886 $w=8.73e-07 $l=3.7e-07 $layer=LI1_cond $X=4.56 $Y=1.342
+ $X2=4.19 $Y2=1.342
r40 18 28 1.53371 $w=8.73e-07 $l=1.1e-07 $layer=LI1_cond $X=4.08 $Y=1.342
+ $X2=4.19 $Y2=1.342
r41 16 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.06 $Y=1.575
+ $X2=4.06 $Y2=1.815
r42 15 27 49.9064 $w=3.7e-07 $l=3.2e-07 $layer=POLY_cond $X=4.17 $Y=1.39
+ $X2=4.17 $Y2=1.07
r43 15 16 49.8761 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.17 $Y=1.39
+ $X2=4.17 $Y2=1.575
r44 14 27 14.8159 $w=3.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.17 $Y=0.975
+ $X2=4.17 $Y2=1.07
r45 6 17 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.11 $Y=1.94
+ $X2=4.11 $Y2=1.815
r46 6 8 116.644 $w=2.5e-07 $l=6.05e-07 $layer=POLY_cond $X=4.11 $Y=1.94 $X2=4.11
+ $Y2=2.545
r47 1 14 25.6283 $w=3.7e-07 $l=1.5e-07 $layer=POLY_cond $X=4.1 $Y=0.825 $X2=4.1
+ $Y2=0.975
r48 1 11 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.28 $Y=0.825 $X2=4.28
+ $Y2=0.495
r49 1 3 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.92 $Y=0.825 $X2=3.92
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_LP%VPWR 1 2 11 15 17 21 23 32 36
r35 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r36 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 30 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r38 29 30 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r39 27 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 26 29 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r41 26 27 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 24 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.83 $Y2=3.33
r43 24 26 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 23 35 4.4922 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.21 $Y=3.33
+ $X2=4.505 $Y2=3.33
r45 23 29 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.21 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 21 30 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=4.08 $Y2=3.33
r47 21 27 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 17 20 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.375 $Y=2.19
+ $X2=4.375 $Y2=2.9
r49 15 35 3.27398 $w=3.3e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.375 $Y=3.245
+ $X2=4.505 $Y2=3.33
r50 15 20 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.375 $Y=3.245
+ $X2=4.375 $Y2=2.9
r51 11 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.83 $Y=2.19 $X2=0.83
+ $Y2=2.9
r52 9 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=3.245 $X2=0.83
+ $Y2=3.33
r53 9 14 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.83 $Y=3.245
+ $X2=0.83 $Y2=2.9
r54 2 20 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.235
+ $Y=2.045 $X2=4.375 $Y2=2.9
r55 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.235
+ $Y=2.045 $X2=4.375 $Y2=2.19
r56 1 14 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=2.045 $X2=0.83 $Y2=2.9
r57 1 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=2.045 $X2=0.83 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_LP%Y 1 2 3 10 13 15 18 19 20 21 22 23 24 46
c59 20 0 6.63748e-20 $X=2.16 $Y=1.295
r60 46 75 1.51047 $w=7.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.035
+ $X2=1.955 $Y2=0.95
r61 24 65 1.91679 $w=7.78e-07 $l=1.25e-07 $layer=LI1_cond $X=1.955 $Y=2.775
+ $X2=1.955 $Y2=2.9
r62 23 24 5.67371 $w=7.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.955 $Y=2.405
+ $X2=1.955 $Y2=2.775
r63 23 57 3.29688 $w=7.78e-07 $l=2.15e-07 $layer=LI1_cond $X=1.955 $Y=2.405
+ $X2=1.955 $Y2=2.19
r64 22 57 2.37682 $w=7.78e-07 $l=1.55e-07 $layer=LI1_cond $X=1.955 $Y=2.035
+ $X2=1.955 $Y2=2.19
r65 21 22 5.67371 $w=7.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.955 $Y=1.665
+ $X2=1.955 $Y2=2.035
r66 20 21 5.67371 $w=7.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.955 $Y=1.295
+ $X2=1.955 $Y2=1.665
r67 20 46 3.98693 $w=7.78e-07 $l=2.6e-07 $layer=LI1_cond $X=1.955 $Y=1.295
+ $X2=1.955 $Y2=1.035
r68 19 75 0.440115 $w=6.93e-07 $l=2.5e-08 $layer=LI1_cond $X=1.955 $Y=0.925
+ $X2=1.955 $Y2=0.95
r69 18 19 6.51371 $w=6.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.955 $Y=0.555
+ $X2=1.955 $Y2=0.925
r70 18 68 1.05628 $w=6.93e-07 $l=6e-08 $layer=LI1_cond $X=1.955 $Y=0.555
+ $X2=1.955 $Y2=0.495
r71 15 17 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.705 $Y=0.495
+ $X2=3.705 $Y2=0.725
r72 13 17 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.625 $Y=0.865
+ $X2=3.625 $Y2=0.725
r73 11 75 9.25536 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=2.345 $Y=0.95
+ $X2=1.955 $Y2=0.95
r74 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.54 $Y=0.95
+ $X2=3.625 $Y2=0.865
r75 10 11 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=3.54 $Y=0.95
+ $X2=2.345 $Y2=0.95
r76 3 65 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.035
+ $Y=2.045 $X2=2.18 $Y2=2.9
r77 3 57 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.035
+ $Y=2.045 $X2=2.18 $Y2=2.19
r78 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.565
+ $Y=0.285 $X2=3.705 $Y2=0.495
r79 1 68 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.9
+ $Y=0.285 $X2=2.04 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_LP%VGND 1 2 3 12 16 18 20 23 24 25 27 39 47 51
r57 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r58 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r60 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r61 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r62 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r63 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r64 39 50 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.565
+ $Y2=0
r65 39 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.08
+ $Y2=0
r66 38 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r67 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 35 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r69 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r70 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r71 32 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r72 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r73 30 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r74 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r75 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r76 27 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.72
+ $Y2=0
r77 25 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r78 25 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r79 23 37 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.665 $Y=0 $X2=2.64
+ $Y2=0
r80 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.665 $Y=0 $X2=2.83
+ $Y2=0
r81 22 41 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.995 $Y=0 $X2=3.12
+ $Y2=0
r82 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.995 $Y=0 $X2=2.83
+ $Y2=0
r83 18 50 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=4.495 $Y=0.085
+ $X2=4.565 $Y2=0
r84 18 20 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.495 $Y=0.085
+ $X2=4.495 $Y2=0.495
r85 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.83 $Y=0.085
+ $X2=2.83 $Y2=0
r86 14 16 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.83 $Y=0.085
+ $X2=2.83 $Y2=0.475
r87 10 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r88 10 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.455
r89 3 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.285 $X2=4.495 $Y2=0.495
r90 2 16 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=2.69
+ $Y=0.285 $X2=2.83 $Y2=0.475
r91 1 12 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.285 $X2=1.22 $Y2=0.455
.ends

