# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand2_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nand2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.430000 1.425000 5.780000 1.760000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.415000 3.505000 1.595000 ;
        RECT 1.815000 1.595000 3.505000 1.605000 ;
        RECT 1.815000 1.605000 2.825000 1.760000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  3.973200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.765000 1.635000 1.930000 ;
        RECT 0.595000 1.930000 6.185000 1.935000 ;
        RECT 0.595000 1.935000 0.785000 3.075000 ;
        RECT 1.455000 1.935000 6.185000 1.945000 ;
        RECT 1.455000 1.945000 3.365000 2.100000 ;
        RECT 1.455000 2.100000 1.645000 3.075000 ;
        RECT 2.315000 2.100000 2.505000 3.075000 ;
        RECT 3.125000 1.775000 4.260000 1.930000 ;
        RECT 3.175000 2.100000 3.365000 3.075000 ;
        RECT 3.965000 0.595000 4.295000 1.085000 ;
        RECT 3.965000 1.085000 6.220000 1.155000 ;
        RECT 3.965000 1.155000 7.115000 1.255000 ;
        RECT 3.965000 1.255000 4.260000 1.775000 ;
        RECT 4.035000 1.945000 6.185000 2.100000 ;
        RECT 4.035000 2.100000 4.260000 3.075000 ;
        RECT 4.930000 2.100000 5.260000 3.075000 ;
        RECT 4.965000 0.595000 5.295000 1.075000 ;
        RECT 4.965000 1.075000 6.220000 1.085000 ;
        RECT 5.950000 1.255000 7.115000 1.500000 ;
        RECT 5.950000 1.500000 7.055000 1.925000 ;
        RECT 5.950000 1.925000 6.185000 1.930000 ;
        RECT 5.950000 2.100000 6.185000 3.075000 ;
        RECT 5.965000 0.605000 6.220000 1.075000 ;
        RECT 6.785000 0.605000 7.115000 1.155000 ;
        RECT 6.855000 1.925000 7.055000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.095000  0.305000 0.355000 1.075000 ;
      RECT 0.095000  1.075000 3.795000 1.245000 ;
      RECT 0.095000  1.820000 0.425000 3.245000 ;
      RECT 0.525000  0.085000 0.855000 0.905000 ;
      RECT 0.955000  2.105000 1.285000 3.245000 ;
      RECT 1.025000  0.305000 1.205000 1.075000 ;
      RECT 1.385000  0.085000 1.715000 0.905000 ;
      RECT 1.815000  2.270000 2.145000 3.245000 ;
      RECT 1.885000  0.305000 2.075000 1.075000 ;
      RECT 2.245000  0.085000 2.575000 0.905000 ;
      RECT 2.675000  2.270000 3.005000 3.245000 ;
      RECT 2.745000  0.305000 2.935000 1.075000 ;
      RECT 3.105000  0.085000 3.435000 0.905000 ;
      RECT 3.535000  2.115000 3.865000 3.245000 ;
      RECT 3.605000  0.255000 7.545000 0.425000 ;
      RECT 3.605000  0.425000 3.795000 1.075000 ;
      RECT 4.430000  2.270000 4.760000 3.245000 ;
      RECT 4.465000  0.425000 4.795000 0.915000 ;
      RECT 5.430000  2.270000 5.760000 3.245000 ;
      RECT 5.465000  0.425000 7.545000 0.435000 ;
      RECT 5.465000  0.435000 5.795000 0.905000 ;
      RECT 6.355000  2.095000 6.685000 3.245000 ;
      RECT 6.390000  0.435000 6.615000 0.985000 ;
      RECT 7.275000  1.815000 7.485000 3.245000 ;
      RECT 7.285000  0.435000 7.545000 1.190000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__nand2_8
