* File: sky130_fd_sc_lp__o22ai_lp.spice
* Created: Wed Sep  2 10:20:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22ai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o22ai_lp  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_70_101#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1533 PD=0.7 PS=1.57 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.3
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1004 N_A_70_101#_M1004_d N_B2_M1004_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_70_101#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1491 AS=0.0756 PD=1.13 PS=0.78 NRD=47.136 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_70_101#_M1002_d N_A1_M1002_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1491 PD=1.41 PS=1.13 NRD=0 NRS=75.708 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_169_419# N_B1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g A_169_419# VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.12 PD=1.32 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1006 A_381_419# N_A2_M1006_g N_Y_M1000_d VPB PHIGHVT L=0.25 W=1 AD=0.305
+ AS=0.16 PD=1.61 PS=1.32 NRD=49.2303 NRS=7.8603 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_381_419# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.305 PD=2.57 PS=1.61 NRD=0 NRS=49.2303 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o22ai_lp.pxi.spice"
*
.ends
*
*
