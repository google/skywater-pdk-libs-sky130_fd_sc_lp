* File: sky130_fd_sc_lp__o41a_0.pxi.spice
* Created: Fri Aug 28 11:19:00 2020
* 
x_PM_SKY130_FD_SC_LP__O41A_0%A_80_21# N_A_80_21#_M1007_s N_A_80_21#_M1005_d
+ N_A_80_21#_M1003_g N_A_80_21#_c_90_n N_A_80_21#_M1010_g N_A_80_21#_c_92_n
+ N_A_80_21#_c_93_n N_A_80_21#_c_94_n N_A_80_21#_c_95_n N_A_80_21#_c_96_n
+ N_A_80_21#_c_101_n N_A_80_21#_c_102_n N_A_80_21#_c_97_n N_A_80_21#_c_103_n
+ N_A_80_21#_c_104_n N_A_80_21#_c_98_n PM_SKY130_FD_SC_LP__O41A_0%A_80_21#
x_PM_SKY130_FD_SC_LP__O41A_0%B1 N_B1_M1005_g N_B1_M1007_g N_B1_c_164_n
+ N_B1_c_165_n B1 B1 N_B1_c_167_n PM_SKY130_FD_SC_LP__O41A_0%B1
x_PM_SKY130_FD_SC_LP__O41A_0%A4 N_A4_c_210_n N_A4_M1009_g N_A4_M1006_g
+ N_A4_c_212_n N_A4_c_216_n A4 A4 A4 PM_SKY130_FD_SC_LP__O41A_0%A4
x_PM_SKY130_FD_SC_LP__O41A_0%A3 N_A3_M1000_g N_A3_c_263_n N_A3_M1008_g
+ N_A3_c_265_n A3 A3 A3 A3 A3 N_A3_c_262_n A3 PM_SKY130_FD_SC_LP__O41A_0%A3
x_PM_SKY130_FD_SC_LP__O41A_0%A2 N_A2_c_314_n N_A2_M1004_g N_A2_M1011_g
+ N_A2_c_315_n N_A2_c_316_n N_A2_c_317_n N_A2_c_322_n A2 A2 A2 A2 A2
+ N_A2_c_319_n PM_SKY130_FD_SC_LP__O41A_0%A2
x_PM_SKY130_FD_SC_LP__O41A_0%A1 N_A1_M1002_g N_A1_c_376_n N_A1_M1001_g
+ N_A1_c_371_n N_A1_c_372_n N_A1_c_378_n N_A1_c_373_n A1 A1 A1 N_A1_c_374_n
+ N_A1_c_375_n PM_SKY130_FD_SC_LP__O41A_0%A1
x_PM_SKY130_FD_SC_LP__O41A_0%X N_X_M1003_s N_X_M1010_s X X X X X X X N_X_c_408_n
+ X PM_SKY130_FD_SC_LP__O41A_0%X
x_PM_SKY130_FD_SC_LP__O41A_0%VPWR N_VPWR_M1010_d N_VPWR_M1001_d N_VPWR_c_425_n
+ N_VPWR_c_426_n N_VPWR_c_427_n VPWR N_VPWR_c_428_n N_VPWR_c_429_n
+ N_VPWR_c_424_n PM_SKY130_FD_SC_LP__O41A_0%VPWR
x_PM_SKY130_FD_SC_LP__O41A_0%VGND N_VGND_M1003_d N_VGND_M1009_d N_VGND_M1004_d
+ N_VGND_c_463_n N_VGND_c_464_n N_VGND_c_465_n VGND N_VGND_c_466_n
+ N_VGND_c_467_n N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n
+ N_VGND_c_472_n N_VGND_c_473_n PM_SKY130_FD_SC_LP__O41A_0%VGND
x_PM_SKY130_FD_SC_LP__O41A_0%A_319_51# N_A_319_51#_M1007_d N_A_319_51#_M1000_d
+ N_A_319_51#_M1002_d N_A_319_51#_c_519_n N_A_319_51#_c_520_n
+ N_A_319_51#_c_521_n N_A_319_51#_c_522_n N_A_319_51#_c_523_n
+ N_A_319_51#_c_524_n N_A_319_51#_c_525_n PM_SKY130_FD_SC_LP__O41A_0%A_319_51#
cc_1 VNB N_A_80_21#_c_90_n 0.0255823f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.248
cc_2 VNB N_A_80_21#_M1010_g 0.0126842f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.735
cc_3 VNB N_A_80_21#_c_92_n 0.0249134f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.435
cc_4 VNB N_A_80_21#_c_93_n 0.0035744f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.93
cc_5 VNB N_A_80_21#_c_94_n 0.022919f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.93
cc_6 VNB N_A_80_21#_c_95_n 0.0199243f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.825
cc_7 VNB N_A_80_21#_c_96_n 0.0019577f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.825
cc_8 VNB N_A_80_21#_c_97_n 0.00686921f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=0.465
cc_9 VNB N_A_80_21#_c_98_n 0.0223774f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=0.765
cc_10 VNB N_B1_M1007_g 0.0387087f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_11 VNB N_B1_c_164_n 0.0394909f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.435
cc_12 VNB N_B1_c_165_n 0.00554256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB B1 0.00307629f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.435
cc_14 VNB N_B1_c_167_n 0.0279677f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.93
cc_15 VNB N_A4_c_210_n 0.0335881f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=0.255
cc_16 VNB N_A4_M1009_g 0.0345784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A4_c_212_n 0.00121392f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=0.952
cc_18 VNB A4 0.0122268f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.435
cc_19 VNB N_A3_M1000_g 0.0552985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A3 0.00679558f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.435
cc_21 VNB N_A3_c_262_n 0.0125454f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=2.13
cc_22 VNB N_A2_c_314_n 0.0157893f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=0.255
cc_23 VNB N_A2_c_315_n 0.0171924f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.435
cc_24 VNB N_A2_c_316_n 0.0179534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A2_c_317_n 0.0158624f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.435
cc_26 VNB A2 0.00545533f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.045
cc_27 VNB N_A2_c_319_n 0.0163876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_M1002_g 0.0236936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A1_c_371_n 0.00176288f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_30 VNB N_A1_c_372_n 0.0387856f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.735
cc_31 VNB N_A1_c_373_n 0.0220464f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.93
cc_32 VNB N_A1_c_374_n 0.0481334f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=0.465
cc_33 VNB N_A1_c_375_n 0.00111806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_408_n 0.0674516f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=2.13
cc_35 VNB N_VPWR_c_424_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.317 $Y2=2.735
cc_36 VNB N_VGND_c_463_n 0.00709303f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.435
cc_37 VNB N_VGND_c_464_n 0.00530857f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.435
cc_38 VNB N_VGND_c_465_n 8.38565e-19 $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.93
cc_39 VNB N_VGND_c_466_n 0.0153306f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=2.13
cc_40 VNB N_VGND_c_467_n 0.0317031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_468_n 0.0148645f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=2.735
cc_42 VNB N_VGND_c_469_n 0.01735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_470_n 0.22235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_471_n 0.00510715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_472_n 0.00536127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_473_n 0.00460914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_319_51#_c_519_n 0.00210838f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.435
cc_48 VNB N_A_319_51#_c_520_n 0.00799154f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.735
cc_49 VNB N_A_319_51#_c_521_n 0.00398942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_319_51#_c_522_n 3.02314e-19 $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.045
cc_51 VNB N_A_319_51#_c_523_n 0.0123718f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.93
cc_52 VNB N_A_319_51#_c_524_n 0.0160869f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=2.13
cc_53 VNB N_A_319_51#_c_525_n 0.00403366f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=0.74
cc_54 VPB N_A_80_21#_M1010_g 0.0571079f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.735
cc_55 VPB N_A_80_21#_c_93_n 0.0070212f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.93
cc_56 VPB N_A_80_21#_c_101_n 0.0179027f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=2.13
cc_57 VPB N_A_80_21#_c_102_n 0.00396682f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=2.13
cc_58 VPB N_A_80_21#_c_103_n 0.00525465f $X=-0.19 $Y=1.655 $X2=1.317 $Y2=2.395
cc_59 VPB N_A_80_21#_c_104_n 0.0170794f $X=-0.19 $Y=1.655 $X2=1.825 $Y2=2.56
cc_60 VPB N_B1_M1005_g 0.0514368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_B1_c_165_n 0.0126313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB B1 0.00256015f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=1.435
cc_63 VPB N_A4_M1006_g 0.0306419f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_64 VPB N_A4_c_212_n 0.0212464f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=0.952
cc_65 VPB N_A4_c_216_n 0.0163166f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=1.248
cc_66 VPB A4 0.0173276f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.435
cc_67 VPB N_A3_c_263_n 0.0174887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A3_M1008_g 0.0216336f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_69 VPB N_A3_c_265_n 0.0208556f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=1.248
cc_70 VPB A3 0.00215221f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.435
cc_71 VPB A3 0.00125529f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A3_c_262_n 0.00277799f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=2.13
cc_73 VPB A3 0.00146039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A2_M1011_g 0.0342926f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_75 VPB N_A2_c_317_n 0.00580292f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=1.435
cc_76 VPB N_A2_c_322_n 0.0153238f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=0.91
cc_77 VPB A2 0.00564092f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.045
cc_78 VPB N_A1_c_376_n 0.0208272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A1_c_371_n 0.0318589f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_80 VPB N_A1_c_378_n 0.028933f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=0.91
cc_81 VPB N_A1_c_375_n 0.022765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_X_c_408_n 0.0395782f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=2.13
cc_83 VPB X 0.0425462f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=0.765
cc_84 VPB N_VPWR_c_425_n 0.0041898f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=1.248
cc_85 VPB N_VPWR_c_426_n 0.0130188f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.735
cc_86 VPB N_VPWR_c_427_n 0.0362773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_428_n 0.062527f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=0.93
cc_88 VPB N_VPWR_c_429_n 0.0246311f $X=-0.19 $Y=1.655 $X2=1.305 $Y2=0.465
cc_89 VPB N_VPWR_c_424_n 0.0786356f $X=-0.19 $Y=1.655 $X2=1.317 $Y2=2.735
cc_90 N_A_80_21#_c_101_n N_B1_M1005_g 0.0152254f $X=1.21 $Y=2.13 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_103_n N_B1_M1005_g 0.00724152f $X=1.317 $Y=2.395 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_104_n N_B1_M1005_g 8.7871e-19 $X=1.825 $Y=2.56 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_93_n N_B1_M1007_g 8.00885e-19 $X=0.61 $Y=0.93 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_94_n N_B1_M1007_g 0.00473976f $X=0.61 $Y=0.93 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_95_n N_B1_M1007_g 0.00260668f $X=1.14 $Y=0.825 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_97_n N_B1_M1007_g 0.00184158f $X=1.305 $Y=0.465 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_90_n N_B1_c_164_n 0.0094249f $X=0.587 $Y=1.248 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_93_n N_B1_c_164_n 0.00136741f $X=0.61 $Y=0.93 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_95_n N_B1_c_164_n 0.00630228f $X=1.14 $Y=0.825 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_101_n N_B1_c_165_n 9.9843e-19 $X=1.21 $Y=2.13 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_90_n B1 0.00133507f $X=0.587 $Y=1.248 $X2=0 $Y2=0
cc_102 N_A_80_21#_M1010_g B1 5.02998e-19 $X=0.66 $Y=2.735 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_93_n B1 0.044529f $X=0.61 $Y=0.93 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_95_n B1 0.0279053f $X=1.14 $Y=0.825 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_101_n B1 0.0244278f $X=1.21 $Y=2.13 $X2=0 $Y2=0
cc_106 N_A_80_21#_M1010_g N_B1_c_167_n 0.0479714f $X=0.66 $Y=2.735 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_92_n N_B1_c_167_n 0.0094249f $X=0.587 $Y=1.435 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_93_n N_B1_c_167_n 0.00655606f $X=0.61 $Y=0.93 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_101_n N_A4_M1006_g 3.97932e-19 $X=1.21 $Y=2.13 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_103_n N_A4_M1006_g 0.00429293f $X=1.317 $Y=2.395 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_104_n N_A4_M1006_g 0.0134628f $X=1.825 $Y=2.56 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_101_n N_A4_c_216_n 2.97048e-19 $X=1.21 $Y=2.13 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_104_n N_A4_c_216_n 0.00116387f $X=1.825 $Y=2.56 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_101_n A4 0.0153213f $X=1.21 $Y=2.13 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_104_n A4 0.0343856f $X=1.825 $Y=2.56 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_104_n N_A3_M1008_g 0.00236678f $X=1.825 $Y=2.56 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_104_n A3 0.015946f $X=1.825 $Y=2.56 $X2=0 $Y2=0
cc_118 N_A_80_21#_M1010_g N_X_c_408_n 0.011008f $X=0.66 $Y=2.735 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_93_n N_X_c_408_n 0.0889025f $X=0.61 $Y=0.93 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_96_n N_X_c_408_n 0.014009f $X=0.775 $Y=0.825 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_102_n N_X_c_408_n 0.0148239f $X=0.775 $Y=2.13 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_98_n N_X_c_408_n 0.0224918f $X=0.587 $Y=0.765 $X2=0 $Y2=0
cc_123 N_A_80_21#_M1010_g X 6.80668e-19 $X=0.66 $Y=2.735 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_102_n X 0.00121296f $X=0.775 $Y=2.13 $X2=0 $Y2=0
cc_125 N_A_80_21#_M1010_g N_VPWR_c_425_n 0.0126905f $X=0.66 $Y=2.735 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_101_n N_VPWR_c_425_n 0.021102f $X=1.21 $Y=2.13 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_102_n N_VPWR_c_425_n 0.00549266f $X=0.775 $Y=2.13 $X2=0
+ $Y2=0
cc_128 N_A_80_21#_c_104_n N_VPWR_c_425_n 0.0272393f $X=1.825 $Y=2.56 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_104_n N_VPWR_c_428_n 0.0554647f $X=1.825 $Y=2.56 $X2=0 $Y2=0
cc_130 N_A_80_21#_M1010_g N_VPWR_c_429_n 0.00452967f $X=0.66 $Y=2.735 $X2=0
+ $Y2=0
cc_131 N_A_80_21#_M1010_g N_VPWR_c_424_n 0.00897084f $X=0.66 $Y=2.735 $X2=0
+ $Y2=0
cc_132 N_A_80_21#_c_104_n N_VPWR_c_424_n 0.0301936f $X=1.825 $Y=2.56 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_94_n N_VGND_c_463_n 0.0014678f $X=0.61 $Y=0.93 $X2=0 $Y2=0
cc_134 N_A_80_21#_c_95_n N_VGND_c_463_n 0.00633428f $X=1.14 $Y=0.825 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_96_n N_VGND_c_463_n 0.0192456f $X=0.775 $Y=0.825 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_97_n N_VGND_c_463_n 0.0155938f $X=1.305 $Y=0.465 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_98_n N_VGND_c_463_n 0.0108284f $X=0.587 $Y=0.765 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_98_n N_VGND_c_466_n 0.00486043f $X=0.587 $Y=0.765 $X2=0
+ $Y2=0
cc_139 N_A_80_21#_c_95_n N_VGND_c_467_n 0.00419647f $X=1.14 $Y=0.825 $X2=0 $Y2=0
cc_140 N_A_80_21#_c_97_n N_VGND_c_467_n 0.0148312f $X=1.305 $Y=0.465 $X2=0 $Y2=0
cc_141 N_A_80_21#_c_95_n N_VGND_c_470_n 0.00783252f $X=1.14 $Y=0.825 $X2=0 $Y2=0
cc_142 N_A_80_21#_c_96_n N_VGND_c_470_n 0.00104841f $X=0.775 $Y=0.825 $X2=0
+ $Y2=0
cc_143 N_A_80_21#_c_97_n N_VGND_c_470_n 0.0112882f $X=1.305 $Y=0.465 $X2=0 $Y2=0
cc_144 N_A_80_21#_c_98_n N_VGND_c_470_n 0.00931325f $X=0.587 $Y=0.765 $X2=0
+ $Y2=0
cc_145 N_A_80_21#_c_95_n N_A_319_51#_c_519_n 0.00516766f $X=1.14 $Y=0.825 $X2=0
+ $Y2=0
cc_146 N_A_80_21#_c_97_n N_A_319_51#_c_519_n 0.00514425f $X=1.305 $Y=0.465 $X2=0
+ $Y2=0
cc_147 N_A_80_21#_c_95_n N_A_319_51#_c_521_n 0.0102993f $X=1.14 $Y=0.825 $X2=0
+ $Y2=0
cc_148 N_B1_c_164_n N_A4_c_210_n 0.00457862f $X=1.52 $Y=1.155 $X2=-0.19
+ $Y2=-0.245
cc_149 B1 N_A4_c_210_n 5.47243e-19 $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_150 N_B1_c_167_n N_A4_c_210_n 0.00779278f $X=1.18 $Y=1.245 $X2=-0.19
+ $Y2=-0.245
cc_151 N_B1_M1007_g N_A4_M1009_g 0.0277566f $X=1.52 $Y=0.465 $X2=0 $Y2=0
cc_152 B1 N_A4_M1009_g 2.37268e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_153 N_B1_M1005_g N_A4_c_212_n 0.00495217f $X=1.09 $Y=2.735 $X2=0 $Y2=0
cc_154 N_B1_c_165_n N_A4_c_212_n 0.00319495f $X=1.18 $Y=1.75 $X2=0 $Y2=0
cc_155 B1 N_A4_c_212_n 3.01812e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B1_M1005_g A4 0.00520455f $X=1.09 $Y=2.735 $X2=0 $Y2=0
cc_157 N_B1_c_164_n A4 0.0010485f $X=1.52 $Y=1.155 $X2=0 $Y2=0
cc_158 B1 A4 0.0449013f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_159 N_B1_c_167_n A4 0.004639f $X=1.18 $Y=1.245 $X2=0 $Y2=0
cc_160 N_B1_M1005_g N_VPWR_c_425_n 0.0123681f $X=1.09 $Y=2.735 $X2=0 $Y2=0
cc_161 N_B1_M1005_g N_VPWR_c_428_n 0.00452967f $X=1.09 $Y=2.735 $X2=0 $Y2=0
cc_162 N_B1_M1005_g N_VPWR_c_424_n 0.00914997f $X=1.09 $Y=2.735 $X2=0 $Y2=0
cc_163 N_B1_M1007_g N_VGND_c_463_n 0.00313089f $X=1.52 $Y=0.465 $X2=0 $Y2=0
cc_164 N_B1_M1007_g N_VGND_c_467_n 0.00565115f $X=1.52 $Y=0.465 $X2=0 $Y2=0
cc_165 N_B1_M1007_g N_VGND_c_470_n 0.0119838f $X=1.52 $Y=0.465 $X2=0 $Y2=0
cc_166 N_B1_M1007_g N_A_319_51#_c_519_n 0.00104844f $X=1.52 $Y=0.465 $X2=0 $Y2=0
cc_167 N_B1_M1007_g N_A_319_51#_c_521_n 0.00295961f $X=1.52 $Y=0.465 $X2=0 $Y2=0
cc_168 N_A4_c_210_n N_A3_M1000_g 0.0138311f $X=1.95 $Y=1.145 $X2=0 $Y2=0
cc_169 N_A4_M1009_g N_A3_M1000_g 0.0324742f $X=1.95 $Y=0.465 $X2=0 $Y2=0
cc_170 A4 N_A3_M1000_g 0.00751359f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A4_M1006_g N_A3_c_263_n 0.0138311f $X=2.04 $Y=2.735 $X2=0 $Y2=0
cc_172 N_A4_M1006_g N_A3_M1008_g 0.0391864f $X=2.04 $Y=2.735 $X2=0 $Y2=0
cc_173 N_A4_c_216_n N_A3_c_265_n 0.0138311f $X=1.95 $Y=2.14 $X2=0 $Y2=0
cc_174 N_A4_c_210_n A3 3.95908e-19 $X=1.95 $Y=1.145 $X2=0 $Y2=0
cc_175 A4 A3 0.0894897f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_176 N_A4_M1006_g A3 0.002604f $X=2.04 $Y=2.735 $X2=0 $Y2=0
cc_177 A4 A3 3.02879e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A4_c_212_n N_A3_c_262_n 0.0138311f $X=1.95 $Y=1.975 $X2=0 $Y2=0
cc_179 N_A4_c_216_n A3 3.95908e-19 $X=1.95 $Y=2.14 $X2=0 $Y2=0
cc_180 N_A4_M1006_g N_VPWR_c_428_n 0.00509964f $X=2.04 $Y=2.735 $X2=0 $Y2=0
cc_181 N_A4_M1006_g N_VPWR_c_424_n 0.0106686f $X=2.04 $Y=2.735 $X2=0 $Y2=0
cc_182 N_A4_M1009_g N_VGND_c_464_n 0.00316278f $X=1.95 $Y=0.465 $X2=0 $Y2=0
cc_183 N_A4_M1009_g N_VGND_c_467_n 0.00565115f $X=1.95 $Y=0.465 $X2=0 $Y2=0
cc_184 N_A4_M1009_g N_VGND_c_470_n 0.00606107f $X=1.95 $Y=0.465 $X2=0 $Y2=0
cc_185 N_A4_M1009_g N_A_319_51#_c_519_n 0.00187378f $X=1.95 $Y=0.465 $X2=0 $Y2=0
cc_186 N_A4_c_210_n N_A_319_51#_c_520_n 4.95131e-19 $X=1.95 $Y=1.145 $X2=0 $Y2=0
cc_187 N_A4_M1009_g N_A_319_51#_c_520_n 0.0115286f $X=1.95 $Y=0.465 $X2=0 $Y2=0
cc_188 A4 N_A_319_51#_c_520_n 0.0298848f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A4_c_210_n N_A_319_51#_c_521_n 4.23004e-19 $X=1.95 $Y=1.145 $X2=0 $Y2=0
cc_190 A4 N_A_319_51#_c_521_n 0.0238659f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_191 N_A3_M1000_g N_A2_c_314_n 0.0183009f $X=2.4 $Y=0.465 $X2=-0.19 $Y2=-0.245
cc_192 N_A3_c_263_n N_A2_M1011_g 0.0134635f $X=2.49 $Y=2.205 $X2=0 $Y2=0
cc_193 N_A3_M1008_g N_A2_M1011_g 0.0393186f $X=2.49 $Y=2.735 $X2=0 $Y2=0
cc_194 A3 N_A2_c_315_n 5.26526e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_195 N_A3_M1000_g N_A2_c_316_n 0.0175616f $X=2.4 $Y=0.465 $X2=0 $Y2=0
cc_196 A3 N_A2_c_316_n 0.0041812f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A3_c_262_n N_A2_c_317_n 0.0134635f $X=2.49 $Y=1.7 $X2=0 $Y2=0
cc_198 N_A3_c_265_n N_A2_c_322_n 0.0134635f $X=2.49 $Y=2.04 $X2=0 $Y2=0
cc_199 A3 N_A2_c_322_n 0.0041812f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_200 N_A3_M1000_g A2 2.98365e-19 $X=2.4 $Y=0.465 $X2=0 $Y2=0
cc_201 N_A3_M1008_g A2 5.38103e-19 $X=2.49 $Y=2.735 $X2=0 $Y2=0
cc_202 A3 A2 0.133417f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A3_c_262_n A2 5.8708e-19 $X=2.49 $Y=1.7 $X2=0 $Y2=0
cc_204 A3 N_A2_c_319_n 0.0041812f $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_205 N_A3_M1008_g N_VPWR_c_428_n 0.00428854f $X=2.49 $Y=2.735 $X2=0 $Y2=0
cc_206 A3 N_VPWR_c_428_n 0.0079931f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_207 N_A3_M1008_g N_VPWR_c_424_n 0.00713902f $X=2.49 $Y=2.735 $X2=0 $Y2=0
cc_208 A3 N_VPWR_c_424_n 0.0100245f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_209 A3 A_513_483# 0.00644262f $X=2.555 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_210 N_A3_M1000_g N_VGND_c_464_n 0.00170612f $X=2.4 $Y=0.465 $X2=0 $Y2=0
cc_211 N_A3_M1000_g N_VGND_c_465_n 5.47085e-19 $X=2.4 $Y=0.465 $X2=0 $Y2=0
cc_212 N_A3_M1000_g N_VGND_c_468_n 0.00565115f $X=2.4 $Y=0.465 $X2=0 $Y2=0
cc_213 N_A3_M1000_g N_VGND_c_470_n 0.00606107f $X=2.4 $Y=0.465 $X2=0 $Y2=0
cc_214 N_A3_M1000_g N_A_319_51#_c_520_n 0.0141253f $X=2.4 $Y=0.465 $X2=0 $Y2=0
cc_215 A3 N_A_319_51#_c_520_n 0.00606289f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_216 N_A3_M1000_g N_A_319_51#_c_522_n 3.39864e-19 $X=2.4 $Y=0.465 $X2=0 $Y2=0
cc_217 A3 N_A_319_51#_c_523_n 0.00255469f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_218 N_A3_M1000_g N_A_319_51#_c_525_n 0.00181792f $X=2.4 $Y=0.465 $X2=0 $Y2=0
cc_219 A3 N_A_319_51#_c_525_n 0.0221017f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A3_c_262_n N_A_319_51#_c_525_n 5.87827e-19 $X=2.49 $Y=1.7 $X2=0 $Y2=0
cc_221 N_A2_c_314_n N_A1_M1002_g 0.0113297f $X=2.83 $Y=0.785 $X2=0 $Y2=0
cc_222 N_A2_c_315_n N_A1_M1002_g 0.00755947f $X=2.94 $Y=0.86 $X2=0 $Y2=0
cc_223 N_A2_M1011_g N_A1_c_371_n 0.00612947f $X=2.94 $Y=2.735 $X2=0 $Y2=0
cc_224 N_A2_c_322_n N_A1_c_371_n 0.0136568f $X=3.03 $Y=1.915 $X2=0 $Y2=0
cc_225 N_A2_c_316_n N_A1_c_372_n 0.00755947f $X=3.03 $Y=1.245 $X2=0 $Y2=0
cc_226 N_A2_M1011_g N_A1_c_378_n 0.0621967f $X=2.94 $Y=2.735 $X2=0 $Y2=0
cc_227 A2 N_A1_c_378_n 0.00757238f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A2_c_317_n N_A1_c_373_n 0.0136568f $X=3.03 $Y=1.75 $X2=0 $Y2=0
cc_229 N_A2_c_316_n N_A1_c_374_n 0.00756606f $X=3.03 $Y=1.245 $X2=0 $Y2=0
cc_230 A2 N_A1_c_374_n 0.00602621f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_231 N_A2_c_319_n N_A1_c_374_n 0.0136568f $X=3.03 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A2_M1011_g N_A1_c_375_n 2.51687e-19 $X=2.94 $Y=2.735 $X2=0 $Y2=0
cc_233 N_A2_c_316_n N_A1_c_375_n 7.09425e-19 $X=3.03 $Y=1.245 $X2=0 $Y2=0
cc_234 A2 N_A1_c_375_n 0.0714065f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_235 N_A2_c_319_n N_A1_c_375_n 8.27053e-19 $X=3.03 $Y=1.41 $X2=0 $Y2=0
cc_236 A2 N_VPWR_c_427_n 0.0199313f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_237 N_A2_M1011_g N_VPWR_c_428_n 0.00464216f $X=2.94 $Y=2.735 $X2=0 $Y2=0
cc_238 A2 N_VPWR_c_428_n 0.0061079f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_239 N_A2_M1011_g N_VPWR_c_424_n 0.00802727f $X=2.94 $Y=2.735 $X2=0 $Y2=0
cc_240 A2 N_VPWR_c_424_n 0.0084671f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_241 A2 A_603_483# 0.00139886f $X=3.035 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_242 N_A2_c_314_n N_VGND_c_465_n 0.00607213f $X=2.83 $Y=0.785 $X2=0 $Y2=0
cc_243 N_A2_c_315_n N_VGND_c_465_n 5.34923e-19 $X=2.94 $Y=0.86 $X2=0 $Y2=0
cc_244 N_A2_c_314_n N_VGND_c_468_n 0.00402217f $X=2.83 $Y=0.785 $X2=0 $Y2=0
cc_245 N_A2_c_314_n N_VGND_c_470_n 0.0048345f $X=2.83 $Y=0.785 $X2=0 $Y2=0
cc_246 N_A2_c_314_n N_A_319_51#_c_522_n 3.39743e-19 $X=2.83 $Y=0.785 $X2=0 $Y2=0
cc_247 N_A2_c_314_n N_A_319_51#_c_523_n 0.00679759f $X=2.83 $Y=0.785 $X2=0 $Y2=0
cc_248 N_A2_c_315_n N_A_319_51#_c_523_n 0.0136989f $X=2.94 $Y=0.86 $X2=0 $Y2=0
cc_249 A2 N_A_319_51#_c_523_n 0.0149804f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_250 N_A2_c_319_n N_A_319_51#_c_523_n 9.16327e-19 $X=3.03 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A2_c_315_n N_A_319_51#_c_525_n 0.00225451f $X=2.94 $Y=0.86 $X2=0 $Y2=0
cc_252 N_A2_c_316_n N_A_319_51#_c_525_n 0.00100484f $X=3.03 $Y=1.245 $X2=0 $Y2=0
cc_253 N_A1_c_376_n N_VPWR_c_427_n 0.00554652f $X=3.3 $Y=2.305 $X2=0 $Y2=0
cc_254 N_A1_c_378_n N_VPWR_c_427_n 0.00594547f $X=3.48 $Y=2.23 $X2=0 $Y2=0
cc_255 N_A1_c_375_n N_VPWR_c_427_n 0.0217528f $X=3.57 $Y=1.12 $X2=0 $Y2=0
cc_256 N_A1_c_376_n N_VPWR_c_428_n 0.00543892f $X=3.3 $Y=2.305 $X2=0 $Y2=0
cc_257 N_A1_c_376_n N_VPWR_c_424_n 0.010909f $X=3.3 $Y=2.305 $X2=0 $Y2=0
cc_258 N_A1_M1002_g N_VGND_c_465_n 0.00845829f $X=3.3 $Y=0.465 $X2=0 $Y2=0
cc_259 N_A1_M1002_g N_VGND_c_469_n 0.00402217f $X=3.3 $Y=0.465 $X2=0 $Y2=0
cc_260 N_A1_M1002_g N_VGND_c_470_n 0.00572361f $X=3.3 $Y=0.465 $X2=0 $Y2=0
cc_261 N_A1_c_372_n N_VGND_c_470_n 7.93082e-19 $X=3.57 $Y=1.005 $X2=0 $Y2=0
cc_262 N_A1_M1002_g N_A_319_51#_c_523_n 0.0107966f $X=3.3 $Y=0.465 $X2=0 $Y2=0
cc_263 N_A1_c_372_n N_A_319_51#_c_523_n 0.0191729f $X=3.57 $Y=1.005 $X2=0 $Y2=0
cc_264 N_A1_c_375_n N_A_319_51#_c_523_n 0.02496f $X=3.57 $Y=1.12 $X2=0 $Y2=0
cc_265 N_A1_M1002_g N_A_319_51#_c_524_n 8.85348e-19 $X=3.3 $Y=0.465 $X2=0 $Y2=0
cc_266 X N_VPWR_c_425_n 0.0263629f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_267 X N_VPWR_c_429_n 0.0305294f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_268 X N_VPWR_c_424_n 0.0175251f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_269 N_X_c_408_n N_VGND_c_466_n 0.0174138f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_270 N_X_M1003_s N_VGND_c_470_n 0.00371907f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_271 N_X_c_408_n N_VGND_c_470_n 0.0103698f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_272 N_VGND_c_467_n N_A_319_51#_c_519_n 0.0114775f $X=2.035 $Y=0 $X2=0 $Y2=0
cc_273 N_VGND_c_470_n N_A_319_51#_c_519_n 0.00961075f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_274 N_VGND_c_464_n N_A_319_51#_c_520_n 0.0183233f $X=2.18 $Y=0.465 $X2=0
+ $Y2=0
cc_275 N_VGND_c_470_n N_A_319_51#_c_520_n 0.0109853f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_468_n N_A_319_51#_c_522_n 0.0111962f $X=2.9 $Y=0 $X2=0 $Y2=0
cc_277 N_VGND_c_470_n N_A_319_51#_c_522_n 0.00922527f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_465_n N_A_319_51#_c_523_n 0.0206863f $X=3.065 $Y=0.415 $X2=0
+ $Y2=0
cc_279 N_VGND_c_468_n N_A_319_51#_c_523_n 0.00245473f $X=2.9 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_469_n N_A_319_51#_c_523_n 0.00245473f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_470_n N_A_319_51#_c_523_n 0.00919364f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_469_n N_A_319_51#_c_524_n 0.0155705f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_470_n N_A_319_51#_c_524_n 0.0114514f $X=3.6 $Y=0 $X2=0 $Y2=0
