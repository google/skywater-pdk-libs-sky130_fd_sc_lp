* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
X0 VPWR a_27_101# a_196_464# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VGND a_573_535# a_709_411# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 a_709_411# a_196_464# a_1252_451# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_27_101# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VPWR RESET_B a_1399_473# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1252_451# a_27_101# a_1399_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_483_78# D a_318_535# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_318_535# a_196_464# a_573_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_811_119# a_709_411# a_883_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 Q a_1836_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND a_27_101# a_196_464# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1252_451# a_196_464# a_1357_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_27_101# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_573_535# a_196_464# a_811_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1399_473# a_1252_451# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_1399_125# a_1399_473# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_318_535# a_27_101# a_573_535# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_1836_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VGND a_1836_47# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VPWR a_573_535# a_709_411# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 a_1593_125# a_1252_451# a_1399_473# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1836_47# a_1252_451# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VGND RESET_B a_483_78# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR RESET_B a_573_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_1836_47# a_1252_451# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 VGND RESET_B a_1593_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_883_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_709_411# a_27_101# a_1252_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X28 a_573_535# a_27_101# a_667_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_667_535# a_709_411# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 a_1357_535# a_1399_473# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_318_535# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VPWR D a_318_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 Q a_1836_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
