* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND a_33_367# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_223_367# a_33_367# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 Y a_33_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_223_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR A2 a_223_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR A1 a_223_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VGND a_33_367# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 Y a_33_367# a_223_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_223_367# a_33_367# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 Y a_33_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_223_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_33_367# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VPWR A1 a_223_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_223_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_33_367# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 Y a_33_367# a_223_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VPWR A2 a_223_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_223_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
