* NGSPICE file created from sky130_fd_sc_lp__clkbuf_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__clkbuf_2 A VGND VNB VPB VPWR X
M1000 VPWR a_27_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=7.497e+11p pd=6.23e+06u as=3.528e+11p ps=3.08e+06u
M1001 X a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.52e+11p ps=2.88e+06u
M1002 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 X a_27_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_27_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_27_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

