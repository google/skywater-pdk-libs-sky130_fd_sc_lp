* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_49_47# a_462_21# a_218_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND a_218_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_218_367# B2 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_49_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VPWR a_462_21# a_218_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR A1_N a_462_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_218_367# a_462_21# a_49_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_462_21# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR a_218_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_132_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 X a_218_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VPWR B1 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND a_218_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_218_367# a_462_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_462_21# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR a_218_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 X a_218_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_768_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 X a_218_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 X a_218_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VGND B2 a_49_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 VGND A1_N a_768_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_132_367# B2 a_218_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 VPWR A2_N a_462_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_768_47# A2_N a_462_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_49_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_462_21# A2_N a_768_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 VGND B1 a_49_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
