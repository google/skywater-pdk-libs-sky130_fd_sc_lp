* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 X a_110_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND A1 a_1223_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_825_119# S0 a_27_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_80_293# S1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_196_125# a_859_351# a_1381_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_110_125# S1 a_196_125# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VGND S0 a_859_351# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND A3 a_825_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_27_125# a_80_293# a_110_125# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_27_125# a_859_351# a_983_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_80_293# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_196_125# S0 a_1400_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_975_419# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VPWR A3 a_817_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_817_419# a_859_351# a_27_125# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_110_125# a_80_293# a_196_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_983_119# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_125# S1 a_110_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_110_125# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VPWR A1 a_1223_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_1223_419# a_859_351# a_196_125# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 a_27_125# S0 a_975_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 VPWR S0 a_859_351# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 VGND a_110_125# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_1223_119# S0 a_196_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_1400_419# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 X a_110_125# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_1381_119# A0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
