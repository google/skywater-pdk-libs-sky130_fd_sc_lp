* File: sky130_fd_sc_lp__a21oi_lp.spice
* Created: Fri Aug 28 09:51:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21oi_lp.pex.spice"
.subckt sky130_fd_sc_lp__a21oi_lp  VNB VPB A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1002 A_132_47# N_A2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_A1_M1006_g A_132_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 A_324_47# N_B1_M1003_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0882 PD=0.63 PS=0.84 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g A_324_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_31_409#_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_A_31_409#_M1001_d N_A1_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_A_31_409#_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX7_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__a21oi_lp.pxi.spice"
*
.ends
*
*
