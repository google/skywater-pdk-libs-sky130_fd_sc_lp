* File: sky130_fd_sc_lp__and4_1.spice
* Created: Fri Aug 28 10:07:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4_1.pex.spice"
.subckt sky130_fd_sc_lp__and4_1  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1001 A_123_47# N_A_M1001_g N_A_40_47#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.1113 PD=0.75 PS=1.37 NRD=31.428 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1002 A_219_47# N_B_M1002_g A_123_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0693 PD=0.81 PS=0.75 NRD=39.996 NRS=31.428 M=1 R=2.8 SA=75000.7
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 A_327_47# N_C_M1006_g A_219_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=39.996 M=1 R=2.8 SA=75001.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_D_M1000_g A_327_47# VNB NSHORT L=0.15 W=0.42 AD=0.0945
+ AS=0.0819 PD=0.82 PS=0.81 NRD=19.992 NRS=39.996 M=1 R=2.8 SA=75001.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_40_47#_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.189 PD=2.21 PS=1.64 NRD=0 NRS=3.564 M=1 R=5.6 SA=75001.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_A_40_47#_M1008_d N_A_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_A_40_47#_M1008_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0924 AS=0.0819 PD=0.86 PS=0.81 NRD=0 NRS=28.1316 M=1 R=2.8 SA=75000.7
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1009 N_A_40_47#_M1009_d N_C_M1009_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0924 PD=0.7 PS=0.86 NRD=0 NRS=75.0373 M=1 R=2.8 SA=75001.3
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_D_M1004_g N_A_40_47#_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.122325 AS=0.0588 PD=0.9475 PS=0.7 NRD=110.812 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1007 N_X_M1007_d N_A_40_47#_M1007_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.366975 PD=3.05 PS=2.8425 NRD=0 NRS=0 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_60 VPB 0 1.96611e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__and4_1.pxi.spice"
*
.ends
*
*
