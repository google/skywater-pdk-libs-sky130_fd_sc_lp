* File: sky130_fd_sc_lp__sdfsbp_lp.spice
* Created: Wed Sep  2 10:35:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfsbp_lp.pex.spice"
.subckt sky130_fd_sc_lp__sdfsbp_lp  VNB VPB SCE D SCD CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1023 A_138_47# N_SCE_M1023_g N_A_27_409#_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_SCE_M1007_g A_138_47# VNB NSHORT L=0.15 W=0.42 AD=0.1218
+ AS=0.0504 PD=1 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1015 A_362_47# N_A_27_409#_M1015_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1218 PD=0.66 PS=1 NRD=18.564 NRS=85.704 M=1 R=2.8 SA=75001.3
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1016 N_A_352_409#_M1016_d N_D_M1016_g A_362_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1032 A_526_47# N_SCE_M1032_g N_A_352_409#_M1016_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_SCD_M1033_g A_526_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1042 A_848_113# N_CLK_M1042_g N_A_761_113#_M1042_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_CLK_M1006_g A_848_113# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1040 A_1006_113# N_A_761_113#_M1040_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1039 N_A_987_409#_M1039_d N_A_761_113#_M1039_g A_1006_113# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1043 N_A_1201_419#_M1043_d N_A_761_113#_M1043_g N_A_352_409#_M1043_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.093975 AS=0.1197 PD=0.99 PS=1.41 NRD=24.276 NRS=0
+ M=1 R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1018 A_1381_125# N_A_987_409#_M1018_g N_A_1201_419#_M1043_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.093975 PD=0.63 PS=0.99 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_1423_99#_M1011_g A_1381_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.2196 AS=0.0441 PD=2.04 PS=0.63 NRD=133.668 NRS=14.28 M=1 R=2.8 SA=75000.8
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1001 A_1729_125# N_A_1201_419#_M1001_g N_A_1423_99#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_SET_B_M1037_g A_1729_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=11.424 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1002 A_1915_125# N_A_1201_419#_M1002_g N_VGND_M1037_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=19.992 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1022 N_A_2019_419#_M1022_d N_A_987_409#_M1022_g A_1915_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.167725 AS=0.0819 PD=1.31 PS=0.81 NRD=67.14 NRS=39.996 M=1 R=2.8
+ SA=75001.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1028 A_2172_66# N_A_761_113#_M1028_g N_A_2019_419#_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.167725 PD=0.66 PS=1.31 NRD=18.564 NRS=22.848 M=1 R=2.8
+ SA=75000.9 SB=75001 A=0.063 P=1.14 MULT=1
MM1029 A_2250_66# N_A_2220_40#_M1029_g A_2172_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.04515 AS=0.0504 PD=0.635 PS=0.66 NRD=14.988 NRS=18.564 M=1 R=2.8
+ SA=75001.3 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1048 N_VGND_M1048_d N_SET_B_M1048_g A_2250_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.04515 PD=1.41 PS=0.635 NRD=0 NRS=14.988 M=1 R=2.8 SA=75001.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 A_2524_57# N_A_2019_419#_M1013_g N_A_2220_40#_M1013_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_2019_419#_M1014_g A_2524_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1036 A_2682_57# N_A_2019_419#_M1036_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1038 N_Q_N_M1038_d N_A_2019_419#_M1038_g A_2682_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1044 A_2951_74# N_A_2019_419#_M1044_g N_A_2865_74#_M1044_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_A_2019_419#_M1030_g A_2951_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_3109_74# N_A_2865_74#_M1003_g N_VGND_M1030_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1041 N_Q_M1041_d N_A_2865_74#_M1041_g A_3109_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_SCE_M1010_g N_A_27_409#_M1010_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1045 N_A_352_409#_M1045_d N_A_27_409#_M1045_g N_A_245_409#_M1045_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1031 A_458_409# N_D_M1031_g N_A_352_409#_M1045_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.14 PD=1.24 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1046 N_VPWR_M1046_d N_SCE_M1046_g A_458_409# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1024 N_A_245_409#_M1024_d N_SCD_M1024_g N_VPWR_M1046_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1047 N_VPWR_M1047_d N_CLK_M1047_g N_A_761_113#_M1047_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1034 N_A_987_409#_M1034_d N_A_761_113#_M1034_g N_VPWR_M1047_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.275 AS=0.14 PD=2.55 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1008 N_A_1201_419#_M1008_d N_A_987_409#_M1008_g N_A_352_409#_M1008_s VPB
+ PHIGHVT L=0.25 W=1 AD=0.305 AS=0.275 PD=1.61 PS=2.55 NRD=65.01 NRS=0 M=1 R=4
+ SA=125000 SB=125006 A=0.25 P=2.5 MULT=1
MM1020 A_1373_419# N_A_761_113#_M1020_g N_A_1201_419#_M1008_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.305 PD=1.28 PS=1.61 NRD=16.7253 NRS=0 M=1 R=4 SA=125001
+ SB=125006 A=0.25 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_1423_99#_M1004_g A_1373_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.325 AS=0.14 PD=1.65 PS=1.28 NRD=72.8703 NRS=16.7253 M=1 R=4 SA=125002
+ SB=125005 A=0.25 P=2.5 MULT=1
MM1026 N_A_1423_99#_M1026_d N_A_1201_419#_M1026_g N_VPWR_M1004_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.325 PD=1.28 PS=1.65 NRD=0 NRS=0 M=1 R=4 SA=125002
+ SB=125004 A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_SET_B_M1005_g N_A_1423_99#_M1026_d VPB PHIGHVT L=0.25
+ W=1 AD=0.265 AS=0.14 PD=1.53 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125004
+ A=0.25 P=2.5 MULT=1
MM1025 A_1921_419# N_A_1201_419#_M1025_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.265 PD=1.24 PS=1.53 NRD=12.7853 NRS=49.2303 M=1 R=4 SA=125004
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1000 N_A_2019_419#_M1000_d N_A_761_113#_M1000_g A_1921_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.31 AS=0.12 PD=1.62 PS=1.24 NRD=26.5753 NRS=12.7853 M=1 R=4 SA=125004
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1035 A_2193_419# N_A_987_409#_M1035_g N_A_2019_419#_M1000_d VPB PHIGHVT L=0.25
+ W=1 AD=0.16 AS=0.31 PD=1.32 PS=1.62 NRD=20.6653 NRS=40.3653 M=1 R=4 SA=125005
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1021 N_VPWR_M1021_d N_A_2220_40#_M1021_g A_2193_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.225 AS=0.16 PD=1.45 PS=1.32 NRD=0 NRS=20.6653 M=1 R=4 SA=125006 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1027 N_A_2019_419#_M1027_d N_SET_B_M1027_g N_VPWR_M1021_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.225 PD=2.57 PS=1.45 NRD=0 NRS=33.4703 M=1 R=4 SA=125006
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_A_2019_419#_M1012_g N_A_2220_40#_M1012_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.225 AS=0.28 PD=1.45 PS=2.56 NRD=33.4703 NRS=0 M=1 R=4
+ SA=125000 SB=125001 A=0.25 P=2.5 MULT=1
MM1017 N_Q_N_M1017_d N_A_2019_419#_M1017_g N_VPWR_M1012_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.225 PD=2.57 PS=1.45 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A_2019_419#_M1009_g N_A_2865_74#_M1009_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1019 N_Q_M1019_d N_A_2865_74#_M1019_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX49_noxref VNB VPB NWDIODE A=31.1455 P=37.13
c_330 VPB 0 3.86737e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfsbp_lp.pxi.spice"
*
.ends
*
*
