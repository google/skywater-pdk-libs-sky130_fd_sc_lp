* File: sky130_fd_sc_lp__einvp_1.pex.spice
* Created: Fri Aug 28 10:33:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVP_1%A 3 7 9 10 16
c28 3 0 8.15599e-20 $X=0.565 $Y=0.655
r29 14 16 26.6261 $w=3.53e-07 $l=1.95e-07 $layer=POLY_cond $X=0.37 $Y=1.51
+ $X2=0.565 $Y2=1.51
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.46 $X2=0.37 $Y2=1.46
r31 10 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=1.46
r32 9 15 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.46
r33 5 16 22.5297 $w=3.53e-07 $l=2.85832e-07 $layer=POLY_cond $X=0.73 $Y=1.725
+ $X2=0.565 $Y2=1.51
r34 5 7 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=0.73 $Y=1.725
+ $X2=0.73 $Y2=2.5
r35 1 16 22.8335 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.565 $Y=1.295
+ $X2=0.565 $Y2=1.51
r36 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.565 $Y=1.295
+ $X2=0.565 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_1%A_207_302# 1 2 9 11 15 17 19 23 25
c41 23 0 1.07708e-19 $X=1.2 $Y=1.675
c42 11 0 2.64593e-20 $X=1.7 $Y=1.775
r43 23 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.675
+ $X2=1.2 $Y2=1.84
r44 22 25 10.0436 $w=3.03e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=1.712
+ $X2=1.415 $Y2=1.712
r45 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.675 $X2=1.2 $Y2=1.675
r46 17 19 33.7501 $w=2.78e-07 $l=8.2e-07 $layer=LI1_cond $X=2.135 $Y=1.685
+ $X2=2.135 $Y2=0.865
r47 13 17 16.6364 $w=1.78e-07 $l=2.7e-07 $layer=LI1_cond $X=1.865 $Y=1.775
+ $X2=2.135 $Y2=1.775
r48 13 15 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.865 $Y=1.865
+ $X2=1.865 $Y2=2.215
r49 11 13 10.1667 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=1.775
+ $X2=1.865 $Y2=1.775
r50 11 25 17.5606 $w=1.78e-07 $l=2.85e-07 $layer=LI1_cond $X=1.7 $Y=1.775
+ $X2=1.415 $Y2=1.775
r51 9 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.11 $Y=2.5 $X2=1.11
+ $Y2=1.84
r52 2 15 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=1.725 $Y=2
+ $X2=1.865 $Y2=2.215
r53 1 19 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.655 $X2=2.11 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_1%TE 1 3 5 8 10 12 13 14 18 24 28
c42 28 0 3.49599e-20 $X=1.705 $Y=1.285
c43 24 0 8.15599e-20 $X=1.585 $Y=1.285
r44 24 28 1.51847 $w=2.1e-07 $l=1.2e-07 $layer=LI1_cond $X=1.585 $Y=1.285
+ $X2=1.705 $Y2=1.285
r45 17 20 14.2284 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=1.65 $Y=1.332
+ $X2=1.74 $Y2=1.332
r46 17 18 32.4387 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.65 $Y=1.332
+ $X2=1.575 $Y2=1.332
r47 14 28 0.480185 $w=2.38e-07 $l=1e-08 $layer=LI1_cond $X=1.705 $Y=1.295
+ $X2=1.705 $Y2=1.285
r48 14 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.35 $X2=1.74 $Y2=1.35
r49 13 24 20.3333 $w=2.08e-07 $l=3.85e-07 $layer=LI1_cond $X=1.2 $Y=1.285
+ $X2=1.585 $Y2=1.285
r50 10 20 21.3427 $w=3.65e-07 $l=1.35e-07 $layer=POLY_cond $X=1.875 $Y=1.332
+ $X2=1.74 $Y2=1.332
r51 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.875 $Y=1.15
+ $X2=1.875 $Y2=0.865
r52 6 17 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=1.65 $Y=1.515
+ $X2=1.65 $Y2=1.332
r53 6 8 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.65 $Y=1.515
+ $X2=1.65 $Y2=2.21
r54 5 18 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.03 $Y=1.225
+ $X2=1.575 $Y2=1.225
r55 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.955 $Y=1.15
+ $X2=1.03 $Y2=1.225
r56 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.955 $Y=1.15
+ $X2=0.955 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_1%Z 1 2 7 8 9 10 11 12 13 38 46
r30 46 47 5.17831 $w=5.13e-07 $l=7.5e-08 $layer=LI1_cond $X=0.607 $Y=2.035
+ $X2=0.607 $Y2=1.96
r31 29 50 2.13668 $w=5.13e-07 $l=9.2e-08 $layer=LI1_cond $X=0.607 $Y=2.217
+ $X2=0.607 $Y2=2.125
r32 13 35 2.32248 $w=5.13e-07 $l=1e-07 $layer=LI1_cond $X=0.607 $Y=2.775
+ $X2=0.607 $Y2=2.875
r33 12 13 8.59318 $w=5.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.607 $Y=2.405
+ $X2=0.607 $Y2=2.775
r34 12 29 4.36627 $w=5.13e-07 $l=1.88e-07 $layer=LI1_cond $X=0.607 $Y=2.405
+ $X2=0.607 $Y2=2.217
r35 11 50 1.97411 $w=5.13e-07 $l=8.5e-08 $layer=LI1_cond $X=0.607 $Y=2.04
+ $X2=0.607 $Y2=2.125
r36 11 46 0.116124 $w=5.13e-07 $l=5e-09 $layer=LI1_cond $X=0.607 $Y=2.04
+ $X2=0.607 $Y2=2.035
r37 11 47 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=0.745 $Y=1.955
+ $X2=0.745 $Y2=1.96
r38 10 11 13.9254 $w=2.38e-07 $l=2.9e-07 $layer=LI1_cond $X=0.745 $Y=1.665
+ $X2=0.745 $Y2=1.955
r39 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.665
r40 9 44 12.2447 $w=2.38e-07 $l=2.55e-07 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.04
r41 8 44 7.33173 $w=6.78e-07 $l=1.15e-07 $layer=LI1_cond $X=0.525 $Y=0.925
+ $X2=0.525 $Y2=1.04
r42 7 8 6.50807 $w=6.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.525 $Y=0.555
+ $X2=0.525 $Y2=0.925
r43 7 38 3.07814 $w=6.78e-07 $l=1.75e-07 $layer=LI1_cond $X=0.525 $Y=0.555
+ $X2=0.525 $Y2=0.38
r44 2 50 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.37 $Y=2
+ $X2=0.515 $Y2=2.125
r45 2 35 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.37 $Y=2
+ $X2=0.515 $Y2=2.875
r46 1 38 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.225
+ $Y=0.235 $X2=0.35 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_1%VPWR 1 6 10 12 19 20 23
r21 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r22 17 23 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.53 $Y=3.33
+ $X2=1.345 $Y2=3.33
r23 17 19 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.53 $Y=3.33
+ $X2=2.16 $Y2=3.33
r24 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r25 12 23 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=1.345 $Y2=3.33
r26 12 14 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 10 20 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 10 15 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 10 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r30 6 9 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.345 $Y=2.14 $X2=1.345
+ $Y2=2.48
r31 4 23 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.345 $Y=3.245
+ $X2=1.345 $Y2=3.33
r32 4 9 23.8275 $w=3.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.345 $Y=3.245
+ $X2=1.345 $Y2=2.48
r33 1 9 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=1.185 $Y=2
+ $X2=1.325 $Y2=2.48
r34 1 6 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=1.185 $Y=2
+ $X2=1.365 $Y2=2.14
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_1%VGND 1 6 12 14 21 22 25
c22 6 0 9.92069e-20 $X=1.17 $Y=0.38
r23 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r24 22 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r25 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r26 19 25 14.5423 $w=1.7e-07 $l=3.95e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.43
+ $Y2=0
r27 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=2.16
+ $Y2=0
r28 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r29 14 25 14.5423 $w=1.7e-07 $l=3.95e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.43
+ $Y2=0
r30 14 16 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.72
+ $Y2=0
r31 12 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r32 12 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r33 12 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r34 8 10 0.378506 $w=7.88e-07 $l=2.5e-08 $layer=LI1_cond $X=1.43 $Y=0.845
+ $X2=1.43 $Y2=0.87
r35 6 8 7.04021 $w=7.88e-07 $l=4.65e-07 $layer=LI1_cond $X=1.43 $Y=0.38 $X2=1.43
+ $Y2=0.845
r36 4 25 3.10749 $w=7.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.43 $Y=0.085 $X2=1.43
+ $Y2=0
r37 4 6 4.46637 $w=7.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.43 $Y=0.085
+ $X2=1.43 $Y2=0.38
r38 1 10 182 $w=1.7e-07 $l=8.96256e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.66 $Y2=0.87
r39 1 8 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.17 $Y2=0.845
r40 1 6 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.17 $Y2=0.38
.ends

