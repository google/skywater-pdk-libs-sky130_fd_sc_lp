* File: sky130_fd_sc_lp__ha_lp.pxi.spice
* Created: Fri Aug 28 10:36:44 2020
* 
x_PM_SKY130_FD_SC_LP__HA_LP%A_83_153# N_A_83_153#_M1005_s N_A_83_153#_M1013_d
+ N_A_83_153#_M1008_g N_A_83_153#_c_117_n N_A_83_153#_M1006_g
+ N_A_83_153#_M1004_g N_A_83_153#_c_112_n N_A_83_153#_c_113_n
+ N_A_83_153#_c_120_n N_A_83_153#_c_121_n N_A_83_153#_c_114_n
+ N_A_83_153#_c_122_n N_A_83_153#_c_123_n N_A_83_153#_c_115_n
+ PM_SKY130_FD_SC_LP__HA_LP%A_83_153#
x_PM_SKY130_FD_SC_LP__HA_LP%A_296_286# N_A_296_286#_M1003_s N_A_296_286#_M1000_d
+ N_A_296_286#_c_180_n N_A_296_286#_M1013_g N_A_296_286#_M1005_g
+ N_A_296_286#_M1002_g N_A_296_286#_M1012_g N_A_296_286#_M1014_g
+ N_A_296_286#_c_185_n N_A_296_286#_c_186_n N_A_296_286#_c_187_n
+ N_A_296_286#_c_188_n N_A_296_286#_c_189_n N_A_296_286#_c_190_n
+ N_A_296_286#_c_214_p N_A_296_286#_c_191_n N_A_296_286#_c_192_n
+ N_A_296_286#_c_193_n N_A_296_286#_c_194_n PM_SKY130_FD_SC_LP__HA_LP%A_296_286#
x_PM_SKY130_FD_SC_LP__HA_LP%B N_B_M1009_g N_B_M1010_g N_B_M1000_g N_B_M1003_g
+ N_B_c_312_n N_B_c_313_n N_B_c_314_n N_B_c_315_n N_B_c_316_n N_B_c_317_n
+ N_B_c_326_n N_B_c_318_n N_B_c_319_n N_B_c_328_n B B N_B_c_320_n N_B_c_321_n
+ PM_SKY130_FD_SC_LP__HA_LP%B
x_PM_SKY130_FD_SC_LP__HA_LP%A N_A_c_421_n N_A_M1015_g N_A_M1007_g N_A_c_422_n
+ N_A_c_423_n N_A_c_424_n N_A_c_425_n N_A_M1011_g N_A_M1001_g N_A_c_428_n
+ N_A_c_429_n N_A_c_430_n A N_A_c_432_n N_A_c_433_n PM_SKY130_FD_SC_LP__HA_LP%A
x_PM_SKY130_FD_SC_LP__HA_LP%SUM N_SUM_M1008_s N_SUM_M1004_s N_SUM_c_519_n
+ N_SUM_c_520_n N_SUM_c_521_n N_SUM_c_522_n SUM SUM SUM SUM SUM SUM SUM
+ PM_SKY130_FD_SC_LP__HA_LP%SUM
x_PM_SKY130_FD_SC_LP__HA_LP%VPWR N_VPWR_M1004_d N_VPWR_M1007_d N_VPWR_M1011_d
+ N_VPWR_c_546_n N_VPWR_c_547_n N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n
+ VPWR N_VPWR_c_551_n N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_545_n
+ N_VPWR_c_555_n N_VPWR_c_556_n PM_SKY130_FD_SC_LP__HA_LP%VPWR
x_PM_SKY130_FD_SC_LP__HA_LP%COUT N_COUT_M1014_d N_COUT_M1012_d COUT COUT COUT
+ COUT COUT COUT COUT COUT COUT PM_SKY130_FD_SC_LP__HA_LP%COUT
x_PM_SKY130_FD_SC_LP__HA_LP%VGND N_VGND_M1006_d N_VGND_M1009_d N_VGND_M1001_d
+ N_VGND_c_632_n N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n
+ N_VGND_c_637_n N_VGND_c_638_n VGND N_VGND_c_639_n N_VGND_c_640_n
+ N_VGND_c_641_n N_VGND_c_642_n PM_SKY130_FD_SC_LP__HA_LP%VGND
x_PM_SKY130_FD_SC_LP__HA_LP%A_369_47# N_A_369_47#_M1005_d N_A_369_47#_M1015_d
+ N_A_369_47#_c_704_n N_A_369_47#_c_705_n N_A_369_47#_c_706_n
+ N_A_369_47#_c_707_n PM_SKY130_FD_SC_LP__HA_LP%A_369_47#
cc_1 VNB N_A_83_153#_M1008_g 0.033018f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.105
cc_2 VNB N_A_83_153#_M1006_g 0.0274667f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.105
cc_3 VNB N_A_83_153#_c_112_n 0.00480765f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.73
cc_4 VNB N_A_83_153#_c_113_n 0.0174957f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.565
cc_5 VNB N_A_83_153#_c_114_n 0.00562723f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.455
cc_6 VNB N_A_83_153#_c_115_n 0.0153959f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.747
cc_7 VNB N_A_296_286#_c_180_n 0.0584164f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.78
cc_8 VNB N_A_296_286#_M1013_g 0.00654836f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.105
cc_9 VNB N_A_296_286#_M1005_g 0.0379846f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.565
cc_10 VNB N_A_296_286#_M1002_g 0.0187693f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.93
cc_11 VNB N_A_296_286#_M1014_g 0.0214479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_296_286#_c_185_n 0.030609f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.565
cc_13 VNB N_A_296_286#_c_186_n 0.0076012f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.24
cc_14 VNB N_A_296_286#_c_187_n 0.0114917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_296_286#_c_188_n 0.00736018f $X=-0.19 $Y=-0.245 $X2=1.415
+ $Y2=0.455
cc_16 VNB N_A_296_286#_c_189_n 0.00913354f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.73
cc_17 VNB N_A_296_286#_c_190_n 0.00474208f $X=-0.19 $Y=-0.245 $X2=1.075
+ $Y2=1.747
cc_18 VNB N_A_296_286#_c_191_n 0.00239799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_296_286#_c_192_n 0.00244365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_296_286#_c_193_n 0.00121962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_296_286#_c_194_n 0.0406207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_312_n 0.0145113f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=2.595
cc_23 VNB N_B_c_313_n 0.0110673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_314_n 0.0136719f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.73
cc_25 VNB N_B_c_315_n 0.0118105f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.73
cc_26 VNB N_B_c_316_n 0.00244759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_c_317_n 0.00973743f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=0.645
cc_28 VNB N_B_c_318_n 0.00147759f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.24
cc_29 VNB N_B_c_319_n 0.00819918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_c_320_n 0.041387f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.747
cc_31 VNB N_B_c_321_n 0.019019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_c_421_n 0.014915f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=0.235
cc_33 VNB N_A_c_422_n 0.029446f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.855
cc_34 VNB N_A_c_423_n 0.0620698f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.855
cc_35 VNB N_A_c_424_n 0.00997868f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.565
cc_36 VNB N_A_c_425_n 0.00844595f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.105
cc_37 VNB N_A_M1011_g 0.00101055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_M1001_g 0.027788f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.73
cc_39 VNB N_A_c_428_n 0.0339217f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.565
cc_40 VNB N_A_c_429_n 0.0106014f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=1.81
cc_41 VNB N_A_c_430_n 0.0104385f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.24
cc_42 VNB A 0.00510312f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.24
cc_43 VNB N_A_c_432_n 0.0186105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_c_433_n 0.0366535f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.455
cc_45 VNB SUM 0.0582485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VPWR_c_545_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB COUT 0.0214779f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.78
cc_48 VNB COUT 0.0310683f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.105
cc_49 VNB COUT 0.00629578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_632_n 0.0274706f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.855
cc_51 VNB N_VGND_c_633_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_634_n 0.0129285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_635_n 0.0286359f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.73
cc_54 VNB N_VGND_c_636_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.73
cc_55 VNB N_VGND_c_637_n 0.0281028f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=0.645
cc_56 VNB N_VGND_c_638_n 0.00436742f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.565
cc_57 VNB N_VGND_c_639_n 0.0401383f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.747
cc_58 VNB N_VGND_c_640_n 0.0286359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_641_n 0.311743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_642_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_369_47#_c_704_n 8.85615e-19 $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.105
cc_62 VNB N_A_369_47#_c_705_n 0.00849417f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.855
cc_63 VNB N_A_369_47#_c_706_n 0.00167412f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.855
cc_64 VNB N_A_369_47#_c_707_n 0.00519315f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.105
cc_65 VPB N_A_83_153#_M1008_g 0.00730636f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.105
cc_66 VPB N_A_83_153#_c_117_n 0.0143179f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.855
cc_67 VPB N_A_83_153#_M1004_g 0.0302188f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=2.595
cc_68 VPB N_A_83_153#_c_112_n 0.00121982f $X=-0.19 $Y=1.655 $X2=1.33 $Y2=1.73
cc_69 VPB N_A_83_153#_c_120_n 0.00456174f $X=-0.19 $Y=1.655 $X2=1.705 $Y2=1.81
cc_70 VPB N_A_83_153#_c_121_n 0.00214507f $X=-0.19 $Y=1.655 $X2=1.87 $Y2=2.24
cc_71 VPB N_A_83_153#_c_122_n 0.00143357f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.73
cc_72 VPB N_A_83_153#_c_123_n 0.01249f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.747
cc_73 VPB N_A_83_153#_c_115_n 0.0227742f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=1.747
cc_74 VPB N_A_296_286#_M1013_g 0.0438035f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.105
cc_75 VPB N_A_296_286#_M1012_g 0.0327471f $X=-0.19 $Y=1.655 $X2=1.33 $Y2=1.73
cc_76 VPB N_A_296_286#_c_191_n 0.00272934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_296_286#_c_193_n 0.00156697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_296_286#_c_194_n 0.0300099f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_B_M1010_g 0.02643f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.105
cc_80 VPB N_B_M1000_g 0.0246446f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.855
cc_81 VPB N_B_c_316_n 2.63523e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_B_c_317_n 0.0259324f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=0.645
cc_83 VPB N_B_c_326_n 0.00843334f $X=-0.19 $Y=1.655 $X2=1.705 $Y2=1.81
cc_84 VPB N_B_c_319_n 0.022131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_B_c_328_n 0.00954425f $X=-0.19 $Y=1.655 $X2=1.555 $Y2=0.455
cc_86 VPB N_A_M1007_g 0.0350465f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.105
cc_87 VPB N_A_M1011_g 0.0411556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB A 0.0024888f $X=-0.19 $Y=1.655 $X2=1.87 $Y2=2.24
cc_89 VPB N_A_c_432_n 0.00919891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_SUM_c_519_n 0.00978391f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.78
cc_91 VPB N_SUM_c_520_n 0.0115669f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.105
cc_92 VPB N_SUM_c_521_n 2.81881e-19 $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.105
cc_93 VPB N_SUM_c_522_n 0.0058831f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.855
cc_94 VPB SUM 0.0634731f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_546_n 0.00316754f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.855
cc_96 VPB N_VPWR_c_547_n 0.0028319f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=2.595
cc_97 VPB N_VPWR_c_548_n 0.00978644f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=1.73
cc_98 VPB N_VPWR_c_549_n 0.0236936f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.565
cc_99 VPB N_VPWR_c_550_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.705 $Y2=1.81
cc_100 VPB N_VPWR_c_551_n 0.0309611f $X=-0.19 $Y=1.655 $X2=1.87 $Y2=2.24
cc_101 VPB N_VPWR_c_552_n 0.0391741f $X=-0.19 $Y=1.655 $X2=1.555 $Y2=0.455
cc_102 VPB N_VPWR_c_553_n 0.0205832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_545_n 0.0514784f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_555_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_556_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB COUT 0.0220041f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.105
cc_107 VPB COUT 0.0126523f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.855
cc_108 VPB COUT 0.0339892f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.855
cc_109 N_A_83_153#_M1006_g N_A_296_286#_c_180_n 0.00448499f $X=0.85 $Y=1.105
+ $X2=0 $Y2=0
cc_110 N_A_83_153#_c_113_n N_A_296_286#_c_180_n 0.00892652f $X=1.415 $Y=1.565
+ $X2=0 $Y2=0
cc_111 N_A_83_153#_c_120_n N_A_296_286#_c_180_n 0.00187133f $X=1.705 $Y=1.81
+ $X2=0 $Y2=0
cc_112 N_A_83_153#_c_114_n N_A_296_286#_c_180_n 0.00197032f $X=1.555 $Y=0.455
+ $X2=0 $Y2=0
cc_113 N_A_83_153#_c_113_n N_A_296_286#_M1013_g 2.54706e-19 $X=1.415 $Y=1.565
+ $X2=0 $Y2=0
cc_114 N_A_83_153#_c_120_n N_A_296_286#_M1013_g 0.0233598f $X=1.705 $Y=1.81
+ $X2=0 $Y2=0
cc_115 N_A_83_153#_c_121_n N_A_296_286#_M1013_g 0.0271716f $X=1.87 $Y=2.24 $X2=0
+ $Y2=0
cc_116 N_A_83_153#_c_122_n N_A_296_286#_M1013_g 0.00839561f $X=1.415 $Y=1.73
+ $X2=0 $Y2=0
cc_117 N_A_83_153#_c_115_n N_A_296_286#_M1013_g 0.0309586f $X=1.075 $Y=1.747
+ $X2=0 $Y2=0
cc_118 N_A_83_153#_c_113_n N_A_296_286#_M1005_g 0.011438f $X=1.415 $Y=1.565
+ $X2=0 $Y2=0
cc_119 N_A_83_153#_c_120_n N_A_296_286#_c_185_n 0.00213317f $X=1.705 $Y=1.81
+ $X2=0 $Y2=0
cc_120 N_A_83_153#_c_113_n N_A_296_286#_c_190_n 0.023611f $X=1.415 $Y=1.565
+ $X2=0 $Y2=0
cc_121 N_A_83_153#_c_120_n N_A_296_286#_c_190_n 0.0166268f $X=1.705 $Y=1.81
+ $X2=0 $Y2=0
cc_122 N_A_83_153#_c_121_n N_B_M1010_g 0.0119364f $X=1.87 $Y=2.24 $X2=0 $Y2=0
cc_123 N_A_83_153#_c_120_n N_B_c_316_n 0.0137322f $X=1.705 $Y=1.81 $X2=0 $Y2=0
cc_124 N_A_83_153#_c_121_n N_B_c_316_n 0.00481615f $X=1.87 $Y=2.24 $X2=0 $Y2=0
cc_125 N_A_83_153#_c_120_n N_B_c_317_n 0.00164713f $X=1.705 $Y=1.81 $X2=0 $Y2=0
cc_126 N_A_83_153#_c_121_n N_B_c_317_n 3.63142e-19 $X=1.87 $Y=2.24 $X2=0 $Y2=0
cc_127 N_A_83_153#_c_121_n N_B_c_328_n 0.0136067f $X=1.87 $Y=2.24 $X2=0 $Y2=0
cc_128 N_A_83_153#_c_121_n B 0.0585416f $X=1.87 $Y=2.24 $X2=0 $Y2=0
cc_129 N_A_83_153#_c_113_n N_B_c_320_n 5.10568e-19 $X=1.415 $Y=1.565 $X2=0 $Y2=0
cc_130 N_A_83_153#_c_122_n N_B_c_320_n 6.53315e-19 $X=1.415 $Y=1.73 $X2=0 $Y2=0
cc_131 N_A_83_153#_M1004_g N_SUM_c_521_n 0.00318401f $X=1.075 $Y=2.595 $X2=0
+ $Y2=0
cc_132 N_A_83_153#_M1004_g N_SUM_c_522_n 0.0122919f $X=1.075 $Y=2.595 $X2=0
+ $Y2=0
cc_133 N_A_83_153#_c_112_n N_SUM_c_522_n 0.00423013f $X=1.33 $Y=1.73 $X2=0 $Y2=0
cc_134 N_A_83_153#_c_123_n N_SUM_c_522_n 0.0118225f $X=0.775 $Y=1.747 $X2=0
+ $Y2=0
cc_135 N_A_83_153#_M1008_g SUM 0.0294743f $X=0.49 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A_83_153#_c_117_n SUM 0.00836338f $X=0.565 $Y=1.855 $X2=0 $Y2=0
cc_137 N_A_83_153#_M1006_g SUM 0.00338778f $X=0.85 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A_83_153#_M1004_g SUM 0.0053636f $X=1.075 $Y=2.595 $X2=0 $Y2=0
cc_139 N_A_83_153#_c_112_n SUM 0.012276f $X=1.33 $Y=1.73 $X2=0 $Y2=0
cc_140 N_A_83_153#_M1004_g N_VPWR_c_546_n 0.0269479f $X=1.075 $Y=2.595 $X2=0
+ $Y2=0
cc_141 N_A_83_153#_c_112_n N_VPWR_c_546_n 0.0128325f $X=1.33 $Y=1.73 $X2=0 $Y2=0
cc_142 N_A_83_153#_c_121_n N_VPWR_c_546_n 0.0652318f $X=1.87 $Y=2.24 $X2=0 $Y2=0
cc_143 N_A_83_153#_c_122_n N_VPWR_c_546_n 0.0150688f $X=1.415 $Y=1.73 $X2=0
+ $Y2=0
cc_144 N_A_83_153#_M1004_g N_VPWR_c_551_n 0.0083972f $X=1.075 $Y=2.595 $X2=0
+ $Y2=0
cc_145 N_A_83_153#_c_121_n N_VPWR_c_552_n 0.0197322f $X=1.87 $Y=2.24 $X2=0 $Y2=0
cc_146 N_A_83_153#_M1013_d N_VPWR_c_545_n 0.0102336f $X=1.73 $Y=2.095 $X2=0
+ $Y2=0
cc_147 N_A_83_153#_M1004_g N_VPWR_c_545_n 0.0148618f $X=1.075 $Y=2.595 $X2=0
+ $Y2=0
cc_148 N_A_83_153#_c_121_n N_VPWR_c_545_n 0.012508f $X=1.87 $Y=2.24 $X2=0 $Y2=0
cc_149 N_A_83_153#_M1008_g N_VGND_c_632_n 0.00155482f $X=0.49 $Y=1.105 $X2=0
+ $Y2=0
cc_150 N_A_83_153#_M1006_g N_VGND_c_632_n 0.0134046f $X=0.85 $Y=1.105 $X2=0
+ $Y2=0
cc_151 N_A_83_153#_c_112_n N_VGND_c_632_n 0.016573f $X=1.33 $Y=1.73 $X2=0 $Y2=0
cc_152 N_A_83_153#_c_113_n N_VGND_c_632_n 0.0507925f $X=1.415 $Y=1.565 $X2=0
+ $Y2=0
cc_153 N_A_83_153#_c_114_n N_VGND_c_632_n 0.0295988f $X=1.555 $Y=0.455 $X2=0
+ $Y2=0
cc_154 N_A_83_153#_c_115_n N_VGND_c_632_n 0.00580107f $X=1.075 $Y=1.747 $X2=0
+ $Y2=0
cc_155 N_A_83_153#_M1008_g N_VGND_c_635_n 0.00256407f $X=0.49 $Y=1.105 $X2=0
+ $Y2=0
cc_156 N_A_83_153#_M1006_g N_VGND_c_635_n 0.00247589f $X=0.85 $Y=1.105 $X2=0
+ $Y2=0
cc_157 N_A_83_153#_c_114_n N_VGND_c_637_n 0.0195577f $X=1.555 $Y=0.455 $X2=0
+ $Y2=0
cc_158 N_A_83_153#_M1005_s N_VGND_c_641_n 0.00424294f $X=1.41 $Y=0.235 $X2=0
+ $Y2=0
cc_159 N_A_83_153#_M1008_g N_VGND_c_641_n 0.00336713f $X=0.49 $Y=1.105 $X2=0
+ $Y2=0
cc_160 N_A_83_153#_M1006_g N_VGND_c_641_n 0.00336713f $X=0.85 $Y=1.105 $X2=0
+ $Y2=0
cc_161 N_A_83_153#_c_114_n N_VGND_c_641_n 0.0117965f $X=1.555 $Y=0.455 $X2=0
+ $Y2=0
cc_162 N_A_83_153#_c_113_n N_A_369_47#_c_704_n 0.00478581f $X=1.415 $Y=1.565
+ $X2=0 $Y2=0
cc_163 N_A_83_153#_c_113_n N_A_369_47#_c_706_n 0.00843802f $X=1.415 $Y=1.565
+ $X2=0 $Y2=0
cc_164 N_A_296_286#_M1013_g N_B_M1010_g 0.0182575f $X=1.605 $Y=2.595 $X2=0 $Y2=0
cc_165 N_A_296_286#_c_214_p N_B_M1000_g 0.0118256f $X=3.755 $Y=2.475 $X2=0 $Y2=0
cc_166 N_A_296_286#_c_191_n N_B_M1000_g 4.54206e-19 $X=3.812 $Y=2.31 $X2=0 $Y2=0
cc_167 N_A_296_286#_M1005_g N_B_c_312_n 0.0180266f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_296_286#_c_185_n N_B_c_313_n 4.32653e-19 $X=3.26 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A_296_286#_c_186_n N_B_c_314_n 0.00982331f $X=3.425 $Y=0.835 $X2=0
+ $Y2=0
cc_170 N_A_296_286#_c_188_n N_B_c_314_n 7.32582e-19 $X=3.59 $Y=1.31 $X2=0 $Y2=0
cc_171 N_A_296_286#_c_187_n N_B_c_315_n 0.00712941f $X=3.865 $Y=1.31 $X2=0 $Y2=0
cc_172 N_A_296_286#_c_188_n N_B_c_315_n 0.00712797f $X=3.59 $Y=1.31 $X2=0 $Y2=0
cc_173 N_A_296_286#_M1013_g N_B_c_316_n 8.74748e-19 $X=1.605 $Y=2.595 $X2=0
+ $Y2=0
cc_174 N_A_296_286#_c_185_n N_B_c_316_n 0.0152416f $X=3.26 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A_296_286#_M1013_g N_B_c_317_n 0.00615535f $X=1.605 $Y=2.595 $X2=0
+ $Y2=0
cc_176 N_A_296_286#_c_185_n N_B_c_317_n 0.0012059f $X=3.26 $Y=1.185 $X2=0 $Y2=0
cc_177 N_A_296_286#_M1000_d N_B_c_326_n 4.51091e-19 $X=3.615 $Y=2.095 $X2=0
+ $Y2=0
cc_178 N_A_296_286#_c_214_p N_B_c_326_n 0.00296493f $X=3.755 $Y=2.475 $X2=0
+ $Y2=0
cc_179 N_A_296_286#_c_191_n N_B_c_326_n 0.0124144f $X=3.812 $Y=2.31 $X2=0 $Y2=0
cc_180 N_A_296_286#_c_187_n N_B_c_318_n 0.00599467f $X=3.865 $Y=1.31 $X2=0 $Y2=0
cc_181 N_A_296_286#_c_188_n N_B_c_318_n 0.0140773f $X=3.59 $Y=1.31 $X2=0 $Y2=0
cc_182 N_A_296_286#_c_191_n N_B_c_318_n 0.0254343f $X=3.812 $Y=2.31 $X2=0 $Y2=0
cc_183 N_A_296_286#_c_188_n N_B_c_319_n 0.0021044f $X=3.59 $Y=1.31 $X2=0 $Y2=0
cc_184 N_A_296_286#_c_214_p N_B_c_319_n 2.23083e-19 $X=3.755 $Y=2.475 $X2=0
+ $Y2=0
cc_185 N_A_296_286#_c_191_n N_B_c_319_n 0.00174446f $X=3.812 $Y=2.31 $X2=0 $Y2=0
cc_186 N_A_296_286#_M1013_g B 3.42828e-19 $X=1.605 $Y=2.595 $X2=0 $Y2=0
cc_187 N_A_296_286#_c_180_n N_B_c_320_n 0.0276174f $X=1.605 $Y=1.555 $X2=0 $Y2=0
cc_188 N_A_296_286#_M1005_g N_B_c_320_n 0.00813444f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_296_286#_c_185_n N_B_c_320_n 0.0121357f $X=3.26 $Y=1.185 $X2=0 $Y2=0
cc_190 N_A_296_286#_c_190_n N_B_c_320_n 0.00118325f $X=1.832 $Y=1.185 $X2=0
+ $Y2=0
cc_191 N_A_296_286#_c_187_n N_B_c_321_n 0.00339349f $X=3.865 $Y=1.31 $X2=0 $Y2=0
cc_192 N_A_296_286#_c_188_n N_B_c_321_n 0.00370743f $X=3.59 $Y=1.31 $X2=0 $Y2=0
cc_193 N_A_296_286#_c_191_n N_B_c_321_n 0.00259535f $X=3.812 $Y=2.31 $X2=0 $Y2=0
cc_194 N_A_296_286#_c_214_p N_A_M1007_g 2.38814e-19 $X=3.755 $Y=2.475 $X2=0
+ $Y2=0
cc_195 N_A_296_286#_c_186_n N_A_c_422_n 0.00301528f $X=3.425 $Y=0.835 $X2=0
+ $Y2=0
cc_196 N_A_296_286#_c_186_n N_A_c_423_n 0.00531824f $X=3.425 $Y=0.835 $X2=0
+ $Y2=0
cc_197 N_A_296_286#_c_191_n N_A_c_425_n 0.00463515f $X=3.812 $Y=2.31 $X2=0 $Y2=0
cc_198 N_A_296_286#_c_194_n N_A_c_425_n 0.0246634f $X=4.52 $Y=1.39 $X2=0 $Y2=0
cc_199 N_A_296_286#_M1012_g N_A_M1011_g 0.0238034f $X=4.645 $Y=2.595 $X2=0 $Y2=0
cc_200 N_A_296_286#_c_214_p N_A_M1011_g 0.0174387f $X=3.755 $Y=2.475 $X2=0 $Y2=0
cc_201 N_A_296_286#_c_191_n N_A_M1011_g 0.0182604f $X=3.812 $Y=2.31 $X2=0 $Y2=0
cc_202 N_A_296_286#_M1002_g N_A_M1001_g 0.0109876f $X=4.43 $Y=0.835 $X2=0 $Y2=0
cc_203 N_A_296_286#_c_186_n N_A_M1001_g 0.00147033f $X=3.425 $Y=0.835 $X2=0
+ $Y2=0
cc_204 N_A_296_286#_c_188_n N_A_M1001_g 6.33663e-19 $X=3.59 $Y=1.31 $X2=0 $Y2=0
cc_205 N_A_296_286#_c_185_n N_A_c_428_n 0.00800326f $X=3.26 $Y=1.185 $X2=0 $Y2=0
cc_206 N_A_296_286#_c_189_n N_A_c_429_n 0.00718524f $X=4.355 $Y=1.31 $X2=0 $Y2=0
cc_207 N_A_296_286#_c_191_n N_A_c_429_n 0.00255078f $X=3.812 $Y=2.31 $X2=0 $Y2=0
cc_208 N_A_296_286#_c_192_n N_A_c_429_n 0.00215667f $X=3.95 $Y=1.31 $X2=0 $Y2=0
cc_209 N_A_296_286#_c_193_n N_A_c_429_n 0.0017602f $X=4.52 $Y=1.39 $X2=0 $Y2=0
cc_210 N_A_296_286#_M1002_g N_A_c_430_n 0.0246634f $X=4.43 $Y=0.835 $X2=0 $Y2=0
cc_211 N_A_296_286#_c_189_n N_A_c_430_n 0.0024226f $X=4.355 $Y=1.31 $X2=0 $Y2=0
cc_212 N_A_296_286#_c_192_n N_A_c_430_n 0.00730994f $X=3.95 $Y=1.31 $X2=0 $Y2=0
cc_213 N_A_296_286#_c_185_n A 0.0300438f $X=3.26 $Y=1.185 $X2=0 $Y2=0
cc_214 N_A_296_286#_c_191_n A 0.00478201f $X=3.812 $Y=2.31 $X2=0 $Y2=0
cc_215 N_A_296_286#_c_185_n N_A_c_432_n 0.00183904f $X=3.26 $Y=1.185 $X2=0 $Y2=0
cc_216 N_A_296_286#_c_185_n N_A_c_433_n 0.0125134f $X=3.26 $Y=1.185 $X2=0 $Y2=0
cc_217 N_A_296_286#_c_186_n N_A_c_433_n 0.00411897f $X=3.425 $Y=0.835 $X2=0
+ $Y2=0
cc_218 N_A_296_286#_c_188_n N_A_c_433_n 0.00261331f $X=3.59 $Y=1.31 $X2=0 $Y2=0
cc_219 N_A_296_286#_M1013_g N_VPWR_c_546_n 0.0239034f $X=1.605 $Y=2.595 $X2=0
+ $Y2=0
cc_220 N_A_296_286#_M1012_g N_VPWR_c_548_n 0.0240869f $X=4.645 $Y=2.595 $X2=0
+ $Y2=0
cc_221 N_A_296_286#_c_191_n N_VPWR_c_548_n 0.0739434f $X=3.812 $Y=2.31 $X2=0
+ $Y2=0
cc_222 N_A_296_286#_c_193_n N_VPWR_c_548_n 0.0159219f $X=4.52 $Y=1.39 $X2=0
+ $Y2=0
cc_223 N_A_296_286#_c_194_n N_VPWR_c_548_n 0.00127338f $X=4.52 $Y=1.39 $X2=0
+ $Y2=0
cc_224 N_A_296_286#_c_214_p N_VPWR_c_549_n 0.0251507f $X=3.755 $Y=2.475 $X2=0
+ $Y2=0
cc_225 N_A_296_286#_M1013_g N_VPWR_c_552_n 0.00840199f $X=1.605 $Y=2.595 $X2=0
+ $Y2=0
cc_226 N_A_296_286#_M1012_g N_VPWR_c_553_n 0.00840199f $X=4.645 $Y=2.595 $X2=0
+ $Y2=0
cc_227 N_A_296_286#_M1000_d N_VPWR_c_545_n 0.00223819f $X=3.615 $Y=2.095 $X2=0
+ $Y2=0
cc_228 N_A_296_286#_M1013_g N_VPWR_c_545_n 0.0140219f $X=1.605 $Y=2.595 $X2=0
+ $Y2=0
cc_229 N_A_296_286#_M1012_g N_VPWR_c_545_n 0.0145947f $X=4.645 $Y=2.595 $X2=0
+ $Y2=0
cc_230 N_A_296_286#_c_214_p N_VPWR_c_545_n 0.0162338f $X=3.755 $Y=2.475 $X2=0
+ $Y2=0
cc_231 N_A_296_286#_M1002_g COUT 0.00149616f $X=4.43 $Y=0.835 $X2=0 $Y2=0
cc_232 N_A_296_286#_M1014_g COUT 0.00921475f $X=4.79 $Y=0.835 $X2=0 $Y2=0
cc_233 N_A_296_286#_M1012_g COUT 0.00688566f $X=4.645 $Y=2.595 $X2=0 $Y2=0
cc_234 N_A_296_286#_M1014_g COUT 0.026824f $X=4.79 $Y=0.835 $X2=0 $Y2=0
cc_235 N_A_296_286#_c_193_n COUT 0.0405906f $X=4.52 $Y=1.39 $X2=0 $Y2=0
cc_236 N_A_296_286#_M1012_g COUT 0.00528709f $X=4.645 $Y=2.595 $X2=0 $Y2=0
cc_237 N_A_296_286#_c_194_n COUT 0.00454725f $X=4.52 $Y=1.39 $X2=0 $Y2=0
cc_238 N_A_296_286#_M1012_g COUT 0.0193408f $X=4.645 $Y=2.595 $X2=0 $Y2=0
cc_239 N_A_296_286#_M1014_g COUT 0.00436312f $X=4.79 $Y=0.835 $X2=0 $Y2=0
cc_240 N_A_296_286#_M1005_g N_VGND_c_632_n 0.00350261f $X=1.77 $Y=0.445 $X2=0
+ $Y2=0
cc_241 N_A_296_286#_M1005_g N_VGND_c_633_n 0.00127275f $X=1.77 $Y=0.445 $X2=0
+ $Y2=0
cc_242 N_A_296_286#_M1002_g N_VGND_c_634_n 0.01155f $X=4.43 $Y=0.835 $X2=0 $Y2=0
cc_243 N_A_296_286#_M1014_g N_VGND_c_634_n 0.00149701f $X=4.79 $Y=0.835 $X2=0
+ $Y2=0
cc_244 N_A_296_286#_c_186_n N_VGND_c_634_n 0.0147212f $X=3.425 $Y=0.835 $X2=0
+ $Y2=0
cc_245 N_A_296_286#_c_189_n N_VGND_c_634_n 0.0187484f $X=4.355 $Y=1.31 $X2=0
+ $Y2=0
cc_246 N_A_296_286#_c_193_n N_VGND_c_634_n 0.00193744f $X=4.52 $Y=1.39 $X2=0
+ $Y2=0
cc_247 N_A_296_286#_M1005_g N_VGND_c_637_n 0.00549284f $X=1.77 $Y=0.445 $X2=0
+ $Y2=0
cc_248 N_A_296_286#_c_186_n N_VGND_c_639_n 0.00700594f $X=3.425 $Y=0.835 $X2=0
+ $Y2=0
cc_249 N_A_296_286#_M1002_g N_VGND_c_640_n 0.00345209f $X=4.43 $Y=0.835 $X2=0
+ $Y2=0
cc_250 N_A_296_286#_M1014_g N_VGND_c_640_n 0.00359554f $X=4.79 $Y=0.835 $X2=0
+ $Y2=0
cc_251 N_A_296_286#_M1005_g N_VGND_c_641_n 0.0115186f $X=1.77 $Y=0.445 $X2=0
+ $Y2=0
cc_252 N_A_296_286#_M1002_g N_VGND_c_641_n 0.00394323f $X=4.43 $Y=0.835 $X2=0
+ $Y2=0
cc_253 N_A_296_286#_M1014_g N_VGND_c_641_n 0.00394323f $X=4.79 $Y=0.835 $X2=0
+ $Y2=0
cc_254 N_A_296_286#_c_186_n N_VGND_c_641_n 0.00884652f $X=3.425 $Y=0.835 $X2=0
+ $Y2=0
cc_255 N_A_296_286#_M1005_g N_A_369_47#_c_704_n 0.00678968f $X=1.77 $Y=0.445
+ $X2=0 $Y2=0
cc_256 N_A_296_286#_c_185_n N_A_369_47#_c_705_n 0.0676544f $X=3.26 $Y=1.185
+ $X2=0 $Y2=0
cc_257 N_A_296_286#_c_186_n N_A_369_47#_c_705_n 0.0108599f $X=3.425 $Y=0.835
+ $X2=0 $Y2=0
cc_258 N_A_296_286#_c_180_n N_A_369_47#_c_706_n 0.00108267f $X=1.605 $Y=1.555
+ $X2=0 $Y2=0
cc_259 N_A_296_286#_M1005_g N_A_369_47#_c_706_n 0.00492511f $X=1.77 $Y=0.445
+ $X2=0 $Y2=0
cc_260 N_A_296_286#_c_185_n N_A_369_47#_c_706_n 0.00687281f $X=3.26 $Y=1.185
+ $X2=0 $Y2=0
cc_261 N_A_296_286#_c_190_n N_A_369_47#_c_706_n 0.0131548f $X=1.832 $Y=1.185
+ $X2=0 $Y2=0
cc_262 N_A_296_286#_c_186_n N_A_369_47#_c_707_n 0.00891647f $X=3.425 $Y=0.835
+ $X2=0 $Y2=0
cc_263 N_B_c_312_n N_A_c_421_n 0.011888f $X=2.235 $Y=0.73 $X2=-0.19 $Y2=-0.245
cc_264 N_B_M1010_g N_A_M1007_g 0.0483401f $X=2.34 $Y=2.595 $X2=0 $Y2=0
cc_265 N_B_M1000_g N_A_M1007_g 0.0216282f $X=3.49 $Y=2.595 $X2=0 $Y2=0
cc_266 N_B_c_316_n N_A_M1007_g 5.42054e-19 $X=2.38 $Y=1.77 $X2=0 $Y2=0
cc_267 N_B_c_326_n N_A_M1007_g 0.0222712f $X=3.385 $Y=2.045 $X2=0 $Y2=0
cc_268 N_B_c_318_n N_A_M1007_g 0.00108469f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_269 N_B_c_319_n N_A_M1007_g 0.00666118f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_270 N_B_c_314_n N_A_c_422_n 0.00840908f $X=3.61 $Y=1.12 $X2=0 $Y2=0
cc_271 N_B_c_314_n N_A_c_423_n 0.00895007f $X=3.61 $Y=1.12 $X2=0 $Y2=0
cc_272 N_B_c_318_n N_A_c_425_n 3.91303e-19 $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_273 N_B_c_319_n N_A_c_425_n 0.0205981f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_274 N_B_c_321_n N_A_c_425_n 0.00473862f $X=3.52 $Y=1.605 $X2=0 $Y2=0
cc_275 N_B_M1000_g N_A_M1011_g 0.0234586f $X=3.49 $Y=2.595 $X2=0 $Y2=0
cc_276 N_B_c_326_n N_A_M1011_g 6.45496e-19 $X=3.385 $Y=2.045 $X2=0 $Y2=0
cc_277 N_B_c_314_n N_A_M1001_g 0.0229438f $X=3.61 $Y=1.12 $X2=0 $Y2=0
cc_278 N_B_c_313_n N_A_c_428_n 0.00981916f $X=2.235 $Y=0.88 $X2=0 $Y2=0
cc_279 N_B_c_321_n N_A_c_429_n 0.00792682f $X=3.52 $Y=1.605 $X2=0 $Y2=0
cc_280 N_B_c_315_n N_A_c_430_n 0.0229438f $X=3.61 $Y=1.27 $X2=0 $Y2=0
cc_281 N_B_c_316_n A 0.0101366f $X=2.38 $Y=1.77 $X2=0 $Y2=0
cc_282 N_B_c_317_n A 6.48023e-19 $X=2.38 $Y=1.77 $X2=0 $Y2=0
cc_283 N_B_c_326_n A 0.0296663f $X=3.385 $Y=2.045 $X2=0 $Y2=0
cc_284 N_B_c_318_n A 0.0134199f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_285 N_B_c_319_n A 0.00114562f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_286 N_B_c_320_n A 8.5606e-19 $X=2.37 $Y=1.605 $X2=0 $Y2=0
cc_287 N_B_c_321_n A 0.00159729f $X=3.52 $Y=1.605 $X2=0 $Y2=0
cc_288 N_B_c_316_n N_A_c_432_n 0.00127962f $X=2.38 $Y=1.77 $X2=0 $Y2=0
cc_289 N_B_c_317_n N_A_c_432_n 0.0183542f $X=2.38 $Y=1.77 $X2=0 $Y2=0
cc_290 N_B_c_326_n N_A_c_432_n 0.00178213f $X=3.385 $Y=2.045 $X2=0 $Y2=0
cc_291 N_B_c_319_n N_A_c_432_n 0.00920236f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_292 N_B_c_321_n N_A_c_432_n 0.00410157f $X=3.52 $Y=1.605 $X2=0 $Y2=0
cc_293 N_B_c_314_n N_A_c_433_n 0.00194472f $X=3.61 $Y=1.12 $X2=0 $Y2=0
cc_294 N_B_c_315_n N_A_c_433_n 0.00559129f $X=3.61 $Y=1.27 $X2=0 $Y2=0
cc_295 N_B_c_320_n N_A_c_433_n 0.0206924f $X=2.37 $Y=1.605 $X2=0 $Y2=0
cc_296 N_B_c_326_n N_VPWR_M1007_d 0.00235187f $X=3.385 $Y=2.045 $X2=0 $Y2=0
cc_297 N_B_M1010_g N_VPWR_c_547_n 0.00206564f $X=2.34 $Y=2.595 $X2=0 $Y2=0
cc_298 N_B_M1000_g N_VPWR_c_547_n 0.00369345f $X=3.49 $Y=2.595 $X2=0 $Y2=0
cc_299 N_B_c_326_n N_VPWR_c_547_n 0.0185435f $X=3.385 $Y=2.045 $X2=0 $Y2=0
cc_300 N_B_M1000_g N_VPWR_c_549_n 0.00939541f $X=3.49 $Y=2.595 $X2=0 $Y2=0
cc_301 N_B_M1010_g N_VPWR_c_552_n 0.00656883f $X=2.34 $Y=2.595 $X2=0 $Y2=0
cc_302 B N_VPWR_c_552_n 0.0154026f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_303 N_B_M1010_g N_VPWR_c_545_n 0.00880496f $X=2.34 $Y=2.595 $X2=0 $Y2=0
cc_304 N_B_M1000_g N_VPWR_c_545_n 0.0160662f $X=3.49 $Y=2.595 $X2=0 $Y2=0
cc_305 B N_VPWR_c_545_n 0.0175175f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_306 B A_493_419# 0.00553029f $X=2.555 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_307 N_B_c_312_n N_VGND_c_633_n 0.00880914f $X=2.235 $Y=0.73 $X2=0 $Y2=0
cc_308 N_B_c_313_n N_VGND_c_633_n 0.00175361f $X=2.235 $Y=0.88 $X2=0 $Y2=0
cc_309 N_B_c_314_n N_VGND_c_634_n 0.00174932f $X=3.61 $Y=1.12 $X2=0 $Y2=0
cc_310 N_B_c_312_n N_VGND_c_637_n 0.00366861f $X=2.235 $Y=0.73 $X2=0 $Y2=0
cc_311 N_B_c_312_n N_VGND_c_641_n 0.00445761f $X=2.235 $Y=0.73 $X2=0 $Y2=0
cc_312 N_B_c_314_n N_VGND_c_641_n 9.49986e-19 $X=3.61 $Y=1.12 $X2=0 $Y2=0
cc_313 N_B_c_312_n N_A_369_47#_c_704_n 0.0024433f $X=2.235 $Y=0.73 $X2=0 $Y2=0
cc_314 N_B_c_313_n N_A_369_47#_c_705_n 0.0103551f $X=2.235 $Y=0.88 $X2=0 $Y2=0
cc_315 N_B_c_320_n N_A_369_47#_c_705_n 0.00379903f $X=2.37 $Y=1.605 $X2=0 $Y2=0
cc_316 N_A_M1007_g N_VPWR_c_547_n 0.0189735f $X=2.91 $Y=2.595 $X2=0 $Y2=0
cc_317 N_A_M1011_g N_VPWR_c_548_n 0.012824f $X=4.02 $Y=2.595 $X2=0 $Y2=0
cc_318 N_A_M1011_g N_VPWR_c_549_n 0.00766559f $X=4.02 $Y=2.595 $X2=0 $Y2=0
cc_319 N_A_M1007_g N_VPWR_c_552_n 0.008763f $X=2.91 $Y=2.595 $X2=0 $Y2=0
cc_320 N_A_M1007_g N_VPWR_c_545_n 0.0146671f $X=2.91 $Y=2.595 $X2=0 $Y2=0
cc_321 N_A_M1011_g N_VPWR_c_545_n 0.012151f $X=4.02 $Y=2.595 $X2=0 $Y2=0
cc_322 N_A_c_421_n N_VGND_c_633_n 0.00887799f $X=2.63 $Y=0.73 $X2=0 $Y2=0
cc_323 N_A_c_424_n N_VGND_c_633_n 0.00119802f $X=3.21 $Y=0.18 $X2=0 $Y2=0
cc_324 N_A_c_423_n N_VGND_c_634_n 0.00763335f $X=3.925 $Y=0.18 $X2=0 $Y2=0
cc_325 N_A_M1001_g N_VGND_c_634_n 0.0263522f $X=4 $Y=0.835 $X2=0 $Y2=0
cc_326 N_A_c_430_n N_VGND_c_634_n 0.0019288f $X=4.035 $Y=1.27 $X2=0 $Y2=0
cc_327 N_A_c_421_n N_VGND_c_639_n 0.00366861f $X=2.63 $Y=0.73 $X2=0 $Y2=0
cc_328 N_A_c_424_n N_VGND_c_639_n 0.0329746f $X=3.21 $Y=0.18 $X2=0 $Y2=0
cc_329 N_A_c_428_n N_VGND_c_639_n 4.06432e-19 $X=3.135 $Y=0.805 $X2=0 $Y2=0
cc_330 N_A_c_421_n N_VGND_c_641_n 0.00462685f $X=2.63 $Y=0.73 $X2=0 $Y2=0
cc_331 N_A_c_423_n N_VGND_c_641_n 0.0354687f $X=3.925 $Y=0.18 $X2=0 $Y2=0
cc_332 N_A_c_424_n N_VGND_c_641_n 0.0103206f $X=3.21 $Y=0.18 $X2=0 $Y2=0
cc_333 N_A_c_428_n N_A_369_47#_c_705_n 0.0174048f $X=3.135 $Y=0.805 $X2=0 $Y2=0
cc_334 N_A_c_433_n N_A_369_47#_c_705_n 0.00386159f $X=2.95 $Y=1.45 $X2=0 $Y2=0
cc_335 N_A_c_421_n N_A_369_47#_c_707_n 0.00202399f $X=2.63 $Y=0.73 $X2=0 $Y2=0
cc_336 N_A_c_422_n N_A_369_47#_c_707_n 0.0103108f $X=3.135 $Y=0.73 $X2=0 $Y2=0
cc_337 N_A_c_428_n N_A_369_47#_c_707_n 0.00485727f $X=3.135 $Y=0.805 $X2=0 $Y2=0
cc_338 N_SUM_c_521_n N_VPWR_c_546_n 0.0119061f $X=0.81 $Y=2.865 $X2=0 $Y2=0
cc_339 N_SUM_c_522_n N_VPWR_c_546_n 0.0467494f $X=0.81 $Y=2.24 $X2=0 $Y2=0
cc_340 N_SUM_c_519_n N_VPWR_c_551_n 0.0105177f $X=0.645 $Y=2.95 $X2=0 $Y2=0
cc_341 N_SUM_c_520_n N_VPWR_c_551_n 0.0188383f $X=0.44 $Y=2.95 $X2=0 $Y2=0
cc_342 N_SUM_c_521_n N_VPWR_c_551_n 0.0168436f $X=0.81 $Y=2.865 $X2=0 $Y2=0
cc_343 N_SUM_M1004_s N_VPWR_c_545_n 0.00234032f $X=0.665 $Y=2.095 $X2=0 $Y2=0
cc_344 N_SUM_c_519_n N_VPWR_c_545_n 0.00751049f $X=0.645 $Y=2.95 $X2=0 $Y2=0
cc_345 N_SUM_c_520_n N_VPWR_c_545_n 0.0125692f $X=0.44 $Y=2.95 $X2=0 $Y2=0
cc_346 N_SUM_c_521_n N_VPWR_c_545_n 0.0123863f $X=0.81 $Y=2.865 $X2=0 $Y2=0
cc_347 SUM N_VGND_c_632_n 0.0319957f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_348 SUM N_VGND_c_635_n 0.0107254f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_349 SUM N_VGND_c_641_n 0.0114362f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_350 N_VPWR_c_545_n A_493_419# 0.00396518f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_351 N_VPWR_c_545_n N_COUT_M1012_d 0.0023218f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_352 N_VPWR_c_548_n COUT 0.0664847f $X=4.38 $Y=2.24 $X2=0 $Y2=0
cc_353 N_VPWR_c_553_n COUT 0.0261633f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_354 N_VPWR_c_545_n COUT 0.0161839f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_355 COUT N_VGND_c_634_n 0.0206867f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_356 COUT N_VGND_c_640_n 0.0107024f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_357 COUT N_VGND_c_641_n 0.0114229f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_358 N_VGND_c_641_n N_A_369_47#_M1005_d 0.00253635f $X=5.04 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_359 N_VGND_c_641_n N_A_369_47#_M1015_d 0.00253635f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_637_n N_A_369_47#_c_704_n 0.0144108f $X=2.25 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_641_n N_A_369_47#_c_704_n 0.00947015f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_362 N_VGND_c_633_n N_A_369_47#_c_705_n 0.0194905f $X=2.415 $Y=0.39 $X2=0
+ $Y2=0
cc_363 N_VGND_c_637_n N_A_369_47#_c_705_n 0.00236694f $X=2.25 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_639_n N_A_369_47#_c_705_n 0.00226816f $X=4.05 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_641_n N_A_369_47#_c_705_n 0.00934461f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_639_n N_A_369_47#_c_707_n 0.0163393f $X=4.05 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_641_n N_A_369_47#_c_707_n 0.00958069f $X=5.04 $Y=0 $X2=0 $Y2=0
