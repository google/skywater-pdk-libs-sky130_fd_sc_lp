# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfrtp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.455000 2.820000 1.850000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.310000 0.255000 10.535000 1.065000 ;
        RECT 10.310000 1.065000 11.850000 1.235000 ;
        RECT 10.310000 1.755000 11.850000 1.925000 ;
        RECT 10.310000 1.925000 10.535000 3.075000 ;
        RECT 11.150000 0.255000 11.395000 1.065000 ;
        RECT 11.205000 1.925000 11.395000 3.075000 ;
        RECT 11.680000 1.235000 11.850000 1.755000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.735000 2.255000 5.065000 2.520000 ;
        RECT 4.895000 2.520000 5.065000 2.635000 ;
        RECT 4.895000 2.635000 5.955000 2.785000 ;
        RECT 4.895000 2.785000 7.515000 2.805000 ;
        RECT 5.785000 2.805000 7.515000 2.955000 ;
        RECT 7.345000 1.450000 8.565000 1.620000 ;
        RECT 7.345000 1.620000 7.515000 2.785000 ;
        RECT 8.155000 1.620000 8.565000 2.120000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.200000 0.470000 2.130000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.095000  0.495000  0.355000 0.860000 ;
      RECT  0.095000  0.860000  1.205000 1.030000 ;
      RECT  0.195000  2.300000  0.935000 2.470000 ;
      RECT  0.195000  2.470000  0.455000 2.970000 ;
      RECT  0.525000  0.085000  0.865000 0.690000 ;
      RECT  0.625000  2.640000  0.935000 3.245000 ;
      RECT  0.765000  1.030000  1.205000 1.650000 ;
      RECT  0.765000  1.650000  0.935000 2.300000 ;
      RECT  1.035000  0.290000  2.065000 0.460000 ;
      RECT  1.035000  0.460000  1.205000 0.860000 ;
      RECT  1.105000  1.870000  1.715000 2.085000 ;
      RECT  1.105000  2.085000  3.085000 2.285000 ;
      RECT  1.105000  2.285000  1.385000 2.960000 ;
      RECT  1.385000  0.630000  1.715000 1.870000 ;
      RECT  1.660000  2.455000  3.425000 2.625000 ;
      RECT  1.660000  2.625000  1.920000 3.050000 ;
      RECT  1.895000  0.460000  2.065000 1.085000 ;
      RECT  1.895000  1.085000  2.820000 1.255000 ;
      RECT  2.090000  2.795000  2.420000 3.245000 ;
      RECT  2.235000  0.085000  2.480000 0.915000 ;
      RECT  2.590000  2.625000  2.820000 3.050000 ;
      RECT  2.650000  0.365000  4.310000 0.525000 ;
      RECT  2.650000  0.525000  7.425000 0.535000 ;
      RECT  2.650000  0.535000  2.820000 1.085000 ;
      RECT  2.990000  0.725000  3.250000 1.055000 ;
      RECT  2.990000  1.055000  3.195000 1.745000 ;
      RECT  2.990000  1.745000  3.425000 1.915000 ;
      RECT  2.990000  2.795000  3.765000 3.075000 ;
      RECT  3.255000  1.915000  3.425000 2.455000 ;
      RECT  3.365000  1.235000  3.590000 1.565000 ;
      RECT  3.420000  0.535000  3.590000 1.235000 ;
      RECT  3.595000  2.455000  4.545000 2.625000 ;
      RECT  3.595000  2.625000  3.765000 2.795000 ;
      RECT  3.760000  0.715000  3.960000 0.875000 ;
      RECT  3.760000  0.875000  5.605000 1.045000 ;
      RECT  3.835000  1.215000  4.205000 2.180000 ;
      RECT  3.935000  2.795000  4.150000 3.245000 ;
      RECT  4.140000  0.535000  7.425000 0.695000 ;
      RECT  4.320000  2.625000  4.585000 3.050000 ;
      RECT  4.375000  1.215000  4.705000 1.485000 ;
      RECT  4.375000  1.485000  5.955000 1.655000 ;
      RECT  4.375000  1.655000  4.705000 1.745000 ;
      RECT  4.375000  1.915000  5.605000 2.085000 ;
      RECT  4.375000  2.085000  4.545000 2.455000 ;
      RECT  5.155000  0.085000  5.485000 0.355000 ;
      RECT  5.275000  1.045000  5.605000 1.315000 ;
      RECT  5.275000  1.825000  5.605000 1.915000 ;
      RECT  5.275000  2.975000  5.605000 3.245000 ;
      RECT  5.785000  0.865000  6.145000 1.065000 ;
      RECT  5.785000  1.065000  5.955000 1.485000 ;
      RECT  5.785000  1.655000  5.955000 2.205000 ;
      RECT  5.785000  2.205000  6.150000 2.465000 ;
      RECT  6.125000  1.245000  6.485000 1.415000 ;
      RECT  6.125000  1.415000  6.315000 1.955000 ;
      RECT  6.315000  0.695000  6.485000 1.245000 ;
      RECT  6.330000  2.345000  6.660000 2.615000 ;
      RECT  6.485000  1.595000  6.845000 1.765000 ;
      RECT  6.485000  1.765000  6.660000 2.345000 ;
      RECT  6.655000  0.865000  6.985000 1.100000 ;
      RECT  6.655000  1.100000  8.955000 1.270000 ;
      RECT  6.655000  1.270000  6.845000 1.595000 ;
      RECT  6.830000  1.935000  7.165000 2.195000 ;
      RECT  7.095000  0.255000  7.425000 0.525000 ;
      RECT  7.685000  1.950000  7.945000 2.300000 ;
      RECT  7.685000  2.300000  9.295000 2.470000 ;
      RECT  7.715000  2.640000  8.045000 3.245000 ;
      RECT  7.895000  0.085000  8.225000 0.930000 ;
      RECT  8.365000  2.470000  8.695000 2.815000 ;
      RECT  8.735000  1.270000  8.955000 1.865000 ;
      RECT  8.840000  0.650000  9.295000 0.930000 ;
      RECT  8.875000  2.640000  9.205000 3.245000 ;
      RECT  9.125000  0.930000  9.295000 2.300000 ;
      RECT  9.465000  0.255000  9.710000 1.405000 ;
      RECT  9.465000  1.405000 11.500000 1.585000 ;
      RECT  9.465000  1.585000  9.710000 3.075000 ;
      RECT  9.880000  0.085000 10.140000 1.095000 ;
      RECT  9.880000  1.815000 10.140000 3.245000 ;
      RECT 10.705000  0.085000 10.980000 0.895000 ;
      RECT 10.705000  2.095000 11.035000 3.245000 ;
      RECT 11.565000  0.085000 11.895000 0.895000 ;
      RECT 11.565000  2.095000 11.895000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.950000  1.285000 2.120000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.950000  4.165000 2.120000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  1.950000  7.045000 2.120000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
    LAYER met1 ;
      RECT 1.055000 1.920000 1.345000 1.965000 ;
      RECT 1.055000 1.965000 7.105000 2.105000 ;
      RECT 1.055000 2.105000 1.345000 2.150000 ;
      RECT 3.935000 1.920000 4.225000 1.965000 ;
      RECT 3.935000 2.105000 4.225000 2.150000 ;
      RECT 6.815000 1.920000 7.105000 1.965000 ;
      RECT 6.815000 2.105000 7.105000 2.150000 ;
  END
END sky130_fd_sc_lp__dfrtp_4
END LIBRARY
