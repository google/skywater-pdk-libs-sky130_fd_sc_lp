* File: sky130_fd_sc_lp__or2b_m.pex.spice
* Created: Fri Aug 28 11:22:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2B_M%B_N 5 7 8 9 11 13 14 15 16 17 18 23
c38 9 0 9.48564e-20 $X=0.88 $Y=0.86
r39 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r40 17 18 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=2.035
r41 17 24 1.82927 $w=3.13e-07 $l=5e-08 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=1.615
r42 16 24 11.7074 $w=3.13e-07 $l=3.2e-07 $layer=LI1_cond $X=0.312 $Y=1.295
+ $X2=0.312 $Y2=1.615
r43 14 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.955
+ $X2=0.385 $Y2=1.615
r44 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.955
+ $X2=0.385 $Y2=2.12
r45 13 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.45
+ $X2=0.385 $Y2=1.615
r46 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.88 $Y=0.86 $X2=0.88
+ $Y2=0.54
r47 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.805 $Y=0.935
+ $X2=0.88 $Y2=0.86
r48 7 8 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.805 $Y=0.935
+ $X2=0.55 $Y2=0.935
r49 5 15 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.475 $Y=2.69
+ $X2=0.475 $Y2=2.12
r50 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=1.01
+ $X2=0.55 $Y2=0.935
r51 1 13 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.475 $Y=1.01
+ $X2=0.475 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_M%A_27_496# 1 2 9 12 15 17 18 21 23 24 26 28 29
+ 36 38 40 41
c71 40 0 1.503e-19 $X=1.33 $Y=1.025
r72 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.33
+ $Y=1.025 $X2=1.33 $Y2=1.025
r73 34 36 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=0.665 $Y=0.605
+ $X2=0.745 $Y2=0.605
r74 30 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=0.945
+ $X2=0.745 $Y2=0.945
r75 29 40 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.945
+ $X2=1.33 $Y2=0.945
r76 29 30 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.245 $Y=0.945
+ $X2=0.83 $Y2=0.945
r77 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=1.03
+ $X2=0.745 $Y2=0.945
r78 27 28 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=0.745 $Y=1.03
+ $X2=0.745 $Y2=2.3
r79 26 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.86
+ $X2=0.745 $Y2=0.945
r80 25 36 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.745 $Y=0.71
+ $X2=0.745 $Y2=0.605
r81 25 26 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.745 $Y=0.71
+ $X2=0.745 $Y2=0.86
r82 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.66 $Y=2.385
+ $X2=0.745 $Y2=2.3
r83 23 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=2.385
+ $X2=0.345 $Y2=2.385
r84 19 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.25 $Y=2.47
+ $X2=0.345 $Y2=2.385
r85 19 21 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=0.25 $Y=2.47
+ $X2=0.25 $Y2=2.625
r86 17 41 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.33 $Y=1.38
+ $X2=1.33 $Y2=1.025
r87 17 18 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.35 $Y=1.38
+ $X2=1.35 $Y2=1.53
r88 15 41 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.86
+ $X2=1.33 $Y2=1.025
r89 12 18 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.46 $Y=2.1 $X2=1.46
+ $Y2=1.53
r90 9 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.35 $Y=0.54 $X2=1.35
+ $Y2=0.86
r91 2 21 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.48 $X2=0.26 $Y2=2.625
r92 1 34 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.54
+ $Y=0.33 $X2=0.665 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_M%A 3 7 8 9 10 12 22
c41 12 0 8.30343e-20 $X=1.68 $Y=2.775
c42 9 0 1.33837e-19 $X=1.8 $Y=1.01
c43 7 0 1.79498e-19 $X=1.82 $Y=2.1
r44 19 22 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.6 $Y=2.845
+ $X2=1.82 $Y2=2.845
r45 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=2.845 $X2=1.6 $Y2=2.845
r46 12 20 1.56863 $w=6.08e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=2.625 $X2=1.6
+ $Y2=2.625
r47 10 20 7.84314 $w=6.08e-07 $l=4e-07 $layer=LI1_cond $X=1.2 $Y=2.625 $X2=1.6
+ $Y2=2.625
r48 8 9 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.8 $Y=0.86 $X2=1.8
+ $Y2=1.01
r49 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=1.82 $Y=2.1 $X2=1.82
+ $Y2=1.01
r50 5 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=2.68
+ $X2=1.82 $Y2=2.845
r51 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.82 $Y=2.68 $X2=1.82
+ $Y2=2.1
r52 3 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.78 $Y=0.54 $X2=1.78
+ $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_M%A_224_378# 1 2 8 11 15 16 17 22 24 25 32 34
+ 36 37 39
c62 34 0 1.63035e-19 $X=1.68 $Y=0.945
c63 32 0 9.48564e-20 $X=1.68 $Y=0.575
c64 11 0 8.30343e-20 $X=2.325 $Y=2.1
r65 37 39 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.292 $Y=1.025
+ $X2=2.292 $Y2=0.86
r66 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.27
+ $Y=1.025 $X2=2.27 $Y2=1.025
r67 30 32 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=0.575
+ $X2=1.68 $Y2=0.575
r68 26 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0.945
+ $X2=1.68 $Y2=0.945
r69 25 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=0.945
+ $X2=2.27 $Y2=0.945
r70 25 26 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.185 $Y=0.945
+ $X2=1.765 $Y2=0.945
r71 23 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=1.03 $X2=1.68
+ $Y2=0.945
r72 23 24 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=1.68 $Y=1.03 $X2=1.68
+ $Y2=1.93
r73 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=0.86 $X2=1.68
+ $Y2=0.945
r74 21 32 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.68 $Y=0.68 $X2=1.68
+ $Y2=0.575
r75 21 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=0.68
+ $X2=1.68 $Y2=0.86
r76 17 24 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.595 $Y=2.035
+ $X2=1.68 $Y2=1.93
r77 17 19 18.4848 $w=2.08e-07 $l=3.5e-07 $layer=LI1_cond $X=1.595 $Y=2.035
+ $X2=1.245 $Y2=2.035
r78 15 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.405 $Y=0.54
+ $X2=2.405 $Y2=0.86
r79 11 16 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.325 $Y=2.1
+ $X2=2.325 $Y2=1.53
r80 8 16 39.8853 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=2.292 $Y=1.343
+ $X2=2.292 $Y2=1.53
r81 7 37 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=2.292 $Y=1.047
+ $X2=2.292 $Y2=1.025
r82 7 8 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=2.292 $Y=1.047
+ $X2=2.292 $Y2=1.343
r83 2 19 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.89 $X2=1.245 $Y2=2.035
r84 1 30 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.425
+ $Y=0.33 $X2=1.565 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_M%VPWR 1 2 9 13 15 17 22 29 30 33 36
r31 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.11 $Y2=3.33
r36 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r40 23 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=2.11 $Y2=3.33
r42 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r46 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.11 $Y2=3.33
r50 11 13 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.11 $Y2=2.035
r51 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r52 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.755
r53 2 13 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.89 $X2=2.11 $Y2=2.035
r54 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.48 $X2=0.69 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_M%X 1 2 7 8 9 10 11 12 13 36 43
r15 43 44 2.51975 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.59 $Y=2.035
+ $X2=2.59 $Y2=2
r16 34 36 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=2.59 $Y=2.135 $X2=2.59
+ $Y2=2.165
r17 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.59 $Y=2.405
+ $X2=2.59 $Y2=2.775
r18 12 36 10.2439 $w=2.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.59 $Y=2.405
+ $X2=2.59 $Y2=2.165
r19 11 34 3.20123 $w=2.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.59 $Y=2.06
+ $X2=2.59 $Y2=2.135
r20 11 43 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.59 $Y=2.06
+ $X2=2.59 $Y2=2.035
r21 11 44 1.45933 $w=1.88e-07 $l=2.5e-08 $layer=LI1_cond $X=2.63 $Y=1.975
+ $X2=2.63 $Y2=2
r22 10 11 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=2.63 $Y=1.665
+ $X2=2.63 $Y2=1.975
r23 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.63 $Y=1.295
+ $X2=2.63 $Y2=1.665
r24 8 9 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.63 $Y=0.925 $X2=2.63
+ $Y2=1.295
r25 7 8 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.63 $Y=0.555 $X2=2.63
+ $Y2=0.925
r26 2 36 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.89 $X2=2.56 $Y2=2.165
r27 1 7 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.33 $X2=2.62 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_M%VGND 1 2 9 13 16 17 18 24 30 31 34
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r40 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r41 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.11
+ $Y2=0
r43 28 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.64
+ $Y2=0
r44 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r45 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r46 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.11
+ $Y2=0
r47 24 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.68
+ $Y2=0
r48 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r50 18 22 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r51 16 21 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.72
+ $Y2=0
r52 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.115
+ $Y2=0
r53 15 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.68
+ $Y2=0
r54 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.115
+ $Y2=0
r55 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0
r56 11 13 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.475
r57 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0
r58 7 9 20.5974 $w=2.08e-07 $l=3.9e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.475
r59 2 13 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=1.855
+ $Y=0.33 $X2=2.11 $Y2=0.475
r60 1 9 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.955
+ $Y=0.33 $X2=1.115 $Y2=0.475
.ends

