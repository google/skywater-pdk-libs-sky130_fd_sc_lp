* File: sky130_fd_sc_lp__dlxtp_1.pxi.spice
* Created: Fri Aug 28 10:28:56 2020
* 
x_PM_SKY130_FD_SC_LP__DLXTP_1%D N_D_M1007_g N_D_M1008_g N_D_c_120_n N_D_c_121_n
+ N_D_c_122_n D D N_D_c_124_n PM_SKY130_FD_SC_LP__DLXTP_1%D
x_PM_SKY130_FD_SC_LP__DLXTP_1%GATE N_GATE_M1015_g N_GATE_M1009_g N_GATE_c_153_n
+ N_GATE_c_158_n GATE N_GATE_c_154_n N_GATE_c_155_n
+ PM_SKY130_FD_SC_LP__DLXTP_1%GATE
x_PM_SKY130_FD_SC_LP__DLXTP_1%A_27_425# N_A_27_425#_M1008_s N_A_27_425#_M1007_s
+ N_A_27_425#_M1010_g N_A_27_425#_M1003_g N_A_27_425#_c_196_n
+ N_A_27_425#_c_205_n N_A_27_425#_c_197_n N_A_27_425#_c_198_n
+ N_A_27_425#_c_199_n N_A_27_425#_c_200_n N_A_27_425#_c_201_n
+ N_A_27_425#_c_202_n N_A_27_425#_c_203_n PM_SKY130_FD_SC_LP__DLXTP_1%A_27_425#
x_PM_SKY130_FD_SC_LP__DLXTP_1%A_196_425# N_A_196_425#_M1009_d
+ N_A_196_425#_M1015_d N_A_196_425#_c_290_n N_A_196_425#_c_291_n
+ N_A_196_425#_c_292_n N_A_196_425#_c_280_n N_A_196_425#_c_281_n
+ N_A_196_425#_M1000_g N_A_196_425#_c_294_n N_A_196_425#_M1001_g
+ N_A_196_425#_c_282_n N_A_196_425#_M1012_g N_A_196_425#_M1005_g
+ N_A_196_425#_c_296_n N_A_196_425#_c_297_n N_A_196_425#_c_298_n
+ N_A_196_425#_c_284_n N_A_196_425#_c_285_n N_A_196_425#_c_286_n
+ N_A_196_425#_c_287_n N_A_196_425#_c_288_n N_A_196_425#_c_289_n
+ PM_SKY130_FD_SC_LP__DLXTP_1%A_196_425#
x_PM_SKY130_FD_SC_LP__DLXTP_1%A_317_461# N_A_317_461#_M1001_s
+ N_A_317_461#_M1000_s N_A_317_461#_M1017_g N_A_317_461#_M1004_g
+ N_A_317_461#_c_386_n N_A_317_461#_c_400_n N_A_317_461#_c_387_n
+ N_A_317_461#_c_388_n N_A_317_461#_c_389_n N_A_317_461#_c_393_n
+ N_A_317_461#_c_394_n N_A_317_461#_c_390_n N_A_317_461#_c_391_n
+ PM_SKY130_FD_SC_LP__DLXTP_1%A_317_461#
x_PM_SKY130_FD_SC_LP__DLXTP_1%A_733_99# N_A_733_99#_M1016_d N_A_733_99#_M1013_d
+ N_A_733_99#_M1002_g N_A_733_99#_M1006_g N_A_733_99#_M1014_g
+ N_A_733_99#_M1011_g N_A_733_99#_c_475_n N_A_733_99#_c_476_n
+ N_A_733_99#_c_497_p N_A_733_99#_c_486_n N_A_733_99#_c_487_n
+ N_A_733_99#_c_477_n N_A_733_99#_c_478_n N_A_733_99#_c_479_n
+ N_A_733_99#_c_480_n N_A_733_99#_c_481_n PM_SKY130_FD_SC_LP__DLXTP_1%A_733_99#
x_PM_SKY130_FD_SC_LP__DLXTP_1%A_596_419# N_A_596_419#_M1017_d
+ N_A_596_419#_M1012_d N_A_596_419#_M1016_g N_A_596_419#_M1013_g
+ N_A_596_419#_c_571_n N_A_596_419#_c_597_n N_A_596_419#_c_562_n
+ N_A_596_419#_c_563_n N_A_596_419#_c_569_n N_A_596_419#_c_564_n
+ N_A_596_419#_c_576_n N_A_596_419#_c_565_n
+ PM_SKY130_FD_SC_LP__DLXTP_1%A_596_419#
x_PM_SKY130_FD_SC_LP__DLXTP_1%VPWR N_VPWR_M1007_d N_VPWR_M1000_d N_VPWR_M1006_d
+ N_VPWR_M1011_s N_VPWR_c_643_n N_VPWR_c_644_n N_VPWR_c_645_n N_VPWR_c_646_n
+ N_VPWR_c_647_n VPWR N_VPWR_c_648_n N_VPWR_c_649_n N_VPWR_c_650_n
+ N_VPWR_c_651_n N_VPWR_c_652_n N_VPWR_c_642_n N_VPWR_c_654_n N_VPWR_c_655_n
+ N_VPWR_c_656_n N_VPWR_c_657_n PM_SKY130_FD_SC_LP__DLXTP_1%VPWR
x_PM_SKY130_FD_SC_LP__DLXTP_1%Q N_Q_M1014_d N_Q_M1011_d Q Q Q Q Q Q Q
+ N_Q_c_724_n PM_SKY130_FD_SC_LP__DLXTP_1%Q
x_PM_SKY130_FD_SC_LP__DLXTP_1%VGND N_VGND_M1008_d N_VGND_M1001_d N_VGND_M1002_d
+ N_VGND_M1014_s N_VGND_c_736_n N_VGND_c_737_n N_VGND_c_738_n N_VGND_c_739_n
+ N_VGND_c_740_n N_VGND_c_741_n N_VGND_c_742_n N_VGND_c_743_n VGND
+ N_VGND_c_744_n N_VGND_c_745_n N_VGND_c_746_n N_VGND_c_747_n N_VGND_c_748_n
+ N_VGND_c_749_n PM_SKY130_FD_SC_LP__DLXTP_1%VGND
cc_1 VNB N_D_M1007_g 0.012842f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.445
cc_2 VNB N_D_c_120_n 0.0197284f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.775
cc_3 VNB N_D_c_121_n 0.0236573f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.28
cc_4 VNB N_D_c_122_n 0.0166743f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.445
cc_5 VNB D 0.00981975f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_D_c_124_n 0.0164777f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.94
cc_7 VNB N_GATE_c_153_n 0.0308363f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.775
cc_8 VNB N_GATE_c_154_n 0.0322629f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.94
cc_9 VNB N_GATE_c_155_n 0.019804f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=0.925
cc_10 VNB N_A_27_425#_M1003_g 0.0305267f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_A_27_425#_c_196_n 0.0505284f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.94
cc_12 VNB N_A_27_425#_c_197_n 0.00841565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_425#_c_198_n 0.036445f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.295
cc_14 VNB N_A_27_425#_c_199_n 0.0173993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_425#_c_200_n 0.00401891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_425#_c_201_n 0.00197502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_425#_c_202_n 0.00284392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_425#_c_203_n 0.0292893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_196_425#_c_280_n 0.0112291f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_A_196_425#_c_281_n 0.00989737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_196_425#_c_282_n 0.0913545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_196_425#_M1005_g 0.0364676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_196_425#_c_284_n 0.00936603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_196_425#_c_285_n 0.00611018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_196_425#_c_286_n 0.00382931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_196_425#_c_287_n 0.0705168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_196_425#_c_288_n 0.0432967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_196_425#_c_289_n 0.016225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_317_461#_M1017_g 0.0296372f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.775
cc_30 VNB N_A_317_461#_c_386_n 0.00375431f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=0.925
cc_31 VNB N_A_317_461#_c_387_n 0.0048325f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.295
cc_32 VNB N_A_317_461#_c_388_n 0.00478471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_317_461#_c_389_n 0.00401429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_317_461#_c_390_n 0.00273627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_317_461#_c_391_n 0.0290662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_733_99#_M1002_g 0.0195155f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.775
cc_37 VNB N_A_733_99#_M1011_g 0.00374169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_733_99#_c_475_n 0.00171403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_733_99#_c_476_n 0.0299123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_733_99#_c_477_n 0.0139542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_733_99#_c_478_n 0.00713018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_733_99#_c_479_n 0.0163304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_733_99#_c_480_n 0.0418676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_733_99#_c_481_n 0.0227217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_596_419#_c_562_n 0.00101797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_596_419#_c_563_n 0.0293235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_596_419#_c_564_n 0.00784573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_596_419#_c_565_n 0.022397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VPWR_c_642_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_Q_c_724_n 0.0625851f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=0.94
cc_51 VNB N_VGND_c_736_n 0.00548418f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.94
cc_52 VNB N_VGND_c_737_n 0.0117576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_738_n 0.00812603f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.295
cc_54 VNB N_VGND_c_739_n 0.0190069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_740_n 0.00459895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_741_n 0.00182111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_742_n 0.0336866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_743_n 0.00223823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_744_n 0.0412128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_745_n 0.0164605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_746_n 0.310149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_747_n 0.0251177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_748_n 0.00510987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_749_n 0.00406894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VPB N_D_M1007_g 0.0416242f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.445
cc_66 VPB N_GATE_M1015_g 0.0284786f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.445
cc_67 VPB N_GATE_c_153_n 0.00132584f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.775
cc_68 VPB N_GATE_c_158_n 0.0174564f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_69 VPB N_A_27_425#_M1010_g 0.0396978f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.775
cc_70 VPB N_A_27_425#_c_205_n 0.0459465f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=0.925
cc_71 VPB N_A_27_425#_c_197_n 0.00614842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_27_425#_c_200_n 0.00640089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_27_425#_c_201_n 0.00136665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_27_425#_c_202_n 0.00388536f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_27_425#_c_203_n 0.015263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_196_425#_c_290_n 0.0669131f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.94
cc_77 VPB N_A_196_425#_c_291_n 0.0203042f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.775
cc_78 VPB N_A_196_425#_c_292_n 0.0125997f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.28
cc_79 VPB N_A_196_425#_M1000_g 0.0206147f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.94
cc_80 VPB N_A_196_425#_c_294_n 0.0693088f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=0.925
cc_81 VPB N_A_196_425#_M1012_g 0.0389066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_196_425#_c_296_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A_196_425#_c_297_n 0.0280283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_196_425#_c_298_n 0.0100078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A_196_425#_c_285_n 0.029098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_317_461#_M1004_g 0.0207659f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_87 VPB N_A_317_461#_c_393_n 0.00850144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_317_461#_c_394_n 0.0130939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_317_461#_c_390_n 0.00167697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_317_461#_c_391_n 0.0365086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_733_99#_M1006_g 0.0419411f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_92 VPB N_A_733_99#_M1011_g 0.0265209f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_733_99#_c_475_n 0.00275121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_733_99#_c_476_n 0.0066316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_733_99#_c_486_n 0.00701005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_733_99#_c_487_n 0.0123136f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_733_99#_c_479_n 0.0116256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_596_419#_M1013_g 0.0234406f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_99 VPB N_A_596_419#_c_562_n 0.00103501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_596_419#_c_563_n 0.00632576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_596_419#_c_569_n 0.0102863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_596_419#_c_564_n 0.00342176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_643_n 0.0194513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_644_n 0.00595287f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=0.925
cc_105 VPB N_VPWR_c_645_n 0.021421f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.295
cc_106 VPB N_VPWR_c_646_n 0.00373695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_647_n 0.0108191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_648_n 0.0192959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_649_n 0.0353155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_650_n 0.0461121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_651_n 0.0177657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_652_n 0.0157301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_642_n 0.0980914f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_654_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_655_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_656_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_657_n 0.00484208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_Q_c_724_n 0.0581116f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=0.94
cc_119 N_D_M1007_g N_GATE_c_153_n 0.00603422f $X=0.475 $Y=2.445 $X2=0 $Y2=0
cc_120 N_D_c_121_n N_GATE_c_153_n 0.0170898f $X=0.565 $Y=1.28 $X2=0 $Y2=0
cc_121 N_D_M1007_g N_GATE_c_158_n 0.0240727f $X=0.475 $Y=2.445 $X2=0 $Y2=0
cc_122 D GATE 0.0200506f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_123 N_D_c_124_n GATE 3.2213e-19 $X=0.565 $Y=0.94 $X2=0 $Y2=0
cc_124 D N_GATE_c_154_n 0.00901216f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_125 N_D_c_124_n N_GATE_c_154_n 0.0170898f $X=0.565 $Y=0.94 $X2=0 $Y2=0
cc_126 N_D_c_120_n N_GATE_c_155_n 0.0131883f $X=0.565 $Y=0.775 $X2=0 $Y2=0
cc_127 N_D_c_120_n N_A_27_425#_c_196_n 0.00506492f $X=0.565 $Y=0.775 $X2=0 $Y2=0
cc_128 D N_A_27_425#_c_196_n 0.0513623f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_129 N_D_c_124_n N_A_27_425#_c_196_n 0.023167f $X=0.565 $Y=0.94 $X2=0 $Y2=0
cc_130 N_D_M1007_g N_A_27_425#_c_205_n 0.0121013f $X=0.475 $Y=2.445 $X2=0 $Y2=0
cc_131 N_D_M1007_g N_A_27_425#_c_197_n 0.0188817f $X=0.475 $Y=2.445 $X2=0 $Y2=0
cc_132 N_D_c_122_n N_A_27_425#_c_197_n 0.00123716f $X=0.565 $Y=1.445 $X2=0 $Y2=0
cc_133 D N_A_27_425#_c_197_n 0.0263004f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_134 D N_A_27_425#_c_199_n 0.00300687f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_135 N_D_c_124_n N_A_27_425#_c_199_n 0.003496f $X=0.565 $Y=0.94 $X2=0 $Y2=0
cc_136 N_D_M1007_g N_A_27_425#_c_201_n 0.00108423f $X=0.475 $Y=2.445 $X2=0 $Y2=0
cc_137 D N_A_27_425#_c_201_n 0.0060629f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_138 N_D_M1007_g N_VPWR_c_643_n 0.00313675f $X=0.475 $Y=2.445 $X2=0 $Y2=0
cc_139 N_D_M1007_g N_VPWR_c_648_n 0.00448383f $X=0.475 $Y=2.445 $X2=0 $Y2=0
cc_140 N_D_M1007_g N_VPWR_c_642_n 0.00486331f $X=0.475 $Y=2.445 $X2=0 $Y2=0
cc_141 N_D_c_120_n N_VGND_c_736_n 0.00295506f $X=0.565 $Y=0.775 $X2=0 $Y2=0
cc_142 D N_VGND_c_736_n 0.00766253f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_143 N_D_c_120_n N_VGND_c_746_n 0.00706439f $X=0.565 $Y=0.775 $X2=0 $Y2=0
cc_144 D N_VGND_c_746_n 0.00629597f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_145 N_D_c_120_n N_VGND_c_747_n 0.00575161f $X=0.565 $Y=0.775 $X2=0 $Y2=0
cc_146 N_GATE_c_153_n N_A_27_425#_c_197_n 0.00183681f $X=1.045 $Y=1.685 $X2=0
+ $Y2=0
cc_147 N_GATE_c_158_n N_A_27_425#_c_197_n 0.012158f $X=1.045 $Y=1.76 $X2=0 $Y2=0
cc_148 N_GATE_c_153_n N_A_27_425#_c_198_n 5.99064e-19 $X=1.045 $Y=1.685 $X2=0
+ $Y2=0
cc_149 GATE N_A_27_425#_c_198_n 0.00711312f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_150 N_GATE_c_154_n N_A_27_425#_c_198_n 0.00325241f $X=1.135 $Y=0.94 $X2=0
+ $Y2=0
cc_151 N_GATE_c_153_n N_A_27_425#_c_201_n 0.0136528f $X=1.045 $Y=1.685 $X2=0
+ $Y2=0
cc_152 N_GATE_c_158_n N_A_27_425#_c_201_n 0.00388257f $X=1.045 $Y=1.76 $X2=0
+ $Y2=0
cc_153 GATE N_A_27_425#_c_201_n 0.0058421f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_154 N_GATE_c_154_n N_A_27_425#_c_201_n 7.39378e-19 $X=1.135 $Y=0.94 $X2=0
+ $Y2=0
cc_155 N_GATE_c_155_n N_A_196_425#_c_281_n 0.00774496f $X=1.135 $Y=0.775 $X2=0
+ $Y2=0
cc_156 N_GATE_M1015_g N_A_196_425#_c_297_n 0.00547304f $X=0.905 $Y=2.445 $X2=0
+ $Y2=0
cc_157 N_GATE_c_158_n N_A_196_425#_c_297_n 0.00419494f $X=1.045 $Y=1.76 $X2=0
+ $Y2=0
cc_158 N_GATE_M1015_g N_A_196_425#_c_285_n 0.0185864f $X=0.905 $Y=2.445 $X2=0
+ $Y2=0
cc_159 N_GATE_c_153_n N_A_196_425#_c_285_n 0.0107241f $X=1.045 $Y=1.685 $X2=0
+ $Y2=0
cc_160 GATE N_A_196_425#_c_286_n 0.0101893f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_161 N_GATE_c_154_n N_A_196_425#_c_286_n 0.00421148f $X=1.135 $Y=0.94 $X2=0
+ $Y2=0
cc_162 N_GATE_c_153_n N_A_196_425#_c_287_n 0.015555f $X=1.045 $Y=1.685 $X2=0
+ $Y2=0
cc_163 GATE N_A_196_425#_c_287_n 0.00118118f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_164 N_GATE_c_154_n N_A_196_425#_c_287_n 0.0170072f $X=1.135 $Y=0.94 $X2=0
+ $Y2=0
cc_165 GATE N_A_317_461#_c_386_n 0.00829655f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_166 GATE N_A_317_461#_c_388_n 0.00337371f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_167 N_GATE_M1015_g N_VPWR_c_643_n 0.00313675f $X=0.905 $Y=2.445 $X2=0 $Y2=0
cc_168 N_GATE_M1015_g N_VPWR_c_649_n 0.00448383f $X=0.905 $Y=2.445 $X2=0 $Y2=0
cc_169 N_GATE_M1015_g N_VPWR_c_642_n 0.00486331f $X=0.905 $Y=2.445 $X2=0 $Y2=0
cc_170 N_GATE_c_155_n N_VGND_c_736_n 0.00292652f $X=1.135 $Y=0.775 $X2=0 $Y2=0
cc_171 N_GATE_c_155_n N_VGND_c_742_n 0.00575161f $X=1.135 $Y=0.775 $X2=0 $Y2=0
cc_172 GATE N_VGND_c_746_n 0.00242619f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_173 N_GATE_c_155_n N_VGND_c_746_n 0.00976725f $X=1.135 $Y=0.775 $X2=0 $Y2=0
cc_174 N_A_27_425#_M1010_g N_A_196_425#_M1000_g 0.0152546f $X=2.545 $Y=2.415
+ $X2=0 $Y2=0
cc_175 N_A_27_425#_c_198_n N_A_196_425#_M1000_g 0.00383003f $X=2.22 $Y=1.45
+ $X2=0 $Y2=0
cc_176 N_A_27_425#_M1010_g N_A_196_425#_c_294_n 0.0100658f $X=2.545 $Y=2.415
+ $X2=0 $Y2=0
cc_177 N_A_27_425#_M1003_g N_A_196_425#_c_282_n 0.00869842f $X=2.575 $Y=0.835
+ $X2=0 $Y2=0
cc_178 N_A_27_425#_M1010_g N_A_196_425#_M1012_g 0.051303f $X=2.545 $Y=2.415
+ $X2=0 $Y2=0
cc_179 N_A_27_425#_c_205_n N_A_196_425#_c_297_n 0.00532496f $X=0.26 $Y=2.27
+ $X2=0 $Y2=0
cc_180 N_A_27_425#_c_198_n N_A_196_425#_c_297_n 0.0348949f $X=2.22 $Y=1.45 $X2=0
+ $Y2=0
cc_181 N_A_27_425#_c_201_n N_A_196_425#_c_297_n 0.0190625f $X=1.07 $Y=1.45 $X2=0
+ $Y2=0
cc_182 N_A_27_425#_c_202_n N_A_196_425#_c_297_n 0.00117102f $X=2.35 $Y=1.45
+ $X2=0 $Y2=0
cc_183 N_A_27_425#_c_198_n N_A_196_425#_c_285_n 0.005019f $X=2.22 $Y=1.45 $X2=0
+ $Y2=0
cc_184 N_A_27_425#_c_201_n N_A_196_425#_c_285_n 0.00165491f $X=1.07 $Y=1.45
+ $X2=0 $Y2=0
cc_185 N_A_27_425#_c_198_n N_A_196_425#_c_287_n 0.0167598f $X=2.22 $Y=1.45 $X2=0
+ $Y2=0
cc_186 N_A_27_425#_c_201_n N_A_196_425#_c_287_n 0.00183285f $X=1.07 $Y=1.45
+ $X2=0 $Y2=0
cc_187 N_A_27_425#_c_202_n N_A_196_425#_c_287_n 0.00111629f $X=2.35 $Y=1.45
+ $X2=0 $Y2=0
cc_188 N_A_27_425#_c_203_n N_A_196_425#_c_287_n 0.00721797f $X=2.545 $Y=1.58
+ $X2=0 $Y2=0
cc_189 N_A_27_425#_M1003_g N_A_196_425#_c_288_n 0.0159008f $X=2.575 $Y=0.835
+ $X2=0 $Y2=0
cc_190 N_A_27_425#_c_198_n N_A_196_425#_c_289_n 0.00100381f $X=2.22 $Y=1.45
+ $X2=0 $Y2=0
cc_191 N_A_27_425#_M1003_g N_A_317_461#_M1017_g 0.0316493f $X=2.575 $Y=0.835
+ $X2=0 $Y2=0
cc_192 N_A_27_425#_M1010_g N_A_317_461#_c_400_n 0.014394f $X=2.545 $Y=2.415
+ $X2=0 $Y2=0
cc_193 N_A_27_425#_c_202_n N_A_317_461#_c_400_n 0.00670908f $X=2.35 $Y=1.45
+ $X2=0 $Y2=0
cc_194 N_A_27_425#_c_203_n N_A_317_461#_c_400_n 0.0011187f $X=2.545 $Y=1.58
+ $X2=0 $Y2=0
cc_195 N_A_27_425#_M1003_g N_A_317_461#_c_387_n 0.0162053f $X=2.575 $Y=0.835
+ $X2=0 $Y2=0
cc_196 N_A_27_425#_c_198_n N_A_317_461#_c_387_n 0.0140654f $X=2.22 $Y=1.45 $X2=0
+ $Y2=0
cc_197 N_A_27_425#_c_202_n N_A_317_461#_c_387_n 0.0199538f $X=2.35 $Y=1.45 $X2=0
+ $Y2=0
cc_198 N_A_27_425#_c_203_n N_A_317_461#_c_387_n 0.00238904f $X=2.545 $Y=1.58
+ $X2=0 $Y2=0
cc_199 N_A_27_425#_c_198_n N_A_317_461#_c_388_n 0.0205981f $X=2.22 $Y=1.45 $X2=0
+ $Y2=0
cc_200 N_A_27_425#_M1003_g N_A_317_461#_c_389_n 0.00460096f $X=2.575 $Y=0.835
+ $X2=0 $Y2=0
cc_201 N_A_27_425#_c_202_n N_A_317_461#_c_389_n 0.00233256f $X=2.35 $Y=1.45
+ $X2=0 $Y2=0
cc_202 N_A_27_425#_c_202_n N_A_317_461#_c_393_n 0.00147599f $X=2.35 $Y=1.45
+ $X2=0 $Y2=0
cc_203 N_A_27_425#_c_203_n N_A_317_461#_c_393_n 0.0109837f $X=2.545 $Y=1.58
+ $X2=0 $Y2=0
cc_204 N_A_27_425#_M1010_g N_A_317_461#_c_394_n 7.9747e-19 $X=2.545 $Y=2.415
+ $X2=0 $Y2=0
cc_205 N_A_27_425#_M1003_g N_A_317_461#_c_390_n 0.00142751f $X=2.575 $Y=0.835
+ $X2=0 $Y2=0
cc_206 N_A_27_425#_c_202_n N_A_317_461#_c_390_n 0.0256993f $X=2.35 $Y=1.45 $X2=0
+ $Y2=0
cc_207 N_A_27_425#_c_203_n N_A_317_461#_c_390_n 0.00135814f $X=2.545 $Y=1.58
+ $X2=0 $Y2=0
cc_208 N_A_27_425#_c_202_n N_A_317_461#_c_391_n 2.13601e-19 $X=2.35 $Y=1.45
+ $X2=0 $Y2=0
cc_209 N_A_27_425#_c_203_n N_A_317_461#_c_391_n 0.0423403f $X=2.545 $Y=1.58
+ $X2=0 $Y2=0
cc_210 N_A_27_425#_M1003_g N_A_596_419#_c_571_n 8.9428e-19 $X=2.575 $Y=0.835
+ $X2=0 $Y2=0
cc_211 N_A_27_425#_c_205_n N_VPWR_c_643_n 5.96572e-19 $X=0.26 $Y=2.27 $X2=0
+ $Y2=0
cc_212 N_A_27_425#_c_197_n N_VPWR_c_643_n 0.00932471f $X=0.985 $Y=1.71 $X2=0
+ $Y2=0
cc_213 N_A_27_425#_M1010_g N_VPWR_c_644_n 0.00503307f $X=2.545 $Y=2.415 $X2=0
+ $Y2=0
cc_214 N_A_27_425#_c_205_n N_VPWR_c_648_n 0.00671288f $X=0.26 $Y=2.27 $X2=0
+ $Y2=0
cc_215 N_A_27_425#_M1010_g N_VPWR_c_642_n 9.39239e-19 $X=2.545 $Y=2.415 $X2=0
+ $Y2=0
cc_216 N_A_27_425#_c_205_n N_VPWR_c_642_n 0.00894339f $X=0.26 $Y=2.27 $X2=0
+ $Y2=0
cc_217 N_A_27_425#_M1003_g N_VGND_c_737_n 0.00377767f $X=2.575 $Y=0.835 $X2=0
+ $Y2=0
cc_218 N_A_27_425#_M1003_g N_VGND_c_741_n 0.00624294f $X=2.575 $Y=0.835 $X2=0
+ $Y2=0
cc_219 N_A_27_425#_M1008_s N_VGND_c_746_n 0.00209361f $X=0.275 $Y=0.245 $X2=0
+ $Y2=0
cc_220 N_A_27_425#_M1003_g N_VGND_c_746_n 5.12992e-19 $X=2.575 $Y=0.835 $X2=0
+ $Y2=0
cc_221 N_A_27_425#_c_199_n N_VGND_c_746_n 0.0170908f $X=0.4 $Y=0.44 $X2=0 $Y2=0
cc_222 N_A_27_425#_c_199_n N_VGND_c_747_n 0.0268244f $X=0.4 $Y=0.44 $X2=0 $Y2=0
cc_223 N_A_196_425#_c_282_n N_A_317_461#_M1017_g 0.00903991f $X=3.305 $Y=0.18
+ $X2=0 $Y2=0
cc_224 N_A_196_425#_M1005_g N_A_317_461#_M1017_g 0.0152147f $X=3.38 $Y=0.835
+ $X2=0 $Y2=0
cc_225 N_A_196_425#_M1012_g N_A_317_461#_M1004_g 0.010077f $X=2.905 $Y=2.415
+ $X2=0 $Y2=0
cc_226 N_A_196_425#_c_280_n N_A_317_461#_c_386_n 0.00458785f $X=1.89 $Y=0.44
+ $X2=0 $Y2=0
cc_227 N_A_196_425#_c_284_n N_A_317_461#_c_386_n 0.0134879f $X=2.055 $Y=0.35
+ $X2=0 $Y2=0
cc_228 N_A_196_425#_c_287_n N_A_317_461#_c_386_n 0.00565108f $X=1.525 $Y=1.635
+ $X2=0 $Y2=0
cc_229 N_A_196_425#_M1000_g N_A_317_461#_c_400_n 0.0125622f $X=1.925 $Y=2.625
+ $X2=0 $Y2=0
cc_230 N_A_196_425#_c_294_n N_A_317_461#_c_400_n 0.00426216f $X=2.83 $Y=3.15
+ $X2=0 $Y2=0
cc_231 N_A_196_425#_c_284_n N_A_317_461#_c_387_n 0.00364031f $X=2.055 $Y=0.35
+ $X2=0 $Y2=0
cc_232 N_A_196_425#_c_289_n N_A_317_461#_c_387_n 0.0116257f $X=2.055 $Y=0.515
+ $X2=0 $Y2=0
cc_233 N_A_196_425#_c_287_n N_A_317_461#_c_388_n 0.0040176f $X=1.525 $Y=1.635
+ $X2=0 $Y2=0
cc_234 N_A_196_425#_M1012_g N_A_317_461#_c_393_n 0.00209172f $X=2.905 $Y=2.415
+ $X2=0 $Y2=0
cc_235 N_A_196_425#_c_290_n N_A_317_461#_c_394_n 0.00992908f $X=1.435 $Y=3.075
+ $X2=0 $Y2=0
cc_236 N_A_196_425#_c_291_n N_A_317_461#_c_394_n 0.00373696f $X=1.85 $Y=3.15
+ $X2=0 $Y2=0
cc_237 N_A_196_425#_M1000_g N_A_317_461#_c_394_n 0.00907231f $X=1.925 $Y=2.625
+ $X2=0 $Y2=0
cc_238 N_A_196_425#_c_297_n N_A_317_461#_c_394_n 0.0129189f $X=1.175 $Y=2.135
+ $X2=0 $Y2=0
cc_239 N_A_196_425#_c_298_n N_A_317_461#_c_394_n 0.034346f $X=1.12 $Y=2.27 $X2=0
+ $Y2=0
cc_240 N_A_196_425#_c_285_n N_A_317_461#_c_394_n 7.53215e-19 $X=1.525 $Y=1.8
+ $X2=0 $Y2=0
cc_241 N_A_196_425#_M1012_g N_A_317_461#_c_390_n 0.00214315f $X=2.905 $Y=2.415
+ $X2=0 $Y2=0
cc_242 N_A_196_425#_M1012_g N_A_317_461#_c_391_n 0.00793765f $X=2.905 $Y=2.415
+ $X2=0 $Y2=0
cc_243 N_A_196_425#_M1005_g N_A_317_461#_c_391_n 0.00307587f $X=3.38 $Y=0.835
+ $X2=0 $Y2=0
cc_244 N_A_196_425#_M1005_g N_A_733_99#_M1002_g 0.0428995f $X=3.38 $Y=0.835
+ $X2=0 $Y2=0
cc_245 N_A_196_425#_c_282_n N_A_596_419#_c_571_n 0.00421869f $X=3.305 $Y=0.18
+ $X2=0 $Y2=0
cc_246 N_A_196_425#_M1012_g N_A_596_419#_c_569_n 0.0021189f $X=2.905 $Y=2.415
+ $X2=0 $Y2=0
cc_247 N_A_196_425#_M1012_g N_A_596_419#_c_564_n 8.19215e-19 $X=2.905 $Y=2.415
+ $X2=0 $Y2=0
cc_248 N_A_196_425#_M1005_g N_A_596_419#_c_564_n 0.00573801f $X=3.38 $Y=0.835
+ $X2=0 $Y2=0
cc_249 N_A_196_425#_M1005_g N_A_596_419#_c_576_n 0.00887196f $X=3.38 $Y=0.835
+ $X2=0 $Y2=0
cc_250 N_A_196_425#_c_290_n N_VPWR_c_643_n 0.00683391f $X=1.435 $Y=3.075 $X2=0
+ $Y2=0
cc_251 N_A_196_425#_c_298_n N_VPWR_c_643_n 6.02795e-19 $X=1.12 $Y=2.27 $X2=0
+ $Y2=0
cc_252 N_A_196_425#_M1000_g N_VPWR_c_644_n 0.00894606f $X=1.925 $Y=2.625 $X2=0
+ $Y2=0
cc_253 N_A_196_425#_c_294_n N_VPWR_c_644_n 0.0248871f $X=2.83 $Y=3.15 $X2=0
+ $Y2=0
cc_254 N_A_196_425#_M1012_g N_VPWR_c_644_n 0.006256f $X=2.905 $Y=2.415 $X2=0
+ $Y2=0
cc_255 N_A_196_425#_c_292_n N_VPWR_c_649_n 0.022531f $X=1.51 $Y=3.15 $X2=0 $Y2=0
cc_256 N_A_196_425#_c_298_n N_VPWR_c_649_n 0.00767876f $X=1.12 $Y=2.27 $X2=0
+ $Y2=0
cc_257 N_A_196_425#_c_294_n N_VPWR_c_650_n 0.0213287f $X=2.83 $Y=3.15 $X2=0
+ $Y2=0
cc_258 N_A_196_425#_c_291_n N_VPWR_c_642_n 0.00956062f $X=1.85 $Y=3.15 $X2=0
+ $Y2=0
cc_259 N_A_196_425#_c_292_n N_VPWR_c_642_n 0.0116041f $X=1.51 $Y=3.15 $X2=0
+ $Y2=0
cc_260 N_A_196_425#_c_294_n N_VPWR_c_642_n 0.0266741f $X=2.83 $Y=3.15 $X2=0
+ $Y2=0
cc_261 N_A_196_425#_c_296_n N_VPWR_c_642_n 0.00458911f $X=1.925 $Y=3.15 $X2=0
+ $Y2=0
cc_262 N_A_196_425#_c_298_n N_VPWR_c_642_n 0.0102302f $X=1.12 $Y=2.27 $X2=0
+ $Y2=0
cc_263 N_A_196_425#_c_282_n N_VGND_c_737_n 0.0156385f $X=3.305 $Y=0.18 $X2=0
+ $Y2=0
cc_264 N_A_196_425#_c_284_n N_VGND_c_737_n 0.0136197f $X=2.055 $Y=0.35 $X2=0
+ $Y2=0
cc_265 N_A_196_425#_c_288_n N_VGND_c_737_n 0.00599011f $X=2.055 $Y=0.18 $X2=0
+ $Y2=0
cc_266 N_A_196_425#_c_282_n N_VGND_c_738_n 0.00986715f $X=3.305 $Y=0.18 $X2=0
+ $Y2=0
cc_267 N_A_196_425#_c_282_n N_VGND_c_741_n 0.00203586f $X=3.305 $Y=0.18 $X2=0
+ $Y2=0
cc_268 N_A_196_425#_c_284_n N_VGND_c_741_n 0.001646f $X=2.055 $Y=0.35 $X2=0
+ $Y2=0
cc_269 N_A_196_425#_c_287_n N_VGND_c_741_n 3.58144e-19 $X=1.525 $Y=1.635 $X2=0
+ $Y2=0
cc_270 N_A_196_425#_c_289_n N_VGND_c_741_n 0.00401642f $X=2.055 $Y=0.515 $X2=0
+ $Y2=0
cc_271 N_A_196_425#_c_281_n N_VGND_c_742_n 0.0016819f $X=1.69 $Y=0.44 $X2=0
+ $Y2=0
cc_272 N_A_196_425#_c_284_n N_VGND_c_742_n 0.0504468f $X=2.055 $Y=0.35 $X2=0
+ $Y2=0
cc_273 N_A_196_425#_c_286_n N_VGND_c_742_n 0.0185939f $X=1.272 $Y=0.345 $X2=0
+ $Y2=0
cc_274 N_A_196_425#_c_288_n N_VGND_c_742_n 0.0124291f $X=2.055 $Y=0.18 $X2=0
+ $Y2=0
cc_275 N_A_196_425#_c_282_n N_VGND_c_744_n 0.0320948f $X=3.305 $Y=0.18 $X2=0
+ $Y2=0
cc_276 N_A_196_425#_M1009_d N_VGND_c_746_n 0.00212301f $X=1.12 $Y=0.245 $X2=0
+ $Y2=0
cc_277 N_A_196_425#_c_282_n N_VGND_c_746_n 0.0391074f $X=3.305 $Y=0.18 $X2=0
+ $Y2=0
cc_278 N_A_196_425#_c_284_n N_VGND_c_746_n 0.0284243f $X=2.055 $Y=0.35 $X2=0
+ $Y2=0
cc_279 N_A_196_425#_c_286_n N_VGND_c_746_n 0.011586f $X=1.272 $Y=0.345 $X2=0
+ $Y2=0
cc_280 N_A_196_425#_c_288_n N_VGND_c_746_n 0.0103902f $X=2.055 $Y=0.18 $X2=0
+ $Y2=0
cc_281 N_A_317_461#_M1017_g N_A_733_99#_M1002_g 0.00232903f $X=2.935 $Y=0.835
+ $X2=0 $Y2=0
cc_282 N_A_317_461#_c_391_n N_A_733_99#_M1006_g 0.0590274f $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_283 N_A_317_461#_c_391_n N_A_733_99#_c_475_n 3.71524e-19 $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_284 N_A_317_461#_c_391_n N_A_733_99#_c_476_n 0.00219367f $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_285 N_A_317_461#_c_391_n N_A_733_99#_c_486_n 9.56664e-19 $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_286 N_A_317_461#_M1017_g N_A_596_419#_c_571_n 0.00378663f $X=2.935 $Y=0.835
+ $X2=0 $Y2=0
cc_287 N_A_317_461#_c_390_n N_A_596_419#_c_571_n 0.00354763f $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_288 N_A_317_461#_c_391_n N_A_596_419#_c_571_n 0.00602837f $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_289 N_A_317_461#_M1004_g N_A_596_419#_c_569_n 0.0170529f $X=3.43 $Y=2.305
+ $X2=0 $Y2=0
cc_290 N_A_317_461#_c_393_n N_A_596_419#_c_569_n 0.00139979f $X=2.735 $Y=2.305
+ $X2=0 $Y2=0
cc_291 N_A_317_461#_c_390_n N_A_596_419#_c_569_n 0.00512088f $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_292 N_A_317_461#_c_391_n N_A_596_419#_c_569_n 0.0088047f $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_293 N_A_317_461#_M1017_g N_A_596_419#_c_564_n 0.00312352f $X=2.935 $Y=0.835
+ $X2=0 $Y2=0
cc_294 N_A_317_461#_M1004_g N_A_596_419#_c_564_n 0.00543222f $X=3.43 $Y=2.305
+ $X2=0 $Y2=0
cc_295 N_A_317_461#_c_387_n N_A_596_419#_c_564_n 0.0057591f $X=2.65 $Y=1.1 $X2=0
+ $Y2=0
cc_296 N_A_317_461#_c_389_n N_A_596_419#_c_564_n 0.00776148f $X=2.735 $Y=1.395
+ $X2=0 $Y2=0
cc_297 N_A_317_461#_c_393_n N_A_596_419#_c_564_n 0.0123145f $X=2.735 $Y=2.305
+ $X2=0 $Y2=0
cc_298 N_A_317_461#_c_390_n N_A_596_419#_c_564_n 0.0248987f $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_299 N_A_317_461#_c_391_n N_A_596_419#_c_564_n 0.0170774f $X=3.025 $Y=1.56
+ $X2=0 $Y2=0
cc_300 N_A_317_461#_c_400_n N_VPWR_M1000_d 0.0140042f $X=2.65 $Y=2.39 $X2=0
+ $Y2=0
cc_301 N_A_317_461#_c_400_n N_VPWR_c_644_n 0.0261336f $X=2.65 $Y=2.39 $X2=0
+ $Y2=0
cc_302 N_A_317_461#_c_394_n N_VPWR_c_644_n 0.0223796f $X=1.71 $Y=2.45 $X2=0
+ $Y2=0
cc_303 N_A_317_461#_c_394_n N_VPWR_c_649_n 0.0136977f $X=1.71 $Y=2.45 $X2=0
+ $Y2=0
cc_304 N_A_317_461#_M1004_g N_VPWR_c_650_n 0.00136343f $X=3.43 $Y=2.305 $X2=0
+ $Y2=0
cc_305 N_A_317_461#_M1004_g N_VPWR_c_642_n 0.00128788f $X=3.43 $Y=2.305 $X2=0
+ $Y2=0
cc_306 N_A_317_461#_c_400_n N_VPWR_c_642_n 0.0195535f $X=2.65 $Y=2.39 $X2=0
+ $Y2=0
cc_307 N_A_317_461#_c_394_n N_VPWR_c_642_n 0.0106298f $X=1.71 $Y=2.45 $X2=0
+ $Y2=0
cc_308 N_A_317_461#_c_400_n A_524_419# 0.00145897f $X=2.65 $Y=2.39 $X2=-0.19
+ $Y2=-0.245
cc_309 N_A_317_461#_c_387_n N_VGND_M1001_d 0.00176891f $X=2.65 $Y=1.1 $X2=0
+ $Y2=0
cc_310 N_A_317_461#_M1017_g N_VGND_c_737_n 6.13277e-19 $X=2.935 $Y=0.835 $X2=0
+ $Y2=0
cc_311 N_A_317_461#_M1017_g N_VGND_c_741_n 0.00118999f $X=2.935 $Y=0.835 $X2=0
+ $Y2=0
cc_312 N_A_317_461#_c_387_n N_VGND_c_741_n 0.0188839f $X=2.65 $Y=1.1 $X2=0 $Y2=0
cc_313 N_A_317_461#_M1017_g N_VGND_c_746_n 9.49986e-19 $X=2.935 $Y=0.835 $X2=0
+ $Y2=0
cc_314 N_A_317_461#_c_387_n A_530_125# 0.00403907f $X=2.65 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_315 N_A_733_99#_M1006_g N_A_596_419#_M1013_g 0.0193113f $X=3.79 $Y=2.305
+ $X2=0 $Y2=0
cc_316 N_A_733_99#_c_475_n N_A_596_419#_M1013_g 0.00188269f $X=3.83 $Y=1.35
+ $X2=0 $Y2=0
cc_317 N_A_733_99#_c_497_p N_A_596_419#_M1013_g 0.0128565f $X=4.455 $Y=1.78
+ $X2=0 $Y2=0
cc_318 N_A_733_99#_c_487_n N_A_596_419#_M1013_g 0.00314257f $X=4.55 $Y=2.785
+ $X2=0 $Y2=0
cc_319 N_A_733_99#_c_479_n N_A_596_419#_M1013_g 0.00298797f $X=4.72 $Y=1.565
+ $X2=0 $Y2=0
cc_320 N_A_733_99#_c_480_n N_A_596_419#_M1013_g 0.00115689f $X=5.13 $Y=1.43
+ $X2=0 $Y2=0
cc_321 N_A_733_99#_M1016_d N_A_596_419#_c_597_n 0.00289746f $X=4.355 $Y=0.235
+ $X2=0 $Y2=0
cc_322 N_A_733_99#_M1002_g N_A_596_419#_c_597_n 0.0132635f $X=3.74 $Y=0.835
+ $X2=0 $Y2=0
cc_323 N_A_733_99#_c_475_n N_A_596_419#_c_597_n 0.0226f $X=3.83 $Y=1.35 $X2=0
+ $Y2=0
cc_324 N_A_733_99#_c_476_n N_A_596_419#_c_597_n 0.00112687f $X=3.83 $Y=1.35
+ $X2=0 $Y2=0
cc_325 N_A_733_99#_c_477_n N_A_596_419#_c_597_n 0.0173634f $X=4.72 $Y=1.265
+ $X2=0 $Y2=0
cc_326 N_A_733_99#_c_478_n N_A_596_419#_c_597_n 0.00440359f $X=4.72 $Y=0.455
+ $X2=0 $Y2=0
cc_327 N_A_733_99#_M1016_d N_A_596_419#_c_562_n 7.44962e-19 $X=4.355 $Y=0.235
+ $X2=0 $Y2=0
cc_328 N_A_733_99#_M1002_g N_A_596_419#_c_562_n 0.0010354f $X=3.74 $Y=0.835
+ $X2=0 $Y2=0
cc_329 N_A_733_99#_c_475_n N_A_596_419#_c_562_n 0.0205382f $X=3.83 $Y=1.35 $X2=0
+ $Y2=0
cc_330 N_A_733_99#_c_476_n N_A_596_419#_c_562_n 0.00115062f $X=3.83 $Y=1.35
+ $X2=0 $Y2=0
cc_331 N_A_733_99#_c_497_p N_A_596_419#_c_562_n 0.0149487f $X=4.455 $Y=1.78
+ $X2=0 $Y2=0
cc_332 N_A_733_99#_c_477_n N_A_596_419#_c_562_n 0.0197305f $X=4.72 $Y=1.265
+ $X2=0 $Y2=0
cc_333 N_A_733_99#_c_479_n N_A_596_419#_c_562_n 0.0204677f $X=4.72 $Y=1.565
+ $X2=0 $Y2=0
cc_334 N_A_733_99#_c_475_n N_A_596_419#_c_563_n 0.00114936f $X=3.83 $Y=1.35
+ $X2=0 $Y2=0
cc_335 N_A_733_99#_c_476_n N_A_596_419#_c_563_n 0.0201104f $X=3.83 $Y=1.35 $X2=0
+ $Y2=0
cc_336 N_A_733_99#_c_477_n N_A_596_419#_c_563_n 9.58238e-19 $X=4.72 $Y=1.265
+ $X2=0 $Y2=0
cc_337 N_A_733_99#_c_478_n N_A_596_419#_c_563_n 0.00210243f $X=4.72 $Y=0.455
+ $X2=0 $Y2=0
cc_338 N_A_733_99#_c_479_n N_A_596_419#_c_563_n 0.00554987f $X=4.72 $Y=1.565
+ $X2=0 $Y2=0
cc_339 N_A_733_99#_c_480_n N_A_596_419#_c_563_n 0.0057317f $X=5.13 $Y=1.43 $X2=0
+ $Y2=0
cc_340 N_A_733_99#_c_481_n N_A_596_419#_c_563_n 8.2258e-19 $X=5.162 $Y=1.265
+ $X2=0 $Y2=0
cc_341 N_A_733_99#_M1002_g N_A_596_419#_c_564_n 0.00590274f $X=3.74 $Y=0.835
+ $X2=0 $Y2=0
cc_342 N_A_733_99#_M1006_g N_A_596_419#_c_564_n 0.00392399f $X=3.79 $Y=2.305
+ $X2=0 $Y2=0
cc_343 N_A_733_99#_c_475_n N_A_596_419#_c_564_n 0.0340252f $X=3.83 $Y=1.35 $X2=0
+ $Y2=0
cc_344 N_A_733_99#_c_486_n N_A_596_419#_c_564_n 0.0121549f $X=3.995 $Y=1.78
+ $X2=0 $Y2=0
cc_345 N_A_733_99#_M1002_g N_A_596_419#_c_565_n 0.0181574f $X=3.74 $Y=0.835
+ $X2=0 $Y2=0
cc_346 N_A_733_99#_c_477_n N_A_596_419#_c_565_n 0.00683546f $X=4.72 $Y=1.265
+ $X2=0 $Y2=0
cc_347 N_A_733_99#_c_475_n N_VPWR_M1006_d 2.72261e-19 $X=3.83 $Y=1.35 $X2=0
+ $Y2=0
cc_348 N_A_733_99#_c_497_p N_VPWR_M1006_d 0.0104241f $X=4.455 $Y=1.78 $X2=0
+ $Y2=0
cc_349 N_A_733_99#_c_486_n N_VPWR_M1006_d 2.10259e-19 $X=3.995 $Y=1.78 $X2=0
+ $Y2=0
cc_350 N_A_733_99#_M1006_g N_VPWR_c_645_n 0.00786215f $X=3.79 $Y=2.305 $X2=0
+ $Y2=0
cc_351 N_A_733_99#_c_497_p N_VPWR_c_645_n 0.0186722f $X=4.455 $Y=1.78 $X2=0
+ $Y2=0
cc_352 N_A_733_99#_c_486_n N_VPWR_c_645_n 0.0035384f $X=3.995 $Y=1.78 $X2=0
+ $Y2=0
cc_353 N_A_733_99#_c_487_n N_VPWR_c_645_n 0.0348948f $X=4.55 $Y=2.785 $X2=0
+ $Y2=0
cc_354 N_A_733_99#_M1011_g N_VPWR_c_646_n 0.004243f $X=5.285 $Y=2.465 $X2=0
+ $Y2=0
cc_355 N_A_733_99#_c_487_n N_VPWR_c_646_n 0.021553f $X=4.55 $Y=2.785 $X2=0 $Y2=0
cc_356 N_A_733_99#_c_479_n N_VPWR_c_646_n 0.0241395f $X=4.72 $Y=1.565 $X2=0
+ $Y2=0
cc_357 N_A_733_99#_c_480_n N_VPWR_c_646_n 0.00187069f $X=5.13 $Y=1.43 $X2=0
+ $Y2=0
cc_358 N_A_733_99#_M1011_g N_VPWR_c_647_n 0.0175392f $X=5.285 $Y=2.465 $X2=0
+ $Y2=0
cc_359 N_A_733_99#_c_487_n N_VPWR_c_647_n 0.0571709f $X=4.55 $Y=2.785 $X2=0
+ $Y2=0
cc_360 N_A_733_99#_M1006_g N_VPWR_c_650_n 0.00327927f $X=3.79 $Y=2.305 $X2=0
+ $Y2=0
cc_361 N_A_733_99#_c_487_n N_VPWR_c_651_n 0.0102724f $X=4.55 $Y=2.785 $X2=0
+ $Y2=0
cc_362 N_A_733_99#_M1011_g N_VPWR_c_652_n 0.00564095f $X=5.285 $Y=2.465 $X2=0
+ $Y2=0
cc_363 N_A_733_99#_M1006_g N_VPWR_c_642_n 0.00419962f $X=3.79 $Y=2.305 $X2=0
+ $Y2=0
cc_364 N_A_733_99#_M1011_g N_VPWR_c_642_n 0.0104155f $X=5.285 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_A_733_99#_c_487_n N_VPWR_c_642_n 0.00935454f $X=4.55 $Y=2.785 $X2=0
+ $Y2=0
cc_366 N_A_733_99#_c_477_n N_Q_c_724_n 0.00457333f $X=4.72 $Y=1.265 $X2=0 $Y2=0
cc_367 N_A_733_99#_c_479_n N_Q_c_724_n 0.034843f $X=4.72 $Y=1.565 $X2=0 $Y2=0
cc_368 N_A_733_99#_c_481_n N_Q_c_724_n 0.0252283f $X=5.162 $Y=1.265 $X2=0 $Y2=0
cc_369 N_A_733_99#_M1002_g N_VGND_c_738_n 0.0035653f $X=3.74 $Y=0.835 $X2=0
+ $Y2=0
cc_370 N_A_733_99#_c_478_n N_VGND_c_739_n 0.0224947f $X=4.72 $Y=0.455 $X2=0
+ $Y2=0
cc_371 N_A_733_99#_c_477_n N_VGND_c_740_n 0.0356686f $X=4.72 $Y=1.265 $X2=0
+ $Y2=0
cc_372 N_A_733_99#_c_478_n N_VGND_c_740_n 0.0276101f $X=4.72 $Y=0.455 $X2=0
+ $Y2=0
cc_373 N_A_733_99#_c_479_n N_VGND_c_740_n 0.0171299f $X=4.72 $Y=1.565 $X2=0
+ $Y2=0
cc_374 N_A_733_99#_c_480_n N_VGND_c_740_n 0.00167931f $X=5.13 $Y=1.43 $X2=0
+ $Y2=0
cc_375 N_A_733_99#_c_481_n N_VGND_c_740_n 0.0146134f $X=5.162 $Y=1.265 $X2=0
+ $Y2=0
cc_376 N_A_733_99#_M1002_g N_VGND_c_744_n 0.00415323f $X=3.74 $Y=0.835 $X2=0
+ $Y2=0
cc_377 N_A_733_99#_c_481_n N_VGND_c_745_n 0.00489931f $X=5.162 $Y=1.265 $X2=0
+ $Y2=0
cc_378 N_A_733_99#_M1016_d N_VGND_c_746_n 0.00243792f $X=4.355 $Y=0.235 $X2=0
+ $Y2=0
cc_379 N_A_733_99#_M1002_g N_VGND_c_746_n 0.00469432f $X=3.74 $Y=0.835 $X2=0
+ $Y2=0
cc_380 N_A_733_99#_c_478_n N_VGND_c_746_n 0.0152094f $X=4.72 $Y=0.455 $X2=0
+ $Y2=0
cc_381 N_A_733_99#_c_481_n N_VGND_c_746_n 0.00961693f $X=5.162 $Y=1.265 $X2=0
+ $Y2=0
cc_382 N_A_596_419#_c_569_n N_VPWR_c_644_n 0.00169005f $X=3.18 $Y=2.24 $X2=0
+ $Y2=0
cc_383 N_A_596_419#_M1013_g N_VPWR_c_645_n 0.0156542f $X=4.335 $Y=2.305 $X2=0
+ $Y2=0
cc_384 N_A_596_419#_c_564_n N_VPWR_c_645_n 0.0253108f $X=3.237 $Y=2.075 $X2=0
+ $Y2=0
cc_385 N_A_596_419#_M1013_g N_VPWR_c_647_n 0.0030504f $X=4.335 $Y=2.305 $X2=0
+ $Y2=0
cc_386 N_A_596_419#_c_569_n N_VPWR_c_650_n 0.00998165f $X=3.18 $Y=2.24 $X2=0
+ $Y2=0
cc_387 N_A_596_419#_M1013_g N_VPWR_c_651_n 0.00465077f $X=4.335 $Y=2.305 $X2=0
+ $Y2=0
cc_388 N_A_596_419#_M1013_g N_VPWR_c_642_n 0.00451796f $X=4.335 $Y=2.305 $X2=0
+ $Y2=0
cc_389 N_A_596_419#_c_569_n N_VPWR_c_642_n 0.0139392f $X=3.18 $Y=2.24 $X2=0
+ $Y2=0
cc_390 N_A_596_419#_c_597_n N_VGND_M1002_d 0.0105973f $X=4.205 $Y=0.9 $X2=0
+ $Y2=0
cc_391 N_A_596_419#_c_597_n N_VGND_c_738_n 0.0218635f $X=4.205 $Y=0.9 $X2=0
+ $Y2=0
cc_392 N_A_596_419#_c_565_n N_VGND_c_738_n 0.0132002f $X=4.37 $Y=1.185 $X2=0
+ $Y2=0
cc_393 N_A_596_419#_c_565_n N_VGND_c_739_n 0.00486043f $X=4.37 $Y=1.185 $X2=0
+ $Y2=0
cc_394 N_A_596_419#_c_565_n N_VGND_c_740_n 0.00299613f $X=4.37 $Y=1.185 $X2=0
+ $Y2=0
cc_395 N_A_596_419#_c_571_n N_VGND_c_741_n 0.00182539f $X=3.29 $Y=0.9 $X2=0
+ $Y2=0
cc_396 N_A_596_419#_c_571_n N_VGND_c_746_n 0.00943433f $X=3.29 $Y=0.9 $X2=0
+ $Y2=0
cc_397 N_A_596_419#_c_597_n N_VGND_c_746_n 0.0229653f $X=4.205 $Y=0.9 $X2=0
+ $Y2=0
cc_398 N_A_596_419#_c_576_n N_VGND_c_746_n 0.00569693f $X=3.375 $Y=0.9 $X2=0
+ $Y2=0
cc_399 N_A_596_419#_c_565_n N_VGND_c_746_n 0.00592249f $X=4.37 $Y=1.185 $X2=0
+ $Y2=0
cc_400 N_A_596_419#_c_597_n A_691_125# 0.00566125f $X=4.205 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_401 N_VPWR_c_642_n N_Q_M1011_d 0.00302127f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_402 N_VPWR_c_646_n N_Q_c_724_n 0.0144811f $X=5.06 $Y=2.19 $X2=0 $Y2=0
cc_403 N_VPWR_c_652_n N_Q_c_724_n 0.0192376f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_404 N_VPWR_c_642_n N_Q_c_724_n 0.0111968f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_405 N_Q_c_724_n N_VGND_c_740_n 0.0293631f $X=5.5 $Y=0.46 $X2=0 $Y2=0
cc_406 N_Q_c_724_n N_VGND_c_745_n 0.0164655f $X=5.5 $Y=0.46 $X2=0 $Y2=0
cc_407 N_Q_c_724_n N_VGND_c_746_n 0.0109746f $X=5.5 $Y=0.46 $X2=0 $Y2=0
