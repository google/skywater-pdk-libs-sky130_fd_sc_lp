* File: sky130_fd_sc_lp__maj3_2.pex.spice
* Created: Fri Aug 28 10:43:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MAJ3_2%C 3 7 11 15 19 20 23 24 27 28 29 35 39 45 47
c89 20 0 1.40829e-19 $X=0.605 $Y=1.935
c90 15 0 1.37614e-19 $X=2.725 $Y=0.455
r91 39 47 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=2.07 $X2=2.64
+ $Y2=2.07
r92 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=2.07
+ $X2=2.745 $Y2=2.235
r93 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=2.07
+ $X2=2.745 $Y2=1.905
r94 28 47 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=2.622 $Y=2.07
+ $X2=2.64 $Y2=2.07
r95 28 45 6.08745 $w=3.28e-07 $l=9.7e-08 $layer=LI1_cond $X=2.622 $Y=2.07
+ $X2=2.525 $Y2=2.07
r96 28 29 14.423 $w=3.28e-07 $l=4.13e-07 $layer=LI1_cond $X=2.707 $Y=2.07
+ $X2=3.12 $Y2=2.07
r97 28 39 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=2.707 $Y=2.07
+ $X2=2.69 $Y2=2.07
r98 28 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.745
+ $Y=2.07 $X2=2.745 $Y2=2.07
r99 27 45 114.497 $w=1.68e-07 $l=1.755e-06 $layer=LI1_cond $X=0.77 $Y=2.15
+ $X2=2.525 $Y2=2.15
r100 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.43 $X2=0.605 $Y2=1.43
r101 21 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.605 $Y=2.065
+ $X2=0.77 $Y2=2.15
r102 21 23 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.605 $Y=2.065
+ $X2=0.605 $Y2=1.43
r103 19 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.605 $Y=1.77
+ $X2=0.605 $Y2=1.43
r104 19 20 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.77
+ $X2=0.605 $Y2=1.935
r105 18 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.265
+ $X2=0.605 $Y2=1.43
r106 15 37 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=2.725 $Y=0.455
+ $X2=2.725 $Y2=1.905
r107 11 38 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.685 $Y=2.775
+ $X2=2.685 $Y2=2.235
r108 7 18 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.695 $Y=0.455
+ $X2=0.695 $Y2=1.265
r109 3 20 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.655 $Y=2.775
+ $X2=0.655 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_2%A 3 7 13 17 19 20 21 22 26
r56 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.25
+ $Y=1.38 $X2=1.25 $Y2=1.38
r57 22 27 7.67632 $w=6.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.68 $Y=1.55
+ $X2=1.25 $Y2=1.55
r58 21 27 0.892596 $w=6.68e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=1.55 $X2=1.25
+ $Y2=1.55
r59 19 20 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.065 $Y=2.175
+ $X2=1.065 $Y2=2.325
r60 15 26 31.1986 $w=2.74e-07 $l=2.85832e-07 $layer=POLY_cond $X=1.515 $Y=1.215
+ $X2=1.3 $Y2=1.38
r61 15 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.515 $Y=1.215
+ $X2=1.515 $Y2=0.455
r62 11 26 91.0088 $w=2.74e-07 $l=5.86003e-07 $layer=POLY_cond $X=1.475 $Y=1.885
+ $X2=1.3 $Y2=1.38
r63 11 13 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.475 $Y=1.885
+ $X2=1.475 $Y2=2.775
r64 9 26 91.0088 $w=2.74e-07 $l=6.02993e-07 $layer=POLY_cond $X=1.085 $Y=1.885
+ $X2=1.3 $Y2=1.38
r65 9 19 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.085 $Y=1.885
+ $X2=1.085 $Y2=2.175
r66 5 26 31.1986 $w=2.74e-07 $l=2.85832e-07 $layer=POLY_cond $X=1.085 $Y=1.215
+ $X2=1.3 $Y2=1.38
r67 5 7 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.085 $Y=1.215
+ $X2=1.085 $Y2=0.455
r68 3 20 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.045 $Y=2.775
+ $X2=1.045 $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_2%B 1 3 7 11 15 22 23 26 27
r56 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.145
+ $Y=1.38 $X2=2.145 $Y2=1.38
r57 23 27 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.145 $Y=1.665
+ $X2=2.145 $Y2=1.38
r58 22 26 1.48619 $w=5.4e-07 $l=1.5e-08 $layer=POLY_cond $X=2.1 $Y=1.365 $X2=2.1
+ $Y2=1.38
r59 18 26 35.1732 $w=5.4e-07 $l=3.55e-07 $layer=POLY_cond $X=2.1 $Y=1.735
+ $X2=2.1 $Y2=1.38
r60 5 22 25.3483 $w=5.4e-07 $l=1.5e-07 $layer=POLY_cond $X=2.12 $Y=1.215
+ $X2=2.12 $Y2=1.365
r61 5 15 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.335 $Y=1.215
+ $X2=2.335 $Y2=0.455
r62 5 7 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.905 $Y=1.215
+ $X2=1.905 $Y2=0.455
r63 1 18 25.3483 $w=5.4e-07 $l=1.5e-07 $layer=POLY_cond $X=2.08 $Y=1.885
+ $X2=2.08 $Y2=1.735
r64 1 11 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2.295 $Y=1.885
+ $X2=2.295 $Y2=2.775
r65 1 3 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.865 $Y=1.885
+ $X2=1.865 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_2%A_59_491# 1 2 3 4 15 19 23 27 30 33 35 37 38
+ 41 45 47 50 58 59 63 69
c134 69 0 2.91364e-20 $X=3.665 $Y=1.435
c135 35 0 1.40829e-19 $X=1.915 $Y=2.5
r136 68 69 55.8541 $w=2.33e-07 $l=2.7e-07 $layer=POLY_cond $X=3.395 $Y=1.435
+ $X2=3.665 $Y2=1.435
r137 64 68 27.927 $w=2.33e-07 $l=1.35e-07 $layer=POLY_cond $X=3.26 $Y=1.435
+ $X2=3.395 $Y2=1.435
r138 64 66 5.17167 $w=2.33e-07 $l=2.5e-08 $layer=POLY_cond $X=3.26 $Y=1.435
+ $X2=3.235 $Y2=1.435
r139 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.26
+ $Y=1.45 $X2=3.26 $Y2=1.45
r140 60 63 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.02 $Y=1.45
+ $X2=3.26 $Y2=1.45
r141 57 58 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=2.74
+ $X2=0.605 $Y2=2.74
r142 54 57 4.87632 $w=6.48e-07 $l=2.65e-07 $layer=LI1_cond $X=0.175 $Y=2.74
+ $X2=0.44 $Y2=2.74
r143 50 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=1.285
+ $X2=3.02 $Y2=1.45
r144 49 50 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.02 $Y=1.035
+ $X2=3.02 $Y2=1.285
r145 48 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=0.95
+ $X2=2.12 $Y2=0.95
r146 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.935 $Y=0.95
+ $X2=3.02 $Y2=1.035
r147 47 48 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.935 $Y=0.95
+ $X2=2.285 $Y2=0.95
r148 43 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=0.865
+ $X2=2.12 $Y2=0.95
r149 43 45 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.12 $Y=0.865
+ $X2=2.12 $Y2=0.475
r150 39 41 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.08 $Y=2.585
+ $X2=2.08 $Y2=2.74
r151 37 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0.95
+ $X2=2.12 $Y2=0.95
r152 37 38 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.955 $Y=0.95
+ $X2=0.645 $Y2=0.95
r153 35 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.915 $Y=2.5
+ $X2=2.08 $Y2=2.585
r154 35 58 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.915 $Y=2.5
+ $X2=0.605 $Y2=2.5
r155 31 38 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.48 $Y=0.95
+ $X2=0.645 $Y2=0.95
r156 31 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.48 $Y=0.95
+ $X2=0.175 $Y2=0.95
r157 31 33 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.48 $Y=0.865
+ $X2=0.48 $Y2=0.475
r158 30 54 8.83581 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=0.175 $Y=2.415
+ $X2=0.175 $Y2=2.74
r159 29 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=1.035
+ $X2=0.175 $Y2=0.95
r160 29 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.175 $Y=1.035
+ $X2=0.175 $Y2=2.415
r161 25 69 33.0987 $w=2.33e-07 $l=1.6e-07 $layer=POLY_cond $X=3.825 $Y=1.435
+ $X2=3.665 $Y2=1.435
r162 25 27 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=3.825 $Y=1.435
+ $X2=3.825 $Y2=2.465
r163 21 69 13.0941 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.665 $Y=1.285
+ $X2=3.665 $Y2=1.435
r164 21 23 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.665 $Y=1.285
+ $X2=3.665 $Y2=0.665
r165 17 68 13.0941 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.395 $Y=1.615
+ $X2=3.395 $Y2=1.435
r166 17 19 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=3.395 $Y=1.615
+ $X2=3.395 $Y2=2.465
r167 13 66 13.0941 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.235 $Y=1.285
+ $X2=3.235 $Y2=1.435
r168 13 15 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.235 $Y=1.285
+ $X2=3.235 $Y2=0.665
r169 4 41 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=2.455 $X2=2.08 $Y2=2.74
r170 3 57 600 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_PDIFF $count=1 $X=0.295
+ $Y=2.455 $X2=0.44 $Y2=2.74
r171 2 45 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.245 $X2=2.12 $Y2=0.475
r172 1 33 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=0.335
+ $Y=0.245 $X2=0.48 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_2%VPWR 1 2 3 12 16 18 20 25 26 27 29 41 46 50
r61 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r63 44 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r65 41 49 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=4.137 $Y2=3.33
r66 41 43 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=3.6 $Y2=3.33
r67 40 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r68 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 37 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r71 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.26 $Y2=3.33
r73 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 32 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r75 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.26 $Y2=3.33
r77 29 31 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 27 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r79 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r80 25 39 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.9 $Y2=3.33
r82 24 43 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=3.6 $Y2=3.33
r83 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=2.9 $Y2=3.33
r84 20 23 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=4.08 $Y=1.96
+ $X2=4.08 $Y2=2.93
r85 18 49 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.137 $Y2=3.33
r86 18 23 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.08 $Y2=2.93
r87 14 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=3.245 $X2=2.9
+ $Y2=3.33
r88 14 16 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=2.9 $Y=3.245
+ $X2=2.9 $Y2=2.58
r89 10 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=3.245
+ $X2=1.26 $Y2=3.33
r90 10 12 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.26 $Y=3.245
+ $X2=1.26 $Y2=2.93
r91 3 23 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=1.835 $X2=4.04 $Y2=2.93
r92 3 20 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=1.835 $X2=4.04 $Y2=1.96
r93 2 16 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.76
+ $Y=2.455 $X2=2.9 $Y2=2.58
r94 1 12 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=2.455 $X2=1.26 $Y2=2.93
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_2%X 1 2 9 11 15 16 17 23 29
c36 29 0 1.37614e-19 $X=3.6 $Y=0.925
r37 21 29 1.58663 $w=4.88e-07 $l=6.5e-08 $layer=LI1_cond $X=3.53 $Y=0.86
+ $X2=3.53 $Y2=0.925
r38 17 31 9.57828 $w=4.88e-07 $l=1.7e-07 $layer=LI1_cond $X=3.53 $Y=0.935
+ $X2=3.53 $Y2=1.105
r39 17 29 0.244098 $w=4.88e-07 $l=1e-08 $layer=LI1_cond $X=3.53 $Y=0.935
+ $X2=3.53 $Y2=0.925
r40 17 21 0.244098 $w=4.88e-07 $l=1e-08 $layer=LI1_cond $X=3.53 $Y=0.85 $X2=3.53
+ $Y2=0.86
r41 16 17 7.20088 $w=4.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3.53 $Y=0.555
+ $X2=3.53 $Y2=0.85
r42 16 23 3.05122 $w=4.88e-07 $l=1.25e-07 $layer=LI1_cond $X=3.53 $Y=0.555
+ $X2=3.53 $Y2=0.43
r43 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.69 $Y=1.795
+ $X2=3.69 $Y2=1.105
r44 9 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.61 $Y=1.96
+ $X2=3.61 $Y2=1.795
r45 9 11 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=3.61 $Y=1.96 $X2=3.61
+ $Y2=2.9
r46 2 11 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.835 $X2=3.61 $Y2=2.9
r47 2 9 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.835 $X2=3.61 $Y2=1.96
r48 1 23 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.31
+ $Y=0.245 $X2=3.45 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_2%VGND 1 2 3 12 16 18 20 23 24 25 27 39 44 48
c55 16 0 2.91364e-20 $X=2.94 $Y=0.455
r56 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r57 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r58 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r59 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r60 39 47 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.955 $Y=0 $X2=4.137
+ $Y2=0
r61 39 41 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=0 $X2=3.6
+ $Y2=0
r62 38 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r63 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r64 35 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r65 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r66 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r67 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.3
+ $Y2=0
r68 32 34 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.68
+ $Y2=0
r69 30 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r70 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r71 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.3
+ $Y2=0
r72 27 29 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.24
+ $Y2=0
r73 25 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r74 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r75 23 37 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.64
+ $Y2=0
r76 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.94
+ $Y2=0
r77 22 41 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.6
+ $Y2=0
r78 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=2.94
+ $Y2=0
r79 18 47 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.08 $Y=0.085
+ $X2=4.137 $Y2=0
r80 18 20 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=4.08 $Y=0.085
+ $X2=4.08 $Y2=0.39
r81 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0
r82 14 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0.455
r83 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=0.085 $X2=1.3
+ $Y2=0
r84 10 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.3 $Y=0.085 $X2=1.3
+ $Y2=0.455
r85 3 20 91 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_NDIFF $count=2 $X=3.74
+ $Y=0.245 $X2=4.04 $Y2=0.39
r86 2 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.245 $X2=2.94 $Y2=0.455
r87 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.245 $X2=1.3 $Y2=0.455
.ends

