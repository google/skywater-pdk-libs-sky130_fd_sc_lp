* File: sky130_fd_sc_lp__and3_lp.pex.spice
* Created: Fri Aug 28 10:06:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3_LP%A 1 2 3 5 9 17 18 22 23
c40 1 0 7.37982e-20 $X=0.63 $Y=0.885
r41 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.02 $X2=0.27 $Y2=1.02
r42 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.665
r43 17 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.02
r44 13 22 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.27 $Y=1.375
+ $X2=0.27 $Y2=1.02
r45 11 22 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.27 $Y=0.96 $X2=0.27
+ $Y2=1.02
r46 7 9 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.705 $Y=0.81
+ $X2=0.705 $Y2=0.445
r47 3 13 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.6 $Y=1.45 $X2=0.27
+ $Y2=1.45
r48 3 5 262.119 $w=2.5e-07 $l=1.055e-06 $layer=POLY_cond $X=0.6 $Y=1.525 $X2=0.6
+ $Y2=2.58
r49 2 11 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=0.885
+ $X2=0.27 $Y2=0.96
r50 1 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.63 $Y=0.885
+ $X2=0.705 $Y2=0.81
r51 1 2 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.63 $Y=0.885
+ $X2=0.435 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_LP%B 1 3 7 11 12 15 16
r46 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.13
+ $Y=1.365 $X2=1.13 $Y2=1.365
r47 12 16 9.87808 $w=3.48e-07 $l=3e-07 $layer=LI1_cond $X=1.14 $Y=1.665 $X2=1.14
+ $Y2=1.365
r48 11 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.13 $Y=1.705
+ $X2=1.13 $Y2=1.365
r49 10 15 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.2
+ $X2=1.13 $Y2=1.365
r50 7 10 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.095 $Y=0.445
+ $X2=1.095 $Y2=1.2
r51 1 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.87
+ $X2=1.13 $Y2=1.705
r52 1 3 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.13 $Y=1.87 $X2=1.13
+ $Y2=2.58
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_LP%C 1 3 8 12 15 16 17 18 21 22
c49 1 0 1.11641e-19 $X=1.485 $Y=0.73
r50 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.7
+ $Y=1.365 $X2=1.7 $Y2=1.365
r51 18 22 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.7 $Y=1.665 $X2=1.7
+ $Y2=1.365
r52 16 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.7 $Y=1.705 $X2=1.7
+ $Y2=1.365
r53 16 17 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.705
+ $X2=1.7 $Y2=1.87
r54 15 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.2 $X2=1.7
+ $Y2=1.365
r55 10 12 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.485 $Y=0.805
+ $X2=1.61 $Y2=0.805
r56 8 17 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.66 $Y=2.58 $X2=1.66
+ $Y2=1.87
r57 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.61 $Y=0.88 $X2=1.61
+ $Y2=0.805
r58 4 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.61 $Y=0.88 $X2=1.61
+ $Y2=1.2
r59 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.485 $Y=0.73
+ $X2=1.485 $Y2=0.805
r60 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.485 $Y=0.73 $X2=1.485
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_LP%A_38_416# 1 2 3 12 16 20 26 29 32 35 37 38
+ 40 41 44 54 56 58 59
c102 54 0 7.37982e-20 $X=0.7 $Y=0.47
r103 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.27
+ $Y=1.015 $X2=2.27 $Y2=1.015
r104 52 54 5.90276 $w=4.08e-07 $l=2.1e-07 $layer=LI1_cond $X=0.49 $Y=0.47
+ $X2=0.7 $Y2=0.47
r105 42 44 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.395 $Y=2.22
+ $X2=1.395 $Y2=2.225
r106 41 50 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=2.135
+ $X2=0.7 $Y2=2.135
r107 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.23 $Y=2.135
+ $X2=1.395 $Y2=2.22
r108 40 41 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.23 $Y=2.135
+ $X2=0.785 $Y2=2.135
r109 39 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.935
+ $X2=0.7 $Y2=0.935
r110 38 58 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=0.935
+ $X2=2.27 $Y2=0.935
r111 38 39 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=2.105 $Y=0.935
+ $X2=0.785 $Y2=0.935
r112 37 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.05 $X2=0.7
+ $Y2=2.135
r113 36 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.02 $X2=0.7
+ $Y2=0.935
r114 36 37 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.7 $Y=1.02
+ $X2=0.7 $Y2=2.05
r115 35 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.85 $X2=0.7
+ $Y2=0.935
r116 34 54 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.7 $Y=0.675
+ $X2=0.7 $Y2=0.47
r117 34 35 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.7 $Y=0.675
+ $X2=0.7 $Y2=0.85
r118 30 50 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.335 $Y=2.135
+ $X2=0.7 $Y2=2.135
r119 30 32 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.335 $Y=2.22
+ $X2=0.335 $Y2=2.225
r120 28 59 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.27 $Y=1.355
+ $X2=2.27 $Y2=1.015
r121 28 29 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.355
+ $X2=2.27 $Y2=1.52
r122 25 59 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.27 $Y=0.96
+ $X2=2.27 $Y2=1.015
r123 25 26 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.27 $Y=0.885
+ $X2=2.36 $Y2=0.885
r124 22 25 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2 $Y=0.885 $X2=2.27
+ $Y2=0.885
r125 18 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=0.81
+ $X2=2.36 $Y2=0.885
r126 18 20 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.36 $Y=0.81
+ $X2=2.36 $Y2=0.445
r127 16 29 263.361 $w=2.5e-07 $l=1.06e-06 $layer=POLY_cond $X=2.23 $Y=2.58
+ $X2=2.23 $Y2=1.52
r128 10 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2 $Y=0.81 $X2=2
+ $Y2=0.885
r129 10 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2 $Y=0.81 $X2=2
+ $Y2=0.445
r130 3 44 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.255
+ $Y=2.08 $X2=1.395 $Y2=2.225
r131 2 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.19
+ $Y=2.08 $X2=0.335 $Y2=2.225
r132 1 52 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.345
+ $Y=0.235 $X2=0.49 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_LP%VPWR 1 2 11 15 20 21 22 29 30 33
r37 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 27 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=0.865 $Y2=3.33
r42 24 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 22 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 22 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 20 26 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.76 $Y=3.33 $X2=1.68
+ $Y2=3.33
r46 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.76 $Y=3.33
+ $X2=1.925 $Y2=3.33
r47 19 29 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.09 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=3.33
+ $X2=1.925 $Y2=3.33
r49 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.925 $Y=2.225
+ $X2=1.925 $Y2=2.935
r50 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.925 $Y=3.245
+ $X2=1.925 $Y2=3.33
r51 13 18 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.925 $Y=3.245
+ $X2=1.925 $Y2=2.935
r52 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=3.33
r53 9 11 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=2.565
r54 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.785
+ $Y=2.08 $X2=1.925 $Y2=2.935
r55 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.785
+ $Y=2.08 $X2=1.925 $Y2=2.225
r56 1 11 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=0.725
+ $Y=2.08 $X2=0.865 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_LP%X 1 2 9 12 13 14 15 19
c29 19 0 1.11641e-19 $X=2.615 $Y=0.467
r30 15 19 2.48344 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=0.467
+ $X2=2.615 $Y2=0.467
r31 15 19 0.853661 $w=4.03e-07 $l=3e-08 $layer=LI1_cond $X=2.585 $Y=0.467
+ $X2=2.615 $Y2=0.467
r32 15 24 0.284554 $w=4.03e-07 $l=1e-08 $layer=LI1_cond $X=2.585 $Y=0.467
+ $X2=2.575 $Y2=0.467
r33 14 24 11.809 $w=4.03e-07 $l=4.15e-07 $layer=LI1_cond $X=2.16 $Y=0.467
+ $X2=2.575 $Y2=0.467
r34 12 13 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.557 $Y=2.225
+ $X2=2.557 $Y2=2.06
r35 9 15 5.93104 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=2.7 $Y=0.67 $X2=2.7
+ $Y2=0.467
r36 9 13 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=2.7 $Y=0.67 $X2=2.7
+ $Y2=2.06
r37 2 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=2.08 $X2=2.495 $Y2=2.225
r38 1 24 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.235 $X2=2.575 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_LP%VGND 1 6 8 10 20 21 24
r35 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r36 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r37 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.7
+ $Y2=0
r39 18 20 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.64
+ $Y2=0
r40 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 13 17 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r42 12 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r43 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.7
+ $Y2=0
r45 10 16 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.2
+ $Y2=0
r46 8 25 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r47 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r48 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r49 4 6 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0.44
r50 1 6 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.7 $Y2=0.44
.ends

