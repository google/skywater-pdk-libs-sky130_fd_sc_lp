* File: sky130_fd_sc_lp__sdfstp_1.pex.spice
* Created: Fri Aug 28 11:29:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%SCD 3 7 9 10 11 12 13 17
r30 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.455
+ $Y=1.335 $X2=0.455 $Y2=1.335
r31 13 18 8.4883 $w=4.63e-07 $l=3.3e-07 $layer=LI1_cond $X=0.387 $Y=1.665
+ $X2=0.387 $Y2=1.335
r32 12 18 1.02888 $w=4.63e-07 $l=4e-08 $layer=LI1_cond $X=0.387 $Y=1.295
+ $X2=0.387 $Y2=1.335
r33 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.455 $Y=1.675
+ $X2=0.455 $Y2=1.335
r34 10 11 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.455 $Y=1.675
+ $X2=0.455 $Y2=1.84
r35 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.455 $Y=1.17
+ $X2=0.455 $Y2=1.335
r36 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.545 $Y=0.85
+ $X2=0.545 $Y2=1.17
r37 3 11 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.475 $Y=2.36
+ $X2=0.475 $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%D 3 7 9 10 11 16
r37 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.695
+ $X2=1.355 $Y2=1.86
r38 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.695
+ $X2=1.355 $Y2=1.53
r39 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.355
+ $Y=1.695 $X2=1.355 $Y2=1.695
r40 10 11 17.8443 $w=3.08e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.685
+ $X2=2.16 $Y2=1.685
r41 10 17 12.0821 $w=3.08e-07 $l=3.25e-07 $layer=LI1_cond $X=1.68 $Y=1.685
+ $X2=1.355 $Y2=1.685
r42 9 17 5.76222 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=1.685
+ $X2=1.355 $Y2=1.685
r43 7 18 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.335 $Y=0.85
+ $X2=1.335 $Y2=1.53
r44 3 19 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.265 $Y=2.36 $X2=1.265
+ $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_324_102# 1 2 7 9 10 12 14 17 24 25 26 27
+ 30
c81 30 0 8.09203e-20 $X=3.32 $Y=2.56
r82 28 30 41.2735 $w=2.13e-07 $l=7.7e-07 $layer=LI1_cond $X=3.332 $Y=1.79
+ $X2=3.332 $Y2=2.56
r83 26 28 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.225 $Y=1.705
+ $X2=3.332 $Y2=1.79
r84 26 27 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.225 $Y=1.705
+ $X2=3.025 $Y2=1.705
r85 25 34 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.86 $Y=1.285
+ $X2=2.86 $Y2=1.505
r86 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.86
+ $Y=1.285 $X2=2.86 $Y2=1.285
r87 22 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.895 $Y=1.62
+ $X2=3.025 $Y2=1.705
r88 22 24 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=2.895 $Y=1.62
+ $X2=2.895 $Y2=1.285
r89 21 24 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=2.895 $Y=1.02
+ $X2=2.895 $Y2=1.285
r90 17 21 6.91731 $w=2.1e-07 $l=1.74786e-07 $layer=LI1_cond $X=2.765 $Y=0.915
+ $X2=2.895 $Y2=1.02
r91 17 19 20.3333 $w=2.08e-07 $l=3.85e-07 $layer=LI1_cond $X=2.765 $Y=0.915
+ $X2=2.38 $Y2=0.915
r92 15 16 8.39207 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=1.88 $Y=1.505
+ $X2=1.75 $Y2=1.505
r93 14 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.505
+ $X2=2.86 $Y2=1.505
r94 14 15 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.695 $Y=1.505
+ $X2=1.88 $Y2=1.505
r95 10 16 21.2973 $w=1.9e-07 $l=9.87421e-08 $layer=POLY_cond $X=1.805 $Y=1.58
+ $X2=1.75 $Y2=1.505
r96 10 12 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.805 $Y=1.58
+ $X2=1.805 $Y2=2.36
r97 7 16 87.2552 $w=1.9e-07 $l=3.61455e-07 $layer=POLY_cond $X=1.695 $Y=1.17
+ $X2=1.75 $Y2=1.505
r98 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.695 $Y=1.17
+ $X2=1.695 $Y2=0.85
r99 2 30 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=2.405 $X2=3.32 $Y2=2.56
r100 1 19 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.64 $X2=2.38 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%SCE 3 5 7 8 11 13 16 17 18 21 24 25 28 30
+ 31 34
r89 37 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.78 $Y=0.35
+ $X2=2.78 $Y2=0.515
r90 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=0.35 $X2=2.78 $Y2=0.35
r91 34 37 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.78 $Y=0.195
+ $X2=2.78 $Y2=0.35
r92 31 38 10.4488 $w=3.73e-07 $l=3.4e-07 $layer=LI1_cond $X=3.12 $Y=0.452
+ $X2=2.78 $Y2=0.452
r93 30 38 4.30245 $w=3.73e-07 $l=1.4e-07 $layer=LI1_cond $X=2.64 $Y=0.452
+ $X2=2.78 $Y2=0.452
r94 26 28 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.105 $Y=2.105
+ $X2=3.34 $Y2=2.105
r95 24 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.34 $Y=2.03
+ $X2=3.34 $Y2=2.105
r96 23 24 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=3.34 $Y=0.88
+ $X2=3.34 $Y2=2.03
r97 19 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.105 $Y=2.18
+ $X2=3.105 $Y2=2.105
r98 19 21 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.105 $Y=2.18
+ $X2=3.105 $Y2=2.725
r99 17 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.265 $Y=0.805
+ $X2=3.34 $Y2=0.88
r100 17 18 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.265 $Y=0.805
+ $X2=2.945 $Y2=0.805
r101 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.87 $Y=0.73
+ $X2=2.945 $Y2=0.805
r102 16 39 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.87 $Y=0.73
+ $X2=2.87 $Y2=0.515
r103 14 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.24 $Y=0.195
+ $X2=2.165 $Y2=0.195
r104 13 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=0.195
+ $X2=2.78 $Y2=0.195
r105 13 14 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.615 $Y=0.195
+ $X2=2.24 $Y2=0.195
r106 9 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.165 $Y=0.27
+ $X2=2.165 $Y2=0.195
r107 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.165 $Y=0.27
+ $X2=2.165 $Y2=0.85
r108 7 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.09 $Y=0.195
+ $X2=2.165 $Y2=0.195
r109 7 8 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=2.09 $Y=0.195
+ $X2=0.98 $Y2=0.195
r110 3 5 774.277 $w=1.5e-07 $l=1.51e-06 $layer=POLY_cond $X=0.905 $Y=0.85
+ $X2=0.905 $Y2=2.36
r111 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=0.27
+ $X2=0.98 $Y2=0.195
r112 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.905 $Y=0.27
+ $X2=0.905 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%CLK 3 7 9 10 11 16
c41 16 0 8.09203e-20 $X=4.08 $Y=1.32
r42 16 19 83.3779 $w=4.9e-07 $l=5.05e-07 $layer=POLY_cond $X=4.02 $Y=1.32
+ $X2=4.02 $Y2=1.825
r43 16 18 46.2534 $w=4.9e-07 $l=1.65e-07 $layer=POLY_cond $X=4.02 $Y=1.32
+ $X2=4.02 $Y2=1.155
r44 10 11 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=4.117 $Y=1.295
+ $X2=4.117 $Y2=1.665
r45 10 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.08
+ $Y=1.32 $X2=4.08 $Y2=1.32
r46 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=4.117 $Y=0.925
+ $X2=4.117 $Y2=1.295
r47 7 19 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.19 $Y=2.735
+ $X2=4.19 $Y2=1.825
r48 3 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.85 $Y=0.445
+ $X2=3.85 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_871_47# 1 2 9 13 17 21 23 25 29 34 35 38
+ 39 42 43 44 46 48 49 55 59 61 63 74
c173 61 0 1.0162e-19 $X=9.305 $Y=1.93
c174 48 0 1.35269e-19 $X=7.8 $Y=1.9
c175 46 0 1.76739e-19 $X=7.715 $Y=2.84
c176 44 0 6.84876e-20 $X=7.06 $Y=2.925
r177 73 74 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=9.485 $Y=1.93
+ $X2=9.52 $Y2=1.93
r178 67 68 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.6 $Y=1.68
+ $X2=6.03 $Y2=1.68
r179 62 73 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=9.305 $Y=1.93
+ $X2=9.485 $Y2=1.93
r180 61 63 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=9.305 $Y=1.96
+ $X2=9.14 $Y2=1.96
r181 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.305
+ $Y=1.93 $X2=9.305 $Y2=1.93
r182 55 57 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=4.87 $Y=2.86 $X2=4.87
+ $Y2=2.95
r183 49 52 3.77524 $w=2.88e-07 $l=9.5e-08 $layer=LI1_cond $X=4.515 $Y=0.35
+ $X2=4.515 $Y2=0.445
r184 48 63 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=7.8 $Y=1.9
+ $X2=9.14 $Y2=1.9
r185 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.715 $Y=1.985
+ $X2=7.8 $Y2=1.9
r186 45 46 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=7.715 $Y=1.985
+ $X2=7.715 $Y2=2.84
r187 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.63 $Y=2.925
+ $X2=7.715 $Y2=2.84
r188 43 44 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.63 $Y=2.925
+ $X2=7.06 $Y2=2.925
r189 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.975 $Y=2.84
+ $X2=7.06 $Y2=2.925
r190 41 42 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.975 $Y=2.115
+ $X2=6.975 $Y2=2.84
r191 40 59 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.41 $Y=2.03
+ $X2=6.245 $Y2=2.03
r192 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.89 $Y=2.03
+ $X2=6.975 $Y2=2.115
r193 39 40 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.89 $Y=2.03
+ $X2=6.41 $Y2=2.03
r194 37 59 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.165 $Y=2.115
+ $X2=6.245 $Y2=2.03
r195 37 38 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=6.165 $Y=2.115
+ $X2=6.165 $Y2=2.865
r196 35 68 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.245 $Y=1.68
+ $X2=6.03 $Y2=1.68
r197 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.245
+ $Y=1.68 $X2=6.245 $Y2=1.68
r198 32 59 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.245 $Y=1.945
+ $X2=6.245 $Y2=2.03
r199 32 34 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=6.245 $Y=1.945
+ $X2=6.245 $Y2=1.68
r200 30 67 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.465 $Y=1.68
+ $X2=5.6 $Y2=1.68
r201 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.465
+ $Y=1.68 $X2=5.465 $Y2=1.68
r202 27 29 76.7121 $w=1.78e-07 $l=1.245e-06 $layer=LI1_cond $X=5.46 $Y=0.435
+ $X2=5.46 $Y2=1.68
r203 26 57 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5 $Y=2.95 $X2=4.87
+ $Y2=2.95
r204 25 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.08 $Y=2.95
+ $X2=6.165 $Y2=2.865
r205 25 26 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=6.08 $Y=2.95 $X2=5
+ $Y2=2.95
r206 24 49 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.66 $Y=0.35
+ $X2=4.515 $Y2=0.35
r207 23 27 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.37 $Y=0.35
+ $X2=5.46 $Y2=0.435
r208 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.37 $Y=0.35
+ $X2=4.66 $Y2=0.35
r209 19 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.52 $Y=1.765
+ $X2=9.52 $Y2=1.93
r210 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=9.52 $Y=1.765
+ $X2=9.52 $Y2=0.945
r211 15 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.485 $Y=2.095
+ $X2=9.485 $Y2=1.93
r212 15 17 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.485 $Y=2.095
+ $X2=9.485 $Y2=2.525
r213 11 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.515
+ $X2=6.03 $Y2=1.68
r214 11 13 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=6.03 $Y=1.515
+ $X2=6.03 $Y2=0.495
r215 7 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.6 $Y=1.845
+ $X2=5.6 $Y2=1.68
r216 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.6 $Y=1.845 $X2=5.6
+ $Y2=2.525
r217 2 55 600 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=1 $X=4.695
+ $Y=2.415 $X2=4.835 $Y2=2.86
r218 1 52 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.495 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_1263_31# 1 2 7 9 10 12 13 14 18 19 24 27
+ 31 34 41 44
c78 14 0 1.41102e-19 $X=6.465 $Y=2.13
c79 10 0 6.84876e-20 $X=6.39 $Y=2.205
r80 34 36 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=7.185 $Y=0.825
+ $X2=7.185 $Y2=0.955
r81 29 31 36.5775 $w=2.28e-07 $l=7.3e-07 $layer=LI1_cond $X=7.345 $Y=1.775
+ $X2=7.345 $Y2=2.505
r82 27 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.785 $Y=1.68
+ $X2=6.785 $Y2=1.845
r83 27 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.785 $Y=1.68
+ $X2=6.785 $Y2=1.515
r84 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.785
+ $Y=1.68 $X2=6.785 $Y2=1.68
r85 24 29 6.94918 $w=1.8e-07 $l=1.53542e-07 $layer=LI1_cond $X=7.23 $Y=1.685
+ $X2=7.345 $Y2=1.775
r86 24 26 27.4192 $w=1.78e-07 $l=4.45e-07 $layer=LI1_cond $X=7.23 $Y=1.685
+ $X2=6.785 $Y2=1.685
r87 22 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.635 $Y=0.98
+ $X2=6.725 $Y2=0.98
r88 22 38 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=6.635 $Y=0.98
+ $X2=6.39 $Y2=0.98
r89 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.635
+ $Y=0.98 $X2=6.635 $Y2=0.98
r90 19 36 1.19992 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=7.055 $Y=0.955
+ $X2=7.185 $Y2=0.955
r91 19 21 20.1678 $w=2.38e-07 $l=4.2e-07 $layer=LI1_cond $X=7.055 $Y=0.955
+ $X2=6.635 $Y2=0.955
r92 18 45 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.725 $Y=2.055
+ $X2=6.725 $Y2=1.845
r93 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.725 $Y=1.145
+ $X2=6.725 $Y2=0.98
r94 15 44 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.725 $Y=1.145
+ $X2=6.725 $Y2=1.515
r95 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.65 $Y=2.13
+ $X2=6.725 $Y2=2.055
r96 13 14 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=6.65 $Y=2.13
+ $X2=6.465 $Y2=2.13
r97 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.39 $Y=2.205
+ $X2=6.465 $Y2=2.13
r98 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.39 $Y=2.205
+ $X2=6.39 $Y2=2.525
r99 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.39 $Y=0.815
+ $X2=6.39 $Y2=0.98
r100 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.39 $Y=0.815
+ $X2=6.39 $Y2=0.495
r101 2 31 600 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=7.225
+ $Y=2.315 $X2=7.365 $Y2=2.505
r102 1 34 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=7.095
+ $Y=0.625 $X2=7.22 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_1135_57# 1 2 7 9 11 12 14 17 19 21 23 26
+ 30 33 36 38 43 44 45 54 56
c115 36 0 1.41102e-19 $X=5.815 $Y=2.525
c116 11 0 3.12009e-19 $X=7.235 $Y=2.055
r117 49 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.53 $Y=1.54
+ $X2=8.53 $Y2=1.705
r118 49 56 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.53 $Y=1.54 $X2=8.53
+ $Y2=1.45
r119 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.53
+ $Y=1.54 $X2=8.53 $Y2=1.54
r120 45 48 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=8.53 $Y=1.335
+ $X2=8.53 $Y2=1.54
r121 42 54 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=7.325 $Y=1.33
+ $X2=7.435 $Y2=1.33
r122 42 51 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.325 $Y=1.33
+ $X2=7.235 $Y2=1.33
r123 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.325
+ $Y=1.33 $X2=7.325 $Y2=1.33
r124 39 44 1.34256 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=5.9 $Y=1.335 $X2=5.81
+ $Y2=1.335
r125 39 41 87.803 $w=1.78e-07 $l=1.425e-06 $layer=LI1_cond $X=5.9 $Y=1.335
+ $X2=7.325 $Y2=1.335
r126 38 45 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.365 $Y=1.335
+ $X2=8.53 $Y2=1.335
r127 38 41 64.0808 $w=1.78e-07 $l=1.04e-06 $layer=LI1_cond $X=8.365 $Y=1.335
+ $X2=7.325 $Y2=1.335
r128 34 44 5.16603 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=5.81 $Y=1.425 $X2=5.81
+ $Y2=1.335
r129 34 36 67.7778 $w=1.78e-07 $l=1.1e-06 $layer=LI1_cond $X=5.81 $Y=1.425
+ $X2=5.81 $Y2=2.525
r130 33 44 5.16603 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=5.81 $Y=1.245 $X2=5.81
+ $Y2=1.335
r131 33 43 32.0404 $w=1.78e-07 $l=5.2e-07 $layer=LI1_cond $X=5.81 $Y=1.245
+ $X2=5.81 $Y2=0.725
r132 28 43 5.68054 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=5.82 $Y=0.625
+ $X2=5.82 $Y2=0.725
r133 28 30 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=5.82 $Y=0.625
+ $X2=5.82 $Y2=0.49
r134 24 26 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=7.15 $Y=2.13
+ $X2=7.235 $Y2=2.13
r135 21 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.16 $Y=1.375
+ $X2=9.16 $Y2=0.945
r136 20 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.695 $Y=1.45
+ $X2=8.53 $Y2=1.45
r137 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.085 $Y=1.45
+ $X2=9.16 $Y2=1.375
r138 19 20 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=9.085 $Y=1.45
+ $X2=8.695 $Y2=1.45
r139 17 59 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.44 $Y=2.315
+ $X2=8.44 $Y2=1.705
r140 12 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.435 $Y=1.165
+ $X2=7.435 $Y2=1.33
r141 12 14 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=7.435 $Y=1.165
+ $X2=7.435 $Y2=0.835
r142 11 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.235 $Y=2.055
+ $X2=7.235 $Y2=2.13
r143 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.235 $Y=1.495
+ $X2=7.235 $Y2=1.33
r144 10 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.235 $Y=1.495
+ $X2=7.235 $Y2=2.055
r145 7 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.15 $Y=2.205
+ $X2=7.15 $Y2=2.13
r146 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.15 $Y=2.205
+ $X2=7.15 $Y2=2.525
r147 2 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.675
+ $Y=2.315 $X2=5.815 $Y2=2.525
r148 1 30 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.675
+ $Y=0.285 $X2=5.815 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%SET_B 3 8 11 12 16 18 20 22 23 25 26 28 29
+ 30 31 32 33 34 42 47
c101 25 0 1.65899e-19 $X=11.495 $Y=1.67
r102 42 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.035 $Y=0.35
+ $X2=8.035 $Y2=0.515
r103 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.035
+ $Y=0.35 $X2=8.035 $Y2=0.35
r104 33 34 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=9.84 $Y=0.452
+ $X2=10.32 $Y2=0.452
r105 32 33 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=0.452
+ $X2=9.84 $Y2=0.452
r106 31 32 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=0.452
+ $X2=9.36 $Y2=0.452
r107 30 31 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=0.452
+ $X2=8.88 $Y2=0.452
r108 30 43 11.2171 $w=3.73e-07 $l=3.65e-07 $layer=LI1_cond $X=8.4 $Y=0.452
+ $X2=8.035 $Y2=0.452
r109 29 43 3.53416 $w=3.73e-07 $l=1.15e-07 $layer=LI1_cond $X=7.92 $Y=0.452
+ $X2=8.035 $Y2=0.452
r110 28 34 3.99514 $w=3.73e-07 $l=1.3e-07 $layer=LI1_cond $X=10.45 $Y=0.452
+ $X2=10.32 $Y2=0.452
r111 26 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.495 $Y=1.67
+ $X2=11.495 $Y2=1.835
r112 26 47 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.495 $Y=1.67
+ $X2=11.495 $Y2=1.505
r113 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.495
+ $Y=1.67 $X2=11.495 $Y2=1.67
r114 23 25 53.9141 $w=1.78e-07 $l=8.75e-07 $layer=LI1_cond $X=10.62 $Y=1.675
+ $X2=11.495 $Y2=1.675
r115 22 23 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=10.535 $Y=1.585
+ $X2=10.62 $Y2=1.675
r116 21 28 8.1532 $w=3.75e-07 $l=2.26548e-07 $layer=LI1_cond $X=10.535 $Y=0.64
+ $X2=10.45 $Y2=0.452
r117 21 22 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=10.535 $Y=0.64
+ $X2=10.535 $Y2=1.585
r118 18 19 82.6961 $w=2.04e-07 $l=3.5e-07 $layer=POLY_cond $X=7.595 $Y=1.735
+ $X2=7.945 $Y2=1.735
r119 16 48 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.44 $Y=2.625
+ $X2=11.44 $Y2=1.835
r120 12 20 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.42 $Y=1.245
+ $X2=11.42 $Y2=1.155
r121 12 47 101.065 $w=1.8e-07 $l=2.6e-07 $layer=POLY_cond $X=11.42 $Y=1.245
+ $X2=11.42 $Y2=1.505
r122 11 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.405 $Y=0.835
+ $X2=11.405 $Y2=1.155
r123 8 45 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.945 $Y=0.835
+ $X2=7.945 $Y2=0.515
r124 6 19 10.0333 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.945 $Y=1.555
+ $X2=7.945 $Y2=1.735
r125 6 8 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=7.945 $Y=1.555
+ $X2=7.945 $Y2=0.835
r126 1 18 10.0333 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=7.595 $Y=1.885
+ $X2=7.595 $Y2=1.735
r127 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.595 $Y=1.885
+ $X2=7.595 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_702_47# 1 2 7 9 11 14 16 18 21 22 23 26
+ 30 32 34 36 37 38 41 43 44 47 50 52 53 56 59 60 63 70
c180 59 0 3.05811e-20 $X=4.67 $Y=2.09
c181 34 0 1.0162e-19 $X=10.03 $Y=1.785
c182 14 0 1.88568e-19 $X=4.62 $Y=2.735
r183 69 70 7.82892 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.86 $Y=2.155
+ $X2=4.025 $Y2=2.155
r184 66 69 5.94228 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=2.155
+ $X2=3.86 $Y2=2.155
r185 63 65 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=0.445
+ $X2=3.625 $Y2=0.61
r186 59 70 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=4.67 $Y=2.09
+ $X2=4.025 $Y2=2.09
r187 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.67
+ $Y=2.09 $X2=4.67 $Y2=2.09
r188 56 66 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.695 $Y=1.995
+ $X2=3.695 $Y2=2.155
r189 56 65 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=3.695 $Y=1.995
+ $X2=3.695 $Y2=0.61
r190 51 60 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.67 $Y=2.105
+ $X2=4.67 $Y2=2.09
r191 51 52 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.67 $Y=2.105
+ $X2=4.67 $Y2=2.18
r192 49 60 142.512 $w=3.3e-07 $l=8.15e-07 $layer=POLY_cond $X=4.67 $Y=1.275
+ $X2=4.67 $Y2=2.09
r193 49 50 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.67 $Y=1.275
+ $X2=4.67 $Y2=1.2
r194 45 47 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=4.28 $Y=0.84 $X2=4.58
+ $Y2=0.84
r195 43 54 50.2292 $w=1.59e-07 $l=1.68953e-07 $layer=POLY_cond $X=10.52 $Y=1.875
+ $X2=10.512 $Y2=1.71
r196 43 44 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=10.52 $Y=1.875
+ $X2=10.52 $Y2=3.075
r197 39 54 22.9461 $w=1.59e-07 $l=7.84219e-08 $layer=POLY_cond $X=10.505
+ $Y=1.635 $X2=10.512 $Y2=1.71
r198 39 41 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=10.505 $Y=1.635
+ $X2=10.505 $Y2=0.835
r199 37 54 4.22461 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=10.43 $Y=1.71
+ $X2=10.512 $Y2=1.71
r200 37 38 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=10.43 $Y=1.71
+ $X2=10.105 $Y2=1.71
r201 34 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.03 $Y=1.785
+ $X2=10.105 $Y2=1.71
r202 34 36 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.03 $Y=1.785
+ $X2=10.03 $Y2=2.315
r203 33 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.105 $Y=3.15
+ $X2=6.03 $Y2=3.15
r204 32 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.445 $Y=3.15
+ $X2=10.52 $Y2=3.075
r205 32 33 2225.4 $w=1.5e-07 $l=4.34e-06 $layer=POLY_cond $X=10.445 $Y=3.15
+ $X2=6.105 $Y2=3.15
r206 28 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.03 $Y=3.075
+ $X2=6.03 $Y2=3.15
r207 28 30 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.03 $Y=3.075
+ $X2=6.03 $Y2=2.525
r208 24 26 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=5.6 $Y=1.125
+ $X2=5.6 $Y2=0.495
r209 22 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.955 $Y=3.15
+ $X2=6.03 $Y2=3.15
r210 22 23 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.955 $Y=3.15
+ $X2=5.185 $Y2=3.15
r211 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.11 $Y=3.075
+ $X2=5.185 $Y2=3.15
r212 20 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.11 $Y=2.255
+ $X2=5.11 $Y2=3.075
r213 19 52 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=2.18
+ $X2=4.67 $Y2=2.18
r214 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.035 $Y=2.18
+ $X2=5.11 $Y2=2.255
r215 18 19 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.035 $Y=2.18
+ $X2=4.835 $Y2=2.18
r216 17 50 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.2
+ $X2=4.67 $Y2=1.2
r217 16 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.525 $Y=1.2
+ $X2=5.6 $Y2=1.125
r218 16 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.525 $Y=1.2
+ $X2=4.835 $Y2=1.2
r219 12 52 13.5877 $w=2.4e-07 $l=9.68246e-08 $layer=POLY_cond $X=4.62 $Y=2.255
+ $X2=4.67 $Y2=2.18
r220 12 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.62 $Y=2.255
+ $X2=4.62 $Y2=2.735
r221 11 50 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.58 $Y=1.125
+ $X2=4.67 $Y2=1.2
r222 10 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.58 $Y=0.915
+ $X2=4.58 $Y2=0.84
r223 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.58 $Y=0.915
+ $X2=4.58 $Y2=1.125
r224 7 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.28 $Y=0.765
+ $X2=4.28 $Y2=0.84
r225 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.28 $Y=0.765
+ $X2=4.28 $Y2=0.445
r226 2 69 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.715
+ $Y=2.105 $X2=3.86 $Y2=2.23
r227 1 63 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.51
+ $Y=0.235 $X2=3.635 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_2158_231# 1 2 9 13 14 17 21 23 27 29 31
c68 9 0 1.29862e-19 $X=11.01 $Y=2.625
r69 25 27 53.8545 $w=2.58e-07 $l=1.215e-06 $layer=LI1_cond $X=12.64 $Y=1.415
+ $X2=12.64 $Y2=2.63
r70 24 29 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=12.325 $Y=1.325
+ $X2=12.16 $Y2=1.325
r71 23 25 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=12.51 $Y=1.325
+ $X2=12.64 $Y2=1.415
r72 23 24 11.399 $w=1.78e-07 $l=1.85e-07 $layer=LI1_cond $X=12.51 $Y=1.325
+ $X2=12.325 $Y2=1.325
r73 19 29 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=12.16 $Y=1.235
+ $X2=12.16 $Y2=1.325
r74 19 21 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=12.16 $Y=1.235
+ $X2=12.16 $Y2=0.83
r75 17 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.955 $Y=1.32
+ $X2=10.955 $Y2=1.485
r76 17 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.955 $Y=1.32
+ $X2=10.955 $Y2=1.155
r77 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.955
+ $Y=1.32 $X2=10.955 $Y2=1.32
r78 14 29 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=11.995 $Y=1.325
+ $X2=12.16 $Y2=1.325
r79 14 16 64.0808 $w=1.78e-07 $l=1.04e-06 $layer=LI1_cond $X=11.995 $Y=1.325
+ $X2=10.955 $Y2=1.325
r80 13 31 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.045 $Y=0.835
+ $X2=11.045 $Y2=1.155
r81 9 32 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=11.01 $Y=2.625
+ $X2=11.01 $Y2=1.485
r82 2 27 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=12.465
+ $Y=2.415 $X2=12.605 $Y2=2.63
r83 1 21 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=12.02
+ $Y=0.625 $X2=12.16 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_1912_463# 1 2 3 12 16 18 22 24 26 28 30
+ 31 32 34 36 40 42 46 47 51
c110 47 0 1.65899e-19 $X=12.255 $Y=1.75
c111 34 0 1.29862e-19 $X=10.115 $Y=0.92
r112 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.255
+ $Y=1.75 $X2=12.255 $Y2=1.75
r113 44 46 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=12.215 $Y=1.935
+ $X2=12.215 $Y2=1.75
r114 43 51 4.9928 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=11.76 $Y=2.095
+ $X2=11.64 $Y2=2.095
r115 42 44 6.95106 $w=3.2e-07 $l=2.13542e-07 $layer=LI1_cond $X=12.09 $Y=2.095
+ $X2=12.215 $Y2=1.935
r116 42 43 11.8846 $w=3.18e-07 $l=3.3e-07 $layer=LI1_cond $X=12.09 $Y=2.095
+ $X2=11.76 $Y2=2.095
r117 38 51 1.48997 $w=2.4e-07 $l=1.6e-07 $layer=LI1_cond $X=11.64 $Y=2.255
+ $X2=11.64 $Y2=2.095
r118 38 40 18.0069 $w=2.38e-07 $l=3.75e-07 $layer=LI1_cond $X=11.64 $Y=2.255
+ $X2=11.64 $Y2=2.63
r119 37 50 7.86733 $w=1.8e-07 $l=3.2e-07 $layer=LI1_cond $X=10.28 $Y=2.025
+ $X2=9.96 $Y2=2.025
r120 36 51 4.9928 $w=2.5e-07 $l=1.50997e-07 $layer=LI1_cond $X=11.52 $Y=2.025
+ $X2=11.64 $Y2=2.095
r121 36 37 76.404 $w=1.78e-07 $l=1.24e-06 $layer=LI1_cond $X=11.52 $Y=2.025
+ $X2=10.28 $Y2=2.025
r122 32 50 2.21269 $w=6.4e-07 $l=9e-08 $layer=LI1_cond $X=9.96 $Y=1.935 $X2=9.96
+ $Y2=2.025
r123 32 34 18.9691 $w=6.38e-07 $l=1.015e-06 $layer=LI1_cond $X=9.96 $Y=1.935
+ $X2=9.96 $Y2=0.92
r124 29 47 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=12.277 $Y=2.068
+ $X2=12.277 $Y2=1.75
r125 29 30 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=12.277 $Y=2.068
+ $X2=12.277 $Y2=2.255
r126 27 47 3.70769 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=12.277 $Y=1.725
+ $X2=12.277 $Y2=1.75
r127 27 28 12.5355 $w=2.62e-07 $l=1.42653e-07 $layer=POLY_cond $X=12.277
+ $Y=1.725 $X2=12.167 $Y2=1.65
r128 24 31 20.4101 $w=1.5e-07 $l=7.74597e-08 $layer=POLY_cond $X=13.34 $Y=1.725
+ $X2=13.335 $Y2=1.65
r129 24 26 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=13.34 $Y=1.725
+ $X2=13.34 $Y2=2.155
r130 20 31 20.4101 $w=1.5e-07 $l=7.74597e-08 $layer=POLY_cond $X=13.33 $Y=1.575
+ $X2=13.335 $Y2=1.65
r131 20 22 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=13.33 $Y=1.575
+ $X2=13.33 $Y2=0.975
r132 19 28 13.4976 $w=1.5e-07 $l=2.98e-07 $layer=POLY_cond $X=12.465 $Y=1.65
+ $X2=12.167 $Y2=1.65
r133 18 31 5.30422 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=13.255 $Y=1.65
+ $X2=13.335 $Y2=1.65
r134 18 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=13.255 $Y=1.65
+ $X2=12.465 $Y2=1.65
r135 16 30 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=12.39 $Y=2.625
+ $X2=12.39 $Y2=2.255
r136 10 28 12.5355 $w=2.62e-07 $l=2.56776e-07 $layer=POLY_cond $X=11.945
+ $Y=1.575 $X2=12.167 $Y2=1.65
r137 10 12 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=11.945 $Y=1.575
+ $X2=11.945 $Y2=0.835
r138 3 40 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=11.515
+ $Y=2.415 $X2=11.655 $Y2=2.63
r139 2 50 600 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_PDIFF $count=1 $X=9.56
+ $Y=2.315 $X2=9.815 $Y2=2.02
r140 1 34 91 $w=1.7e-07 $l=6.50999e-07 $layer=licon1_NDIFF $count=2 $X=9.595
+ $Y=0.625 $X2=10.115 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_2598_153# 1 2 9 12 16 20 24 25 27 29
r42 25 30 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=13.822 $Y=1.46
+ $X2=13.822 $Y2=1.625
r43 25 29 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=13.822 $Y=1.46
+ $X2=13.822 $Y2=1.295
r44 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.81
+ $Y=1.46 $X2=13.81 $Y2=1.46
r45 22 27 0.911997 $w=3.3e-07 $l=1.53e-07 $layer=LI1_cond $X=13.255 $Y=1.46
+ $X2=13.102 $Y2=1.46
r46 22 24 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=13.255 $Y=1.46
+ $X2=13.81 $Y2=1.46
r47 18 27 5.7047 $w=2.92e-07 $l=1.65e-07 $layer=LI1_cond $X=13.102 $Y=1.625
+ $X2=13.102 $Y2=1.46
r48 18 20 13.4137 $w=3.03e-07 $l=3.55e-07 $layer=LI1_cond $X=13.102 $Y=1.625
+ $X2=13.102 $Y2=1.98
r49 14 27 5.7047 $w=2.92e-07 $l=1.70895e-07 $layer=LI1_cond $X=13.09 $Y=1.295
+ $X2=13.102 $Y2=1.46
r50 14 16 13.1708 $w=2.78e-07 $l=3.2e-07 $layer=LI1_cond $X=13.09 $Y=1.295
+ $X2=13.09 $Y2=0.975
r51 12 30 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=13.925 $Y=2.465
+ $X2=13.925 $Y2=1.625
r52 9 29 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=13.84 $Y=0.765
+ $X2=13.84 $Y2=1.295
r53 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=13
+ $Y=1.835 $X2=13.125 $Y2=1.98
r54 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=12.99
+ $Y=0.765 $X2=13.115 $Y2=0.975
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_27_408# 1 2 9 11 12 13
r32 13 16 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.02 $Y=2.095 $X2=2.02
+ $Y2=2.195
r33 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=2.095
+ $X2=2.02 $Y2=2.095
r34 11 12 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=1.855 $Y=2.095
+ $X2=0.39 $Y2=2.095
r35 7 12 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=0.242 $Y=2.18
+ $X2=0.39 $Y2=2.095
r36 7 9 0.195329 $w=2.93e-07 $l=5e-09 $layer=LI1_cond $X=0.242 $Y=2.18 $X2=0.242
+ $Y2=2.185
r37 2 16 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=1.88
+ $Y=2.04 $X2=2.02 $Y2=2.195
r38 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.04 $X2=0.26 $Y2=2.185
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 37 41 45 49
+ 53 57 62 63 65 66 67 69 74 82 100 104 111 112 115 118 121 124 127 130
c163 35 0 3.05811e-20 $X=4.405 $Y=2.93
r164 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r165 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r166 124 125 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r167 122 125 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r168 121 122 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r169 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r170 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r171 112 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r172 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r173 109 130 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=13.865 $Y=3.33
+ $X2=13.645 $Y2=3.33
r174 109 111 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.865 $Y=3.33
+ $X2=14.16 $Y2=3.33
r175 108 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r176 108 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.24 $Y2=3.33
r177 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r178 105 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.34 $Y=3.33
+ $X2=12.175 $Y2=3.33
r179 105 107 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=12.34 $Y=3.33
+ $X2=13.2 $Y2=3.33
r180 104 130 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=13.425 $Y=3.33
+ $X2=13.645 $Y2=3.33
r181 104 107 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=13.425 $Y=3.33
+ $X2=13.2 $Y2=3.33
r182 103 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r183 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r184 100 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.01 $Y=3.33
+ $X2=12.175 $Y2=3.33
r185 100 102 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=12.01 $Y=3.33
+ $X2=11.76 $Y2=3.33
r186 99 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r187 98 99 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r188 96 99 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=10.8 $Y2=3.33
r189 95 98 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=10.8 $Y2=3.33
r190 95 96 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r191 93 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r192 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r193 90 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r194 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r195 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r196 87 124 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.72 $Y=3.33
+ $X2=6.58 $Y2=3.33
r197 87 89 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r198 86 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r199 86 119 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r200 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r201 83 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.54 $Y2=3.33
r202 83 85 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r203 82 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.405 $Y2=3.33
r204 82 85 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r205 81 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r206 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r207 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r208 78 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r209 77 80 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r210 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 75 115 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.707 $Y2=3.33
r212 75 77 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r213 74 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=3.33
+ $X2=2.54 $Y2=3.33
r214 74 80 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.375 $Y=3.33
+ $X2=2.16 $Y2=3.33
r215 72 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r216 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r217 69 115 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.707 $Y2=3.33
r218 69 71 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r219 67 93 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.92 $Y2=3.33
r220 67 90 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.96 $Y2=3.33
r221 65 98 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=11.09 $Y=3.33
+ $X2=10.8 $Y2=3.33
r222 65 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.09 $Y=3.33
+ $X2=11.22 $Y2=3.33
r223 64 102 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=11.35 $Y=3.33
+ $X2=11.76 $Y2=3.33
r224 64 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.35 $Y=3.33
+ $X2=11.22 $Y2=3.33
r225 62 92 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=7.97 $Y=3.33 $X2=7.92
+ $Y2=3.33
r226 62 63 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.97 $Y=3.33
+ $X2=8.14 $Y2=3.33
r227 61 95 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.31 $Y=3.33 $X2=8.4
+ $Y2=3.33
r228 61 63 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.31 $Y=3.33
+ $X2=8.14 $Y2=3.33
r229 57 60 12.3102 $w=4.38e-07 $l=4.7e-07 $layer=LI1_cond $X=13.645 $Y=1.98
+ $X2=13.645 $Y2=2.45
r230 55 130 1.73497 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=13.645 $Y=3.245
+ $X2=13.645 $Y2=3.33
r231 55 60 20.8225 $w=4.38e-07 $l=7.95e-07 $layer=LI1_cond $X=13.645 $Y=3.245
+ $X2=13.645 $Y2=2.45
r232 51 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.175 $Y=3.245
+ $X2=12.175 $Y2=3.33
r233 51 53 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=12.175 $Y=3.245
+ $X2=12.175 $Y2=2.63
r234 47 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=3.245
+ $X2=11.22 $Y2=3.33
r235 47 49 27.2597 $w=2.58e-07 $l=6.15e-07 $layer=LI1_cond $X=11.22 $Y=3.245
+ $X2=11.22 $Y2=2.63
r236 43 63 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.14 $Y=3.245
+ $X2=8.14 $Y2=3.33
r237 43 45 33.7259 $w=3.38e-07 $l=9.95e-07 $layer=LI1_cond $X=8.14 $Y=3.245
+ $X2=8.14 $Y2=2.25
r238 39 124 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.58 $Y=3.245
+ $X2=6.58 $Y2=3.33
r239 39 41 29.2227 $w=2.78e-07 $l=7.1e-07 $layer=LI1_cond $X=6.58 $Y=3.245
+ $X2=6.58 $Y2=2.535
r240 38 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.57 $Y=3.33
+ $X2=4.405 $Y2=3.33
r241 37 124 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.44 $Y=3.33
+ $X2=6.58 $Y2=3.33
r242 37 38 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=6.44 $Y=3.33 $X2=4.57
+ $Y2=3.33
r243 33 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=3.245
+ $X2=4.405 $Y2=3.33
r244 33 35 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.405 $Y=3.245
+ $X2=4.405 $Y2=2.93
r245 29 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=3.245
+ $X2=2.54 $Y2=3.33
r246 29 31 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.54 $Y=3.245
+ $X2=2.54 $Y2=2.905
r247 25 115 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=3.245
+ $X2=0.707 $Y2=3.33
r248 25 27 28.5181 $w=2.93e-07 $l=7.3e-07 $layer=LI1_cond $X=0.707 $Y=3.245
+ $X2=0.707 $Y2=2.515
r249 8 60 300 $w=1.7e-07 $l=7.48098e-07 $layer=licon1_PDIFF $count=2 $X=13.415
+ $Y=1.835 $X2=13.71 $Y2=2.45
r250 8 57 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.415
+ $Y=1.835 $X2=13.555 $Y2=1.98
r251 7 53 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=12.05
+ $Y=2.415 $X2=12.175 $Y2=2.63
r252 6 49 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=11.085
+ $Y=2.415 $X2=11.225 $Y2=2.63
r253 5 45 300 $w=1.7e-07 $l=5.06458e-07 $layer=licon1_PDIFF $count=2 $X=7.67
+ $Y=2.315 $X2=8.145 $Y2=2.25
r254 4 41 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=6.465
+ $Y=2.315 $X2=6.605 $Y2=2.535
r255 3 35 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=4.265
+ $Y=2.415 $X2=4.405 $Y2=2.93
r256 2 31 600 $w=1.7e-07 $l=5.59017e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=2.405 $X2=2.54 $Y2=2.905
r257 1 27 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.04 $X2=0.69 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_196_128# 1 2 3 4 15 17 18 19 22 23 26 27
+ 28 30 31 32 33 36 38 42 43 50 52
c148 31 0 1.88568e-19 $X=4.4 $Y=2.58
r149 52 54 9.65982 $w=3.41e-07 $l=2.7e-07 $layer=LI1_cond $X=5.115 $Y=2.492
+ $X2=5.385 $Y2=2.492
r150 48 50 4.43636 $w=1.98e-07 $l=8e-08 $layer=LI1_cond $X=5.035 $Y=0.705
+ $X2=5.115 $Y2=0.705
r151 43 45 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.485 $Y=2.44
+ $X2=4.485 $Y2=2.58
r152 38 40 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.535 $Y=2.47
+ $X2=1.535 $Y2=2.545
r153 36 52 4.81864 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=5.115 $Y=2.295
+ $X2=5.115 $Y2=2.492
r154 35 50 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.115 $Y=0.805
+ $X2=5.115 $Y2=0.705
r155 35 36 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=5.115 $Y=0.805
+ $X2=5.115 $Y2=2.295
r156 34 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=2.44
+ $X2=4.485 $Y2=2.44
r157 33 52 6.10782 $w=3.41e-07 $l=1.07912e-07 $layer=LI1_cond $X=5.03 $Y=2.44
+ $X2=5.115 $Y2=2.492
r158 33 34 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.03 $Y=2.44
+ $X2=4.57 $Y2=2.44
r159 31 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.4 $Y=2.58
+ $X2=4.485 $Y2=2.58
r160 31 32 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.4 $Y=2.58
+ $X2=4.06 $Y2=2.58
r161 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.975 $Y=2.665
+ $X2=4.06 $Y2=2.58
r162 29 30 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.975 $Y=2.665
+ $X2=3.975 $Y2=2.895
r163 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.89 $Y=2.98
+ $X2=3.975 $Y2=2.895
r164 27 28 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=3.89 $Y=2.98
+ $X2=3.055 $Y2=2.98
r165 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.97 $Y=2.895
+ $X2=3.055 $Y2=2.98
r166 25 26 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.97 $Y=2.64
+ $X2=2.97 $Y2=2.895
r167 24 42 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=2.545
+ $X2=2.51 $Y2=2.545
r168 23 25 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.885 $Y=2.545
+ $X2=2.97 $Y2=2.64
r169 23 24 16.9282 $w=1.88e-07 $l=2.9e-07 $layer=LI1_cond $X=2.885 $Y=2.545
+ $X2=2.595 $Y2=2.545
r170 22 42 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.51 $Y=2.45
+ $X2=2.51 $Y2=2.545
r171 21 22 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=2.51 $Y=1.36
+ $X2=2.51 $Y2=2.45
r172 20 40 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=2.545
+ $X2=1.535 $Y2=2.545
r173 19 42 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=2.545
+ $X2=2.51 $Y2=2.545
r174 19 20 42.3206 $w=1.88e-07 $l=7.25e-07 $layer=LI1_cond $X=2.425 $Y=2.545
+ $X2=1.7 $Y2=2.545
r175 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.425 $Y=1.275
+ $X2=2.51 $Y2=1.36
r176 17 18 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2.425 $Y=1.275
+ $X2=1.285 $Y2=1.275
r177 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.12 $Y=1.19
+ $X2=1.285 $Y2=1.275
r178 13 15 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.12 $Y=1.19
+ $X2=1.12 $Y2=0.85
r179 4 54 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=5.26
+ $Y=2.315 $X2=5.385 $Y2=2.525
r180 3 38 600 $w=1.7e-07 $l=5.18411e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.04 $X2=1.535 $Y2=2.47
r181 2 48 182 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.285 $X2=5.035 $Y2=0.7
r182 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.64 $X2=1.12 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_1703_379# 1 2 10 15 16
r33 15 16 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=10.245 $Y=2.455
+ $X2=10.08 $Y2=2.455
r34 10 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=8.655 $Y=2.25
+ $X2=8.655 $Y2=2.37
r35 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.82 $Y=2.37
+ $X2=8.655 $Y2=2.37
r36 8 16 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=8.82 $Y=2.37
+ $X2=10.08 $Y2=2.37
r37 2 15 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=10.105
+ $Y=1.895 $X2=10.245 $Y2=2.43
r38 1 10 300 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=2 $X=8.515
+ $Y=1.895 $X2=8.655 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%A_1810_463# 1 2 7 11 14
r24 14 16 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.175 $Y=2.71
+ $X2=9.175 $Y2=2.88
r25 9 11 6.557 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=10.775 $Y=2.795
+ $X2=10.775 $Y2=2.63
r26 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.34 $Y=2.88
+ $X2=9.175 $Y2=2.88
r27 7 9 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=10.63 $Y=2.88
+ $X2=10.775 $Y2=2.795
r28 7 8 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=10.63 $Y=2.88
+ $X2=9.34 $Y2=2.88
r29 2 11 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=10.67
+ $Y=2.415 $X2=10.795 $Y2=2.63
r30 1 14 600 $w=1.7e-07 $l=4.53211e-07 $layer=licon1_PDIFF $count=1 $X=9.05
+ $Y=2.315 $X2=9.175 $Y2=2.71
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%Q 1 2 7 8 9 10 11 12 13 25 31 41
r18 38 41 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=14.175 $Y=1.99
+ $X2=14.175 $Y2=2.015
r19 23 31 0.147749 $w=3.88e-07 $l=5e-09 $layer=LI1_cond $X=14.12 $Y=0.93
+ $X2=14.12 $Y2=0.925
r20 13 48 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=14.175 $Y=2.775
+ $X2=14.175 $Y2=2.91
r21 12 13 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=14.175 $Y=2.405
+ $X2=14.175 $Y2=2.775
r22 11 38 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=14.175 $Y=1.97
+ $X2=14.175 $Y2=1.99
r23 11 53 5.09803 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=14.175 $Y=1.97
+ $X2=14.175 $Y2=1.85
r24 11 12 14.4055 $w=2.78e-07 $l=3.5e-07 $layer=LI1_cond $X=14.175 $Y=2.055
+ $X2=14.175 $Y2=2.405
r25 11 41 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=14.175 $Y=2.055
+ $X2=14.175 $Y2=2.015
r26 10 53 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=14.19 $Y=1.665
+ $X2=14.19 $Y2=1.85
r27 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=14.19 $Y=1.295
+ $X2=14.19 $Y2=1.665
r28 9 51 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=14.19 $Y=1.295
+ $X2=14.19 $Y2=1.125
r29 8 51 6.06074 $w=3.88e-07 $l=1.55e-07 $layer=LI1_cond $X=14.12 $Y=0.97
+ $X2=14.12 $Y2=1.125
r30 8 23 1.18199 $w=3.88e-07 $l=4e-08 $layer=LI1_cond $X=14.12 $Y=0.97 $X2=14.12
+ $Y2=0.93
r31 8 31 1.18199 $w=3.88e-07 $l=4e-08 $layer=LI1_cond $X=14.12 $Y=0.885
+ $X2=14.12 $Y2=0.925
r32 7 8 9.75144 $w=3.88e-07 $l=3.3e-07 $layer=LI1_cond $X=14.12 $Y=0.555
+ $X2=14.12 $Y2=0.885
r33 7 25 1.92074 $w=3.88e-07 $l=6.5e-08 $layer=LI1_cond $X=14.12 $Y=0.555
+ $X2=14.12 $Y2=0.49
r34 2 48 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=14
+ $Y=1.835 $X2=14.14 $Y2=2.91
r35 2 41 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=14 $Y=1.835
+ $X2=14.14 $Y2=2.015
r36 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.915
+ $Y=0.345 $X2=14.055 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_1%VGND 1 2 3 4 5 6 7 22 24 28 32 36 39 40 42
+ 46 50 55 56 58 59 61 62 63 72 79 88 100 101 107 110 113
r142 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r143 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r144 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r145 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r146 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r147 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=14.16 $Y2=0
r148 98 114 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=11.76 $Y2=0
r149 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r150 95 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.825 $Y=0
+ $X2=11.66 $Y2=0
r151 95 97 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=11.825 $Y=0
+ $X2=13.2 $Y2=0
r152 94 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r153 93 94 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r154 91 94 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=11.28 $Y2=0
r155 90 93 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=11.28 $Y2=0
r156 90 91 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r157 88 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.495 $Y=0
+ $X2=11.66 $Y2=0
r158 88 93 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=11.495 $Y=0
+ $X2=11.28 $Y2=0
r159 87 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r160 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r161 84 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.77 $Y=0
+ $X2=6.605 $Y2=0
r162 84 86 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.77 $Y=0 $X2=7.44
+ $Y2=0
r163 83 111 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r164 83 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r165 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r166 80 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.075
+ $Y2=0
r167 80 82 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.56
+ $Y2=0
r168 79 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.44 $Y=0
+ $X2=6.605 $Y2=0
r169 79 82 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=6.44 $Y=0 $X2=4.56
+ $Y2=0
r170 78 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r171 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r172 75 78 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r173 74 77 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r174 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r175 72 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.95 $Y=0
+ $X2=4.075 $Y2=0
r176 72 77 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.95 $Y=0 $X2=3.6
+ $Y2=0
r177 71 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r178 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r179 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r180 68 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r181 67 70 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r182 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r183 65 104 4.62984 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=0.495 $Y=0
+ $X2=0.247 $Y2=0
r184 65 67 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.495 $Y=0
+ $X2=0.72 $Y2=0
r185 63 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=7.44
+ $Y2=0
r186 63 111 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=6.48
+ $Y2=0
r187 61 97 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=13.4 $Y=0 $X2=13.2
+ $Y2=0
r188 61 62 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=13.4 $Y=0
+ $X2=13.577 $Y2=0
r189 60 100 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=13.755 $Y=0
+ $X2=14.16 $Y2=0
r190 60 62 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=13.755 $Y=0
+ $X2=13.577 $Y2=0
r191 58 86 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.485 $Y=0 $X2=7.44
+ $Y2=0
r192 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=0 $X2=7.57
+ $Y2=0
r193 57 90 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.655 $Y=0
+ $X2=7.92 $Y2=0
r194 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.655 $Y=0 $X2=7.57
+ $Y2=0
r195 55 70 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.68
+ $Y2=0
r196 55 56 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.88
+ $Y2=0
r197 54 74 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.015 $Y=0
+ $X2=2.16 $Y2=0
r198 54 56 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=1.88
+ $Y2=0
r199 50 52 17.8548 $w=3.53e-07 $l=5.5e-07 $layer=LI1_cond $X=13.577 $Y=0.49
+ $X2=13.577 $Y2=1.04
r200 48 62 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=13.577 $Y=0.085
+ $X2=13.577 $Y2=0
r201 48 50 13.1476 $w=3.53e-07 $l=4.05e-07 $layer=LI1_cond $X=13.577 $Y=0.085
+ $X2=13.577 $Y2=0.49
r202 44 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.66 $Y=0.085
+ $X2=11.66 $Y2=0
r203 44 46 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=11.66 $Y=0.085
+ $X2=11.66 $Y2=0.83
r204 40 42 60.4163 $w=1.88e-07 $l=1.035e-06 $layer=LI1_cond $X=7.655 $Y=0.915
+ $X2=8.69 $Y2=0.915
r205 39 40 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.57 $Y=0.82
+ $X2=7.655 $Y2=0.915
r206 38 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.57 $Y=0.085
+ $X2=7.57 $Y2=0
r207 38 39 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=7.57 $Y=0.085
+ $X2=7.57 $Y2=0.82
r208 34 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=0.085
+ $X2=6.605 $Y2=0
r209 34 36 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=6.605 $Y=0.085
+ $X2=6.605 $Y2=0.5
r210 30 107 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=0.085
+ $X2=4.075 $Y2=0
r211 30 32 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=4.075 $Y=0.085
+ $X2=4.075 $Y2=0.445
r212 26 56 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=0.085
+ $X2=1.88 $Y2=0
r213 26 28 32.6526 $w=2.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.88 $Y=0.085
+ $X2=1.88 $Y2=0.85
r214 22 104 3.13634 $w=3.3e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.247 $Y2=0
r215 22 24 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.33 $Y2=0.85
r216 7 52 182 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_NDIFF $count=1 $X=13.405
+ $Y=0.765 $X2=13.565 $Y2=1.04
r217 7 50 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=13.405
+ $Y=0.765 $X2=13.625 $Y2=0.49
r218 6 46 182 $w=1.7e-07 $l=2.80936e-07 $layer=licon1_NDIFF $count=1 $X=11.48
+ $Y=0.625 $X2=11.66 $Y2=0.83
r219 5 42 182 $w=1.7e-07 $l=7.9781e-07 $layer=licon1_NDIFF $count=1 $X=8.02
+ $Y=0.625 $X2=8.69 $Y2=0.905
r220 4 36 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=6.465
+ $Y=0.285 $X2=6.605 $Y2=0.5
r221 3 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.925
+ $Y=0.235 $X2=4.065 $Y2=0.445
r222 2 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.64 $X2=1.91 $Y2=0.85
r223 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.64 $X2=0.33 $Y2=0.85
.ends

