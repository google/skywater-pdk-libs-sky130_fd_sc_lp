* File: sky130_fd_sc_lp__nand4_4.pxi.spice
* Created: Fri Aug 28 10:51:03 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4_4%D N_D_M1001_g N_D_M1000_g N_D_M1011_g N_D_M1012_g
+ N_D_M1023_g N_D_M1019_g N_D_M1031_g N_D_M1027_g D D D D N_D_c_118_n
+ PM_SKY130_FD_SC_LP__NAND4_4%D
x_PM_SKY130_FD_SC_LP__NAND4_4%C N_C_M1006_g N_C_M1002_g N_C_M1009_g N_C_M1007_g
+ N_C_M1018_g N_C_M1016_g N_C_M1030_g N_C_M1028_g C C C N_C_c_197_n N_C_c_191_n
+ N_C_c_192_n PM_SKY130_FD_SC_LP__NAND4_4%C
x_PM_SKY130_FD_SC_LP__NAND4_4%B N_B_M1010_g N_B_M1015_g N_B_M1013_g N_B_M1022_g
+ N_B_M1014_g N_B_M1029_g N_B_M1020_g N_B_M1026_g B B B B N_B_c_285_n
+ N_B_c_286_n PM_SKY130_FD_SC_LP__NAND4_4%B
x_PM_SKY130_FD_SC_LP__NAND4_4%A N_A_M1004_g N_A_c_364_n N_A_M1003_g N_A_M1005_g
+ N_A_c_365_n N_A_M1008_g N_A_M1024_g N_A_c_366_n N_A_M1017_g N_A_M1025_g
+ N_A_c_367_n N_A_M1021_g A A A A N_A_c_363_n PM_SKY130_FD_SC_LP__NAND4_4%A
x_PM_SKY130_FD_SC_LP__NAND4_4%VPWR N_VPWR_M1000_s N_VPWR_M1012_s N_VPWR_M1027_s
+ N_VPWR_M1007_s N_VPWR_M1028_s N_VPWR_M1015_s N_VPWR_M1029_s N_VPWR_M1008_s
+ N_VPWR_M1021_s N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n N_VPWR_c_439_n
+ N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n
+ N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n N_VPWR_c_449_n
+ N_VPWR_c_450_n N_VPWR_c_451_n VPWR N_VPWR_c_452_n N_VPWR_c_453_n
+ N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n
+ N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_435_n
+ PM_SKY130_FD_SC_LP__NAND4_4%VPWR
x_PM_SKY130_FD_SC_LP__NAND4_4%Y N_Y_M1004_s N_Y_M1024_s N_Y_M1000_d N_Y_M1019_d
+ N_Y_M1002_d N_Y_M1016_d N_Y_M1010_d N_Y_M1022_d N_Y_M1003_d N_Y_M1017_d
+ N_Y_c_571_n N_Y_c_584_n N_Y_c_667_n N_Y_c_565_n N_Y_c_566_n N_Y_c_567_n
+ N_Y_c_613_n N_Y_c_594_n N_Y_c_671_n N_Y_c_616_n N_Y_c_675_n N_Y_c_620_n
+ N_Y_c_623_n N_Y_c_679_n N_Y_c_635_n N_Y_c_568_n N_Y_c_644_n N_Y_c_647_n
+ N_Y_c_683_n N_Y_c_572_n N_Y_c_600_n N_Y_c_624_n N_Y_c_626_n N_Y_c_569_n
+ N_Y_c_653_n Y Y Y N_Y_c_578_n N_Y_c_689_n N_Y_c_582_n
+ PM_SKY130_FD_SC_LP__NAND4_4%Y
x_PM_SKY130_FD_SC_LP__NAND4_4%A_27_65# N_A_27_65#_M1001_d N_A_27_65#_M1011_d
+ N_A_27_65#_M1031_d N_A_27_65#_M1009_d N_A_27_65#_M1030_d N_A_27_65#_c_716_n
+ N_A_27_65#_c_717_n N_A_27_65#_c_718_n N_A_27_65#_c_719_n N_A_27_65#_c_720_n
+ N_A_27_65#_c_721_n N_A_27_65#_c_722_n N_A_27_65#_c_779_p N_A_27_65#_c_723_n
+ N_A_27_65#_c_724_n N_A_27_65#_c_725_n N_A_27_65#_c_726_n
+ PM_SKY130_FD_SC_LP__NAND4_4%A_27_65#
x_PM_SKY130_FD_SC_LP__NAND4_4%VGND N_VGND_M1001_s N_VGND_M1023_s N_VGND_c_787_n
+ N_VGND_c_788_n VGND N_VGND_c_789_n N_VGND_c_790_n N_VGND_c_791_n
+ N_VGND_c_792_n N_VGND_c_793_n N_VGND_c_794_n PM_SKY130_FD_SC_LP__NAND4_4%VGND
x_PM_SKY130_FD_SC_LP__NAND4_4%A_454_65# N_A_454_65#_M1006_s N_A_454_65#_M1018_s
+ N_A_454_65#_M1013_d N_A_454_65#_M1020_d N_A_454_65#_c_872_n
+ N_A_454_65#_c_868_n N_A_454_65#_c_869_n N_A_454_65#_c_870_n
+ N_A_454_65#_c_871_n PM_SKY130_FD_SC_LP__NAND4_4%A_454_65#
x_PM_SKY130_FD_SC_LP__NAND4_4%A_843_67# N_A_843_67#_M1013_s N_A_843_67#_M1014_s
+ N_A_843_67#_M1026_s N_A_843_67#_M1005_d N_A_843_67#_M1025_d
+ N_A_843_67#_c_920_n N_A_843_67#_c_943_n N_A_843_67#_c_921_n
+ N_A_843_67#_c_948_n N_A_843_67#_c_922_n N_A_843_67#_c_923_n
+ N_A_843_67#_c_924_n N_A_843_67#_c_925_n PM_SKY130_FD_SC_LP__NAND4_4%A_843_67#
cc_1 VNB N_D_M1001_g 0.0259905f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.745
cc_2 VNB N_D_M1011_g 0.0190925f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.745
cc_3 VNB N_D_M1023_g 0.0190925f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.745
cc_4 VNB N_D_M1031_g 0.0193981f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.745
cc_5 VNB D 0.0146613f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_D_c_118_n 0.0733946f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.51
cc_7 VNB N_C_M1006_g 0.020025f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.745
cc_8 VNB N_C_M1009_g 0.0195018f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.745
cc_9 VNB N_C_M1018_g 0.0194987f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.745
cc_10 VNB N_C_M1030_g 0.0229058f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.745
cc_11 VNB N_C_c_191_n 0.0759819f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=1.51
cc_12 VNB N_C_c_192_n 0.00268666f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=1.51
cc_13 VNB N_B_M1013_g 0.025037f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.745
cc_14 VNB N_B_M1014_g 0.0187462f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.745
cc_15 VNB N_B_M1020_g 0.0187462f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.745
cc_16 VNB N_B_M1026_g 0.0189781f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=2.465
cc_17 VNB N_B_c_285_n 0.0030655f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.587
cc_18 VNB N_B_c_286_n 0.09708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_M1004_g 0.0189739f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.745
cc_20 VNB N_A_M1005_g 0.018742f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.745
cc_21 VNB N_A_M1024_g 0.018742f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.345
cc_22 VNB N_A_M1025_g 0.0262103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB A 0.01294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_c_363_n 0.084631f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.51
cc_25 VNB N_VPWR_c_435_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_565_n 0.00778591f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_27 VNB N_Y_c_566_n 0.0210665f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.51
cc_28 VNB N_Y_c_567_n 0.00134782f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.51
cc_29 VNB N_Y_c_568_n 0.00452057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_569_n 0.00228361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_65#_c_716_n 0.00252407f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.745
cc_32 VNB N_A_27_65#_c_717_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_65#_c_718_n 0.00575994f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=1.675
cc_34 VNB N_A_27_65#_c_719_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_65#_c_720_n 0.0071769f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.745
cc_36 VNB N_A_27_65#_c_721_n 0.00266623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_65#_c_722_n 0.00185825f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_A_27_65#_c_723_n 0.00291153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_65#_c_724_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_65#_c_725_n 0.0013899f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_41 VNB N_A_27_65#_c_726_n 0.00591076f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_42 VNB N_VGND_c_787_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.345
cc_43 VNB N_VGND_c_788_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.675
cc_44 VNB N_VGND_c_789_n 0.0167063f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.345
cc_45 VNB N_VGND_c_790_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=2.465
cc_46 VNB N_VGND_c_791_n 0.152856f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=1.675
cc_47 VNB N_VGND_c_792_n 0.436386f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=2.465
cc_48 VNB N_VGND_c_793_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_49 VNB N_VGND_c_794_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_50 VNB N_A_454_65#_c_868_n 0.00226807f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.345
cc_51 VNB N_A_454_65#_c_869_n 0.00231169f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.745
cc_52 VNB N_A_454_65#_c_870_n 0.00792639f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=2.465
cc_53 VNB N_A_454_65#_c_871_n 0.00231361f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.745
cc_54 VNB N_A_843_67#_c_920_n 0.0122056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_843_67#_c_921_n 0.00271277f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.745
cc_56 VNB N_A_843_67#_c_922_n 0.0119556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_843_67#_c_923_n 0.0298516f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_58 VNB N_A_843_67#_c_924_n 0.00141599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_843_67#_c_925_n 0.00141599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VPB N_D_M1000_g 0.0244533f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_61 VPB N_D_M1012_g 0.0179387f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_62 VPB N_D_M1019_g 0.0179387f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=2.465
cc_63 VPB N_D_M1027_g 0.0203096f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=2.465
cc_64 VPB D 0.0171568f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_65 VPB N_D_c_118_n 0.0140686f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.51
cc_66 VPB N_C_M1002_g 0.0198977f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_67 VPB N_C_M1007_g 0.0179387f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_68 VPB N_C_M1016_g 0.0179264f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=2.465
cc_69 VPB N_C_M1028_g 0.0178593f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=2.465
cc_70 VPB N_C_c_197_n 0.00669616f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.51
cc_71 VPB N_C_c_191_n 0.0189911f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=1.51
cc_72 VPB N_C_c_192_n 0.0030799f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=1.51
cc_73 VPB N_B_M1010_g 0.0180832f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.745
cc_74 VPB N_B_M1015_g 0.0179379f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_75 VPB N_B_M1022_g 0.0179387f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_76 VPB N_B_M1029_g 0.0235869f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=2.465
cc_77 VPB N_B_c_285_n 0.0145041f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.587
cc_78 VPB N_B_c_286_n 0.0301395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_c_364_n 0.0206946f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.675
cc_80 VPB N_A_c_365_n 0.015814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_c_366_n 0.015814f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.745
cc_82 VPB N_A_c_367_n 0.0206946f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.745
cc_83 VPB A 0.018096f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_c_363_n 0.0305773f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.51
cc_85 VPB N_VPWR_c_436_n 0.0124746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_437_n 0.049796f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=2.465
cc_87 VPB N_VPWR_c_438_n 3.28559e-19 $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_88 VPB N_VPWR_c_439_n 0.00437923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_440_n 3.22457e-19 $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.51
cc_90 VPB N_VPWR_c_441_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.245 $Y2=1.51
cc_91 VPB N_VPWR_c_442_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.585 $Y2=1.51
cc_92 VPB N_VPWR_c_443_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=1.51
cc_93 VPB N_VPWR_c_444_n 0.00234818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_445_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.587
cc_95 VPB N_VPWR_c_446_n 0.0135296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_447_n 0.0483636f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=1.587
cc_97 VPB N_VPWR_c_448_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_449_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_450_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_451_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_452_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_453_n 0.0157463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_454_n 0.0156522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_455_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_456_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_457_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_458_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_459_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_460_n 0.0125509f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_461_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_435_n 0.0503333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_Y_c_565_n 0.00146017f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.51
cc_113 N_D_M1031_g N_C_M1006_g 0.0202264f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_114 N_D_M1027_g N_C_M1002_g 0.0341156f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_115 D N_C_c_191_n 2.56089e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_116 N_D_c_118_n N_C_c_191_n 0.0203265f $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_117 D N_C_c_192_n 0.0183154f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_118 N_D_c_118_n N_C_c_192_n 0.00320472f $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_119 N_D_M1000_g N_VPWR_c_437_n 0.00509958f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_120 D N_VPWR_c_437_n 0.0233766f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_121 N_D_M1000_g N_VPWR_c_438_n 6.86223e-19 $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_122 N_D_M1012_g N_VPWR_c_438_n 0.0143756f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_123 N_D_M1019_g N_VPWR_c_438_n 0.0144748f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_124 N_D_M1027_g N_VPWR_c_438_n 7.19937e-19 $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_125 N_D_M1027_g N_VPWR_c_439_n 0.00686811f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_126 N_D_M1000_g N_VPWR_c_452_n 0.00585385f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_127 N_D_M1012_g N_VPWR_c_452_n 0.00486043f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_128 N_D_M1019_g N_VPWR_c_453_n 0.00486043f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_129 N_D_M1027_g N_VPWR_c_453_n 0.0054895f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_130 N_D_M1000_g N_VPWR_c_435_n 0.011499f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_131 N_D_M1012_g N_VPWR_c_435_n 0.00824727f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_132 N_D_M1019_g N_VPWR_c_435_n 0.00824727f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_133 N_D_M1027_g N_VPWR_c_435_n 0.0102908f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_134 N_D_M1027_g N_Y_c_571_n 9.39085e-19 $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_135 N_D_M1027_g N_Y_c_572_n 0.0135461f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_136 D Y 0.0168356f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_137 N_D_c_118_n Y 6.49221e-19 $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_138 N_D_M1027_g Y 0.00140328f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_139 D Y 0.019204f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_140 N_D_c_118_n Y 6.49221e-19 $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_141 N_D_M1012_g N_Y_c_578_n 0.0131606f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_142 N_D_M1019_g N_Y_c_578_n 0.0131057f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_143 D N_Y_c_578_n 0.043132f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_144 N_D_c_118_n N_Y_c_578_n 5.81779e-19 $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_145 N_D_M1027_g N_Y_c_582_n 0.0120398f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_146 N_D_M1001_g N_A_27_65#_c_716_n 0.00354208f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_147 N_D_M1001_g N_A_27_65#_c_717_n 0.0139726f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_148 N_D_M1011_g N_A_27_65#_c_717_n 0.013286f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_149 D N_A_27_65#_c_717_n 0.049286f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_150 N_D_c_118_n N_A_27_65#_c_717_n 0.00267963f $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_151 D N_A_27_65#_c_718_n 0.017673f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_152 N_D_M1011_g N_A_27_65#_c_719_n 8.28776e-19 $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_153 N_D_M1023_g N_A_27_65#_c_719_n 8.28776e-19 $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_154 N_D_M1023_g N_A_27_65#_c_720_n 0.013286f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_155 N_D_M1031_g N_A_27_65#_c_720_n 0.0142283f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_156 D N_A_27_65#_c_720_n 0.0404108f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_157 N_D_c_118_n N_A_27_65#_c_720_n 0.00406698f $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_158 N_D_M1031_g N_A_27_65#_c_722_n 4.90985e-19 $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_159 D N_A_27_65#_c_724_n 0.0160075f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_160 N_D_c_118_n N_A_27_65#_c_724_n 0.00278273f $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_161 N_D_M1001_g N_VGND_c_787_n 0.012533f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_162 N_D_M1011_g N_VGND_c_787_n 0.0102222f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_163 N_D_M1023_g N_VGND_c_787_n 5.123e-19 $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_164 N_D_M1011_g N_VGND_c_788_n 5.123e-19 $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_165 N_D_M1023_g N_VGND_c_788_n 0.0102222f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_166 N_D_M1031_g N_VGND_c_788_n 0.0103482f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_167 N_D_M1001_g N_VGND_c_789_n 0.00414769f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_168 N_D_M1011_g N_VGND_c_790_n 0.00414769f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_169 N_D_M1023_g N_VGND_c_790_n 0.00414769f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_170 N_D_M1031_g N_VGND_c_791_n 0.00414769f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_171 N_D_M1001_g N_VGND_c_792_n 0.00823375f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_172 N_D_M1011_g N_VGND_c_792_n 0.00787505f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_173 N_D_M1023_g N_VGND_c_792_n 0.00787505f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_174 N_D_M1031_g N_VGND_c_792_n 0.0078848f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_175 N_C_M1028_g N_B_M1010_g 0.0359893f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_176 N_C_M1028_g N_B_c_285_n 2.80931e-19 $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_177 N_C_c_191_n N_B_c_286_n 0.0143f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_178 N_C_M1002_g N_VPWR_c_439_n 0.00686811f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_179 N_C_M1002_g N_VPWR_c_440_n 7.32965e-19 $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_180 N_C_M1007_g N_VPWR_c_440_n 0.0151391f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_181 N_C_M1016_g N_VPWR_c_440_n 0.0149593f $X=3.265 $Y=2.465 $X2=0 $Y2=0
cc_182 N_C_M1028_g N_VPWR_c_440_n 6.80491e-19 $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_183 N_C_M1016_g N_VPWR_c_441_n 6.80491e-19 $X=3.265 $Y=2.465 $X2=0 $Y2=0
cc_184 N_C_M1028_g N_VPWR_c_441_n 0.0148681f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_185 N_C_M1016_g N_VPWR_c_448_n 0.00486043f $X=3.265 $Y=2.465 $X2=0 $Y2=0
cc_186 N_C_M1028_g N_VPWR_c_448_n 0.00486043f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_187 N_C_M1002_g N_VPWR_c_454_n 0.00533769f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_188 N_C_M1007_g N_VPWR_c_454_n 0.00486043f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_189 N_C_M1002_g N_VPWR_c_435_n 0.00992019f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_190 N_C_M1007_g N_VPWR_c_435_n 0.00824727f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_191 N_C_M1016_g N_VPWR_c_435_n 0.00824727f $X=3.265 $Y=2.465 $X2=0 $Y2=0
cc_192 N_C_M1028_g N_VPWR_c_435_n 0.00824727f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_193 N_C_M1002_g N_Y_c_571_n 0.013227f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_194 N_C_M1007_g N_Y_c_584_n 0.0122595f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_195 N_C_M1016_g N_Y_c_584_n 0.0122595f $X=3.265 $Y=2.465 $X2=0 $Y2=0
cc_196 N_C_c_197_n N_Y_c_584_n 0.0479354f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_197 N_C_c_191_n N_Y_c_584_n 5.70783e-19 $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_198 N_C_M1016_g N_Y_c_565_n 0.00105613f $X=3.265 $Y=2.465 $X2=0 $Y2=0
cc_199 N_C_M1030_g N_Y_c_565_n 0.00598723f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_200 N_C_M1028_g N_Y_c_565_n 0.00713623f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_201 N_C_c_197_n N_Y_c_565_n 0.0276152f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_202 N_C_c_191_n N_Y_c_565_n 0.00743849f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_203 N_C_M1030_g N_Y_c_567_n 0.00506442f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_204 N_C_M1028_g N_Y_c_594_n 0.0110208f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_205 N_C_c_191_n N_Y_c_594_n 0.00317776f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_206 N_C_M1002_g N_Y_c_572_n 0.0111388f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_207 N_C_c_197_n N_Y_c_572_n 0.00425245f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_208 N_C_c_191_n N_Y_c_572_n 0.00120453f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_209 N_C_c_192_n N_Y_c_572_n 0.0219604f $X=2.385 $Y=1.565 $X2=0 $Y2=0
cc_210 N_C_M1002_g N_Y_c_600_n 0.00103713f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_211 N_C_c_197_n N_Y_c_600_n 0.0202219f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_212 N_C_c_191_n N_Y_c_600_n 6.4545e-19 $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_213 N_C_M1002_g N_Y_c_582_n 7.95991e-19 $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_214 N_C_M1006_g N_A_27_65#_c_720_n 0.00192697f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_215 N_C_M1006_g N_A_27_65#_c_721_n 0.0117888f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_216 N_C_M1009_g N_A_27_65#_c_721_n 0.0111044f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_217 N_C_M1018_g N_A_27_65#_c_723_n 0.0111044f $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_218 N_C_M1030_g N_A_27_65#_c_723_n 0.0106489f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_219 N_C_M1030_g N_A_27_65#_c_726_n 0.00150276f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_220 N_C_M1006_g N_VGND_c_788_n 5.59621e-19 $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_221 N_C_M1006_g N_VGND_c_791_n 0.0030414f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_222 N_C_M1009_g N_VGND_c_791_n 0.0030414f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_223 N_C_M1018_g N_VGND_c_791_n 0.0030414f $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_224 N_C_M1030_g N_VGND_c_791_n 0.0030414f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_225 N_C_M1006_g N_VGND_c_792_n 0.00435814f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_226 N_C_M1009_g N_VGND_c_792_n 0.0043484f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_227 N_C_M1018_g N_VGND_c_792_n 0.0043484f $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_228 N_C_M1030_g N_VGND_c_792_n 0.00483918f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_229 N_C_M1006_g N_A_454_65#_c_872_n 0.00466181f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_230 N_C_M1009_g N_A_454_65#_c_872_n 0.00590281f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_231 N_C_M1018_g N_A_454_65#_c_872_n 5.08406e-19 $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_232 N_C_M1009_g N_A_454_65#_c_868_n 0.00907529f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_233 N_C_M1018_g N_A_454_65#_c_868_n 0.0101078f $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_234 N_C_c_197_n N_A_454_65#_c_868_n 0.0383442f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_235 N_C_c_191_n N_A_454_65#_c_868_n 0.00273579f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_236 N_C_M1006_g N_A_454_65#_c_869_n 0.00253474f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_237 N_C_M1009_g N_A_454_65#_c_869_n 0.00120503f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_238 N_C_c_197_n N_A_454_65#_c_869_n 0.0154921f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_239 N_C_c_191_n N_A_454_65#_c_869_n 0.00281768f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_240 N_C_c_192_n N_A_454_65#_c_869_n 0.0114687f $X=2.385 $Y=1.565 $X2=0 $Y2=0
cc_241 N_C_M1030_g N_A_454_65#_c_870_n 0.014566f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_242 N_C_c_197_n N_A_454_65#_c_870_n 4.77713e-19 $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_243 N_C_c_191_n N_A_454_65#_c_870_n 0.00162676f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_244 N_C_M1009_g N_A_454_65#_c_871_n 5.90645e-19 $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_245 N_C_M1018_g N_A_454_65#_c_871_n 0.00761643f $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_246 N_C_M1030_g N_A_454_65#_c_871_n 0.0169044f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_247 N_C_c_197_n N_A_454_65#_c_871_n 0.0267867f $X=3.285 $Y=1.51 $X2=0 $Y2=0
cc_248 N_C_c_191_n N_A_454_65#_c_871_n 0.00281811f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_249 N_C_M1030_g N_A_843_67#_c_920_n 4.77499e-19 $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_250 N_B_M1026_g N_A_M1004_g 0.0341662f $X=5.865 $Y=0.755 $X2=0 $Y2=0
cc_251 N_B_c_285_n A 0.023354f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_252 N_B_c_286_n A 3.08904e-19 $X=5.865 $Y=1.51 $X2=0 $Y2=0
cc_253 N_B_c_285_n N_A_c_363_n 8.72863e-19 $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_254 N_B_c_286_n N_A_c_363_n 0.0230593f $X=5.865 $Y=1.51 $X2=0 $Y2=0
cc_255 N_B_M1010_g N_VPWR_c_441_n 0.0148681f $X=4.125 $Y=2.465 $X2=0 $Y2=0
cc_256 N_B_M1015_g N_VPWR_c_441_n 6.80491e-19 $X=4.555 $Y=2.465 $X2=0 $Y2=0
cc_257 N_B_M1010_g N_VPWR_c_442_n 6.80491e-19 $X=4.125 $Y=2.465 $X2=0 $Y2=0
cc_258 N_B_M1015_g N_VPWR_c_442_n 0.0149593f $X=4.555 $Y=2.465 $X2=0 $Y2=0
cc_259 N_B_M1022_g N_VPWR_c_442_n 0.0149593f $X=4.985 $Y=2.465 $X2=0 $Y2=0
cc_260 N_B_M1029_g N_VPWR_c_442_n 6.80491e-19 $X=5.415 $Y=2.465 $X2=0 $Y2=0
cc_261 N_B_M1022_g N_VPWR_c_443_n 0.00486043f $X=4.985 $Y=2.465 $X2=0 $Y2=0
cc_262 N_B_M1029_g N_VPWR_c_443_n 0.00486043f $X=5.415 $Y=2.465 $X2=0 $Y2=0
cc_263 N_B_M1022_g N_VPWR_c_444_n 6.94833e-19 $X=4.985 $Y=2.465 $X2=0 $Y2=0
cc_264 N_B_M1029_g N_VPWR_c_444_n 0.0189553f $X=5.415 $Y=2.465 $X2=0 $Y2=0
cc_265 N_B_M1010_g N_VPWR_c_450_n 0.00486043f $X=4.125 $Y=2.465 $X2=0 $Y2=0
cc_266 N_B_M1015_g N_VPWR_c_450_n 0.00486043f $X=4.555 $Y=2.465 $X2=0 $Y2=0
cc_267 N_B_M1010_g N_VPWR_c_435_n 0.00824727f $X=4.125 $Y=2.465 $X2=0 $Y2=0
cc_268 N_B_M1015_g N_VPWR_c_435_n 0.00824727f $X=4.555 $Y=2.465 $X2=0 $Y2=0
cc_269 N_B_M1022_g N_VPWR_c_435_n 0.00824727f $X=4.985 $Y=2.465 $X2=0 $Y2=0
cc_270 N_B_M1029_g N_VPWR_c_435_n 0.00824727f $X=5.415 $Y=2.465 $X2=0 $Y2=0
cc_271 N_B_M1010_g N_Y_c_565_n 0.00204091f $X=4.125 $Y=2.465 $X2=0 $Y2=0
cc_272 N_B_c_285_n N_Y_c_565_n 0.0250521f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_273 N_B_c_286_n N_Y_c_565_n 0.00272329f $X=5.865 $Y=1.51 $X2=0 $Y2=0
cc_274 N_B_M1013_g N_Y_c_566_n 0.0125331f $X=4.575 $Y=0.755 $X2=0 $Y2=0
cc_275 N_B_M1014_g N_Y_c_566_n 0.0104926f $X=5.005 $Y=0.755 $X2=0 $Y2=0
cc_276 N_B_M1020_g N_Y_c_566_n 0.0104926f $X=5.435 $Y=0.755 $X2=0 $Y2=0
cc_277 N_B_M1026_g N_Y_c_566_n 0.0118639f $X=5.865 $Y=0.755 $X2=0 $Y2=0
cc_278 N_B_c_285_n N_Y_c_566_n 0.150146f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_279 N_B_c_286_n N_Y_c_566_n 0.0236123f $X=5.865 $Y=1.51 $X2=0 $Y2=0
cc_280 N_B_M1010_g N_Y_c_613_n 0.0122129f $X=4.125 $Y=2.465 $X2=0 $Y2=0
cc_281 N_B_c_285_n N_Y_c_613_n 0.0159139f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_282 N_B_c_286_n N_Y_c_613_n 2.96829e-19 $X=5.865 $Y=1.51 $X2=0 $Y2=0
cc_283 N_B_M1015_g N_Y_c_616_n 0.0122595f $X=4.555 $Y=2.465 $X2=0 $Y2=0
cc_284 N_B_M1022_g N_Y_c_616_n 0.0122595f $X=4.985 $Y=2.465 $X2=0 $Y2=0
cc_285 N_B_c_285_n N_Y_c_616_n 0.0427276f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_286 N_B_c_286_n N_Y_c_616_n 5.768e-19 $X=5.865 $Y=1.51 $X2=0 $Y2=0
cc_287 N_B_M1029_g N_Y_c_620_n 0.0143f $X=5.415 $Y=2.465 $X2=0 $Y2=0
cc_288 N_B_c_285_n N_Y_c_620_n 0.0509486f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_289 N_B_c_286_n N_Y_c_620_n 0.00287287f $X=5.865 $Y=1.51 $X2=0 $Y2=0
cc_290 N_B_M1026_g N_Y_c_623_n 8.43475e-19 $X=5.865 $Y=0.755 $X2=0 $Y2=0
cc_291 N_B_c_285_n N_Y_c_624_n 0.0153757f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_292 N_B_c_286_n N_Y_c_624_n 6.52992e-19 $X=5.865 $Y=1.51 $X2=0 $Y2=0
cc_293 N_B_c_285_n N_Y_c_626_n 0.0153757f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_294 N_B_c_286_n N_Y_c_626_n 6.51484e-19 $X=5.865 $Y=1.51 $X2=0 $Y2=0
cc_295 N_B_M1013_g N_A_27_65#_c_726_n 9.20079e-19 $X=4.575 $Y=0.755 $X2=0 $Y2=0
cc_296 N_B_M1013_g N_VGND_c_791_n 0.00300112f $X=4.575 $Y=0.755 $X2=0 $Y2=0
cc_297 N_B_M1014_g N_VGND_c_791_n 0.00300112f $X=5.005 $Y=0.755 $X2=0 $Y2=0
cc_298 N_B_M1020_g N_VGND_c_791_n 0.00300112f $X=5.435 $Y=0.755 $X2=0 $Y2=0
cc_299 N_B_M1026_g N_VGND_c_791_n 0.00300112f $X=5.865 $Y=0.755 $X2=0 $Y2=0
cc_300 N_B_M1013_g N_VGND_c_792_n 0.00457098f $X=4.575 $Y=0.755 $X2=0 $Y2=0
cc_301 N_B_M1014_g N_VGND_c_792_n 0.00417108f $X=5.005 $Y=0.755 $X2=0 $Y2=0
cc_302 N_B_M1020_g N_VGND_c_792_n 0.00417108f $X=5.435 $Y=0.755 $X2=0 $Y2=0
cc_303 N_B_M1026_g N_VGND_c_792_n 0.00417887f $X=5.865 $Y=0.755 $X2=0 $Y2=0
cc_304 N_B_M1013_g N_A_454_65#_c_870_n 0.0104719f $X=4.575 $Y=0.755 $X2=0 $Y2=0
cc_305 N_B_M1014_g N_A_454_65#_c_870_n 0.00843134f $X=5.005 $Y=0.755 $X2=0 $Y2=0
cc_306 N_B_M1020_g N_A_454_65#_c_870_n 0.00843134f $X=5.435 $Y=0.755 $X2=0 $Y2=0
cc_307 N_B_M1026_g N_A_454_65#_c_870_n 0.00236045f $X=5.865 $Y=0.755 $X2=0 $Y2=0
cc_308 N_B_M1013_g N_A_843_67#_c_920_n 0.0120693f $X=4.575 $Y=0.755 $X2=0 $Y2=0
cc_309 N_B_M1014_g N_A_843_67#_c_920_n 0.0115903f $X=5.005 $Y=0.755 $X2=0 $Y2=0
cc_310 N_B_M1020_g N_A_843_67#_c_920_n 0.0115545f $X=5.435 $Y=0.755 $X2=0 $Y2=0
cc_311 N_B_M1026_g N_A_843_67#_c_920_n 0.0153553f $X=5.865 $Y=0.755 $X2=0 $Y2=0
cc_312 N_A_c_364_n N_VPWR_c_444_n 0.0189553f $X=6.295 $Y=1.725 $X2=0 $Y2=0
cc_313 N_A_c_365_n N_VPWR_c_444_n 6.94833e-19 $X=6.725 $Y=1.725 $X2=0 $Y2=0
cc_314 N_A_c_364_n N_VPWR_c_445_n 6.80491e-19 $X=6.295 $Y=1.725 $X2=0 $Y2=0
cc_315 N_A_c_365_n N_VPWR_c_445_n 0.0149593f $X=6.725 $Y=1.725 $X2=0 $Y2=0
cc_316 N_A_c_366_n N_VPWR_c_445_n 0.0149593f $X=7.155 $Y=1.725 $X2=0 $Y2=0
cc_317 N_A_c_367_n N_VPWR_c_445_n 6.80491e-19 $X=7.585 $Y=1.725 $X2=0 $Y2=0
cc_318 N_A_c_366_n N_VPWR_c_447_n 7.28867e-19 $X=7.155 $Y=1.725 $X2=0 $Y2=0
cc_319 N_A_c_367_n N_VPWR_c_447_n 0.0202762f $X=7.585 $Y=1.725 $X2=0 $Y2=0
cc_320 A N_VPWR_c_447_n 0.0257069f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_321 N_A_c_363_n N_VPWR_c_447_n 0.00148251f $X=7.585 $Y=1.535 $X2=0 $Y2=0
cc_322 N_A_c_364_n N_VPWR_c_455_n 0.00486043f $X=6.295 $Y=1.725 $X2=0 $Y2=0
cc_323 N_A_c_365_n N_VPWR_c_455_n 0.00486043f $X=6.725 $Y=1.725 $X2=0 $Y2=0
cc_324 N_A_c_366_n N_VPWR_c_456_n 0.00486043f $X=7.155 $Y=1.725 $X2=0 $Y2=0
cc_325 N_A_c_367_n N_VPWR_c_456_n 0.00486043f $X=7.585 $Y=1.725 $X2=0 $Y2=0
cc_326 N_A_c_364_n N_VPWR_c_435_n 0.00824727f $X=6.295 $Y=1.725 $X2=0 $Y2=0
cc_327 N_A_c_365_n N_VPWR_c_435_n 0.00824727f $X=6.725 $Y=1.725 $X2=0 $Y2=0
cc_328 N_A_c_366_n N_VPWR_c_435_n 0.00824727f $X=7.155 $Y=1.725 $X2=0 $Y2=0
cc_329 N_A_c_367_n N_VPWR_c_435_n 0.00824727f $X=7.585 $Y=1.725 $X2=0 $Y2=0
cc_330 N_A_M1004_g N_Y_c_566_n 0.00911783f $X=6.295 $Y=0.755 $X2=0 $Y2=0
cc_331 A N_Y_c_566_n 0.00888173f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_332 N_A_c_364_n N_Y_c_620_n 0.0143f $X=6.295 $Y=1.725 $X2=0 $Y2=0
cc_333 A N_Y_c_620_n 0.0125341f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_334 N_A_M1004_g N_Y_c_623_n 0.00634772f $X=6.295 $Y=0.755 $X2=0 $Y2=0
cc_335 N_A_M1005_g N_Y_c_623_n 0.00621687f $X=6.725 $Y=0.755 $X2=0 $Y2=0
cc_336 N_A_M1024_g N_Y_c_623_n 5.16893e-19 $X=7.155 $Y=0.755 $X2=0 $Y2=0
cc_337 N_A_c_365_n N_Y_c_635_n 0.0122129f $X=6.725 $Y=1.725 $X2=0 $Y2=0
cc_338 N_A_c_366_n N_Y_c_635_n 0.0122595f $X=7.155 $Y=1.725 $X2=0 $Y2=0
cc_339 A N_Y_c_635_n 0.0427275f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_340 N_A_c_363_n N_Y_c_635_n 6.55867e-19 $X=7.585 $Y=1.535 $X2=0 $Y2=0
cc_341 N_A_M1005_g N_Y_c_568_n 0.0091644f $X=6.725 $Y=0.755 $X2=0 $Y2=0
cc_342 N_A_M1024_g N_Y_c_568_n 0.0108465f $X=7.155 $Y=0.755 $X2=0 $Y2=0
cc_343 N_A_M1025_g N_Y_c_568_n 0.00529889f $X=7.585 $Y=0.755 $X2=0 $Y2=0
cc_344 A N_Y_c_568_n 0.0661906f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_345 N_A_c_363_n N_Y_c_568_n 0.00516597f $X=7.585 $Y=1.535 $X2=0 $Y2=0
cc_346 N_A_M1005_g N_Y_c_644_n 5.16893e-19 $X=6.725 $Y=0.755 $X2=0 $Y2=0
cc_347 N_A_M1024_g N_Y_c_644_n 0.00621687f $X=7.155 $Y=0.755 $X2=0 $Y2=0
cc_348 N_A_M1025_g N_Y_c_644_n 0.00522733f $X=7.585 $Y=0.755 $X2=0 $Y2=0
cc_349 A N_Y_c_647_n 0.0153756f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_350 N_A_c_363_n N_Y_c_647_n 7.38452e-19 $X=7.585 $Y=1.535 $X2=0 $Y2=0
cc_351 N_A_M1004_g N_Y_c_569_n 0.00168206f $X=6.295 $Y=0.755 $X2=0 $Y2=0
cc_352 N_A_M1005_g N_Y_c_569_n 0.00168206f $X=6.725 $Y=0.755 $X2=0 $Y2=0
cc_353 A N_Y_c_569_n 0.0274057f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_354 N_A_c_363_n N_Y_c_569_n 0.00262908f $X=7.585 $Y=1.535 $X2=0 $Y2=0
cc_355 A N_Y_c_653_n 0.0153756f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_356 N_A_c_363_n N_Y_c_653_n 7.38452e-19 $X=7.585 $Y=1.535 $X2=0 $Y2=0
cc_357 N_A_M1004_g N_VGND_c_791_n 0.00300112f $X=6.295 $Y=0.755 $X2=0 $Y2=0
cc_358 N_A_M1005_g N_VGND_c_791_n 0.00300112f $X=6.725 $Y=0.755 $X2=0 $Y2=0
cc_359 N_A_M1024_g N_VGND_c_791_n 0.00300112f $X=7.155 $Y=0.755 $X2=0 $Y2=0
cc_360 N_A_M1025_g N_VGND_c_791_n 0.00300112f $X=7.585 $Y=0.755 $X2=0 $Y2=0
cc_361 N_A_M1004_g N_VGND_c_792_n 0.00417887f $X=6.295 $Y=0.755 $X2=0 $Y2=0
cc_362 N_A_M1005_g N_VGND_c_792_n 0.00417108f $X=6.725 $Y=0.755 $X2=0 $Y2=0
cc_363 N_A_M1024_g N_VGND_c_792_n 0.00417108f $X=7.155 $Y=0.755 $X2=0 $Y2=0
cc_364 N_A_M1025_g N_VGND_c_792_n 0.0044832f $X=7.585 $Y=0.755 $X2=0 $Y2=0
cc_365 N_A_M1004_g N_A_843_67#_c_921_n 0.0112649f $X=6.295 $Y=0.755 $X2=0 $Y2=0
cc_366 N_A_M1005_g N_A_843_67#_c_921_n 0.0113115f $X=6.725 $Y=0.755 $X2=0 $Y2=0
cc_367 N_A_M1024_g N_A_843_67#_c_922_n 0.0113115f $X=7.155 $Y=0.755 $X2=0 $Y2=0
cc_368 N_A_M1025_g N_A_843_67#_c_922_n 0.012468f $X=7.585 $Y=0.755 $X2=0 $Y2=0
cc_369 N_A_M1025_g N_A_843_67#_c_923_n 0.00354524f $X=7.585 $Y=0.755 $X2=0 $Y2=0
cc_370 A N_A_843_67#_c_923_n 0.0175666f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A_c_363_n N_A_843_67#_c_923_n 0.00507493f $X=7.585 $Y=1.535 $X2=0 $Y2=0
cc_372 N_VPWR_c_435_n N_Y_M1000_d 0.0041489f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_373 N_VPWR_c_435_n N_Y_M1019_d 0.00380103f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_374 N_VPWR_c_435_n N_Y_M1002_d 0.00380103f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_375 N_VPWR_c_435_n N_Y_M1016_d 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_376 N_VPWR_c_435_n N_Y_M1010_d 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_377 N_VPWR_c_435_n N_Y_M1022_d 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_378 N_VPWR_c_435_n N_Y_M1003_d 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_379 N_VPWR_c_435_n N_Y_M1017_d 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_380 N_VPWR_c_454_n N_Y_c_571_n 0.0163698f $X=2.885 $Y=3.33 $X2=0 $Y2=0
cc_381 N_VPWR_c_435_n N_Y_c_571_n 0.0101905f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_382 N_VPWR_M1007_s N_Y_c_584_n 0.00332836f $X=2.91 $Y=1.835 $X2=0 $Y2=0
cc_383 N_VPWR_c_440_n N_Y_c_584_n 0.0170777f $X=3.05 $Y=2.36 $X2=0 $Y2=0
cc_384 N_VPWR_c_448_n N_Y_c_667_n 0.0124525f $X=3.745 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_c_435_n N_Y_c_667_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_M1028_s N_Y_c_613_n 0.00492819f $X=3.77 $Y=1.835 $X2=0 $Y2=0
cc_387 N_VPWR_c_441_n N_Y_c_594_n 0.0170777f $X=3.91 $Y=2.36 $X2=0 $Y2=0
cc_388 N_VPWR_c_450_n N_Y_c_671_n 0.0124525f $X=4.605 $Y=3.33 $X2=0 $Y2=0
cc_389 N_VPWR_c_435_n N_Y_c_671_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_390 N_VPWR_M1015_s N_Y_c_616_n 0.00332836f $X=4.63 $Y=1.835 $X2=0 $Y2=0
cc_391 N_VPWR_c_442_n N_Y_c_616_n 0.0170777f $X=4.77 $Y=2.36 $X2=0 $Y2=0
cc_392 N_VPWR_c_443_n N_Y_c_675_n 0.0124525f $X=5.465 $Y=3.33 $X2=0 $Y2=0
cc_393 N_VPWR_c_435_n N_Y_c_675_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_394 N_VPWR_M1029_s N_Y_c_620_n 0.0170244f $X=5.49 $Y=1.835 $X2=0 $Y2=0
cc_395 N_VPWR_c_444_n N_Y_c_620_n 0.053689f $X=6.08 $Y=2.36 $X2=0 $Y2=0
cc_396 N_VPWR_c_455_n N_Y_c_679_n 0.0124525f $X=6.775 $Y=3.33 $X2=0 $Y2=0
cc_397 N_VPWR_c_435_n N_Y_c_679_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_398 N_VPWR_M1008_s N_Y_c_635_n 0.00331217f $X=6.8 $Y=1.835 $X2=0 $Y2=0
cc_399 N_VPWR_c_445_n N_Y_c_635_n 0.0170777f $X=6.94 $Y=2.36 $X2=0 $Y2=0
cc_400 N_VPWR_c_456_n N_Y_c_683_n 0.0124525f $X=7.635 $Y=3.33 $X2=0 $Y2=0
cc_401 N_VPWR_c_435_n N_Y_c_683_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_402 N_VPWR_M1027_s N_Y_c_572_n 0.008649f $X=1.89 $Y=1.835 $X2=0 $Y2=0
cc_403 N_VPWR_c_439_n N_Y_c_572_n 0.0265229f $X=2.11 $Y=2.36 $X2=0 $Y2=0
cc_404 N_VPWR_M1012_s N_Y_c_578_n 0.00334509f $X=1.03 $Y=1.835 $X2=0 $Y2=0
cc_405 N_VPWR_c_438_n N_Y_c_578_n 0.0172684f $X=1.17 $Y=2.39 $X2=0 $Y2=0
cc_406 N_VPWR_c_452_n N_Y_c_689_n 0.0136943f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_407 N_VPWR_c_435_n N_Y_c_689_n 0.00866972f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_408 N_VPWR_c_453_n N_Y_c_582_n 0.015688f $X=1.945 $Y=3.33 $X2=0 $Y2=0
cc_409 N_VPWR_c_435_n N_Y_c_582_n 0.00984745f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_410 N_Y_c_566_n N_A_27_65#_M1030_d 0.00186357f $X=6.345 $Y=1.17 $X2=0 $Y2=0
cc_411 N_Y_c_567_n N_A_27_65#_M1030_d 0.00329984f $X=3.8 $Y=1.17 $X2=0 $Y2=0
cc_412 N_Y_c_572_n N_A_27_65#_c_720_n 0.00786592f $X=2.445 $Y=2.005 $X2=0 $Y2=0
cc_413 N_Y_c_566_n N_A_454_65#_M1013_d 0.00176891f $X=6.345 $Y=1.17 $X2=0 $Y2=0
cc_414 N_Y_c_566_n N_A_454_65#_M1020_d 0.00176891f $X=6.345 $Y=1.17 $X2=0 $Y2=0
cc_415 N_Y_c_566_n N_A_454_65#_c_870_n 0.115672f $X=6.345 $Y=1.17 $X2=0 $Y2=0
cc_416 N_Y_c_567_n N_A_454_65#_c_870_n 0.013831f $X=3.8 $Y=1.17 $X2=0 $Y2=0
cc_417 N_Y_c_567_n N_A_454_65#_c_871_n 0.00898376f $X=3.8 $Y=1.17 $X2=0 $Y2=0
cc_418 N_Y_c_566_n N_A_843_67#_M1013_s 0.00294684f $X=6.345 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_419 N_Y_c_566_n N_A_843_67#_M1014_s 0.00176891f $X=6.345 $Y=1.17 $X2=0 $Y2=0
cc_420 N_Y_c_566_n N_A_843_67#_M1026_s 0.00176461f $X=6.345 $Y=1.17 $X2=0 $Y2=0
cc_421 N_Y_c_568_n N_A_843_67#_M1005_d 0.00176461f $X=7.205 $Y=1.17 $X2=0 $Y2=0
cc_422 N_Y_c_566_n N_A_843_67#_c_920_n 0.00359747f $X=6.345 $Y=1.17 $X2=0 $Y2=0
cc_423 N_Y_c_566_n N_A_843_67#_c_943_n 0.0134388f $X=6.345 $Y=1.17 $X2=0 $Y2=0
cc_424 N_Y_M1004_s N_A_843_67#_c_921_n 0.00180746f $X=6.37 $Y=0.335 $X2=0 $Y2=0
cc_425 N_Y_c_566_n N_A_843_67#_c_921_n 0.00280043f $X=6.345 $Y=1.17 $X2=0 $Y2=0
cc_426 N_Y_c_623_n N_A_843_67#_c_921_n 0.0151822f $X=6.51 $Y=0.71 $X2=0 $Y2=0
cc_427 N_Y_c_568_n N_A_843_67#_c_921_n 0.00280043f $X=7.205 $Y=1.17 $X2=0 $Y2=0
cc_428 N_Y_c_568_n N_A_843_67#_c_948_n 0.0134388f $X=7.205 $Y=1.17 $X2=0 $Y2=0
cc_429 N_Y_M1024_s N_A_843_67#_c_922_n 0.00180746f $X=7.23 $Y=0.335 $X2=0 $Y2=0
cc_430 N_Y_c_568_n N_A_843_67#_c_922_n 0.00280043f $X=7.205 $Y=1.17 $X2=0 $Y2=0
cc_431 N_Y_c_644_n N_A_843_67#_c_922_n 0.0151822f $X=7.37 $Y=0.71 $X2=0 $Y2=0
cc_432 N_Y_c_568_n N_A_843_67#_c_923_n 0.00539933f $X=7.205 $Y=1.17 $X2=0 $Y2=0
cc_433 N_A_27_65#_c_717_n N_VGND_M1001_s 0.00176461f $X=1.025 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_434 N_A_27_65#_c_720_n N_VGND_M1023_s 0.00176461f $X=1.885 $Y=1.17 $X2=0
+ $Y2=0
cc_435 N_A_27_65#_c_716_n N_VGND_c_787_n 0.0236214f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_436 N_A_27_65#_c_717_n N_VGND_c_787_n 0.0170777f $X=1.025 $Y=1.17 $X2=0 $Y2=0
cc_437 N_A_27_65#_c_719_n N_VGND_c_787_n 0.0236157f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_438 N_A_27_65#_c_719_n N_VGND_c_788_n 0.0236157f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_439 N_A_27_65#_c_720_n N_VGND_c_788_n 0.0170777f $X=1.885 $Y=1.17 $X2=0 $Y2=0
cc_440 N_A_27_65#_c_722_n N_VGND_c_788_n 0.00915965f $X=2.075 $Y=0.35 $X2=0
+ $Y2=0
cc_441 N_A_27_65#_c_716_n N_VGND_c_789_n 0.0107715f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_442 N_A_27_65#_c_719_n N_VGND_c_790_n 0.0102275f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_443 N_A_27_65#_c_721_n N_VGND_c_791_n 0.0397112f $X=2.745 $Y=0.35 $X2=0 $Y2=0
cc_444 N_A_27_65#_c_722_n N_VGND_c_791_n 0.0128106f $X=2.075 $Y=0.35 $X2=0 $Y2=0
cc_445 N_A_27_65#_c_723_n N_VGND_c_791_n 0.0403449f $X=3.615 $Y=0.35 $X2=0 $Y2=0
cc_446 N_A_27_65#_c_725_n N_VGND_c_791_n 0.0126918f $X=2.84 $Y=0.35 $X2=0 $Y2=0
cc_447 N_A_27_65#_c_726_n N_VGND_c_791_n 0.0208271f $X=3.78 $Y=0.35 $X2=0 $Y2=0
cc_448 N_A_27_65#_c_716_n N_VGND_c_792_n 0.00750444f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_449 N_A_27_65#_c_719_n N_VGND_c_792_n 0.00712543f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_450 N_A_27_65#_c_721_n N_VGND_c_792_n 0.0236582f $X=2.745 $Y=0.35 $X2=0 $Y2=0
cc_451 N_A_27_65#_c_722_n N_VGND_c_792_n 0.0073517f $X=2.075 $Y=0.35 $X2=0 $Y2=0
cc_452 N_A_27_65#_c_723_n N_VGND_c_792_n 0.0240361f $X=3.615 $Y=0.35 $X2=0 $Y2=0
cc_453 N_A_27_65#_c_725_n N_VGND_c_792_n 0.00732706f $X=2.84 $Y=0.35 $X2=0 $Y2=0
cc_454 N_A_27_65#_c_726_n N_VGND_c_792_n 0.0124284f $X=3.78 $Y=0.35 $X2=0 $Y2=0
cc_455 N_A_27_65#_c_721_n N_A_454_65#_M1006_s 0.00176461f $X=2.745 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_456 N_A_27_65#_c_723_n N_A_454_65#_M1018_s 0.00176461f $X=3.615 $Y=0.35 $X2=0
+ $Y2=0
cc_457 N_A_27_65#_c_721_n N_A_454_65#_c_872_n 0.0158608f $X=2.745 $Y=0.35 $X2=0
+ $Y2=0
cc_458 N_A_27_65#_M1009_d N_A_454_65#_c_868_n 0.00176461f $X=2.7 $Y=0.325 $X2=0
+ $Y2=0
cc_459 N_A_27_65#_c_721_n N_A_454_65#_c_868_n 0.00297369f $X=2.745 $Y=0.35 $X2=0
+ $Y2=0
cc_460 N_A_27_65#_c_779_p N_A_454_65#_c_868_n 0.0133685f $X=2.84 $Y=0.7 $X2=0
+ $Y2=0
cc_461 N_A_27_65#_c_723_n N_A_454_65#_c_868_n 0.00298563f $X=3.615 $Y=0.35 $X2=0
+ $Y2=0
cc_462 N_A_27_65#_c_720_n N_A_454_65#_c_869_n 0.00690488f $X=1.885 $Y=1.17 $X2=0
+ $Y2=0
cc_463 N_A_27_65#_M1030_d N_A_454_65#_c_870_n 0.00822145f $X=3.56 $Y=0.325 $X2=0
+ $Y2=0
cc_464 N_A_27_65#_c_723_n N_A_454_65#_c_870_n 0.00463083f $X=3.615 $Y=0.35 $X2=0
+ $Y2=0
cc_465 N_A_27_65#_c_726_n N_A_454_65#_c_870_n 0.0230135f $X=3.78 $Y=0.35 $X2=0
+ $Y2=0
cc_466 N_A_27_65#_c_723_n N_A_454_65#_c_871_n 0.0158608f $X=3.615 $Y=0.35 $X2=0
+ $Y2=0
cc_467 N_A_27_65#_c_726_n N_A_843_67#_c_920_n 0.0195142f $X=3.78 $Y=0.35 $X2=0
+ $Y2=0
cc_468 N_VGND_c_791_n N_A_454_65#_c_870_n 0.00368137f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_792_n N_A_454_65#_c_870_n 0.0100985f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_470 N_VGND_c_791_n N_A_843_67#_c_920_n 0.10479f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_471 N_VGND_c_792_n N_A_843_67#_c_920_n 0.0646156f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_472 N_VGND_c_791_n N_A_843_67#_c_921_n 0.0374727f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_792_n N_A_843_67#_c_921_n 0.0234973f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_474 N_VGND_c_791_n N_A_843_67#_c_922_n 0.0540166f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_475 N_VGND_c_792_n N_A_843_67#_c_922_n 0.033508f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_476 N_VGND_c_791_n N_A_843_67#_c_924_n 0.0120354f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_477 N_VGND_c_792_n N_A_843_67#_c_924_n 0.00730317f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_478 N_VGND_c_791_n N_A_843_67#_c_925_n 0.0120354f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_479 N_VGND_c_792_n N_A_843_67#_c_925_n 0.00730317f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_480 N_A_454_65#_c_870_n N_A_843_67#_M1013_s 0.00546004f $X=5.65 $Y=0.83
+ $X2=-0.19 $Y2=-0.245
cc_481 N_A_454_65#_c_870_n N_A_843_67#_M1014_s 0.00335727f $X=5.65 $Y=0.83 $X2=0
+ $Y2=0
cc_482 N_A_454_65#_M1013_d N_A_843_67#_c_920_n 0.00180013f $X=4.65 $Y=0.335
+ $X2=0 $Y2=0
cc_483 N_A_454_65#_M1020_d N_A_843_67#_c_920_n 0.00180013f $X=5.51 $Y=0.335
+ $X2=0 $Y2=0
cc_484 N_A_454_65#_c_870_n N_A_843_67#_c_920_n 0.0870117f $X=5.65 $Y=0.83 $X2=0
+ $Y2=0
