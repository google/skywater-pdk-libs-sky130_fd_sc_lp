* File: sky130_fd_sc_lp__o2111ai_lp.pex.spice
* Created: Wed Sep  2 10:13:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111AI_LP%D1 3 7 11 12 13 16 17
c37 17 0 1.15577e-20 $X=0.67 $Y=1.07
c38 3 0 1.06792e-19 $X=0.68 $Y=2.545
r39 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.67
+ $Y=1.07 $X2=0.67 $Y2=1.07
r40 13 17 8.10312 $w=3.18e-07 $l=2.25e-07 $layer=LI1_cond $X=0.675 $Y=1.295
+ $X2=0.675 $Y2=1.07
r41 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.67 $Y=1.41
+ $X2=0.67 $Y2=1.07
r42 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=1.41
+ $X2=0.67 $Y2=1.575
r43 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=0.905
+ $X2=0.67 $Y2=1.07
r44 7 10 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.76 $Y=0.495
+ $X2=0.76 $Y2=0.905
r45 3 12 241 $w=2.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.68 $Y=2.545 $X2=0.68
+ $Y2=1.575
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_LP%C1 3 5 7 11 12 13 14 19
c49 12 0 6.50813e-20 $X=1.2 $Y=0.555
c50 7 0 1.01005e-19 $X=1.21 $Y=2.545
c51 3 0 1.15577e-20 $X=1.15 $Y=0.495
r52 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.21
+ $Y=1.08 $X2=1.21 $Y2=1.08
r53 14 20 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.21 $Y=1.295
+ $X2=1.21 $Y2=1.08
r54 13 20 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.21 $Y=0.925
+ $X2=1.21 $Y2=1.08
r55 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.21 $Y=0.555
+ $X2=1.21 $Y2=0.925
r56 11 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.21 $Y=1.42
+ $X2=1.21 $Y2=1.08
r57 10 19 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.21 $Y=0.915
+ $X2=1.21 $Y2=1.08
r58 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.21 $Y=1.585
+ $X2=1.21 $Y2=1.42
r59 5 7 238.515 $w=2.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.21 $Y=1.585 $X2=1.21
+ $Y2=2.545
r60 3 10 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.15 $Y=0.495
+ $X2=1.15 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_LP%B1 3 7 11 12 13 14 18
c42 12 0 2.73319e-20 $X=1.75 $Y=1.795
c43 7 0 1.93845e-19 $X=1.76 $Y=2.545
r44 13 14 12.7108 $w=3.38e-07 $l=3.75e-07 $layer=LI1_cond $X=1.735 $Y=1.29
+ $X2=1.735 $Y2=1.665
r45 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.75
+ $Y=1.29 $X2=1.75 $Y2=1.29
r46 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.75 $Y=1.63
+ $X2=1.75 $Y2=1.29
r47 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.63
+ $X2=1.75 $Y2=1.795
r48 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.125
+ $X2=1.75 $Y2=1.29
r49 7 12 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.76 $Y=2.545 $X2=1.76
+ $Y2=1.795
r50 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.66 $Y=0.495
+ $X2=1.66 $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_LP%A2 3 5 7 11 12 13 17 18
c41 17 0 1.77943e-19 $X=2.29 $Y=1.29
r42 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.29 $X2=2.29 $Y2=1.29
r43 12 13 7.13789 $w=6.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.435 $Y=1.295
+ $X2=2.435 $Y2=1.665
r44 12 18 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=2.435 $Y=1.295
+ $X2=2.435 $Y2=1.29
r45 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.29 $Y=1.63
+ $X2=2.29 $Y2=1.29
r46 10 17 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.125
+ $X2=2.29 $Y2=1.29
r47 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.795
+ $X2=2.29 $Y2=1.63
r48 5 7 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.29 $Y=1.795 $X2=2.29
+ $Y2=2.545
r49 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.23 $Y=0.495
+ $X2=2.23 $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_LP%A1 3 7 9 10 17
c29 9 0 1.77943e-19 $X=3.12 $Y=1.295
r30 15 17 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.79 $Y=1.345 $X2=3.09
+ $Y2=1.345
r31 13 15 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.77 $Y=1.345 $X2=2.79
+ $Y2=1.345
r32 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.665
r33 9 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.345 $X2=3.09 $Y2=1.345
r34 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.18
+ $X2=2.77 $Y2=1.345
r35 5 7 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.77 $Y=1.18 $X2=2.77
+ $Y2=0.495
r36 1 15 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.51
+ $X2=2.79 $Y2=1.345
r37 1 3 257.149 $w=2.5e-07 $l=1.035e-06 $layer=POLY_cond $X=2.79 $Y=1.51
+ $X2=2.79 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_LP%VPWR 1 2 3 10 12 16 18 20 25 26 27 33 45
r41 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r46 33 44 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=3.125 $Y2=3.33
r47 33 38 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 32 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 29 41 4.50438 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=0.58 $Y=3.33 $X2=0.29
+ $Y2=3.33
r51 29 31 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=0.58 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 27 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 27 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 27 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 25 31 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.31 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=3.33
+ $X2=1.475 $Y2=3.33
r57 24 35 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.64 $Y=3.33 $X2=1.68
+ $Y2=3.33
r58 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.64 $Y=3.33
+ $X2=1.475 $Y2=3.33
r59 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.055 $Y=2.19
+ $X2=3.055 $Y2=2.9
r60 18 44 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.055 $Y=3.245
+ $X2=3.125 $Y2=3.33
r61 18 23 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.055 $Y=3.245
+ $X2=3.055 $Y2=2.9
r62 14 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=3.245
+ $X2=1.475 $Y2=3.33
r63 14 16 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=1.475 $Y=3.245
+ $X2=1.475 $Y2=2.49
r64 10 41 3.26179 $w=3.3e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.415 $Y=3.245
+ $X2=0.29 $Y2=3.33
r65 10 12 33.7002 $w=3.28e-07 $l=9.65e-07 $layer=LI1_cond $X=0.415 $Y=3.245
+ $X2=0.415 $Y2=2.28
r66 3 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.915
+ $Y=2.045 $X2=3.055 $Y2=2.9
r67 3 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.915
+ $Y=2.045 $X2=3.055 $Y2=2.19
r68 2 16 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=1.335
+ $Y=2.045 $X2=1.475 $Y2=2.49
r69 1 12 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=0.27
+ $Y=2.045 $X2=0.415 $Y2=2.28
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_LP%Y 1 2 3 10 11 14 18 22 27 30 31 32 33 50
c58 27 0 2.73319e-20 $X=0.945 $Y=1.85
c59 18 0 4.17108e-20 $X=1.86 $Y=2.06
c60 14 0 1.93845e-19 $X=0.945 $Y=2.19
c61 10 0 1.01005e-19 $X=0.78 $Y=1.85
r62 38 45 5.34566 $w=2.1e-07 $l=2.3e-07 $layer=LI1_cond $X=0.23 $Y=0.725
+ $X2=0.23 $Y2=0.495
r63 32 33 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.665
r64 31 32 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=0.925
+ $X2=0.23 $Y2=1.295
r65 31 38 10.5628 $w=2.08e-07 $l=2e-07 $layer=LI1_cond $X=0.23 $Y=0.925 $X2=0.23
+ $Y2=0.725
r66 30 50 7.93052 $w=4.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.24 $Y=0.495
+ $X2=0.545 $Y2=0.495
r67 30 45 0.260017 $w=4.58e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=0.495
+ $X2=0.23 $Y2=0.495
r68 27 29 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.945 $Y=1.85
+ $X2=0.945 $Y2=2.06
r69 26 33 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=0.23 $Y=1.765 $X2=0.23
+ $Y2=1.665
r70 22 24 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.025 $Y=2.19
+ $X2=2.025 $Y2=2.9
r71 20 22 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.025 $Y=2.145
+ $X2=2.025 $Y2=2.19
r72 19 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.11 $Y=2.06
+ $X2=0.945 $Y2=2.06
r73 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.86 $Y=2.06
+ $X2=2.025 $Y2=2.145
r74 18 19 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.86 $Y=2.06
+ $X2=1.11 $Y2=2.06
r75 14 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.945 $Y=2.19
+ $X2=0.945 $Y2=2.9
r76 12 29 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.945 $Y=2.145
+ $X2=0.945 $Y2=2.06
r77 12 14 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.945 $Y=2.145
+ $X2=0.945 $Y2=2.19
r78 11 26 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.335 $Y=1.85
+ $X2=0.23 $Y2=1.765
r79 10 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=1.85
+ $X2=0.945 $Y2=1.85
r80 10 11 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.78 $Y=1.85
+ $X2=0.335 $Y2=1.85
r81 3 24 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.885
+ $Y=2.045 $X2=2.025 $Y2=2.9
r82 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.885
+ $Y=2.045 $X2=2.025 $Y2=2.19
r83 2 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.805
+ $Y=2.045 $X2=0.945 $Y2=2.9
r84 2 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.805
+ $Y=2.045 $X2=0.945 $Y2=2.19
r85 1 50 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.4
+ $Y=0.285 $X2=0.545 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_LP%A_347_57# 1 2 9 11 12 15
r27 13 15 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.985 $Y=0.775
+ $X2=2.985 $Y2=0.495
r28 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.82 $Y=0.86
+ $X2=2.985 $Y2=0.775
r29 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.82 $Y=0.86 $X2=2.13
+ $Y2=0.86
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.965 $Y=0.775
+ $X2=2.13 $Y2=0.86
r31 7 9 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.965 $Y=0.775
+ $X2=1.965 $Y2=0.495
r32 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.845
+ $Y=0.285 $X2=2.985 $Y2=0.495
r33 1 9 182 $w=1.7e-07 $l=3.18119e-07 $layer=licon1_NDIFF $count=1 $X=1.735
+ $Y=0.285 $X2=1.965 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_LP%VGND 1 6 9 10 11 21 22
r29 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r30 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r31 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r32 14 18 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r33 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r34 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r35 11 15 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r36 9 18 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.16
+ $Y2=0
r37 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.475
+ $Y2=0
r38 8 21 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r39 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.475
+ $Y2=0
r40 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0
r41 4 6 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0.43
r42 1 6 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.285 $X2=2.475 $Y2=0.43
.ends

