* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__isobufsrc_4 A SLEEP VGND VNB VPB VPWR X
X0 a_245_367# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 X a_60_47# a_245_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_60_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 X a_60_47# a_245_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR SLEEP a_245_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND a_60_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VPWR SLEEP a_245_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_245_367# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_60_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_245_367# a_60_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 X a_60_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_245_367# a_60_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 X a_60_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VGND a_60_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
