* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 VPWR a_808_463# a_936_333# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 Q a_2431_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_1406_69# a_864_255# a_1593_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_225_50# a_35_74# a_308_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_380_50# a_864_255# a_808_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1809_119# a_1406_69# a_1635_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_490_468# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VPWR RESET_B a_808_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_936_333# a_864_255# a_1406_69# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_512_81# SCD a_225_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_332_468# D a_380_50# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VGND CLK a_864_255# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_380_50# a_756_265# a_808_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_2431_47# a_1406_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VGND a_808_463# a_936_333# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 VPWR RESET_B a_1635_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_808_463# a_756_265# a_991_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_308_50# D a_380_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_225_50# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_756_265# a_864_255# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_1569_534# a_1635_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_2431_47# a_1406_69# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR CLK a_864_255# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_35_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_380_50# a_35_74# a_490_468# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_35_74# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND a_2431_47# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_808_463# a_864_255# a_894_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_894_463# a_936_333# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 Q a_2431_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 a_380_50# SCE a_512_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_936_333# a_756_265# a_1406_69# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 a_1635_21# a_1406_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 VPWR a_2431_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 a_1085_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_991_119# a_936_333# a_1085_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_1593_113# a_1635_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VPWR SCE a_332_468# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X38 VGND RESET_B a_1809_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1406_69# a_756_265# a_1569_534# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X40 VPWR RESET_B a_380_50# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X41 a_756_265# a_864_255# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
