* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a211o_m A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VGND B1 a_82_483# VNB nshort w=420000u l=150000u
+  ad=5.145e+11p pd=4.13e+06u as=2.289e+11p ps=2.77e+06u
M1001 a_322_145# A2 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1002 VPWR A2 a_225_389# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.289e+11p ps=2.77e+06u
M1003 a_480_389# B1 a_225_389# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_82_483# C1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_82_483# C1 a_480_389# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 VPWR a_82_483# X VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 VGND a_82_483# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 a_225_389# A1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_82_483# A1 a_322_145# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
