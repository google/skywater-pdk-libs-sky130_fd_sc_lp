* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
X0 VPWR a_1039_367# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 GCLK a_1039_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_33_47# a_78_269# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_258_81# a_300_55# a_78_269# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1039_367# a_33_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 GCLK a_1039_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_416_81# a_33_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_300_55# a_284_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_78_269# a_300_55# a_422_465# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_300_55# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_422_465# a_33_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_242_465# a_284_367# a_78_269# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 VPWR CLK a_1039_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VGND CLK a_1002_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_33_47# a_78_269# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND GATE a_258_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_78_269# a_284_367# a_416_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_300_55# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_1002_133# a_33_47# a_1039_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_1039_367# GCLK VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VPWR GATE a_242_465# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VPWR a_300_55# a_284_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
