# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand4_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nand4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.220000 1.425000 8.005000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.980000 1.425000 6.010000 1.750000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.425000 3.450000 1.750000 ;
        RECT 2.200000 1.380000 3.450000 1.425000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.425000 1.765000 1.750000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.292800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.920000 7.465000 2.090000 ;
        RECT 0.610000 2.090000 1.765000 2.120000 ;
        RECT 0.610000 2.120000 0.835000 3.075000 ;
        RECT 1.505000 2.120000 1.765000 3.075000 ;
        RECT 2.445000 2.090000 2.715000 3.075000 ;
        RECT 3.385000 2.090000 3.575000 3.075000 ;
        RECT 3.630000 1.085000 7.535000 1.255000 ;
        RECT 3.630000 1.255000 3.800000 1.920000 ;
        RECT 4.245000 2.090000 4.435000 3.075000 ;
        RECT 5.105000 2.090000 5.295000 3.075000 ;
        RECT 6.345000 0.625000 6.675000 1.085000 ;
        RECT 6.415000 2.090000 6.605000 3.075000 ;
        RECT 7.205000 0.625000 7.535000 1.085000 ;
        RECT 7.275000 2.090000 7.465000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.145000  1.920000 0.440000 3.245000 ;
      RECT 0.155000  0.305000 0.355000 1.085000 ;
      RECT 0.155000  1.085000 2.075000 1.255000 ;
      RECT 0.525000  0.085000 0.855000 0.915000 ;
      RECT 1.005000  2.290000 1.335000 3.245000 ;
      RECT 1.025000  0.305000 1.215000 1.085000 ;
      RECT 1.385000  0.085000 1.715000 0.915000 ;
      RECT 1.885000  0.265000 3.945000 0.435000 ;
      RECT 1.885000  0.435000 2.075000 1.085000 ;
      RECT 1.945000  2.260000 2.275000 3.245000 ;
      RECT 2.245000  0.605000 2.575000 1.035000 ;
      RECT 2.245000  1.035000 3.435000 1.205000 ;
      RECT 2.745000  0.435000 2.935000 0.865000 ;
      RECT 2.885000  2.260000 3.215000 3.245000 ;
      RECT 3.105000  0.605000 3.435000 0.745000 ;
      RECT 3.105000  0.745000 5.815000 0.915000 ;
      RECT 3.105000  0.915000 3.435000 1.035000 ;
      RECT 3.615000  0.435000 3.945000 0.565000 ;
      RECT 3.745000  2.260000 4.075000 3.245000 ;
      RECT 4.195000  0.275000 7.965000 0.445000 ;
      RECT 4.195000  0.445000 6.175000 0.575000 ;
      RECT 4.605000  2.260000 4.935000 3.245000 ;
      RECT 5.465000  2.260000 6.245000 3.245000 ;
      RECT 5.985000  0.575000 6.175000 0.915000 ;
      RECT 6.775000  2.260000 7.105000 3.245000 ;
      RECT 6.845000  0.445000 7.035000 0.915000 ;
      RECT 7.635000  1.920000 7.965000 3.245000 ;
      RECT 7.705000  0.445000 7.965000 1.195000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__nand4_4
END LIBRARY
