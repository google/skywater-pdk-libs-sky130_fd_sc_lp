* File: sky130_fd_sc_lp__and3_1.spice
* Created: Wed Sep  2 09:31:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and3_1.pex.spice"
.subckt sky130_fd_sc_lp__and3_1  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_149_53# N_A_M1002_g N_A_61_367#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1113 PD=0.66 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1006 A_227_53# N_B_M1006_g A_149_53# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0504 PD=0.81 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_C_M1004_g A_227_53# VNB NSHORT L=0.15 W=0.42 AD=0.0994
+ AS=0.0819 PD=0.856667 PS=0.81 NRD=25.704 NRS=39.996 M=1 R=2.8 SA=75001.1
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_61_367#_M1001_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1988 PD=2.21 PS=1.71333 NRD=0 NRS=10.704 M=1 R=5.6 SA=75001
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_61_367#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.1113 PD=0.72 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_61_367#_M1007_d N_B_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.07455 AS=0.063 PD=0.775 PS=0.72 NRD=9.3772 NRS=9.3772 M=1 R=2.8
+ SA=75000.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_A_61_367#_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.122325 AS=0.07455 PD=0.9475 PS=0.775 NRD=100.844 NRS=25.7873 M=1 R=2.8
+ SA=75001.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_61_367#_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.366975 PD=3.05 PS=2.8425 NRD=0 NRS=7.289 M=1 R=8.4 SA=75000.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__and3_1.pxi.spice"
*
.ends
*
*
