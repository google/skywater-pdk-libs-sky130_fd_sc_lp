* NGSPICE file created from sky130_fd_sc_lp__o211ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=8.253e+11p pd=6.35e+06u as=1.2537e+12p ps=7.03e+06u
M1001 VGND A1 a_27_47# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=5.502e+11p ps=4.67e+06u
M1002 a_27_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y C1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_326_47# B1 a_27_47# VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1005 Y C1 a_326_47# VNB nshort w=840000u l=150000u
+  ad=5.082e+11p pd=2.89e+06u as=0p ps=0u
M1006 Y A2 a_110_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1007 a_110_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

