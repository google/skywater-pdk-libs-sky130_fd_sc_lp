* File: sky130_fd_sc_lp__and2_m.pex.spice
* Created: Wed Sep  2 09:30:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2_M%A 3 5 7 9 10
c24 9 0 6.54564e-20 $X=0.24 $Y=1.295
r25 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.46 $X2=0.35 $Y2=1.46
r26 10 15 8.43753 $w=2.78e-07 $l=2.05e-07 $layer=LI1_cond $X=0.295 $Y=1.665
+ $X2=0.295 $Y2=1.46
r27 9 15 6.79118 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.295 $Y=1.295
+ $X2=0.295 $Y2=1.46
r28 5 14 57.1555 $w=4.23e-07 $l=3.88034e-07 $layer=POLY_cond $X=0.585 $Y=1.775
+ $X2=0.422 $Y2=1.46
r29 5 7 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.585 $Y=1.775
+ $X2=0.585 $Y2=2.195
r30 1 14 40.0633 $w=4.23e-07 $l=2.04316e-07 $layer=POLY_cond $X=0.51 $Y=1.295
+ $X2=0.422 $Y2=1.46
r31 1 3 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.51 $Y=1.295 $X2=0.51
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_M%B 4 7 11 13 14 18 19
c29 19 0 1.58809e-19 $X=0.96 $Y=0.43
c30 11 0 6.54564e-20 $X=1.015 $Y=1.31
c31 7 0 4.4852e-21 $X=1.015 $Y=2.195
r32 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=0.43
+ $X2=0.96 $Y2=0.595
r33 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=0.43 $X2=0.96 $Y2=0.43
r34 14 19 7.37564 $w=3.73e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=0.452
+ $X2=0.96 $Y2=0.452
r35 13 14 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=0.452
+ $X2=0.72 $Y2=0.452
r36 9 11 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.87 $Y=1.31
+ $X2=1.015 $Y2=1.31
r37 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.015 $Y=1.385
+ $X2=1.015 $Y2=1.31
r38 5 7 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.015 $Y=1.385
+ $X2=1.015 $Y2=2.195
r39 4 21 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.87 $Y=0.915
+ $X2=0.87 $Y2=0.595
r40 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.87 $Y=1.235 $X2=0.87
+ $Y2=1.31
r41 2 4 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.87 $Y=1.235 $X2=0.87
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_M%A_34_141# 1 2 7 11 14 15 21 26
c47 11 0 1.58809e-19 $X=1.445 $Y=0.915
r48 24 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.78 $Y=2.94 $X2=0.78
+ $Y2=2.85
r49 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.78
+ $Y=2.94 $X2=0.78 $Y2=2.94
r50 21 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.78 $Y=2.26
+ $X2=0.78 $Y2=2.94
r51 19 21 42.9547 $w=3.28e-07 $l=1.23e-06 $layer=LI1_cond $X=0.78 $Y=1.03
+ $X2=0.78 $Y2=2.26
r52 15 19 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=0.615 $Y=0.925
+ $X2=0.78 $Y2=1.03
r53 15 17 16.9004 $w=2.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.615 $Y=0.925
+ $X2=0.295 $Y2=0.925
r54 11 14 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=1.445 $Y=0.915
+ $X2=1.445 $Y2=2.195
r55 9 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.445 $Y=2.775
+ $X2=1.445 $Y2=2.195
r56 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=2.85
+ $X2=0.78 $Y2=2.85
r57 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.37 $Y=2.85
+ $X2=1.445 $Y2=2.775
r58 7 8 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=1.37 $Y=2.85
+ $X2=0.945 $Y2=2.85
r59 2 21 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.985 $X2=0.8 $Y2=2.26
r60 1 17 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.705 $X2=0.295 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_M%VPWR 1 2 7 9 11 15 17 21 22 28
c29 22 0 4.4852e-21 $X=1.68 $Y=3.33
r30 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r31 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 22 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 19 28 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.23 $Y2=3.33
r35 19 21 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 17 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r37 17 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 13 28 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r39 13 15 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.26
r40 12 25 3.64968 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=3.33 $X2=0.19
+ $Y2=3.33
r41 11 28 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=1.23 $Y2=3.33
r42 11 12 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=0.38 $Y2=3.33
r43 7 25 3.26551 $w=2.1e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.19 $Y2=3.33
r44 7 9 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.26
r45 2 15 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.985 $X2=1.23 $Y2=2.26
r46 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.985 $X2=0.275 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_M%X 1 2 7 8 9 10 11 12 13
r10 12 13 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.67 $Y=2.405
+ $X2=1.67 $Y2=2.775
r11 12 34 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.67 $Y=2.405
+ $X2=1.67 $Y2=2.26
r12 11 34 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=1.67 $Y=2.035
+ $X2=1.67 $Y2=2.26
r13 10 11 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=2.035
r14 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.67 $Y=1.295
+ $X2=1.67 $Y2=1.665
r15 8 9 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=1.67 $Y=0.85 $X2=1.67
+ $Y2=1.295
r16 7 8 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.67 $Y=0.555
+ $X2=1.67 $Y2=0.85
r17 2 34 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.985 $X2=1.66 $Y2=2.26
r18 1 8 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.705 $X2=1.66 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_M%VGND 1 7 8 11 12 13 23 24
r25 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r26 21 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r27 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r28 16 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r29 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r30 13 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r31 13 17 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r32 11 20 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.2
+ $Y2=0
r33 11 12 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.31
+ $Y2=0
r34 10 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.68
+ $Y2=0
r35 10 12 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.31
+ $Y2=0
r36 7 8 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.26 $Y=0.985
+ $X2=1.26 $Y2=0.82
r37 4 12 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=0.085 $X2=1.31
+ $Y2=0
r38 4 8 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.31 $Y=0.085
+ $X2=1.31 $Y2=0.82
r39 1 7 182 $w=1.7e-07 $l=4.01279e-07 $layer=licon1_NDIFF $count=1 $X=0.945
+ $Y=0.705 $X2=1.23 $Y2=0.985
.ends

