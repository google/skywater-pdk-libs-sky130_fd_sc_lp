* File: sky130_fd_sc_lp__o32a_1.spice
* Created: Wed Sep  2 10:25:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32a_1.pex.spice"
.subckt sky130_fd_sc_lp__o32a_1  VNB VPB A1 A2 A3 B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_88_269#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1386 AS=0.2394 PD=1.17 PS=2.25 NRD=3.564 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1006 N_A_250_69#_M1006_d N_A1_M1006_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1386 PD=1.12 PS=1.17 NRD=0 NRS=3.564 M=1 R=5.6 SA=75000.7
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_250_69#_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1003 N_A_250_69#_M1003_d N_A3_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2604 PD=1.12 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_88_269#_M1000_d N_B2_M1000_g N_A_250_69#_M1003_d VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=6.42 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1011 N_A_250_69#_M1011_d N_B1_M1011_g N_A_88_269#_M1000_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2604 AS=0.147 PD=2.3 PS=1.19 NRD=3.564 NRS=3.564 M=1 R=5.6
+ SA=75002.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_A_88_269#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.25515 AS=0.3591 PD=1.665 PS=3.09 NRD=9.3772 NRS=3.1126 M=1 R=8.4
+ SA=75000.2 SB=75002.8 A=0.189 P=2.82 MULT=1
MM1010 A_264_367# N_A1_M1010_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.25515 PD=1.58 PS=1.665 NRD=16.4101 NRS=10.1455 M=1 R=8.4
+ SA=75000.8 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1008 A_358_367# N_A2_M1008_g A_264_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.1953
+ AS=0.2016 PD=1.57 PS=1.58 NRD=15.6221 NRS=16.4101 M=1 R=8.4 SA=75001.2
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1007 N_A_88_269#_M1007_d N_A3_M1007_g A_358_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.1953 PD=1.88 PS=1.57 NRD=0 NRS=15.6221 M=1 R=8.4 SA=75001.7
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1002 A_604_367# N_B2_M1002_g N_A_88_269#_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3906 PD=1.47 PS=1.88 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_B1_M1005_g A_604_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75002.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o32a_1.pxi.spice"
*
.ends
*
*
