* File: sky130_fd_sc_lp__or4bb_1.pex.spice
* Created: Wed Sep  2 10:33:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4BB_1%C_N 3 7 9 10 11 12 13 17
c40 17 0 1.54048e-19 $X=0.53 $Y=0.93
c41 12 0 1.26363e-19 $X=0.72 $Y=0.925
r42 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.53
+ $Y=0.93 $X2=0.53 $Y2=0.93
r43 13 18 9.00141 $w=4.83e-07 $l=3.65e-07 $layer=LI1_cond $X=0.677 $Y=1.295
+ $X2=0.677 $Y2=0.93
r44 12 18 0.123307 $w=4.83e-07 $l=5e-09 $layer=LI1_cond $X=0.677 $Y=0.925
+ $X2=0.677 $Y2=0.93
r45 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.53 $Y=1.27
+ $X2=0.53 $Y2=0.93
r46 10 11 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.27
+ $X2=0.53 $Y2=1.435
r47 9 17 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=0.765
+ $X2=0.53 $Y2=0.93
r48 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.55 $Y=0.445 $X2=0.55
+ $Y2=0.765
r49 3 11 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=0.475 $Y=2.885
+ $X2=0.475 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_1%D_N 3 7 12 13 14 18 20
c40 12 0 1.26363e-19 $X=0.995 $Y=1.585
r41 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=2.22
+ $X2=0.955 $Y2=2.385
r42 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=2.22
+ $X2=0.955 $Y2=2.055
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.955
+ $Y=2.22 $X2=0.955 $Y2=2.22
r44 14 19 5.80276 $w=5.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.2 $Y=2.297
+ $X2=0.955 $Y2=2.297
r45 13 19 5.56591 $w=5.03e-07 $l=2.35e-07 $layer=LI1_cond $X=0.72 $Y=2.297
+ $X2=0.955 $Y2=2.297
r46 12 20 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.01 $Y=1.585 $X2=1.01
+ $Y2=2.055
r47 11 12 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.995 $Y=1.435
+ $X2=0.995 $Y2=1.585
r48 7 11 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=0.98 $Y=0.445
+ $X2=0.98 $Y2=1.435
r49 3 21 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.905 $Y=2.885
+ $X2=0.905 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_1%A_196_535# 1 2 8 10 13 16 21 27 28 32 39 40
+ 47
c70 39 0 9.78455e-20 $X=1.695 $Y=0.93
r71 40 47 47.6426 $w=4.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.767 $Y=0.93
+ $X2=1.767 $Y2=0.765
r72 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.695
+ $Y=0.93 $X2=1.695 $Y2=0.93
r73 30 39 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.225 $Y=0.86
+ $X2=1.695 $Y2=0.86
r74 30 32 14.0854 $w=2.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.225 $Y=0.775
+ $X2=1.225 $Y2=0.445
r75 28 42 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.62 $Y=2.92
+ $X2=1.415 $Y2=2.92
r76 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=2.92 $X2=1.62 $Y2=2.92
r77 24 27 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=1.12 $Y=2.885 $X2=1.62
+ $Y2=2.885
r78 14 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2 $Y=1.435 $X2=2
+ $Y2=1.36
r79 14 16 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2 $Y=1.435 $X2=2
+ $Y2=2.165
r80 13 47 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.93 $Y=0.445
+ $X2=1.93 $Y2=0.765
r81 10 21 119.474 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.767 $Y=1.36 $X2=2
+ $Y2=1.36
r82 10 18 180.494 $w=1.5e-07 $l=3.52e-07 $layer=POLY_cond $X=1.767 $Y=1.36
+ $X2=1.415 $Y2=1.36
r83 9 40 8.43012 $w=4.75e-07 $l=7.2e-08 $layer=POLY_cond $X=1.767 $Y=1.002
+ $X2=1.767 $Y2=0.93
r84 9 10 33.1351 $w=4.75e-07 $l=2.83e-07 $layer=POLY_cond $X=1.767 $Y=1.002
+ $X2=1.767 $Y2=1.285
r85 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=2.755
+ $X2=1.415 $Y2=2.92
r86 7 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.415 $Y=1.435
+ $X2=1.415 $Y2=1.36
r87 7 8 676.851 $w=1.5e-07 $l=1.32e-06 $layer=POLY_cond $X=1.415 $Y=1.435
+ $X2=1.415 $Y2=2.755
r88 2 24 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.675 $X2=1.12 $Y2=2.885
r89 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.055
+ $Y=0.235 $X2=1.195 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_1%A_27_535# 1 2 9 14 16 17 19 22 29 31 33 34
+ 35 38
c81 17 0 9.78455e-20 $X=2.345 $Y=0.915
r82 34 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=1.63
+ $X2=2.45 $Y2=1.795
r83 34 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=1.63
+ $X2=2.45 $Y2=1.465
r84 33 35 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.45 $Y=1.665
+ $X2=2.285 $Y2=1.665
r85 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.45
+ $Y=1.63 $X2=2.45 $Y2=1.63
r86 26 29 5.85368 $w=3.13e-07 $l=1.6e-07 $layer=LI1_cond $X=0.175 $Y=0.437
+ $X2=0.335 $Y2=0.437
r87 25 31 2.43474 $w=1.8e-07 $l=1.53e-07 $layer=LI1_cond $X=0.39 $Y=1.705
+ $X2=0.237 $Y2=1.705
r88 25 35 116.763 $w=1.78e-07 $l=1.895e-06 $layer=LI1_cond $X=0.39 $Y=1.705
+ $X2=2.285 $Y2=1.705
r89 20 31 4.00459 $w=2.42e-07 $l=9e-08 $layer=LI1_cond $X=0.237 $Y=1.795
+ $X2=0.237 $Y2=1.705
r90 20 22 41.1857 $w=3.03e-07 $l=1.09e-06 $layer=LI1_cond $X=0.237 $Y=1.795
+ $X2=0.237 $Y2=2.885
r91 19 31 4.00459 $w=2.42e-07 $l=1.16962e-07 $layer=LI1_cond $X=0.175 $Y=1.615
+ $X2=0.237 $Y2=1.705
r92 18 26 4.01183 $w=1.8e-07 $l=1.58e-07 $layer=LI1_cond $X=0.175 $Y=0.595
+ $X2=0.175 $Y2=0.437
r93 18 19 62.8485 $w=1.78e-07 $l=1.02e-06 $layer=LI1_cond $X=0.175 $Y=0.595
+ $X2=0.175 $Y2=1.615
r94 17 38 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.36 $Y=0.915
+ $X2=2.36 $Y2=1.465
r95 16 17 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.345 $Y=0.765
+ $X2=2.345 $Y2=0.915
r96 14 39 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.36 $Y=2.165
+ $X2=2.36 $Y2=1.795
r97 9 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.36 $Y=0.445
+ $X2=2.36 $Y2=0.765
r98 2 22 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.675 $X2=0.26 $Y2=2.885
r99 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.235 $X2=0.335 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_1%B 3 6 8 11 12 13
c36 11 0 1.7683e-19 $X=2.81 $Y=0.93
r37 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=0.93
+ $X2=2.81 $Y2=1.095
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=0.93
+ $X2=2.81 $Y2=0.765
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=0.93 $X2=2.81 $Y2=0.93
r40 8 12 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=2.64 $Y=0.902
+ $X2=2.81 $Y2=0.902
r41 6 14 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.9 $Y=2.165 $X2=2.9
+ $Y2=1.095
r42 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.83 $Y=0.445
+ $X2=2.83 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_1%A 3 6 7 9 11 23
c37 23 0 3.62896e-20 $X=3.26 $Y=2.91
r38 20 23 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.04 $Y=2.91
+ $X2=3.26 $Y2=2.91
r39 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=2.91 $X2=3.04 $Y2=2.91
r40 11 21 1.38676 $w=6.88e-07 $l=8e-08 $layer=LI1_cond $X=3.12 $Y=2.65 $X2=3.04
+ $Y2=2.65
r41 9 21 6.93379 $w=6.88e-07 $l=4e-07 $layer=LI1_cond $X=2.64 $Y=2.65 $X2=3.04
+ $Y2=2.65
r42 7 9 8.32055 $w=6.88e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.65 $X2=2.64
+ $Y2=2.65
r43 3 6 881.957 $w=1.5e-07 $l=1.72e-06 $layer=POLY_cond $X=3.26 $Y=0.445
+ $X2=3.26 $Y2=2.165
r44 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=2.745
+ $X2=3.26 $Y2=2.91
r45 1 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.26 $Y=2.745 $X2=3.26
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_1%A_332_391# 1 2 3 12 16 17 21 24 26 28 29 31
+ 32 34 40 45 48
c91 21 0 1.7683e-19 $X=2.145 $Y=0.445
c92 17 0 3.62896e-20 $X=2.795 $Y=2.05
r93 43 45 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.045 $Y=0.445
+ $X2=3.24 $Y2=0.445
r94 39 41 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.88 $Y=1.36
+ $X2=3.24 $Y2=1.36
r95 39 40 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=1.36
+ $X2=2.795 $Y2=1.36
r96 34 37 4.90855 $w=2.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.755 $Y=2.05
+ $X2=1.755 $Y2=2.165
r97 32 49 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.732 $Y=1.36
+ $X2=3.732 $Y2=1.525
r98 32 48 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.732 $Y=1.36
+ $X2=3.732 $Y2=1.195
r99 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.71
+ $Y=1.36 $X2=3.71 $Y2=1.36
r100 29 41 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=1.36
+ $X2=3.24 $Y2=1.36
r101 29 31 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.325 $Y=1.36
+ $X2=3.71 $Y2=1.36
r102 28 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=1.195
+ $X2=3.24 $Y2=1.36
r103 27 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0.61
+ $X2=3.24 $Y2=0.445
r104 27 28 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.24 $Y=0.61
+ $X2=3.24 $Y2=1.195
r105 25 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=1.525
+ $X2=2.88 $Y2=1.36
r106 25 26 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.88 $Y=1.525
+ $X2=2.88 $Y2=1.965
r107 24 40 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.26 $Y=1.28
+ $X2=2.795 $Y2=1.28
r108 19 24 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.145 $Y=1.195
+ $X2=2.26 $Y2=1.28
r109 19 21 37.5797 $w=2.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.145 $Y=1.195
+ $X2=2.145 $Y2=0.445
r110 18 34 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.89 $Y=2.05
+ $X2=1.755 $Y2=2.05
r111 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.795 $Y=2.05
+ $X2=2.88 $Y2=1.965
r112 17 18 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.795 $Y=2.05
+ $X2=1.89 $Y2=2.05
r113 16 48 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.845 $Y=0.655
+ $X2=3.845 $Y2=1.195
r114 12 49 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.785 $Y=2.465
+ $X2=3.785 $Y2=1.525
r115 3 37 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.66
+ $Y=1.955 $X2=1.785 $Y2=2.165
r116 2 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.905
+ $Y=0.235 $X2=3.045 $Y2=0.445
r117 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.145 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
r42 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r44 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 27 39 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.82 $Y=3.33 $X2=0.69
+ $Y2=3.33
r50 27 29 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 22 39 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.69
+ $Y2=3.33
r54 22 24 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r55 20 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 20 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 18 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 18 19 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.525 $Y2=3.33
r59 17 35 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 17 19 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=3.525 $Y2=3.33
r61 13 16 18.8232 $w=2.98e-07 $l=4.9e-07 $layer=LI1_cond $X=3.525 $Y=1.98
+ $X2=3.525 $Y2=2.47
r62 11 19 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=3.245
+ $X2=3.525 $Y2=3.33
r63 11 16 29.7714 $w=2.98e-07 $l=7.75e-07 $layer=LI1_cond $X=3.525 $Y=3.245
+ $X2=3.525 $Y2=2.47
r64 7 39 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r65 7 9 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.885
r66 2 16 300 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=2 $X=3.335
+ $Y=1.955 $X2=3.57 $Y2=2.47
r67 2 13 600 $w=1.7e-07 $l=2.47184e-07 $layer=licon1_PDIFF $count=1 $X=3.335
+ $Y=1.955 $X2=3.57 $Y2=1.98
r68 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.675 $X2=0.69 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_1%X 1 2 9 13 15 16 17 18 24
r17 17 18 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.1 $Y=1.295 $X2=4.1
+ $Y2=1.665
r18 16 17 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.1 $Y=0.925 $X2=4.1
+ $Y2=1.295
r19 15 16 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.1 $Y=0.555 $X2=4.1
+ $Y2=0.925
r20 15 24 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.1 $Y=0.555
+ $X2=4.1 $Y2=0.42
r21 14 18 6.40246 $w=2.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.1 $Y=1.815 $X2=4.1
+ $Y2=1.665
r22 13 14 6.1139 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=4.065 $Y=1.98
+ $X2=4.065 $Y2=1.815
r23 7 13 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=4.065 $Y=1.985
+ $X2=4.065 $Y2=1.98
r24 7 9 31.3532 $w=3.38e-07 $l=9.25e-07 $layer=LI1_cond $X=4.065 $Y=1.985
+ $X2=4.065 $Y2=2.91
r25 2 13 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=1.835 $X2=4 $Y2=1.98
r26 2 9 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=1.835 $X2=4 $Y2=2.91
r27 1 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.92
+ $Y=0.235 $X2=4.06 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_1%VGND 1 2 3 4 17 21 25 29 33 35 40 45 52 53
+ 56 59 62 65
c74 17 0 1.54048e-19 $X=0.765 $Y=0.43
r75 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r76 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r77 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r78 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r79 53 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r80 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r81 50 65 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.645
+ $Y2=0
r82 50 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=4.08
+ $Y2=0
r83 49 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r84 49 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r85 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r86 46 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=2.595
+ $Y2=0
r87 46 48 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=3.12
+ $Y2=0
r88 45 65 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.645
+ $Y2=0
r89 45 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.12
+ $Y2=0
r90 41 59 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.705
+ $Y2=0
r91 41 43 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=2.16
+ $Y2=0
r92 40 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.595
+ $Y2=0
r93 40 43 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.16
+ $Y2=0
r94 39 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r95 39 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r96 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r97 36 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=0.795
+ $Y2=0
r98 36 38 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=1.2
+ $Y2=0
r99 35 59 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=1.705
+ $Y2=0
r100 35 38 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=1.2
+ $Y2=0
r101 33 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r102 33 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r103 33 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r104 29 31 18.4391 $w=2.98e-07 $l=4.8e-07 $layer=LI1_cond $X=3.645 $Y=0.38
+ $X2=3.645 $Y2=0.86
r105 27 65 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=0.085
+ $X2=3.645 $Y2=0
r106 27 29 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=3.645 $Y=0.085
+ $X2=3.645 $Y2=0.38
r107 23 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0
r108 23 25 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0.445
r109 19 59 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.085
+ $X2=1.705 $Y2=0
r110 19 21 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=1.705 $Y=0.085
+ $X2=1.705 $Y2=0.44
r111 15 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r112 15 17 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.43
r113 4 31 182 $w=1.7e-07 $l=7.58288e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.235 $X2=3.63 $Y2=0.86
r114 4 29 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.235 $X2=3.595 $Y2=0.38
r115 3 25 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.235 $X2=2.595 $Y2=0.445
r116 2 21 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.235 $X2=1.715 $Y2=0.44
r117 1 17 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.235 $X2=0.765 $Y2=0.43
.ends

