* File: sky130_fd_sc_lp__dfbbn_2.spice
* Created: Wed Sep  2 09:43:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfbbn_2.pex.spice"
.subckt sky130_fd_sc_lp__dfbbn_2  VNB VPB CLK_N D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK_N	CLK_N
* VPB	VPB
* VNB	VNB
MM1025 N_A_113_57#_M1025_d N_CLK_N_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_113_57#_M1002_g N_A_223_119#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.16275 AS=0.1176 PD=1.195 PS=1.4 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_463_449#_M1012_d N_D_M1012_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.16275 PD=0.7 PS=1.195 NRD=0 NRS=118.56 M=1 R=2.8 SA=75001.1
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_549_449#_M1013_d N_A_223_119#_M1013_g N_A_463_449#_M1012_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.110625 AS=0.0588 PD=0.97 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1041 A_705_104# N_A_113_57#_M1041_g N_A_549_449#_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.110625 PD=0.84 PS=0.97 NRD=44.28 NRS=32.856 M=1 R=2.8
+ SA=75001.9 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_A_789_78#_M1037_g A_705_104# VNB NSHORT L=0.15 W=0.42
+ AD=0.202947 AS=0.0882 PD=1.17679 PS=0.84 NRD=39.996 NRS=44.28 M=1 R=2.8
+ SA=75002.4 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1017 N_A_1018_60#_M1017_d N_SET_B_M1017_g N_VGND_M1037_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0912 AS=0.309253 PD=0.925 PS=1.79321 NRD=0 NRS=80.616 M=1
+ R=4.26667 SA=75002.5 SB=75001 A=0.096 P=1.58 MULT=1
MM1010 N_A_789_78#_M1010_d N_A_549_449#_M1010_g N_A_1018_60#_M1017_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1845 AS=0.0912 PD=1.405 PS=0.925 NRD=43.74 NRS=0.936 M=1
+ R=4.26667 SA=75002.9 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1003 N_A_1018_60#_M1003_d N_A_1191_21#_M1003_g N_A_789_78#_M1010_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1845 PD=1.85 PS=1.405 NRD=0 NRS=14.052 M=1
+ R=4.26667 SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1043 A_1447_119# N_A_789_78#_M1043_g N_VGND_M1043_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1152 AS=0.1824 PD=1 PS=1.85 NRD=23.436 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1019 N_A_1542_428#_M1019_d N_A_113_57#_M1019_g A_1447_119# VNB NSHORT L=0.15
+ W=0.64 AD=0.219955 AS=0.1152 PD=1.49132 PS=1 NRD=44.052 NRS=23.436 M=1
+ R=4.26667 SA=75000.7 SB=75002 A=0.096 P=1.58 MULT=1
MM1015 A_1698_163# N_A_223_119#_M1015_g N_A_1542_428#_M1019_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.144345 PD=0.66 PS=0.978679 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.5 SB=75002 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_1746_137#_M1000_g A_1698_163# VNB NSHORT L=0.15 W=0.42
+ AD=0.117877 AS=0.0504 PD=0.923208 PS=0.66 NRD=52.848 NRS=18.564 M=1 R=2.8
+ SA=75001.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1031 N_A_1911_119#_M1031_d N_SET_B_M1031_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0944 AS=0.179623 PD=0.935 PS=1.40679 NRD=2.808 NRS=12.18 M=1
+ R=4.26667 SA=75001.8 SB=75001 A=0.096 P=1.58 MULT=1
MM1004 N_A_1746_137#_M1004_d N_A_1542_428#_M1004_g N_A_1911_119#_M1031_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.177775 AS=0.0944 PD=1.335 PS=0.935 NRD=14.988 NRS=0
+ M=1 R=4.26667 SA=75002.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1038 N_A_1911_119#_M1038_d N_A_1191_21#_M1038_g N_A_1746_137#_M1004_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1888 AS=0.177775 PD=1.87 PS=1.335 NRD=1.872
+ NRS=14.988 M=1 R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_RESET_B_M1001_g N_A_1191_21#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_Q_N_M1008_d N_A_1746_137#_M1008_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1806 PD=1.12 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1028 N_Q_N_M1008_d N_A_1746_137#_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1032 N_VGND_M1032_d N_A_1746_137#_M1032_g N_A_2618_131#_M1032_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1018 N_Q_M1018_d N_A_2618_131#_M1018_g N_VGND_M1032_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1806 PD=1.12 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1033 N_Q_M1018_d N_A_2618_131#_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2352 PD=1.12 PS=2.24 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1034 N_A_113_57#_M1034_d N_CLK_N_M1034_g N_VPWR_M1034_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.2336 PD=1.85 PS=2.01 NRD=0 NRS=24.6053 M=1 R=4.26667
+ SA=75000.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1035 N_VPWR_M1035_d N_A_113_57#_M1035_g N_A_223_119#_M1035_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.175275 AS=0.1824 PD=1.3766 PS=1.85 NRD=24.6053 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75004.8 A=0.096 P=1.58 MULT=1
MM1042 N_A_463_449#_M1042_d N_D_M1042_g N_VPWR_M1035_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.115025 PD=0.7 PS=0.903396 NRD=0 NRS=66.8224 M=1 R=2.8
+ SA=75000.9 SB=75006.5 A=0.063 P=1.14 MULT=1
MM1023 N_A_549_449#_M1023_d N_A_113_57#_M1023_g N_A_463_449#_M1042_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1365 AS=0.0588 PD=1.07 PS=0.7 NRD=173.537 NRS=0 M=1 R=2.8
+ SA=75001.3 SB=75006.1 A=0.063 P=1.14 MULT=1
MM1030 A_709_449# N_A_223_119#_M1030_g N_A_549_449#_M1023_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.084 AS=0.1365 PD=0.82 PS=1.07 NRD=68.0044 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75005.3 A=0.063 P=1.14 MULT=1
MM1039 N_VPWR_M1039_d N_A_789_78#_M1039_g A_709_449# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.202617 AS=0.084 PD=1.33 PS=0.82 NRD=200.467 NRS=68.0044 M=1 R=2.8
+ SA=75002.6 SB=75004.8 A=0.063 P=1.14 MULT=1
MM1024 N_A_789_78#_M1024_d N_SET_B_M1024_g N_VPWR_M1039_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1176 AS=0.405233 PD=1.12 PS=2.66 NRD=0 NRS=100.234 M=1 R=5.6
+ SA=75002 SB=75003.3 A=0.126 P=1.98 MULT=1
MM1040 A_1119_379# N_A_549_449#_M1040_g N_A_789_78#_M1024_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=29.3136 NRS=0 M=1 R=5.6
+ SA=75002.4 SB=75002.9 A=0.126 P=1.98 MULT=1
MM1036 N_VPWR_M1036_d N_A_1191_21#_M1036_g A_1119_379# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.4116 AS=0.1512 PD=1.82 PS=1.2 NRD=36.3465 NRS=29.3136 M=1 R=5.6
+ SA=75002.9 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1005 A_1447_379# N_A_789_78#_M1005_g N_VPWR_M1036_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.157937 AS=0.4116 PD=1.41 PS=1.82 NRD=31.1851 NRS=127.814 M=1 R=5.6
+ SA=75004.1 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1020 N_A_1542_428#_M1020_d N_A_223_119#_M1020_g A_1447_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1799 AS=0.157937 PD=1.6 PS=1.41 NRD=0 NRS=31.1851 M=1 R=5.6
+ SA=75003.8 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1016 A_1644_506# N_A_113_57#_M1016_g N_A_1542_428#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.14595 AS=0.08995 PD=1.115 PS=0.8 NRD=137.191 NRS=74.6433 M=1 R=2.8
+ SA=75003.1 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_1746_137#_M1021_g A_1644_506# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1232 AS=0.14595 PD=0.956667 PS=1.115 NRD=147.73 NRS=137.191 M=1
+ R=2.8 SA=75003.9 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1014 N_A_1746_137#_M1014_d N_SET_B_M1014_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1176 AS=0.2464 PD=1.12 PS=1.91333 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1022 A_2048_428# N_A_1542_428#_M1022_g N_A_1746_137#_M1014_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.0882 AS=0.1176 PD=1.05 PS=1.12 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75002.9 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_A_1191_21#_M1009_g A_2048_428# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1026 N_VPWR_M1026_d N_RESET_B_M1026_g N_A_1191_21#_M1026_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.137128 AS=0.1792 PD=1.09137 PS=1.84 NRD=49.0136 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1026_d N_A_1746_137#_M1011_g N_Q_N_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.269972 AS=0.1764 PD=2.14863 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1029 N_VPWR_M1029_d N_A_1746_137#_M1029_g N_Q_N_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3717 AS=0.1764 PD=3.11 PS=1.54 NRD=1.5563 NRS=0 M=1 R=8.4
+ SA=75000.9 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_1746_137#_M1006_g N_A_2618_131#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.137128 AS=0.1824 PD=1.09137 PS=1.85 NRD=25.3933 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1007 N_Q_M1007_d N_A_2618_131#_M1007_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.269972 PD=1.54 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_Q_M1007_d N_A_2618_131#_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3528 PD=1.54 PS=3.08 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX44_noxref VNB VPB NWDIODE A=28.713 P=34.5
c_160 VNB 0 3.81024e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dfbbn_2.pxi.spice"
*
.ends
*
*
