# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__o221ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o221ai_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.420000 3.270000 1.755000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 1.310000 2.280000 1.760000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.210000 1.290000 1.410000 ;
        RECT 1.105000 1.410000 1.290000 1.760000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 1.930000 3.275000 2.140000 ;
        RECT 2.955000 2.140000 3.275000 2.945000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.920000 0.585000 2.150000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.280000 0.365000 1.580000 ;
        RECT 0.095000 1.580000 0.935000 1.750000 ;
        RECT 0.185000 2.320000 1.795000 2.490000 ;
        RECT 0.185000 2.490000 0.445000 3.000000 ;
        RECT 0.765000 1.750000 0.935000 2.320000 ;
        RECT 1.465000 2.490000 1.795000 2.990000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.360000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 3.550000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.545000  0.280000 0.835000 0.615000 ;
      RECT 0.545000  0.615000 0.715000 0.870000 ;
      RECT 0.545000  0.870000 1.635000 0.875000 ;
      RECT 0.545000  0.875000 3.075000 1.040000 ;
      RECT 0.615000  2.660000 0.945000 3.245000 ;
      RECT 1.005000  0.280000 1.285000 0.530000 ;
      RECT 1.005000  0.530000 2.600000 0.700000 ;
      RECT 1.465000  0.085000 2.135000 0.360000 ;
      RECT 1.465000  1.040000 3.075000 1.045000 ;
      RECT 2.315000  0.280000 2.600000 0.530000 ;
      RECT 2.365000  2.330000 2.695000 3.245000 ;
      RECT 2.770000  0.280000 3.075000 0.875000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__o221ai_0
END LIBRARY
