* File: sky130_fd_sc_lp__sleep_pargate_plv_14.pxi.spice
* Created: Wed Sep  2 10:37:33 2020
* 
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_14%SLEEP N_SLEEP_c_32_n N_SLEEP_M1000_g
+ N_SLEEP_c_33_n N_SLEEP_M1001_g N_SLEEP_c_34_n SLEEP SLEEP SLEEP SLEEP SLEEP
+ N_SLEEP_c_36_n N_SLEEP_c_37_n PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_14%SLEEP
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_14%VIRTPWR N_VIRTPWR_M1000_d
+ N_VIRTPWR_M1001_d N_VIRTPWR_c_74_n N_VIRTPWR_c_75_n VIRTPWR N_VIRTPWR_c_76_n
+ N_VIRTPWR_c_77_n N_VIRTPWR_c_78_n N_VIRTPWR_c_79_n N_VIRTPWR_c_80_n
+ N_VIRTPWR_c_81_n N_VIRTPWR_c_82_n N_VIRTPWR_c_69_n N_VIRTPWR_c_84_n
+ N_VIRTPWR_c_70_n N_VIRTPWR_c_71_n N_VIRTPWR_c_72_n VIRTPWR N_VIRTPWR_c_73_n
+ PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_14%VIRTPWR
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_14%VPWR N_VPWR_M1000_s VPWR
+ N_VPWR_c_157_n N_VPWR_c_158_n N_VPWR_c_191_n N_VPWR_c_196_n N_VPWR_c_201_n
+ N_VPWR_c_166_n N_VPWR_c_156_n PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_14%VPWR
cc_1 noxref_1 SLEEP 0.0599664f $X=-0.19 $Y=-0.007 $X2=8.315 $Y2=0.84
cc_2 noxref_1 VIRTPWR 0.105802f $X=-0.19 $Y=-0.007 $X2=8.315 $Y2=1.21
cc_3 noxref_1 N_VIRTPWR_c_69_n 0.0836651f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_4 noxref_1 N_VIRTPWR_c_70_n 0.0786895f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_5 noxref_1 N_VIRTPWR_c_71_n 0.0386646f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_6 noxref_1 N_VIRTPWR_c_72_n 0.0386646f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_7 noxref_1 N_VIRTPWR_c_73_n 0.0386646f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_8 noxref_1 N_VPWR_c_156_n 0.672577f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_9 VPB N_SLEEP_c_32_n 0.0222395f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=2.325
cc_10 VPB N_SLEEP_c_33_n 0.045835f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=2.755
cc_11 VPB N_SLEEP_c_34_n 0.0108874f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=2.325
cc_12 VPB SLEEP 0.030975f $X=-0.19 $Y=1.655 $X2=8.315 $Y2=0.84
cc_13 VPB N_SLEEP_c_36_n 0.0602836f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=1.985
cc_14 VPB N_SLEEP_c_37_n 0.0240095f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=2.665
cc_15 VPB N_VIRTPWR_c_74_n 0.0130323f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=2.25
cc_16 VPB N_VIRTPWR_c_75_n 0.0357155f $X=-0.19 $Y=1.655 $X2=8.315 $Y2=0.84
cc_17 VPB N_VIRTPWR_c_76_n 0.15875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_18 VPB N_VIRTPWR_c_77_n 0.00830421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_19 VPB N_VIRTPWR_c_78_n 0.00830421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_20 VPB N_VIRTPWR_c_79_n 0.00830421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_21 VPB N_VIRTPWR_c_80_n 0.00855727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_VIRTPWR_c_81_n 0.121651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_23 VPB N_VIRTPWR_c_82_n 0.0329627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_24 VPB N_VIRTPWR_c_69_n 0.0405705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 VPB N_VIRTPWR_c_84_n 0.0130323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_VIRTPWR_c_70_n 0.0404102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_157_n 0.00214921f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=1.985
cc_28 VPB N_VPWR_c_158_n 0.00210523f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=2.665
cc_29 VPB N_VPWR_c_156_n 0.124448f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 N_SLEEP_c_33_n N_VIRTPWR_c_74_n 0.0158929f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_31 N_SLEEP_c_33_n N_VIRTPWR_c_75_n 0.00259154f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_32 N_SLEEP_c_32_n N_VIRTPWR_c_77_n 0.00539584f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_33 N_SLEEP_c_33_n N_VIRTPWR_c_77_n 0.00539584f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_34 N_SLEEP_c_32_n N_VIRTPWR_c_78_n 0.00539584f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_35 N_SLEEP_c_33_n N_VIRTPWR_c_78_n 0.00539584f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_36 N_SLEEP_c_32_n N_VIRTPWR_c_79_n 0.00539584f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_37 N_SLEEP_c_33_n N_VIRTPWR_c_79_n 0.00539584f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_38 N_SLEEP_c_32_n N_VIRTPWR_c_80_n 0.00539734f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_39 N_SLEEP_c_33_n N_VIRTPWR_c_80_n 0.00539734f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_40 N_SLEEP_c_32_n N_VIRTPWR_c_81_n 0.0119829f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_41 SLEEP N_VIRTPWR_c_81_n 0.0112305f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_42 N_SLEEP_c_36_n N_VIRTPWR_c_81_n 0.00525497f $X=8.42 $Y=1.985 $X2=0 $Y2=0
cc_43 N_SLEEP_c_33_n N_VIRTPWR_c_82_n 0.00576677f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_44 SLEEP N_VIRTPWR_c_82_n 0.0165417f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_45 N_SLEEP_c_33_n N_VIRTPWR_c_69_n 0.0037323f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_46 SLEEP N_VIRTPWR_c_69_n 0.0123629f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_47 N_SLEEP_c_33_n N_VIRTPWR_c_70_n 0.00224979f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_48 N_SLEEP_c_32_n N_VPWR_c_157_n 0.010275f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_49 N_SLEEP_c_33_n N_VPWR_c_157_n 0.010275f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_50 SLEEP N_VPWR_c_157_n 0.0107074f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_51 N_SLEEP_c_37_n N_VPWR_c_157_n 0.00207026f $X=8.42 $Y=2.665 $X2=0 $Y2=0
cc_52 N_SLEEP_c_32_n N_VPWR_c_158_n 0.00731714f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_53 N_SLEEP_c_33_n N_VPWR_c_158_n 0.00246406f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_54 SLEEP N_VPWR_c_166_n 0.0033926f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_55 N_SLEEP_c_32_n N_VPWR_c_156_n 0.00722775f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_56 N_SLEEP_c_33_n N_VPWR_c_156_n 0.00984441f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_57 SLEEP N_VPWR_c_156_n 0.106016f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_58 N_SLEEP_c_36_n N_VPWR_c_156_n 0.00617994f $X=8.42 $Y=1.985 $X2=0 $Y2=0
cc_59 N_SLEEP_c_37_n N_VPWR_c_156_n 0.00118998f $X=8.42 $Y=2.665 $X2=0 $Y2=0
cc_60 N_VIRTPWR_c_77_n N_VPWR_M1000_s 4.84807e-19 $X=2.34 $Y=2.11 $X2=-0.19
+ $Y2=-0.007
cc_61 N_VIRTPWR_c_78_n N_VPWR_M1000_s 4.84807e-19 $X=3.895 $Y=2.11 $X2=-0.19
+ $Y2=-0.007
cc_62 N_VIRTPWR_c_79_n N_VPWR_M1000_s 4.84807e-19 $X=5.45 $Y=2.11 $X2=-0.19
+ $Y2=-0.007
cc_63 N_VIRTPWR_c_80_n N_VPWR_M1000_s 4.85041e-19 $X=7.005 $Y=2.11 $X2=-0.19
+ $Y2=-0.007
cc_64 N_VIRTPWR_c_74_n N_VPWR_c_157_n 0.262559f $X=1.342 $Y=3.127 $X2=0 $Y2=0
cc_65 N_VIRTPWR_c_77_n N_VPWR_c_157_n 0.0346616f $X=2.34 $Y=2.11 $X2=0 $Y2=0
cc_66 N_VIRTPWR_c_78_n N_VPWR_c_157_n 0.0346616f $X=3.895 $Y=2.11 $X2=0 $Y2=0
cc_67 N_VIRTPWR_c_79_n N_VPWR_c_157_n 0.0346616f $X=5.45 $Y=2.11 $X2=0 $Y2=0
cc_68 N_VIRTPWR_c_80_n N_VPWR_c_157_n 0.0356496f $X=7.005 $Y=2.11 $X2=0 $Y2=0
cc_69 N_VIRTPWR_c_81_n N_VPWR_c_157_n 0.258116f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_70 N_VIRTPWR_c_69_n N_VPWR_c_157_n 0.00290716f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_71 N_VIRTPWR_c_70_n N_VPWR_c_157_n 0.00285709f $X=1.845 $Y=3.33 $X2=0 $Y2=0
cc_72 N_VIRTPWR_c_71_n N_VPWR_c_157_n 0.0012824f $X=3.4 $Y=3.33 $X2=0 $Y2=0
cc_73 N_VIRTPWR_c_72_n N_VPWR_c_157_n 0.0012824f $X=4.955 $Y=3.33 $X2=0 $Y2=0
cc_74 N_VIRTPWR_c_73_n N_VPWR_c_157_n 0.0012824f $X=6.51 $Y=3.33 $X2=0 $Y2=0
cc_75 N_VIRTPWR_c_74_n N_VPWR_c_158_n 0.00538617f $X=1.342 $Y=3.127 $X2=0 $Y2=0
cc_76 N_VIRTPWR_c_77_n N_VPWR_c_158_n 0.0219135f $X=2.34 $Y=2.11 $X2=0 $Y2=0
cc_77 N_VIRTPWR_c_81_n N_VPWR_c_158_n 0.0145601f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_78 N_VIRTPWR_c_70_n N_VPWR_c_158_n 0.0256157f $X=1.845 $Y=3.33 $X2=0 $Y2=0
cc_79 N_VIRTPWR_c_76_n N_VPWR_c_191_n 0.0065368f $X=7.768 $Y=3.127 $X2=0 $Y2=0
cc_80 N_VIRTPWR_c_77_n N_VPWR_c_191_n 0.0219135f $X=2.34 $Y=2.11 $X2=0 $Y2=0
cc_81 N_VIRTPWR_c_78_n N_VPWR_c_191_n 0.0219135f $X=3.895 $Y=2.11 $X2=0 $Y2=0
cc_82 N_VIRTPWR_c_81_n N_VPWR_c_191_n 0.0145601f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_83 N_VIRTPWR_c_71_n N_VPWR_c_191_n 0.0224574f $X=3.4 $Y=3.33 $X2=0 $Y2=0
cc_84 N_VIRTPWR_c_76_n N_VPWR_c_196_n 0.0065368f $X=7.768 $Y=3.127 $X2=0 $Y2=0
cc_85 N_VIRTPWR_c_78_n N_VPWR_c_196_n 0.0219135f $X=3.895 $Y=2.11 $X2=0 $Y2=0
cc_86 N_VIRTPWR_c_79_n N_VPWR_c_196_n 0.0219135f $X=5.45 $Y=2.11 $X2=0 $Y2=0
cc_87 N_VIRTPWR_c_81_n N_VPWR_c_196_n 0.0145601f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_88 N_VIRTPWR_c_72_n N_VPWR_c_196_n 0.0224574f $X=4.955 $Y=3.33 $X2=0 $Y2=0
cc_89 N_VIRTPWR_c_76_n N_VPWR_c_201_n 0.0065368f $X=7.768 $Y=3.127 $X2=0 $Y2=0
cc_90 N_VIRTPWR_c_79_n N_VPWR_c_201_n 0.0219135f $X=5.45 $Y=2.11 $X2=0 $Y2=0
cc_91 N_VIRTPWR_c_80_n N_VPWR_c_201_n 0.0219152f $X=7.005 $Y=2.11 $X2=0 $Y2=0
cc_92 N_VIRTPWR_c_81_n N_VPWR_c_201_n 0.0145601f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_93 N_VIRTPWR_c_73_n N_VPWR_c_201_n 0.0224574f $X=6.51 $Y=3.33 $X2=0 $Y2=0
cc_94 N_VIRTPWR_c_76_n N_VPWR_c_166_n 0.00538617f $X=7.768 $Y=3.127 $X2=0 $Y2=0
cc_95 N_VIRTPWR_c_80_n N_VPWR_c_166_n 0.0219152f $X=7.005 $Y=2.11 $X2=0 $Y2=0
cc_96 N_VIRTPWR_c_81_n N_VPWR_c_166_n 0.0145601f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_97 N_VIRTPWR_c_69_n N_VPWR_c_166_n 0.0256157f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_98 N_VIRTPWR_c_74_n N_VPWR_c_156_n 0.00611837f $X=1.342 $Y=3.127 $X2=0 $Y2=0
cc_99 VIRTPWR N_VPWR_c_156_n 0.224849f $X=0 $Y=3.085 $X2=0 $Y2=0
cc_100 N_VIRTPWR_c_76_n N_VPWR_c_156_n 0.0186573f $X=7.768 $Y=3.127 $X2=0 $Y2=0
cc_101 N_VIRTPWR_c_77_n N_VPWR_c_156_n 0.198826f $X=2.34 $Y=2.11 $X2=0 $Y2=0
cc_102 N_VIRTPWR_c_78_n N_VPWR_c_156_n 0.198826f $X=3.895 $Y=2.11 $X2=0 $Y2=0
cc_103 N_VIRTPWR_c_79_n N_VPWR_c_156_n 0.198826f $X=5.45 $Y=2.11 $X2=0 $Y2=0
cc_104 N_VIRTPWR_c_80_n N_VPWR_c_156_n 0.203254f $X=7.005 $Y=2.11 $X2=0 $Y2=0
cc_105 N_VIRTPWR_c_81_n N_VPWR_c_156_n 0.119244f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_106 N_VIRTPWR_c_69_n N_VPWR_c_156_n 0.227442f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_107 N_VIRTPWR_c_84_n N_VPWR_c_156_n 0.00787277f $X=8.055 $Y=3.127 $X2=0 $Y2=0
cc_108 N_VIRTPWR_c_70_n N_VPWR_c_156_n 0.212348f $X=1.845 $Y=3.33 $X2=0 $Y2=0
cc_109 N_VIRTPWR_c_71_n N_VPWR_c_156_n 0.0980574f $X=3.4 $Y=3.33 $X2=0 $Y2=0
cc_110 N_VIRTPWR_c_72_n N_VPWR_c_156_n 0.0980574f $X=4.955 $Y=3.33 $X2=0 $Y2=0
cc_111 N_VIRTPWR_c_73_n N_VPWR_c_156_n 0.0980574f $X=6.51 $Y=3.33 $X2=0 $Y2=0
