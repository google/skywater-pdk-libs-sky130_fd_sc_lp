* File: sky130_fd_sc_lp__a31oi_0.spice
* Created: Wed Sep  2 09:26:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a31oi_0.pex.spice"
.subckt sky130_fd_sc_lp__a31oi_0  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1002 A_123_47# N_A3_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1113 PD=0.66 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1007 A_201_47# N_A2_M1007_g A_123_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g A_201_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=21.42 NRS=18.564 M=1 R=2.8 SA=75001 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0882 PD=1.37 PS=0.84 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_110_473#_M1005_d N_A3_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_110_473#_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_A_110_473#_M1006_d N_A1_M1006_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_110_473#_M1006_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
c_54 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a31oi_0.pxi.spice"
*
.ends
*
*
