# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux2_lp2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__mux2_lp2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.810000 2.315000 1.145000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.515000 2.665000 1.845000 ;
        RECT 2.495000 0.905000 3.235000 1.235000 ;
        RECT 2.495000 1.235000 2.665000 1.515000 ;
        RECT 3.005000 0.440000 3.235000 0.905000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.845000 1.475000 4.195000 1.805000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.265000 0.450000 2.520000 ;
        RECT 0.115000 2.520000 0.445000 3.025000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.630000  0.905000 1.590000 1.235000 ;
      RECT 0.645000  2.765000 0.975000 3.245000 ;
      RECT 0.910000  0.085000 1.240000 0.725000 ;
      RECT 0.910000  1.515000 1.240000 2.415000 ;
      RECT 0.910000  2.415000 3.915000 2.585000 ;
      RECT 1.420000  0.345000 2.825000 0.515000 ;
      RECT 1.420000  0.515000 1.590000 0.905000 ;
      RECT 1.420000  1.235000 1.590000 2.065000 ;
      RECT 1.420000  2.065000 2.325000 2.235000 ;
      RECT 2.495000  0.515000 2.825000 0.725000 ;
      RECT 3.055000  2.765000 3.385000 3.245000 ;
      RECT 3.425000  0.085000 3.755000 0.725000 ;
      RECT 3.585000  1.985000 4.545000 2.155000 ;
      RECT 3.585000  2.155000 3.915000 2.415000 ;
      RECT 3.585000  2.585000 3.915000 3.025000 ;
      RECT 4.215000  0.265000 4.545000 0.725000 ;
      RECT 4.375000  0.725000 4.545000 1.985000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__mux2_lp2
END LIBRARY
