* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
X0 VGND CI a_239_135# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_878_41# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_239_135# a_814_384# a_84_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_84_21# a_1022_362# a_630_100# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_84_21# a_1022_362# a_239_135# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 a_814_384# B a_1930_367# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 COUT a_413_34# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_1930_367# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_630_100# a_814_384# a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_1022_362# B a_1741_367# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 VGND A a_2229_269# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_413_34# a_1022_362# a_239_135# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_413_34# a_1022_362# a_878_41# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_1930_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_1022_362# B a_1930_367# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_878_41# a_814_384# a_413_34# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VPWR a_239_135# a_630_100# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_814_384# B a_1741_367# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 SUM a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_1741_367# a_2229_269# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 a_239_135# a_814_384# a_413_34# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_1741_367# a_878_41# a_1022_362# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 VPWR A a_2229_269# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VPWR CI a_239_135# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_1930_367# a_878_41# a_814_384# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_1741_367# a_2229_269# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 SUM a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 COUT a_413_34# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_1741_367# a_878_41# a_814_384# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X29 VGND a_239_135# a_630_100# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 a_1930_367# a_878_41# a_1022_362# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X31 a_878_41# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
