# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o21ba_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o21ba_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.015000 1.415000 4.345000 1.675000 ;
        RECT 4.075000 1.675000 4.345000 2.310000 ;
        RECT 4.075000 2.310000 5.605000 2.500000 ;
        RECT 5.435000 1.415000 5.860000 1.645000 ;
        RECT 5.435000 1.645000 5.605000 2.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.920000 1.415000 5.250000 1.760000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.200000 0.865000 1.750000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.920000 1.205000 1.930000 ;
        RECT 0.625000 1.930000 2.255000 2.260000 ;
        RECT 1.035000 0.255000 1.285000 1.075000 ;
        RECT 1.035000 1.075000 2.145000 1.245000 ;
        RECT 1.035000 1.245000 1.205000 1.920000 ;
        RECT 1.955000 0.255000 2.145000 1.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.085000  0.255000 0.425000 1.030000 ;
      RECT 0.085000  1.030000 0.260000 1.920000 ;
      RECT 0.085000  1.920000 0.455000 2.430000 ;
      RECT 0.085000  2.430000 2.595000 2.610000 ;
      RECT 0.085000  2.610000 0.465000 3.075000 ;
      RECT 0.595000  0.085000 0.865000 1.030000 ;
      RECT 0.635000  2.780000 0.965000 3.245000 ;
      RECT 1.375000  1.415000 2.485000 1.605000 ;
      RECT 1.455000  0.085000 1.785000 0.905000 ;
      RECT 1.495000  2.780000 1.825000 3.245000 ;
      RECT 2.315000  0.085000 2.645000 0.905000 ;
      RECT 2.315000  1.075000 4.695000 1.245000 ;
      RECT 2.315000  1.245000 2.485000 1.415000 ;
      RECT 2.360000  2.780000 3.035000 3.245000 ;
      RECT 2.425000  1.775000 3.010000 1.945000 ;
      RECT 2.425000  1.945000 2.595000 2.430000 ;
      RECT 2.680000  1.415000 3.010000 1.775000 ;
      RECT 2.765000  2.115000 3.035000 2.780000 ;
      RECT 2.835000  0.265000 4.185000 0.435000 ;
      RECT 2.835000  0.435000 3.175000 0.905000 ;
      RECT 3.205000  1.245000 3.425000 3.075000 ;
      RECT 3.345000  0.605000 3.675000 1.075000 ;
      RECT 3.595000  1.815000 3.905000 2.785000 ;
      RECT 3.595000  2.785000 4.265000 3.245000 ;
      RECT 3.855000  0.435000 4.185000 0.725000 ;
      RECT 3.855000  0.725000 5.055000 0.895000 ;
      RECT 4.355000  0.085000 4.695000 0.555000 ;
      RECT 4.435000  2.670000 5.495000 3.000000 ;
      RECT 4.525000  1.245000 4.695000 1.930000 ;
      RECT 4.525000  1.930000 5.125000 2.140000 ;
      RECT 4.865000  0.295000 5.055000 0.725000 ;
      RECT 4.865000  0.895000 5.055000 1.075000 ;
      RECT 4.865000  1.075000 6.005000 1.245000 ;
      RECT 5.225000  0.085000 5.555000 0.905000 ;
      RECT 5.735000  0.305000 6.005000 1.075000 ;
      RECT 5.775000  1.815000 6.025000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__o21ba_4
END LIBRARY
